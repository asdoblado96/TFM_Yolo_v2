LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_8_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_8_WROM;

ARCHITECTURE RTL OF L8_8_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"001100001",
  1=>"011110101",
  2=>"111011001",
  3=>"111011010",
  4=>"010000101",
  5=>"000110010",
  6=>"000011101",
  7=>"111100001",
  8=>"110110110",
  9=>"000000001",
  10=>"010001000",
  11=>"101101010",
  12=>"101111100",
  13=>"001110010",
  14=>"000011100",
  15=>"010101110",
  16=>"110110011",
  17=>"101111100",
  18=>"011001111",
  19=>"001110010",
  20=>"000010101",
  21=>"001111110",
  22=>"001000110",
  23=>"001001000",
  24=>"011001000",
  25=>"111101001",
  26=>"100011001",
  27=>"100100000",
  28=>"000100110",
  29=>"000100111",
  30=>"010110001",
  31=>"001001011",
  32=>"111110111",
  33=>"000000001",
  34=>"101001101",
  35=>"111100101",
  36=>"000101011",
  37=>"010110111",
  38=>"011010000",
  39=>"000010110",
  40=>"111101101",
  41=>"100000101",
  42=>"000111011",
  43=>"001001011",
  44=>"101001101",
  45=>"100001101",
  46=>"111010010",
  47=>"111100100",
  48=>"101010100",
  49=>"111100111",
  50=>"011110110",
  51=>"111010001",
  52=>"110001110",
  53=>"011100110",
  54=>"001000000",
  55=>"010010111",
  56=>"111001011",
  57=>"000001011",
  58=>"010001001",
  59=>"000000000",
  60=>"110101111",
  61=>"110100100",
  62=>"101111101",
  63=>"001000011",
  64=>"111011101",
  65=>"000000011",
  66=>"111111011",
  67=>"111100010",
  68=>"110111100",
  69=>"101100110",
  70=>"001100111",
  71=>"101010000",
  72=>"000101000",
  73=>"111100010",
  74=>"000000100",
  75=>"011100111",
  76=>"101111101",
  77=>"011101100",
  78=>"100000111",
  79=>"011111111",
  80=>"111101101",
  81=>"111110111",
  82=>"110010001",
  83=>"100001010",
  84=>"110010001",
  85=>"110111110",
  86=>"111110101",
  87=>"101001000",
  88=>"001000001",
  89=>"001111010",
  90=>"000100101",
  91=>"111010010",
  92=>"000000100",
  93=>"101111011",
  94=>"001010110",
  95=>"010111110",
  96=>"100001110",
  97=>"000110100",
  98=>"010011100",
  99=>"100010010",
  100=>"010110110",
  101=>"100000011",
  102=>"010111010",
  103=>"001000010",
  104=>"011100010",
  105=>"000000111",
  106=>"010010101",
  107=>"001011110",
  108=>"010000101",
  109=>"110110000",
  110=>"100001001",
  111=>"100000010",
  112=>"000010000",
  113=>"101111000",
  114=>"111001110",
  115=>"010101000",
  116=>"010000000",
  117=>"110111000",
  118=>"001001110",
  119=>"011101110",
  120=>"011010111",
  121=>"101001011",
  122=>"000010011",
  123=>"000010001",
  124=>"000101001",
  125=>"111110011",
  126=>"100001110",
  127=>"010010111",
  128=>"011000101",
  129=>"111111101",
  130=>"011000000",
  131=>"011001100",
  132=>"101010101",
  133=>"001011111",
  134=>"010100100",
  135=>"001101011",
  136=>"001000111",
  137=>"100110101",
  138=>"001000000",
  139=>"101101111",
  140=>"111101000",
  141=>"011000010",
  142=>"011011010",
  143=>"011000001",
  144=>"111101101",
  145=>"100000100",
  146=>"110111110",
  147=>"001010010",
  148=>"111111011",
  149=>"010001000",
  150=>"000111110",
  151=>"000111010",
  152=>"000011010",
  153=>"111000111",
  154=>"011111111",
  155=>"010010000",
  156=>"001001011",
  157=>"001110100",
  158=>"011101011",
  159=>"101101110",
  160=>"111100001",
  161=>"010010010",
  162=>"100100000",
  163=>"010001000",
  164=>"110111101",
  165=>"101001000",
  166=>"000111100",
  167=>"001000100",
  168=>"101001110",
  169=>"110001011",
  170=>"011101011",
  171=>"110001011",
  172=>"010110001",
  173=>"011110101",
  174=>"010110011",
  175=>"100101000",
  176=>"111111111",
  177=>"000100010",
  178=>"111011000",
  179=>"110011110",
  180=>"110010000",
  181=>"010001000",
  182=>"010101000",
  183=>"000101001",
  184=>"110100101",
  185=>"100001000",
  186=>"001101011",
  187=>"100100010",
  188=>"011011000",
  189=>"111100000",
  190=>"000000010",
  191=>"000000010",
  192=>"110000001",
  193=>"011011110",
  194=>"100000101",
  195=>"000100111",
  196=>"011100101",
  197=>"101101110",
  198=>"000111001",
  199=>"001011111",
  200=>"100110110",
  201=>"011010110",
  202=>"011000101",
  203=>"111011011",
  204=>"101000011",
  205=>"000101100",
  206=>"110100000",
  207=>"011010110",
  208=>"111001000",
  209=>"010101100",
  210=>"001010011",
  211=>"000010000",
  212=>"010000011",
  213=>"001010011",
  214=>"010000110",
  215=>"111000111",
  216=>"110001110",
  217=>"110000000",
  218=>"101001100",
  219=>"001111100",
  220=>"111011010",
  221=>"101100110",
  222=>"101101110",
  223=>"111111110",
  224=>"000111011",
  225=>"110111111",
  226=>"001011110",
  227=>"101110000",
  228=>"110111000",
  229=>"011000101",
  230=>"010100110",
  231=>"010010110",
  232=>"011100000",
  233=>"101001101",
  234=>"000000100",
  235=>"011001101",
  236=>"010000000",
  237=>"101001000",
  238=>"101110010",
  239=>"111111111",
  240=>"111111011",
  241=>"000110100",
  242=>"000001110",
  243=>"010010101",
  244=>"000000101",
  245=>"101000000",
  246=>"100011010",
  247=>"000001010",
  248=>"101001011",
  249=>"111101010",
  250=>"000111010",
  251=>"001111111",
  252=>"011000101",
  253=>"001011000",
  254=>"111111010",
  255=>"001011111",
  256=>"001010111",
  257=>"001010100",
  258=>"100110111",
  259=>"011100101",
  260=>"111011011",
  261=>"010110101",
  262=>"000000101",
  263=>"010100010",
  264=>"011101001",
  265=>"111100101",
  266=>"001101111",
  267=>"100100101",
  268=>"001111001",
  269=>"110000100",
  270=>"110001111",
  271=>"111000110",
  272=>"100111110",
  273=>"010011111",
  274=>"111000000",
  275=>"100111101",
  276=>"110110011",
  277=>"101111100",
  278=>"101001110",
  279=>"011100101",
  280=>"101100100",
  281=>"011110011",
  282=>"000010010",
  283=>"001010011",
  284=>"101100011",
  285=>"101000111",
  286=>"010000110",
  287=>"111001110",
  288=>"000010111",
  289=>"100100001",
  290=>"101100100",
  291=>"110111110",
  292=>"010111101",
  293=>"110100000",
  294=>"001110011",
  295=>"111110011",
  296=>"100101010",
  297=>"000110000",
  298=>"001000110",
  299=>"100111011",
  300=>"111000011",
  301=>"110101001",
  302=>"111101111",
  303=>"101010011",
  304=>"001010011",
  305=>"000010110",
  306=>"111110110",
  307=>"100010100",
  308=>"000110111",
  309=>"011001110",
  310=>"010101110",
  311=>"000101111",
  312=>"010010001",
  313=>"101100000",
  314=>"001000000",
  315=>"110111111",
  316=>"010100000",
  317=>"001110110",
  318=>"001100011",
  319=>"011111111",
  320=>"011000000",
  321=>"011000001",
  322=>"000010110",
  323=>"110010100",
  324=>"001010111",
  325=>"100111011",
  326=>"111100101",
  327=>"111000100",
  328=>"011111010",
  329=>"010101001",
  330=>"010110100",
  331=>"110010110",
  332=>"111111001",
  333=>"110110011",
  334=>"001001111",
  335=>"100011101",
  336=>"100001100",
  337=>"101000110",
  338=>"001101101",
  339=>"100011100",
  340=>"000111000",
  341=>"111110100",
  342=>"111011010",
  343=>"001010101",
  344=>"100010101",
  345=>"000111110",
  346=>"100001110",
  347=>"110100001",
  348=>"000010001",
  349=>"011011000",
  350=>"110011000",
  351=>"000011010",
  352=>"110110101",
  353=>"010101110",
  354=>"010011111",
  355=>"100010011",
  356=>"100101000",
  357=>"011000111",
  358=>"111001101",
  359=>"110111001",
  360=>"010110100",
  361=>"000111001",
  362=>"010111000",
  363=>"100100101",
  364=>"111001000",
  365=>"001111110",
  366=>"110111010",
  367=>"000001100",
  368=>"110111110",
  369=>"110001001",
  370=>"010110100",
  371=>"111101111",
  372=>"100001000",
  373=>"000111101",
  374=>"011011000",
  375=>"101011111",
  376=>"000100100",
  377=>"110000001",
  378=>"111000111",
  379=>"111111100",
  380=>"001011110",
  381=>"111011010",
  382=>"110011000",
  383=>"100001110",
  384=>"111111101",
  385=>"000011100",
  386=>"001001110",
  387=>"101101011",
  388=>"001101111",
  389=>"000111000",
  390=>"010001011",
  391=>"000101100",
  392=>"001011010",
  393=>"110100010",
  394=>"110100011",
  395=>"110110100",
  396=>"100110110",
  397=>"000100110",
  398=>"010111011",
  399=>"101111011",
  400=>"101011101",
  401=>"100000001",
  402=>"000101010",
  403=>"000110011",
  404=>"000100000",
  405=>"011000110",
  406=>"000010001",
  407=>"001101111",
  408=>"010001101",
  409=>"111001101",
  410=>"101111001",
  411=>"110100111",
  412=>"101101011",
  413=>"100101011",
  414=>"101111011",
  415=>"000001000",
  416=>"001001111",
  417=>"101100110",
  418=>"010111101",
  419=>"001000001",
  420=>"001011011",
  421=>"001100011",
  422=>"000100101",
  423=>"010111001",
  424=>"001010100",
  425=>"011110000",
  426=>"111010000",
  427=>"001010111",
  428=>"100000101",
  429=>"101010101",
  430=>"111100111",
  431=>"101100100",
  432=>"100100010",
  433=>"110001000",
  434=>"111001110",
  435=>"011001100",
  436=>"010011110",
  437=>"000011110",
  438=>"111011110",
  439=>"001100111",
  440=>"101101000",
  441=>"100101101",
  442=>"010111111",
  443=>"011111111",
  444=>"011111111",
  445=>"000000110",
  446=>"100100101",
  447=>"001000101",
  448=>"010000011",
  449=>"001110111",
  450=>"101111010",
  451=>"110010110",
  452=>"001001010",
  453=>"111010011",
  454=>"100000101",
  455=>"111001000",
  456=>"110101100",
  457=>"101001110",
  458=>"000000100",
  459=>"000101110",
  460=>"000111101",
  461=>"000001001",
  462=>"101110100",
  463=>"100101001",
  464=>"111100011",
  465=>"100010010",
  466=>"111111000",
  467=>"011101111",
  468=>"010110100",
  469=>"000011110",
  470=>"101100010",
  471=>"110011000",
  472=>"001001111",
  473=>"011100001",
  474=>"100100001",
  475=>"010110001",
  476=>"111100101",
  477=>"111000000",
  478=>"000000111",
  479=>"110110010",
  480=>"111111111",
  481=>"010101000",
  482=>"010010010",
  483=>"001110101",
  484=>"010010000",
  485=>"001011111",
  486=>"110100000",
  487=>"000000001",
  488=>"111011000",
  489=>"011001110",
  490=>"001101010",
  491=>"101011101",
  492=>"111000001",
  493=>"100000011",
  494=>"100010110",
  495=>"011000010",
  496=>"111010100",
  497=>"100100100",
  498=>"001101010",
  499=>"000111111",
  500=>"101001111",
  501=>"010110111",
  502=>"010110111",
  503=>"001000111",
  504=>"110100111",
  505=>"100011101",
  506=>"011110111",
  507=>"110001101",
  508=>"110111000",
  509=>"001111100",
  510=>"110011110",
  511=>"000000100",
  512=>"010011111",
  513=>"110100111",
  514=>"101010111",
  515=>"000011001",
  516=>"110101100",
  517=>"001111000",
  518=>"110110101",
  519=>"000000110",
  520=>"001001000",
  521=>"011110100",
  522=>"011011100",
  523=>"011000001",
  524=>"110010110",
  525=>"010110001",
  526=>"001001010",
  527=>"111110110",
  528=>"011010011",
  529=>"111101110",
  530=>"010001011",
  531=>"010001001",
  532=>"010010000",
  533=>"001011000",
  534=>"001111011",
  535=>"010000001",
  536=>"110110110",
  537=>"001010010",
  538=>"010100001",
  539=>"010001010",
  540=>"000101000",
  541=>"011111010",
  542=>"101010000",
  543=>"110011111",
  544=>"010000000",
  545=>"101010001",
  546=>"001000011",
  547=>"000111011",
  548=>"001110100",
  549=>"100101111",
  550=>"101001000",
  551=>"100100100",
  552=>"011010011",
  553=>"100111011",
  554=>"010011111",
  555=>"101001111",
  556=>"010110010",
  557=>"101001101",
  558=>"010011010",
  559=>"011111101",
  560=>"011111111",
  561=>"010111000",
  562=>"011111000",
  563=>"011100011",
  564=>"111100100",
  565=>"111111000",
  566=>"100000000",
  567=>"101101010",
  568=>"100011111",
  569=>"111101010",
  570=>"000011000",
  571=>"111010111",
  572=>"000100110",
  573=>"010101011",
  574=>"111011000",
  575=>"000111001",
  576=>"011110000",
  577=>"011111100",
  578=>"001101100",
  579=>"000110111",
  580=>"000101011",
  581=>"111101010",
  582=>"101111000",
  583=>"100001111",
  584=>"001011101",
  585=>"110111011",
  586=>"000110101",
  587=>"011001001",
  588=>"011000111",
  589=>"110111110",
  590=>"001110010",
  591=>"011011110",
  592=>"010011101",
  593=>"000111000",
  594=>"100010111",
  595=>"010110111",
  596=>"000111000",
  597=>"100001001",
  598=>"010000010",
  599=>"001000001",
  600=>"100111101",
  601=>"101010001",
  602=>"101101000",
  603=>"000000000",
  604=>"010110101",
  605=>"001000111",
  606=>"010101111",
  607=>"101011011",
  608=>"101110010",
  609=>"100000100",
  610=>"000000001",
  611=>"011111000",
  612=>"111011101",
  613=>"110001101",
  614=>"000001010",
  615=>"101001001",
  616=>"110011011",
  617=>"010001111",
  618=>"011110100",
  619=>"010000000",
  620=>"100111100",
  621=>"011001001",
  622=>"010001101",
  623=>"001101111",
  624=>"111101011",
  625=>"111111101",
  626=>"111100110",
  627=>"101011100",
  628=>"111000110",
  629=>"110110100",
  630=>"100111101",
  631=>"011101000",
  632=>"101101011",
  633=>"101010110",
  634=>"000111100",
  635=>"110001101",
  636=>"111100111",
  637=>"101101101",
  638=>"100111011",
  639=>"011010101",
  640=>"110110001",
  641=>"000011110",
  642=>"100100000",
  643=>"101101110",
  644=>"000011010",
  645=>"100011010",
  646=>"101101010",
  647=>"111110010",
  648=>"100011110",
  649=>"000010101",
  650=>"111101110",
  651=>"010010111",
  652=>"011100110",
  653=>"111001011",
  654=>"000110001",
  655=>"001010001",
  656=>"010000011",
  657=>"110111010",
  658=>"111010011",
  659=>"011101010",
  660=>"011011111",
  661=>"011100000",
  662=>"111111110",
  663=>"001101110",
  664=>"011110000",
  665=>"000011001",
  666=>"011001110",
  667=>"001110000",
  668=>"101001001",
  669=>"010010110",
  670=>"000010000",
  671=>"110100001",
  672=>"010011110",
  673=>"111110000",
  674=>"010000111",
  675=>"000111101",
  676=>"111100000",
  677=>"100011000",
  678=>"011100100",
  679=>"000010110",
  680=>"101010001",
  681=>"011011010",
  682=>"011111111",
  683=>"010110010",
  684=>"001000000",
  685=>"000000111",
  686=>"111010100",
  687=>"111001110",
  688=>"011110100",
  689=>"111111011",
  690=>"111100100",
  691=>"001000110",
  692=>"100000111",
  693=>"111101100",
  694=>"101011001",
  695=>"110111000",
  696=>"011001100",
  697=>"110101011",
  698=>"101101111",
  699=>"100100111",
  700=>"101000001",
  701=>"000101011",
  702=>"111011100",
  703=>"000011001",
  704=>"110010000",
  705=>"111010101",
  706=>"101011011",
  707=>"011000111",
  708=>"010010000",
  709=>"100011010",
  710=>"101001001",
  711=>"011000101",
  712=>"111100001",
  713=>"101001010",
  714=>"111100010",
  715=>"111110101",
  716=>"111010100",
  717=>"100110010",
  718=>"010101011",
  719=>"000110101",
  720=>"011111101",
  721=>"100000100",
  722=>"000110010",
  723=>"000110101",
  724=>"100100001",
  725=>"001010010",
  726=>"111001010",
  727=>"010000000",
  728=>"001000010",
  729=>"010100000",
  730=>"110111000",
  731=>"011100101",
  732=>"101111000",
  733=>"001010010",
  734=>"001100100",
  735=>"111001111",
  736=>"010111101",
  737=>"100011100",
  738=>"000101001",
  739=>"011111100",
  740=>"011100010",
  741=>"011011001",
  742=>"000110101",
  743=>"000111010",
  744=>"110101001",
  745=>"011011011",
  746=>"001011000",
  747=>"101001011",
  748=>"000101000",
  749=>"100110110",
  750=>"010111000",
  751=>"111100111",
  752=>"001100100",
  753=>"011001111",
  754=>"111111000",
  755=>"010110111",
  756=>"100010101",
  757=>"111000011",
  758=>"011100000",
  759=>"000111011",
  760=>"111110001",
  761=>"100110100",
  762=>"001111001",
  763=>"100010000",
  764=>"010110101",
  765=>"100010100",
  766=>"101001101",
  767=>"010110110",
  768=>"101000101",
  769=>"010001100",
  770=>"100011111",
  771=>"100001111",
  772=>"001101100",
  773=>"001110100",
  774=>"111001101",
  775=>"001101000",
  776=>"000011001",
  777=>"001010001",
  778=>"010010111",
  779=>"101101010",
  780=>"000111000",
  781=>"111011011",
  782=>"110000001",
  783=>"011000000",
  784=>"111000010",
  785=>"000001110",
  786=>"000000111",
  787=>"111100011",
  788=>"101100111",
  789=>"110000111",
  790=>"000111100",
  791=>"011000010",
  792=>"100000101",
  793=>"000110110",
  794=>"001110111",
  795=>"110100000",
  796=>"110011000",
  797=>"101111000",
  798=>"110000100",
  799=>"011101101",
  800=>"000111000",
  801=>"001010101",
  802=>"111001010",
  803=>"100001000",
  804=>"011110001",
  805=>"101011101",
  806=>"001100010",
  807=>"000111101",
  808=>"111010010",
  809=>"010100100",
  810=>"101010101",
  811=>"011000100",
  812=>"111111110",
  813=>"110101110",
  814=>"010001101",
  815=>"010010011",
  816=>"100011001",
  817=>"110111001",
  818=>"100110011",
  819=>"010011011",
  820=>"001110110",
  821=>"111010110",
  822=>"100100110",
  823=>"101000010",
  824=>"101001100",
  825=>"000010101",
  826=>"100111111",
  827=>"100110110",
  828=>"111111100",
  829=>"111011111",
  830=>"101101100",
  831=>"110100001",
  832=>"000100111",
  833=>"100001111",
  834=>"111101001",
  835=>"011000011",
  836=>"010011110",
  837=>"100111111",
  838=>"110111011",
  839=>"001011010",
  840=>"000101111",
  841=>"111101111",
  842=>"100111100",
  843=>"001001101",
  844=>"111010011",
  845=>"111001111",
  846=>"011101001",
  847=>"011011110",
  848=>"010111101",
  849=>"001000011",
  850=>"101101110",
  851=>"001111100",
  852=>"100110101",
  853=>"100011000",
  854=>"111100111",
  855=>"011001010",
  856=>"000110001",
  857=>"100111001",
  858=>"101010110",
  859=>"010001000",
  860=>"100100100",
  861=>"011001110",
  862=>"010110110",
  863=>"010000111",
  864=>"101111000",
  865=>"011000001",
  866=>"100110001",
  867=>"100111100",
  868=>"000000010",
  869=>"001010111",
  870=>"010111110",
  871=>"110001010",
  872=>"111110000",
  873=>"110110111",
  874=>"000100100",
  875=>"110110101",
  876=>"011011110",
  877=>"000010110",
  878=>"100000011",
  879=>"110010000",
  880=>"111101001",
  881=>"011111010",
  882=>"110101100",
  883=>"011000100",
  884=>"100110100",
  885=>"100101100",
  886=>"110011111",
  887=>"110001111",
  888=>"010000000",
  889=>"100011010",
  890=>"011111110",
  891=>"101000110",
  892=>"110011100",
  893=>"111010111",
  894=>"110101000",
  895=>"011101000",
  896=>"001111111",
  897=>"011100110",
  898=>"100101000",
  899=>"111011001",
  900=>"111000100",
  901=>"010010101",
  902=>"101000010",
  903=>"001110000",
  904=>"000101110",
  905=>"100011010",
  906=>"000100010",
  907=>"111111111",
  908=>"011010100",
  909=>"011111001",
  910=>"001111100",
  911=>"101100101",
  912=>"010001101",
  913=>"001010111",
  914=>"000011011",
  915=>"110010010",
  916=>"001111111",
  917=>"010010110",
  918=>"000011010",
  919=>"110000110",
  920=>"100011111",
  921=>"010001111",
  922=>"000110110",
  923=>"001001000",
  924=>"100000111",
  925=>"000000000",
  926=>"011000110",
  927=>"101111110",
  928=>"101111110",
  929=>"100010100",
  930=>"001011000",
  931=>"111000110",
  932=>"111101111",
  933=>"001101111",
  934=>"011111111",
  935=>"111001001",
  936=>"010001000",
  937=>"111011000",
  938=>"110101100",
  939=>"100010000",
  940=>"111000111",
  941=>"001100011",
  942=>"000011111",
  943=>"111010111",
  944=>"111010010",
  945=>"100100101",
  946=>"111010111",
  947=>"000011111",
  948=>"101001010",
  949=>"010010111",
  950=>"100101011",
  951=>"001001101",
  952=>"101111000",
  953=>"001001010",
  954=>"100001111",
  955=>"101010010",
  956=>"110100001",
  957=>"000110110",
  958=>"001111001",
  959=>"001101010",
  960=>"101011111",
  961=>"001000011",
  962=>"000000000",
  963=>"001001111",
  964=>"111101101",
  965=>"011000010",
  966=>"100001111",
  967=>"111101000",
  968=>"001100101",
  969=>"100111001",
  970=>"110101001",
  971=>"010110011",
  972=>"101011111",
  973=>"110110100",
  974=>"010010000",
  975=>"010100000",
  976=>"111111101",
  977=>"000101001",
  978=>"010001000",
  979=>"000010000",
  980=>"010101101",
  981=>"111100101",
  982=>"110101011",
  983=>"100001110",
  984=>"011001110",
  985=>"010100000",
  986=>"010110010",
  987=>"110101010",
  988=>"010011101",
  989=>"101001000",
  990=>"100101000",
  991=>"011110110",
  992=>"110001110",
  993=>"001000111",
  994=>"111000110",
  995=>"011111110",
  996=>"001001001",
  997=>"011000011",
  998=>"000011001",
  999=>"110101111",
  1000=>"111000111",
  1001=>"011100011",
  1002=>"110010011",
  1003=>"011001011",
  1004=>"111010000",
  1005=>"001000010",
  1006=>"000011111",
  1007=>"000011111",
  1008=>"111000100",
  1009=>"111110101",
  1010=>"110010100",
  1011=>"111111011",
  1012=>"001111101",
  1013=>"101110100",
  1014=>"000000010",
  1015=>"101111100",
  1016=>"111000001",
  1017=>"110100111",
  1018=>"110100111",
  1019=>"011111100",
  1020=>"010100010",
  1021=>"101000101",
  1022=>"110100100",
  1023=>"000001001",
  1024=>"001110101",
  1025=>"011011111",
  1026=>"101000000",
  1027=>"010001001",
  1028=>"001001100",
  1029=>"000110110",
  1030=>"101110001",
  1031=>"001101100",
  1032=>"101001001",
  1033=>"011110001",
  1034=>"010111111",
  1035=>"100110001",
  1036=>"001110001",
  1037=>"100111111",
  1038=>"000100010",
  1039=>"000111011",
  1040=>"101111001",
  1041=>"110011111",
  1042=>"011000111",
  1043=>"111001110",
  1044=>"111111100",
  1045=>"100100110",
  1046=>"111100000",
  1047=>"111101111",
  1048=>"010010111",
  1049=>"110111100",
  1050=>"100101101",
  1051=>"111011010",
  1052=>"100010011",
  1053=>"000101101",
  1054=>"001011001",
  1055=>"110000100",
  1056=>"111110101",
  1057=>"111111101",
  1058=>"111101001",
  1059=>"011010001",
  1060=>"100000010",
  1061=>"000110110",
  1062=>"110000111",
  1063=>"010101011",
  1064=>"010011000",
  1065=>"100010000",
  1066=>"110100000",
  1067=>"100001011",
  1068=>"010110010",
  1069=>"100000000",
  1070=>"100010101",
  1071=>"000111010",
  1072=>"000000100",
  1073=>"111011010",
  1074=>"100111111",
  1075=>"010000010",
  1076=>"000101001",
  1077=>"001100011",
  1078=>"010100010",
  1079=>"010000110",
  1080=>"011000001",
  1081=>"111110010",
  1082=>"011111111",
  1083=>"011100101",
  1084=>"010011111",
  1085=>"110000010",
  1086=>"100011000",
  1087=>"111100100",
  1088=>"111111101",
  1089=>"100111000",
  1090=>"000000111",
  1091=>"011001111",
  1092=>"000001101",
  1093=>"100010000",
  1094=>"101000010",
  1095=>"101001110",
  1096=>"100001100",
  1097=>"001000111",
  1098=>"010101010",
  1099=>"100010011",
  1100=>"101001011",
  1101=>"000111001",
  1102=>"101001001",
  1103=>"001000000",
  1104=>"110010011",
  1105=>"010010110",
  1106=>"001010111",
  1107=>"110001000",
  1108=>"100100110",
  1109=>"001110111",
  1110=>"000001100",
  1111=>"010100101",
  1112=>"000001001",
  1113=>"111110100",
  1114=>"110101110",
  1115=>"011011100",
  1116=>"001110001",
  1117=>"100100111",
  1118=>"000100110",
  1119=>"000000011",
  1120=>"100110100",
  1121=>"110001110",
  1122=>"111101010",
  1123=>"011001011",
  1124=>"101101011",
  1125=>"000100110",
  1126=>"011101111",
  1127=>"101010000",
  1128=>"100000111",
  1129=>"110000011",
  1130=>"100101010",
  1131=>"001111100",
  1132=>"010111011",
  1133=>"011010001",
  1134=>"101000100",
  1135=>"110110111",
  1136=>"011000100",
  1137=>"010111010",
  1138=>"110111001",
  1139=>"000000111",
  1140=>"101101111",
  1141=>"101101111",
  1142=>"000001111",
  1143=>"100000110",
  1144=>"111001101",
  1145=>"111001100",
  1146=>"110101110",
  1147=>"100001100",
  1148=>"110000000",
  1149=>"110010011",
  1150=>"001000111",
  1151=>"011101011",
  1152=>"010010000",
  1153=>"011010101",
  1154=>"011100010",
  1155=>"100110100",
  1156=>"000011011",
  1157=>"011010101",
  1158=>"100000110",
  1159=>"010110101",
  1160=>"100011010",
  1161=>"101001100",
  1162=>"010000001",
  1163=>"010100011",
  1164=>"110001101",
  1165=>"111111000",
  1166=>"000000001",
  1167=>"000101010",
  1168=>"000010110",
  1169=>"100110011",
  1170=>"110001101",
  1171=>"001111011",
  1172=>"011001010",
  1173=>"011101001",
  1174=>"110110010",
  1175=>"100111010",
  1176=>"110010010",
  1177=>"111111101",
  1178=>"011100110",
  1179=>"100101101",
  1180=>"000010000",
  1181=>"101101110",
  1182=>"100010010",
  1183=>"111001111",
  1184=>"100111010",
  1185=>"001100101",
  1186=>"110010111",
  1187=>"101001101",
  1188=>"000011000",
  1189=>"111011101",
  1190=>"110000110",
  1191=>"101110101",
  1192=>"100111111",
  1193=>"111101011",
  1194=>"111001111",
  1195=>"011110111",
  1196=>"001011010",
  1197=>"110101101",
  1198=>"010010101",
  1199=>"010100000",
  1200=>"000001101",
  1201=>"110010000",
  1202=>"011101001",
  1203=>"100001010",
  1204=>"111110010",
  1205=>"010100110",
  1206=>"101111110",
  1207=>"110010100",
  1208=>"010011101",
  1209=>"111010010",
  1210=>"001001011",
  1211=>"000010001",
  1212=>"010010011",
  1213=>"010011000",
  1214=>"011110000",
  1215=>"000101010",
  1216=>"000110010",
  1217=>"100001111",
  1218=>"111010010",
  1219=>"111010011",
  1220=>"101101101",
  1221=>"000000010",
  1222=>"010111001",
  1223=>"111101011",
  1224=>"111101110",
  1225=>"000001001",
  1226=>"010011101",
  1227=>"001010001",
  1228=>"011111100",
  1229=>"010000101",
  1230=>"001001011",
  1231=>"010011100",
  1232=>"011000110",
  1233=>"100101111",
  1234=>"010000000",
  1235=>"001100010",
  1236=>"000000111",
  1237=>"100100000",
  1238=>"011011100",
  1239=>"101000010",
  1240=>"010100001",
  1241=>"001100000",
  1242=>"010111111",
  1243=>"100100000",
  1244=>"101011010",
  1245=>"110100000",
  1246=>"101000111",
  1247=>"101000000",
  1248=>"111000100",
  1249=>"100011001",
  1250=>"011111100",
  1251=>"001000000",
  1252=>"111011011",
  1253=>"111111011",
  1254=>"111110100",
  1255=>"101001100",
  1256=>"110111101",
  1257=>"111001001",
  1258=>"001100100",
  1259=>"001011110",
  1260=>"101000010",
  1261=>"011100100",
  1262=>"011100110",
  1263=>"001001010",
  1264=>"111111011",
  1265=>"000011011",
  1266=>"001001000",
  1267=>"001011010",
  1268=>"010000011",
  1269=>"010101000",
  1270=>"010011001",
  1271=>"111011011",
  1272=>"111100010",
  1273=>"101011111",
  1274=>"101101100",
  1275=>"000100010",
  1276=>"010111101",
  1277=>"010100100",
  1278=>"011111110",
  1279=>"011001011",
  1280=>"001100001",
  1281=>"111101010",
  1282=>"001010100",
  1283=>"110001111",
  1284=>"011000000",
  1285=>"101101101",
  1286=>"000111001",
  1287=>"010110101",
  1288=>"101011010",
  1289=>"100000011",
  1290=>"110100100",
  1291=>"010100110",
  1292=>"111111100",
  1293=>"101001111",
  1294=>"010111110",
  1295=>"001010100",
  1296=>"000001101",
  1297=>"011000011",
  1298=>"101100111",
  1299=>"011011101",
  1300=>"111001101",
  1301=>"000000010",
  1302=>"010111110",
  1303=>"001010000",
  1304=>"011001111",
  1305=>"001010000",
  1306=>"111000111",
  1307=>"000101110",
  1308=>"000000010",
  1309=>"110110000",
  1310=>"110110101",
  1311=>"101101101",
  1312=>"010000010",
  1313=>"101001111",
  1314=>"011101111",
  1315=>"000011001",
  1316=>"101010100",
  1317=>"110010111",
  1318=>"000011111",
  1319=>"100100110",
  1320=>"100100101",
  1321=>"110111011",
  1322=>"010101100",
  1323=>"011010111",
  1324=>"001010110",
  1325=>"001101010",
  1326=>"000000011",
  1327=>"010111001",
  1328=>"111111111",
  1329=>"111101001",
  1330=>"000001000",
  1331=>"011100000",
  1332=>"000011100",
  1333=>"010101010",
  1334=>"101001101",
  1335=>"010100001",
  1336=>"101110111",
  1337=>"100000111",
  1338=>"110010000",
  1339=>"011001000",
  1340=>"101011010",
  1341=>"011000001",
  1342=>"010111001",
  1343=>"100100000",
  1344=>"000110011",
  1345=>"101110110",
  1346=>"011111010",
  1347=>"000100100",
  1348=>"110001010",
  1349=>"100010111",
  1350=>"000000101",
  1351=>"011001001",
  1352=>"011100111",
  1353=>"010110000",
  1354=>"111110101",
  1355=>"000101100",
  1356=>"101001101",
  1357=>"101001110",
  1358=>"011110101",
  1359=>"111101010",
  1360=>"000101110",
  1361=>"001110000",
  1362=>"000010100",
  1363=>"110101101",
  1364=>"100101110",
  1365=>"001010111",
  1366=>"110001101",
  1367=>"000011111",
  1368=>"001101111",
  1369=>"100000111",
  1370=>"101001111",
  1371=>"000110101",
  1372=>"010011101",
  1373=>"101001101",
  1374=>"100101101",
  1375=>"110100101",
  1376=>"011000101",
  1377=>"100000011",
  1378=>"111111101",
  1379=>"101000011",
  1380=>"110001100",
  1381=>"011110100",
  1382=>"000000111",
  1383=>"001111000",
  1384=>"111001000",
  1385=>"111100111",
  1386=>"000010110",
  1387=>"010010011",
  1388=>"001011010",
  1389=>"111011011",
  1390=>"000010111",
  1391=>"001101101",
  1392=>"010001100",
  1393=>"100000000",
  1394=>"101001001",
  1395=>"010111100",
  1396=>"010111111",
  1397=>"001011100",
  1398=>"100100111",
  1399=>"000010101",
  1400=>"100000101",
  1401=>"111001110",
  1402=>"111101111",
  1403=>"110000011",
  1404=>"000101111",
  1405=>"000110000",
  1406=>"011010111",
  1407=>"100001110",
  1408=>"000000011",
  1409=>"100101111",
  1410=>"111100011",
  1411=>"011000010",
  1412=>"100011000",
  1413=>"010110001",
  1414=>"111011100",
  1415=>"101010011",
  1416=>"001000000",
  1417=>"111111000",
  1418=>"010010100",
  1419=>"000000010",
  1420=>"010001011",
  1421=>"001000000",
  1422=>"000000011",
  1423=>"000101010",
  1424=>"010010101",
  1425=>"011010010",
  1426=>"100011110",
  1427=>"001101100",
  1428=>"100010111",
  1429=>"001101100",
  1430=>"011010010",
  1431=>"010000100",
  1432=>"100101011",
  1433=>"101000010",
  1434=>"010111101",
  1435=>"000010001",
  1436=>"000101110",
  1437=>"011111111",
  1438=>"001010101",
  1439=>"000101110",
  1440=>"010110010",
  1441=>"001000100",
  1442=>"000100010",
  1443=>"110101110",
  1444=>"100111101",
  1445=>"000100100",
  1446=>"110001101",
  1447=>"000001111",
  1448=>"000110001",
  1449=>"010101111",
  1450=>"111000111",
  1451=>"010111010",
  1452=>"110101101",
  1453=>"011100000",
  1454=>"101100000",
  1455=>"100000111",
  1456=>"111110111",
  1457=>"010000000",
  1458=>"010101011",
  1459=>"001110011",
  1460=>"100100101",
  1461=>"100011010",
  1462=>"101101011",
  1463=>"001111100",
  1464=>"000101001",
  1465=>"001001000",
  1466=>"111101011",
  1467=>"111111011",
  1468=>"010111100",
  1469=>"101000111",
  1470=>"110101011",
  1471=>"110110010",
  1472=>"100100000",
  1473=>"110011101",
  1474=>"100000101",
  1475=>"101000000",
  1476=>"111110111",
  1477=>"000011000",
  1478=>"110111011",
  1479=>"000101100",
  1480=>"111001001",
  1481=>"011001010",
  1482=>"100111111",
  1483=>"011101000",
  1484=>"001000111",
  1485=>"100100010",
  1486=>"001010001",
  1487=>"010010000",
  1488=>"010100000",
  1489=>"100001111",
  1490=>"101001010",
  1491=>"110000010",
  1492=>"100100001",
  1493=>"101011011",
  1494=>"001110010",
  1495=>"010001100",
  1496=>"000001011",
  1497=>"110100010",
  1498=>"111001010",
  1499=>"000011100",
  1500=>"100111010",
  1501=>"100111110",
  1502=>"001110110",
  1503=>"110110000",
  1504=>"111001001",
  1505=>"011001111",
  1506=>"011000000",
  1507=>"001000000",
  1508=>"100001010",
  1509=>"101000100",
  1510=>"000111000",
  1511=>"000001110",
  1512=>"111110101",
  1513=>"001010100",
  1514=>"101110001",
  1515=>"000010011",
  1516=>"000111000",
  1517=>"000010011",
  1518=>"110010100",
  1519=>"011010110",
  1520=>"010010100",
  1521=>"011001001",
  1522=>"110110100",
  1523=>"011010100",
  1524=>"010100001",
  1525=>"101000000",
  1526=>"000000101",
  1527=>"011001101",
  1528=>"000000110",
  1529=>"100110001",
  1530=>"111001111",
  1531=>"000001010",
  1532=>"010001100",
  1533=>"111110010",
  1534=>"000001010",
  1535=>"000001110",
  1536=>"101100011",
  1537=>"101100111",
  1538=>"110101110",
  1539=>"001010110",
  1540=>"000010010",
  1541=>"101001110",
  1542=>"011100100",
  1543=>"110000000",
  1544=>"000011100",
  1545=>"111101111",
  1546=>"000101101",
  1547=>"011100100",
  1548=>"111000000",
  1549=>"011010100",
  1550=>"100000011",
  1551=>"010110111",
  1552=>"011011001",
  1553=>"110110110",
  1554=>"010000011",
  1555=>"111110101",
  1556=>"000001011",
  1557=>"010110011",
  1558=>"000000110",
  1559=>"001000010",
  1560=>"010101000",
  1561=>"110011101",
  1562=>"100000110",
  1563=>"001111111",
  1564=>"110001100",
  1565=>"011111010",
  1566=>"110100111",
  1567=>"111110100",
  1568=>"111000101",
  1569=>"101011111",
  1570=>"111001000",
  1571=>"111100000",
  1572=>"111101011",
  1573=>"010101100",
  1574=>"000110011",
  1575=>"000101010",
  1576=>"001101100",
  1577=>"010101011",
  1578=>"101001000",
  1579=>"111111001",
  1580=>"011001101",
  1581=>"001011110",
  1582=>"111111000",
  1583=>"111000001",
  1584=>"111001000",
  1585=>"000101110",
  1586=>"011001110",
  1587=>"111000111",
  1588=>"100010011",
  1589=>"001100110",
  1590=>"101011101",
  1591=>"000101100",
  1592=>"011101101",
  1593=>"000010000",
  1594=>"001110100",
  1595=>"010011100",
  1596=>"001010110",
  1597=>"001101100",
  1598=>"111010110",
  1599=>"111000100",
  1600=>"110010100",
  1601=>"100101001",
  1602=>"100111000",
  1603=>"011111010",
  1604=>"001010110",
  1605=>"101011111",
  1606=>"101101011",
  1607=>"010111101",
  1608=>"101011001",
  1609=>"100100101",
  1610=>"000001001",
  1611=>"011011101",
  1612=>"100001011",
  1613=>"100001100",
  1614=>"001011110",
  1615=>"111000101",
  1616=>"010111010",
  1617=>"010101101",
  1618=>"101010001",
  1619=>"001101000",
  1620=>"001010010",
  1621=>"010101110",
  1622=>"100000001",
  1623=>"011010111",
  1624=>"000000000",
  1625=>"010010111",
  1626=>"110011010",
  1627=>"111011101",
  1628=>"110011101",
  1629=>"101111111",
  1630=>"011101101",
  1631=>"011011010",
  1632=>"001101010",
  1633=>"110110010",
  1634=>"000010111",
  1635=>"101100101",
  1636=>"100111101",
  1637=>"110001001",
  1638=>"101011000",
  1639=>"101110000",
  1640=>"001100000",
  1641=>"010000111",
  1642=>"100000100",
  1643=>"001111110",
  1644=>"010000101",
  1645=>"000001000",
  1646=>"100011111",
  1647=>"111100000",
  1648=>"000000001",
  1649=>"011000111",
  1650=>"101000101",
  1651=>"100111111",
  1652=>"100000011",
  1653=>"100001110",
  1654=>"101001011",
  1655=>"100100101",
  1656=>"110101011",
  1657=>"100010100",
  1658=>"000100011",
  1659=>"111011110",
  1660=>"011010110",
  1661=>"100011011",
  1662=>"011001110",
  1663=>"100100111",
  1664=>"101100101",
  1665=>"111000000",
  1666=>"101111010",
  1667=>"001010111",
  1668=>"011110100",
  1669=>"010000110",
  1670=>"101001000",
  1671=>"000101101",
  1672=>"101001111",
  1673=>"100000100",
  1674=>"111000011",
  1675=>"110010111",
  1676=>"001001101",
  1677=>"010110010",
  1678=>"100111111",
  1679=>"011000000",
  1680=>"100110001",
  1681=>"001101101",
  1682=>"001100010",
  1683=>"011110000",
  1684=>"111011001",
  1685=>"010100010",
  1686=>"001111111",
  1687=>"111000110",
  1688=>"000000100",
  1689=>"101110000",
  1690=>"001111110",
  1691=>"011000111",
  1692=>"101010010",
  1693=>"001111000",
  1694=>"110101110",
  1695=>"001111101",
  1696=>"101100011",
  1697=>"101001101",
  1698=>"000001010",
  1699=>"000010110",
  1700=>"000100100",
  1701=>"110001101",
  1702=>"001011111",
  1703=>"011010010",
  1704=>"001001010",
  1705=>"010001110",
  1706=>"010011101",
  1707=>"010101101",
  1708=>"111101000",
  1709=>"110001001",
  1710=>"011000111",
  1711=>"111111001",
  1712=>"100001011",
  1713=>"110101000",
  1714=>"010101110",
  1715=>"110111110",
  1716=>"101001011",
  1717=>"000000001",
  1718=>"011010100",
  1719=>"010000011",
  1720=>"101101010",
  1721=>"000010110",
  1722=>"010110101",
  1723=>"010000101",
  1724=>"000101011",
  1725=>"100111001",
  1726=>"000101010",
  1727=>"100010010",
  1728=>"101011100",
  1729=>"010110011",
  1730=>"111001111",
  1731=>"011011100",
  1732=>"111111010",
  1733=>"001011100",
  1734=>"110111001",
  1735=>"101011011",
  1736=>"111001101",
  1737=>"101110100",
  1738=>"111111001",
  1739=>"000100001",
  1740=>"111111011",
  1741=>"001101111",
  1742=>"000101110",
  1743=>"011011101",
  1744=>"111110110",
  1745=>"101110010",
  1746=>"101101001",
  1747=>"001100000",
  1748=>"011100101",
  1749=>"101111101",
  1750=>"100010001",
  1751=>"011001011",
  1752=>"001000111",
  1753=>"011100010",
  1754=>"011110010",
  1755=>"100111011",
  1756=>"111011011",
  1757=>"010111011",
  1758=>"100001110",
  1759=>"110101011",
  1760=>"110001111",
  1761=>"101010100",
  1762=>"100111001",
  1763=>"000100001",
  1764=>"010010100",
  1765=>"101011000",
  1766=>"110101010",
  1767=>"111000100",
  1768=>"111110011",
  1769=>"111010000",
  1770=>"000100000",
  1771=>"110110101",
  1772=>"001011100",
  1773=>"001100011",
  1774=>"010100001",
  1775=>"000000010",
  1776=>"110111001",
  1777=>"111011000",
  1778=>"100010000",
  1779=>"000110010",
  1780=>"111101111",
  1781=>"000011110",
  1782=>"101011001",
  1783=>"100000101",
  1784=>"110001010",
  1785=>"100001110",
  1786=>"111010011",
  1787=>"000100000",
  1788=>"110000000",
  1789=>"000010011",
  1790=>"101110111",
  1791=>"001000101",
  1792=>"100000111",
  1793=>"011110001",
  1794=>"011101111",
  1795=>"010100111",
  1796=>"100111111",
  1797=>"101111101",
  1798=>"011000111",
  1799=>"010111100",
  1800=>"100010011",
  1801=>"100110010",
  1802=>"011011010",
  1803=>"111101111",
  1804=>"110100010",
  1805=>"001110110",
  1806=>"100101001",
  1807=>"010010000",
  1808=>"101010110",
  1809=>"011011001",
  1810=>"010110001",
  1811=>"010100111",
  1812=>"001110001",
  1813=>"111110100",
  1814=>"111110111",
  1815=>"111101111",
  1816=>"101100000",
  1817=>"101001011",
  1818=>"000001111",
  1819=>"010111100",
  1820=>"000011010",
  1821=>"110001010",
  1822=>"100110110",
  1823=>"110101110",
  1824=>"000001000",
  1825=>"011010101",
  1826=>"010000111",
  1827=>"001111001",
  1828=>"100001011",
  1829=>"010010100",
  1830=>"000100001",
  1831=>"101100110",
  1832=>"111000111",
  1833=>"001001100",
  1834=>"100101110",
  1835=>"011010001",
  1836=>"110101000",
  1837=>"010010010",
  1838=>"010001001",
  1839=>"101000011",
  1840=>"000000010",
  1841=>"101000010",
  1842=>"000011000",
  1843=>"011101100",
  1844=>"110100000",
  1845=>"011101111",
  1846=>"100001100",
  1847=>"011010111",
  1848=>"011111011",
  1849=>"010100110",
  1850=>"100100001",
  1851=>"111110010",
  1852=>"110001010",
  1853=>"011000001",
  1854=>"011011000",
  1855=>"001101001",
  1856=>"101000111",
  1857=>"110100010",
  1858=>"000000000",
  1859=>"000100100",
  1860=>"100101010",
  1861=>"001001111",
  1862=>"110101100",
  1863=>"111011010",
  1864=>"010100010",
  1865=>"010010000",
  1866=>"010100010",
  1867=>"001000001",
  1868=>"110000101",
  1869=>"111000011",
  1870=>"110101111",
  1871=>"001111000",
  1872=>"000000000",
  1873=>"101001100",
  1874=>"111111011",
  1875=>"111111101",
  1876=>"000110101",
  1877=>"101101100",
  1878=>"000111100",
  1879=>"011001101",
  1880=>"110001101",
  1881=>"011001101",
  1882=>"011111001",
  1883=>"010110011",
  1884=>"001011001",
  1885=>"101001111",
  1886=>"011000010",
  1887=>"110101001",
  1888=>"010000011",
  1889=>"101011001",
  1890=>"011001111",
  1891=>"100011100",
  1892=>"001100010",
  1893=>"000110000",
  1894=>"111001101",
  1895=>"011000011",
  1896=>"001101010",
  1897=>"100111101",
  1898=>"110000010",
  1899=>"000100011",
  1900=>"101011010",
  1901=>"010100010",
  1902=>"011111111",
  1903=>"011110110",
  1904=>"000100001",
  1905=>"000110001",
  1906=>"101101000",
  1907=>"110011110",
  1908=>"110011101",
  1909=>"111100011",
  1910=>"101110000",
  1911=>"101100100",
  1912=>"100101111",
  1913=>"101111010",
  1914=>"110000000",
  1915=>"100111011",
  1916=>"001000100",
  1917=>"011100001",
  1918=>"010100011",
  1919=>"110111101",
  1920=>"010111110",
  1921=>"111110111",
  1922=>"110110000",
  1923=>"110001011",
  1924=>"100100110",
  1925=>"111011001",
  1926=>"101111011",
  1927=>"101111011",
  1928=>"111100101",
  1929=>"010101100",
  1930=>"001000111",
  1931=>"011000010",
  1932=>"101011011",
  1933=>"110101111",
  1934=>"100010011",
  1935=>"010001111",
  1936=>"010000010",
  1937=>"001111010",
  1938=>"100000011",
  1939=>"100111011",
  1940=>"011101111",
  1941=>"001111011",
  1942=>"010111011",
  1943=>"110100010",
  1944=>"010110011",
  1945=>"110010110",
  1946=>"111011111",
  1947=>"101010000",
  1948=>"001000110",
  1949=>"101111101",
  1950=>"010011010",
  1951=>"101101011",
  1952=>"100101101",
  1953=>"110001001",
  1954=>"100110000",
  1955=>"001010111",
  1956=>"110010000",
  1957=>"001100100",
  1958=>"011011111",
  1959=>"000011011",
  1960=>"101100001",
  1961=>"111110011",
  1962=>"100001111",
  1963=>"000111001",
  1964=>"011100001",
  1965=>"111011010",
  1966=>"011111001",
  1967=>"110001101",
  1968=>"000010111",
  1969=>"000110111",
  1970=>"010000010",
  1971=>"101111101",
  1972=>"110001011",
  1973=>"001011011",
  1974=>"110110010",
  1975=>"001111100",
  1976=>"001110111",
  1977=>"000110011",
  1978=>"001001101",
  1979=>"000111001",
  1980=>"110111011",
  1981=>"000010100",
  1982=>"111100011",
  1983=>"000111011",
  1984=>"101010100",
  1985=>"101110010",
  1986=>"001100111",
  1987=>"100101111",
  1988=>"100001111",
  1989=>"110110100",
  1990=>"001100011",
  1991=>"000000001",
  1992=>"110000001",
  1993=>"100110110",
  1994=>"010011101",
  1995=>"110000100",
  1996=>"110101100",
  1997=>"001100000",
  1998=>"101000110",
  1999=>"110001011",
  2000=>"100010100",
  2001=>"000100011",
  2002=>"001110001",
  2003=>"100101100",
  2004=>"110000011",
  2005=>"100111000",
  2006=>"110101000",
  2007=>"110110010",
  2008=>"000110000",
  2009=>"111111110",
  2010=>"110100111",
  2011=>"001101101",
  2012=>"010010110",
  2013=>"111101111",
  2014=>"011110010",
  2015=>"000000000",
  2016=>"000110100",
  2017=>"110000000",
  2018=>"011011010",
  2019=>"011111001",
  2020=>"000110001",
  2021=>"001110100",
  2022=>"000100000",
  2023=>"101000001",
  2024=>"101010001",
  2025=>"001101001",
  2026=>"001110110",
  2027=>"111001010",
  2028=>"110001100",
  2029=>"100111011",
  2030=>"111001111",
  2031=>"111111010",
  2032=>"100011000",
  2033=>"100010010",
  2034=>"000000110",
  2035=>"100100000",
  2036=>"000001010",
  2037=>"000110101",
  2038=>"111111101",
  2039=>"011000011",
  2040=>"101101110",
  2041=>"111010101",
  2042=>"110010010",
  2043=>"111011000",
  2044=>"001011110",
  2045=>"000011001",
  2046=>"010101100",
  2047=>"011011001",
  2048=>"001110110",
  2049=>"110111011",
  2050=>"011000010",
  2051=>"101001010",
  2052=>"000010110",
  2053=>"001011001",
  2054=>"100000101",
  2055=>"111101000",
  2056=>"101110010",
  2057=>"110110011",
  2058=>"110101001",
  2059=>"010101100",
  2060=>"111001010",
  2061=>"111010101",
  2062=>"010010100",
  2063=>"011000000",
  2064=>"110001110",
  2065=>"111010101",
  2066=>"111010101",
  2067=>"100001000",
  2068=>"000011011",
  2069=>"011111111",
  2070=>"101000000",
  2071=>"011011101",
  2072=>"100010011",
  2073=>"000101100",
  2074=>"011111110",
  2075=>"111111110",
  2076=>"101000100",
  2077=>"001000010",
  2078=>"101010000",
  2079=>"010100011",
  2080=>"101111001",
  2081=>"101010000",
  2082=>"101110101",
  2083=>"011100001",
  2084=>"000001000",
  2085=>"011111000",
  2086=>"000010010",
  2087=>"001111011",
  2088=>"000111100",
  2089=>"111111111",
  2090=>"010000101",
  2091=>"001010011",
  2092=>"101010010",
  2093=>"101001001",
  2094=>"000111011",
  2095=>"111011011",
  2096=>"010100011",
  2097=>"100100100",
  2098=>"111001101",
  2099=>"100010001",
  2100=>"101000000",
  2101=>"100100101",
  2102=>"101010010",
  2103=>"010001110",
  2104=>"010011011",
  2105=>"110010010",
  2106=>"001011110",
  2107=>"010010100",
  2108=>"111011011",
  2109=>"011001111",
  2110=>"001010100",
  2111=>"000011100",
  2112=>"100011100",
  2113=>"001000011",
  2114=>"100110110",
  2115=>"110000000",
  2116=>"001001000",
  2117=>"010001001",
  2118=>"110110011",
  2119=>"111011101",
  2120=>"000101000",
  2121=>"110001101",
  2122=>"000010111",
  2123=>"100110111",
  2124=>"010011000",
  2125=>"100000011",
  2126=>"001100110",
  2127=>"111101100",
  2128=>"111110110",
  2129=>"011001111",
  2130=>"001100110",
  2131=>"011101000",
  2132=>"001101110",
  2133=>"101110000",
  2134=>"100011000",
  2135=>"100000000",
  2136=>"010100110",
  2137=>"110111110",
  2138=>"101001110",
  2139=>"001000000",
  2140=>"101101100",
  2141=>"101100001",
  2142=>"111011010",
  2143=>"001001001",
  2144=>"000010100",
  2145=>"010011111",
  2146=>"101110111",
  2147=>"011010000",
  2148=>"000011000",
  2149=>"100111010",
  2150=>"101001000",
  2151=>"011000000",
  2152=>"100011100",
  2153=>"011110101",
  2154=>"000111111",
  2155=>"110000100",
  2156=>"011001010",
  2157=>"011111011",
  2158=>"010011001",
  2159=>"001011001",
  2160=>"101010100",
  2161=>"111010000",
  2162=>"001100101",
  2163=>"001000001",
  2164=>"001010010",
  2165=>"100111101",
  2166=>"110100000",
  2167=>"100111001",
  2168=>"011101010",
  2169=>"011111001",
  2170=>"010100000",
  2171=>"001100001",
  2172=>"111010111",
  2173=>"010010010",
  2174=>"101101010",
  2175=>"001110000",
  2176=>"111000000",
  2177=>"111000110",
  2178=>"110100110",
  2179=>"100110001",
  2180=>"100101100",
  2181=>"100010110",
  2182=>"100110011",
  2183=>"001001001",
  2184=>"010010000",
  2185=>"111000000",
  2186=>"000100101",
  2187=>"011111100",
  2188=>"011010111",
  2189=>"010101101",
  2190=>"010111101",
  2191=>"011110100",
  2192=>"011001011",
  2193=>"011011010",
  2194=>"001010010",
  2195=>"111110000",
  2196=>"000111001",
  2197=>"111000000",
  2198=>"111000010",
  2199=>"100001101",
  2200=>"010001110",
  2201=>"110111110",
  2202=>"001110010",
  2203=>"001110111",
  2204=>"110110000",
  2205=>"101011100",
  2206=>"000110000",
  2207=>"111000101",
  2208=>"110100100",
  2209=>"001010001",
  2210=>"011010010",
  2211=>"000000000",
  2212=>"001001111",
  2213=>"011101111",
  2214=>"010010010",
  2215=>"011001001",
  2216=>"001100101",
  2217=>"001010101",
  2218=>"100000111",
  2219=>"010010001",
  2220=>"100011111",
  2221=>"011100001",
  2222=>"100100110",
  2223=>"011000011",
  2224=>"011110110",
  2225=>"001111000",
  2226=>"001101110",
  2227=>"100100000",
  2228=>"100000101",
  2229=>"000110101",
  2230=>"001110101",
  2231=>"011111110",
  2232=>"100011110",
  2233=>"100111001",
  2234=>"000011100",
  2235=>"100111111",
  2236=>"010111010",
  2237=>"101010001",
  2238=>"000110100",
  2239=>"010100110",
  2240=>"010110111",
  2241=>"111100011",
  2242=>"110110001",
  2243=>"100010011",
  2244=>"100000011",
  2245=>"001011011",
  2246=>"010101100",
  2247=>"111001111",
  2248=>"011111000",
  2249=>"001110001",
  2250=>"011101011",
  2251=>"011111001",
  2252=>"011010001",
  2253=>"011101110",
  2254=>"000111101",
  2255=>"110111000",
  2256=>"101001101",
  2257=>"111100101",
  2258=>"101110000",
  2259=>"110010011",
  2260=>"111111101",
  2261=>"010000111",
  2262=>"011010000",
  2263=>"100000010",
  2264=>"101110111",
  2265=>"110110110",
  2266=>"001111100",
  2267=>"011010001",
  2268=>"101000111",
  2269=>"001111100",
  2270=>"011010000",
  2271=>"111111001",
  2272=>"111011101",
  2273=>"000100110",
  2274=>"001011111",
  2275=>"110000110",
  2276=>"000100001",
  2277=>"111111110",
  2278=>"001101001",
  2279=>"010100000",
  2280=>"110101001",
  2281=>"001111110",
  2282=>"110000010",
  2283=>"010010100",
  2284=>"101001000",
  2285=>"000001100",
  2286=>"101001110",
  2287=>"001101101",
  2288=>"111100001",
  2289=>"001011010",
  2290=>"001010011",
  2291=>"000100110",
  2292=>"101001001",
  2293=>"011000010",
  2294=>"111000100",
  2295=>"010010001",
  2296=>"011000111",
  2297=>"100110110",
  2298=>"111101110",
  2299=>"001100011",
  2300=>"111111100",
  2301=>"100000110",
  2302=>"010100001",
  2303=>"011010110",
  2304=>"011001101",
  2305=>"001001011",
  2306=>"101010011",
  2307=>"100100010",
  2308=>"101100010",
  2309=>"101011100",
  2310=>"101011101",
  2311=>"111001000",
  2312=>"100000111",
  2313=>"011101010",
  2314=>"111010111",
  2315=>"101010010",
  2316=>"110011100",
  2317=>"100000010",
  2318=>"101000011",
  2319=>"101011010",
  2320=>"001111100",
  2321=>"000101010",
  2322=>"100110001",
  2323=>"111111101",
  2324=>"110101101",
  2325=>"111001011",
  2326=>"011000101",
  2327=>"010001010",
  2328=>"110100100",
  2329=>"001011010",
  2330=>"000011110",
  2331=>"001011100",
  2332=>"010100010",
  2333=>"000011000",
  2334=>"010111010",
  2335=>"100000000",
  2336=>"110110000",
  2337=>"110011111",
  2338=>"010001100",
  2339=>"010011001",
  2340=>"000001100",
  2341=>"111011000",
  2342=>"110100001",
  2343=>"001110100",
  2344=>"001111111",
  2345=>"111100000",
  2346=>"101101101",
  2347=>"001001001",
  2348=>"111111010",
  2349=>"010000010",
  2350=>"011111100",
  2351=>"000001111",
  2352=>"010101100",
  2353=>"111101000",
  2354=>"100011111",
  2355=>"110111000",
  2356=>"011011001",
  2357=>"000000000",
  2358=>"110100000",
  2359=>"001001111",
  2360=>"011100000",
  2361=>"101101011",
  2362=>"111010000",
  2363=>"111010011",
  2364=>"110010110",
  2365=>"010110100",
  2366=>"101010100",
  2367=>"111110110",
  2368=>"100011111",
  2369=>"101001101",
  2370=>"100110111",
  2371=>"000001100",
  2372=>"111010000",
  2373=>"010011110",
  2374=>"000000010",
  2375=>"111101111",
  2376=>"001101111",
  2377=>"000001000",
  2378=>"100011010",
  2379=>"000100111",
  2380=>"001111011",
  2381=>"100110110",
  2382=>"101000101",
  2383=>"100011000",
  2384=>"101011101",
  2385=>"000001010",
  2386=>"010011010",
  2387=>"010000011",
  2388=>"010100011",
  2389=>"101111010",
  2390=>"110010001",
  2391=>"100100111",
  2392=>"111010011",
  2393=>"001000100",
  2394=>"101001111",
  2395=>"001101010",
  2396=>"000100110",
  2397=>"101100011",
  2398=>"100101000",
  2399=>"011110010",
  2400=>"111000110",
  2401=>"100011110",
  2402=>"000001001",
  2403=>"111101111",
  2404=>"000101000",
  2405=>"111011000",
  2406=>"010011111",
  2407=>"010100100",
  2408=>"001100100",
  2409=>"111110010",
  2410=>"111101110",
  2411=>"011010101",
  2412=>"011100000",
  2413=>"100001010",
  2414=>"110010100",
  2415=>"100000001",
  2416=>"100100001",
  2417=>"000011011",
  2418=>"101110111",
  2419=>"110110100",
  2420=>"001010001",
  2421=>"101110111",
  2422=>"111101010",
  2423=>"001010010",
  2424=>"010000000",
  2425=>"000001011",
  2426=>"111100111",
  2427=>"010000110",
  2428=>"111101100",
  2429=>"000000101",
  2430=>"111111001",
  2431=>"010000010",
  2432=>"001010010",
  2433=>"010100101",
  2434=>"101000101",
  2435=>"100001100",
  2436=>"110110001",
  2437=>"000110100",
  2438=>"000100000",
  2439=>"011100101",
  2440=>"101101001",
  2441=>"000001000",
  2442=>"110111101",
  2443=>"110111011",
  2444=>"000100111",
  2445=>"100111000",
  2446=>"100000100",
  2447=>"001100101",
  2448=>"001011010",
  2449=>"111000010",
  2450=>"100001000",
  2451=>"001001101",
  2452=>"100100101",
  2453=>"000000001",
  2454=>"101010110",
  2455=>"001010100",
  2456=>"111001100",
  2457=>"000110100",
  2458=>"111101001",
  2459=>"000111101",
  2460=>"110010100",
  2461=>"011010110",
  2462=>"110100110",
  2463=>"101100000",
  2464=>"101100101",
  2465=>"111110010",
  2466=>"101011111",
  2467=>"010000001",
  2468=>"001111000",
  2469=>"100001001",
  2470=>"000000011",
  2471=>"010000101",
  2472=>"110101101",
  2473=>"000010011",
  2474=>"001000010",
  2475=>"100101000",
  2476=>"111100001",
  2477=>"101110110",
  2478=>"000011111",
  2479=>"110111111",
  2480=>"110000001",
  2481=>"110010000",
  2482=>"010011001",
  2483=>"010100110",
  2484=>"111110110",
  2485=>"000100111",
  2486=>"111100011",
  2487=>"010111001",
  2488=>"110111101",
  2489=>"101000001",
  2490=>"101000010",
  2491=>"001110001",
  2492=>"100011110",
  2493=>"100100011",
  2494=>"000101000",
  2495=>"110111101",
  2496=>"001010010",
  2497=>"001110011",
  2498=>"100011000",
  2499=>"111101100",
  2500=>"100000011",
  2501=>"001001011",
  2502=>"011010011",
  2503=>"110111111",
  2504=>"111111011",
  2505=>"100100110",
  2506=>"011100001",
  2507=>"101111011",
  2508=>"010110001",
  2509=>"110111110",
  2510=>"010000110",
  2511=>"101001000",
  2512=>"111000000",
  2513=>"111011000",
  2514=>"100100100",
  2515=>"011100000",
  2516=>"111110010",
  2517=>"011110110",
  2518=>"000101000",
  2519=>"001110011",
  2520=>"100111000",
  2521=>"000000011",
  2522=>"001010000",
  2523=>"100110000",
  2524=>"111111110",
  2525=>"010010000",
  2526=>"011101111",
  2527=>"010110010",
  2528=>"100101101",
  2529=>"000011110",
  2530=>"100111000",
  2531=>"100110100",
  2532=>"001010010",
  2533=>"111010011",
  2534=>"110010000",
  2535=>"111000001",
  2536=>"001101001",
  2537=>"110000010",
  2538=>"000000110",
  2539=>"010000011",
  2540=>"111010110",
  2541=>"110001101",
  2542=>"100100110",
  2543=>"001111010",
  2544=>"110111111",
  2545=>"000011000",
  2546=>"100010111",
  2547=>"101000000",
  2548=>"101010001",
  2549=>"111011111",
  2550=>"100100101",
  2551=>"111100110",
  2552=>"110111110",
  2553=>"000101101",
  2554=>"000111000",
  2555=>"011000110",
  2556=>"100101111",
  2557=>"010010111",
  2558=>"100101100",
  2559=>"010010011",
  2560=>"100101101",
  2561=>"000110011",
  2562=>"101000001",
  2563=>"001010001",
  2564=>"000000100",
  2565=>"101101101",
  2566=>"000101000",
  2567=>"101110110",
  2568=>"001011100",
  2569=>"010010110",
  2570=>"000111101",
  2571=>"001001011",
  2572=>"010001111",
  2573=>"101011010",
  2574=>"011010101",
  2575=>"101011111",
  2576=>"010001111",
  2577=>"011100000",
  2578=>"101010001",
  2579=>"101010100",
  2580=>"000000001",
  2581=>"100111101",
  2582=>"001000110",
  2583=>"010001101",
  2584=>"010001101",
  2585=>"001111101",
  2586=>"110100111",
  2587=>"100101000",
  2588=>"000100100",
  2589=>"011100001",
  2590=>"000111011",
  2591=>"010010001",
  2592=>"101001111",
  2593=>"001111111",
  2594=>"111000110",
  2595=>"000100101",
  2596=>"001101111",
  2597=>"110000011",
  2598=>"111110010",
  2599=>"000001000",
  2600=>"001011011",
  2601=>"011010100",
  2602=>"101010111",
  2603=>"100110111",
  2604=>"001000011",
  2605=>"001100101",
  2606=>"111100101",
  2607=>"101011100",
  2608=>"001010111",
  2609=>"000001110",
  2610=>"001010101",
  2611=>"110001100",
  2612=>"000000000",
  2613=>"111111001",
  2614=>"001010111",
  2615=>"011101100",
  2616=>"100011010",
  2617=>"010101110",
  2618=>"100100011",
  2619=>"111000011",
  2620=>"010000110",
  2621=>"000010000",
  2622=>"110001110",
  2623=>"100100000",
  2624=>"101101111",
  2625=>"000111010",
  2626=>"100000010",
  2627=>"111111011",
  2628=>"000010000",
  2629=>"011100110",
  2630=>"100001011",
  2631=>"101110011",
  2632=>"000000000",
  2633=>"110010010",
  2634=>"010011111",
  2635=>"110110111",
  2636=>"001111110",
  2637=>"000000000",
  2638=>"111111111",
  2639=>"111001111",
  2640=>"010011000",
  2641=>"110110100",
  2642=>"011001111",
  2643=>"001011101",
  2644=>"000011111",
  2645=>"011010111",
  2646=>"000011100",
  2647=>"110001010",
  2648=>"010110110",
  2649=>"011000110",
  2650=>"101010010",
  2651=>"000001100",
  2652=>"010000000",
  2653=>"111101110",
  2654=>"110000100",
  2655=>"010100011",
  2656=>"011001100",
  2657=>"111100110",
  2658=>"101010101",
  2659=>"100111001",
  2660=>"000011110",
  2661=>"100000101",
  2662=>"100001011",
  2663=>"100100000",
  2664=>"101000001",
  2665=>"001111101",
  2666=>"100000011",
  2667=>"100111010",
  2668=>"100101011",
  2669=>"011101110",
  2670=>"110100001",
  2671=>"011111000",
  2672=>"110111011",
  2673=>"100100111",
  2674=>"101101100",
  2675=>"101101010",
  2676=>"101111101",
  2677=>"000111000",
  2678=>"100011111",
  2679=>"111110001",
  2680=>"100000110",
  2681=>"101100000",
  2682=>"100100001",
  2683=>"101110101",
  2684=>"010000001",
  2685=>"100100101",
  2686=>"111100000",
  2687=>"100100011",
  2688=>"001010011",
  2689=>"111001010",
  2690=>"000000011",
  2691=>"011001110",
  2692=>"000000000",
  2693=>"100101001",
  2694=>"010001100",
  2695=>"001010011",
  2696=>"001011010",
  2697=>"111101001",
  2698=>"100111110",
  2699=>"100110110",
  2700=>"100111000",
  2701=>"111101101",
  2702=>"010101100",
  2703=>"110100110",
  2704=>"111111001",
  2705=>"001111001",
  2706=>"001000100",
  2707=>"110010101",
  2708=>"010100111",
  2709=>"001001000",
  2710=>"101011010",
  2711=>"111111011",
  2712=>"100000000",
  2713=>"001100111",
  2714=>"000010000",
  2715=>"101010101",
  2716=>"001101111",
  2717=>"110100000",
  2718=>"001111001",
  2719=>"011101111",
  2720=>"000000000",
  2721=>"101000000",
  2722=>"010110111",
  2723=>"000000110",
  2724=>"001101111",
  2725=>"000011111",
  2726=>"111111110",
  2727=>"001000011",
  2728=>"010110101",
  2729=>"100010000",
  2730=>"101010100",
  2731=>"011010100",
  2732=>"111100001",
  2733=>"010011110",
  2734=>"010101001",
  2735=>"101101101",
  2736=>"100111111",
  2737=>"001111111",
  2738=>"100110111",
  2739=>"001110111",
  2740=>"101110100",
  2741=>"001011001",
  2742=>"100110000",
  2743=>"101100110",
  2744=>"000011110",
  2745=>"100101110",
  2746=>"110100011",
  2747=>"111010111",
  2748=>"010111101",
  2749=>"111110101",
  2750=>"000011101",
  2751=>"100111100",
  2752=>"010010110",
  2753=>"111001100",
  2754=>"111011100",
  2755=>"010110001",
  2756=>"001101011",
  2757=>"111001111",
  2758=>"000111101",
  2759=>"001110001",
  2760=>"011101111",
  2761=>"101001011",
  2762=>"111010010",
  2763=>"101100001",
  2764=>"110100011",
  2765=>"011110100",
  2766=>"010110011",
  2767=>"011110001",
  2768=>"111111011",
  2769=>"111010001",
  2770=>"101011110",
  2771=>"011000110",
  2772=>"001100100",
  2773=>"011010111",
  2774=>"000000100",
  2775=>"011000000",
  2776=>"110011001",
  2777=>"011010000",
  2778=>"000100010",
  2779=>"010010000",
  2780=>"000111111",
  2781=>"110010101",
  2782=>"101101010",
  2783=>"000010101",
  2784=>"100110111",
  2785=>"001111011",
  2786=>"101011001",
  2787=>"100110101",
  2788=>"001100101",
  2789=>"000001000",
  2790=>"101001111",
  2791=>"110110011",
  2792=>"001010001",
  2793=>"011110010",
  2794=>"010100111",
  2795=>"001010100",
  2796=>"011000000",
  2797=>"010100110",
  2798=>"100111111",
  2799=>"110010110",
  2800=>"111101011",
  2801=>"001000101",
  2802=>"100000100",
  2803=>"001001011",
  2804=>"110101111",
  2805=>"010001110",
  2806=>"111011001",
  2807=>"101010001",
  2808=>"000001010",
  2809=>"000001101",
  2810=>"101101001",
  2811=>"110001100",
  2812=>"110011001",
  2813=>"010001101",
  2814=>"100000010",
  2815=>"111111010",
  2816=>"100100001",
  2817=>"101110001",
  2818=>"001111000",
  2819=>"010110011",
  2820=>"010010010",
  2821=>"011000000",
  2822=>"011111110",
  2823=>"000010010",
  2824=>"101000000",
  2825=>"000111011",
  2826=>"110001001",
  2827=>"011011010",
  2828=>"100001011",
  2829=>"111100100",
  2830=>"111010101",
  2831=>"001101101",
  2832=>"001100101",
  2833=>"010110111",
  2834=>"100110010",
  2835=>"101100001",
  2836=>"000000001",
  2837=>"010001010",
  2838=>"100101101",
  2839=>"011010011",
  2840=>"001110001",
  2841=>"011111101",
  2842=>"101001000",
  2843=>"100011110",
  2844=>"011100000",
  2845=>"101111110",
  2846=>"000111110",
  2847=>"101111001",
  2848=>"110100101",
  2849=>"011001111",
  2850=>"101111011",
  2851=>"011100000",
  2852=>"011100000",
  2853=>"000111001",
  2854=>"010110001",
  2855=>"110101001",
  2856=>"110010100",
  2857=>"100110100",
  2858=>"111010001",
  2859=>"101110011",
  2860=>"100100111",
  2861=>"011001100",
  2862=>"001101000",
  2863=>"101100011",
  2864=>"000100110",
  2865=>"111110011",
  2866=>"101010110",
  2867=>"011110100",
  2868=>"000011011",
  2869=>"010011111",
  2870=>"110011100",
  2871=>"010001000",
  2872=>"001011111",
  2873=>"100001001",
  2874=>"111111110",
  2875=>"111101101",
  2876=>"100001110",
  2877=>"110110000",
  2878=>"011001101",
  2879=>"111001010",
  2880=>"000100011",
  2881=>"100001011",
  2882=>"111000010",
  2883=>"011110110",
  2884=>"111101110",
  2885=>"010111100",
  2886=>"100000100",
  2887=>"011111100",
  2888=>"001111110",
  2889=>"111001000",
  2890=>"111110001",
  2891=>"000010000",
  2892=>"000101100",
  2893=>"100100011",
  2894=>"011111110",
  2895=>"000000100",
  2896=>"010000110",
  2897=>"101110101",
  2898=>"001100110",
  2899=>"101111000",
  2900=>"001101110",
  2901=>"000101101",
  2902=>"111010101",
  2903=>"100100110",
  2904=>"000110111",
  2905=>"001000101",
  2906=>"101111110",
  2907=>"101001100",
  2908=>"101000000",
  2909=>"011010010",
  2910=>"001001000",
  2911=>"110110100",
  2912=>"000011000",
  2913=>"101101001",
  2914=>"001101101",
  2915=>"100001011",
  2916=>"010001111",
  2917=>"110111000",
  2918=>"111001000",
  2919=>"111011101",
  2920=>"000010000",
  2921=>"011100001",
  2922=>"001001101",
  2923=>"001001001",
  2924=>"110011011",
  2925=>"110011000",
  2926=>"110001011",
  2927=>"011111101",
  2928=>"100010000",
  2929=>"110111110",
  2930=>"011001011",
  2931=>"111001010",
  2932=>"010001000",
  2933=>"111100100",
  2934=>"000111101",
  2935=>"001110000",
  2936=>"111000100",
  2937=>"110011011",
  2938=>"101110111",
  2939=>"110110011",
  2940=>"111100000",
  2941=>"010011110",
  2942=>"001111000",
  2943=>"110011110",
  2944=>"011000100",
  2945=>"101001001",
  2946=>"101110011",
  2947=>"110000110",
  2948=>"000111101",
  2949=>"100011111",
  2950=>"011010010",
  2951=>"000110000",
  2952=>"110011011",
  2953=>"011111010",
  2954=>"011110111",
  2955=>"101111000",
  2956=>"100001101",
  2957=>"011001011",
  2958=>"111111001",
  2959=>"010001110",
  2960=>"111101011",
  2961=>"000111110",
  2962=>"101100111",
  2963=>"011111001",
  2964=>"001000001",
  2965=>"010011111",
  2966=>"000101000",
  2967=>"010010111",
  2968=>"001111000",
  2969=>"100100101",
  2970=>"000010010",
  2971=>"110011000",
  2972=>"100100100",
  2973=>"001000010",
  2974=>"000000011",
  2975=>"110011000",
  2976=>"001011110",
  2977=>"000111110",
  2978=>"001001000",
  2979=>"010101000",
  2980=>"111011001",
  2981=>"100001111",
  2982=>"111100011",
  2983=>"111010110",
  2984=>"101001100",
  2985=>"000011000",
  2986=>"110011011",
  2987=>"000011111",
  2988=>"101011001",
  2989=>"101011001",
  2990=>"000111010",
  2991=>"010100110",
  2992=>"111000010",
  2993=>"001001000",
  2994=>"010011100",
  2995=>"001000011",
  2996=>"011101000",
  2997=>"001000010",
  2998=>"111111110",
  2999=>"101101001",
  3000=>"010010110",
  3001=>"001011100",
  3002=>"010000011",
  3003=>"100000111",
  3004=>"111011111",
  3005=>"000001011",
  3006=>"011010001",
  3007=>"110110100",
  3008=>"011100011",
  3009=>"111111111",
  3010=>"011100010",
  3011=>"000100100",
  3012=>"100110111",
  3013=>"011111110",
  3014=>"110001011",
  3015=>"001001101",
  3016=>"101000011",
  3017=>"000101100",
  3018=>"010010001",
  3019=>"001001111",
  3020=>"000010110",
  3021=>"000010111",
  3022=>"010100100",
  3023=>"110010100",
  3024=>"101010101",
  3025=>"111000100",
  3026=>"010110110",
  3027=>"010110000",
  3028=>"000111101",
  3029=>"011101010",
  3030=>"010001101",
  3031=>"111100011",
  3032=>"111010001",
  3033=>"000010101",
  3034=>"101001100",
  3035=>"101111010",
  3036=>"001000100",
  3037=>"011111110",
  3038=>"010000010",
  3039=>"001010011",
  3040=>"011111010",
  3041=>"000000100",
  3042=>"000000000",
  3043=>"110101101",
  3044=>"011101111",
  3045=>"101000101",
  3046=>"000111111",
  3047=>"001000011",
  3048=>"010000000",
  3049=>"110100110",
  3050=>"001011100",
  3051=>"110101010",
  3052=>"101100111",
  3053=>"101011011",
  3054=>"001010011",
  3055=>"001111101",
  3056=>"111011001",
  3057=>"100101011",
  3058=>"001011101",
  3059=>"111111001",
  3060=>"001111011",
  3061=>"110100101",
  3062=>"000011100",
  3063=>"100101110",
  3064=>"011111111",
  3065=>"011100000",
  3066=>"110000100",
  3067=>"110010001",
  3068=>"101101001",
  3069=>"000000000",
  3070=>"111110010",
  3071=>"011110100",
  3072=>"111110101",
  3073=>"100010111",
  3074=>"011011010",
  3075=>"001100010",
  3076=>"101011100",
  3077=>"100100011",
  3078=>"101010100",
  3079=>"001000100",
  3080=>"110010001",
  3081=>"000001000",
  3082=>"101100110",
  3083=>"110101001",
  3084=>"011100010",
  3085=>"111001000",
  3086=>"010111110",
  3087=>"011001001",
  3088=>"111110111",
  3089=>"010100101",
  3090=>"001100011",
  3091=>"101110011",
  3092=>"000000001",
  3093=>"111111100",
  3094=>"110000100",
  3095=>"000010001",
  3096=>"000000101",
  3097=>"111000011",
  3098=>"111110011",
  3099=>"110111110",
  3100=>"011111000",
  3101=>"100000000",
  3102=>"001000000",
  3103=>"100000101",
  3104=>"111000011",
  3105=>"001100111",
  3106=>"011011110",
  3107=>"110111101",
  3108=>"011111101",
  3109=>"101100011",
  3110=>"001000100",
  3111=>"111001101",
  3112=>"011010100",
  3113=>"100010001",
  3114=>"011111111",
  3115=>"001000000",
  3116=>"000000000",
  3117=>"010111111",
  3118=>"011110101",
  3119=>"100111001",
  3120=>"111100000",
  3121=>"010010010",
  3122=>"100001101",
  3123=>"001011111",
  3124=>"111110100",
  3125=>"100100011",
  3126=>"101011111",
  3127=>"001000100",
  3128=>"000101101",
  3129=>"010101010",
  3130=>"010010111",
  3131=>"010001010",
  3132=>"010000011",
  3133=>"000111101",
  3134=>"001011011",
  3135=>"000011110",
  3136=>"100011101",
  3137=>"101000011",
  3138=>"101001001",
  3139=>"100001010",
  3140=>"011100101",
  3141=>"111101111",
  3142=>"100001001",
  3143=>"110011010",
  3144=>"000101000",
  3145=>"110001101",
  3146=>"101001111",
  3147=>"010001110",
  3148=>"101110000",
  3149=>"111110001",
  3150=>"110010110",
  3151=>"111101001",
  3152=>"001110100",
  3153=>"100110001",
  3154=>"011100001",
  3155=>"101010011",
  3156=>"101101011",
  3157=>"010000001",
  3158=>"001000010",
  3159=>"001100000",
  3160=>"100111110",
  3161=>"100111011",
  3162=>"110111111",
  3163=>"111000001",
  3164=>"001111110",
  3165=>"010110101",
  3166=>"011011010",
  3167=>"100010000",
  3168=>"010101101",
  3169=>"111100110",
  3170=>"001010000",
  3171=>"001001011",
  3172=>"011111000",
  3173=>"110100000",
  3174=>"100001000",
  3175=>"110111110",
  3176=>"010100100",
  3177=>"011010010",
  3178=>"101110100",
  3179=>"111100011",
  3180=>"000011111",
  3181=>"100010010",
  3182=>"111101011",
  3183=>"010010001",
  3184=>"011110000",
  3185=>"100111100",
  3186=>"001011111",
  3187=>"001101110",
  3188=>"000111010",
  3189=>"000011111",
  3190=>"010111111",
  3191=>"001011101",
  3192=>"010011010",
  3193=>"010111001",
  3194=>"111010101",
  3195=>"110001101",
  3196=>"010000011",
  3197=>"111001000",
  3198=>"000110010",
  3199=>"001111011",
  3200=>"100010001",
  3201=>"110010110",
  3202=>"110100011",
  3203=>"110111111",
  3204=>"000111111",
  3205=>"000001000",
  3206=>"111100000",
  3207=>"011100010",
  3208=>"101000111",
  3209=>"001010010",
  3210=>"010110000",
  3211=>"101100101",
  3212=>"010110100",
  3213=>"011011010",
  3214=>"011110101",
  3215=>"111101111",
  3216=>"111010010",
  3217=>"101011100",
  3218=>"011111100",
  3219=>"010111100",
  3220=>"110011110",
  3221=>"010011001",
  3222=>"000000100",
  3223=>"011110001",
  3224=>"111100110",
  3225=>"111001100",
  3226=>"110110010",
  3227=>"010001100",
  3228=>"011001100",
  3229=>"100100100",
  3230=>"010001000",
  3231=>"000000011",
  3232=>"101101100",
  3233=>"101000001",
  3234=>"000000101",
  3235=>"100100101",
  3236=>"010000101",
  3237=>"010111110",
  3238=>"111100100",
  3239=>"000001100",
  3240=>"001010110",
  3241=>"110011110",
  3242=>"110011100",
  3243=>"101111110",
  3244=>"010000000",
  3245=>"101011010",
  3246=>"000010011",
  3247=>"100101000",
  3248=>"011111111",
  3249=>"011010001",
  3250=>"111001101",
  3251=>"101111010",
  3252=>"001010001",
  3253=>"001000001",
  3254=>"000111110",
  3255=>"011000000",
  3256=>"100011000",
  3257=>"111101111",
  3258=>"010000010",
  3259=>"111000110",
  3260=>"100100000",
  3261=>"010110000",
  3262=>"011110001",
  3263=>"101001100",
  3264=>"000110100",
  3265=>"100111101",
  3266=>"111110001",
  3267=>"011111101",
  3268=>"101110110",
  3269=>"100000000",
  3270=>"000110000",
  3271=>"010000100",
  3272=>"000011100",
  3273=>"010011011",
  3274=>"101111010",
  3275=>"110100000",
  3276=>"111010101",
  3277=>"111001011",
  3278=>"111101001",
  3279=>"100000101",
  3280=>"101110101",
  3281=>"000000100",
  3282=>"001001100",
  3283=>"101101010",
  3284=>"101011101",
  3285=>"101110000",
  3286=>"110011111",
  3287=>"001110000",
  3288=>"100100110",
  3289=>"100101001",
  3290=>"000000100",
  3291=>"000000011",
  3292=>"100111110",
  3293=>"111010110",
  3294=>"100111011",
  3295=>"110110110",
  3296=>"101010101",
  3297=>"011110001",
  3298=>"100100011",
  3299=>"110110000",
  3300=>"100101010",
  3301=>"110011011",
  3302=>"111100111",
  3303=>"000010111",
  3304=>"111001001",
  3305=>"010001100",
  3306=>"001101111",
  3307=>"000000011",
  3308=>"000110011",
  3309=>"110010101",
  3310=>"100111101",
  3311=>"111010111",
  3312=>"000000000",
  3313=>"010000000",
  3314=>"100110010",
  3315=>"010010110",
  3316=>"100010000",
  3317=>"100000010",
  3318=>"101100111",
  3319=>"101001001",
  3320=>"100111011",
  3321=>"101111001",
  3322=>"100101001",
  3323=>"010110100",
  3324=>"010000100",
  3325=>"000000110",
  3326=>"101001111",
  3327=>"010011110",
  3328=>"010110100",
  3329=>"110110100",
  3330=>"111010101",
  3331=>"010011011",
  3332=>"010111001",
  3333=>"011001000",
  3334=>"101101000",
  3335=>"011011011",
  3336=>"010101100",
  3337=>"111011011",
  3338=>"111010010",
  3339=>"010011000",
  3340=>"001011111",
  3341=>"010110001",
  3342=>"111110111",
  3343=>"110000001",
  3344=>"000110000",
  3345=>"010001111",
  3346=>"111001000",
  3347=>"111010101",
  3348=>"010011111",
  3349=>"001000111",
  3350=>"110001000",
  3351=>"001011010",
  3352=>"100101001",
  3353=>"100001111",
  3354=>"010000001",
  3355=>"001100101",
  3356=>"101000001",
  3357=>"010111001",
  3358=>"111100111",
  3359=>"101001100",
  3360=>"110000011",
  3361=>"000110010",
  3362=>"101010111",
  3363=>"101111000",
  3364=>"011011101",
  3365=>"010010010",
  3366=>"011111111",
  3367=>"000011101",
  3368=>"110011101",
  3369=>"101110110",
  3370=>"111100101",
  3371=>"111001010",
  3372=>"001010110",
  3373=>"111100000",
  3374=>"000000001",
  3375=>"111001011",
  3376=>"011000001",
  3377=>"111110011",
  3378=>"111100011",
  3379=>"010100111",
  3380=>"110110101",
  3381=>"100011000",
  3382=>"010110010",
  3383=>"011011011",
  3384=>"001110000",
  3385=>"101000011",
  3386=>"001111110",
  3387=>"001001011",
  3388=>"110111011",
  3389=>"001011100",
  3390=>"011100101",
  3391=>"010100100",
  3392=>"100010001",
  3393=>"000101010",
  3394=>"101010100",
  3395=>"111010000",
  3396=>"110010101",
  3397=>"111101111",
  3398=>"101001100",
  3399=>"001010100",
  3400=>"001110010",
  3401=>"001000000",
  3402=>"100001101",
  3403=>"010010000",
  3404=>"011100100",
  3405=>"110001101",
  3406=>"100001111",
  3407=>"001001000",
  3408=>"000010000",
  3409=>"111011100",
  3410=>"110100111",
  3411=>"111110101",
  3412=>"010100111",
  3413=>"100111101",
  3414=>"011111111",
  3415=>"110101000",
  3416=>"000010000",
  3417=>"000010011",
  3418=>"010010011",
  3419=>"010000000",
  3420=>"111111010",
  3421=>"000000111",
  3422=>"111111101",
  3423=>"000101000",
  3424=>"101011111",
  3425=>"111011001",
  3426=>"101000001",
  3427=>"001000011",
  3428=>"100110101",
  3429=>"000011001",
  3430=>"011010101",
  3431=>"100111110",
  3432=>"100101011",
  3433=>"011101100",
  3434=>"110111100",
  3435=>"001011110",
  3436=>"010101101",
  3437=>"011011101",
  3438=>"100010110",
  3439=>"111111111",
  3440=>"101001000",
  3441=>"011000011",
  3442=>"101110111",
  3443=>"010001000",
  3444=>"000110101",
  3445=>"100111111",
  3446=>"100110001",
  3447=>"111010000",
  3448=>"110000000",
  3449=>"100100010",
  3450=>"010110011",
  3451=>"011101001",
  3452=>"110000000",
  3453=>"101001000",
  3454=>"101011001",
  3455=>"110111101",
  3456=>"001100101",
  3457=>"001000010",
  3458=>"101101010",
  3459=>"000010101",
  3460=>"001110001",
  3461=>"110111100",
  3462=>"010111111",
  3463=>"111010101",
  3464=>"000110001",
  3465=>"100101110",
  3466=>"111000110",
  3467=>"000010010",
  3468=>"001111011",
  3469=>"001101001",
  3470=>"111100000",
  3471=>"010100101",
  3472=>"100011001",
  3473=>"111111011",
  3474=>"000111101",
  3475=>"001110001",
  3476=>"000101111",
  3477=>"000010011",
  3478=>"110110110",
  3479=>"000101111",
  3480=>"111010010",
  3481=>"001000010",
  3482=>"110010010",
  3483=>"000011010",
  3484=>"000101011",
  3485=>"110100100",
  3486=>"000010000",
  3487=>"000110001",
  3488=>"010100101",
  3489=>"000101000",
  3490=>"101000100",
  3491=>"010110110",
  3492=>"000111010",
  3493=>"001111000",
  3494=>"110110001",
  3495=>"011011011",
  3496=>"110011000",
  3497=>"011001101",
  3498=>"000001000",
  3499=>"101010110",
  3500=>"010110001",
  3501=>"111101111",
  3502=>"011101110",
  3503=>"011011111",
  3504=>"101001100",
  3505=>"101000001",
  3506=>"110111101",
  3507=>"111011000",
  3508=>"001011010",
  3509=>"001100000",
  3510=>"010101010",
  3511=>"101111010",
  3512=>"011000100",
  3513=>"000000000",
  3514=>"000101010",
  3515=>"110100111",
  3516=>"101001000",
  3517=>"011010000",
  3518=>"010110100",
  3519=>"101010111",
  3520=>"111010110",
  3521=>"111011000",
  3522=>"011111001",
  3523=>"001000100",
  3524=>"011110110",
  3525=>"010100010",
  3526=>"110000010",
  3527=>"011100011",
  3528=>"110110010",
  3529=>"010010001",
  3530=>"000010100",
  3531=>"011010010",
  3532=>"010011100",
  3533=>"011100001",
  3534=>"000000000",
  3535=>"011001001",
  3536=>"001111111",
  3537=>"111111000",
  3538=>"001000001",
  3539=>"111111000",
  3540=>"110110111",
  3541=>"010101011",
  3542=>"011110100",
  3543=>"011011101",
  3544=>"111100110",
  3545=>"011001011",
  3546=>"111010001",
  3547=>"110110010",
  3548=>"000101110",
  3549=>"001011010",
  3550=>"110110000",
  3551=>"001111000",
  3552=>"010001010",
  3553=>"101010101",
  3554=>"100001110",
  3555=>"010100101",
  3556=>"110000000",
  3557=>"000001011",
  3558=>"100110100",
  3559=>"000111001",
  3560=>"101101000",
  3561=>"011101100",
  3562=>"011011110",
  3563=>"101011011",
  3564=>"110111010",
  3565=>"100010100",
  3566=>"010000110",
  3567=>"011001111",
  3568=>"010011110",
  3569=>"110000011",
  3570=>"000111111",
  3571=>"111110000",
  3572=>"100000101",
  3573=>"110110100",
  3574=>"011000000",
  3575=>"001001110",
  3576=>"010111110",
  3577=>"011001011",
  3578=>"000100111",
  3579=>"110111011",
  3580=>"101000001",
  3581=>"111101101",
  3582=>"000110011",
  3583=>"000000111",
  3584=>"000100101",
  3585=>"011001111",
  3586=>"110101001",
  3587=>"111000100",
  3588=>"110010010",
  3589=>"100000110",
  3590=>"010100110",
  3591=>"010101011",
  3592=>"011110000",
  3593=>"100000110",
  3594=>"100011010",
  3595=>"000100000",
  3596=>"011101111",
  3597=>"001001101",
  3598=>"101000100",
  3599=>"011001100",
  3600=>"101000010",
  3601=>"011011100",
  3602=>"110110001",
  3603=>"001011001",
  3604=>"001110011",
  3605=>"000111001",
  3606=>"000110011",
  3607=>"001110001",
  3608=>"101101101",
  3609=>"101000000",
  3610=>"000000001",
  3611=>"010001111",
  3612=>"010000001",
  3613=>"111100110",
  3614=>"111001101",
  3615=>"011000000",
  3616=>"001101100",
  3617=>"101010110",
  3618=>"001011011",
  3619=>"010101101",
  3620=>"010000010",
  3621=>"111010101",
  3622=>"001011011",
  3623=>"011100011",
  3624=>"100111111",
  3625=>"111100000",
  3626=>"110111111",
  3627=>"111001110",
  3628=>"100001011",
  3629=>"110011011",
  3630=>"100100001",
  3631=>"001100100",
  3632=>"101011010",
  3633=>"000111011",
  3634=>"100001111",
  3635=>"111001010",
  3636=>"100000000",
  3637=>"111100011",
  3638=>"100100011",
  3639=>"110010111",
  3640=>"110111100",
  3641=>"111100001",
  3642=>"010110001",
  3643=>"111000000",
  3644=>"010101100",
  3645=>"101111010",
  3646=>"000110010",
  3647=>"000110011",
  3648=>"001111000",
  3649=>"100010111",
  3650=>"111010101",
  3651=>"001101100",
  3652=>"001100011",
  3653=>"010000011",
  3654=>"010011110",
  3655=>"011000111",
  3656=>"000000111",
  3657=>"011100101",
  3658=>"111110100",
  3659=>"100001010",
  3660=>"010011110",
  3661=>"010101000",
  3662=>"100000110",
  3663=>"011000000",
  3664=>"101100101",
  3665=>"000100010",
  3666=>"011111101",
  3667=>"100101001",
  3668=>"101011100",
  3669=>"110100101",
  3670=>"010110000",
  3671=>"001111100",
  3672=>"011110011",
  3673=>"011011100",
  3674=>"011010010",
  3675=>"110100101",
  3676=>"000101100",
  3677=>"111101110",
  3678=>"000111010",
  3679=>"000010111",
  3680=>"100011110",
  3681=>"011110010",
  3682=>"111001010",
  3683=>"001110010",
  3684=>"110010001",
  3685=>"011001001",
  3686=>"000111011",
  3687=>"110110010",
  3688=>"001100010",
  3689=>"001001001",
  3690=>"001010110",
  3691=>"011110111",
  3692=>"000100001",
  3693=>"000010111",
  3694=>"111111101",
  3695=>"100010101",
  3696=>"010100101",
  3697=>"111100001",
  3698=>"011100011",
  3699=>"000010000",
  3700=>"010011100",
  3701=>"010110010",
  3702=>"011001100",
  3703=>"010000100",
  3704=>"101000110",
  3705=>"000010000",
  3706=>"101100111",
  3707=>"000010101",
  3708=>"011000011",
  3709=>"010100110",
  3710=>"011111101",
  3711=>"001000100",
  3712=>"111101101",
  3713=>"111001111",
  3714=>"111000001",
  3715=>"110110100",
  3716=>"001000010",
  3717=>"000011100",
  3718=>"110011111",
  3719=>"110110100",
  3720=>"110011111",
  3721=>"000000001",
  3722=>"000011011",
  3723=>"000011001",
  3724=>"000010000",
  3725=>"011000111",
  3726=>"000000000",
  3727=>"110101001",
  3728=>"110110111",
  3729=>"000110000",
  3730=>"111001011",
  3731=>"010001000",
  3732=>"000001110",
  3733=>"100011111",
  3734=>"101010011",
  3735=>"011001010",
  3736=>"000100000",
  3737=>"100110001",
  3738=>"111111100",
  3739=>"111100110",
  3740=>"101001011",
  3741=>"110111001",
  3742=>"001101011",
  3743=>"101100100",
  3744=>"000011000",
  3745=>"100001001",
  3746=>"011011011",
  3747=>"010001101",
  3748=>"000001010",
  3749=>"100001100",
  3750=>"110010110",
  3751=>"000101000",
  3752=>"101100010",
  3753=>"110101010",
  3754=>"010111110",
  3755=>"101110110",
  3756=>"111001100",
  3757=>"011100010",
  3758=>"111000011",
  3759=>"100110001",
  3760=>"110110110",
  3761=>"011111011",
  3762=>"000111010",
  3763=>"101000100",
  3764=>"001110101",
  3765=>"001011110",
  3766=>"001001010",
  3767=>"000011011",
  3768=>"001000000",
  3769=>"110110011",
  3770=>"010110100",
  3771=>"100010001",
  3772=>"100001001",
  3773=>"000001001",
  3774=>"100000000",
  3775=>"111011111",
  3776=>"100111111",
  3777=>"100110110",
  3778=>"001101010",
  3779=>"010110011",
  3780=>"011101011",
  3781=>"000010000",
  3782=>"110010110",
  3783=>"001000101",
  3784=>"000011100",
  3785=>"111010010",
  3786=>"111011110",
  3787=>"000111010",
  3788=>"000000000",
  3789=>"111110111",
  3790=>"010101100",
  3791=>"001100000",
  3792=>"000101010",
  3793=>"010101001",
  3794=>"110110110",
  3795=>"010101100",
  3796=>"100011011",
  3797=>"110011001",
  3798=>"100100010",
  3799=>"010001011",
  3800=>"000000010",
  3801=>"001001001",
  3802=>"111111011",
  3803=>"001101010",
  3804=>"000011111",
  3805=>"100011000",
  3806=>"010001111",
  3807=>"011011110",
  3808=>"010000100",
  3809=>"010110010",
  3810=>"100011100",
  3811=>"100111000",
  3812=>"010100101",
  3813=>"001011001",
  3814=>"001010111",
  3815=>"011100011",
  3816=>"011010111",
  3817=>"101001011",
  3818=>"000110000",
  3819=>"011110111",
  3820=>"001001000",
  3821=>"001101011",
  3822=>"011010110",
  3823=>"001011101",
  3824=>"110111110",
  3825=>"110010010",
  3826=>"010000100",
  3827=>"000011110",
  3828=>"011000110",
  3829=>"010111111",
  3830=>"000010010",
  3831=>"100001110",
  3832=>"110110101",
  3833=>"100101111",
  3834=>"011100111",
  3835=>"011110000",
  3836=>"100001101",
  3837=>"010001110",
  3838=>"001010100",
  3839=>"000011101",
  3840=>"011001100",
  3841=>"011101110",
  3842=>"100001001",
  3843=>"111101001",
  3844=>"001011010",
  3845=>"110111010",
  3846=>"101110111",
  3847=>"000001011",
  3848=>"001110111",
  3849=>"110110100",
  3850=>"011001011",
  3851=>"100011011",
  3852=>"011100111",
  3853=>"010011100",
  3854=>"101100111",
  3855=>"111111111",
  3856=>"010101100",
  3857=>"101000010",
  3858=>"001101101",
  3859=>"110011011",
  3860=>"010111010",
  3861=>"011111111",
  3862=>"101001011",
  3863=>"100001110",
  3864=>"001011011",
  3865=>"000101100",
  3866=>"111111101",
  3867=>"011100101",
  3868=>"011011110",
  3869=>"001011000",
  3870=>"100110100",
  3871=>"001110000",
  3872=>"101010101",
  3873=>"000000010",
  3874=>"001110000",
  3875=>"100111010",
  3876=>"101010101",
  3877=>"010010110",
  3878=>"000001011",
  3879=>"100011000",
  3880=>"111110001",
  3881=>"111101101",
  3882=>"000110100",
  3883=>"101011110",
  3884=>"110110010",
  3885=>"000100000",
  3886=>"100010110",
  3887=>"000010001",
  3888=>"111100001",
  3889=>"100010110",
  3890=>"010100110",
  3891=>"001100101",
  3892=>"001011011",
  3893=>"101110111",
  3894=>"001010001",
  3895=>"110001010",
  3896=>"000110111",
  3897=>"100110110",
  3898=>"001101000",
  3899=>"000100001",
  3900=>"110010110",
  3901=>"001000011",
  3902=>"101000010",
  3903=>"100100001",
  3904=>"110101111",
  3905=>"111110010",
  3906=>"000100011",
  3907=>"001011010",
  3908=>"101101110",
  3909=>"100110001",
  3910=>"110100110",
  3911=>"111010000",
  3912=>"100100101",
  3913=>"010111011",
  3914=>"000000000",
  3915=>"111100100",
  3916=>"011001011",
  3917=>"010101010",
  3918=>"100000000",
  3919=>"111110110",
  3920=>"010110001",
  3921=>"110100111",
  3922=>"100011111",
  3923=>"100110011",
  3924=>"010010111",
  3925=>"100111110",
  3926=>"101110011",
  3927=>"011000011",
  3928=>"111101011",
  3929=>"011010001",
  3930=>"011001100",
  3931=>"111101001",
  3932=>"011110001",
  3933=>"100111100",
  3934=>"110110011",
  3935=>"011010010",
  3936=>"000101111",
  3937=>"001001110",
  3938=>"010101011",
  3939=>"000010100",
  3940=>"000011000",
  3941=>"101101110",
  3942=>"110110010",
  3943=>"010000001",
  3944=>"101100010",
  3945=>"010101111",
  3946=>"101100010",
  3947=>"011010011",
  3948=>"010100100",
  3949=>"100001011",
  3950=>"001100010",
  3951=>"011101011",
  3952=>"010110101",
  3953=>"101000101",
  3954=>"111110011",
  3955=>"000001111",
  3956=>"000000001",
  3957=>"111110100",
  3958=>"010100010",
  3959=>"001110000",
  3960=>"001010000",
  3961=>"110100010",
  3962=>"010111010",
  3963=>"110111011",
  3964=>"111101001",
  3965=>"000110010",
  3966=>"100100011",
  3967=>"110001111",
  3968=>"000000100",
  3969=>"001001001",
  3970=>"110000010",
  3971=>"010110001",
  3972=>"011010001",
  3973=>"100001010",
  3974=>"000011101",
  3975=>"101010000",
  3976=>"100111110",
  3977=>"110010001",
  3978=>"110001010",
  3979=>"100010000",
  3980=>"010001111",
  3981=>"111111100",
  3982=>"111110001",
  3983=>"111011000",
  3984=>"111011100",
  3985=>"101110111",
  3986=>"000010101",
  3987=>"110001110",
  3988=>"011101011",
  3989=>"001011001",
  3990=>"001011000",
  3991=>"001111001",
  3992=>"000111010",
  3993=>"001001111",
  3994=>"001101110",
  3995=>"000001000",
  3996=>"110110011",
  3997=>"000101011",
  3998=>"001010110",
  3999=>"101011011",
  4000=>"000000001",
  4001=>"001110101",
  4002=>"101010010",
  4003=>"101001100",
  4004=>"100001100",
  4005=>"010110100",
  4006=>"000001110",
  4007=>"111000010",
  4008=>"010010110",
  4009=>"100001010",
  4010=>"010001111",
  4011=>"101100011",
  4012=>"010101100",
  4013=>"111100111",
  4014=>"100010000",
  4015=>"011001111",
  4016=>"110110000",
  4017=>"001001011",
  4018=>"010100100",
  4019=>"000011000",
  4020=>"001100000",
  4021=>"001110011",
  4022=>"000100110",
  4023=>"010100101",
  4024=>"111110010",
  4025=>"101001010",
  4026=>"111111010",
  4027=>"100001001",
  4028=>"010100110",
  4029=>"101100110",
  4030=>"101110010",
  4031=>"011000001",
  4032=>"011010011",
  4033=>"000011010",
  4034=>"011110111",
  4035=>"000000001",
  4036=>"000110100",
  4037=>"010110010",
  4038=>"101110100",
  4039=>"111011010",
  4040=>"100101000",
  4041=>"000010100",
  4042=>"101010000",
  4043=>"101000001",
  4044=>"001101101",
  4045=>"000000000",
  4046=>"100100000",
  4047=>"101101111",
  4048=>"010010110",
  4049=>"100000100",
  4050=>"010000011",
  4051=>"111011110",
  4052=>"101100001",
  4053=>"000100111",
  4054=>"111011101",
  4055=>"000000000",
  4056=>"111100010",
  4057=>"000100011",
  4058=>"111110000",
  4059=>"111001001",
  4060=>"000111111",
  4061=>"010000000",
  4062=>"100011000",
  4063=>"100101110",
  4064=>"011111010",
  4065=>"101011111",
  4066=>"111100001",
  4067=>"000000001",
  4068=>"011001111",
  4069=>"101100000",
  4070=>"000100010",
  4071=>"001000001",
  4072=>"010000010",
  4073=>"110001010",
  4074=>"011000101",
  4075=>"111101010",
  4076=>"100101001",
  4077=>"111101101",
  4078=>"100110010",
  4079=>"000111011",
  4080=>"000011011",
  4081=>"111101101",
  4082=>"100010000",
  4083=>"000000000",
  4084=>"110001101",
  4085=>"011010101",
  4086=>"111111111",
  4087=>"000100101",
  4088=>"101011101",
  4089=>"110101001",
  4090=>"101100110",
  4091=>"000011110",
  4092=>"110110111",
  4093=>"111011000",
  4094=>"001000101",
  4095=>"101101010",
  4096=>"001001010",
  4097=>"001010100",
  4098=>"101111000",
  4099=>"111011111",
  4100=>"101000101",
  4101=>"100011110",
  4102=>"100110101",
  4103=>"011001000",
  4104=>"110101101",
  4105=>"010000100",
  4106=>"010100101",
  4107=>"111101010",
  4108=>"101111111",
  4109=>"011011111",
  4110=>"100110011",
  4111=>"101101010",
  4112=>"101100111",
  4113=>"000001100",
  4114=>"000010000",
  4115=>"001110101",
  4116=>"010101001",
  4117=>"100000110",
  4118=>"110001100",
  4119=>"011001110",
  4120=>"001011000",
  4121=>"010111010",
  4122=>"110111111",
  4123=>"000000110",
  4124=>"010110101",
  4125=>"100101011",
  4126=>"100001100",
  4127=>"001101000",
  4128=>"011000001",
  4129=>"010110001",
  4130=>"110000001",
  4131=>"101111010",
  4132=>"000100001",
  4133=>"111011111",
  4134=>"011110001",
  4135=>"111111110",
  4136=>"101110000",
  4137=>"000110100",
  4138=>"110111011",
  4139=>"011011100",
  4140=>"101101110",
  4141=>"011010101",
  4142=>"000000111",
  4143=>"111011101",
  4144=>"100000111",
  4145=>"001100001",
  4146=>"001011110",
  4147=>"011100000",
  4148=>"010100111",
  4149=>"010100101",
  4150=>"001110101",
  4151=>"111011011",
  4152=>"001101101",
  4153=>"001010100",
  4154=>"011110110",
  4155=>"011101010",
  4156=>"010011010",
  4157=>"010100000",
  4158=>"111110001",
  4159=>"111101010",
  4160=>"110101011",
  4161=>"000000001",
  4162=>"111100110",
  4163=>"111010000",
  4164=>"000010001",
  4165=>"001000101",
  4166=>"011111000",
  4167=>"000011100",
  4168=>"011010001",
  4169=>"110001000",
  4170=>"101010000",
  4171=>"000111111",
  4172=>"000000100",
  4173=>"111000010",
  4174=>"100100100",
  4175=>"011011100",
  4176=>"011110110",
  4177=>"101110100",
  4178=>"001111010",
  4179=>"011001000",
  4180=>"000100101",
  4181=>"100010010",
  4182=>"100001110",
  4183=>"010010011",
  4184=>"110000111",
  4185=>"111010010",
  4186=>"000010100",
  4187=>"111101010",
  4188=>"111111110",
  4189=>"011100010",
  4190=>"000101110",
  4191=>"001000011",
  4192=>"000110111",
  4193=>"111000000",
  4194=>"010000011",
  4195=>"001010101",
  4196=>"001111011",
  4197=>"000100110",
  4198=>"100111001",
  4199=>"000000110",
  4200=>"000000111",
  4201=>"111011001",
  4202=>"000000111",
  4203=>"011011001",
  4204=>"111110011",
  4205=>"000101010",
  4206=>"010011111",
  4207=>"111111011",
  4208=>"110100111",
  4209=>"010000011",
  4210=>"101111101",
  4211=>"011100010",
  4212=>"001111010",
  4213=>"001001111",
  4214=>"101100001",
  4215=>"111100101",
  4216=>"001010100",
  4217=>"100001010",
  4218=>"000011101",
  4219=>"111111100",
  4220=>"011111111",
  4221=>"000101111",
  4222=>"100101101",
  4223=>"100000111",
  4224=>"010001100",
  4225=>"111011000",
  4226=>"010010000",
  4227=>"010101001",
  4228=>"101001001",
  4229=>"001101011",
  4230=>"011111010",
  4231=>"101100100",
  4232=>"100010011",
  4233=>"000000100",
  4234=>"101000000",
  4235=>"001101111",
  4236=>"100100001",
  4237=>"111111111",
  4238=>"011110000",
  4239=>"001001010",
  4240=>"011000011",
  4241=>"000011011",
  4242=>"111000000",
  4243=>"011001011",
  4244=>"010011111",
  4245=>"110001010",
  4246=>"011011001",
  4247=>"010100111",
  4248=>"001111011",
  4249=>"110010101",
  4250=>"000011101",
  4251=>"010001100",
  4252=>"000000000",
  4253=>"100111010",
  4254=>"100000100",
  4255=>"001110101",
  4256=>"110011010",
  4257=>"111010101",
  4258=>"110100000",
  4259=>"110010010",
  4260=>"110110011",
  4261=>"101001011",
  4262=>"100110011",
  4263=>"101111100",
  4264=>"110001010",
  4265=>"111000101",
  4266=>"001011000",
  4267=>"001010101",
  4268=>"100110101",
  4269=>"001000101",
  4270=>"101100011",
  4271=>"001110101",
  4272=>"010000100",
  4273=>"001101010",
  4274=>"001010100",
  4275=>"101101111",
  4276=>"100010011",
  4277=>"000010010",
  4278=>"111110101",
  4279=>"000001011",
  4280=>"010101001",
  4281=>"100010111",
  4282=>"100101101",
  4283=>"101111101",
  4284=>"001110001",
  4285=>"011011101",
  4286=>"110111010",
  4287=>"000111111",
  4288=>"111111010",
  4289=>"100100001",
  4290=>"110110000",
  4291=>"100110110",
  4292=>"001111110",
  4293=>"010010010",
  4294=>"101011011",
  4295=>"101011111",
  4296=>"000111111",
  4297=>"001010111",
  4298=>"111001111",
  4299=>"001110011",
  4300=>"000101111",
  4301=>"001010111",
  4302=>"011000101",
  4303=>"111101010",
  4304=>"011111101",
  4305=>"110100111",
  4306=>"001000110",
  4307=>"110111011",
  4308=>"001110001",
  4309=>"110000010",
  4310=>"010100100",
  4311=>"111011111",
  4312=>"000011010",
  4313=>"010111011",
  4314=>"000011101",
  4315=>"111001010",
  4316=>"010001101",
  4317=>"000101001",
  4318=>"101111011",
  4319=>"100100110",
  4320=>"101101101",
  4321=>"000010100",
  4322=>"000010111",
  4323=>"100001111",
  4324=>"100111110",
  4325=>"101110100",
  4326=>"001111111",
  4327=>"000101000",
  4328=>"010111111",
  4329=>"110010011",
  4330=>"111011111",
  4331=>"011011111",
  4332=>"110110111",
  4333=>"110100111",
  4334=>"010000010",
  4335=>"110000100",
  4336=>"110111000",
  4337=>"001000001",
  4338=>"100100001",
  4339=>"111001000",
  4340=>"001111010",
  4341=>"001010101",
  4342=>"110101100",
  4343=>"011110101",
  4344=>"110110110",
  4345=>"101110101",
  4346=>"100001101",
  4347=>"100011100",
  4348=>"001000111",
  4349=>"101101100",
  4350=>"100101100",
  4351=>"100000110",
  4352=>"100000010",
  4353=>"011110001",
  4354=>"010111110",
  4355=>"111110100",
  4356=>"110011100",
  4357=>"111001110",
  4358=>"110001000",
  4359=>"011111111",
  4360=>"000001100",
  4361=>"101111111",
  4362=>"100010001",
  4363=>"110001011",
  4364=>"000010001",
  4365=>"000011110",
  4366=>"110000111",
  4367=>"000011010",
  4368=>"001100000",
  4369=>"101001111",
  4370=>"101011000",
  4371=>"111010111",
  4372=>"011110100",
  4373=>"011010110",
  4374=>"100011111",
  4375=>"000111001",
  4376=>"110111010",
  4377=>"110101111",
  4378=>"100111100",
  4379=>"111101101",
  4380=>"110000000",
  4381=>"000100000",
  4382=>"111100001",
  4383=>"101011011",
  4384=>"001101000",
  4385=>"101000111",
  4386=>"011001100",
  4387=>"011101000",
  4388=>"011011010",
  4389=>"011101100",
  4390=>"001001100",
  4391=>"011110001",
  4392=>"101010011",
  4393=>"101011100",
  4394=>"010001010",
  4395=>"010011111",
  4396=>"010011111",
  4397=>"101111000",
  4398=>"110011100",
  4399=>"100000111",
  4400=>"000001100",
  4401=>"001110110",
  4402=>"100000111",
  4403=>"000000101",
  4404=>"001101110",
  4405=>"110111110",
  4406=>"001101100",
  4407=>"001111111",
  4408=>"000110011",
  4409=>"000111001",
  4410=>"100001110",
  4411=>"111001001",
  4412=>"010111000",
  4413=>"010001010",
  4414=>"001101001",
  4415=>"011100000",
  4416=>"101110010",
  4417=>"001000001",
  4418=>"010000001",
  4419=>"001000001",
  4420=>"101101101",
  4421=>"001101000",
  4422=>"010101010",
  4423=>"000010001",
  4424=>"000000101",
  4425=>"100111001",
  4426=>"110100000",
  4427=>"011000011",
  4428=>"101000010",
  4429=>"010110010",
  4430=>"111001001",
  4431=>"000101111",
  4432=>"011011110",
  4433=>"010001010",
  4434=>"010001000",
  4435=>"000100000",
  4436=>"001001110",
  4437=>"000001100",
  4438=>"110100111",
  4439=>"001000010",
  4440=>"011110100",
  4441=>"011111001",
  4442=>"011010001",
  4443=>"110111001",
  4444=>"101011110",
  4445=>"010000010",
  4446=>"101001111",
  4447=>"000010100",
  4448=>"011001100",
  4449=>"000000110",
  4450=>"000011110",
  4451=>"000000000",
  4452=>"001110110",
  4453=>"100001101",
  4454=>"001100010",
  4455=>"101101110",
  4456=>"100101111",
  4457=>"000110011",
  4458=>"000001101",
  4459=>"111010001",
  4460=>"100010010",
  4461=>"111000100",
  4462=>"000010111",
  4463=>"110011010",
  4464=>"001001011",
  4465=>"011001101",
  4466=>"101100011",
  4467=>"111010100",
  4468=>"111001011",
  4469=>"000101011",
  4470=>"110011011",
  4471=>"010000001",
  4472=>"010011110",
  4473=>"111001111",
  4474=>"111110111",
  4475=>"110001011",
  4476=>"010010001",
  4477=>"110100010",
  4478=>"001001011",
  4479=>"000000000",
  4480=>"100101010",
  4481=>"011001001",
  4482=>"111111011",
  4483=>"101011110",
  4484=>"001000001",
  4485=>"000000101",
  4486=>"110000000",
  4487=>"011000100",
  4488=>"111100001",
  4489=>"110001001",
  4490=>"000110111",
  4491=>"001010111",
  4492=>"000110010",
  4493=>"100101100",
  4494=>"010000001",
  4495=>"100110000",
  4496=>"001000110",
  4497=>"010110000",
  4498=>"111111011",
  4499=>"101101111",
  4500=>"111000010",
  4501=>"101001101",
  4502=>"000000011",
  4503=>"101101010",
  4504=>"110110111",
  4505=>"000000111",
  4506=>"010011110",
  4507=>"111100100",
  4508=>"001110101",
  4509=>"010011110",
  4510=>"011111000",
  4511=>"100001001",
  4512=>"110101101",
  4513=>"010000111",
  4514=>"000101001",
  4515=>"011101001",
  4516=>"100111000",
  4517=>"001110100",
  4518=>"101011011",
  4519=>"111101100",
  4520=>"100101111",
  4521=>"111010001",
  4522=>"000111010",
  4523=>"111011101",
  4524=>"100000010",
  4525=>"110111101",
  4526=>"100001000",
  4527=>"101010101",
  4528=>"010000011",
  4529=>"100100001",
  4530=>"010000011",
  4531=>"000011110",
  4532=>"110111101",
  4533=>"010101100",
  4534=>"011110111",
  4535=>"001111001",
  4536=>"100100100",
  4537=>"101100001",
  4538=>"110100101",
  4539=>"000000011",
  4540=>"001011101",
  4541=>"011111110",
  4542=>"101111010",
  4543=>"111100110",
  4544=>"110111001",
  4545=>"110110010",
  4546=>"010000001",
  4547=>"010011110",
  4548=>"000111100",
  4549=>"000010010",
  4550=>"000000011",
  4551=>"001101011",
  4552=>"001110001",
  4553=>"011000100",
  4554=>"010011110",
  4555=>"111001001",
  4556=>"111101011",
  4557=>"010100000",
  4558=>"010110110",
  4559=>"100011101",
  4560=>"011001111",
  4561=>"100111111",
  4562=>"111111010",
  4563=>"101100110",
  4564=>"010000100",
  4565=>"011011110",
  4566=>"011001101",
  4567=>"010101110",
  4568=>"001001000",
  4569=>"101101011",
  4570=>"000001100",
  4571=>"111011101",
  4572=>"001011110",
  4573=>"011000010",
  4574=>"100000100",
  4575=>"000100110",
  4576=>"111101000",
  4577=>"101100000",
  4578=>"001111000",
  4579=>"000110000",
  4580=>"000001110",
  4581=>"110010000",
  4582=>"111011110",
  4583=>"110010100",
  4584=>"011111110",
  4585=>"011110000",
  4586=>"010111010",
  4587=>"001011000",
  4588=>"110000000",
  4589=>"001111000",
  4590=>"100001101",
  4591=>"001001110",
  4592=>"010001110",
  4593=>"010000000",
  4594=>"100101110",
  4595=>"001000110",
  4596=>"111110100",
  4597=>"001001110",
  4598=>"100100111",
  4599=>"011000100",
  4600=>"110001011",
  4601=>"001100100",
  4602=>"010111110",
  4603=>"010110110",
  4604=>"001000010",
  4605=>"100010011",
  4606=>"000010001",
  4607=>"011111111",
  4608=>"000111011",
  4609=>"001000110",
  4610=>"000110111",
  4611=>"110011110",
  4612=>"110001011",
  4613=>"000111100",
  4614=>"101111110",
  4615=>"001100000",
  4616=>"111100011",
  4617=>"011111000",
  4618=>"100111111",
  4619=>"111010010",
  4620=>"000001100",
  4621=>"111100100",
  4622=>"010010100",
  4623=>"100010101",
  4624=>"000001100",
  4625=>"000010000",
  4626=>"110010100",
  4627=>"111111100",
  4628=>"110101011",
  4629=>"101001101",
  4630=>"011111000",
  4631=>"110010011",
  4632=>"010111111",
  4633=>"000101010",
  4634=>"010110000",
  4635=>"101000110",
  4636=>"010100100",
  4637=>"000110011",
  4638=>"100100001",
  4639=>"101100000",
  4640=>"101111111",
  4641=>"000001110",
  4642=>"101000000",
  4643=>"001101001",
  4644=>"011001111",
  4645=>"000111000",
  4646=>"100010111",
  4647=>"000001101",
  4648=>"010001101",
  4649=>"111100000",
  4650=>"010100011",
  4651=>"110101000",
  4652=>"011100101",
  4653=>"101001000",
  4654=>"000001001",
  4655=>"000100100",
  4656=>"110011111",
  4657=>"000110101",
  4658=>"101000001",
  4659=>"111001000",
  4660=>"001110101",
  4661=>"100110011",
  4662=>"111000111",
  4663=>"011111100",
  4664=>"111101101",
  4665=>"110101110",
  4666=>"111011000",
  4667=>"010111100",
  4668=>"001111011",
  4669=>"101011000",
  4670=>"111011100",
  4671=>"010101111",
  4672=>"000100100",
  4673=>"000010001",
  4674=>"100000100",
  4675=>"110000010",
  4676=>"110110000",
  4677=>"111110110",
  4678=>"101100000",
  4679=>"000101100",
  4680=>"011100011",
  4681=>"110001101",
  4682=>"110110001",
  4683=>"101010010",
  4684=>"100001100",
  4685=>"000011110",
  4686=>"010111000",
  4687=>"001011011",
  4688=>"010010000",
  4689=>"111100010",
  4690=>"000011011",
  4691=>"000101011",
  4692=>"100110110",
  4693=>"011110000",
  4694=>"100001101",
  4695=>"100001000",
  4696=>"111101111",
  4697=>"111010000",
  4698=>"000011110",
  4699=>"010110100",
  4700=>"000000101",
  4701=>"000001110",
  4702=>"110001000",
  4703=>"011110110",
  4704=>"110111000",
  4705=>"101100100",
  4706=>"000110111",
  4707=>"100001101",
  4708=>"101111011",
  4709=>"010011010",
  4710=>"010100010",
  4711=>"001110110",
  4712=>"001000010",
  4713=>"000001000",
  4714=>"101000001",
  4715=>"000011100",
  4716=>"011111100",
  4717=>"111110111",
  4718=>"101101110",
  4719=>"011110101",
  4720=>"011100111",
  4721=>"101001010",
  4722=>"111000111",
  4723=>"100010010",
  4724=>"100101011",
  4725=>"000000100",
  4726=>"011010000",
  4727=>"111000110",
  4728=>"000001111",
  4729=>"010110111",
  4730=>"100111100",
  4731=>"110000101",
  4732=>"110100100",
  4733=>"110110010",
  4734=>"000000010",
  4735=>"110000110",
  4736=>"011110110",
  4737=>"011000000",
  4738=>"110110011",
  4739=>"011000010",
  4740=>"111111011",
  4741=>"110000101",
  4742=>"011111111",
  4743=>"100101111",
  4744=>"101111100",
  4745=>"010111110",
  4746=>"111110111",
  4747=>"111101011",
  4748=>"011010010",
  4749=>"101001110",
  4750=>"000101111",
  4751=>"010110000",
  4752=>"001001110",
  4753=>"101110111",
  4754=>"000101001",
  4755=>"111100011",
  4756=>"010000000",
  4757=>"110000100",
  4758=>"011001111",
  4759=>"010001010",
  4760=>"011110110",
  4761=>"100011111",
  4762=>"110000000",
  4763=>"110010111",
  4764=>"100001100",
  4765=>"100011111",
  4766=>"101011101",
  4767=>"110010100",
  4768=>"110000000",
  4769=>"100110100",
  4770=>"010110010",
  4771=>"000000000",
  4772=>"111111101",
  4773=>"011011100",
  4774=>"101111011",
  4775=>"011000101",
  4776=>"101001011",
  4777=>"110100101",
  4778=>"001001110",
  4779=>"011001110",
  4780=>"001000010",
  4781=>"010011110",
  4782=>"011000000",
  4783=>"011000010",
  4784=>"011101000",
  4785=>"000010110",
  4786=>"101011101",
  4787=>"100010010",
  4788=>"111011010",
  4789=>"000001101",
  4790=>"110110111",
  4791=>"110000110",
  4792=>"111010111",
  4793=>"100010000",
  4794=>"111111011",
  4795=>"000010001",
  4796=>"001000000",
  4797=>"010011000",
  4798=>"000011000",
  4799=>"111100000",
  4800=>"111111100",
  4801=>"000110011",
  4802=>"110100010",
  4803=>"100110100",
  4804=>"010100110",
  4805=>"001100111",
  4806=>"110000101",
  4807=>"010000010",
  4808=>"010001000",
  4809=>"000101010",
  4810=>"000010111",
  4811=>"111011010",
  4812=>"111110101",
  4813=>"100110000",
  4814=>"101011010",
  4815=>"110100111",
  4816=>"101000001",
  4817=>"101110101",
  4818=>"000101100",
  4819=>"110011010",
  4820=>"000001000",
  4821=>"011100010",
  4822=>"111010010",
  4823=>"111100000",
  4824=>"001111111",
  4825=>"111111011",
  4826=>"111111111",
  4827=>"110000100",
  4828=>"010010100",
  4829=>"010111101",
  4830=>"011010101",
  4831=>"100100001",
  4832=>"010110111",
  4833=>"001001101",
  4834=>"100100001",
  4835=>"001011001",
  4836=>"101010010",
  4837=>"011111000",
  4838=>"110111111",
  4839=>"111111011",
  4840=>"000000100",
  4841=>"101110011",
  4842=>"110100001",
  4843=>"110001100",
  4844=>"000111011",
  4845=>"010110111",
  4846=>"011011001",
  4847=>"000110100",
  4848=>"110001001",
  4849=>"100000001",
  4850=>"110100010",
  4851=>"010110111",
  4852=>"100110100",
  4853=>"100101110",
  4854=>"110001100",
  4855=>"111111101",
  4856=>"101001100",
  4857=>"111111111",
  4858=>"110100101",
  4859=>"110110001",
  4860=>"011001111",
  4861=>"000110110",
  4862=>"110100111",
  4863=>"010101100",
  4864=>"001111101",
  4865=>"010111000",
  4866=>"010000110",
  4867=>"000000000",
  4868=>"110001010",
  4869=>"010100100",
  4870=>"010001110",
  4871=>"010010010",
  4872=>"110111010",
  4873=>"010110011",
  4874=>"011111001",
  4875=>"000010111",
  4876=>"100110011",
  4877=>"011100110",
  4878=>"000001101",
  4879=>"110111000",
  4880=>"001010001",
  4881=>"001111110",
  4882=>"111000111",
  4883=>"011000011",
  4884=>"110101000",
  4885=>"001110010",
  4886=>"110110101",
  4887=>"100100010",
  4888=>"101111100",
  4889=>"010001010",
  4890=>"101001001",
  4891=>"000111011",
  4892=>"000001010",
  4893=>"001110111",
  4894=>"001001100",
  4895=>"000011101",
  4896=>"010001010",
  4897=>"100000011",
  4898=>"010100000",
  4899=>"110111001",
  4900=>"101011101",
  4901=>"000100010",
  4902=>"111110100",
  4903=>"111111011",
  4904=>"000101001",
  4905=>"000111000",
  4906=>"010101011",
  4907=>"000101001",
  4908=>"110000000",
  4909=>"010111100",
  4910=>"010010110",
  4911=>"111110111",
  4912=>"110110011",
  4913=>"010000101",
  4914=>"000110000",
  4915=>"111101011",
  4916=>"010010000",
  4917=>"101000110",
  4918=>"100011010",
  4919=>"101011111",
  4920=>"100010010",
  4921=>"010010111",
  4922=>"111011010",
  4923=>"101111111",
  4924=>"101110101",
  4925=>"000000100",
  4926=>"101100101",
  4927=>"110011000",
  4928=>"001000100",
  4929=>"000011011",
  4930=>"010010001",
  4931=>"000111011",
  4932=>"100010100",
  4933=>"000011111",
  4934=>"010011000",
  4935=>"001011110",
  4936=>"101010001",
  4937=>"011000001",
  4938=>"100101100",
  4939=>"011111010",
  4940=>"100000010",
  4941=>"110111111",
  4942=>"111110010",
  4943=>"110010100",
  4944=>"110011011",
  4945=>"010001000",
  4946=>"000001000",
  4947=>"010111110",
  4948=>"000111000",
  4949=>"111011000",
  4950=>"000110010",
  4951=>"011010111",
  4952=>"000101011",
  4953=>"011000111",
  4954=>"001010001",
  4955=>"010001101",
  4956=>"010110100",
  4957=>"000001010",
  4958=>"111100100",
  4959=>"000110011",
  4960=>"001111000",
  4961=>"000011000",
  4962=>"010101011",
  4963=>"110100011",
  4964=>"011110111",
  4965=>"001001101",
  4966=>"101111101",
  4967=>"000111100",
  4968=>"010101111",
  4969=>"111010100",
  4970=>"001000100",
  4971=>"000000101",
  4972=>"000000000",
  4973=>"111110001",
  4974=>"111001111",
  4975=>"110100011",
  4976=>"110001111",
  4977=>"101001001",
  4978=>"100110100",
  4979=>"001001101",
  4980=>"010011001",
  4981=>"011101100",
  4982=>"100001101",
  4983=>"100110111",
  4984=>"000100100",
  4985=>"010000101",
  4986=>"100110101",
  4987=>"101011011",
  4988=>"000000001",
  4989=>"000011000",
  4990=>"010000010",
  4991=>"001100110",
  4992=>"001100100",
  4993=>"010000001",
  4994=>"111100111",
  4995=>"100010100",
  4996=>"101111101",
  4997=>"000001101",
  4998=>"011111010",
  4999=>"110001000",
  5000=>"001100000",
  5001=>"000100011",
  5002=>"111010001",
  5003=>"000100000",
  5004=>"100000000",
  5005=>"000000101",
  5006=>"011011010",
  5007=>"001001101",
  5008=>"010111000",
  5009=>"110011111",
  5010=>"000010010",
  5011=>"010111111",
  5012=>"101111001",
  5013=>"010101101",
  5014=>"100110100",
  5015=>"101010000",
  5016=>"110010111",
  5017=>"101000001",
  5018=>"000101010",
  5019=>"110111001",
  5020=>"010110100",
  5021=>"101101110",
  5022=>"101010010",
  5023=>"100010011",
  5024=>"100110010",
  5025=>"010000000",
  5026=>"101000010",
  5027=>"101100111",
  5028=>"100011010",
  5029=>"110110011",
  5030=>"100010010",
  5031=>"000110000",
  5032=>"000001111",
  5033=>"100101100",
  5034=>"111010111",
  5035=>"000001110",
  5036=>"101010101",
  5037=>"011110101",
  5038=>"100100101",
  5039=>"000001001",
  5040=>"101101001",
  5041=>"011010101",
  5042=>"001000110",
  5043=>"101011000",
  5044=>"100010110",
  5045=>"110001000",
  5046=>"100100101",
  5047=>"011100010",
  5048=>"101111011",
  5049=>"101101000",
  5050=>"010101100",
  5051=>"000001011",
  5052=>"100101011",
  5053=>"010101010",
  5054=>"111111111",
  5055=>"001001011",
  5056=>"101011000",
  5057=>"001110001",
  5058=>"111010101",
  5059=>"111001010",
  5060=>"000011011",
  5061=>"111011110",
  5062=>"111000111",
  5063=>"110111101",
  5064=>"010110001",
  5065=>"000010001",
  5066=>"000010110",
  5067=>"101010100",
  5068=>"110110000",
  5069=>"101010100",
  5070=>"011100001",
  5071=>"001001111",
  5072=>"011010010",
  5073=>"000010001",
  5074=>"001100110",
  5075=>"010000011",
  5076=>"010101001",
  5077=>"001110001",
  5078=>"101010011",
  5079=>"111101101",
  5080=>"100100111",
  5081=>"100100011",
  5082=>"111011111",
  5083=>"111010111",
  5084=>"100101110",
  5085=>"111101101",
  5086=>"001011010",
  5087=>"000111001",
  5088=>"110010110",
  5089=>"000011010",
  5090=>"100000100",
  5091=>"000000001",
  5092=>"010110010",
  5093=>"010111110",
  5094=>"010011001",
  5095=>"110111111",
  5096=>"001101111",
  5097=>"011000100",
  5098=>"010101101",
  5099=>"100111001",
  5100=>"011001111",
  5101=>"001001001",
  5102=>"000111110",
  5103=>"001011110",
  5104=>"011010010",
  5105=>"101100000",
  5106=>"110001011",
  5107=>"010001100",
  5108=>"000101101",
  5109=>"101101110",
  5110=>"011110010",
  5111=>"011000111",
  5112=>"001001000",
  5113=>"001010010",
  5114=>"110011001",
  5115=>"011000100",
  5116=>"001011000",
  5117=>"001010100",
  5118=>"000000000",
  5119=>"101110001",
  5120=>"110000110",
  5121=>"000010000",
  5122=>"111001101",
  5123=>"001000001",
  5124=>"000011111",
  5125=>"110101000",
  5126=>"101001000",
  5127=>"101010001",
  5128=>"011111100",
  5129=>"101001101",
  5130=>"001100011",
  5131=>"100011001",
  5132=>"001100111",
  5133=>"111111001",
  5134=>"010011100",
  5135=>"101011001",
  5136=>"000100111",
  5137=>"000110001",
  5138=>"001010111",
  5139=>"111000101",
  5140=>"110011110",
  5141=>"100001000",
  5142=>"000000000",
  5143=>"011011010",
  5144=>"100001101",
  5145=>"011000110",
  5146=>"100100101",
  5147=>"111000000",
  5148=>"011110101",
  5149=>"110101000",
  5150=>"111100110",
  5151=>"101001101",
  5152=>"001011011",
  5153=>"111010001",
  5154=>"001110100",
  5155=>"101011111",
  5156=>"110100011",
  5157=>"110100110",
  5158=>"011101000",
  5159=>"011110111",
  5160=>"001001101",
  5161=>"101110101",
  5162=>"000000100",
  5163=>"001000100",
  5164=>"000101000",
  5165=>"010011001",
  5166=>"010000000",
  5167=>"010110010",
  5168=>"011100110",
  5169=>"000010000",
  5170=>"010100011",
  5171=>"101000111",
  5172=>"000111011",
  5173=>"101110011",
  5174=>"010001111",
  5175=>"000111100",
  5176=>"011101100",
  5177=>"011111000",
  5178=>"101100110",
  5179=>"000001010",
  5180=>"011100001",
  5181=>"100000110",
  5182=>"010011100",
  5183=>"001111011",
  5184=>"101100100",
  5185=>"011010000",
  5186=>"000001000",
  5187=>"000111111",
  5188=>"101001001",
  5189=>"001110011",
  5190=>"001100101",
  5191=>"011110000",
  5192=>"000111001",
  5193=>"000111101",
  5194=>"000101001",
  5195=>"011011100",
  5196=>"000011010",
  5197=>"111110101",
  5198=>"100111101",
  5199=>"100111011",
  5200=>"001100000",
  5201=>"011010111",
  5202=>"000110010",
  5203=>"101000000",
  5204=>"110110110",
  5205=>"101001001",
  5206=>"100100111",
  5207=>"111011111",
  5208=>"000100011",
  5209=>"000101111",
  5210=>"011111110",
  5211=>"000110111",
  5212=>"000101101",
  5213=>"011101100",
  5214=>"010001111",
  5215=>"010011011",
  5216=>"011011101",
  5217=>"100101111",
  5218=>"111010011",
  5219=>"100101000",
  5220=>"001011000",
  5221=>"100100000",
  5222=>"110100000",
  5223=>"111010010",
  5224=>"011010110",
  5225=>"110000000",
  5226=>"101100000",
  5227=>"101101010",
  5228=>"101111001",
  5229=>"000111101",
  5230=>"011010001",
  5231=>"001010110",
  5232=>"110010000",
  5233=>"101000011",
  5234=>"110111110",
  5235=>"111100110",
  5236=>"001001110",
  5237=>"000000001",
  5238=>"111011011",
  5239=>"000111010",
  5240=>"000100110",
  5241=>"010010111",
  5242=>"010101110",
  5243=>"001100111",
  5244=>"010010111",
  5245=>"111011010",
  5246=>"011010011",
  5247=>"010110100",
  5248=>"010101101",
  5249=>"000101111",
  5250=>"000010000",
  5251=>"000001100",
  5252=>"101011111",
  5253=>"110111011",
  5254=>"110101000",
  5255=>"111001111",
  5256=>"110001010",
  5257=>"100011100",
  5258=>"000000100",
  5259=>"100100100",
  5260=>"110110101",
  5261=>"110011000",
  5262=>"001000110",
  5263=>"101110010",
  5264=>"010011011",
  5265=>"000110011",
  5266=>"010101101",
  5267=>"000000001",
  5268=>"011101011",
  5269=>"011100110",
  5270=>"000101010",
  5271=>"011001001",
  5272=>"000110101",
  5273=>"100010010",
  5274=>"010000010",
  5275=>"110111010",
  5276=>"100111110",
  5277=>"100010000",
  5278=>"100101001",
  5279=>"101111011",
  5280=>"100011010",
  5281=>"001110111",
  5282=>"000111110",
  5283=>"000011010",
  5284=>"000101010",
  5285=>"110110110",
  5286=>"010100001",
  5287=>"011110111",
  5288=>"100011001",
  5289=>"110110111",
  5290=>"101100111",
  5291=>"110000101",
  5292=>"001001001",
  5293=>"000101011",
  5294=>"110000010",
  5295=>"111000000",
  5296=>"111011101",
  5297=>"011010001",
  5298=>"101000101",
  5299=>"101000100",
  5300=>"100000001",
  5301=>"001010000",
  5302=>"111010101",
  5303=>"001010000",
  5304=>"101010010",
  5305=>"100110111",
  5306=>"011111100",
  5307=>"111001010",
  5308=>"001011011",
  5309=>"100000001",
  5310=>"011101000",
  5311=>"101111011",
  5312=>"000010011",
  5313=>"001001011",
  5314=>"011011111",
  5315=>"110010011",
  5316=>"101111100",
  5317=>"011011011",
  5318=>"001000000",
  5319=>"100010010",
  5320=>"000111111",
  5321=>"101100001",
  5322=>"010100110",
  5323=>"001010001",
  5324=>"111101111",
  5325=>"010100011",
  5326=>"011111001",
  5327=>"111000100",
  5328=>"000001100",
  5329=>"100011001",
  5330=>"101111001",
  5331=>"110000011",
  5332=>"001101110",
  5333=>"100001001",
  5334=>"111101100",
  5335=>"011110000",
  5336=>"001111000",
  5337=>"010111101",
  5338=>"000001000",
  5339=>"011001001",
  5340=>"101110000",
  5341=>"101111101",
  5342=>"101001011",
  5343=>"001100101",
  5344=>"001011111",
  5345=>"100001111",
  5346=>"110001011",
  5347=>"010010100",
  5348=>"111110011",
  5349=>"110000100",
  5350=>"110111101",
  5351=>"111011110",
  5352=>"101111101",
  5353=>"000001111",
  5354=>"000000100",
  5355=>"001001011",
  5356=>"000011001",
  5357=>"011000000",
  5358=>"001100010",
  5359=>"011000000",
  5360=>"010010101",
  5361=>"110110001",
  5362=>"000010010",
  5363=>"101101001",
  5364=>"001100000",
  5365=>"001010100",
  5366=>"111100110",
  5367=>"011100100",
  5368=>"001111111",
  5369=>"101010111",
  5370=>"011111111",
  5371=>"001110011",
  5372=>"101100100",
  5373=>"000101011",
  5374=>"100111101",
  5375=>"111100101",
  5376=>"111010010",
  5377=>"010110000",
  5378=>"010110010",
  5379=>"100000001",
  5380=>"000110001",
  5381=>"000101101",
  5382=>"010110000",
  5383=>"111000001",
  5384=>"000011000",
  5385=>"000100001",
  5386=>"011100001",
  5387=>"111110110",
  5388=>"101100001",
  5389=>"001010100",
  5390=>"011001000",
  5391=>"010000011",
  5392=>"010101100",
  5393=>"001100111",
  5394=>"001011000",
  5395=>"001011001",
  5396=>"101011100",
  5397=>"001110110",
  5398=>"010101111",
  5399=>"011110111",
  5400=>"100100100",
  5401=>"011001000",
  5402=>"001110000",
  5403=>"001010010",
  5404=>"001011010",
  5405=>"010011100",
  5406=>"011011011",
  5407=>"010101111",
  5408=>"001001101",
  5409=>"100111010",
  5410=>"011111110",
  5411=>"100110100",
  5412=>"101010001",
  5413=>"010011001",
  5414=>"010111100",
  5415=>"101011010",
  5416=>"011111100",
  5417=>"111110011",
  5418=>"100000101",
  5419=>"110010110",
  5420=>"010010000",
  5421=>"000101101",
  5422=>"010100001",
  5423=>"000010101",
  5424=>"000001100",
  5425=>"101100010",
  5426=>"011001000",
  5427=>"110110111",
  5428=>"010110111",
  5429=>"100000010",
  5430=>"101101010",
  5431=>"101111110",
  5432=>"101000011",
  5433=>"111000010",
  5434=>"011100100",
  5435=>"111001110",
  5436=>"101111011",
  5437=>"011101111",
  5438=>"101001100",
  5439=>"111111100",
  5440=>"100111001",
  5441=>"101101101",
  5442=>"000011110",
  5443=>"101100101",
  5444=>"111100001",
  5445=>"110110100",
  5446=>"100001100",
  5447=>"000101110",
  5448=>"000101111",
  5449=>"111101110",
  5450=>"011010111",
  5451=>"000000000",
  5452=>"010110110",
  5453=>"000111100",
  5454=>"101000010",
  5455=>"101010110",
  5456=>"100011000",
  5457=>"011111000",
  5458=>"100011110",
  5459=>"000100110",
  5460=>"000100011",
  5461=>"101000001",
  5462=>"101000000",
  5463=>"111100011",
  5464=>"000001000",
  5465=>"110001010",
  5466=>"000010110",
  5467=>"100010111",
  5468=>"101110001",
  5469=>"111111011",
  5470=>"010101010",
  5471=>"110100110",
  5472=>"010011111",
  5473=>"110101001",
  5474=>"100111111",
  5475=>"101111010",
  5476=>"001111010",
  5477=>"010101110",
  5478=>"100001000",
  5479=>"100111111",
  5480=>"110111100",
  5481=>"000010001",
  5482=>"001010011",
  5483=>"010101110",
  5484=>"101001001",
  5485=>"111010101",
  5486=>"011111101",
  5487=>"101100100",
  5488=>"000011111",
  5489=>"111110111",
  5490=>"010001100",
  5491=>"010000100",
  5492=>"101011110",
  5493=>"100110000",
  5494=>"001000001",
  5495=>"111101101",
  5496=>"011110101",
  5497=>"101010110",
  5498=>"001110110",
  5499=>"100110001",
  5500=>"010011001",
  5501=>"000000000",
  5502=>"010111100",
  5503=>"000110011",
  5504=>"110010101",
  5505=>"001101110",
  5506=>"011110101",
  5507=>"110100110",
  5508=>"100010100",
  5509=>"000111001",
  5510=>"110001100",
  5511=>"011000000",
  5512=>"111111110",
  5513=>"100110101",
  5514=>"001000001",
  5515=>"100110010",
  5516=>"111101011",
  5517=>"110010101",
  5518=>"000101111",
  5519=>"010011010",
  5520=>"000101001",
  5521=>"000011001",
  5522=>"000100000",
  5523=>"001001100",
  5524=>"111110001",
  5525=>"010110111",
  5526=>"001000010",
  5527=>"001100110",
  5528=>"101100110",
  5529=>"011010000",
  5530=>"011110100",
  5531=>"001000110",
  5532=>"010011011",
  5533=>"010011011",
  5534=>"000100110",
  5535=>"111010011",
  5536=>"100001111",
  5537=>"010101000",
  5538=>"001010001",
  5539=>"011011001",
  5540=>"011000101",
  5541=>"000000010",
  5542=>"010011111",
  5543=>"100111010",
  5544=>"101011111",
  5545=>"111000000",
  5546=>"001110101",
  5547=>"100101011",
  5548=>"110110010",
  5549=>"101101001",
  5550=>"111010100",
  5551=>"011011001",
  5552=>"110001011",
  5553=>"001111000",
  5554=>"100010111",
  5555=>"000000011",
  5556=>"000010000",
  5557=>"100110101",
  5558=>"011111011",
  5559=>"000101101",
  5560=>"110011000",
  5561=>"000000111",
  5562=>"010001000",
  5563=>"011001000",
  5564=>"100111001",
  5565=>"110000100",
  5566=>"011010110",
  5567=>"100110111",
  5568=>"010001000",
  5569=>"000010001",
  5570=>"111010101",
  5571=>"111101110",
  5572=>"101100011",
  5573=>"011011010",
  5574=>"110010101",
  5575=>"111111100",
  5576=>"111011110",
  5577=>"000100001",
  5578=>"001001110",
  5579=>"101100101",
  5580=>"001011000",
  5581=>"011000011",
  5582=>"110001001",
  5583=>"010000000",
  5584=>"011000010",
  5585=>"011110001",
  5586=>"001110011",
  5587=>"100110010",
  5588=>"000111111",
  5589=>"111111010",
  5590=>"110101110",
  5591=>"111100111",
  5592=>"101010111",
  5593=>"111011101",
  5594=>"101101011",
  5595=>"000010010",
  5596=>"111011000",
  5597=>"111101110",
  5598=>"001011111",
  5599=>"100000000",
  5600=>"110100111",
  5601=>"100100000",
  5602=>"110011000",
  5603=>"000001001",
  5604=>"111011101",
  5605=>"011000011",
  5606=>"101100111",
  5607=>"001000010",
  5608=>"001010000",
  5609=>"100001010",
  5610=>"000010011",
  5611=>"101000000",
  5612=>"000000011",
  5613=>"011010000",
  5614=>"100101110",
  5615=>"110001011",
  5616=>"110100101",
  5617=>"011100101",
  5618=>"110010111",
  5619=>"000100110",
  5620=>"111110101",
  5621=>"101001100",
  5622=>"110110110",
  5623=>"001000110",
  5624=>"001101000",
  5625=>"100100110",
  5626=>"111010000",
  5627=>"100101011",
  5628=>"111101101",
  5629=>"110000101",
  5630=>"010100101",
  5631=>"110110111",
  5632=>"001110010",
  5633=>"010011000",
  5634=>"100011100",
  5635=>"100001000",
  5636=>"111000000",
  5637=>"011001010",
  5638=>"101001010",
  5639=>"010111010",
  5640=>"110011100",
  5641=>"010100000",
  5642=>"000001010",
  5643=>"001001101",
  5644=>"111000011",
  5645=>"100000001",
  5646=>"111001111",
  5647=>"111001000",
  5648=>"110100011",
  5649=>"110000100",
  5650=>"001100101",
  5651=>"010101100",
  5652=>"001110011",
  5653=>"011010111",
  5654=>"101110100",
  5655=>"111111110",
  5656=>"010001100",
  5657=>"111011110",
  5658=>"000110011",
  5659=>"000111110",
  5660=>"000100100",
  5661=>"000011111",
  5662=>"111100111",
  5663=>"101110111",
  5664=>"011001111",
  5665=>"010001111",
  5666=>"100101011",
  5667=>"010110110",
  5668=>"110101101",
  5669=>"110011101",
  5670=>"001000010",
  5671=>"110100010",
  5672=>"010001010",
  5673=>"001110110",
  5674=>"000111111",
  5675=>"111101000",
  5676=>"111010011",
  5677=>"001001001",
  5678=>"000101001",
  5679=>"000001111",
  5680=>"011101100",
  5681=>"011101011",
  5682=>"101100000",
  5683=>"001011111",
  5684=>"010000100",
  5685=>"000011101",
  5686=>"010011010",
  5687=>"110000001",
  5688=>"110101100",
  5689=>"001100011",
  5690=>"111011111",
  5691=>"101110000",
  5692=>"101101000",
  5693=>"000000001",
  5694=>"110011110",
  5695=>"011111110",
  5696=>"010101000",
  5697=>"011101010",
  5698=>"110000111",
  5699=>"000010101",
  5700=>"101010011",
  5701=>"010010111",
  5702=>"100011111",
  5703=>"110011000",
  5704=>"010000111",
  5705=>"100010000",
  5706=>"101010000",
  5707=>"010100101",
  5708=>"110110010",
  5709=>"101101111",
  5710=>"111000111",
  5711=>"101000001",
  5712=>"101000010",
  5713=>"001011111",
  5714=>"001100000",
  5715=>"100101100",
  5716=>"101001011",
  5717=>"000111011",
  5718=>"100101001",
  5719=>"010110011",
  5720=>"010111011",
  5721=>"011000000",
  5722=>"011010101",
  5723=>"100100100",
  5724=>"000011100",
  5725=>"000001011",
  5726=>"001110000",
  5727=>"001110111",
  5728=>"111110001",
  5729=>"101011000",
  5730=>"011111110",
  5731=>"110010100",
  5732=>"001100111",
  5733=>"100100100",
  5734=>"010001000",
  5735=>"111110001",
  5736=>"000011010",
  5737=>"101001000",
  5738=>"010101101",
  5739=>"010101110",
  5740=>"100011101",
  5741=>"011000100",
  5742=>"111010111",
  5743=>"100101000",
  5744=>"101110101",
  5745=>"110010111",
  5746=>"000111010",
  5747=>"010110001",
  5748=>"110000111",
  5749=>"100101101",
  5750=>"101010111",
  5751=>"111100000",
  5752=>"001101010",
  5753=>"000111001",
  5754=>"110110011",
  5755=>"110010000",
  5756=>"100000000",
  5757=>"110000011",
  5758=>"011110010",
  5759=>"110111010",
  5760=>"101110000",
  5761=>"110101001",
  5762=>"001010110",
  5763=>"011000100",
  5764=>"000101111",
  5765=>"111010101",
  5766=>"000011010",
  5767=>"011011101",
  5768=>"011011010",
  5769=>"011111010",
  5770=>"000000100",
  5771=>"001000010",
  5772=>"011101010",
  5773=>"000100110",
  5774=>"111111000",
  5775=>"010001001",
  5776=>"111110110",
  5777=>"111001000",
  5778=>"010100101",
  5779=>"001001010",
  5780=>"000110110",
  5781=>"001001101",
  5782=>"110101000",
  5783=>"010100011",
  5784=>"000101011",
  5785=>"011000101",
  5786=>"010100010",
  5787=>"000001100",
  5788=>"011001010",
  5789=>"100000100",
  5790=>"010000111",
  5791=>"001100001",
  5792=>"010000111",
  5793=>"110010101",
  5794=>"100101000",
  5795=>"011110101",
  5796=>"010011000",
  5797=>"111110101",
  5798=>"110111000",
  5799=>"100000010",
  5800=>"100011100",
  5801=>"010000001",
  5802=>"100010111",
  5803=>"001001011",
  5804=>"001101010",
  5805=>"010011010",
  5806=>"111111010",
  5807=>"000001010",
  5808=>"111001100",
  5809=>"011101010",
  5810=>"010010111",
  5811=>"011011111",
  5812=>"000011011",
  5813=>"101000010",
  5814=>"001001100",
  5815=>"100011011",
  5816=>"001111101",
  5817=>"001011001",
  5818=>"101110001",
  5819=>"001111001",
  5820=>"011010100",
  5821=>"001011111",
  5822=>"101100001",
  5823=>"110010011",
  5824=>"111111111",
  5825=>"000000101",
  5826=>"010000100",
  5827=>"100111000",
  5828=>"000011110",
  5829=>"111000000",
  5830=>"001100011",
  5831=>"110100101",
  5832=>"101000111",
  5833=>"100000010",
  5834=>"001001000",
  5835=>"100001010",
  5836=>"010010001",
  5837=>"111111001",
  5838=>"010011101",
  5839=>"000010000",
  5840=>"100111011",
  5841=>"000111000",
  5842=>"110111101",
  5843=>"111110000",
  5844=>"000000000",
  5845=>"000011111",
  5846=>"000101000",
  5847=>"110111101",
  5848=>"011000000",
  5849=>"010111100",
  5850=>"000101011",
  5851=>"110110010",
  5852=>"110101011",
  5853=>"011110111",
  5854=>"110111111",
  5855=>"110110000",
  5856=>"010000010",
  5857=>"010101011",
  5858=>"100111110",
  5859=>"101010101",
  5860=>"011010011",
  5861=>"000101010",
  5862=>"111010111",
  5863=>"100101101",
  5864=>"100101110",
  5865=>"000111000",
  5866=>"100111101",
  5867=>"010010001",
  5868=>"101111101",
  5869=>"111000101",
  5870=>"010000101",
  5871=>"100000101",
  5872=>"111011110",
  5873=>"100111011",
  5874=>"000001011",
  5875=>"101011000",
  5876=>"110010011",
  5877=>"111101101",
  5878=>"011000110",
  5879=>"010110110",
  5880=>"011011111",
  5881=>"010100001",
  5882=>"110000100",
  5883=>"101001001",
  5884=>"101100010",
  5885=>"000100001",
  5886=>"011010010",
  5887=>"000111111",
  5888=>"001000010",
  5889=>"111000110",
  5890=>"110100001",
  5891=>"100100100",
  5892=>"110010101",
  5893=>"000000010",
  5894=>"010011100",
  5895=>"000010100",
  5896=>"111000100",
  5897=>"111001000",
  5898=>"001011101",
  5899=>"111011101",
  5900=>"110100100",
  5901=>"111010000",
  5902=>"010110111",
  5903=>"111001000",
  5904=>"100111111",
  5905=>"000000100",
  5906=>"110001010",
  5907=>"001011111",
  5908=>"111111101",
  5909=>"011101110",
  5910=>"101001111",
  5911=>"100001111",
  5912=>"000000011",
  5913=>"110110101",
  5914=>"111011001",
  5915=>"100111011",
  5916=>"101011110",
  5917=>"100100001",
  5918=>"110110001",
  5919=>"110100111",
  5920=>"000101111",
  5921=>"010011011",
  5922=>"011110011",
  5923=>"000011001",
  5924=>"111111110",
  5925=>"011101010",
  5926=>"000101011",
  5927=>"010101100",
  5928=>"010001011",
  5929=>"111000111",
  5930=>"000000111",
  5931=>"010000000",
  5932=>"001001001",
  5933=>"001000101",
  5934=>"001111111",
  5935=>"100111111",
  5936=>"100011011",
  5937=>"011110101",
  5938=>"001010111",
  5939=>"111001011",
  5940=>"001110000",
  5941=>"101100010",
  5942=>"111111000",
  5943=>"001110001",
  5944=>"110011101",
  5945=>"011000011",
  5946=>"100101100",
  5947=>"101100101",
  5948=>"000100001",
  5949=>"001001010",
  5950=>"010011101",
  5951=>"011010011",
  5952=>"111000000",
  5953=>"000100111",
  5954=>"011010010",
  5955=>"001110000",
  5956=>"100110001",
  5957=>"010111111",
  5958=>"110100110",
  5959=>"101110111",
  5960=>"000100001",
  5961=>"011111101",
  5962=>"000111001",
  5963=>"001011010",
  5964=>"010100111",
  5965=>"111001110",
  5966=>"011001101",
  5967=>"010110011",
  5968=>"000110110",
  5969=>"111111010",
  5970=>"010101011",
  5971=>"101001001",
  5972=>"101110101",
  5973=>"001010110",
  5974=>"110000011",
  5975=>"100110000",
  5976=>"010101110",
  5977=>"110010001",
  5978=>"100101010",
  5979=>"000000111",
  5980=>"111101110",
  5981=>"110010110",
  5982=>"010001101",
  5983=>"010001000",
  5984=>"100100010",
  5985=>"011111100",
  5986=>"000000111",
  5987=>"111100000",
  5988=>"110111101",
  5989=>"101110000",
  5990=>"111001011",
  5991=>"011010000",
  5992=>"010000100",
  5993=>"110010010",
  5994=>"110011000",
  5995=>"011010100",
  5996=>"001010111",
  5997=>"111000010",
  5998=>"010000101",
  5999=>"000000010",
  6000=>"010000100",
  6001=>"010111101",
  6002=>"110101010",
  6003=>"110111010",
  6004=>"011110100",
  6005=>"100110100",
  6006=>"010100100",
  6007=>"100001101",
  6008=>"000010000",
  6009=>"001111111",
  6010=>"000001000",
  6011=>"001101101",
  6012=>"101010001",
  6013=>"110011111",
  6014=>"000110000",
  6015=>"001100100",
  6016=>"101110111",
  6017=>"111011110",
  6018=>"111101010",
  6019=>"010001011",
  6020=>"001100011",
  6021=>"000100010",
  6022=>"010101110",
  6023=>"001000101",
  6024=>"010001100",
  6025=>"110010100",
  6026=>"000000001",
  6027=>"010010010",
  6028=>"000001001",
  6029=>"000100010",
  6030=>"101010010",
  6031=>"101111010",
  6032=>"001111001",
  6033=>"111101001",
  6034=>"111100111",
  6035=>"010011111",
  6036=>"010001010",
  6037=>"001100110",
  6038=>"101000000",
  6039=>"000111100",
  6040=>"100101011",
  6041=>"000111101",
  6042=>"111001011",
  6043=>"011110110",
  6044=>"010000000",
  6045=>"010000100",
  6046=>"100110001",
  6047=>"100110111",
  6048=>"001111101",
  6049=>"011010010",
  6050=>"100011000",
  6051=>"001000000",
  6052=>"101101100",
  6053=>"010010101",
  6054=>"001011000",
  6055=>"000100110",
  6056=>"001110111",
  6057=>"111110101",
  6058=>"101110111",
  6059=>"001000001",
  6060=>"000010010",
  6061=>"010010000",
  6062=>"101010010",
  6063=>"011101111",
  6064=>"001010001",
  6065=>"100101110",
  6066=>"110010001",
  6067=>"001101010",
  6068=>"101111110",
  6069=>"001110101",
  6070=>"001101000",
  6071=>"010100010",
  6072=>"011110000",
  6073=>"001101100",
  6074=>"001110111",
  6075=>"011000011",
  6076=>"111110010",
  6077=>"000011000",
  6078=>"001011010",
  6079=>"101000010",
  6080=>"110111000",
  6081=>"000111110",
  6082=>"010001011",
  6083=>"101010111",
  6084=>"101110001",
  6085=>"000100011",
  6086=>"001101100",
  6087=>"011000100",
  6088=>"100001000",
  6089=>"000001101",
  6090=>"101001101",
  6091=>"100100011",
  6092=>"111010110",
  6093=>"101000000",
  6094=>"111101110",
  6095=>"001101000",
  6096=>"111100010",
  6097=>"111000001",
  6098=>"011011111",
  6099=>"100111010",
  6100=>"001110001",
  6101=>"101000100",
  6102=>"001000001",
  6103=>"111001100",
  6104=>"000111100",
  6105=>"011110000",
  6106=>"000011010",
  6107=>"110011111",
  6108=>"011111001",
  6109=>"111000011",
  6110=>"011110010",
  6111=>"011101111",
  6112=>"110000101",
  6113=>"110100001",
  6114=>"101000100",
  6115=>"000011110",
  6116=>"111010111",
  6117=>"100000001",
  6118=>"100010000",
  6119=>"001001101",
  6120=>"100001110",
  6121=>"100011011",
  6122=>"100010100",
  6123=>"001000110",
  6124=>"000011000",
  6125=>"000101100",
  6126=>"000111101",
  6127=>"110001101",
  6128=>"011110111",
  6129=>"000111011",
  6130=>"011110011",
  6131=>"000101111",
  6132=>"110111000",
  6133=>"111011011",
  6134=>"100111100",
  6135=>"010111101",
  6136=>"100000010",
  6137=>"000111000",
  6138=>"001110101",
  6139=>"100101000",
  6140=>"101001101",
  6141=>"010010100",
  6142=>"100101001",
  6143=>"100001100",
  6144=>"110111011",
  6145=>"101100000",
  6146=>"100101101",
  6147=>"000001100",
  6148=>"100111101",
  6149=>"111000000",
  6150=>"011000010",
  6151=>"010101100",
  6152=>"000000011",
  6153=>"001111011",
  6154=>"100000011",
  6155=>"111011110",
  6156=>"001100001",
  6157=>"111001001",
  6158=>"110010001",
  6159=>"001101010",
  6160=>"000011110",
  6161=>"111101010",
  6162=>"011101101",
  6163=>"111101000",
  6164=>"111001010",
  6165=>"001101001",
  6166=>"110101010",
  6167=>"110001110",
  6168=>"100100010",
  6169=>"011110010",
  6170=>"001011001",
  6171=>"111011001",
  6172=>"111101000",
  6173=>"101101100",
  6174=>"111010011",
  6175=>"000110010",
  6176=>"100111110",
  6177=>"001110011",
  6178=>"100001100",
  6179=>"011101001",
  6180=>"011001111",
  6181=>"010101010",
  6182=>"100011001",
  6183=>"101100001",
  6184=>"000100001",
  6185=>"111100011",
  6186=>"111110001",
  6187=>"111010101",
  6188=>"101100101",
  6189=>"011110101",
  6190=>"100010010",
  6191=>"010000111",
  6192=>"011111011",
  6193=>"000100100",
  6194=>"110011010",
  6195=>"010111011",
  6196=>"011001010",
  6197=>"110101010",
  6198=>"100111111",
  6199=>"100001001",
  6200=>"011001100",
  6201=>"110110010",
  6202=>"100110111",
  6203=>"010011001",
  6204=>"010000000",
  6205=>"001101101",
  6206=>"000001101",
  6207=>"010111100",
  6208=>"111101011",
  6209=>"011100001",
  6210=>"111111101",
  6211=>"110001000",
  6212=>"100011010",
  6213=>"100001011",
  6214=>"111101110",
  6215=>"010111000",
  6216=>"111100100",
  6217=>"110010100",
  6218=>"011101110",
  6219=>"000010001",
  6220=>"100000111",
  6221=>"100000011",
  6222=>"110101001",
  6223=>"110000111",
  6224=>"100111101",
  6225=>"111010111",
  6226=>"101001111",
  6227=>"100001111",
  6228=>"001011101",
  6229=>"010111000",
  6230=>"001000110",
  6231=>"010111100",
  6232=>"100000100",
  6233=>"100111111",
  6234=>"000100001",
  6235=>"100110001",
  6236=>"001011010",
  6237=>"010000101",
  6238=>"101010110",
  6239=>"100110000",
  6240=>"011110110",
  6241=>"010101011",
  6242=>"000010111",
  6243=>"100101101",
  6244=>"011010111",
  6245=>"011100001",
  6246=>"011011010",
  6247=>"111000110",
  6248=>"011101010",
  6249=>"100011100",
  6250=>"100010101",
  6251=>"111100010",
  6252=>"000011010",
  6253=>"010101111",
  6254=>"001001101",
  6255=>"010101010",
  6256=>"101001000",
  6257=>"011101001",
  6258=>"101100011",
  6259=>"100110111",
  6260=>"000100111",
  6261=>"001011000",
  6262=>"000100100",
  6263=>"001110000",
  6264=>"110000000",
  6265=>"000011110",
  6266=>"110010001",
  6267=>"000011111",
  6268=>"101000110",
  6269=>"001000110",
  6270=>"100111110",
  6271=>"100101101",
  6272=>"111100111",
  6273=>"001100001",
  6274=>"101010111",
  6275=>"111011010",
  6276=>"111111011",
  6277=>"000000111",
  6278=>"100010001",
  6279=>"010001011",
  6280=>"111111111",
  6281=>"011001001",
  6282=>"011110000",
  6283=>"101100100",
  6284=>"100101000",
  6285=>"111011010",
  6286=>"110010100",
  6287=>"111111001",
  6288=>"010010100",
  6289=>"100001101",
  6290=>"101111100",
  6291=>"011010011",
  6292=>"000001001",
  6293=>"000010011",
  6294=>"100101110",
  6295=>"110111100",
  6296=>"011001000",
  6297=>"101011110",
  6298=>"001101111",
  6299=>"110101010",
  6300=>"010001011",
  6301=>"000000000",
  6302=>"011010001",
  6303=>"010010000",
  6304=>"100010111",
  6305=>"001101000",
  6306=>"111000001",
  6307=>"011110001",
  6308=>"111100101",
  6309=>"000110000",
  6310=>"000000001",
  6311=>"110101110",
  6312=>"100011001",
  6313=>"110101100",
  6314=>"111101110",
  6315=>"101110011",
  6316=>"000011100",
  6317=>"001110010",
  6318=>"110011100",
  6319=>"101110111",
  6320=>"100110000",
  6321=>"000100101",
  6322=>"001010010",
  6323=>"010000000",
  6324=>"010101000",
  6325=>"100000000",
  6326=>"110101100",
  6327=>"011100001",
  6328=>"111101011",
  6329=>"011110110",
  6330=>"111101011",
  6331=>"110000101",
  6332=>"000000011",
  6333=>"011110000",
  6334=>"011000011",
  6335=>"110001011",
  6336=>"111001110",
  6337=>"000000000",
  6338=>"100001110",
  6339=>"101011101",
  6340=>"000100011",
  6341=>"011111111",
  6342=>"111001011",
  6343=>"111100010",
  6344=>"011011110",
  6345=>"111110011",
  6346=>"011111101",
  6347=>"100010100",
  6348=>"101110011",
  6349=>"010000000",
  6350=>"010111011",
  6351=>"011001001",
  6352=>"111010010",
  6353=>"101001100",
  6354=>"010011011",
  6355=>"010101001",
  6356=>"111110010",
  6357=>"101010010",
  6358=>"001000101",
  6359=>"111011001",
  6360=>"011111011",
  6361=>"101101111",
  6362=>"011110011",
  6363=>"010101010",
  6364=>"000110001",
  6365=>"100000111",
  6366=>"001001001",
  6367=>"101011000",
  6368=>"011001111",
  6369=>"011010111",
  6370=>"101111000",
  6371=>"111101100",
  6372=>"001001000",
  6373=>"000010100",
  6374=>"010001000",
  6375=>"010000001",
  6376=>"101011001",
  6377=>"110011101",
  6378=>"110101000",
  6379=>"101000001",
  6380=>"001101110",
  6381=>"101111111",
  6382=>"111110011",
  6383=>"001100100",
  6384=>"001110000",
  6385=>"111000011",
  6386=>"000000101",
  6387=>"000000011",
  6388=>"111101010",
  6389=>"010111111",
  6390=>"000100110",
  6391=>"111111001",
  6392=>"111010001",
  6393=>"000011010",
  6394=>"001010001",
  6395=>"110101001",
  6396=>"101010100",
  6397=>"001000010",
  6398=>"011011101",
  6399=>"011101111",
  6400=>"110001101",
  6401=>"110100111",
  6402=>"101000000",
  6403=>"110010011",
  6404=>"010011110",
  6405=>"001101110",
  6406=>"110010011",
  6407=>"101001111",
  6408=>"000101100",
  6409=>"011001101",
  6410=>"100100011",
  6411=>"011110011",
  6412=>"000011101",
  6413=>"111111010",
  6414=>"011010010",
  6415=>"011010001",
  6416=>"110110001",
  6417=>"000010001",
  6418=>"101110100",
  6419=>"000000101",
  6420=>"110111100",
  6421=>"101111011",
  6422=>"101110101",
  6423=>"110111101",
  6424=>"111100101",
  6425=>"000101100",
  6426=>"011111100",
  6427=>"010100111",
  6428=>"111101000",
  6429=>"111000000",
  6430=>"100000100",
  6431=>"101011110",
  6432=>"110111000",
  6433=>"100100101",
  6434=>"000010011",
  6435=>"000001001",
  6436=>"111100100",
  6437=>"101101101",
  6438=>"011110110",
  6439=>"100000001",
  6440=>"001000000",
  6441=>"001101101",
  6442=>"010000110",
  6443=>"110100011",
  6444=>"001001000",
  6445=>"010110100",
  6446=>"000110100",
  6447=>"010100010",
  6448=>"000000100",
  6449=>"101001011",
  6450=>"110110101",
  6451=>"011001011",
  6452=>"101001010",
  6453=>"101110010",
  6454=>"010110000",
  6455=>"011100111",
  6456=>"011011011",
  6457=>"110100100",
  6458=>"011010011",
  6459=>"101100010",
  6460=>"010000110",
  6461=>"011010100",
  6462=>"110001011",
  6463=>"011110101",
  6464=>"101000000",
  6465=>"010111000",
  6466=>"110011100",
  6467=>"001101011",
  6468=>"111001010",
  6469=>"111111111",
  6470=>"111110110",
  6471=>"001011011",
  6472=>"111001010",
  6473=>"011100100",
  6474=>"110100100",
  6475=>"000001101",
  6476=>"001111011",
  6477=>"011101111",
  6478=>"101010010",
  6479=>"110111111",
  6480=>"111110101",
  6481=>"001000101",
  6482=>"101111011",
  6483=>"110001101",
  6484=>"111000000",
  6485=>"100101111",
  6486=>"101101110",
  6487=>"101000111",
  6488=>"001111101",
  6489=>"001111110",
  6490=>"111101110",
  6491=>"111000010",
  6492=>"100111101",
  6493=>"010000100",
  6494=>"101100110",
  6495=>"010010001",
  6496=>"110001010",
  6497=>"110000111",
  6498=>"100000000",
  6499=>"011000111",
  6500=>"101110001",
  6501=>"000101010",
  6502=>"010100011",
  6503=>"101000000",
  6504=>"110110110",
  6505=>"010101111",
  6506=>"011000100",
  6507=>"000011001",
  6508=>"111101011",
  6509=>"111111010",
  6510=>"010110100",
  6511=>"010101101",
  6512=>"000011010",
  6513=>"110101010",
  6514=>"111011111",
  6515=>"001011101",
  6516=>"001110010",
  6517=>"111110110",
  6518=>"000111110",
  6519=>"101001100",
  6520=>"010000101",
  6521=>"101111011",
  6522=>"000110101",
  6523=>"000110110",
  6524=>"101110011",
  6525=>"000101100",
  6526=>"000000010",
  6527=>"011011101",
  6528=>"110100111",
  6529=>"011000100",
  6530=>"110100100",
  6531=>"000000110",
  6532=>"110010000",
  6533=>"110100000",
  6534=>"111101010",
  6535=>"011110100",
  6536=>"010000111",
  6537=>"001110001",
  6538=>"000010001",
  6539=>"000100000",
  6540=>"011010001",
  6541=>"111001011",
  6542=>"011010101",
  6543=>"111101110",
  6544=>"101110110",
  6545=>"011000001",
  6546=>"100111110",
  6547=>"110110101",
  6548=>"000110111",
  6549=>"001010010",
  6550=>"010001011",
  6551=>"001011000",
  6552=>"100000001",
  6553=>"000001111",
  6554=>"001010011",
  6555=>"100001111",
  6556=>"111110011",
  6557=>"010101100",
  6558=>"101101001",
  6559=>"000011011",
  6560=>"011010011",
  6561=>"000000101",
  6562=>"100110100",
  6563=>"101110010",
  6564=>"010001010",
  6565=>"110100000",
  6566=>"110110000",
  6567=>"101011001",
  6568=>"101001000",
  6569=>"100110101",
  6570=>"010000011",
  6571=>"111110011",
  6572=>"000110000",
  6573=>"001100010",
  6574=>"010001000",
  6575=>"100011010",
  6576=>"100101000",
  6577=>"011000000",
  6578=>"001110010",
  6579=>"100100001",
  6580=>"111100001",
  6581=>"111110111",
  6582=>"011011110",
  6583=>"100101011",
  6584=>"001010110",
  6585=>"110010011",
  6586=>"011011001",
  6587=>"100010000",
  6588=>"111000010",
  6589=>"111110000",
  6590=>"100011001",
  6591=>"101001010",
  6592=>"111011001",
  6593=>"011000001",
  6594=>"011110110",
  6595=>"111101110",
  6596=>"000001011",
  6597=>"001001000",
  6598=>"111101100",
  6599=>"001010101",
  6600=>"110010100",
  6601=>"001011010",
  6602=>"001000000",
  6603=>"011000000",
  6604=>"100011000",
  6605=>"111010100",
  6606=>"110110000",
  6607=>"000101110",
  6608=>"011000110",
  6609=>"110001001",
  6610=>"011000011",
  6611=>"111100111",
  6612=>"100000101",
  6613=>"110001010",
  6614=>"110101001",
  6615=>"010011010",
  6616=>"110110101",
  6617=>"110111110",
  6618=>"110100100",
  6619=>"100111111",
  6620=>"100000011",
  6621=>"110101010",
  6622=>"110111011",
  6623=>"101010100",
  6624=>"111110001",
  6625=>"101000001",
  6626=>"100101011",
  6627=>"001011010",
  6628=>"110011010",
  6629=>"000010000",
  6630=>"011101011",
  6631=>"011000010",
  6632=>"010000110",
  6633=>"000000101",
  6634=>"101101011",
  6635=>"101011011",
  6636=>"011001100",
  6637=>"000101100",
  6638=>"011111011",
  6639=>"101110010",
  6640=>"001011110",
  6641=>"100011000",
  6642=>"010100110",
  6643=>"010101010",
  6644=>"001000111",
  6645=>"000101001",
  6646=>"011000010",
  6647=>"101100111",
  6648=>"100111010",
  6649=>"100010011",
  6650=>"010100101",
  6651=>"010011011",
  6652=>"011101010",
  6653=>"110110110",
  6654=>"001100010",
  6655=>"100101101",
  6656=>"000001111",
  6657=>"100011100",
  6658=>"000000011",
  6659=>"011010100",
  6660=>"000110101",
  6661=>"010100100",
  6662=>"011111001",
  6663=>"011110111",
  6664=>"011001000",
  6665=>"101100110",
  6666=>"010100101",
  6667=>"100100110",
  6668=>"101011101",
  6669=>"101110011",
  6670=>"001001100",
  6671=>"100110011",
  6672=>"110100001",
  6673=>"000101100",
  6674=>"001101111",
  6675=>"110011111",
  6676=>"111110010",
  6677=>"001001011",
  6678=>"011110100",
  6679=>"111110100",
  6680=>"111011101",
  6681=>"100010101",
  6682=>"010000011",
  6683=>"000101100",
  6684=>"100010000",
  6685=>"101110100",
  6686=>"100111101",
  6687=>"000001111",
  6688=>"000100010",
  6689=>"110110011",
  6690=>"100011100",
  6691=>"101000100",
  6692=>"100001001",
  6693=>"101010110",
  6694=>"000000010",
  6695=>"001111110",
  6696=>"010000011",
  6697=>"111010110",
  6698=>"110001111",
  6699=>"101110111",
  6700=>"110101010",
  6701=>"001011100",
  6702=>"101010111",
  6703=>"000000100",
  6704=>"000101111",
  6705=>"011001011",
  6706=>"010010100",
  6707=>"111101110",
  6708=>"110111110",
  6709=>"000000100",
  6710=>"100100110",
  6711=>"110101101",
  6712=>"101111100",
  6713=>"001000110",
  6714=>"100100010",
  6715=>"111011001",
  6716=>"101001110",
  6717=>"101110110",
  6718=>"110010011",
  6719=>"110010010",
  6720=>"010000100",
  6721=>"000000001",
  6722=>"001101111",
  6723=>"000111110",
  6724=>"001110010",
  6725=>"101011010",
  6726=>"001110101",
  6727=>"100011111",
  6728=>"100011101",
  6729=>"000111101",
  6730=>"100000100",
  6731=>"001001000",
  6732=>"111100000",
  6733=>"001110100",
  6734=>"010010010",
  6735=>"011010011",
  6736=>"110010100",
  6737=>"100000001",
  6738=>"111011001",
  6739=>"010010011",
  6740=>"000000100",
  6741=>"011111110",
  6742=>"111010111",
  6743=>"000101010",
  6744=>"000100100",
  6745=>"001111000",
  6746=>"100010111",
  6747=>"010010101",
  6748=>"100010010",
  6749=>"111100101",
  6750=>"010001111",
  6751=>"010011001",
  6752=>"110010101",
  6753=>"001011111",
  6754=>"000010110",
  6755=>"101110011",
  6756=>"011101100",
  6757=>"000001110",
  6758=>"111000100",
  6759=>"000101101",
  6760=>"111001001",
  6761=>"111111110",
  6762=>"010010011",
  6763=>"010000010",
  6764=>"110010001",
  6765=>"111111010",
  6766=>"100111010",
  6767=>"000000111",
  6768=>"010111111",
  6769=>"111111110",
  6770=>"011010101",
  6771=>"000101000",
  6772=>"011111000",
  6773=>"001001110",
  6774=>"111111101",
  6775=>"011111110",
  6776=>"000100101",
  6777=>"010111100",
  6778=>"110000000",
  6779=>"111001000",
  6780=>"110000110",
  6781=>"010000011",
  6782=>"011011001",
  6783=>"001011110",
  6784=>"101100011",
  6785=>"110000010",
  6786=>"100011001",
  6787=>"000011010",
  6788=>"000011000",
  6789=>"101110100",
  6790=>"001010110",
  6791=>"111100101",
  6792=>"110101101",
  6793=>"100010110",
  6794=>"000110101",
  6795=>"101110100",
  6796=>"010000010",
  6797=>"011010011",
  6798=>"100010001",
  6799=>"100110001",
  6800=>"110101101",
  6801=>"010010010",
  6802=>"111001101",
  6803=>"101000111",
  6804=>"111100011",
  6805=>"101010001",
  6806=>"011000000",
  6807=>"000011101",
  6808=>"000000100",
  6809=>"100111110",
  6810=>"101110110",
  6811=>"000011011",
  6812=>"100111010",
  6813=>"000000001",
  6814=>"000001100",
  6815=>"110110100",
  6816=>"011010110",
  6817=>"101000111",
  6818=>"110001010",
  6819=>"011100111",
  6820=>"101110100",
  6821=>"101010011",
  6822=>"101010100",
  6823=>"000110011",
  6824=>"110100000",
  6825=>"110000000",
  6826=>"101001011",
  6827=>"001010110",
  6828=>"110111001",
  6829=>"101111001",
  6830=>"001000011",
  6831=>"100100001",
  6832=>"001000101",
  6833=>"001010001",
  6834=>"000011111",
  6835=>"111011010",
  6836=>"011000010",
  6837=>"010111110",
  6838=>"011100010",
  6839=>"110001100",
  6840=>"101000000",
  6841=>"100011101",
  6842=>"011011111",
  6843=>"011110111",
  6844=>"100000101",
  6845=>"000011100",
  6846=>"011100101",
  6847=>"001111001",
  6848=>"010010011",
  6849=>"011110011",
  6850=>"010110111",
  6851=>"001100111",
  6852=>"001001001",
  6853=>"000000000",
  6854=>"110110011",
  6855=>"010010001",
  6856=>"001110010",
  6857=>"001010000",
  6858=>"111001001",
  6859=>"111111110",
  6860=>"110000111",
  6861=>"110111111",
  6862=>"000100011",
  6863=>"000000000",
  6864=>"100110111",
  6865=>"010001111",
  6866=>"100101011",
  6867=>"000110010",
  6868=>"010111111",
  6869=>"001100010",
  6870=>"011011010",
  6871=>"110110001",
  6872=>"000011111",
  6873=>"010110110",
  6874=>"111011110",
  6875=>"010101000",
  6876=>"001101011",
  6877=>"001001001",
  6878=>"110110010",
  6879=>"100001011",
  6880=>"100010101",
  6881=>"110001111",
  6882=>"101001101",
  6883=>"111001100",
  6884=>"000011001",
  6885=>"011011101",
  6886=>"101111001",
  6887=>"010101101",
  6888=>"101000110",
  6889=>"000110001",
  6890=>"011111101",
  6891=>"101010111",
  6892=>"111111100",
  6893=>"111111101",
  6894=>"100010001",
  6895=>"000101010",
  6896=>"100010101",
  6897=>"100010000",
  6898=>"101011010",
  6899=>"010001100",
  6900=>"101010010",
  6901=>"110101011",
  6902=>"000000000",
  6903=>"101011101",
  6904=>"000000101",
  6905=>"110111111",
  6906=>"100100101",
  6907=>"100000011",
  6908=>"010011011",
  6909=>"010001001",
  6910=>"111010101",
  6911=>"000000011",
  6912=>"111001111",
  6913=>"111001010",
  6914=>"000101011",
  6915=>"001000001",
  6916=>"000010110",
  6917=>"011100010",
  6918=>"111100011",
  6919=>"111000100",
  6920=>"101111101",
  6921=>"100001001",
  6922=>"001100000",
  6923=>"101111000",
  6924=>"111000001",
  6925=>"111111111",
  6926=>"110000001",
  6927=>"100011100",
  6928=>"001100101",
  6929=>"010100111",
  6930=>"010110011",
  6931=>"000011111",
  6932=>"100111110",
  6933=>"011111010",
  6934=>"011010110",
  6935=>"011000010",
  6936=>"110010010",
  6937=>"110101111",
  6938=>"001100010",
  6939=>"110101101",
  6940=>"000100000",
  6941=>"101111001",
  6942=>"011101101",
  6943=>"100011110",
  6944=>"011111111",
  6945=>"010100101",
  6946=>"010001110",
  6947=>"110110001",
  6948=>"010100001",
  6949=>"111000000",
  6950=>"100111011",
  6951=>"101000111",
  6952=>"001100001",
  6953=>"100110110",
  6954=>"110001101",
  6955=>"001100100",
  6956=>"110011000",
  6957=>"001100010",
  6958=>"010010011",
  6959=>"010100000",
  6960=>"111101111",
  6961=>"001110110",
  6962=>"000001000",
  6963=>"111100000",
  6964=>"110110011",
  6965=>"101011010",
  6966=>"011000111",
  6967=>"111011001",
  6968=>"010011010",
  6969=>"001100010",
  6970=>"110111110",
  6971=>"111000100",
  6972=>"111111000",
  6973=>"000111110",
  6974=>"100010001",
  6975=>"101110001",
  6976=>"001010011",
  6977=>"100001011",
  6978=>"110000111",
  6979=>"001100001",
  6980=>"100101001",
  6981=>"101010100",
  6982=>"110100111",
  6983=>"101000100",
  6984=>"100111011",
  6985=>"101101110",
  6986=>"000111101",
  6987=>"111010010",
  6988=>"011101011",
  6989=>"100011001",
  6990=>"010010110",
  6991=>"000001111",
  6992=>"011001111",
  6993=>"101001000",
  6994=>"000100100",
  6995=>"101001010",
  6996=>"101111011",
  6997=>"010111111",
  6998=>"000100111",
  6999=>"101111011",
  7000=>"000010111",
  7001=>"000110010",
  7002=>"010000000",
  7003=>"010101000",
  7004=>"000001101",
  7005=>"100000010",
  7006=>"101100000",
  7007=>"100010101",
  7008=>"111100111",
  7009=>"010100001",
  7010=>"110000010",
  7011=>"001110111",
  7012=>"101010111",
  7013=>"001000011",
  7014=>"111001011",
  7015=>"111101111",
  7016=>"010100101",
  7017=>"110100010",
  7018=>"100111101",
  7019=>"011110010",
  7020=>"001000001",
  7021=>"111111010",
  7022=>"111111011",
  7023=>"110000101",
  7024=>"011010111",
  7025=>"101000010",
  7026=>"010101010",
  7027=>"000100001",
  7028=>"000001101",
  7029=>"010000101",
  7030=>"110011101",
  7031=>"111011101",
  7032=>"000101010",
  7033=>"000000011",
  7034=>"000101011",
  7035=>"111001110",
  7036=>"011001100",
  7037=>"110011011",
  7038=>"110010000",
  7039=>"011101101",
  7040=>"111101100",
  7041=>"010100111",
  7042=>"111101110",
  7043=>"000010000",
  7044=>"101001000",
  7045=>"000100101",
  7046=>"010011100",
  7047=>"111000000",
  7048=>"000110011",
  7049=>"111010110",
  7050=>"000000011",
  7051=>"000111000",
  7052=>"100011011",
  7053=>"111001111",
  7054=>"100010000",
  7055=>"011101100",
  7056=>"000000000",
  7057=>"111100011",
  7058=>"100001010",
  7059=>"111010000",
  7060=>"000101100",
  7061=>"100011110",
  7062=>"110110111",
  7063=>"001100111",
  7064=>"101111000",
  7065=>"101111010",
  7066=>"000010001",
  7067=>"000111011",
  7068=>"010000000",
  7069=>"101001110",
  7070=>"111000110",
  7071=>"001101010",
  7072=>"000000100",
  7073=>"111010010",
  7074=>"110110011",
  7075=>"111101101",
  7076=>"100001011",
  7077=>"000100110",
  7078=>"001101000",
  7079=>"111101010",
  7080=>"111001111",
  7081=>"111111111",
  7082=>"101101010",
  7083=>"001011111",
  7084=>"011110011",
  7085=>"000101111",
  7086=>"001011011",
  7087=>"111010011",
  7088=>"100101011",
  7089=>"111101000",
  7090=>"000111001",
  7091=>"010001011",
  7092=>"110000001",
  7093=>"111010010",
  7094=>"011110110",
  7095=>"000011111",
  7096=>"111010011",
  7097=>"001100011",
  7098=>"001111101",
  7099=>"000111010",
  7100=>"010100011",
  7101=>"111111001",
  7102=>"110000111",
  7103=>"001101111",
  7104=>"001000111",
  7105=>"001001010",
  7106=>"100010010",
  7107=>"100011011",
  7108=>"100011001",
  7109=>"010001110",
  7110=>"111000111",
  7111=>"100110100",
  7112=>"010001010",
  7113=>"000010000",
  7114=>"001100010",
  7115=>"111100000",
  7116=>"111011101",
  7117=>"101111111",
  7118=>"011011010",
  7119=>"111111101",
  7120=>"111110110",
  7121=>"101111000",
  7122=>"011011010",
  7123=>"101010011",
  7124=>"100010111",
  7125=>"101000111",
  7126=>"111111011",
  7127=>"100100010",
  7128=>"010010011",
  7129=>"010000101",
  7130=>"110110100",
  7131=>"010001000",
  7132=>"100011100",
  7133=>"000101010",
  7134=>"100110100",
  7135=>"110001011",
  7136=>"011010110",
  7137=>"001000000",
  7138=>"111111010",
  7139=>"111010000",
  7140=>"111011011",
  7141=>"111101000",
  7142=>"010000111",
  7143=>"110100110",
  7144=>"001111010",
  7145=>"001001101",
  7146=>"101110111",
  7147=>"000000010",
  7148=>"110010011",
  7149=>"111011001",
  7150=>"100111011",
  7151=>"110111101",
  7152=>"001001110",
  7153=>"011000000",
  7154=>"100011100",
  7155=>"111001000",
  7156=>"101000011",
  7157=>"001010001",
  7158=>"000111001",
  7159=>"010010111",
  7160=>"101011111",
  7161=>"001001011",
  7162=>"110111000",
  7163=>"111000101",
  7164=>"000101110",
  7165=>"101111110",
  7166=>"111101101",
  7167=>"111100001",
  7168=>"001010000",
  7169=>"100011111",
  7170=>"110010000",
  7171=>"001111000",
  7172=>"100001001",
  7173=>"010000001",
  7174=>"001110110",
  7175=>"110100110",
  7176=>"100101101",
  7177=>"100101010",
  7178=>"110111100",
  7179=>"011001010",
  7180=>"010001010",
  7181=>"101111010",
  7182=>"101111010",
  7183=>"100001101",
  7184=>"010000000",
  7185=>"001000010",
  7186=>"100100111",
  7187=>"000011100",
  7188=>"000011011",
  7189=>"001011110",
  7190=>"110101100",
  7191=>"111111100",
  7192=>"110100011",
  7193=>"101000010",
  7194=>"111010101",
  7195=>"110111001",
  7196=>"010001111",
  7197=>"010010110",
  7198=>"111101100",
  7199=>"000011010",
  7200=>"111110001",
  7201=>"001100010",
  7202=>"001001111",
  7203=>"000101110",
  7204=>"011101011",
  7205=>"110100010",
  7206=>"001111100",
  7207=>"001101001",
  7208=>"011101011",
  7209=>"101100011",
  7210=>"010101100",
  7211=>"010010110",
  7212=>"000010100",
  7213=>"111111100",
  7214=>"010111001",
  7215=>"110100000",
  7216=>"001111010",
  7217=>"000000100",
  7218=>"010100000",
  7219=>"111011101",
  7220=>"100111010",
  7221=>"100101000",
  7222=>"011111001",
  7223=>"001110011",
  7224=>"001011000",
  7225=>"111111110",
  7226=>"110011101",
  7227=>"000000110",
  7228=>"111100000",
  7229=>"111000101",
  7230=>"001010001",
  7231=>"001010111",
  7232=>"001101010",
  7233=>"001110101",
  7234=>"110101101",
  7235=>"101111000",
  7236=>"001011010",
  7237=>"001101011",
  7238=>"000100001",
  7239=>"010001101",
  7240=>"100011101",
  7241=>"000011011",
  7242=>"000000100",
  7243=>"110001100",
  7244=>"101111110",
  7245=>"111001110",
  7246=>"111100110",
  7247=>"110010001",
  7248=>"100000110",
  7249=>"111111101",
  7250=>"001000011",
  7251=>"110110011",
  7252=>"111111111",
  7253=>"110100010",
  7254=>"000000000",
  7255=>"101001100",
  7256=>"111011000",
  7257=>"100111001",
  7258=>"111110010",
  7259=>"100010110",
  7260=>"110111111",
  7261=>"000011100",
  7262=>"101000110",
  7263=>"001010011",
  7264=>"010111111",
  7265=>"111111111",
  7266=>"110111010",
  7267=>"100111101",
  7268=>"100100001",
  7269=>"011110010",
  7270=>"101111100",
  7271=>"101001110",
  7272=>"100001001",
  7273=>"100110111",
  7274=>"100100001",
  7275=>"110100111",
  7276=>"101001111",
  7277=>"100100000",
  7278=>"011000011",
  7279=>"111111111",
  7280=>"000111110",
  7281=>"010101000",
  7282=>"110111111",
  7283=>"100011110",
  7284=>"000011001",
  7285=>"110111100",
  7286=>"101110011",
  7287=>"000111111",
  7288=>"011101110",
  7289=>"111110001",
  7290=>"000001100",
  7291=>"110011110",
  7292=>"111111110",
  7293=>"110110011",
  7294=>"011111011",
  7295=>"010001000",
  7296=>"101011000",
  7297=>"110010110",
  7298=>"000011110",
  7299=>"011011010",
  7300=>"000010110",
  7301=>"111010010",
  7302=>"001001100",
  7303=>"010010000",
  7304=>"011110110",
  7305=>"000011000",
  7306=>"101000010",
  7307=>"110110101",
  7308=>"011010100",
  7309=>"001001100",
  7310=>"111001100",
  7311=>"111110001",
  7312=>"111110010",
  7313=>"110110111",
  7314=>"100110011",
  7315=>"010011010",
  7316=>"010010110",
  7317=>"111000101",
  7318=>"111111110",
  7319=>"101000110",
  7320=>"000001100",
  7321=>"100111010",
  7322=>"000100001",
  7323=>"000101100",
  7324=>"101101001",
  7325=>"100111001",
  7326=>"010010000",
  7327=>"000111111",
  7328=>"111010101",
  7329=>"010001001",
  7330=>"111100101",
  7331=>"011100111",
  7332=>"100100000",
  7333=>"011110101",
  7334=>"101111000",
  7335=>"111100101",
  7336=>"000000010",
  7337=>"111011000",
  7338=>"111110111",
  7339=>"011000010",
  7340=>"000100011",
  7341=>"011000100",
  7342=>"011100100",
  7343=>"000111010",
  7344=>"001101000",
  7345=>"000001000",
  7346=>"100110000",
  7347=>"101001000",
  7348=>"111100011",
  7349=>"110011000",
  7350=>"100100101",
  7351=>"000101000",
  7352=>"101001100",
  7353=>"001111111",
  7354=>"000011110",
  7355=>"100110100",
  7356=>"011101011",
  7357=>"111101001",
  7358=>"010000010",
  7359=>"100101001",
  7360=>"001000100",
  7361=>"111111000",
  7362=>"111100101",
  7363=>"111010000",
  7364=>"100101110",
  7365=>"010010000",
  7366=>"111111000",
  7367=>"000111100",
  7368=>"000010011",
  7369=>"000010101",
  7370=>"000011100",
  7371=>"100000111",
  7372=>"111101101",
  7373=>"101100010",
  7374=>"111001101",
  7375=>"111001000",
  7376=>"000001010",
  7377=>"011000010",
  7378=>"111000011",
  7379=>"000011111",
  7380=>"000010000",
  7381=>"000101011",
  7382=>"011010011",
  7383=>"111111101",
  7384=>"101110100",
  7385=>"111101011",
  7386=>"011011101",
  7387=>"111110001",
  7388=>"000010101",
  7389=>"101011100",
  7390=>"000010100",
  7391=>"000101000",
  7392=>"001000111",
  7393=>"101111011",
  7394=>"011010110",
  7395=>"011101100",
  7396=>"101000111",
  7397=>"001000010",
  7398=>"011111110",
  7399=>"000011111",
  7400=>"001111100",
  7401=>"101101110",
  7402=>"000010110",
  7403=>"010001110",
  7404=>"100110111",
  7405=>"000101111",
  7406=>"101001001",
  7407=>"100111011",
  7408=>"000100011",
  7409=>"111010110",
  7410=>"001110010",
  7411=>"111101100",
  7412=>"000010001",
  7413=>"111001001",
  7414=>"000010011",
  7415=>"010001100",
  7416=>"100100001",
  7417=>"101011101",
  7418=>"011101111",
  7419=>"101100010",
  7420=>"001010101",
  7421=>"000000101",
  7422=>"011100111",
  7423=>"001010011",
  7424=>"001001100",
  7425=>"001110000",
  7426=>"100000111",
  7427=>"001111010",
  7428=>"010011100",
  7429=>"101111000",
  7430=>"010000101",
  7431=>"101110001",
  7432=>"101000100",
  7433=>"111011001",
  7434=>"111110001",
  7435=>"100101001",
  7436=>"100001101",
  7437=>"010000111",
  7438=>"100111111",
  7439=>"000010010",
  7440=>"101000111",
  7441=>"100101010",
  7442=>"110111111",
  7443=>"001101101",
  7444=>"111110011",
  7445=>"110000001",
  7446=>"101110000",
  7447=>"010110001",
  7448=>"100001100",
  7449=>"111011001",
  7450=>"101111001",
  7451=>"011100010",
  7452=>"000101000",
  7453=>"111000011",
  7454=>"001100001",
  7455=>"100100110",
  7456=>"111111001",
  7457=>"111001010",
  7458=>"100111111",
  7459=>"111101010",
  7460=>"001111101",
  7461=>"001011101",
  7462=>"010011100",
  7463=>"110011110",
  7464=>"000000110",
  7465=>"111110110",
  7466=>"111100110",
  7467=>"001001000",
  7468=>"110100010",
  7469=>"011101000",
  7470=>"111100000",
  7471=>"010101001",
  7472=>"101010111",
  7473=>"101011100",
  7474=>"001110011",
  7475=>"100100100",
  7476=>"001001001",
  7477=>"001011100",
  7478=>"010100001",
  7479=>"111101111",
  7480=>"100010001",
  7481=>"110111110",
  7482=>"011001100",
  7483=>"001011001",
  7484=>"001001011",
  7485=>"100010101",
  7486=>"010110110",
  7487=>"101011111",
  7488=>"111010110",
  7489=>"100111110",
  7490=>"011111110",
  7491=>"111001000",
  7492=>"010111111",
  7493=>"111010101",
  7494=>"010110000",
  7495=>"001101111",
  7496=>"110001101",
  7497=>"001101010",
  7498=>"110001010",
  7499=>"111101111",
  7500=>"000010101",
  7501=>"110000111",
  7502=>"000001010",
  7503=>"101110011",
  7504=>"000000001",
  7505=>"110000001",
  7506=>"000101100",
  7507=>"000111111",
  7508=>"000000000",
  7509=>"000111000",
  7510=>"000100101",
  7511=>"011111000",
  7512=>"011011111",
  7513=>"001100111",
  7514=>"001110100",
  7515=>"000101001",
  7516=>"001111100",
  7517=>"001100101",
  7518=>"111110001",
  7519=>"010000101",
  7520=>"110100110",
  7521=>"010110111",
  7522=>"100010000",
  7523=>"100000011",
  7524=>"000110000",
  7525=>"111110100",
  7526=>"100011101",
  7527=>"111110111",
  7528=>"010010111",
  7529=>"011111010",
  7530=>"011011111",
  7531=>"100110100",
  7532=>"101101010",
  7533=>"100001101",
  7534=>"011010111",
  7535=>"101000000",
  7536=>"101001000",
  7537=>"110100001",
  7538=>"111111111",
  7539=>"101110110",
  7540=>"101111001",
  7541=>"011010100",
  7542=>"011001000",
  7543=>"010111101",
  7544=>"101001000",
  7545=>"101101100",
  7546=>"101000101",
  7547=>"110010011",
  7548=>"010111011",
  7549=>"000011100",
  7550=>"001010001",
  7551=>"000101011",
  7552=>"101111111",
  7553=>"011000010",
  7554=>"100000000",
  7555=>"010111111",
  7556=>"111001010",
  7557=>"111101110",
  7558=>"110011100",
  7559=>"100111101",
  7560=>"000011010",
  7561=>"001110101",
  7562=>"111011101",
  7563=>"001001001",
  7564=>"110110000",
  7565=>"000101001",
  7566=>"001110011",
  7567=>"001111010",
  7568=>"000000100",
  7569=>"111000000",
  7570=>"000011001",
  7571=>"100010011",
  7572=>"100000011",
  7573=>"011101000",
  7574=>"101100111",
  7575=>"011010101",
  7576=>"000100000",
  7577=>"011101011",
  7578=>"110100011",
  7579=>"101000011",
  7580=>"001100001",
  7581=>"011000010",
  7582=>"110010010",
  7583=>"010110111",
  7584=>"111101001",
  7585=>"111101011",
  7586=>"110001011",
  7587=>"110010000",
  7588=>"111010100",
  7589=>"010010001",
  7590=>"100101011",
  7591=>"011101100",
  7592=>"100000100",
  7593=>"100001000",
  7594=>"000001000",
  7595=>"110010101",
  7596=>"010110011",
  7597=>"000110111",
  7598=>"011011110",
  7599=>"000100111",
  7600=>"111111101",
  7601=>"000100001",
  7602=>"001010100",
  7603=>"101011101",
  7604=>"000001011",
  7605=>"100011111",
  7606=>"110100101",
  7607=>"101011011",
  7608=>"001001111",
  7609=>"011101010",
  7610=>"001011101",
  7611=>"111011101",
  7612=>"010100101",
  7613=>"100100000",
  7614=>"000110011",
  7615=>"010000110",
  7616=>"011101111",
  7617=>"010000110",
  7618=>"101111101",
  7619=>"010010110",
  7620=>"001111011",
  7621=>"011100100",
  7622=>"000100000",
  7623=>"000111111",
  7624=>"001010000",
  7625=>"011101010",
  7626=>"001001000",
  7627=>"001100101",
  7628=>"011100010",
  7629=>"100110001",
  7630=>"111111101",
  7631=>"100101011",
  7632=>"010111011",
  7633=>"000011010",
  7634=>"100111111",
  7635=>"011000100",
  7636=>"111111110",
  7637=>"011101011",
  7638=>"100110010",
  7639=>"010001001",
  7640=>"111000010",
  7641=>"111110001",
  7642=>"100010101",
  7643=>"111111011",
  7644=>"011011010",
  7645=>"001010101",
  7646=>"110010001",
  7647=>"001011101",
  7648=>"111101001",
  7649=>"101111010",
  7650=>"011000001",
  7651=>"000110000",
  7652=>"001011100",
  7653=>"101111111",
  7654=>"100000101",
  7655=>"110110011",
  7656=>"010110101",
  7657=>"011001000",
  7658=>"110101001",
  7659=>"111110111",
  7660=>"111100011",
  7661=>"010001101",
  7662=>"100000000",
  7663=>"001100111",
  7664=>"010111100",
  7665=>"000000111",
  7666=>"110101011",
  7667=>"100110100",
  7668=>"110110101",
  7669=>"110110110",
  7670=>"000011000",
  7671=>"000000100",
  7672=>"001000101",
  7673=>"010000110",
  7674=>"101011000",
  7675=>"101000110",
  7676=>"110110001",
  7677=>"110010111",
  7678=>"110110011",
  7679=>"011111111",
  7680=>"100010011",
  7681=>"111110000",
  7682=>"100011100",
  7683=>"010100010",
  7684=>"011001000",
  7685=>"100011111",
  7686=>"011100110",
  7687=>"111111110",
  7688=>"000001000",
  7689=>"110011100",
  7690=>"001100001",
  7691=>"010011111",
  7692=>"001011011",
  7693=>"011011101",
  7694=>"101001110",
  7695=>"101010111",
  7696=>"101001100",
  7697=>"100000101",
  7698=>"100111000",
  7699=>"100101011",
  7700=>"011100101",
  7701=>"011111001",
  7702=>"110101011",
  7703=>"100001001",
  7704=>"110110110",
  7705=>"011010100",
  7706=>"000110001",
  7707=>"001011000",
  7708=>"010101010",
  7709=>"000101000",
  7710=>"000001110",
  7711=>"011001010",
  7712=>"111001101",
  7713=>"000111110",
  7714=>"111000000",
  7715=>"100000110",
  7716=>"011111100",
  7717=>"000011111",
  7718=>"000010110",
  7719=>"111000001",
  7720=>"010110111",
  7721=>"011010000",
  7722=>"111111101",
  7723=>"101101111",
  7724=>"101110111",
  7725=>"100101100",
  7726=>"111000000",
  7727=>"110010001",
  7728=>"000011010",
  7729=>"110011010",
  7730=>"010110100",
  7731=>"011111001",
  7732=>"100101101",
  7733=>"111010000",
  7734=>"001000100",
  7735=>"001111111",
  7736=>"010011111",
  7737=>"010011011",
  7738=>"101100000",
  7739=>"110101100",
  7740=>"110001101",
  7741=>"111001000",
  7742=>"110110101",
  7743=>"011001001",
  7744=>"000110010",
  7745=>"001010111",
  7746=>"101111010",
  7747=>"000000100",
  7748=>"110010000",
  7749=>"001001010",
  7750=>"000000000",
  7751=>"000010000",
  7752=>"101111010",
  7753=>"011111100",
  7754=>"100011000",
  7755=>"001111010",
  7756=>"100110111",
  7757=>"100101111",
  7758=>"010100000",
  7759=>"011100000",
  7760=>"111011100",
  7761=>"001000001",
  7762=>"111011011",
  7763=>"011100000",
  7764=>"001011010",
  7765=>"111101001",
  7766=>"110100101",
  7767=>"001111001",
  7768=>"000001110",
  7769=>"000010000",
  7770=>"100001001",
  7771=>"011111111",
  7772=>"101111010",
  7773=>"001100001",
  7774=>"001110111",
  7775=>"101010111",
  7776=>"011100100",
  7777=>"100011011",
  7778=>"010001101",
  7779=>"100100100",
  7780=>"101010101",
  7781=>"001010011",
  7782=>"111010111",
  7783=>"001101010",
  7784=>"001110110",
  7785=>"010101000",
  7786=>"100101011",
  7787=>"101011000",
  7788=>"001001010",
  7789=>"111001001",
  7790=>"000001101",
  7791=>"111111100",
  7792=>"011001100",
  7793=>"000011100",
  7794=>"110110000",
  7795=>"000001001",
  7796=>"100101011",
  7797=>"011000101",
  7798=>"011011111",
  7799=>"000000010",
  7800=>"101101011",
  7801=>"110111110",
  7802=>"100011011",
  7803=>"010111100",
  7804=>"001010001",
  7805=>"101011100",
  7806=>"001111000",
  7807=>"110101001",
  7808=>"000000010",
  7809=>"100111100",
  7810=>"010010100",
  7811=>"000011010",
  7812=>"001110001",
  7813=>"110110101",
  7814=>"110001000",
  7815=>"000101111",
  7816=>"001011000",
  7817=>"101010101",
  7818=>"000110110",
  7819=>"000100001",
  7820=>"010000110",
  7821=>"000001101",
  7822=>"010101110",
  7823=>"010000011",
  7824=>"000110110",
  7825=>"100011100",
  7826=>"011101000",
  7827=>"101010101",
  7828=>"000000011",
  7829=>"001011001",
  7830=>"010000011",
  7831=>"011101111",
  7832=>"001111100",
  7833=>"011011001",
  7834=>"100010000",
  7835=>"001001101",
  7836=>"011000000",
  7837=>"111101010",
  7838=>"101001100",
  7839=>"110000010",
  7840=>"110010000",
  7841=>"100110100",
  7842=>"101011001",
  7843=>"010100000",
  7844=>"101111011",
  7845=>"001101101",
  7846=>"000101010",
  7847=>"001001111",
  7848=>"110000010",
  7849=>"111110110",
  7850=>"011011000",
  7851=>"110011001",
  7852=>"101000111",
  7853=>"111011001",
  7854=>"000011100",
  7855=>"001011000",
  7856=>"111010111",
  7857=>"110010000",
  7858=>"100011110",
  7859=>"101110000",
  7860=>"000010100",
  7861=>"101001011",
  7862=>"100110011",
  7863=>"100111000",
  7864=>"111110110",
  7865=>"001110001",
  7866=>"000001101",
  7867=>"111111110",
  7868=>"000010010",
  7869=>"011010100",
  7870=>"010101111",
  7871=>"110010100",
  7872=>"101011011",
  7873=>"001110011",
  7874=>"101011010",
  7875=>"101100110",
  7876=>"110000100",
  7877=>"000111110",
  7878=>"000111111",
  7879=>"001010011",
  7880=>"111111111",
  7881=>"000111000",
  7882=>"001000011",
  7883=>"111010101",
  7884=>"111011110",
  7885=>"010000001",
  7886=>"100110010",
  7887=>"110101101",
  7888=>"111111101",
  7889=>"110000100",
  7890=>"000001011",
  7891=>"011000100",
  7892=>"010011010",
  7893=>"000101111",
  7894=>"010001001",
  7895=>"000001000",
  7896=>"111110111",
  7897=>"100010110",
  7898=>"111001010",
  7899=>"000011001",
  7900=>"001001100",
  7901=>"100010111",
  7902=>"110111001",
  7903=>"010001011",
  7904=>"100100001",
  7905=>"000010011",
  7906=>"000001001",
  7907=>"111111111",
  7908=>"110101100",
  7909=>"100110001",
  7910=>"100100000",
  7911=>"001011101",
  7912=>"100001001",
  7913=>"101101011",
  7914=>"000110010",
  7915=>"001001011",
  7916=>"101010111",
  7917=>"101010110",
  7918=>"011110001",
  7919=>"000111111",
  7920=>"111100110",
  7921=>"011001011",
  7922=>"011111010",
  7923=>"111000000",
  7924=>"101110110",
  7925=>"110101101",
  7926=>"101000001",
  7927=>"110110101",
  7928=>"010100110",
  7929=>"010001111",
  7930=>"010000111",
  7931=>"011111111",
  7932=>"101001111",
  7933=>"110110011",
  7934=>"000101011",
  7935=>"110110101",
  7936=>"000000011",
  7937=>"111011010",
  7938=>"000001001",
  7939=>"010000010",
  7940=>"010001101",
  7941=>"000101101",
  7942=>"001001000",
  7943=>"111010101",
  7944=>"010000110",
  7945=>"110011001",
  7946=>"100101011",
  7947=>"101101010",
  7948=>"000110000",
  7949=>"100111110",
  7950=>"100011000",
  7951=>"010001000",
  7952=>"100000010",
  7953=>"010110000",
  7954=>"111011001",
  7955=>"110000101",
  7956=>"001100100",
  7957=>"010011001",
  7958=>"111111100",
  7959=>"010101000",
  7960=>"111001001",
  7961=>"001101110",
  7962=>"000010101",
  7963=>"111111011",
  7964=>"010100110",
  7965=>"010100001",
  7966=>"100111101",
  7967=>"010110000",
  7968=>"111001001",
  7969=>"100101000",
  7970=>"001100101",
  7971=>"111100101",
  7972=>"011001000",
  7973=>"000101111",
  7974=>"110111101",
  7975=>"100010001",
  7976=>"110010101",
  7977=>"000000110",
  7978=>"111000111",
  7979=>"011110100",
  7980=>"010110100",
  7981=>"100011110",
  7982=>"111011110",
  7983=>"111110111",
  7984=>"101001001",
  7985=>"011000000",
  7986=>"101111000",
  7987=>"010011000",
  7988=>"011010000",
  7989=>"101010101",
  7990=>"111111000",
  7991=>"011011110",
  7992=>"110110010",
  7993=>"011110111",
  7994=>"010010010",
  7995=>"010011110",
  7996=>"101100000",
  7997=>"010010001",
  7998=>"001111110",
  7999=>"111100111",
  8000=>"001100110",
  8001=>"110111100",
  8002=>"000000001",
  8003=>"111101101",
  8004=>"101010111",
  8005=>"000000111",
  8006=>"110101101",
  8007=>"011011111",
  8008=>"100100111",
  8009=>"010011010",
  8010=>"000001000",
  8011=>"011101110",
  8012=>"010111111",
  8013=>"111111110",
  8014=>"001110101",
  8015=>"001110101",
  8016=>"111111001",
  8017=>"000011101",
  8018=>"010101011",
  8019=>"111011000",
  8020=>"101011111",
  8021=>"111001011",
  8022=>"101111101",
  8023=>"001100110",
  8024=>"100111001",
  8025=>"111110000",
  8026=>"100011011",
  8027=>"000100100",
  8028=>"111100111",
  8029=>"110110000",
  8030=>"100001101",
  8031=>"111110010",
  8032=>"100000110",
  8033=>"100001110",
  8034=>"100110010",
  8035=>"011101001",
  8036=>"011001101",
  8037=>"010110010",
  8038=>"011100001",
  8039=>"101100110",
  8040=>"010101001",
  8041=>"000110101",
  8042=>"000101000",
  8043=>"111101011",
  8044=>"000110000",
  8045=>"010011001",
  8046=>"111011111",
  8047=>"111111111",
  8048=>"011001011",
  8049=>"000111111",
  8050=>"111101011",
  8051=>"000100100",
  8052=>"110011110",
  8053=>"001000110",
  8054=>"011111011",
  8055=>"010111100",
  8056=>"100101000",
  8057=>"101111001",
  8058=>"010111011",
  8059=>"011100000",
  8060=>"111101111",
  8061=>"100101101",
  8062=>"111111100",
  8063=>"000111010",
  8064=>"001010100",
  8065=>"010001010",
  8066=>"111110110",
  8067=>"110111101",
  8068=>"111101000",
  8069=>"110001110",
  8070=>"111111100",
  8071=>"010011000",
  8072=>"101001001",
  8073=>"111011001",
  8074=>"111100001",
  8075=>"000000000",
  8076=>"111100101",
  8077=>"110101010",
  8078=>"010001000",
  8079=>"111000110",
  8080=>"111111101",
  8081=>"100100010",
  8082=>"001000001",
  8083=>"000010010",
  8084=>"111000101",
  8085=>"010000001",
  8086=>"010110000",
  8087=>"011000011",
  8088=>"100111001",
  8089=>"101001001",
  8090=>"001010011",
  8091=>"100111110",
  8092=>"110000101",
  8093=>"101011000",
  8094=>"010110000",
  8095=>"010011100",
  8096=>"001110100",
  8097=>"001000001",
  8098=>"001011010",
  8099=>"011011000",
  8100=>"101101110",
  8101=>"000000011",
  8102=>"100010001",
  8103=>"010100010",
  8104=>"000111111",
  8105=>"100001100",
  8106=>"111101101",
  8107=>"001101010",
  8108=>"110111111",
  8109=>"111110101",
  8110=>"001111111",
  8111=>"000001100",
  8112=>"010100111",
  8113=>"110010111",
  8114=>"110001010",
  8115=>"011100001",
  8116=>"011010111",
  8117=>"101000100",
  8118=>"011101011",
  8119=>"111001101",
  8120=>"100101011",
  8121=>"100111101",
  8122=>"001001001",
  8123=>"110111110",
  8124=>"111000101",
  8125=>"110001101",
  8126=>"111101111",
  8127=>"000101111",
  8128=>"100110011",
  8129=>"111011011",
  8130=>"001110000",
  8131=>"100100001",
  8132=>"101011100",
  8133=>"001000000",
  8134=>"011101100",
  8135=>"100111110",
  8136=>"010000011",
  8137=>"111100011",
  8138=>"001000100",
  8139=>"011011100",
  8140=>"011011001",
  8141=>"100101011",
  8142=>"111111101",
  8143=>"011010010",
  8144=>"111000011",
  8145=>"001110101",
  8146=>"011000000",
  8147=>"110100111",
  8148=>"111011110",
  8149=>"111111111",
  8150=>"010111000",
  8151=>"111110000",
  8152=>"100000101",
  8153=>"110101100",
  8154=>"101000111",
  8155=>"111011110",
  8156=>"110000110",
  8157=>"011010000",
  8158=>"001111100",
  8159=>"110101000",
  8160=>"110000100",
  8161=>"110010010",
  8162=>"000000101",
  8163=>"101011110",
  8164=>"111011111",
  8165=>"000000100",
  8166=>"100011011",
  8167=>"100100111",
  8168=>"101100010",
  8169=>"100010111",
  8170=>"101010111",
  8171=>"100000111",
  8172=>"101000001",
  8173=>"001011010",
  8174=>"100000001",
  8175=>"011110110",
  8176=>"101111100",
  8177=>"000001001",
  8178=>"100011111",
  8179=>"000100100",
  8180=>"010101100",
  8181=>"010000000",
  8182=>"111010100",
  8183=>"011100000",
  8184=>"111010110",
  8185=>"101101000",
  8186=>"101010101",
  8187=>"001000001",
  8188=>"111100110",
  8189=>"101111010",
  8190=>"101001111",
  8191=>"000111110",
  8192=>"110000100",
  8193=>"111100111",
  8194=>"011010111",
  8195=>"101110000",
  8196=>"001010010",
  8197=>"100011000",
  8198=>"010001100",
  8199=>"011111001",
  8200=>"010101110",
  8201=>"011100101",
  8202=>"100100011",
  8203=>"000001111",
  8204=>"111110110",
  8205=>"100100101",
  8206=>"011100101",
  8207=>"111011111",
  8208=>"000011010",
  8209=>"100001100",
  8210=>"000011101",
  8211=>"110100110",
  8212=>"111000011",
  8213=>"010100100",
  8214=>"111011101",
  8215=>"100111100",
  8216=>"011001011",
  8217=>"101111111",
  8218=>"100011111",
  8219=>"111111111",
  8220=>"100011010",
  8221=>"100010100",
  8222=>"100100110",
  8223=>"111000011",
  8224=>"010011111",
  8225=>"111010100",
  8226=>"100100111",
  8227=>"110111111",
  8228=>"000100111",
  8229=>"000111110",
  8230=>"110001110",
  8231=>"111000100",
  8232=>"010100000",
  8233=>"100101111",
  8234=>"111001010",
  8235=>"110100000",
  8236=>"000100110",
  8237=>"010001011",
  8238=>"001011100",
  8239=>"101110110",
  8240=>"010101010",
  8241=>"100100010",
  8242=>"000001001",
  8243=>"001011111",
  8244=>"011101101",
  8245=>"101011101",
  8246=>"001100010",
  8247=>"101111000",
  8248=>"110111110",
  8249=>"100011010",
  8250=>"101000010",
  8251=>"111011010",
  8252=>"000111000",
  8253=>"001100100",
  8254=>"000100001",
  8255=>"110011110",
  8256=>"010000010",
  8257=>"011101100",
  8258=>"111100011",
  8259=>"101100110",
  8260=>"100011110",
  8261=>"100001000",
  8262=>"000000111",
  8263=>"001101111",
  8264=>"111101100",
  8265=>"010101110",
  8266=>"011100111",
  8267=>"110001111",
  8268=>"100010000",
  8269=>"000100100",
  8270=>"100111001",
  8271=>"011111110",
  8272=>"001010110",
  8273=>"001001000",
  8274=>"101100010",
  8275=>"111110100",
  8276=>"101011011",
  8277=>"100101111",
  8278=>"010010010",
  8279=>"001011100",
  8280=>"101011001",
  8281=>"101001110",
  8282=>"011110000",
  8283=>"110000000",
  8284=>"010111000",
  8285=>"001100110",
  8286=>"100000010",
  8287=>"111000100",
  8288=>"000101011",
  8289=>"111011010",
  8290=>"001110011",
  8291=>"101010000",
  8292=>"001010001",
  8293=>"000010110",
  8294=>"011010000",
  8295=>"111101101",
  8296=>"101100010",
  8297=>"011101000",
  8298=>"100000100",
  8299=>"101100001",
  8300=>"100101001",
  8301=>"100001001",
  8302=>"001110001",
  8303=>"111000110",
  8304=>"101100100",
  8305=>"000011110",
  8306=>"001000011",
  8307=>"011111100",
  8308=>"100010100",
  8309=>"000111001",
  8310=>"011110110",
  8311=>"000101001",
  8312=>"010111100",
  8313=>"010011011",
  8314=>"110101011",
  8315=>"011000000",
  8316=>"000111111",
  8317=>"011110110",
  8318=>"011101000",
  8319=>"011001110",
  8320=>"000010000",
  8321=>"000001000",
  8322=>"010010000",
  8323=>"010001011",
  8324=>"010000001",
  8325=>"011010100",
  8326=>"100000011",
  8327=>"100110110",
  8328=>"001100001",
  8329=>"111110000",
  8330=>"010100000",
  8331=>"010010000",
  8332=>"010010000",
  8333=>"011110000",
  8334=>"000110100",
  8335=>"101011111",
  8336=>"100110010",
  8337=>"111000110",
  8338=>"001000001",
  8339=>"111100111",
  8340=>"000010010",
  8341=>"000101011",
  8342=>"111011100",
  8343=>"111110101",
  8344=>"111111111",
  8345=>"010100101",
  8346=>"100100100",
  8347=>"100001110",
  8348=>"101001100",
  8349=>"010001100",
  8350=>"110100000",
  8351=>"101000000",
  8352=>"110010000",
  8353=>"001100111",
  8354=>"000010001",
  8355=>"110110111",
  8356=>"111101011",
  8357=>"111110100",
  8358=>"000111011",
  8359=>"000100000",
  8360=>"000000001",
  8361=>"111110110",
  8362=>"010010100",
  8363=>"000110001",
  8364=>"010111100",
  8365=>"000111101",
  8366=>"000000110",
  8367=>"110001111",
  8368=>"010100110",
  8369=>"110010100",
  8370=>"010000010",
  8371=>"001111101",
  8372=>"100011001",
  8373=>"111110001",
  8374=>"101001111",
  8375=>"010111110",
  8376=>"101000010",
  8377=>"111011110",
  8378=>"110011000",
  8379=>"101010000",
  8380=>"100110011",
  8381=>"101000001",
  8382=>"101100111",
  8383=>"001011110",
  8384=>"110010111",
  8385=>"111110101",
  8386=>"011011010",
  8387=>"000010001",
  8388=>"101011011",
  8389=>"111001110",
  8390=>"101000011",
  8391=>"000000110",
  8392=>"011001100",
  8393=>"000110111",
  8394=>"101101101",
  8395=>"001000101",
  8396=>"010000010",
  8397=>"110100111",
  8398=>"010010010",
  8399=>"111000111",
  8400=>"001100000",
  8401=>"000011001",
  8402=>"000100010",
  8403=>"110000001",
  8404=>"001111110",
  8405=>"111011100",
  8406=>"011100011",
  8407=>"011101011",
  8408=>"010101001",
  8409=>"001000011",
  8410=>"000000110",
  8411=>"101000000",
  8412=>"001101010",
  8413=>"010100010",
  8414=>"110010110",
  8415=>"000101010",
  8416=>"100101100",
  8417=>"110011000",
  8418=>"001010100",
  8419=>"010000011",
  8420=>"110010011",
  8421=>"100111111",
  8422=>"101111001",
  8423=>"001010001",
  8424=>"001001000",
  8425=>"011110101",
  8426=>"010011100",
  8427=>"011010100",
  8428=>"100010001",
  8429=>"100010110",
  8430=>"010101000",
  8431=>"001100101",
  8432=>"000110000",
  8433=>"011101111",
  8434=>"101110100",
  8435=>"101101101",
  8436=>"010011001",
  8437=>"000001000",
  8438=>"111111011",
  8439=>"111110110",
  8440=>"100111000",
  8441=>"010000000",
  8442=>"010111100",
  8443=>"100010100",
  8444=>"010011011",
  8445=>"110010001",
  8446=>"000000101",
  8447=>"010011100",
  8448=>"011001101",
  8449=>"110011001",
  8450=>"000001111",
  8451=>"000101011",
  8452=>"000111001",
  8453=>"100111101",
  8454=>"111100101",
  8455=>"111010110",
  8456=>"110111101",
  8457=>"000010111",
  8458=>"000001111",
  8459=>"000110101",
  8460=>"101100101",
  8461=>"010111111",
  8462=>"000101011",
  8463=>"011001000",
  8464=>"011110000",
  8465=>"000011110",
  8466=>"010100100",
  8467=>"101000100",
  8468=>"011100101",
  8469=>"101011011",
  8470=>"001101000",
  8471=>"110000110",
  8472=>"011100111",
  8473=>"111011111",
  8474=>"111011011",
  8475=>"110001010",
  8476=>"000011101",
  8477=>"101010010",
  8478=>"000101001",
  8479=>"001000110",
  8480=>"000010100",
  8481=>"100100101",
  8482=>"111101110",
  8483=>"110111000",
  8484=>"010111100",
  8485=>"001100000",
  8486=>"011100100",
  8487=>"110110010",
  8488=>"101111000",
  8489=>"110011011",
  8490=>"001100010",
  8491=>"001010100",
  8492=>"110010110",
  8493=>"111111101",
  8494=>"001011001",
  8495=>"100101000",
  8496=>"011000100",
  8497=>"101000110",
  8498=>"110011011",
  8499=>"000001000",
  8500=>"101011100",
  8501=>"001011101",
  8502=>"100111001",
  8503=>"010111011",
  8504=>"011111101",
  8505=>"001000011",
  8506=>"000011110",
  8507=>"001111001",
  8508=>"001110110",
  8509=>"111111111",
  8510=>"000000010",
  8511=>"001101100",
  8512=>"100010111",
  8513=>"111111101",
  8514=>"001000001",
  8515=>"110010100",
  8516=>"000010000",
  8517=>"001001110",
  8518=>"010110000",
  8519=>"000100100",
  8520=>"000100001",
  8521=>"000010110",
  8522=>"011001110",
  8523=>"001000000",
  8524=>"100001000",
  8525=>"111001110",
  8526=>"110000110",
  8527=>"110011000",
  8528=>"110000000",
  8529=>"110001101",
  8530=>"001011100",
  8531=>"001110111",
  8532=>"010000011",
  8533=>"110010000",
  8534=>"111000111",
  8535=>"011111010",
  8536=>"110101010",
  8537=>"010110010",
  8538=>"001000101",
  8539=>"101100100",
  8540=>"001101101",
  8541=>"100001101",
  8542=>"101010101",
  8543=>"000010000",
  8544=>"100101011",
  8545=>"000100100",
  8546=>"111000110",
  8547=>"001010101",
  8548=>"110100101",
  8549=>"011000011",
  8550=>"111001011",
  8551=>"111011010",
  8552=>"110010011",
  8553=>"001000101",
  8554=>"101010101",
  8555=>"001001111",
  8556=>"100100010",
  8557=>"111100000",
  8558=>"000100101",
  8559=>"111011000",
  8560=>"100011101",
  8561=>"110010010",
  8562=>"101000111",
  8563=>"100010110",
  8564=>"010010010",
  8565=>"110111111",
  8566=>"010011011",
  8567=>"111110101",
  8568=>"010100101",
  8569=>"011110111",
  8570=>"001010100",
  8571=>"101110001",
  8572=>"110101011",
  8573=>"001011011",
  8574=>"001000101",
  8575=>"000111110",
  8576=>"101111000",
  8577=>"000101000",
  8578=>"100101111",
  8579=>"111100110",
  8580=>"001100001",
  8581=>"001001010",
  8582=>"111011011",
  8583=>"111000101",
  8584=>"100110101",
  8585=>"100100110",
  8586=>"110111010",
  8587=>"010001000",
  8588=>"110010111",
  8589=>"110010001",
  8590=>"011001001",
  8591=>"111101011",
  8592=>"100001001",
  8593=>"010101111",
  8594=>"010010011",
  8595=>"011111011",
  8596=>"111010011",
  8597=>"000000101",
  8598=>"111111010",
  8599=>"011110100",
  8600=>"010100101",
  8601=>"000101011",
  8602=>"001000000",
  8603=>"110101111",
  8604=>"010010010",
  8605=>"000110001",
  8606=>"111111110",
  8607=>"101000111",
  8608=>"001000111",
  8609=>"111101001",
  8610=>"100011111",
  8611=>"111011110",
  8612=>"100000011",
  8613=>"111011001",
  8614=>"000000100",
  8615=>"101110100",
  8616=>"010110001",
  8617=>"011010011",
  8618=>"111100110",
  8619=>"011110100",
  8620=>"011110100",
  8621=>"110111010",
  8622=>"010111010",
  8623=>"111011110",
  8624=>"101001010",
  8625=>"010011101",
  8626=>"000100111",
  8627=>"000101001",
  8628=>"100010001",
  8629=>"010000011",
  8630=>"000001001",
  8631=>"111101110",
  8632=>"011111011",
  8633=>"000011010",
  8634=>"100001010",
  8635=>"010010010",
  8636=>"011110010",
  8637=>"001010001",
  8638=>"011010000",
  8639=>"100100100",
  8640=>"010010010",
  8641=>"000000100",
  8642=>"011001001",
  8643=>"001110110",
  8644=>"001011011",
  8645=>"111110001",
  8646=>"010101110",
  8647=>"010010011",
  8648=>"001001111",
  8649=>"111010111",
  8650=>"000110000",
  8651=>"010000000",
  8652=>"100011000",
  8653=>"111000101",
  8654=>"101010001",
  8655=>"001101001",
  8656=>"011011110",
  8657=>"110100000",
  8658=>"100010010",
  8659=>"100101010",
  8660=>"000001000",
  8661=>"111000010",
  8662=>"110111101",
  8663=>"010111000",
  8664=>"011010011",
  8665=>"111100111",
  8666=>"000110001",
  8667=>"100101011",
  8668=>"110001111",
  8669=>"011110011",
  8670=>"010010111",
  8671=>"111111011",
  8672=>"111010011",
  8673=>"010111000",
  8674=>"011011110",
  8675=>"000001111",
  8676=>"111100100",
  8677=>"100111010",
  8678=>"011000100",
  8679=>"100011100",
  8680=>"110000101",
  8681=>"110110100",
  8682=>"110000000",
  8683=>"001011000",
  8684=>"110000010",
  8685=>"100010000",
  8686=>"011111001",
  8687=>"011000111",
  8688=>"000001001",
  8689=>"011100100",
  8690=>"010001100",
  8691=>"101000000",
  8692=>"011101101",
  8693=>"101011011",
  8694=>"010001001",
  8695=>"010000001",
  8696=>"111111010",
  8697=>"101000000",
  8698=>"000011011",
  8699=>"111111000",
  8700=>"010000010",
  8701=>"000001000",
  8702=>"100010011",
  8703=>"110000001",
  8704=>"010000100",
  8705=>"110000010",
  8706=>"001010010",
  8707=>"001101011",
  8708=>"110000001",
  8709=>"110101100",
  8710=>"111100111",
  8711=>"000010111",
  8712=>"110001100",
  8713=>"010110000",
  8714=>"010110000",
  8715=>"010111111",
  8716=>"100011110",
  8717=>"111111010",
  8718=>"111001000",
  8719=>"010011011",
  8720=>"001101001",
  8721=>"000111011",
  8722=>"000010111",
  8723=>"101010100",
  8724=>"000010010",
  8725=>"000001011",
  8726=>"011111100",
  8727=>"100101000",
  8728=>"110000001",
  8729=>"001000101",
  8730=>"100110010",
  8731=>"110010010",
  8732=>"010010101",
  8733=>"100100010",
  8734=>"001101100",
  8735=>"011001111",
  8736=>"011010010",
  8737=>"110111111",
  8738=>"010011010",
  8739=>"101011010",
  8740=>"111010110",
  8741=>"001001011",
  8742=>"100011001",
  8743=>"101011100",
  8744=>"011110110",
  8745=>"001101001",
  8746=>"101000000",
  8747=>"100011001",
  8748=>"011101011",
  8749=>"111010000",
  8750=>"001001000",
  8751=>"000110100",
  8752=>"001101111",
  8753=>"011101010",
  8754=>"010101100",
  8755=>"011110011",
  8756=>"110110010",
  8757=>"010010100",
  8758=>"011100100",
  8759=>"011101011",
  8760=>"000000010",
  8761=>"100001100",
  8762=>"100100110",
  8763=>"101011110",
  8764=>"101111111",
  8765=>"100100000",
  8766=>"001111111",
  8767=>"001000111",
  8768=>"101000011",
  8769=>"111000111",
  8770=>"101100100",
  8771=>"101110100",
  8772=>"011100100",
  8773=>"100110000",
  8774=>"001010000",
  8775=>"001101011",
  8776=>"010101110",
  8777=>"001101110",
  8778=>"111101011",
  8779=>"011100011",
  8780=>"111001100",
  8781=>"011110010",
  8782=>"100001000",
  8783=>"101011000",
  8784=>"010010100",
  8785=>"000000110",
  8786=>"000111101",
  8787=>"111111100",
  8788=>"110010001",
  8789=>"010101010",
  8790=>"001011101",
  8791=>"111111111",
  8792=>"111101101",
  8793=>"101011011",
  8794=>"001110010",
  8795=>"110010000",
  8796=>"101001111",
  8797=>"100001011",
  8798=>"100001011",
  8799=>"101011100",
  8800=>"101001110",
  8801=>"010100011",
  8802=>"010110010",
  8803=>"011010001",
  8804=>"011010010",
  8805=>"111101110",
  8806=>"110000001",
  8807=>"010111101",
  8808=>"000000100",
  8809=>"000111111",
  8810=>"101101111",
  8811=>"101010011",
  8812=>"011100010",
  8813=>"011011000",
  8814=>"000111100",
  8815=>"000010010",
  8816=>"100101100",
  8817=>"010101001",
  8818=>"111010100",
  8819=>"100010011",
  8820=>"101111011",
  8821=>"111010000",
  8822=>"110011111",
  8823=>"100010011",
  8824=>"101010100",
  8825=>"010111010",
  8826=>"110000010",
  8827=>"101111001",
  8828=>"010001010",
  8829=>"000111000",
  8830=>"000000010",
  8831=>"110100110",
  8832=>"100010100",
  8833=>"000110101",
  8834=>"000000010",
  8835=>"111110111",
  8836=>"100111011",
  8837=>"101000100",
  8838=>"111000010",
  8839=>"000001101",
  8840=>"110001110",
  8841=>"011001011",
  8842=>"111111000",
  8843=>"111000000",
  8844=>"011111011",
  8845=>"110111001",
  8846=>"010001110",
  8847=>"110011000",
  8848=>"101101101",
  8849=>"001000010",
  8850=>"010010010",
  8851=>"000111010",
  8852=>"010001010",
  8853=>"111101100",
  8854=>"111100111",
  8855=>"111100101",
  8856=>"010000000",
  8857=>"101011110",
  8858=>"111111101",
  8859=>"000011000",
  8860=>"111010011",
  8861=>"100001101",
  8862=>"111101110",
  8863=>"111001110",
  8864=>"011001110",
  8865=>"010000111",
  8866=>"011101010",
  8867=>"110111110",
  8868=>"101110110",
  8869=>"100011000",
  8870=>"001100101",
  8871=>"000000001",
  8872=>"001100101",
  8873=>"010110000",
  8874=>"000001110",
  8875=>"001010110",
  8876=>"000011000",
  8877=>"011110000",
  8878=>"000001000",
  8879=>"001100000",
  8880=>"101010010",
  8881=>"110110000",
  8882=>"101111101",
  8883=>"110111000",
  8884=>"010110110",
  8885=>"110001100",
  8886=>"010101000",
  8887=>"111000011",
  8888=>"101100101",
  8889=>"111101110",
  8890=>"100010110",
  8891=>"111100010",
  8892=>"111001110",
  8893=>"001101101",
  8894=>"010100100",
  8895=>"000101001",
  8896=>"010011001",
  8897=>"000001101",
  8898=>"111010000",
  8899=>"100100010",
  8900=>"100111011",
  8901=>"011001011",
  8902=>"010010111",
  8903=>"000001111",
  8904=>"111110001",
  8905=>"001111100",
  8906=>"111110001",
  8907=>"000110000",
  8908=>"100100101",
  8909=>"010110110",
  8910=>"110110111",
  8911=>"000101110",
  8912=>"100100100",
  8913=>"101101000",
  8914=>"011001000",
  8915=>"011000100",
  8916=>"001110111",
  8917=>"011001000",
  8918=>"010000111",
  8919=>"111000111",
  8920=>"111000001",
  8921=>"010000100",
  8922=>"100111111",
  8923=>"011010000",
  8924=>"111011000",
  8925=>"000101010",
  8926=>"000011001",
  8927=>"000000001",
  8928=>"011001000",
  8929=>"011100110",
  8930=>"100011100",
  8931=>"001111110",
  8932=>"011010110",
  8933=>"101011101",
  8934=>"101101001",
  8935=>"011101001",
  8936=>"010010010",
  8937=>"100110101",
  8938=>"001110100",
  8939=>"010000000",
  8940=>"000111000",
  8941=>"111001111",
  8942=>"010100101",
  8943=>"101111010",
  8944=>"101010100",
  8945=>"000000110",
  8946=>"011010100",
  8947=>"000100111",
  8948=>"100010101",
  8949=>"111100110",
  8950=>"101110100",
  8951=>"011001010",
  8952=>"000000111",
  8953=>"010111000",
  8954=>"001100101",
  8955=>"011100000",
  8956=>"101001110",
  8957=>"010001110",
  8958=>"001001000",
  8959=>"000111001",
  8960=>"011001101",
  8961=>"101001110",
  8962=>"100111000",
  8963=>"111101111",
  8964=>"000000000",
  8965=>"010000111",
  8966=>"110101010",
  8967=>"111110111",
  8968=>"100010101",
  8969=>"111111100",
  8970=>"100100010",
  8971=>"111010011",
  8972=>"111100000",
  8973=>"000011010",
  8974=>"100011110",
  8975=>"000101110",
  8976=>"010100110",
  8977=>"111111010",
  8978=>"111111011",
  8979=>"110110000",
  8980=>"101110011",
  8981=>"011110000",
  8982=>"100001101",
  8983=>"000010010",
  8984=>"111001100",
  8985=>"001010000",
  8986=>"000101110",
  8987=>"100110110",
  8988=>"100100110",
  8989=>"011100000",
  8990=>"010111110",
  8991=>"101010011",
  8992=>"111011011",
  8993=>"000010100",
  8994=>"011010011",
  8995=>"111110110",
  8996=>"111000100",
  8997=>"000000000",
  8998=>"010000100",
  8999=>"111011111",
  9000=>"111000110",
  9001=>"110111000",
  9002=>"110010010",
  9003=>"111010000",
  9004=>"100101110",
  9005=>"010000101",
  9006=>"111111101",
  9007=>"010100110",
  9008=>"011101110",
  9009=>"011001110",
  9010=>"110111100",
  9011=>"100011001",
  9012=>"101101100",
  9013=>"001001011",
  9014=>"000000010",
  9015=>"111001101",
  9016=>"100100100",
  9017=>"010011001",
  9018=>"101000111",
  9019=>"000000001",
  9020=>"111101101",
  9021=>"001010010",
  9022=>"001010011",
  9023=>"101110101",
  9024=>"111010000",
  9025=>"000111011",
  9026=>"100010111",
  9027=>"000011001",
  9028=>"100010000",
  9029=>"011110111",
  9030=>"110101101",
  9031=>"001000001",
  9032=>"100101110",
  9033=>"110110110",
  9034=>"010101010",
  9035=>"110110101",
  9036=>"000111100",
  9037=>"100101000",
  9038=>"010000011",
  9039=>"100000110",
  9040=>"010010001",
  9041=>"011110100",
  9042=>"001101100",
  9043=>"010011000",
  9044=>"110111010",
  9045=>"011110111",
  9046=>"101101100",
  9047=>"111010000",
  9048=>"001100001",
  9049=>"010111001",
  9050=>"000101000",
  9051=>"010110010",
  9052=>"101111110",
  9053=>"000011100",
  9054=>"011101011",
  9055=>"000010000",
  9056=>"001010101",
  9057=>"100111011",
  9058=>"111011010",
  9059=>"101000000",
  9060=>"000011010",
  9061=>"001101111",
  9062=>"010111100",
  9063=>"001010000",
  9064=>"001111100",
  9065=>"111010111",
  9066=>"011010011",
  9067=>"011100001",
  9068=>"000011111",
  9069=>"000101110",
  9070=>"100101110",
  9071=>"001101111",
  9072=>"100011100",
  9073=>"101001000",
  9074=>"010010011",
  9075=>"110101110",
  9076=>"001000010",
  9077=>"000110001",
  9078=>"000101001",
  9079=>"101010101",
  9080=>"010000101",
  9081=>"101110010",
  9082=>"111111011",
  9083=>"010110011",
  9084=>"011011001",
  9085=>"000000101",
  9086=>"111110111",
  9087=>"111001000",
  9088=>"010111100",
  9089=>"000111001",
  9090=>"111011100",
  9091=>"101000110",
  9092=>"110010010",
  9093=>"000110011",
  9094=>"110100000",
  9095=>"110101011",
  9096=>"001101101",
  9097=>"000000001",
  9098=>"000001110",
  9099=>"111100011",
  9100=>"011000000",
  9101=>"000111101",
  9102=>"000110001",
  9103=>"101000111",
  9104=>"001110001",
  9105=>"000000101",
  9106=>"010010011",
  9107=>"101001100",
  9108=>"001110010",
  9109=>"011010000",
  9110=>"101010011",
  9111=>"111010111",
  9112=>"000000010",
  9113=>"100111100",
  9114=>"000100100",
  9115=>"101101010",
  9116=>"100110111",
  9117=>"001110010",
  9118=>"001010000",
  9119=>"010101110",
  9120=>"110000010",
  9121=>"010110100",
  9122=>"110011100",
  9123=>"010111101",
  9124=>"010000000",
  9125=>"110010011",
  9126=>"000000001",
  9127=>"011000001",
  9128=>"011001101",
  9129=>"111101101",
  9130=>"011111101",
  9131=>"000110110",
  9132=>"011010101",
  9133=>"000001001",
  9134=>"110100001",
  9135=>"011000111",
  9136=>"000000010",
  9137=>"111111110",
  9138=>"111010001",
  9139=>"100000000",
  9140=>"101011101",
  9141=>"011111000",
  9142=>"100110111",
  9143=>"001010001",
  9144=>"110011011",
  9145=>"111000111",
  9146=>"011110000",
  9147=>"000011001",
  9148=>"010111010",
  9149=>"000001111",
  9150=>"001010001",
  9151=>"000101110",
  9152=>"101001000",
  9153=>"011010010",
  9154=>"000001010",
  9155=>"010010111",
  9156=>"011010001",
  9157=>"111011011",
  9158=>"101100100",
  9159=>"001100000",
  9160=>"010101000",
  9161=>"110111110",
  9162=>"001011000",
  9163=>"110101000",
  9164=>"111001110",
  9165=>"111100011",
  9166=>"101110010",
  9167=>"010011010",
  9168=>"010111110",
  9169=>"111100001",
  9170=>"111110001",
  9171=>"011100110",
  9172=>"000100001",
  9173=>"100010011",
  9174=>"000001100",
  9175=>"010000101",
  9176=>"001110010",
  9177=>"011000111",
  9178=>"001000001",
  9179=>"000101101",
  9180=>"100011101",
  9181=>"010100001",
  9182=>"110100010",
  9183=>"111011011",
  9184=>"110111110",
  9185=>"010100000",
  9186=>"000110011",
  9187=>"010110001",
  9188=>"000011000",
  9189=>"111001101",
  9190=>"100110100",
  9191=>"100101110",
  9192=>"101001110",
  9193=>"001101011",
  9194=>"100100000",
  9195=>"001011110",
  9196=>"010111011",
  9197=>"000111110",
  9198=>"011001000",
  9199=>"110001000",
  9200=>"000000100",
  9201=>"111001111",
  9202=>"010111110",
  9203=>"100011101",
  9204=>"010001010",
  9205=>"100110101",
  9206=>"100111010",
  9207=>"110111111",
  9208=>"110111000",
  9209=>"001011000",
  9210=>"110100101",
  9211=>"111110110",
  9212=>"001011110",
  9213=>"001110011",
  9214=>"011101110",
  9215=>"011000001",
  9216=>"100001101",
  9217=>"010001100",
  9218=>"110111101",
  9219=>"100100001",
  9220=>"101100111",
  9221=>"101001010",
  9222=>"111101000",
  9223=>"000000111",
  9224=>"010111011",
  9225=>"001111010",
  9226=>"011001000",
  9227=>"101101000",
  9228=>"110110100",
  9229=>"011111010",
  9230=>"000110101",
  9231=>"010000001",
  9232=>"101110001",
  9233=>"011101110",
  9234=>"000001011",
  9235=>"000010100",
  9236=>"100000011",
  9237=>"011110111",
  9238=>"000001010",
  9239=>"101100110",
  9240=>"100100100",
  9241=>"110100101",
  9242=>"010111011",
  9243=>"101000011",
  9244=>"011111101",
  9245=>"011111010",
  9246=>"111101100",
  9247=>"010111100",
  9248=>"100000010",
  9249=>"111010000",
  9250=>"000000000",
  9251=>"100011111",
  9252=>"100100000",
  9253=>"111111010",
  9254=>"100010001",
  9255=>"011101000",
  9256=>"000001110",
  9257=>"100100100",
  9258=>"011011100",
  9259=>"100011111",
  9260=>"111001111",
  9261=>"110011100",
  9262=>"101101101",
  9263=>"010000000",
  9264=>"110111111",
  9265=>"111100000",
  9266=>"000110010",
  9267=>"011010011",
  9268=>"011000110",
  9269=>"101011001",
  9270=>"000100010",
  9271=>"000001111",
  9272=>"111111010",
  9273=>"010001110",
  9274=>"011000001",
  9275=>"010111000",
  9276=>"111110000",
  9277=>"010001010",
  9278=>"001110000",
  9279=>"101110001",
  9280=>"111011011",
  9281=>"011000001",
  9282=>"101111011",
  9283=>"000111010",
  9284=>"110110010",
  9285=>"100000000",
  9286=>"101000011",
  9287=>"000100111",
  9288=>"101111000",
  9289=>"010101111",
  9290=>"101001110",
  9291=>"011001011",
  9292=>"011110110",
  9293=>"001011100",
  9294=>"100101100",
  9295=>"001000010",
  9296=>"011000001",
  9297=>"100110111",
  9298=>"110111101",
  9299=>"100110100",
  9300=>"001011111",
  9301=>"000000101",
  9302=>"110001110",
  9303=>"000100010",
  9304=>"001010101",
  9305=>"101100110",
  9306=>"010111101",
  9307=>"010001001",
  9308=>"000010001",
  9309=>"100011111",
  9310=>"100101010",
  9311=>"110000000",
  9312=>"001100001",
  9313=>"101100101",
  9314=>"000111000",
  9315=>"001100010",
  9316=>"010010000",
  9317=>"101101111",
  9318=>"110000100",
  9319=>"100100110",
  9320=>"001010110",
  9321=>"111001110",
  9322=>"100001101",
  9323=>"111100100",
  9324=>"111110010",
  9325=>"001001000",
  9326=>"100011010",
  9327=>"100110111",
  9328=>"011000100",
  9329=>"100000010",
  9330=>"001000100",
  9331=>"011101101",
  9332=>"101000001",
  9333=>"110111101",
  9334=>"111011111",
  9335=>"110011000",
  9336=>"110000000",
  9337=>"110110110",
  9338=>"011011010",
  9339=>"000010110",
  9340=>"101101010",
  9341=>"000001001",
  9342=>"010101111",
  9343=>"000100000",
  9344=>"100111111",
  9345=>"100000010",
  9346=>"111010000",
  9347=>"101101010",
  9348=>"111011100",
  9349=>"001101100",
  9350=>"101000100",
  9351=>"100010101",
  9352=>"000111111",
  9353=>"001000111",
  9354=>"111000011",
  9355=>"000011010",
  9356=>"101000011",
  9357=>"110110010",
  9358=>"010001001",
  9359=>"110010001",
  9360=>"100000111",
  9361=>"101001001",
  9362=>"010101111",
  9363=>"001110101",
  9364=>"101111101",
  9365=>"001000001",
  9366=>"111110110",
  9367=>"000100010",
  9368=>"111110011",
  9369=>"101111100",
  9370=>"101101001",
  9371=>"111100010",
  9372=>"101100101",
  9373=>"000111010",
  9374=>"100111110",
  9375=>"010000101",
  9376=>"000100000",
  9377=>"100100001",
  9378=>"010010001",
  9379=>"100000010",
  9380=>"111111111",
  9381=>"001111011",
  9382=>"101001011",
  9383=>"101011010",
  9384=>"011010010",
  9385=>"110010001",
  9386=>"110101111",
  9387=>"000000111",
  9388=>"010000011",
  9389=>"011011010",
  9390=>"001101000",
  9391=>"001010001",
  9392=>"111001001",
  9393=>"111001111",
  9394=>"000011010",
  9395=>"100110100",
  9396=>"011010000",
  9397=>"110101110",
  9398=>"100001110",
  9399=>"111011110",
  9400=>"001100011",
  9401=>"011101111",
  9402=>"001100100",
  9403=>"001100000",
  9404=>"110100001",
  9405=>"010000000",
  9406=>"111101011",
  9407=>"100110001",
  9408=>"011101010",
  9409=>"100110101",
  9410=>"000001001",
  9411=>"110110111",
  9412=>"000111111",
  9413=>"101101001",
  9414=>"010011000",
  9415=>"110100111",
  9416=>"100000011",
  9417=>"100100101",
  9418=>"010111101",
  9419=>"001011000",
  9420=>"111111000",
  9421=>"101010010",
  9422=>"001011111",
  9423=>"100111111",
  9424=>"110100010",
  9425=>"100000101",
  9426=>"100000100",
  9427=>"110110101",
  9428=>"110110011",
  9429=>"101010110",
  9430=>"111000111",
  9431=>"100100001",
  9432=>"010001011",
  9433=>"110101010",
  9434=>"101110100",
  9435=>"101111101",
  9436=>"001011000",
  9437=>"111011101",
  9438=>"010101010",
  9439=>"111101111",
  9440=>"010010111",
  9441=>"110010001",
  9442=>"111001110",
  9443=>"100010011",
  9444=>"111010110",
  9445=>"010001110",
  9446=>"100101000",
  9447=>"010010011",
  9448=>"010110111",
  9449=>"100001011",
  9450=>"110101001",
  9451=>"010111010",
  9452=>"010101001",
  9453=>"110000100",
  9454=>"111010110",
  9455=>"111111100",
  9456=>"011001110",
  9457=>"011000000",
  9458=>"111100011",
  9459=>"111000011",
  9460=>"110110000",
  9461=>"101110100",
  9462=>"110110011",
  9463=>"010110010",
  9464=>"000111011",
  9465=>"100111011",
  9466=>"011001110",
  9467=>"101101001",
  9468=>"001111111",
  9469=>"010000010",
  9470=>"100000001",
  9471=>"011110001",
  9472=>"100110101",
  9473=>"000100101",
  9474=>"101001001",
  9475=>"000000111",
  9476=>"111010110",
  9477=>"010011001",
  9478=>"001000010",
  9479=>"100111101",
  9480=>"101111111",
  9481=>"110100100",
  9482=>"011011101",
  9483=>"011000101",
  9484=>"110011011",
  9485=>"100001110",
  9486=>"001110111",
  9487=>"100010100",
  9488=>"011010011",
  9489=>"001111010",
  9490=>"110000110",
  9491=>"110011000",
  9492=>"010110000",
  9493=>"011001110",
  9494=>"110110000",
  9495=>"001110100",
  9496=>"011110101",
  9497=>"010100100",
  9498=>"010111010",
  9499=>"111100010",
  9500=>"110010101",
  9501=>"010011101",
  9502=>"000000110",
  9503=>"010011001",
  9504=>"100101001",
  9505=>"010011011",
  9506=>"110110110",
  9507=>"100010011",
  9508=>"011101000",
  9509=>"110001111",
  9510=>"011001101",
  9511=>"100110010",
  9512=>"111000010",
  9513=>"010111100",
  9514=>"011010101",
  9515=>"010000100",
  9516=>"010011111",
  9517=>"001111000",
  9518=>"010011001",
  9519=>"100100011",
  9520=>"001100100",
  9521=>"000011111",
  9522=>"000011101",
  9523=>"011111110",
  9524=>"100011000",
  9525=>"001111000",
  9526=>"000001100",
  9527=>"010010111",
  9528=>"000100001",
  9529=>"110010010",
  9530=>"010010000",
  9531=>"111100000",
  9532=>"101000110",
  9533=>"111011101",
  9534=>"111110100",
  9535=>"111111001",
  9536=>"110100101",
  9537=>"010001001",
  9538=>"101000110",
  9539=>"110101111",
  9540=>"100101100",
  9541=>"101011000",
  9542=>"111111000",
  9543=>"110111011",
  9544=>"100000010",
  9545=>"100110111",
  9546=>"010111111",
  9547=>"010111000",
  9548=>"001100001",
  9549=>"111101111",
  9550=>"000000100",
  9551=>"001011001",
  9552=>"110001111",
  9553=>"101001100",
  9554=>"010001010",
  9555=>"101110100",
  9556=>"000111011",
  9557=>"110010001",
  9558=>"001101011",
  9559=>"011110101",
  9560=>"101100000",
  9561=>"010010101",
  9562=>"000000100",
  9563=>"100100011",
  9564=>"110100101",
  9565=>"010100001",
  9566=>"100100110",
  9567=>"100000111",
  9568=>"111101100",
  9569=>"101101100",
  9570=>"000101011",
  9571=>"001010000",
  9572=>"111011100",
  9573=>"110110111",
  9574=>"011010100",
  9575=>"000000001",
  9576=>"010001100",
  9577=>"111100000",
  9578=>"100101111",
  9579=>"010110101",
  9580=>"110110101",
  9581=>"010101101",
  9582=>"110100110",
  9583=>"010101011",
  9584=>"101111110",
  9585=>"000000110",
  9586=>"110111000",
  9587=>"111101011",
  9588=>"000011101",
  9589=>"110000000",
  9590=>"001000110",
  9591=>"101100110",
  9592=>"000101000",
  9593=>"110111001",
  9594=>"001001010",
  9595=>"000011111",
  9596=>"001110110",
  9597=>"000010001",
  9598=>"100011010",
  9599=>"100110000",
  9600=>"000111110",
  9601=>"010111010",
  9602=>"100011001",
  9603=>"101011000",
  9604=>"100100001",
  9605=>"101000110",
  9606=>"011110111",
  9607=>"010100100",
  9608=>"101100101",
  9609=>"011001010",
  9610=>"110011100",
  9611=>"100001100",
  9612=>"000100000",
  9613=>"011100101",
  9614=>"100000111",
  9615=>"101101011",
  9616=>"001010011",
  9617=>"100100111",
  9618=>"000101010",
  9619=>"010101100",
  9620=>"001110001",
  9621=>"000001101",
  9622=>"100100001",
  9623=>"110001011",
  9624=>"110000101",
  9625=>"101100001",
  9626=>"010100110",
  9627=>"010011010",
  9628=>"000101100",
  9629=>"011010111",
  9630=>"100110111",
  9631=>"111001100",
  9632=>"010000000",
  9633=>"111110111",
  9634=>"001001101",
  9635=>"111001110",
  9636=>"000010110",
  9637=>"111100000",
  9638=>"101100010",
  9639=>"011010100",
  9640=>"101001110",
  9641=>"101000011",
  9642=>"101010000",
  9643=>"111111110",
  9644=>"110110011",
  9645=>"101100101",
  9646=>"011101100",
  9647=>"001110011",
  9648=>"001101001",
  9649=>"010011110",
  9650=>"000101101",
  9651=>"010011111",
  9652=>"011000000",
  9653=>"000010011",
  9654=>"010110000",
  9655=>"111001111",
  9656=>"000000000",
  9657=>"110100110",
  9658=>"000000111",
  9659=>"010010000",
  9660=>"101001111",
  9661=>"111111110",
  9662=>"010100000",
  9663=>"111011011",
  9664=>"111000010",
  9665=>"010110010",
  9666=>"001011100",
  9667=>"100101111",
  9668=>"000000100",
  9669=>"100000000",
  9670=>"100001010",
  9671=>"001101010",
  9672=>"110110101",
  9673=>"001001101",
  9674=>"111111110",
  9675=>"010101001",
  9676=>"111100100",
  9677=>"101010110",
  9678=>"101000000",
  9679=>"001110100",
  9680=>"101010101",
  9681=>"001111111",
  9682=>"100000101",
  9683=>"000101110",
  9684=>"100111000",
  9685=>"110110101",
  9686=>"000110010",
  9687=>"101100000",
  9688=>"100000011",
  9689=>"110110110",
  9690=>"001110111",
  9691=>"101001000",
  9692=>"010011011",
  9693=>"111111101",
  9694=>"110011111",
  9695=>"110101011",
  9696=>"011110111",
  9697=>"000000111",
  9698=>"001101101",
  9699=>"101101000",
  9700=>"110100100",
  9701=>"011000111",
  9702=>"011000100",
  9703=>"011100110",
  9704=>"011111111",
  9705=>"101010111",
  9706=>"110001111",
  9707=>"110010001",
  9708=>"110001000",
  9709=>"010000000",
  9710=>"110011100",
  9711=>"100010011",
  9712=>"101010111",
  9713=>"111111101",
  9714=>"111110000",
  9715=>"000001100",
  9716=>"000110110",
  9717=>"010100100",
  9718=>"100111000",
  9719=>"111101111",
  9720=>"000101100",
  9721=>"110101011",
  9722=>"011011101",
  9723=>"100000011",
  9724=>"001110111",
  9725=>"010110000",
  9726=>"110111110",
  9727=>"000000010",
  9728=>"110111001",
  9729=>"111111100",
  9730=>"001100111",
  9731=>"001100110",
  9732=>"101110110",
  9733=>"000111101",
  9734=>"110101000",
  9735=>"110110000",
  9736=>"001100011",
  9737=>"101011100",
  9738=>"110001011",
  9739=>"110010101",
  9740=>"000111101",
  9741=>"000001000",
  9742=>"001001001",
  9743=>"101001011",
  9744=>"000111110",
  9745=>"101111110",
  9746=>"100011111",
  9747=>"111010101",
  9748=>"000001010",
  9749=>"010000101",
  9750=>"001011101",
  9751=>"110000111",
  9752=>"000010000",
  9753=>"011010101",
  9754=>"111001011",
  9755=>"110000101",
  9756=>"101011011",
  9757=>"000000001",
  9758=>"111100010",
  9759=>"011010101",
  9760=>"101010110",
  9761=>"001111000",
  9762=>"101111010",
  9763=>"110001100",
  9764=>"000000010",
  9765=>"101010101",
  9766=>"011100111",
  9767=>"111110100",
  9768=>"110000100",
  9769=>"001010111",
  9770=>"011100110",
  9771=>"100001000",
  9772=>"111100000",
  9773=>"111110010",
  9774=>"100101101",
  9775=>"111101001",
  9776=>"000101001",
  9777=>"101111001",
  9778=>"100101111",
  9779=>"001010000",
  9780=>"010001101",
  9781=>"110111101",
  9782=>"000111011",
  9783=>"001000101",
  9784=>"000011001",
  9785=>"101000100",
  9786=>"001101100",
  9787=>"011001011",
  9788=>"110100111",
  9789=>"001011011",
  9790=>"001011110",
  9791=>"101011110",
  9792=>"101100000",
  9793=>"111010000",
  9794=>"000010100",
  9795=>"011011000",
  9796=>"101100100",
  9797=>"011011111",
  9798=>"110001111",
  9799=>"101010001",
  9800=>"010001101",
  9801=>"010010111",
  9802=>"010010001",
  9803=>"000110110",
  9804=>"111001110",
  9805=>"000111001",
  9806=>"001001000",
  9807=>"101010100",
  9808=>"111010111",
  9809=>"011111100",
  9810=>"110001111",
  9811=>"001001001",
  9812=>"010011011",
  9813=>"000100011",
  9814=>"100101011",
  9815=>"010101011",
  9816=>"010011001",
  9817=>"010000101",
  9818=>"010110010",
  9819=>"111010011",
  9820=>"100111110",
  9821=>"100001100",
  9822=>"001100110",
  9823=>"011110101",
  9824=>"100110111",
  9825=>"101111110",
  9826=>"101001000",
  9827=>"001110111",
  9828=>"001110010",
  9829=>"000001000",
  9830=>"111011101",
  9831=>"100110100",
  9832=>"110011100",
  9833=>"101100101",
  9834=>"010010011",
  9835=>"101001001",
  9836=>"011010110",
  9837=>"000110110",
  9838=>"011100100",
  9839=>"110010000",
  9840=>"000101000",
  9841=>"000101000",
  9842=>"001011000",
  9843=>"101111001",
  9844=>"111001010",
  9845=>"010100110",
  9846=>"010100010",
  9847=>"111110010",
  9848=>"001001101",
  9849=>"010001010",
  9850=>"101010100",
  9851=>"111011100",
  9852=>"111000101",
  9853=>"010010110",
  9854=>"111110010",
  9855=>"011101001",
  9856=>"111011100",
  9857=>"110001111",
  9858=>"000100111",
  9859=>"001001110",
  9860=>"110010001",
  9861=>"010010101",
  9862=>"101011111",
  9863=>"010110110",
  9864=>"010100101",
  9865=>"010110010",
  9866=>"011101010",
  9867=>"011111101",
  9868=>"110100011",
  9869=>"001000011",
  9870=>"000001100",
  9871=>"011110001",
  9872=>"111010111",
  9873=>"111111110",
  9874=>"100100001",
  9875=>"110001101",
  9876=>"100110000",
  9877=>"000011010",
  9878=>"101010001",
  9879=>"001110011",
  9880=>"100110110",
  9881=>"001101011",
  9882=>"100000000",
  9883=>"010010001",
  9884=>"000110000",
  9885=>"101001100",
  9886=>"111111111",
  9887=>"010100000",
  9888=>"100101011",
  9889=>"110111000",
  9890=>"111111010",
  9891=>"010101101",
  9892=>"100011001",
  9893=>"101100101",
  9894=>"101111000",
  9895=>"100101000",
  9896=>"011111111",
  9897=>"010000000",
  9898=>"001000000",
  9899=>"111010010",
  9900=>"100000001",
  9901=>"101110111",
  9902=>"101111001",
  9903=>"000101110",
  9904=>"000000001",
  9905=>"111001000",
  9906=>"101011010",
  9907=>"011100000",
  9908=>"010010101",
  9909=>"001001101",
  9910=>"111100110",
  9911=>"110101001",
  9912=>"110011101",
  9913=>"100110010",
  9914=>"011101001",
  9915=>"011101000",
  9916=>"100111110",
  9917=>"010001000",
  9918=>"111010010",
  9919=>"011011111",
  9920=>"011111111",
  9921=>"010110100",
  9922=>"111011101",
  9923=>"110111100",
  9924=>"010001011",
  9925=>"111111010",
  9926=>"000110110",
  9927=>"101110111",
  9928=>"101110001",
  9929=>"010111011",
  9930=>"110101001",
  9931=>"101000010",
  9932=>"000001101",
  9933=>"000011110",
  9934=>"010010001",
  9935=>"110001100",
  9936=>"010001001",
  9937=>"001110110",
  9938=>"000111011",
  9939=>"110000101",
  9940=>"100100000",
  9941=>"111101010",
  9942=>"000001001",
  9943=>"101011111",
  9944=>"011001001",
  9945=>"101011011",
  9946=>"000010100",
  9947=>"011010011",
  9948=>"110111101",
  9949=>"011011100",
  9950=>"110111001",
  9951=>"100110110",
  9952=>"010101011",
  9953=>"111001001",
  9954=>"001001111",
  9955=>"100010000",
  9956=>"011101110",
  9957=>"010111111",
  9958=>"001100001",
  9959=>"000110111",
  9960=>"000010010",
  9961=>"101011011",
  9962=>"010011110",
  9963=>"100011010",
  9964=>"011110011",
  9965=>"000001011",
  9966=>"101011000",
  9967=>"101111101",
  9968=>"110111110",
  9969=>"101110010",
  9970=>"011001000",
  9971=>"011110000",
  9972=>"100110111",
  9973=>"110000011",
  9974=>"001100001",
  9975=>"100100011",
  9976=>"010000111",
  9977=>"110101011",
  9978=>"011000000",
  9979=>"000001110",
  9980=>"001101011",
  9981=>"010000000",
  9982=>"011111100",
  9983=>"011110000",
  9984=>"011111001",
  9985=>"010101011",
  9986=>"101000110",
  9987=>"101000001",
  9988=>"110111011",
  9989=>"011110010",
  9990=>"111110001",
  9991=>"001000110",
  9992=>"111001110",
  9993=>"110010100",
  9994=>"110000001",
  9995=>"110010010",
  9996=>"111001100",
  9997=>"011011111",
  9998=>"001101100",
  9999=>"010011000",
  10000=>"100001011",
  10001=>"111000010",
  10002=>"011110101",
  10003=>"100000001",
  10004=>"111000000",
  10005=>"010110010",
  10006=>"111101101",
  10007=>"100111001",
  10008=>"100100010",
  10009=>"101110000",
  10010=>"110110001",
  10011=>"110100000",
  10012=>"010000011",
  10013=>"001101011",
  10014=>"000011110",
  10015=>"110001011",
  10016=>"001011000",
  10017=>"110110110",
  10018=>"101000011",
  10019=>"010001000",
  10020=>"001000011",
  10021=>"111110011",
  10022=>"001000101",
  10023=>"001000110",
  10024=>"011000010",
  10025=>"100100000",
  10026=>"101011001",
  10027=>"000101000",
  10028=>"101110111",
  10029=>"010000110",
  10030=>"111001101",
  10031=>"100110110",
  10032=>"001000011",
  10033=>"110010101",
  10034=>"001110110",
  10035=>"001110011",
  10036=>"111000100",
  10037=>"100100000",
  10038=>"101100101",
  10039=>"100010001",
  10040=>"100001111",
  10041=>"000010011",
  10042=>"001000110",
  10043=>"000001101",
  10044=>"010000001",
  10045=>"100001001",
  10046=>"001110000",
  10047=>"010000000",
  10048=>"111100000",
  10049=>"011100100",
  10050=>"110100100",
  10051=>"001110111",
  10052=>"000101101",
  10053=>"111010111",
  10054=>"101001001",
  10055=>"111011111",
  10056=>"001001000",
  10057=>"011110010",
  10058=>"010100011",
  10059=>"001111101",
  10060=>"010111101",
  10061=>"010101010",
  10062=>"000111000",
  10063=>"011101010",
  10064=>"101111111",
  10065=>"000111110",
  10066=>"001100101",
  10067=>"000001010",
  10068=>"101111110",
  10069=>"101011110",
  10070=>"010100110",
  10071=>"011111001",
  10072=>"100100100",
  10073=>"110100011",
  10074=>"000110101",
  10075=>"110000000",
  10076=>"101111011",
  10077=>"110010000",
  10078=>"101010111",
  10079=>"100010000",
  10080=>"111000010",
  10081=>"000010100",
  10082=>"011001111",
  10083=>"000101000",
  10084=>"001101100",
  10085=>"011010101",
  10086=>"110000110",
  10087=>"001011101",
  10088=>"110110110",
  10089=>"110011000",
  10090=>"011100101",
  10091=>"001111111",
  10092=>"000011000",
  10093=>"000000000",
  10094=>"111111111",
  10095=>"011011101",
  10096=>"010111101",
  10097=>"010011101",
  10098=>"110100001",
  10099=>"001110101",
  10100=>"101101110",
  10101=>"100000110",
  10102=>"110101111",
  10103=>"110101101",
  10104=>"011001110",
  10105=>"101101111",
  10106=>"101101110",
  10107=>"000100011",
  10108=>"110111111",
  10109=>"111100110",
  10110=>"111111110",
  10111=>"001100100",
  10112=>"011001011",
  10113=>"001000011",
  10114=>"011011000",
  10115=>"000111100",
  10116=>"001101110",
  10117=>"110110001",
  10118=>"101011000",
  10119=>"110011110",
  10120=>"101011001",
  10121=>"011010111",
  10122=>"010111011",
  10123=>"111110111",
  10124=>"000111111",
  10125=>"110000110",
  10126=>"000000111",
  10127=>"010110110",
  10128=>"100001010",
  10129=>"100110000",
  10130=>"010111011",
  10131=>"101110010",
  10132=>"100100110",
  10133=>"000100100",
  10134=>"101101001",
  10135=>"101101011",
  10136=>"011010100",
  10137=>"100110000",
  10138=>"001010110",
  10139=>"010011101",
  10140=>"100110110",
  10141=>"100110111",
  10142=>"101110111",
  10143=>"111101101",
  10144=>"101110001",
  10145=>"100101100",
  10146=>"100111001",
  10147=>"111010001",
  10148=>"001100010",
  10149=>"110010010",
  10150=>"101110101",
  10151=>"001001000",
  10152=>"011011011",
  10153=>"101001111",
  10154=>"101100111",
  10155=>"011011010",
  10156=>"010000110",
  10157=>"110001001",
  10158=>"010000000",
  10159=>"111001000",
  10160=>"011100101",
  10161=>"010000100",
  10162=>"001001101",
  10163=>"100111100",
  10164=>"001010011",
  10165=>"001100000",
  10166=>"000011011",
  10167=>"000010111",
  10168=>"110100111",
  10169=>"001101001",
  10170=>"111011100",
  10171=>"110010000",
  10172=>"111010110",
  10173=>"111110000",
  10174=>"110010111",
  10175=>"100001001",
  10176=>"001000011",
  10177=>"001101110",
  10178=>"001010000",
  10179=>"001000111",
  10180=>"100010001",
  10181=>"000101101",
  10182=>"110011001",
  10183=>"010111000",
  10184=>"101100110",
  10185=>"101000111",
  10186=>"011100000",
  10187=>"111011100",
  10188=>"000010011",
  10189=>"100111110",
  10190=>"010000001",
  10191=>"101000011",
  10192=>"000111110",
  10193=>"101100010",
  10194=>"111110111",
  10195=>"110011010",
  10196=>"111000100",
  10197=>"011100011",
  10198=>"010101001",
  10199=>"101110101",
  10200=>"001001010",
  10201=>"100111100",
  10202=>"110100000",
  10203=>"000000011",
  10204=>"010001010",
  10205=>"010010110",
  10206=>"001100100",
  10207=>"011011000",
  10208=>"100000011",
  10209=>"111011100",
  10210=>"100000001",
  10211=>"110111010",
  10212=>"000001100",
  10213=>"111111111",
  10214=>"100110110",
  10215=>"110100100",
  10216=>"111101010",
  10217=>"110110010",
  10218=>"010100100",
  10219=>"000110010",
  10220=>"000100111",
  10221=>"001110100",
  10222=>"111011100",
  10223=>"101011101",
  10224=>"101011101",
  10225=>"011010110",
  10226=>"001101011",
  10227=>"011100111",
  10228=>"111001010",
  10229=>"110101001",
  10230=>"110111110",
  10231=>"001001010",
  10232=>"110000100",
  10233=>"011101001",
  10234=>"111000001",
  10235=>"100111000",
  10236=>"010010010",
  10237=>"011111101",
  10238=>"100000100",
  10239=>"100110110",
  10240=>"101001011",
  10241=>"101100110",
  10242=>"001011110",
  10243=>"100100110",
  10244=>"011011011",
  10245=>"011111011",
  10246=>"001001000",
  10247=>"011000110",
  10248=>"011000100",
  10249=>"101100001",
  10250=>"001001111",
  10251=>"001110101",
  10252=>"001010010",
  10253=>"101010010",
  10254=>"011100011",
  10255=>"110110010",
  10256=>"001010011",
  10257=>"010100100",
  10258=>"100111100",
  10259=>"010111001",
  10260=>"111001100",
  10261=>"110110010",
  10262=>"100010101",
  10263=>"010011011",
  10264=>"110101111",
  10265=>"000000110",
  10266=>"000100110",
  10267=>"111111101",
  10268=>"001001010",
  10269=>"111010011",
  10270=>"111111100",
  10271=>"111101000",
  10272=>"010101001",
  10273=>"011010101",
  10274=>"101111001",
  10275=>"111010001",
  10276=>"000101111",
  10277=>"100010000",
  10278=>"110010010",
  10279=>"110001000",
  10280=>"011100111",
  10281=>"001110011",
  10282=>"001011111",
  10283=>"111100011",
  10284=>"000010100",
  10285=>"010000111",
  10286=>"011000010",
  10287=>"011111010",
  10288=>"111100100",
  10289=>"000111111",
  10290=>"100100101",
  10291=>"011101001",
  10292=>"100000101",
  10293=>"011001000",
  10294=>"100110000",
  10295=>"011111000",
  10296=>"000011110",
  10297=>"101001101",
  10298=>"110110111",
  10299=>"010100101",
  10300=>"100011101",
  10301=>"011000000",
  10302=>"010000110",
  10303=>"010110010",
  10304=>"000111110",
  10305=>"000010101",
  10306=>"110100100",
  10307=>"000000100",
  10308=>"000001110",
  10309=>"000100010",
  10310=>"010111100",
  10311=>"111111101",
  10312=>"110101101",
  10313=>"000000010",
  10314=>"010000111",
  10315=>"010101011",
  10316=>"001000010",
  10317=>"000100011",
  10318=>"110010010",
  10319=>"001000101",
  10320=>"001000101",
  10321=>"110011101",
  10322=>"100110110",
  10323=>"101100010",
  10324=>"001101001",
  10325=>"100111110",
  10326=>"101010110",
  10327=>"011100000",
  10328=>"000010011",
  10329=>"111101101",
  10330=>"000000110",
  10331=>"001100011",
  10332=>"000001110",
  10333=>"100100000",
  10334=>"000111011",
  10335=>"110001101",
  10336=>"110000000",
  10337=>"101000000",
  10338=>"111111011",
  10339=>"111111010",
  10340=>"010110101",
  10341=>"101111110",
  10342=>"110001011",
  10343=>"110010001",
  10344=>"011010011",
  10345=>"111100001",
  10346=>"100010110",
  10347=>"111001000",
  10348=>"000011111",
  10349=>"110011001",
  10350=>"110011001",
  10351=>"111010011",
  10352=>"001011110",
  10353=>"000011001",
  10354=>"011101100",
  10355=>"011010111",
  10356=>"111111111",
  10357=>"101000000",
  10358=>"100100101",
  10359=>"110101010",
  10360=>"010100010",
  10361=>"111110001",
  10362=>"000110011",
  10363=>"001111101",
  10364=>"010000111",
  10365=>"000100100",
  10366=>"011001111",
  10367=>"001000110",
  10368=>"111101100",
  10369=>"011001001",
  10370=>"100001111",
  10371=>"001101001",
  10372=>"110011100",
  10373=>"000101010",
  10374=>"101110001",
  10375=>"011010010",
  10376=>"011001101",
  10377=>"000011010",
  10378=>"100011010",
  10379=>"100001111",
  10380=>"000000100",
  10381=>"111010001",
  10382=>"100010111",
  10383=>"110110101",
  10384=>"101110100",
  10385=>"100000101",
  10386=>"001100000",
  10387=>"111001101",
  10388=>"000011011",
  10389=>"000000101",
  10390=>"100101001",
  10391=>"100000110",
  10392=>"011011100",
  10393=>"110101101",
  10394=>"110010110",
  10395=>"011000101",
  10396=>"011111110",
  10397=>"111101110",
  10398=>"110010110",
  10399=>"111110100",
  10400=>"110101100",
  10401=>"101001100",
  10402=>"110111001",
  10403=>"110000000",
  10404=>"100010110",
  10405=>"011101110",
  10406=>"000100000",
  10407=>"111101101",
  10408=>"111100110",
  10409=>"011010010",
  10410=>"111010001",
  10411=>"000111111",
  10412=>"001100100",
  10413=>"100011101",
  10414=>"001110001",
  10415=>"110110000",
  10416=>"001101111",
  10417=>"100000000",
  10418=>"100000111",
  10419=>"000000110",
  10420=>"111010001",
  10421=>"110100011",
  10422=>"100101011",
  10423=>"101011000",
  10424=>"011100001",
  10425=>"110101010",
  10426=>"101100100",
  10427=>"001100101",
  10428=>"000101011",
  10429=>"100101111",
  10430=>"010101011",
  10431=>"110011011",
  10432=>"011111110",
  10433=>"110101111",
  10434=>"011000000",
  10435=>"101011001",
  10436=>"001110101",
  10437=>"100001011",
  10438=>"010100101",
  10439=>"110101001",
  10440=>"111000010",
  10441=>"011000011",
  10442=>"110100111",
  10443=>"111000011",
  10444=>"001000011",
  10445=>"010000100",
  10446=>"101111000",
  10447=>"100110011",
  10448=>"010000111",
  10449=>"110010000",
  10450=>"100000001",
  10451=>"101010011",
  10452=>"011000001",
  10453=>"101110001",
  10454=>"101000001",
  10455=>"111000100",
  10456=>"111101011",
  10457=>"101010110",
  10458=>"011010110",
  10459=>"000101000",
  10460=>"010100100",
  10461=>"001101000",
  10462=>"001100001",
  10463=>"011010011",
  10464=>"001100111",
  10465=>"011000011",
  10466=>"011010010",
  10467=>"100001001",
  10468=>"011101110",
  10469=>"110101001",
  10470=>"111101001",
  10471=>"001110110",
  10472=>"101100110",
  10473=>"101010010",
  10474=>"001101000",
  10475=>"111010111",
  10476=>"100010000",
  10477=>"000010111",
  10478=>"001111100",
  10479=>"110011000",
  10480=>"000111101",
  10481=>"010100010",
  10482=>"001101110",
  10483=>"110101000",
  10484=>"001110000",
  10485=>"010100111",
  10486=>"000111010",
  10487=>"110111010",
  10488=>"011101110",
  10489=>"011110010",
  10490=>"111000110",
  10491=>"111010000",
  10492=>"001011111",
  10493=>"111101100",
  10494=>"011001110",
  10495=>"011111000",
  10496=>"010101000",
  10497=>"001001001",
  10498=>"101111001",
  10499=>"111100001",
  10500=>"000010011",
  10501=>"110111010",
  10502=>"010010111",
  10503=>"001001000",
  10504=>"010100011",
  10505=>"010110111",
  10506=>"000000001",
  10507=>"010101011",
  10508=>"011010100",
  10509=>"011000111",
  10510=>"010000010",
  10511=>"110101101",
  10512=>"011001111",
  10513=>"101111111",
  10514=>"111110000",
  10515=>"000111010",
  10516=>"001100101",
  10517=>"010110111",
  10518=>"011111100",
  10519=>"110011111",
  10520=>"101101100",
  10521=>"011101110",
  10522=>"010011010",
  10523=>"101100100",
  10524=>"010110110",
  10525=>"000100100",
  10526=>"101010010",
  10527=>"000110010",
  10528=>"110111001",
  10529=>"101110100",
  10530=>"001111100",
  10531=>"101100011",
  10532=>"111100110",
  10533=>"110011000",
  10534=>"010001000",
  10535=>"001101110",
  10536=>"100101000",
  10537=>"101110101",
  10538=>"101100011",
  10539=>"000101000",
  10540=>"101011101",
  10541=>"101011011",
  10542=>"111110011",
  10543=>"000000110",
  10544=>"110110001",
  10545=>"101110110",
  10546=>"011100111",
  10547=>"000001000",
  10548=>"111111010",
  10549=>"101101001",
  10550=>"110001101",
  10551=>"110000101",
  10552=>"111011000",
  10553=>"110110110",
  10554=>"111011010",
  10555=>"110000101",
  10556=>"100001011",
  10557=>"110000111",
  10558=>"010000011",
  10559=>"010001000",
  10560=>"010111010",
  10561=>"001000001",
  10562=>"111100101",
  10563=>"110110110",
  10564=>"111100000",
  10565=>"110110001",
  10566=>"000011101",
  10567=>"001010000",
  10568=>"010010001",
  10569=>"100000000",
  10570=>"000011110",
  10571=>"010110000",
  10572=>"010000010",
  10573=>"101101010",
  10574=>"110011101",
  10575=>"001010110",
  10576=>"100100101",
  10577=>"010000101",
  10578=>"001000101",
  10579=>"101000001",
  10580=>"110011010",
  10581=>"100010000",
  10582=>"011010010",
  10583=>"110101101",
  10584=>"010100110",
  10585=>"000010100",
  10586=>"111101010",
  10587=>"101110111",
  10588=>"101101010",
  10589=>"101110111",
  10590=>"110111110",
  10591=>"011110010",
  10592=>"010001001",
  10593=>"010100100",
  10594=>"011110010",
  10595=>"101001111",
  10596=>"011011111",
  10597=>"100000010",
  10598=>"011100010",
  10599=>"000001001",
  10600=>"110110100",
  10601=>"000001101",
  10602=>"000111111",
  10603=>"110000110",
  10604=>"110011010",
  10605=>"110111000",
  10606=>"011100111",
  10607=>"000100100",
  10608=>"001001001",
  10609=>"000011000",
  10610=>"111001110",
  10611=>"111111100",
  10612=>"111011000",
  10613=>"000011111",
  10614=>"101000110",
  10615=>"111100000",
  10616=>"100001010",
  10617=>"110110010",
  10618=>"110001001",
  10619=>"100101000",
  10620=>"100001001",
  10621=>"111010010",
  10622=>"110101101",
  10623=>"000000101",
  10624=>"100011010",
  10625=>"000100011",
  10626=>"111100111",
  10627=>"000000000",
  10628=>"010100110",
  10629=>"010101101",
  10630=>"000111001",
  10631=>"100110000",
  10632=>"011111110",
  10633=>"000000000",
  10634=>"000011010",
  10635=>"111100010",
  10636=>"000000011",
  10637=>"101100001",
  10638=>"111111101",
  10639=>"111011010",
  10640=>"001001100",
  10641=>"000010111",
  10642=>"101010101",
  10643=>"001011110",
  10644=>"110111010",
  10645=>"010111000",
  10646=>"100111010",
  10647=>"011010100",
  10648=>"010111111",
  10649=>"101011111",
  10650=>"010000011",
  10651=>"110011101",
  10652=>"010010110",
  10653=>"011110001",
  10654=>"001010001",
  10655=>"011111110",
  10656=>"111101101",
  10657=>"001111011",
  10658=>"000000000",
  10659=>"111011110",
  10660=>"000001101",
  10661=>"111000111",
  10662=>"011100010",
  10663=>"000010001",
  10664=>"001111101",
  10665=>"010010111",
  10666=>"101000000",
  10667=>"010001000",
  10668=>"111101000",
  10669=>"001110000",
  10670=>"111000111",
  10671=>"000100111",
  10672=>"001110101",
  10673=>"110101011",
  10674=>"000001001",
  10675=>"101001001",
  10676=>"011111001",
  10677=>"110111110",
  10678=>"101000011",
  10679=>"010110110",
  10680=>"011001111",
  10681=>"010001010",
  10682=>"000001101",
  10683=>"110000011",
  10684=>"000110101",
  10685=>"111001010",
  10686=>"011110010",
  10687=>"110011100",
  10688=>"001110000",
  10689=>"000101000",
  10690=>"110000001",
  10691=>"000000100",
  10692=>"110001110",
  10693=>"100111000",
  10694=>"011101010",
  10695=>"110110010",
  10696=>"100110010",
  10697=>"010001100",
  10698=>"100011110",
  10699=>"111010000",
  10700=>"111111111",
  10701=>"111101011",
  10702=>"001011010",
  10703=>"101110000",
  10704=>"001010111",
  10705=>"100110010",
  10706=>"101001011",
  10707=>"100110010",
  10708=>"010111001",
  10709=>"011010000",
  10710=>"000110110",
  10711=>"000101001",
  10712=>"100111110",
  10713=>"101101101",
  10714=>"011101100",
  10715=>"101000001",
  10716=>"011101101",
  10717=>"101011110",
  10718=>"100001100",
  10719=>"110101101",
  10720=>"111100010",
  10721=>"101101001",
  10722=>"000010101",
  10723=>"001011101",
  10724=>"000001111",
  10725=>"000000011",
  10726=>"100011110",
  10727=>"111111000",
  10728=>"111100111",
  10729=>"100110011",
  10730=>"110010101",
  10731=>"100101110",
  10732=>"001100111",
  10733=>"011010111",
  10734=>"110110100",
  10735=>"100000000",
  10736=>"011101100",
  10737=>"101101010",
  10738=>"011110110",
  10739=>"000100001",
  10740=>"110110110",
  10741=>"010100011",
  10742=>"011110010",
  10743=>"001001110",
  10744=>"100100001",
  10745=>"000000100",
  10746=>"101000000",
  10747=>"100010011",
  10748=>"111000101",
  10749=>"101100010",
  10750=>"001101100",
  10751=>"000000010",
  10752=>"011000000",
  10753=>"011100001",
  10754=>"000100011",
  10755=>"111001101",
  10756=>"100001100",
  10757=>"010011011",
  10758=>"101110010",
  10759=>"110111110",
  10760=>"110111011",
  10761=>"100110000",
  10762=>"001000111",
  10763=>"010000111",
  10764=>"011111000",
  10765=>"101100010",
  10766=>"000011100",
  10767=>"111111010",
  10768=>"001110011",
  10769=>"101010011",
  10770=>"001110000",
  10771=>"010110010",
  10772=>"001000101",
  10773=>"110100110",
  10774=>"010111001",
  10775=>"110101010",
  10776=>"101010110",
  10777=>"000001110",
  10778=>"011000001",
  10779=>"110100010",
  10780=>"101011010",
  10781=>"101010010",
  10782=>"111100101",
  10783=>"000101000",
  10784=>"110111010",
  10785=>"110101001",
  10786=>"010101101",
  10787=>"010101000",
  10788=>"110011010",
  10789=>"110100101",
  10790=>"001010110",
  10791=>"111000010",
  10792=>"011111011",
  10793=>"011000100",
  10794=>"001010010",
  10795=>"101001100",
  10796=>"100011011",
  10797=>"110101110",
  10798=>"000011010",
  10799=>"010000011",
  10800=>"001111001",
  10801=>"100000010",
  10802=>"111111000",
  10803=>"011011011",
  10804=>"110000100",
  10805=>"110011010",
  10806=>"111100100",
  10807=>"011010011",
  10808=>"010100011",
  10809=>"110001101",
  10810=>"010001100",
  10811=>"010011010",
  10812=>"011110011",
  10813=>"101110110",
  10814=>"100001011",
  10815=>"010000101",
  10816=>"110111110",
  10817=>"101100001",
  10818=>"000000110",
  10819=>"111011001",
  10820=>"010001101",
  10821=>"111000111",
  10822=>"000010111",
  10823=>"100000111",
  10824=>"001001001",
  10825=>"101111000",
  10826=>"010001110",
  10827=>"101010000",
  10828=>"001111011",
  10829=>"111101001",
  10830=>"100001111",
  10831=>"101000100",
  10832=>"001100101",
  10833=>"100101001",
  10834=>"001111110",
  10835=>"010001101",
  10836=>"011110100",
  10837=>"001111011",
  10838=>"011011011",
  10839=>"100110001",
  10840=>"100011111",
  10841=>"000001100",
  10842=>"000101010",
  10843=>"001011010",
  10844=>"001100100",
  10845=>"101100010",
  10846=>"110100001",
  10847=>"101100110",
  10848=>"010000001",
  10849=>"000110110",
  10850=>"100101011",
  10851=>"011010101",
  10852=>"001101011",
  10853=>"011101100",
  10854=>"000000110",
  10855=>"010011100",
  10856=>"100111100",
  10857=>"110100000",
  10858=>"001110010",
  10859=>"110011000",
  10860=>"000100100",
  10861=>"001010011",
  10862=>"111111011",
  10863=>"101001010",
  10864=>"110011010",
  10865=>"011101100",
  10866=>"100011111",
  10867=>"101100100",
  10868=>"001111110",
  10869=>"000111101",
  10870=>"011011110",
  10871=>"001011000",
  10872=>"111000110",
  10873=>"110110111",
  10874=>"110100001",
  10875=>"100000000",
  10876=>"000011011",
  10877=>"001011001",
  10878=>"001000010",
  10879=>"111111000",
  10880=>"001111000",
  10881=>"000111110",
  10882=>"101001100",
  10883=>"100110000",
  10884=>"000100001",
  10885=>"101101100",
  10886=>"000011111",
  10887=>"100111010",
  10888=>"000000000",
  10889=>"010111101",
  10890=>"101000100",
  10891=>"001011111",
  10892=>"000100010",
  10893=>"110101011",
  10894=>"111011000",
  10895=>"110000111",
  10896=>"100111000",
  10897=>"100000000",
  10898=>"010000100",
  10899=>"000111000",
  10900=>"011000111",
  10901=>"011010100",
  10902=>"001011101",
  10903=>"010101110",
  10904=>"001000110",
  10905=>"000101110",
  10906=>"000010011",
  10907=>"010101001",
  10908=>"101110000",
  10909=>"110101011",
  10910=>"110000111",
  10911=>"101010110",
  10912=>"010110001",
  10913=>"010111000",
  10914=>"001101111",
  10915=>"110110001",
  10916=>"000000001",
  10917=>"000000101",
  10918=>"110000001",
  10919=>"000100000",
  10920=>"001100011",
  10921=>"001000101",
  10922=>"111110110",
  10923=>"111000001",
  10924=>"000001110",
  10925=>"001100100",
  10926=>"000110010",
  10927=>"000000000",
  10928=>"101100001",
  10929=>"110110101",
  10930=>"011001100",
  10931=>"111111100",
  10932=>"010001101",
  10933=>"101101011",
  10934=>"101101000",
  10935=>"001000111",
  10936=>"101001010",
  10937=>"110001001",
  10938=>"001111000",
  10939=>"110000100",
  10940=>"110100010",
  10941=>"001100111",
  10942=>"111001011",
  10943=>"110000101",
  10944=>"111011111",
  10945=>"101100001",
  10946=>"010110011",
  10947=>"101110001",
  10948=>"110111001",
  10949=>"110010111",
  10950=>"001111001",
  10951=>"001000000",
  10952=>"111111010",
  10953=>"010110100",
  10954=>"000011111",
  10955=>"011111010",
  10956=>"110111101",
  10957=>"000010100",
  10958=>"101101001",
  10959=>"100010010",
  10960=>"110111101",
  10961=>"000010001",
  10962=>"001100000",
  10963=>"111111001",
  10964=>"111101111",
  10965=>"011100101",
  10966=>"100011100",
  10967=>"111011001",
  10968=>"110110111",
  10969=>"001000110",
  10970=>"001110101",
  10971=>"001011111",
  10972=>"001000110",
  10973=>"001010000",
  10974=>"100000010",
  10975=>"001110111",
  10976=>"110001010",
  10977=>"011010000",
  10978=>"100111110",
  10979=>"100111101",
  10980=>"000100010",
  10981=>"100001000",
  10982=>"010011001",
  10983=>"001011010",
  10984=>"101010010",
  10985=>"000110001",
  10986=>"100001001",
  10987=>"110111010",
  10988=>"000111011",
  10989=>"010011100",
  10990=>"100000110",
  10991=>"101100101",
  10992=>"101010100",
  10993=>"111100010",
  10994=>"010001001",
  10995=>"001000111",
  10996=>"111001110",
  10997=>"010001101",
  10998=>"010001100",
  10999=>"111011011",
  11000=>"111011001",
  11001=>"110100000",
  11002=>"100111101",
  11003=>"000000110",
  11004=>"010010011",
  11005=>"011100111",
  11006=>"110011110",
  11007=>"001001100",
  11008=>"001100111",
  11009=>"101100110",
  11010=>"110011001",
  11011=>"111010111",
  11012=>"000101111",
  11013=>"100100110",
  11014=>"110000010",
  11015=>"011110111",
  11016=>"101000011",
  11017=>"010100111",
  11018=>"010001000",
  11019=>"110000011",
  11020=>"011001111",
  11021=>"110001110",
  11022=>"010111000",
  11023=>"100000011",
  11024=>"101100101",
  11025=>"100100101",
  11026=>"100000111",
  11027=>"111010000",
  11028=>"101001100",
  11029=>"010011000",
  11030=>"010000100",
  11031=>"001011000",
  11032=>"001101100",
  11033=>"000011000",
  11034=>"101101111",
  11035=>"010110100",
  11036=>"011001001",
  11037=>"001010110",
  11038=>"101010001",
  11039=>"101111010",
  11040=>"000000110",
  11041=>"100000100",
  11042=>"000111110",
  11043=>"100000000",
  11044=>"101100110",
  11045=>"000001001",
  11046=>"011111001",
  11047=>"000111110",
  11048=>"010111110",
  11049=>"111111001",
  11050=>"111100010",
  11051=>"101110000",
  11052=>"000001110",
  11053=>"110010010",
  11054=>"110111000",
  11055=>"011010000",
  11056=>"000100000",
  11057=>"011000111",
  11058=>"010110011",
  11059=>"100000100",
  11060=>"000001000",
  11061=>"000111000",
  11062=>"011011101",
  11063=>"011110001",
  11064=>"110010010",
  11065=>"110000000",
  11066=>"010000010",
  11067=>"010011001",
  11068=>"100000011",
  11069=>"110100000",
  11070=>"110110110",
  11071=>"000001100",
  11072=>"110001100",
  11073=>"110100000",
  11074=>"011001111",
  11075=>"110001010",
  11076=>"000000110",
  11077=>"011001000",
  11078=>"101110111",
  11079=>"111111011",
  11080=>"011011011",
  11081=>"000100110",
  11082=>"011001111",
  11083=>"010000001",
  11084=>"101101011",
  11085=>"101010111",
  11086=>"001111001",
  11087=>"001000010",
  11088=>"100101101",
  11089=>"110100100",
  11090=>"010100111",
  11091=>"010111001",
  11092=>"101001100",
  11093=>"001001111",
  11094=>"110010111",
  11095=>"010101111",
  11096=>"010010000",
  11097=>"110001001",
  11098=>"000001000",
  11099=>"010111101",
  11100=>"111000011",
  11101=>"010000100",
  11102=>"111110110",
  11103=>"101100001",
  11104=>"110001110",
  11105=>"100010101",
  11106=>"100100011",
  11107=>"111111111",
  11108=>"010001010",
  11109=>"101000110",
  11110=>"000111110",
  11111=>"011000100",
  11112=>"011000010",
  11113=>"001010001",
  11114=>"001101001",
  11115=>"111101101",
  11116=>"101110000",
  11117=>"010001011",
  11118=>"100000100",
  11119=>"011001001",
  11120=>"110100010",
  11121=>"100110111",
  11122=>"011000011",
  11123=>"110001110",
  11124=>"010110101",
  11125=>"001100010",
  11126=>"110111100",
  11127=>"100100011",
  11128=>"011010001",
  11129=>"110010101",
  11130=>"100110011",
  11131=>"001100111",
  11132=>"100000011",
  11133=>"000000000",
  11134=>"100000111",
  11135=>"111110110",
  11136=>"101010000",
  11137=>"001101101",
  11138=>"101110010",
  11139=>"110100100",
  11140=>"110001111",
  11141=>"000001110",
  11142=>"110111111",
  11143=>"010110100",
  11144=>"110001101",
  11145=>"001100111",
  11146=>"010100010",
  11147=>"111000111",
  11148=>"100110111",
  11149=>"100110000",
  11150=>"000000001",
  11151=>"010010000",
  11152=>"001101000",
  11153=>"001010000",
  11154=>"101111110",
  11155=>"011001001",
  11156=>"101000010",
  11157=>"000101111",
  11158=>"010100101",
  11159=>"111000011",
  11160=>"011001100",
  11161=>"100011101",
  11162=>"110111110",
  11163=>"110100011",
  11164=>"001011110",
  11165=>"101101110",
  11166=>"101011011",
  11167=>"110000010",
  11168=>"101010100",
  11169=>"001100101",
  11170=>"111011111",
  11171=>"110011111",
  11172=>"010011001",
  11173=>"000011110",
  11174=>"000101001",
  11175=>"100000001",
  11176=>"000110111",
  11177=>"100001000",
  11178=>"000100111",
  11179=>"001000001",
  11180=>"111011101",
  11181=>"111111100",
  11182=>"001111010",
  11183=>"100110010",
  11184=>"100001011",
  11185=>"110001100",
  11186=>"100110001",
  11187=>"001101111",
  11188=>"111110111",
  11189=>"111010011",
  11190=>"010001011",
  11191=>"011000100",
  11192=>"000101010",
  11193=>"011001101",
  11194=>"011000101",
  11195=>"001000001",
  11196=>"011111001",
  11197=>"010101001",
  11198=>"110010001",
  11199=>"101111011",
  11200=>"111011011",
  11201=>"011110001",
  11202=>"011000010",
  11203=>"110100101",
  11204=>"011111011",
  11205=>"010001011",
  11206=>"111100001",
  11207=>"000101011",
  11208=>"011101110",
  11209=>"011011100",
  11210=>"001101100",
  11211=>"111111000",
  11212=>"110000101",
  11213=>"000100001",
  11214=>"000011001",
  11215=>"110110010",
  11216=>"101101111",
  11217=>"001110011",
  11218=>"110111111",
  11219=>"100001110",
  11220=>"111010011",
  11221=>"011011010",
  11222=>"000100001",
  11223=>"011010111",
  11224=>"101101011",
  11225=>"110111111",
  11226=>"010011111",
  11227=>"110110001",
  11228=>"100011011",
  11229=>"110111101",
  11230=>"110010111",
  11231=>"011110001",
  11232=>"100001011",
  11233=>"001101001",
  11234=>"000100101",
  11235=>"101000100",
  11236=>"010001000",
  11237=>"101111011",
  11238=>"000111101",
  11239=>"100111100",
  11240=>"111111010",
  11241=>"111101101",
  11242=>"011111100",
  11243=>"111110000",
  11244=>"101101011",
  11245=>"101101100",
  11246=>"111011010",
  11247=>"011000001",
  11248=>"110101100",
  11249=>"100110101",
  11250=>"000000111",
  11251=>"010111010",
  11252=>"111101001",
  11253=>"011110101",
  11254=>"000100100",
  11255=>"101000101",
  11256=>"001110100",
  11257=>"110111101",
  11258=>"101100100",
  11259=>"010111110",
  11260=>"101000001",
  11261=>"001010110",
  11262=>"110010010",
  11263=>"001110111",
  11264=>"101111111",
  11265=>"101000011",
  11266=>"000100010",
  11267=>"110101100",
  11268=>"001101101",
  11269=>"010000111",
  11270=>"001111001",
  11271=>"110100110",
  11272=>"101111001",
  11273=>"011101110",
  11274=>"110100110",
  11275=>"000100000",
  11276=>"000100001",
  11277=>"101110011",
  11278=>"111110000",
  11279=>"110101010",
  11280=>"101001001",
  11281=>"010000111",
  11282=>"010100000",
  11283=>"100011100",
  11284=>"100010110",
  11285=>"110100001",
  11286=>"000100000",
  11287=>"101010001",
  11288=>"101100110",
  11289=>"000111101",
  11290=>"110110110",
  11291=>"100110010",
  11292=>"110010101",
  11293=>"000011111",
  11294=>"100100111",
  11295=>"010000111",
  11296=>"000010010",
  11297=>"001100110",
  11298=>"010101011",
  11299=>"010000001",
  11300=>"111000000",
  11301=>"100000000",
  11302=>"010101101",
  11303=>"010000010",
  11304=>"010111011",
  11305=>"101001001",
  11306=>"011001001",
  11307=>"101111110",
  11308=>"010110111",
  11309=>"000110111",
  11310=>"001001001",
  11311=>"110111110",
  11312=>"010110010",
  11313=>"001010100",
  11314=>"101010001",
  11315=>"001100111",
  11316=>"010000001",
  11317=>"101011001",
  11318=>"001010100",
  11319=>"100100111",
  11320=>"011001101",
  11321=>"111010001",
  11322=>"110010110",
  11323=>"110111010",
  11324=>"010011100",
  11325=>"010000000",
  11326=>"101000010",
  11327=>"010001010",
  11328=>"101110010",
  11329=>"000110010",
  11330=>"001001010",
  11331=>"011110011",
  11332=>"011110101",
  11333=>"011010011",
  11334=>"000000111",
  11335=>"010000101",
  11336=>"100111111",
  11337=>"101001000",
  11338=>"101101000",
  11339=>"100001100",
  11340=>"111001011",
  11341=>"100010111",
  11342=>"111100100",
  11343=>"110100111",
  11344=>"010010110",
  11345=>"010001010",
  11346=>"110100011",
  11347=>"010110101",
  11348=>"001100110",
  11349=>"100011010",
  11350=>"000101000",
  11351=>"010001110",
  11352=>"011101110",
  11353=>"111100101",
  11354=>"111111001",
  11355=>"011010000",
  11356=>"101011000",
  11357=>"001110010",
  11358=>"000110111",
  11359=>"000000001",
  11360=>"100110000",
  11361=>"111011010",
  11362=>"000010111",
  11363=>"011011101",
  11364=>"100110111",
  11365=>"001110001",
  11366=>"100000000",
  11367=>"111101101",
  11368=>"010101101",
  11369=>"111101010",
  11370=>"111110101",
  11371=>"100001100",
  11372=>"111010101",
  11373=>"110100001",
  11374=>"001000010",
  11375=>"000100000",
  11376=>"000001011",
  11377=>"000001111",
  11378=>"000011000",
  11379=>"111111110",
  11380=>"101110011",
  11381=>"100101010",
  11382=>"011011101",
  11383=>"100111100",
  11384=>"111000001",
  11385=>"000100001",
  11386=>"100010111",
  11387=>"010010110",
  11388=>"010111001",
  11389=>"100101100",
  11390=>"110101000",
  11391=>"000101001",
  11392=>"101111101",
  11393=>"101011110",
  11394=>"011101110",
  11395=>"100011000",
  11396=>"101011001",
  11397=>"000000111",
  11398=>"010111100",
  11399=>"011101011",
  11400=>"010111011",
  11401=>"011101011",
  11402=>"111000111",
  11403=>"100001101",
  11404=>"001010100",
  11405=>"111001001",
  11406=>"001111110",
  11407=>"111011110",
  11408=>"110100110",
  11409=>"011001110",
  11410=>"010100000",
  11411=>"101010011",
  11412=>"001111001",
  11413=>"011100111",
  11414=>"000010100",
  11415=>"011000001",
  11416=>"111100110",
  11417=>"000000000",
  11418=>"000011000",
  11419=>"101001101",
  11420=>"011100100",
  11421=>"100011001",
  11422=>"110111001",
  11423=>"100101010",
  11424=>"000100000",
  11425=>"110111100",
  11426=>"001001011",
  11427=>"011001001",
  11428=>"100100110",
  11429=>"000001101",
  11430=>"010110011",
  11431=>"101110100",
  11432=>"011010110",
  11433=>"001000000",
  11434=>"101001101",
  11435=>"111101110",
  11436=>"101011010",
  11437=>"010111101",
  11438=>"110011100",
  11439=>"101101010",
  11440=>"011111111",
  11441=>"001001100",
  11442=>"000011010",
  11443=>"100000010",
  11444=>"000111001",
  11445=>"010000110",
  11446=>"110110011",
  11447=>"100001111",
  11448=>"000010101",
  11449=>"000111111",
  11450=>"111011011",
  11451=>"001010101",
  11452=>"110000010",
  11453=>"001011000",
  11454=>"010001100",
  11455=>"101111011",
  11456=>"100111011",
  11457=>"101010111",
  11458=>"010110001",
  11459=>"001110110",
  11460=>"111110101",
  11461=>"111010100",
  11462=>"011000000",
  11463=>"101101011",
  11464=>"000000111",
  11465=>"010000110",
  11466=>"001111100",
  11467=>"011100010",
  11468=>"001011100",
  11469=>"110001010",
  11470=>"000010010",
  11471=>"011100010",
  11472=>"000100100",
  11473=>"010001100",
  11474=>"101011100",
  11475=>"011000010",
  11476=>"111011011",
  11477=>"011110111",
  11478=>"100111011",
  11479=>"001001011",
  11480=>"100100101",
  11481=>"110101100",
  11482=>"100110001",
  11483=>"000100011",
  11484=>"101101000",
  11485=>"110011100",
  11486=>"010101100",
  11487=>"110001000",
  11488=>"000100111",
  11489=>"110100010",
  11490=>"111100111",
  11491=>"101111100",
  11492=>"101111110",
  11493=>"001110001",
  11494=>"000101000",
  11495=>"000110010",
  11496=>"000010000",
  11497=>"000011111",
  11498=>"101111001",
  11499=>"111010000",
  11500=>"000111011",
  11501=>"100110010",
  11502=>"001010100",
  11503=>"000000100",
  11504=>"111010100",
  11505=>"111001101",
  11506=>"101000010",
  11507=>"001011000",
  11508=>"010001001",
  11509=>"110010011",
  11510=>"010110010",
  11511=>"110101010",
  11512=>"010000010",
  11513=>"110101110",
  11514=>"010111010",
  11515=>"110011100",
  11516=>"001000110",
  11517=>"110111010",
  11518=>"010010110",
  11519=>"000111001",
  11520=>"100011111",
  11521=>"010111011",
  11522=>"000001101",
  11523=>"011101110",
  11524=>"110011110",
  11525=>"110011100",
  11526=>"101000001",
  11527=>"001110100",
  11528=>"011101001",
  11529=>"010010110",
  11530=>"001000110",
  11531=>"100001101",
  11532=>"110000100",
  11533=>"111011111",
  11534=>"000101100",
  11535=>"101111101",
  11536=>"110101011",
  11537=>"110011101",
  11538=>"001011001",
  11539=>"101010101",
  11540=>"100011101",
  11541=>"000000110",
  11542=>"100110000",
  11543=>"100111001",
  11544=>"010110100",
  11545=>"010011000",
  11546=>"101100011",
  11547=>"000101111",
  11548=>"111011100",
  11549=>"011100100",
  11550=>"110110110",
  11551=>"000000110",
  11552=>"000110011",
  11553=>"010101111",
  11554=>"000111111",
  11555=>"000011001",
  11556=>"101110111",
  11557=>"010010000",
  11558=>"001110011",
  11559=>"001000100",
  11560=>"001010110",
  11561=>"001001100",
  11562=>"111000000",
  11563=>"001101011",
  11564=>"100101000",
  11565=>"101111001",
  11566=>"001011010",
  11567=>"101010010",
  11568=>"001001001",
  11569=>"101110010",
  11570=>"101110010",
  11571=>"011110101",
  11572=>"000001010",
  11573=>"000100110",
  11574=>"111100101",
  11575=>"110000111",
  11576=>"001001000",
  11577=>"111111000",
  11578=>"100100110",
  11579=>"000001100",
  11580=>"110101110",
  11581=>"101000010",
  11582=>"011000000",
  11583=>"111100000",
  11584=>"110011011",
  11585=>"011110110",
  11586=>"000110111",
  11587=>"011110111",
  11588=>"000110000",
  11589=>"101111011",
  11590=>"111111000",
  11591=>"000000111",
  11592=>"010001000",
  11593=>"010011110",
  11594=>"111100111",
  11595=>"010011000",
  11596=>"101011010",
  11597=>"110010111",
  11598=>"000111111",
  11599=>"111010001",
  11600=>"001001100",
  11601=>"100001100",
  11602=>"111011101",
  11603=>"000001111",
  11604=>"110000111",
  11605=>"101101110",
  11606=>"100001000",
  11607=>"100101001",
  11608=>"111011110",
  11609=>"101101000",
  11610=>"011110100",
  11611=>"000000101",
  11612=>"000110001",
  11613=>"001010001",
  11614=>"010001111",
  11615=>"111110101",
  11616=>"011110000",
  11617=>"100010000",
  11618=>"110011000",
  11619=>"000001011",
  11620=>"001110110",
  11621=>"000101011",
  11622=>"010000001",
  11623=>"001010001",
  11624=>"001110110",
  11625=>"111101100",
  11626=>"011000000",
  11627=>"001010101",
  11628=>"010000110",
  11629=>"011010110",
  11630=>"000001100",
  11631=>"100100001",
  11632=>"101110100",
  11633=>"101000100",
  11634=>"000110111",
  11635=>"110000011",
  11636=>"000000010",
  11637=>"001010100",
  11638=>"000101111",
  11639=>"001010011",
  11640=>"100101011",
  11641=>"101001101",
  11642=>"100101001",
  11643=>"100011101",
  11644=>"001101010",
  11645=>"000011111",
  11646=>"001110010",
  11647=>"100101000",
  11648=>"001111110",
  11649=>"000000000",
  11650=>"011010101",
  11651=>"110111000",
  11652=>"000110111",
  11653=>"110001010",
  11654=>"001000100",
  11655=>"011010001",
  11656=>"110010010",
  11657=>"011000011",
  11658=>"101111110",
  11659=>"101001111",
  11660=>"000000011",
  11661=>"111011010",
  11662=>"101110101",
  11663=>"001101000",
  11664=>"111101011",
  11665=>"010000000",
  11666=>"110110110",
  11667=>"011111001",
  11668=>"100111000",
  11669=>"000100000",
  11670=>"111001010",
  11671=>"101100111",
  11672=>"101000100",
  11673=>"100100101",
  11674=>"010111001",
  11675=>"001001100",
  11676=>"011111110",
  11677=>"101010101",
  11678=>"111111110",
  11679=>"011110000",
  11680=>"001000111",
  11681=>"111000000",
  11682=>"010001111",
  11683=>"000011001",
  11684=>"001100111",
  11685=>"011100111",
  11686=>"110111001",
  11687=>"111110110",
  11688=>"110000110",
  11689=>"001000000",
  11690=>"000101100",
  11691=>"011010101",
  11692=>"000101100",
  11693=>"000101100",
  11694=>"111010111",
  11695=>"010100000",
  11696=>"001001100",
  11697=>"111100010",
  11698=>"101111010",
  11699=>"110111100",
  11700=>"111110100",
  11701=>"101010100",
  11702=>"001110010",
  11703=>"110000100",
  11704=>"100001001",
  11705=>"000010011",
  11706=>"111110101",
  11707=>"111010100",
  11708=>"111011011",
  11709=>"110100000",
  11710=>"100010101",
  11711=>"101010111",
  11712=>"001111001",
  11713=>"110110110",
  11714=>"100100110",
  11715=>"100000000",
  11716=>"101111101",
  11717=>"100101010",
  11718=>"100100110",
  11719=>"001110100",
  11720=>"100011111",
  11721=>"010001000",
  11722=>"000110011",
  11723=>"110100000",
  11724=>"111011100",
  11725=>"111110001",
  11726=>"011010000",
  11727=>"111101110",
  11728=>"011011010",
  11729=>"010010100",
  11730=>"000000001",
  11731=>"010010001",
  11732=>"100101011",
  11733=>"101000111",
  11734=>"101000110",
  11735=>"001110011",
  11736=>"000101101",
  11737=>"011010110",
  11738=>"010110011",
  11739=>"100001001",
  11740=>"100101000",
  11741=>"000110100",
  11742=>"111101001",
  11743=>"100000111",
  11744=>"100010111",
  11745=>"100110000",
  11746=>"011010010",
  11747=>"000000001",
  11748=>"010010000",
  11749=>"011110011",
  11750=>"101010010",
  11751=>"111000101",
  11752=>"110101100",
  11753=>"110110001",
  11754=>"111000100",
  11755=>"011011011",
  11756=>"101101010",
  11757=>"000011010",
  11758=>"110111111",
  11759=>"111010110",
  11760=>"011010001",
  11761=>"001010111",
  11762=>"100010101",
  11763=>"110001000",
  11764=>"011010101",
  11765=>"101110011",
  11766=>"011011011",
  11767=>"110000001",
  11768=>"000010100",
  11769=>"111110111",
  11770=>"001011101",
  11771=>"101101011",
  11772=>"000011011",
  11773=>"101011001",
  11774=>"001010110",
  11775=>"100000100",
  11776=>"111100010",
  11777=>"011101101",
  11778=>"000011111",
  11779=>"110101000",
  11780=>"111110011",
  11781=>"111011000",
  11782=>"010100100",
  11783=>"011000000",
  11784=>"111001010",
  11785=>"001100110",
  11786=>"100100110",
  11787=>"001011010",
  11788=>"111000100",
  11789=>"011100111",
  11790=>"000001110",
  11791=>"111011101",
  11792=>"011001010",
  11793=>"000110001",
  11794=>"100010111",
  11795=>"011011011",
  11796=>"111100000",
  11797=>"101101100",
  11798=>"110001001",
  11799=>"011001101",
  11800=>"000101111",
  11801=>"110110001",
  11802=>"101000001",
  11803=>"101100010",
  11804=>"100111110",
  11805=>"110011000",
  11806=>"111010000",
  11807=>"001100100",
  11808=>"000001000",
  11809=>"011100010",
  11810=>"001100000",
  11811=>"101011011",
  11812=>"000110001",
  11813=>"110001100",
  11814=>"110010010",
  11815=>"000101010",
  11816=>"001111001",
  11817=>"011011100",
  11818=>"000100000",
  11819=>"111011011",
  11820=>"101111110",
  11821=>"010101101",
  11822=>"100001111",
  11823=>"110110001",
  11824=>"000110100",
  11825=>"110011111",
  11826=>"010110110",
  11827=>"001101000",
  11828=>"001010100",
  11829=>"011001100",
  11830=>"011000111",
  11831=>"101101110",
  11832=>"110110111",
  11833=>"011110111",
  11834=>"111010101",
  11835=>"110111101",
  11836=>"010101101",
  11837=>"010110001",
  11838=>"100000101",
  11839=>"100000100",
  11840=>"110000110",
  11841=>"101011100",
  11842=>"100010101",
  11843=>"110110110",
  11844=>"100011100",
  11845=>"111111111",
  11846=>"001000010",
  11847=>"011101110",
  11848=>"011101110",
  11849=>"010111101",
  11850=>"001000110",
  11851=>"010011101",
  11852=>"101110110",
  11853=>"100000111",
  11854=>"101010000",
  11855=>"001011111",
  11856=>"110001000",
  11857=>"101000000",
  11858=>"010100001",
  11859=>"010010110",
  11860=>"011001011",
  11861=>"010000000",
  11862=>"111101010",
  11863=>"001111000",
  11864=>"100001100",
  11865=>"100000111",
  11866=>"000011000",
  11867=>"000101110",
  11868=>"110101110",
  11869=>"101100111",
  11870=>"011100010",
  11871=>"110101000",
  11872=>"000001111",
  11873=>"101000010",
  11874=>"011111100",
  11875=>"100110011",
  11876=>"100100100",
  11877=>"100011000",
  11878=>"011100111",
  11879=>"001010111",
  11880=>"101001010",
  11881=>"001000010",
  11882=>"010000110",
  11883=>"000000000",
  11884=>"111110000",
  11885=>"100000010",
  11886=>"011100101",
  11887=>"100010001",
  11888=>"011100001",
  11889=>"111111111",
  11890=>"101011000",
  11891=>"100010000",
  11892=>"001000011",
  11893=>"100010110",
  11894=>"111100011",
  11895=>"111100101",
  11896=>"000000110",
  11897=>"000101111",
  11898=>"000010000",
  11899=>"001110000",
  11900=>"101010010",
  11901=>"100110010",
  11902=>"011101111",
  11903=>"001000101",
  11904=>"000000011",
  11905=>"101101101",
  11906=>"100001000",
  11907=>"011110000",
  11908=>"110110011",
  11909=>"110010001",
  11910=>"100110111",
  11911=>"110100011",
  11912=>"000111001",
  11913=>"001000101",
  11914=>"110110110",
  11915=>"010110010",
  11916=>"110001010",
  11917=>"001000010",
  11918=>"110010011",
  11919=>"111110001",
  11920=>"111001100",
  11921=>"011011110",
  11922=>"110001011",
  11923=>"010011111",
  11924=>"110110111",
  11925=>"100010000",
  11926=>"000010000",
  11927=>"110111011",
  11928=>"000100000",
  11929=>"011011101",
  11930=>"001001010",
  11931=>"111010011",
  11932=>"111110100",
  11933=>"101001001",
  11934=>"101000100",
  11935=>"011111000",
  11936=>"101011111",
  11937=>"001100001",
  11938=>"100100001",
  11939=>"011100011",
  11940=>"001110110",
  11941=>"001111100",
  11942=>"010111101",
  11943=>"110111011",
  11944=>"110000101",
  11945=>"000001100",
  11946=>"011010101",
  11947=>"100011010",
  11948=>"101011001",
  11949=>"000110111",
  11950=>"110101010",
  11951=>"001100010",
  11952=>"100111100",
  11953=>"110101100",
  11954=>"000000010",
  11955=>"110111000",
  11956=>"011110101",
  11957=>"100110001",
  11958=>"111000001",
  11959=>"111011111",
  11960=>"001101100",
  11961=>"011100000",
  11962=>"010001001",
  11963=>"000101010",
  11964=>"010100000",
  11965=>"100110100",
  11966=>"110110110",
  11967=>"000110100",
  11968=>"110011110",
  11969=>"000101101",
  11970=>"101111111",
  11971=>"111010011",
  11972=>"100011101",
  11973=>"010010110",
  11974=>"111010110",
  11975=>"100111000",
  11976=>"111111000",
  11977=>"111110011",
  11978=>"011011011",
  11979=>"011010011",
  11980=>"100011011",
  11981=>"001010110",
  11982=>"001101010",
  11983=>"010010010",
  11984=>"010100011",
  11985=>"001011001",
  11986=>"110011011",
  11987=>"110101110",
  11988=>"101100011",
  11989=>"000111010",
  11990=>"010100110",
  11991=>"110000110",
  11992=>"000010000",
  11993=>"011010101",
  11994=>"101111111",
  11995=>"111111110",
  11996=>"101101010",
  11997=>"001101001",
  11998=>"101010000",
  11999=>"000101111",
  12000=>"111000010",
  12001=>"000110010",
  12002=>"110001110",
  12003=>"001000101",
  12004=>"101001101",
  12005=>"010000111",
  12006=>"100111111",
  12007=>"110010101",
  12008=>"111010101",
  12009=>"110001000",
  12010=>"011010110",
  12011=>"110001001",
  12012=>"111011100",
  12013=>"110011111",
  12014=>"100000001",
  12015=>"111101111",
  12016=>"011100101",
  12017=>"101011100",
  12018=>"100101101",
  12019=>"011101010",
  12020=>"011011011",
  12021=>"100101010",
  12022=>"100110000",
  12023=>"010001100",
  12024=>"010000100",
  12025=>"100000010",
  12026=>"111101001",
  12027=>"111011001",
  12028=>"101011011",
  12029=>"101111101",
  12030=>"001101100",
  12031=>"011101110",
  12032=>"000000001",
  12033=>"111111000",
  12034=>"111010111",
  12035=>"100000100",
  12036=>"111100001",
  12037=>"111001111",
  12038=>"010001110",
  12039=>"000100010",
  12040=>"101001000",
  12041=>"110111110",
  12042=>"101010010",
  12043=>"111111101",
  12044=>"001001111",
  12045=>"011111111",
  12046=>"100110010",
  12047=>"101011000",
  12048=>"010000001",
  12049=>"110100001",
  12050=>"111100001",
  12051=>"010010101",
  12052=>"101101000",
  12053=>"000001011",
  12054=>"000000011",
  12055=>"100000111",
  12056=>"100100110",
  12057=>"000000101",
  12058=>"101000000",
  12059=>"001010001",
  12060=>"100110001",
  12061=>"110001011",
  12062=>"010110011",
  12063=>"100010010",
  12064=>"110111110",
  12065=>"000101110",
  12066=>"000010011",
  12067=>"101110001",
  12068=>"111011010",
  12069=>"011100001",
  12070=>"011001101",
  12071=>"000000100",
  12072=>"111101101",
  12073=>"101111011",
  12074=>"010111000",
  12075=>"001010010",
  12076=>"000010001",
  12077=>"111110110",
  12078=>"110100000",
  12079=>"100000010",
  12080=>"111100111",
  12081=>"111011001",
  12082=>"011111110",
  12083=>"111010100",
  12084=>"010010111",
  12085=>"001001010",
  12086=>"011001111",
  12087=>"000111111",
  12088=>"011111110",
  12089=>"000001010",
  12090=>"001010100",
  12091=>"101001110",
  12092=>"100111010",
  12093=>"100001110",
  12094=>"001011010",
  12095=>"001100001",
  12096=>"001001001",
  12097=>"110001110",
  12098=>"100111111",
  12099=>"100100011",
  12100=>"110110010",
  12101=>"100001011",
  12102=>"011011001",
  12103=>"000101011",
  12104=>"000010110",
  12105=>"100011110",
  12106=>"011101110",
  12107=>"110000101",
  12108=>"101110011",
  12109=>"100000101",
  12110=>"110000010",
  12111=>"001011011",
  12112=>"110001111",
  12113=>"111001000",
  12114=>"111100111",
  12115=>"011000111",
  12116=>"011000111",
  12117=>"101110110",
  12118=>"011011101",
  12119=>"111111010",
  12120=>"011110011",
  12121=>"101100100",
  12122=>"000111001",
  12123=>"111110001",
  12124=>"100111010",
  12125=>"001001101",
  12126=>"011100010",
  12127=>"001011111",
  12128=>"110110001",
  12129=>"110001000",
  12130=>"001000010",
  12131=>"011111110",
  12132=>"001010001",
  12133=>"001010000",
  12134=>"111111110",
  12135=>"011111111",
  12136=>"101000000",
  12137=>"011001011",
  12138=>"100101001",
  12139=>"011011100",
  12140=>"000100111",
  12141=>"110100000",
  12142=>"111110001",
  12143=>"011010101",
  12144=>"000011110",
  12145=>"010011100",
  12146=>"111111010",
  12147=>"100011010",
  12148=>"001101010",
  12149=>"101010001",
  12150=>"101111101",
  12151=>"000010010",
  12152=>"011111000",
  12153=>"001001101",
  12154=>"011110110",
  12155=>"111000100",
  12156=>"110110110",
  12157=>"111100000",
  12158=>"110110010",
  12159=>"011011010",
  12160=>"111011001",
  12161=>"111101100",
  12162=>"111010110",
  12163=>"000011100",
  12164=>"001010101",
  12165=>"001001001",
  12166=>"000101110",
  12167=>"110001000",
  12168=>"011100111",
  12169=>"111000011",
  12170=>"111010000",
  12171=>"100000000",
  12172=>"101010000",
  12173=>"000110111",
  12174=>"000100000",
  12175=>"111100101",
  12176=>"101001001",
  12177=>"100111011",
  12178=>"100111011",
  12179=>"000000101",
  12180=>"101110001",
  12181=>"101111100",
  12182=>"010110010",
  12183=>"110010011",
  12184=>"111011101",
  12185=>"000110101",
  12186=>"011101111",
  12187=>"100100001",
  12188=>"100110101",
  12189=>"100111100",
  12190=>"000100000",
  12191=>"001111110",
  12192=>"011000011",
  12193=>"100000101",
  12194=>"111110110",
  12195=>"000100110",
  12196=>"110010001",
  12197=>"100010110",
  12198=>"001000001",
  12199=>"111111110",
  12200=>"110001000",
  12201=>"100000110",
  12202=>"001000101",
  12203=>"010001110",
  12204=>"001100001",
  12205=>"101101111",
  12206=>"100000111",
  12207=>"101001110",
  12208=>"001100000",
  12209=>"010011110",
  12210=>"101100000",
  12211=>"000001110",
  12212=>"001111110",
  12213=>"111100110",
  12214=>"111011100",
  12215=>"001000101",
  12216=>"111000001",
  12217=>"011111111",
  12218=>"100100101",
  12219=>"111111100",
  12220=>"001010111",
  12221=>"101110100",
  12222=>"111111001",
  12223=>"111000100",
  12224=>"001011111",
  12225=>"101010111",
  12226=>"110110110",
  12227=>"100111011",
  12228=>"001001001",
  12229=>"000000111",
  12230=>"101110011",
  12231=>"110011001",
  12232=>"000111001",
  12233=>"101001110",
  12234=>"111110100",
  12235=>"001001101",
  12236=>"001010100",
  12237=>"000110100",
  12238=>"000110010",
  12239=>"110111101",
  12240=>"001111111",
  12241=>"010010000",
  12242=>"110101001",
  12243=>"011111101",
  12244=>"000001111",
  12245=>"010000011",
  12246=>"101000010",
  12247=>"101001101",
  12248=>"101110110",
  12249=>"000000110",
  12250=>"011100000",
  12251=>"111110001",
  12252=>"000101101",
  12253=>"000111001",
  12254=>"000000000",
  12255=>"001111000",
  12256=>"001100011",
  12257=>"001000101",
  12258=>"011111000",
  12259=>"011011000",
  12260=>"011011000",
  12261=>"101000101",
  12262=>"100011001",
  12263=>"111100101",
  12264=>"100110011",
  12265=>"010111010",
  12266=>"011110000",
  12267=>"000001110",
  12268=>"001000001",
  12269=>"111011111",
  12270=>"110001111",
  12271=>"101011111",
  12272=>"100111110",
  12273=>"110110010",
  12274=>"110101010",
  12275=>"101100101",
  12276=>"101000111",
  12277=>"111100011",
  12278=>"110111101",
  12279=>"100100010",
  12280=>"100111110",
  12281=>"110100011",
  12282=>"111100100",
  12283=>"011001000",
  12284=>"010011000",
  12285=>"011101100",
  12286=>"100101010",
  12287=>"001110101",
  12288=>"010011010",
  12289=>"001011011",
  12290=>"000100111",
  12291=>"011111001",
  12292=>"010011110",
  12293=>"000100011",
  12294=>"011010110",
  12295=>"100000100",
  12296=>"000101001",
  12297=>"101111111",
  12298=>"100110100",
  12299=>"111001011",
  12300=>"111110000",
  12301=>"011000100",
  12302=>"110010110",
  12303=>"000000011",
  12304=>"001000011",
  12305=>"001001101",
  12306=>"110001001",
  12307=>"001101110",
  12308=>"111100110",
  12309=>"000100001",
  12310=>"001111100",
  12311=>"011011101",
  12312=>"011001100",
  12313=>"010111010",
  12314=>"011010011",
  12315=>"110110001",
  12316=>"001010110",
  12317=>"101111000",
  12318=>"111010100",
  12319=>"101011001",
  12320=>"100111110",
  12321=>"011100011",
  12322=>"001100010",
  12323=>"000101000",
  12324=>"011001100",
  12325=>"100110110",
  12326=>"011001111",
  12327=>"001011001",
  12328=>"001000010",
  12329=>"111011011",
  12330=>"111011000",
  12331=>"100100111",
  12332=>"011000111",
  12333=>"011000110",
  12334=>"010111110",
  12335=>"010111011",
  12336=>"110000000",
  12337=>"101101000",
  12338=>"111010110",
  12339=>"010011001",
  12340=>"100110111",
  12341=>"011110110",
  12342=>"001001010",
  12343=>"100101001",
  12344=>"010001011",
  12345=>"100100001",
  12346=>"011010110",
  12347=>"010100111",
  12348=>"110101111",
  12349=>"000101001",
  12350=>"100101000",
  12351=>"111001101",
  12352=>"110110110",
  12353=>"101001000",
  12354=>"010101001",
  12355=>"110010110",
  12356=>"011111101",
  12357=>"111000111",
  12358=>"000001001",
  12359=>"011011010",
  12360=>"101100101",
  12361=>"011100000",
  12362=>"101111001",
  12363=>"000001010",
  12364=>"011110011",
  12365=>"110101101",
  12366=>"110101000",
  12367=>"110001100",
  12368=>"110100101",
  12369=>"011111101",
  12370=>"101111110",
  12371=>"110101010",
  12372=>"010110101",
  12373=>"111110110",
  12374=>"111001000",
  12375=>"110111111",
  12376=>"101010110",
  12377=>"100101111",
  12378=>"110011000",
  12379=>"011000111",
  12380=>"100101110",
  12381=>"101111101",
  12382=>"000111000",
  12383=>"010101001",
  12384=>"000100010",
  12385=>"111011000",
  12386=>"000100101",
  12387=>"010111111",
  12388=>"000100001",
  12389=>"110010011",
  12390=>"010111101",
  12391=>"010000110",
  12392=>"111101101",
  12393=>"010101101",
  12394=>"110000010",
  12395=>"001101100",
  12396=>"010000010",
  12397=>"011001000",
  12398=>"111110110",
  12399=>"101110010",
  12400=>"100001010",
  12401=>"100101001",
  12402=>"010101001",
  12403=>"100001110",
  12404=>"010101111",
  12405=>"101111010",
  12406=>"110101011",
  12407=>"101010000",
  12408=>"001101010",
  12409=>"111110001",
  12410=>"111100010",
  12411=>"000001010",
  12412=>"011111011",
  12413=>"100100011",
  12414=>"100010010",
  12415=>"000010000",
  12416=>"011100000",
  12417=>"110100000",
  12418=>"100000111",
  12419=>"010011110",
  12420=>"000000101",
  12421=>"000100100",
  12422=>"001101011",
  12423=>"110110001",
  12424=>"001110000",
  12425=>"001001000",
  12426=>"101000111",
  12427=>"100010101",
  12428=>"110110000",
  12429=>"000011101",
  12430=>"011011011",
  12431=>"001000000",
  12432=>"110110000",
  12433=>"011100001",
  12434=>"010001001",
  12435=>"110101101",
  12436=>"011011001",
  12437=>"011011101",
  12438=>"001011010",
  12439=>"110000111",
  12440=>"000101000",
  12441=>"011101101",
  12442=>"001000010",
  12443=>"001101001",
  12444=>"111010100",
  12445=>"110101110",
  12446=>"111011010",
  12447=>"110111111",
  12448=>"110011000",
  12449=>"011010110",
  12450=>"000110011",
  12451=>"011101110",
  12452=>"011011000",
  12453=>"111001010",
  12454=>"010011010",
  12455=>"111011000",
  12456=>"111110010",
  12457=>"100000110",
  12458=>"111000101",
  12459=>"110010100",
  12460=>"001111100",
  12461=>"101101101",
  12462=>"100110001",
  12463=>"111100110",
  12464=>"000101100",
  12465=>"011011101",
  12466=>"100000010",
  12467=>"001110010",
  12468=>"100110111",
  12469=>"000011111",
  12470=>"101110100",
  12471=>"101100111",
  12472=>"100010101",
  12473=>"011001100",
  12474=>"111011111",
  12475=>"010111011",
  12476=>"011010011",
  12477=>"011011010",
  12478=>"111111110",
  12479=>"010001111",
  12480=>"011110101",
  12481=>"101000110",
  12482=>"110111001",
  12483=>"111101101",
  12484=>"100111011",
  12485=>"111111111",
  12486=>"111111000",
  12487=>"000010101",
  12488=>"101010111",
  12489=>"100100101",
  12490=>"001001101",
  12491=>"110101001",
  12492=>"100101010",
  12493=>"000110000",
  12494=>"001110011",
  12495=>"011110000",
  12496=>"001000000",
  12497=>"010110000",
  12498=>"010010011",
  12499=>"010011100",
  12500=>"010001111",
  12501=>"011101101",
  12502=>"111100100",
  12503=>"001001111",
  12504=>"000110101",
  12505=>"111010110",
  12506=>"011110011",
  12507=>"100111001",
  12508=>"101011100",
  12509=>"100001000",
  12510=>"001011100",
  12511=>"101111111",
  12512=>"010110011",
  12513=>"001110011",
  12514=>"001110001",
  12515=>"111001011",
  12516=>"111011010",
  12517=>"011100111",
  12518=>"010110101",
  12519=>"110101111",
  12520=>"010110010",
  12521=>"101011101",
  12522=>"111010000",
  12523=>"001111010",
  12524=>"101010001",
  12525=>"011011100",
  12526=>"001011010",
  12527=>"111100100",
  12528=>"111101000",
  12529=>"110011000",
  12530=>"111001100",
  12531=>"001010010",
  12532=>"101010100",
  12533=>"111100100",
  12534=>"001101011",
  12535=>"100000111",
  12536=>"000001101",
  12537=>"101001000",
  12538=>"100000100",
  12539=>"001111010",
  12540=>"101101110",
  12541=>"001001011",
  12542=>"110010101",
  12543=>"100100100",
  12544=>"110111100",
  12545=>"001000001",
  12546=>"100011111",
  12547=>"110111111",
  12548=>"001000010",
  12549=>"111100001",
  12550=>"101100111",
  12551=>"101011000",
  12552=>"111001111",
  12553=>"111111011",
  12554=>"010001111",
  12555=>"100111110",
  12556=>"011011100",
  12557=>"010001100",
  12558=>"000110010",
  12559=>"101100111",
  12560=>"110101010",
  12561=>"101011000",
  12562=>"100001101",
  12563=>"100101100",
  12564=>"111001100",
  12565=>"011100111",
  12566=>"000011110",
  12567=>"000000111",
  12568=>"111100101",
  12569=>"110101110",
  12570=>"000011110",
  12571=>"110000011",
  12572=>"110111010",
  12573=>"100000110",
  12574=>"000001111",
  12575=>"001000010",
  12576=>"000111100",
  12577=>"010011010",
  12578=>"010100101",
  12579=>"010011101",
  12580=>"011111000",
  12581=>"100000100",
  12582=>"000110010",
  12583=>"111000000",
  12584=>"101011000",
  12585=>"111111000",
  12586=>"010100110",
  12587=>"010100011",
  12588=>"011101000",
  12589=>"010101111",
  12590=>"000111100",
  12591=>"001101111",
  12592=>"000111100",
  12593=>"101010001",
  12594=>"101010001",
  12595=>"101101110",
  12596=>"111101100",
  12597=>"011111111",
  12598=>"100110111",
  12599=>"000100001",
  12600=>"000101011",
  12601=>"011111001",
  12602=>"010001110",
  12603=>"101100011",
  12604=>"110000001",
  12605=>"100011111",
  12606=>"001001011",
  12607=>"110010101",
  12608=>"111110101",
  12609=>"101111000",
  12610=>"001111011",
  12611=>"110010000",
  12612=>"000010100",
  12613=>"000000001",
  12614=>"000011100",
  12615=>"111001001",
  12616=>"110101101",
  12617=>"010100110",
  12618=>"101010010",
  12619=>"001100101",
  12620=>"100100110",
  12621=>"111011101",
  12622=>"001101001",
  12623=>"100011011",
  12624=>"001101100",
  12625=>"101001010",
  12626=>"100010111",
  12627=>"001010110",
  12628=>"101110011",
  12629=>"110010000",
  12630=>"010000101",
  12631=>"110000000",
  12632=>"000000101",
  12633=>"011111101",
  12634=>"110111100",
  12635=>"000001010",
  12636=>"011000111",
  12637=>"001001110",
  12638=>"111111011",
  12639=>"101111011",
  12640=>"001011001",
  12641=>"111000111",
  12642=>"011011011",
  12643=>"101110010",
  12644=>"001001101",
  12645=>"001001110",
  12646=>"101001011",
  12647=>"000100010",
  12648=>"111011100",
  12649=>"110110110",
  12650=>"000110011",
  12651=>"101110001",
  12652=>"001001001",
  12653=>"111101101",
  12654=>"000011000",
  12655=>"111111000",
  12656=>"110000111",
  12657=>"101100101",
  12658=>"000111000",
  12659=>"111110000",
  12660=>"110011100",
  12661=>"101111110",
  12662=>"100011101",
  12663=>"011111000",
  12664=>"011010011",
  12665=>"010101100",
  12666=>"101001000",
  12667=>"100000111",
  12668=>"110101001",
  12669=>"010000000",
  12670=>"000100010",
  12671=>"101111000",
  12672=>"111110001",
  12673=>"100010001",
  12674=>"100110111",
  12675=>"110111100",
  12676=>"011110000",
  12677=>"000111011",
  12678=>"010000001",
  12679=>"010110111",
  12680=>"011001100",
  12681=>"001110101",
  12682=>"000111111",
  12683=>"101100011",
  12684=>"001100001",
  12685=>"101100100",
  12686=>"101101010",
  12687=>"101101110",
  12688=>"101000000",
  12689=>"101111000",
  12690=>"111110100",
  12691=>"110101111",
  12692=>"110000100",
  12693=>"101100100",
  12694=>"010111110",
  12695=>"000011011",
  12696=>"111110011",
  12697=>"101101000",
  12698=>"111110011",
  12699=>"001011110",
  12700=>"110011000",
  12701=>"011110010",
  12702=>"000010110",
  12703=>"001000010",
  12704=>"011101011",
  12705=>"110111101",
  12706=>"100011111",
  12707=>"110110101",
  12708=>"110011001",
  12709=>"101001111",
  12710=>"000000111",
  12711=>"010111010",
  12712=>"111110111",
  12713=>"111011011",
  12714=>"111010010",
  12715=>"110010111",
  12716=>"001111111",
  12717=>"010000001",
  12718=>"000001110",
  12719=>"111010011",
  12720=>"011101011",
  12721=>"010011010",
  12722=>"000101110",
  12723=>"111111011",
  12724=>"110011111",
  12725=>"000010110",
  12726=>"011111111",
  12727=>"010000011",
  12728=>"010111111",
  12729=>"010100111",
  12730=>"000000100",
  12731=>"010101011",
  12732=>"111011011",
  12733=>"011111100",
  12734=>"001001101",
  12735=>"001100110",
  12736=>"110111010",
  12737=>"001011011",
  12738=>"101100000",
  12739=>"100010000",
  12740=>"111010100",
  12741=>"001001010",
  12742=>"001011111",
  12743=>"110111010",
  12744=>"101110110",
  12745=>"010010101",
  12746=>"101011001",
  12747=>"110111001",
  12748=>"111110100",
  12749=>"000011110",
  12750=>"101001110",
  12751=>"101010110",
  12752=>"011011011",
  12753=>"111011011",
  12754=>"011101001",
  12755=>"111000000",
  12756=>"010101011",
  12757=>"011010000",
  12758=>"010011101",
  12759=>"010111110",
  12760=>"111001100",
  12761=>"011001010",
  12762=>"011010001",
  12763=>"110101110",
  12764=>"000111110",
  12765=>"001000000",
  12766=>"010110101",
  12767=>"100100101",
  12768=>"111111001",
  12769=>"100110011",
  12770=>"000000001",
  12771=>"001011010",
  12772=>"100001100",
  12773=>"001110010",
  12774=>"001101111",
  12775=>"111001000",
  12776=>"110111110",
  12777=>"110000001",
  12778=>"101111000",
  12779=>"010100110",
  12780=>"011111111",
  12781=>"111010001",
  12782=>"101111101",
  12783=>"011000001",
  12784=>"111101101",
  12785=>"101111110",
  12786=>"100101001",
  12787=>"100100101",
  12788=>"011001111",
  12789=>"000001000",
  12790=>"111010001",
  12791=>"111101000",
  12792=>"000110010",
  12793=>"101111011",
  12794=>"000001110",
  12795=>"001001100",
  12796=>"101010110",
  12797=>"110001010",
  12798=>"000100000",
  12799=>"000001000",
  12800=>"011111000",
  12801=>"111011010",
  12802=>"001101101",
  12803=>"001111111",
  12804=>"011010110",
  12805=>"110100110",
  12806=>"010000011",
  12807=>"011110101",
  12808=>"001101111",
  12809=>"000011110",
  12810=>"100101011",
  12811=>"110110011",
  12812=>"000011010",
  12813=>"010001001",
  12814=>"000100110",
  12815=>"011000101",
  12816=>"100000111",
  12817=>"001100101",
  12818=>"000000010",
  12819=>"111001100",
  12820=>"110000010",
  12821=>"111011101",
  12822=>"111101011",
  12823=>"001101111",
  12824=>"111100000",
  12825=>"100010101",
  12826=>"110111101",
  12827=>"000110010",
  12828=>"001011011",
  12829=>"100001111",
  12830=>"000010110",
  12831=>"100110010",
  12832=>"011110111",
  12833=>"110001100",
  12834=>"111111100",
  12835=>"001010011",
  12836=>"111101111",
  12837=>"111001111",
  12838=>"001011100",
  12839=>"001011000",
  12840=>"001101101",
  12841=>"001001010",
  12842=>"110111100",
  12843=>"010011001",
  12844=>"000110011",
  12845=>"001000110",
  12846=>"001000000",
  12847=>"101001100",
  12848=>"100001001",
  12849=>"110001100",
  12850=>"011100110",
  12851=>"001101101",
  12852=>"111001100",
  12853=>"001011111",
  12854=>"111100000",
  12855=>"011000000",
  12856=>"101010111",
  12857=>"010010001",
  12858=>"111100111",
  12859=>"110100110",
  12860=>"110101011",
  12861=>"010001000",
  12862=>"011010100",
  12863=>"011000101",
  12864=>"101010011",
  12865=>"011000110",
  12866=>"010011000",
  12867=>"011001100",
  12868=>"110001110",
  12869=>"000110110",
  12870=>"110000100",
  12871=>"011111001",
  12872=>"000110001",
  12873=>"001010101",
  12874=>"010100110",
  12875=>"000011001",
  12876=>"111111001",
  12877=>"111111101",
  12878=>"010000101",
  12879=>"100001110",
  12880=>"100000010",
  12881=>"100000010",
  12882=>"101100101",
  12883=>"000111001",
  12884=>"111101000",
  12885=>"111000110",
  12886=>"110111110",
  12887=>"000001011",
  12888=>"000001000",
  12889=>"001000100",
  12890=>"000111011",
  12891=>"101000110",
  12892=>"111111110",
  12893=>"010001110",
  12894=>"100111110",
  12895=>"011001010",
  12896=>"100100110",
  12897=>"111111000",
  12898=>"101000110",
  12899=>"110000001",
  12900=>"001111000",
  12901=>"101100100",
  12902=>"001100101",
  12903=>"000010001",
  12904=>"111010010",
  12905=>"011011010",
  12906=>"110111110",
  12907=>"111010000",
  12908=>"000001011",
  12909=>"000010010",
  12910=>"000101001",
  12911=>"111101110",
  12912=>"110000000",
  12913=>"111101110",
  12914=>"101111011",
  12915=>"010100010",
  12916=>"011001001",
  12917=>"000001110",
  12918=>"000011110",
  12919=>"110000011",
  12920=>"111111110",
  12921=>"010011101",
  12922=>"100100010",
  12923=>"111110111",
  12924=>"110011001",
  12925=>"100010100",
  12926=>"100001111",
  12927=>"110000000",
  12928=>"110011001",
  12929=>"000101101",
  12930=>"111001011",
  12931=>"000001100",
  12932=>"101001111",
  12933=>"011000001",
  12934=>"010111110",
  12935=>"111101111",
  12936=>"101011111",
  12937=>"001000011",
  12938=>"110100000",
  12939=>"111100101",
  12940=>"001111110",
  12941=>"010101011",
  12942=>"110111100",
  12943=>"010101100",
  12944=>"111011110",
  12945=>"001011010",
  12946=>"000010111",
  12947=>"011100110",
  12948=>"001111010",
  12949=>"100011101",
  12950=>"010101011",
  12951=>"100111100",
  12952=>"000100001",
  12953=>"100001010",
  12954=>"011100000",
  12955=>"100001000",
  12956=>"011111111",
  12957=>"011011010",
  12958=>"111111100",
  12959=>"001010000",
  12960=>"100110001",
  12961=>"011011110",
  12962=>"010111000",
  12963=>"001000001",
  12964=>"011011000",
  12965=>"011001101",
  12966=>"001000111",
  12967=>"001000010",
  12968=>"111101110",
  12969=>"010111111",
  12970=>"111110111",
  12971=>"001111110",
  12972=>"111011111",
  12973=>"110110000",
  12974=>"011001111",
  12975=>"111110000",
  12976=>"110000111",
  12977=>"101101101",
  12978=>"111000101",
  12979=>"110111110",
  12980=>"110000000",
  12981=>"011100111",
  12982=>"111100100",
  12983=>"110100111",
  12984=>"001000101",
  12985=>"001000001",
  12986=>"101011011",
  12987=>"111011001",
  12988=>"101011011",
  12989=>"000100001",
  12990=>"101100001",
  12991=>"111100100",
  12992=>"010010000",
  12993=>"001001110",
  12994=>"111111111",
  12995=>"100011111",
  12996=>"110010100",
  12997=>"110110110",
  12998=>"111000010",
  12999=>"001111101",
  13000=>"011110110",
  13001=>"101110111",
  13002=>"000010110",
  13003=>"001111000",
  13004=>"001110110",
  13005=>"100000101",
  13006=>"100001110",
  13007=>"011000011",
  13008=>"111101110",
  13009=>"000000101",
  13010=>"010000100",
  13011=>"110110001",
  13012=>"000011111",
  13013=>"001111111",
  13014=>"010111111",
  13015=>"001000101",
  13016=>"011110110",
  13017=>"110101100",
  13018=>"010001001",
  13019=>"011001101",
  13020=>"100111110",
  13021=>"101101001",
  13022=>"111011010",
  13023=>"000100010",
  13024=>"111101111",
  13025=>"001110111",
  13026=>"001101111",
  13027=>"001010001",
  13028=>"111111011",
  13029=>"101001111",
  13030=>"111111001",
  13031=>"000110100",
  13032=>"011100010",
  13033=>"111110100",
  13034=>"110000010",
  13035=>"101100100",
  13036=>"110011100",
  13037=>"010001001",
  13038=>"101111110",
  13039=>"101000001",
  13040=>"110001000",
  13041=>"110001101",
  13042=>"110110101",
  13043=>"100000101",
  13044=>"000000111",
  13045=>"011101101",
  13046=>"111100011",
  13047=>"011000111",
  13048=>"100000011",
  13049=>"111111111",
  13050=>"010100010",
  13051=>"100101101",
  13052=>"001110111",
  13053=>"011101000",
  13054=>"110111011",
  13055=>"001000001",
  13056=>"111010011",
  13057=>"111000010",
  13058=>"111110000",
  13059=>"000110000",
  13060=>"001101000",
  13061=>"010011101",
  13062=>"100000000",
  13063=>"111101001",
  13064=>"010011100",
  13065=>"010110001",
  13066=>"110111001",
  13067=>"010111100",
  13068=>"000111010",
  13069=>"111100100",
  13070=>"110110110",
  13071=>"001110011",
  13072=>"101011100",
  13073=>"011010001",
  13074=>"010000110",
  13075=>"101111100",
  13076=>"010100000",
  13077=>"010110100",
  13078=>"001001101",
  13079=>"111101001",
  13080=>"110111001",
  13081=>"101110110",
  13082=>"010001000",
  13083=>"111111111",
  13084=>"101000000",
  13085=>"000100100",
  13086=>"001000101",
  13087=>"010110101",
  13088=>"111001111",
  13089=>"111000000",
  13090=>"010010010",
  13091=>"110111111",
  13092=>"011110000",
  13093=>"101011110",
  13094=>"000011010",
  13095=>"000110101",
  13096=>"110000101",
  13097=>"000101100",
  13098=>"110011000",
  13099=>"100011110",
  13100=>"111110000",
  13101=>"111001010",
  13102=>"111110010",
  13103=>"101001111",
  13104=>"011111111",
  13105=>"000110111",
  13106=>"111010111",
  13107=>"010000111",
  13108=>"010100010",
  13109=>"100001111",
  13110=>"101011011",
  13111=>"000000100",
  13112=>"100110011",
  13113=>"010100110",
  13114=>"010111010",
  13115=>"010101101",
  13116=>"001100011",
  13117=>"110110001",
  13118=>"000111000",
  13119=>"000110000",
  13120=>"110001101",
  13121=>"101100111",
  13122=>"110111110",
  13123=>"000000110",
  13124=>"001000111",
  13125=>"000000000",
  13126=>"100100010",
  13127=>"101010110",
  13128=>"010111011",
  13129=>"000100100",
  13130=>"011100101",
  13131=>"011100011",
  13132=>"111100110",
  13133=>"110000000",
  13134=>"011010111",
  13135=>"100110100",
  13136=>"110101110",
  13137=>"000011111",
  13138=>"011101001",
  13139=>"111000110",
  13140=>"011100000",
  13141=>"001000001",
  13142=>"111110100",
  13143=>"010000100",
  13144=>"111010111",
  13145=>"000110111",
  13146=>"111010101",
  13147=>"111000010",
  13148=>"010110110",
  13149=>"101010000",
  13150=>"110010010",
  13151=>"011111111",
  13152=>"100010000",
  13153=>"111001111",
  13154=>"101110100",
  13155=>"010101110",
  13156=>"011100000",
  13157=>"111110011",
  13158=>"100100001",
  13159=>"110000000",
  13160=>"011111110",
  13161=>"111000000",
  13162=>"001101010",
  13163=>"010010001",
  13164=>"110101110",
  13165=>"110010101",
  13166=>"000001111",
  13167=>"101110101",
  13168=>"101010011",
  13169=>"100000100",
  13170=>"110110000",
  13171=>"111111011",
  13172=>"111111001",
  13173=>"111001000",
  13174=>"101111001",
  13175=>"011111010",
  13176=>"010010111",
  13177=>"111100110",
  13178=>"100100010",
  13179=>"101000101",
  13180=>"110110111",
  13181=>"111011101",
  13182=>"111001110",
  13183=>"100100111",
  13184=>"111111010",
  13185=>"000100101",
  13186=>"100111011",
  13187=>"110101011",
  13188=>"101100000",
  13189=>"000111010",
  13190=>"010101010",
  13191=>"001110111",
  13192=>"110101010",
  13193=>"000101000",
  13194=>"111110111",
  13195=>"101110110",
  13196=>"011110000",
  13197=>"100011011",
  13198=>"101111001",
  13199=>"001010010",
  13200=>"010111110",
  13201=>"101001111",
  13202=>"001000111",
  13203=>"010000011",
  13204=>"111100110",
  13205=>"010110101",
  13206=>"100100000",
  13207=>"100011000",
  13208=>"110100101",
  13209=>"010111010",
  13210=>"010000000",
  13211=>"101011101",
  13212=>"101001011",
  13213=>"111011101",
  13214=>"000000011",
  13215=>"100110110",
  13216=>"110110110",
  13217=>"000011011",
  13218=>"110101110",
  13219=>"110010001",
  13220=>"001001010",
  13221=>"000011110",
  13222=>"000111110",
  13223=>"000101110",
  13224=>"111110010",
  13225=>"101011001",
  13226=>"100010111",
  13227=>"011000000",
  13228=>"001001100",
  13229=>"001101000",
  13230=>"110110101",
  13231=>"000001111",
  13232=>"110101111",
  13233=>"000010110",
  13234=>"000001110",
  13235=>"011000001",
  13236=>"010000101",
  13237=>"000101111",
  13238=>"001000010",
  13239=>"001100000",
  13240=>"110001011",
  13241=>"100101010",
  13242=>"001101010",
  13243=>"111010111",
  13244=>"001001100",
  13245=>"000000000",
  13246=>"000001000",
  13247=>"010001100",
  13248=>"000100110",
  13249=>"000000100",
  13250=>"000110000",
  13251=>"001011010",
  13252=>"111011101",
  13253=>"100010111",
  13254=>"110001100",
  13255=>"110001100",
  13256=>"001001001",
  13257=>"010100100",
  13258=>"000110100",
  13259=>"111010010",
  13260=>"010000001",
  13261=>"000001110",
  13262=>"101010111",
  13263=>"000010100",
  13264=>"000110100",
  13265=>"110111011",
  13266=>"011001111",
  13267=>"101001000",
  13268=>"001111111",
  13269=>"110100000",
  13270=>"101100111",
  13271=>"101100101",
  13272=>"000010101",
  13273=>"110011001",
  13274=>"011100101",
  13275=>"111110001",
  13276=>"011100010",
  13277=>"000000000",
  13278=>"010111111",
  13279=>"111000001",
  13280=>"101100000",
  13281=>"111111101",
  13282=>"110000100",
  13283=>"110101011",
  13284=>"100111100",
  13285=>"101011001",
  13286=>"111110100",
  13287=>"000000001",
  13288=>"000110010",
  13289=>"000011010",
  13290=>"110101011",
  13291=>"011010101",
  13292=>"101110110",
  13293=>"110101001",
  13294=>"100000110",
  13295=>"101111111",
  13296=>"111100010",
  13297=>"001011010",
  13298=>"110101101",
  13299=>"010111001",
  13300=>"011111111",
  13301=>"111101001",
  13302=>"111011010",
  13303=>"010100100",
  13304=>"011100100",
  13305=>"101000101",
  13306=>"100100001",
  13307=>"111101010",
  13308=>"110001010",
  13309=>"001011110",
  13310=>"111101101",
  13311=>"011010001",
  13312=>"000001100",
  13313=>"110111001",
  13314=>"111010011",
  13315=>"000100100",
  13316=>"001101100",
  13317=>"101001111",
  13318=>"010001000",
  13319=>"011101100",
  13320=>"010111111",
  13321=>"001110011",
  13322=>"001011101",
  13323=>"001001010",
  13324=>"011011110",
  13325=>"000100111",
  13326=>"101101010",
  13327=>"000001011",
  13328=>"110110111",
  13329=>"011011000",
  13330=>"111111110",
  13331=>"011000101",
  13332=>"000100110",
  13333=>"100110111",
  13334=>"000000101",
  13335=>"101101010",
  13336=>"111110010",
  13337=>"001100010",
  13338=>"111111001",
  13339=>"101100110",
  13340=>"001000010",
  13341=>"000111000",
  13342=>"001001001",
  13343=>"011011101",
  13344=>"111111111",
  13345=>"101010010",
  13346=>"011000100",
  13347=>"001100111",
  13348=>"011000011",
  13349=>"111011111",
  13350=>"000011011",
  13351=>"001000100",
  13352=>"110000111",
  13353=>"000011000",
  13354=>"100000100",
  13355=>"001010001",
  13356=>"000001000",
  13357=>"101011000",
  13358=>"101100010",
  13359=>"100010110",
  13360=>"100001111",
  13361=>"011101010",
  13362=>"101111001",
  13363=>"110100000",
  13364=>"011101100",
  13365=>"111100001",
  13366=>"111011001",
  13367=>"110110111",
  13368=>"101111100",
  13369=>"000000011",
  13370=>"110111101",
  13371=>"100000110",
  13372=>"001010101",
  13373=>"100010001",
  13374=>"000110101",
  13375=>"001110111",
  13376=>"101001010",
  13377=>"000100000",
  13378=>"000011100",
  13379=>"110101001",
  13380=>"010001000",
  13381=>"100110011",
  13382=>"100011100",
  13383=>"011101001",
  13384=>"111100111",
  13385=>"010011000",
  13386=>"111010110",
  13387=>"010010000",
  13388=>"001101010",
  13389=>"010101011",
  13390=>"111110001",
  13391=>"101101000",
  13392=>"101100011",
  13393=>"110000000",
  13394=>"011001011",
  13395=>"001010010",
  13396=>"011111101",
  13397=>"111101000",
  13398=>"010010010",
  13399=>"001011001",
  13400=>"101110010",
  13401=>"000101001",
  13402=>"010111000",
  13403=>"001000001",
  13404=>"110000111",
  13405=>"000110000",
  13406=>"000111100",
  13407=>"100001110",
  13408=>"110000101",
  13409=>"001001000",
  13410=>"011010110",
  13411=>"001001111",
  13412=>"110010001",
  13413=>"000111011",
  13414=>"001111001",
  13415=>"011111100",
  13416=>"111111100",
  13417=>"111010101",
  13418=>"000001111",
  13419=>"101001100",
  13420=>"111110101",
  13421=>"110100111",
  13422=>"111011010",
  13423=>"100010110",
  13424=>"000001000",
  13425=>"111011010",
  13426=>"011110100",
  13427=>"000000111",
  13428=>"010011100",
  13429=>"000001010",
  13430=>"101100100",
  13431=>"001000100",
  13432=>"000000010",
  13433=>"001110010",
  13434=>"011100011",
  13435=>"000011010",
  13436=>"001100111",
  13437=>"100011101",
  13438=>"001101000",
  13439=>"111111110",
  13440=>"110000110",
  13441=>"111111011",
  13442=>"110000000",
  13443=>"110111100",
  13444=>"010001101",
  13445=>"100000110",
  13446=>"011011100",
  13447=>"010010101",
  13448=>"001011000",
  13449=>"101000101",
  13450=>"010001111",
  13451=>"100110010",
  13452=>"001011010",
  13453=>"111101111",
  13454=>"001011100",
  13455=>"110010001",
  13456=>"101010000",
  13457=>"100111001",
  13458=>"110011001",
  13459=>"001000101",
  13460=>"011111000",
  13461=>"000110111",
  13462=>"100100001",
  13463=>"101110111",
  13464=>"100110000",
  13465=>"000000110",
  13466=>"101011101",
  13467=>"011011010",
  13468=>"000001011",
  13469=>"000011001",
  13470=>"111001001",
  13471=>"111111100",
  13472=>"011100111",
  13473=>"010000110",
  13474=>"100110001",
  13475=>"000001010",
  13476=>"011000001",
  13477=>"000010000",
  13478=>"010010001",
  13479=>"000110010",
  13480=>"010100010",
  13481=>"111000000",
  13482=>"111001110",
  13483=>"111101001",
  13484=>"111110110",
  13485=>"001000100",
  13486=>"100111110",
  13487=>"111111010",
  13488=>"001000010",
  13489=>"001101111",
  13490=>"110010100",
  13491=>"111111110",
  13492=>"111000110",
  13493=>"010010011",
  13494=>"000111111",
  13495=>"110101000",
  13496=>"100111010",
  13497=>"001001001",
  13498=>"110100100",
  13499=>"111100101",
  13500=>"101011100",
  13501=>"100000011",
  13502=>"011010010",
  13503=>"110111011",
  13504=>"011101110",
  13505=>"010110101",
  13506=>"111001110",
  13507=>"011100111",
  13508=>"110110110",
  13509=>"011010110",
  13510=>"101111111",
  13511=>"001110111",
  13512=>"011010111",
  13513=>"110001000",
  13514=>"010010110",
  13515=>"101110011",
  13516=>"111111111",
  13517=>"010101100",
  13518=>"010010001",
  13519=>"111000011",
  13520=>"110110110",
  13521=>"101010001",
  13522=>"000010001",
  13523=>"000100001",
  13524=>"011100001",
  13525=>"001000101",
  13526=>"100011100",
  13527=>"110101110",
  13528=>"000010000",
  13529=>"010010001",
  13530=>"000010111",
  13531=>"000010010",
  13532=>"010010101",
  13533=>"101100010",
  13534=>"011100111",
  13535=>"110010001",
  13536=>"010001001",
  13537=>"001011011",
  13538=>"001000100",
  13539=>"001110001",
  13540=>"100010110",
  13541=>"000000000",
  13542=>"100000001",
  13543=>"100101000",
  13544=>"110000011",
  13545=>"100001100",
  13546=>"010110110",
  13547=>"000000001",
  13548=>"011011011",
  13549=>"100110000",
  13550=>"001001100",
  13551=>"101000000",
  13552=>"001000001",
  13553=>"000100010",
  13554=>"001100101",
  13555=>"001001000",
  13556=>"010010011",
  13557=>"101000111",
  13558=>"100010010",
  13559=>"001001110",
  13560=>"010010111",
  13561=>"001001010",
  13562=>"110001000",
  13563=>"111011010",
  13564=>"111000110",
  13565=>"011011011",
  13566=>"010100111",
  13567=>"011101111",
  13568=>"100110110",
  13569=>"100000010",
  13570=>"111001011",
  13571=>"110101000",
  13572=>"001101100",
  13573=>"011000000",
  13574=>"100001000",
  13575=>"100111101",
  13576=>"000101001",
  13577=>"110011001",
  13578=>"001110111",
  13579=>"000110101",
  13580=>"110010011",
  13581=>"111100111",
  13582=>"111101010",
  13583=>"011010110",
  13584=>"111001111",
  13585=>"010001101",
  13586=>"101111110",
  13587=>"100111001",
  13588=>"110100101",
  13589=>"001011000",
  13590=>"011000100",
  13591=>"011110110",
  13592=>"111001111",
  13593=>"010001000",
  13594=>"100100101",
  13595=>"111000001",
  13596=>"011000110",
  13597=>"100100000",
  13598=>"100101000",
  13599=>"101001111",
  13600=>"000000110",
  13601=>"001100110",
  13602=>"000111000",
  13603=>"100001111",
  13604=>"111010100",
  13605=>"101011011",
  13606=>"011011010",
  13607=>"100111111",
  13608=>"000101010",
  13609=>"011000110",
  13610=>"111110001",
  13611=>"000110100",
  13612=>"001111010",
  13613=>"100000101",
  13614=>"000000110",
  13615=>"110011000",
  13616=>"010011111",
  13617=>"111100000",
  13618=>"000101011",
  13619=>"100000000",
  13620=>"101000010",
  13621=>"010100111",
  13622=>"101101000",
  13623=>"111101010",
  13624=>"100000000",
  13625=>"001101111",
  13626=>"001010101",
  13627=>"101110111",
  13628=>"100000110",
  13629=>"000101000",
  13630=>"000000010",
  13631=>"011011001",
  13632=>"001100000",
  13633=>"101000110",
  13634=>"010100000",
  13635=>"111111010",
  13636=>"010101000",
  13637=>"011001111",
  13638=>"110100010",
  13639=>"100111000",
  13640=>"111101000",
  13641=>"100101110",
  13642=>"100010011",
  13643=>"010010010",
  13644=>"111011011",
  13645=>"111011011",
  13646=>"101011010",
  13647=>"101111010",
  13648=>"111010110",
  13649=>"110100001",
  13650=>"111101010",
  13651=>"100011101",
  13652=>"000010000",
  13653=>"001011110",
  13654=>"111001011",
  13655=>"001111100",
  13656=>"101000001",
  13657=>"100100101",
  13658=>"110010011",
  13659=>"110000011",
  13660=>"101110110",
  13661=>"101110000",
  13662=>"010001010",
  13663=>"000011010",
  13664=>"011111101",
  13665=>"110010111",
  13666=>"001011010",
  13667=>"100001110",
  13668=>"100101110",
  13669=>"000110111",
  13670=>"101100011",
  13671=>"000000101",
  13672=>"110001101",
  13673=>"110101001",
  13674=>"100001011",
  13675=>"101101101",
  13676=>"011000010",
  13677=>"101111110",
  13678=>"001010000",
  13679=>"111110001",
  13680=>"111011001",
  13681=>"101011110",
  13682=>"011000000",
  13683=>"111100010",
  13684=>"011010111",
  13685=>"010100011",
  13686=>"010110000",
  13687=>"110000000",
  13688=>"010111100",
  13689=>"001111001",
  13690=>"011111011",
  13691=>"011001001",
  13692=>"011110011",
  13693=>"100011010",
  13694=>"110101000",
  13695=>"010101111",
  13696=>"000001011",
  13697=>"011010110",
  13698=>"100100000",
  13699=>"100101000",
  13700=>"010000111",
  13701=>"101000010",
  13702=>"101000110",
  13703=>"001010001",
  13704=>"111110110",
  13705=>"100010100",
  13706=>"100001101",
  13707=>"011010000",
  13708=>"001110010",
  13709=>"110001000",
  13710=>"001100000",
  13711=>"001110011",
  13712=>"001110111",
  13713=>"001001100",
  13714=>"011000010",
  13715=>"100110001",
  13716=>"100110111",
  13717=>"001101100",
  13718=>"011000010",
  13719=>"111111100",
  13720=>"101100001",
  13721=>"001001011",
  13722=>"001111101",
  13723=>"011011000",
  13724=>"011010010",
  13725=>"110100110",
  13726=>"100010001",
  13727=>"010111101",
  13728=>"101001001",
  13729=>"101110100",
  13730=>"000101011",
  13731=>"000001100",
  13732=>"110100010",
  13733=>"010010010",
  13734=>"000101101",
  13735=>"100101011",
  13736=>"111100110",
  13737=>"110010111",
  13738=>"001011010",
  13739=>"010101010",
  13740=>"100000010",
  13741=>"100000001",
  13742=>"001000001",
  13743=>"001101110",
  13744=>"111010010",
  13745=>"011011001",
  13746=>"011100011",
  13747=>"011011010",
  13748=>"010010110",
  13749=>"111110010",
  13750=>"000001011",
  13751=>"110011101",
  13752=>"101010100",
  13753=>"101010100",
  13754=>"000000001",
  13755=>"001111101",
  13756=>"111110100",
  13757=>"110000010",
  13758=>"111101011",
  13759=>"000110110",
  13760=>"100100100",
  13761=>"001001111",
  13762=>"001101001",
  13763=>"110111101",
  13764=>"000000011",
  13765=>"000000101",
  13766=>"110000101",
  13767=>"000110001",
  13768=>"010011110",
  13769=>"000000000",
  13770=>"110000100",
  13771=>"001100010",
  13772=>"001100011",
  13773=>"000010000",
  13774=>"110000101",
  13775=>"001001010",
  13776=>"000100010",
  13777=>"010010000",
  13778=>"001011100",
  13779=>"111111010",
  13780=>"111101010",
  13781=>"011100000",
  13782=>"101111010",
  13783=>"011001011",
  13784=>"011001001",
  13785=>"111111010",
  13786=>"101011001",
  13787=>"111101111",
  13788=>"000000100",
  13789=>"011111111",
  13790=>"001110111",
  13791=>"111111000",
  13792=>"001111000",
  13793=>"010100100",
  13794=>"111110000",
  13795=>"011011001",
  13796=>"110111110",
  13797=>"010011000",
  13798=>"111111100",
  13799=>"001010010",
  13800=>"010011010",
  13801=>"111110000",
  13802=>"010110010",
  13803=>"011101100",
  13804=>"100001101",
  13805=>"011101010",
  13806=>"001011001",
  13807=>"110111111",
  13808=>"111000111",
  13809=>"000111110",
  13810=>"010010101",
  13811=>"001101001",
  13812=>"101011000",
  13813=>"110000111",
  13814=>"110011101",
  13815=>"110011110",
  13816=>"000100100",
  13817=>"111001000",
  13818=>"000110011",
  13819=>"101001111",
  13820=>"000001111",
  13821=>"000110111",
  13822=>"101111011",
  13823=>"011000001",
  13824=>"111101100",
  13825=>"110110111",
  13826=>"001000101",
  13827=>"011101000",
  13828=>"010110010",
  13829=>"111000000",
  13830=>"001000010",
  13831=>"100010010",
  13832=>"100101111",
  13833=>"110000010",
  13834=>"001101110",
  13835=>"011000000",
  13836=>"110110011",
  13837=>"110101010",
  13838=>"111001000",
  13839=>"100110010",
  13840=>"111001100",
  13841=>"111100110",
  13842=>"110110000",
  13843=>"101111000",
  13844=>"010001000",
  13845=>"101011000",
  13846=>"011111000",
  13847=>"110110001",
  13848=>"001001000",
  13849=>"011011100",
  13850=>"010101101",
  13851=>"001110101",
  13852=>"111001000",
  13853=>"110100110",
  13854=>"100011000",
  13855=>"000100100",
  13856=>"011011011",
  13857=>"000001110",
  13858=>"001111011",
  13859=>"100100111",
  13860=>"010000000",
  13861=>"011000100",
  13862=>"111101000",
  13863=>"011101101",
  13864=>"010010000",
  13865=>"101110111",
  13866=>"001001100",
  13867=>"001100000",
  13868=>"010110011",
  13869=>"101011110",
  13870=>"000000101",
  13871=>"001011000",
  13872=>"111010001",
  13873=>"111011010",
  13874=>"111101001",
  13875=>"111011001",
  13876=>"000001110",
  13877=>"010011000",
  13878=>"110011111",
  13879=>"100101110",
  13880=>"011101110",
  13881=>"111111010",
  13882=>"010010000",
  13883=>"001000010",
  13884=>"110000001",
  13885=>"110010010",
  13886=>"101000110",
  13887=>"010111000",
  13888=>"011100000",
  13889=>"011110111",
  13890=>"011101010",
  13891=>"110011110",
  13892=>"011010010",
  13893=>"000011100",
  13894=>"001001001",
  13895=>"010111110",
  13896=>"001110111",
  13897=>"100101010",
  13898=>"001110001",
  13899=>"000111000",
  13900=>"100111110",
  13901=>"001100000",
  13902=>"000001010",
  13903=>"001111010",
  13904=>"101011010",
  13905=>"000111110",
  13906=>"101110111",
  13907=>"010000011",
  13908=>"010000111",
  13909=>"000110010",
  13910=>"001011100",
  13911=>"001110000",
  13912=>"000000000",
  13913=>"000001001",
  13914=>"101101100",
  13915=>"001101110",
  13916=>"001100011",
  13917=>"101001000",
  13918=>"101011001",
  13919=>"100110001",
  13920=>"111100111",
  13921=>"101101011",
  13922=>"011110001",
  13923=>"000000111",
  13924=>"101110110",
  13925=>"101100100",
  13926=>"110110100",
  13927=>"011011011",
  13928=>"000000000",
  13929=>"101000010",
  13930=>"110000101",
  13931=>"101001100",
  13932=>"011001011",
  13933=>"001000100",
  13934=>"111010111",
  13935=>"111110000",
  13936=>"110110000",
  13937=>"000100111",
  13938=>"111001000",
  13939=>"000001101",
  13940=>"101010111",
  13941=>"100111101",
  13942=>"111010010",
  13943=>"011100100",
  13944=>"111100100",
  13945=>"001010011",
  13946=>"111000010",
  13947=>"001000011",
  13948=>"000000011",
  13949=>"000010000",
  13950=>"000110100",
  13951=>"111100101",
  13952=>"001011001",
  13953=>"100011011",
  13954=>"111011001",
  13955=>"001000110",
  13956=>"100111001",
  13957=>"111000011",
  13958=>"111100111",
  13959=>"100100010",
  13960=>"110111000",
  13961=>"010110101",
  13962=>"011110110",
  13963=>"010001011",
  13964=>"111100001",
  13965=>"001001010",
  13966=>"111110100",
  13967=>"110000100",
  13968=>"000100010",
  13969=>"011000111",
  13970=>"110001010",
  13971=>"011111010",
  13972=>"100001100",
  13973=>"101100101",
  13974=>"000100011",
  13975=>"110001111",
  13976=>"100110100",
  13977=>"010011101",
  13978=>"100100001",
  13979=>"000000010",
  13980=>"011100101",
  13981=>"000011011",
  13982=>"110011001",
  13983=>"111110100",
  13984=>"001001001",
  13985=>"111000110",
  13986=>"100011011",
  13987=>"100010011",
  13988=>"001011101",
  13989=>"000110000",
  13990=>"001100110",
  13991=>"100000100",
  13992=>"000111010",
  13993=>"011111010",
  13994=>"111000111",
  13995=>"100110000",
  13996=>"100010000",
  13997=>"100101100",
  13998=>"010111000",
  13999=>"001001111",
  14000=>"000100101",
  14001=>"000101010",
  14002=>"100101010",
  14003=>"001010000",
  14004=>"110000100",
  14005=>"010101111",
  14006=>"000001000",
  14007=>"011011010",
  14008=>"101110010",
  14009=>"001010101",
  14010=>"100010111",
  14011=>"001111000",
  14012=>"010010000",
  14013=>"001011010",
  14014=>"001000001",
  14015=>"000100111",
  14016=>"101111000",
  14017=>"010101110",
  14018=>"100010100",
  14019=>"111110011",
  14020=>"100011001",
  14021=>"000100011",
  14022=>"011000000",
  14023=>"001001001",
  14024=>"010101010",
  14025=>"001000011",
  14026=>"011111001",
  14027=>"100001100",
  14028=>"000110101",
  14029=>"000101011",
  14030=>"011000011",
  14031=>"011001000",
  14032=>"110000011",
  14033=>"000100110",
  14034=>"110100000",
  14035=>"110000000",
  14036=>"110010111",
  14037=>"100000101",
  14038=>"110011111",
  14039=>"100010001",
  14040=>"011010000",
  14041=>"110111111",
  14042=>"000100101",
  14043=>"101101111",
  14044=>"100100001",
  14045=>"001100110",
  14046=>"111111100",
  14047=>"100111110",
  14048=>"001000111",
  14049=>"000001100",
  14050=>"111010001",
  14051=>"111001011",
  14052=>"001010010",
  14053=>"011111110",
  14054=>"010110001",
  14055=>"011000001",
  14056=>"001111110",
  14057=>"111101111",
  14058=>"110111011",
  14059=>"000100110",
  14060=>"001000000",
  14061=>"111000101",
  14062=>"101001111",
  14063=>"101110110",
  14064=>"010110001",
  14065=>"011001000",
  14066=>"110100100",
  14067=>"011011100",
  14068=>"010100010",
  14069=>"111111111",
  14070=>"011110100",
  14071=>"011110011",
  14072=>"101011000",
  14073=>"100100101",
  14074=>"111001111",
  14075=>"100110000",
  14076=>"101011000",
  14077=>"011000001",
  14078=>"101010000",
  14079=>"010110011",
  14080=>"011000101",
  14081=>"110011110",
  14082=>"001000110",
  14083=>"001100101",
  14084=>"100011110",
  14085=>"000010001",
  14086=>"110111111",
  14087=>"111100111",
  14088=>"100001000",
  14089=>"111001100",
  14090=>"111010100",
  14091=>"101101001",
  14092=>"111000011",
  14093=>"111111111",
  14094=>"111010101",
  14095=>"111111011",
  14096=>"000111101",
  14097=>"011010000",
  14098=>"001110111",
  14099=>"011011011",
  14100=>"001101101",
  14101=>"101001001",
  14102=>"000000110",
  14103=>"111010010",
  14104=>"101111100",
  14105=>"011011001",
  14106=>"101110111",
  14107=>"011001000",
  14108=>"111110010",
  14109=>"100010110",
  14110=>"100101010",
  14111=>"110111001",
  14112=>"000100101",
  14113=>"001001110",
  14114=>"100100111",
  14115=>"100111011",
  14116=>"000011111",
  14117=>"101011000",
  14118=>"001000111",
  14119=>"000011101",
  14120=>"011010010",
  14121=>"101011100",
  14122=>"000111010",
  14123=>"010100110",
  14124=>"110110110",
  14125=>"001011110",
  14126=>"000101100",
  14127=>"010010011",
  14128=>"100010101",
  14129=>"001111101",
  14130=>"000010111",
  14131=>"010101011",
  14132=>"111011101",
  14133=>"011100010",
  14134=>"000110011",
  14135=>"000010100",
  14136=>"011110111",
  14137=>"111010010",
  14138=>"101010111",
  14139=>"000011001",
  14140=>"101111001",
  14141=>"011001011",
  14142=>"111000011",
  14143=>"000010110",
  14144=>"110000101",
  14145=>"100110101",
  14146=>"001001001",
  14147=>"010100010",
  14148=>"110011001",
  14149=>"001010001",
  14150=>"010101010",
  14151=>"011000101",
  14152=>"011000110",
  14153=>"000101011",
  14154=>"001101000",
  14155=>"010000001",
  14156=>"001111011",
  14157=>"011011010",
  14158=>"101110011",
  14159=>"110001000",
  14160=>"111011000",
  14161=>"001010111",
  14162=>"001000111",
  14163=>"110001010",
  14164=>"001001011",
  14165=>"000101000",
  14166=>"101100101",
  14167=>"100011111",
  14168=>"011000001",
  14169=>"000000101",
  14170=>"111010110",
  14171=>"000000110",
  14172=>"010111101",
  14173=>"001101110",
  14174=>"101000001",
  14175=>"000010010",
  14176=>"010011010",
  14177=>"000010010",
  14178=>"001011000",
  14179=>"101100010",
  14180=>"011010001",
  14181=>"001010010",
  14182=>"100101110",
  14183=>"001101110",
  14184=>"000010010",
  14185=>"000010110",
  14186=>"010010000",
  14187=>"110100011",
  14188=>"111100101",
  14189=>"001110000",
  14190=>"001001011",
  14191=>"111100111",
  14192=>"100110001",
  14193=>"100110001",
  14194=>"101101011",
  14195=>"111001010",
  14196=>"101001011",
  14197=>"000100010",
  14198=>"100001011",
  14199=>"100110000",
  14200=>"000001101",
  14201=>"011110110",
  14202=>"101111011",
  14203=>"000110111",
  14204=>"000010000",
  14205=>"111000110",
  14206=>"100011001",
  14207=>"110011101",
  14208=>"110111010",
  14209=>"110000111",
  14210=>"111101000",
  14211=>"000110000",
  14212=>"010011110",
  14213=>"101000011",
  14214=>"101001111",
  14215=>"001101110",
  14216=>"111110010",
  14217=>"110100110",
  14218=>"110001101",
  14219=>"010000000",
  14220=>"110101110",
  14221=>"111001101",
  14222=>"000111000",
  14223=>"011100111",
  14224=>"010111100",
  14225=>"110111111",
  14226=>"011010000",
  14227=>"111001000",
  14228=>"010011101",
  14229=>"010101001",
  14230=>"011011011",
  14231=>"100100001",
  14232=>"011100111",
  14233=>"100000010",
  14234=>"010000000",
  14235=>"010110110",
  14236=>"001100101",
  14237=>"011110011",
  14238=>"101100000",
  14239=>"111110110",
  14240=>"001111101",
  14241=>"111101001",
  14242=>"001111010",
  14243=>"000000000",
  14244=>"110011010",
  14245=>"110101111",
  14246=>"010101110",
  14247=>"011011111",
  14248=>"110110001",
  14249=>"000010111",
  14250=>"110010000",
  14251=>"111100101",
  14252=>"011100110",
  14253=>"101000100",
  14254=>"100100110",
  14255=>"111110000",
  14256=>"000001001",
  14257=>"101111010",
  14258=>"001100100",
  14259=>"111011001",
  14260=>"000110010",
  14261=>"111110111",
  14262=>"101010110",
  14263=>"000001011",
  14264=>"101010100",
  14265=>"001101000",
  14266=>"110010110",
  14267=>"001110011",
  14268=>"010101101",
  14269=>"110010011",
  14270=>"000000100",
  14271=>"101101100",
  14272=>"110101100",
  14273=>"100110111",
  14274=>"101111111",
  14275=>"111101111",
  14276=>"100001011",
  14277=>"100000100",
  14278=>"111111001",
  14279=>"111101000",
  14280=>"000000000",
  14281=>"101011010",
  14282=>"111110110",
  14283=>"100100010",
  14284=>"000001101",
  14285=>"000000000",
  14286=>"000100001",
  14287=>"000110010",
  14288=>"111111110",
  14289=>"111001100",
  14290=>"010100010",
  14291=>"101100010",
  14292=>"001001100",
  14293=>"111010111",
  14294=>"011001001",
  14295=>"000011001",
  14296=>"101001100",
  14297=>"000001110",
  14298=>"010011110",
  14299=>"111010101",
  14300=>"110100001",
  14301=>"010000011",
  14302=>"101111110",
  14303=>"110000000",
  14304=>"001100111",
  14305=>"100111110",
  14306=>"110010101",
  14307=>"111010101",
  14308=>"001001011",
  14309=>"100001100",
  14310=>"111011000",
  14311=>"111100000",
  14312=>"010111101",
  14313=>"110110010",
  14314=>"110000011",
  14315=>"001101000",
  14316=>"011010100",
  14317=>"101001000",
  14318=>"100110111",
  14319=>"001101010",
  14320=>"001101101",
  14321=>"011000000",
  14322=>"110000110",
  14323=>"000100000",
  14324=>"110010000",
  14325=>"101010000",
  14326=>"000100101",
  14327=>"001010010",
  14328=>"010111010",
  14329=>"111001010",
  14330=>"110100010",
  14331=>"111101010",
  14332=>"100011010",
  14333=>"100011010",
  14334=>"100010010",
  14335=>"100010000",
  14336=>"001010010",
  14337=>"001001101",
  14338=>"011101100",
  14339=>"011111010",
  14340=>"100100000",
  14341=>"011110101",
  14342=>"001101111",
  14343=>"000110010",
  14344=>"011000111",
  14345=>"010110101",
  14346=>"101011111",
  14347=>"010001001",
  14348=>"001000001",
  14349=>"100100000",
  14350=>"001100110",
  14351=>"111111001",
  14352=>"110110100",
  14353=>"011001010",
  14354=>"011101011",
  14355=>"111101110",
  14356=>"111100011",
  14357=>"100011100",
  14358=>"110011101",
  14359=>"011010001",
  14360=>"001100010",
  14361=>"101000000",
  14362=>"011101011",
  14363=>"111000010",
  14364=>"110011101",
  14365=>"011010011",
  14366=>"100110100",
  14367=>"110110110",
  14368=>"010011001",
  14369=>"100010110",
  14370=>"011000100",
  14371=>"011000100",
  14372=>"001010000",
  14373=>"001101010",
  14374=>"100111010",
  14375=>"110011110",
  14376=>"100100101",
  14377=>"000011110",
  14378=>"000111110",
  14379=>"000000101",
  14380=>"011000110",
  14381=>"111111001",
  14382=>"111000111",
  14383=>"011001100",
  14384=>"011000001",
  14385=>"101001101",
  14386=>"110001001",
  14387=>"000000011",
  14388=>"011000010",
  14389=>"110111100",
  14390=>"100100011",
  14391=>"010001100",
  14392=>"000001010",
  14393=>"110111100",
  14394=>"101110110",
  14395=>"110001011",
  14396=>"101010111",
  14397=>"101100100",
  14398=>"011110011",
  14399=>"100110001",
  14400=>"000001100",
  14401=>"010010010",
  14402=>"001000010",
  14403=>"100011111",
  14404=>"110101001",
  14405=>"111111100",
  14406=>"100100101",
  14407=>"001010010",
  14408=>"011100000",
  14409=>"011001001",
  14410=>"100100010",
  14411=>"000010011",
  14412=>"000001111",
  14413=>"110110101",
  14414=>"010000111",
  14415=>"011001010",
  14416=>"111101011",
  14417=>"001111000",
  14418=>"011001111",
  14419=>"110011010",
  14420=>"001110111",
  14421=>"010010011",
  14422=>"110010110",
  14423=>"011100010",
  14424=>"011111101",
  14425=>"001010110",
  14426=>"110100110",
  14427=>"100010010",
  14428=>"100000110",
  14429=>"100011110",
  14430=>"101001000",
  14431=>"111000001",
  14432=>"111111011",
  14433=>"111101100",
  14434=>"000000010",
  14435=>"011111110",
  14436=>"110111000",
  14437=>"001000101",
  14438=>"010000010",
  14439=>"100011010",
  14440=>"011111100",
  14441=>"010010100",
  14442=>"000100100",
  14443=>"001111110",
  14444=>"100100000",
  14445=>"111111101",
  14446=>"010101101",
  14447=>"000100100",
  14448=>"001010110",
  14449=>"111111111",
  14450=>"010100111",
  14451=>"011010101",
  14452=>"000010101",
  14453=>"101011101",
  14454=>"100001001",
  14455=>"101000111",
  14456=>"111111101",
  14457=>"010100111",
  14458=>"100100111",
  14459=>"110101110",
  14460=>"011010001",
  14461=>"100010011",
  14462=>"000011110",
  14463=>"001101010",
  14464=>"100010001",
  14465=>"101011100",
  14466=>"010111110",
  14467=>"111111001",
  14468=>"111000101",
  14469=>"000001111",
  14470=>"100101100",
  14471=>"101011111",
  14472=>"000000011",
  14473=>"011101110",
  14474=>"011001100",
  14475=>"010010011",
  14476=>"110011000",
  14477=>"000011111",
  14478=>"111000001",
  14479=>"010010001",
  14480=>"000011100",
  14481=>"000010110",
  14482=>"101000110",
  14483=>"110101011",
  14484=>"101101001",
  14485=>"011011100",
  14486=>"011011100",
  14487=>"001111010",
  14488=>"010100001",
  14489=>"000001010",
  14490=>"011011011",
  14491=>"101110010",
  14492=>"000010001",
  14493=>"111110101",
  14494=>"101000101",
  14495=>"000011000",
  14496=>"001111101",
  14497=>"111111000",
  14498=>"010110001",
  14499=>"011011010",
  14500=>"100000001",
  14501=>"011001000",
  14502=>"101010100",
  14503=>"111000010",
  14504=>"101101101",
  14505=>"011100001",
  14506=>"001000010",
  14507=>"010100001",
  14508=>"000011100",
  14509=>"000111000",
  14510=>"001000010",
  14511=>"000110111",
  14512=>"110111001",
  14513=>"111101101",
  14514=>"110010010",
  14515=>"001000101",
  14516=>"000001100",
  14517=>"000100111",
  14518=>"000011000",
  14519=>"000001011",
  14520=>"010101110",
  14521=>"111011001",
  14522=>"100010101",
  14523=>"011000011",
  14524=>"100101101",
  14525=>"100111100",
  14526=>"110100100",
  14527=>"011110011",
  14528=>"001101001",
  14529=>"101101001",
  14530=>"010100011",
  14531=>"111111010",
  14532=>"001110110",
  14533=>"000000010",
  14534=>"100101011",
  14535=>"111010111",
  14536=>"101011001",
  14537=>"101100110",
  14538=>"111101111",
  14539=>"110010110",
  14540=>"100010010",
  14541=>"111100101",
  14542=>"010000011",
  14543=>"110100010",
  14544=>"011100011",
  14545=>"110100000",
  14546=>"000001001",
  14547=>"100111100",
  14548=>"111001011",
  14549=>"101000001",
  14550=>"010111111",
  14551=>"011010010",
  14552=>"100010011",
  14553=>"100100101",
  14554=>"100110111",
  14555=>"110111101",
  14556=>"011101111",
  14557=>"111100101",
  14558=>"110100101",
  14559=>"110010110",
  14560=>"110011001",
  14561=>"011001111",
  14562=>"010101011",
  14563=>"111101111",
  14564=>"011001000",
  14565=>"010100101",
  14566=>"111111011",
  14567=>"101000111",
  14568=>"010001110",
  14569=>"111100001",
  14570=>"001111000",
  14571=>"111010000",
  14572=>"000101010",
  14573=>"000011101",
  14574=>"111101011",
  14575=>"010100101",
  14576=>"000001110",
  14577=>"000001000",
  14578=>"100001101",
  14579=>"010010101",
  14580=>"100101111",
  14581=>"111101000",
  14582=>"011010000",
  14583=>"000110010",
  14584=>"011101101",
  14585=>"000000110",
  14586=>"011001011",
  14587=>"000001000",
  14588=>"111010101",
  14589=>"000000101",
  14590=>"111111001",
  14591=>"001001101",
  14592=>"001100001",
  14593=>"100001101",
  14594=>"010110101",
  14595=>"001101011",
  14596=>"100101001",
  14597=>"011000001",
  14598=>"001010100",
  14599=>"100010100",
  14600=>"011101101",
  14601=>"110100101",
  14602=>"101111001",
  14603=>"110000110",
  14604=>"011000001",
  14605=>"110010111",
  14606=>"010000000",
  14607=>"111100110",
  14608=>"000100001",
  14609=>"010000010",
  14610=>"111100011",
  14611=>"011010110",
  14612=>"111101001",
  14613=>"010101010",
  14614=>"000101000",
  14615=>"011111011",
  14616=>"111001011",
  14617=>"000010000",
  14618=>"101011100",
  14619=>"101010001",
  14620=>"001101001",
  14621=>"101000101",
  14622=>"000010000",
  14623=>"100001000",
  14624=>"000101111",
  14625=>"001010001",
  14626=>"101010001",
  14627=>"001001101",
  14628=>"000000000",
  14629=>"000100100",
  14630=>"110101100",
  14631=>"011100000",
  14632=>"110111111",
  14633=>"000100010",
  14634=>"100010111",
  14635=>"010001100",
  14636=>"000000110",
  14637=>"010111000",
  14638=>"101000001",
  14639=>"111101110",
  14640=>"000010110",
  14641=>"010001001",
  14642=>"000010110",
  14643=>"111010001",
  14644=>"110101011",
  14645=>"000010101",
  14646=>"110001111",
  14647=>"111111101",
  14648=>"000011011",
  14649=>"101101000",
  14650=>"001101110",
  14651=>"110000100",
  14652=>"101100110",
  14653=>"010111111",
  14654=>"000010100",
  14655=>"101011110",
  14656=>"101001010",
  14657=>"000010110",
  14658=>"110101111",
  14659=>"100100101",
  14660=>"011101100",
  14661=>"000110000",
  14662=>"111000001",
  14663=>"110011001",
  14664=>"010111000",
  14665=>"001100101",
  14666=>"000110010",
  14667=>"101110000",
  14668=>"100001001",
  14669=>"000100000",
  14670=>"110101011",
  14671=>"100100101",
  14672=>"100111111",
  14673=>"000011101",
  14674=>"011100010",
  14675=>"011001100",
  14676=>"110110111",
  14677=>"000010010",
  14678=>"110101111",
  14679=>"001110110",
  14680=>"011000111",
  14681=>"110001001",
  14682=>"010101010",
  14683=>"110001001",
  14684=>"010110101",
  14685=>"000010010",
  14686=>"010010000",
  14687=>"001001111",
  14688=>"110101001",
  14689=>"010010101",
  14690=>"111010110",
  14691=>"100000000",
  14692=>"001001010",
  14693=>"011010011",
  14694=>"011100010",
  14695=>"011101100",
  14696=>"000111000",
  14697=>"110100110",
  14698=>"101001100",
  14699=>"111101011",
  14700=>"001100000",
  14701=>"111011010",
  14702=>"101110000",
  14703=>"000111100",
  14704=>"000100001",
  14705=>"000000100",
  14706=>"000011100",
  14707=>"100110000",
  14708=>"010110101",
  14709=>"110111001",
  14710=>"011110001",
  14711=>"000010110",
  14712=>"000111000",
  14713=>"011101110",
  14714=>"111110000",
  14715=>"010010110",
  14716=>"000010000",
  14717=>"111011010",
  14718=>"110110101",
  14719=>"000111000",
  14720=>"101100110",
  14721=>"011101000",
  14722=>"001110101",
  14723=>"001010101",
  14724=>"001010001",
  14725=>"000000111",
  14726=>"111100010",
  14727=>"100111010",
  14728=>"110111111",
  14729=>"001100111",
  14730=>"110011100",
  14731=>"011111100",
  14732=>"001100000",
  14733=>"111011010",
  14734=>"000010101",
  14735=>"101011110",
  14736=>"000011001",
  14737=>"101100111",
  14738=>"110001000",
  14739=>"001001011",
  14740=>"010100001",
  14741=>"001011111",
  14742=>"010011011",
  14743=>"101100000",
  14744=>"111010101",
  14745=>"010010000",
  14746=>"100110101",
  14747=>"000011111",
  14748=>"010100111",
  14749=>"000001000",
  14750=>"010101010",
  14751=>"000100010",
  14752=>"010010110",
  14753=>"000001100",
  14754=>"000101001",
  14755=>"000000110",
  14756=>"000000111",
  14757=>"011101001",
  14758=>"111111011",
  14759=>"011010001",
  14760=>"010000110",
  14761=>"010001010",
  14762=>"010001110",
  14763=>"101110110",
  14764=>"111011011",
  14765=>"101111110",
  14766=>"011111000",
  14767=>"100101101",
  14768=>"111101010",
  14769=>"001010101",
  14770=>"111101100",
  14771=>"100111001",
  14772=>"101111110",
  14773=>"110110101",
  14774=>"101110101",
  14775=>"001010110",
  14776=>"001001111",
  14777=>"111101110",
  14778=>"111111101",
  14779=>"011001110",
  14780=>"000110000",
  14781=>"000101011",
  14782=>"101110110",
  14783=>"001100110",
  14784=>"000101101",
  14785=>"100001110",
  14786=>"000110111",
  14787=>"111111000",
  14788=>"100101111",
  14789=>"101100101",
  14790=>"000100000",
  14791=>"011011000",
  14792=>"101011111",
  14793=>"000111000",
  14794=>"011010110",
  14795=>"100100000",
  14796=>"000010100",
  14797=>"111100110",
  14798=>"101000000",
  14799=>"011010001",
  14800=>"100011111",
  14801=>"100101101",
  14802=>"111010101",
  14803=>"110110111",
  14804=>"101001110",
  14805=>"011101000",
  14806=>"100001110",
  14807=>"110100000",
  14808=>"100101000",
  14809=>"111100010",
  14810=>"010101101",
  14811=>"010101010",
  14812=>"001000011",
  14813=>"001101100",
  14814=>"110100000",
  14815=>"100000100",
  14816=>"111010011",
  14817=>"101001010",
  14818=>"010010000",
  14819=>"010101010",
  14820=>"001010010",
  14821=>"100110000",
  14822=>"110000111",
  14823=>"010100110",
  14824=>"010111110",
  14825=>"011110110",
  14826=>"000110001",
  14827=>"100000111",
  14828=>"110100010",
  14829=>"110111010",
  14830=>"001111001",
  14831=>"011100000",
  14832=>"110101000",
  14833=>"100101000",
  14834=>"001110001",
  14835=>"111010011",
  14836=>"011100101",
  14837=>"001000000",
  14838=>"111111000",
  14839=>"010001010",
  14840=>"011110001",
  14841=>"110110111",
  14842=>"010000110",
  14843=>"001100000",
  14844=>"011110111",
  14845=>"101111000",
  14846=>"010000110",
  14847=>"000000001",
  14848=>"101101000",
  14849=>"000001100",
  14850=>"100011111",
  14851=>"100100011",
  14852=>"111011001",
  14853=>"000000101",
  14854=>"001100010",
  14855=>"000001101",
  14856=>"001010100",
  14857=>"011001010",
  14858=>"000110011",
  14859=>"110101111",
  14860=>"001011111",
  14861=>"101111100",
  14862=>"000001111",
  14863=>"101111010",
  14864=>"010100101",
  14865=>"011010000",
  14866=>"000001111",
  14867=>"101000000",
  14868=>"100110100",
  14869=>"011101100",
  14870=>"100111110",
  14871=>"101000100",
  14872=>"000000110",
  14873=>"100000000",
  14874=>"010010001",
  14875=>"010100000",
  14876=>"000000010",
  14877=>"100001010",
  14878=>"110100100",
  14879=>"001100111",
  14880=>"100100000",
  14881=>"110000001",
  14882=>"111000111",
  14883=>"100110110",
  14884=>"010110100",
  14885=>"101010010",
  14886=>"111010000",
  14887=>"101001110",
  14888=>"100000110",
  14889=>"000011000",
  14890=>"111110010",
  14891=>"110101000",
  14892=>"000100100",
  14893=>"111000010",
  14894=>"011100100",
  14895=>"101111110",
  14896=>"011100000",
  14897=>"110110101",
  14898=>"100111011",
  14899=>"010000111",
  14900=>"001011110",
  14901=>"100101101",
  14902=>"101100110",
  14903=>"000110101",
  14904=>"011011101",
  14905=>"000101010",
  14906=>"111110101",
  14907=>"010001000",
  14908=>"011000000",
  14909=>"000111111",
  14910=>"101101110",
  14911=>"110100110",
  14912=>"111101000",
  14913=>"011110111",
  14914=>"101111010",
  14915=>"011101000",
  14916=>"001010010",
  14917=>"011100100",
  14918=>"100111110",
  14919=>"011110111",
  14920=>"010000001",
  14921=>"101110010",
  14922=>"001111010",
  14923=>"000011110",
  14924=>"001111111",
  14925=>"000001111",
  14926=>"101001000",
  14927=>"000001000",
  14928=>"001101111",
  14929=>"001111000",
  14930=>"000101010",
  14931=>"011101011",
  14932=>"000001101",
  14933=>"111101000",
  14934=>"000110000",
  14935=>"011010001",
  14936=>"011111111",
  14937=>"010000110",
  14938=>"101101111",
  14939=>"111010101",
  14940=>"010000010",
  14941=>"110000101",
  14942=>"011110011",
  14943=>"111100011",
  14944=>"000000101",
  14945=>"100010101",
  14946=>"111111011",
  14947=>"111011101",
  14948=>"110000111",
  14949=>"001000100",
  14950=>"101000011",
  14951=>"100101101",
  14952=>"101101000",
  14953=>"100011101",
  14954=>"010100000",
  14955=>"011011110",
  14956=>"101001101",
  14957=>"010001011",
  14958=>"111100010",
  14959=>"011000010",
  14960=>"100110010",
  14961=>"110000001",
  14962=>"111100111",
  14963=>"111011000",
  14964=>"111111011",
  14965=>"010000100",
  14966=>"010010011",
  14967=>"000111010",
  14968=>"010001000",
  14969=>"000000010",
  14970=>"100110000",
  14971=>"011011110",
  14972=>"001111110",
  14973=>"001011111",
  14974=>"111111101",
  14975=>"101110001",
  14976=>"000001011",
  14977=>"011100100",
  14978=>"101111000",
  14979=>"011001111",
  14980=>"110101000",
  14981=>"000110000",
  14982=>"111001101",
  14983=>"100000000",
  14984=>"010001100",
  14985=>"001100001",
  14986=>"111100110",
  14987=>"101011100",
  14988=>"000001010",
  14989=>"001000011",
  14990=>"000101010",
  14991=>"000110001",
  14992=>"011001001",
  14993=>"111011100",
  14994=>"011010011",
  14995=>"000001111",
  14996=>"111000101",
  14997=>"100101101",
  14998=>"111101010",
  14999=>"100010000",
  15000=>"101111110",
  15001=>"110010101",
  15002=>"111001011",
  15003=>"101110101",
  15004=>"101110000",
  15005=>"100011110",
  15006=>"001011110",
  15007=>"101111111",
  15008=>"000010110",
  15009=>"001000001",
  15010=>"101001111",
  15011=>"111111110",
  15012=>"100011001",
  15013=>"001000100",
  15014=>"010111000",
  15015=>"111110101",
  15016=>"100110110",
  15017=>"000101100",
  15018=>"010110100",
  15019=>"100100111",
  15020=>"111111001",
  15021=>"110111000",
  15022=>"110010001",
  15023=>"000000100",
  15024=>"011100010",
  15025=>"000111110",
  15026=>"001111110",
  15027=>"101000100",
  15028=>"111010101",
  15029=>"111010100",
  15030=>"101010101",
  15031=>"100001000",
  15032=>"010010011",
  15033=>"101101101",
  15034=>"000100000",
  15035=>"100001110",
  15036=>"111000001",
  15037=>"000000001",
  15038=>"100101100",
  15039=>"100000111",
  15040=>"011101100",
  15041=>"010000001",
  15042=>"101111011",
  15043=>"011100101",
  15044=>"100110011",
  15045=>"011001101",
  15046=>"001000111",
  15047=>"000110011",
  15048=>"010100010",
  15049=>"001010100",
  15050=>"101101101",
  15051=>"111111001",
  15052=>"011101101",
  15053=>"110110111",
  15054=>"010111100",
  15055=>"111111001",
  15056=>"001011010",
  15057=>"000001000",
  15058=>"011110011",
  15059=>"100100000",
  15060=>"000010001",
  15061=>"000110000",
  15062=>"000000001",
  15063=>"101100010",
  15064=>"110001110",
  15065=>"110101100",
  15066=>"010100001",
  15067=>"100100110",
  15068=>"000000000",
  15069=>"011000010",
  15070=>"110000101",
  15071=>"101011001",
  15072=>"101001011",
  15073=>"000110101",
  15074=>"010000010",
  15075=>"000010011",
  15076=>"001011110",
  15077=>"010011010",
  15078=>"111110100",
  15079=>"111000100",
  15080=>"001001000",
  15081=>"010011001",
  15082=>"100111101",
  15083=>"110011011",
  15084=>"101101111",
  15085=>"100011011",
  15086=>"001000001",
  15087=>"000011100",
  15088=>"111000100",
  15089=>"101011011",
  15090=>"010000110",
  15091=>"101110100",
  15092=>"111111111",
  15093=>"001011111",
  15094=>"110000100",
  15095=>"100000101",
  15096=>"011001011",
  15097=>"100000011",
  15098=>"101111010",
  15099=>"000000001",
  15100=>"010101001",
  15101=>"000110010",
  15102=>"110000111",
  15103=>"100011111",
  15104=>"101010000",
  15105=>"011111110",
  15106=>"011010011",
  15107=>"110111110",
  15108=>"100011000",
  15109=>"100000111",
  15110=>"010110011",
  15111=>"101101001",
  15112=>"100000001",
  15113=>"000001111",
  15114=>"111100010",
  15115=>"010111100",
  15116=>"100011010",
  15117=>"001100100",
  15118=>"110010111",
  15119=>"101101011",
  15120=>"010000000",
  15121=>"010111110",
  15122=>"001100110",
  15123=>"011000101",
  15124=>"011111110",
  15125=>"110011011",
  15126=>"111111001",
  15127=>"110011111",
  15128=>"010100011",
  15129=>"111111000",
  15130=>"001011010",
  15131=>"000111011",
  15132=>"110011001",
  15133=>"000110010",
  15134=>"100001001",
  15135=>"110101010",
  15136=>"011110111",
  15137=>"010110011",
  15138=>"001110101",
  15139=>"111101110",
  15140=>"110100111",
  15141=>"000101001",
  15142=>"110111111",
  15143=>"111010101",
  15144=>"110101011",
  15145=>"100000111",
  15146=>"100101000",
  15147=>"110000010",
  15148=>"111100001",
  15149=>"011101001",
  15150=>"100001000",
  15151=>"110111010",
  15152=>"010110011",
  15153=>"111110110",
  15154=>"111101111",
  15155=>"111010111",
  15156=>"110010001",
  15157=>"101001001",
  15158=>"100101011",
  15159=>"000000010",
  15160=>"101101111",
  15161=>"110101110",
  15162=>"111100000",
  15163=>"010110001",
  15164=>"011110001",
  15165=>"100100110",
  15166=>"100000011",
  15167=>"110011011",
  15168=>"000011011",
  15169=>"000101011",
  15170=>"001101101",
  15171=>"100010100",
  15172=>"100011010",
  15173=>"011000100",
  15174=>"010110000",
  15175=>"100010110",
  15176=>"000110110",
  15177=>"111110110",
  15178=>"101101101",
  15179=>"001000101",
  15180=>"110001100",
  15181=>"111001111",
  15182=>"110010001",
  15183=>"011111011",
  15184=>"000100111",
  15185=>"100001111",
  15186=>"011100100",
  15187=>"110000010",
  15188=>"001111001",
  15189=>"001101101",
  15190=>"011000010",
  15191=>"000011111",
  15192=>"010000100",
  15193=>"010110110",
  15194=>"001101101",
  15195=>"000110101",
  15196=>"010001001",
  15197=>"011101110",
  15198=>"001011010",
  15199=>"110010000",
  15200=>"011111011",
  15201=>"000010011",
  15202=>"001000100",
  15203=>"011110010",
  15204=>"101100011",
  15205=>"001000110",
  15206=>"010101011",
  15207=>"100100111",
  15208=>"101100011",
  15209=>"111100000",
  15210=>"010000000",
  15211=>"111100110",
  15212=>"100011111",
  15213=>"110001000",
  15214=>"000100101",
  15215=>"111001010",
  15216=>"111101110",
  15217=>"110100000",
  15218=>"011101010",
  15219=>"111100101",
  15220=>"110100001",
  15221=>"001111001",
  15222=>"110100001",
  15223=>"011111000",
  15224=>"101001000",
  15225=>"111100100",
  15226=>"000110111",
  15227=>"111110111",
  15228=>"000110000",
  15229=>"011101110",
  15230=>"111001100",
  15231=>"010110100",
  15232=>"111011111",
  15233=>"001010011",
  15234=>"111100111",
  15235=>"010111011",
  15236=>"000100110",
  15237=>"100010000",
  15238=>"001011100",
  15239=>"100110101",
  15240=>"010011001",
  15241=>"100111100",
  15242=>"010111100",
  15243=>"010000001",
  15244=>"011111001",
  15245=>"111101001",
  15246=>"101001011",
  15247=>"100000001",
  15248=>"101101000",
  15249=>"100100101",
  15250=>"010000100",
  15251=>"110111100",
  15252=>"000100000",
  15253=>"111000111",
  15254=>"111100101",
  15255=>"111101101",
  15256=>"001101000",
  15257=>"000111000",
  15258=>"101101011",
  15259=>"110101111",
  15260=>"111010000",
  15261=>"010101001",
  15262=>"101101101",
  15263=>"000111111",
  15264=>"100001000",
  15265=>"111000001",
  15266=>"111001100",
  15267=>"111111111",
  15268=>"101010111",
  15269=>"101011001",
  15270=>"001100010",
  15271=>"010100111",
  15272=>"011001011",
  15273=>"010011111",
  15274=>"011110010",
  15275=>"111000001",
  15276=>"011100101",
  15277=>"000010010",
  15278=>"110101000",
  15279=>"110110100",
  15280=>"001110000",
  15281=>"001001011",
  15282=>"000010111",
  15283=>"010111111",
  15284=>"100110101",
  15285=>"000010110",
  15286=>"100001101",
  15287=>"110001101",
  15288=>"001100011",
  15289=>"110111000",
  15290=>"001110001",
  15291=>"010100110",
  15292=>"101001000",
  15293=>"111101101",
  15294=>"101111000",
  15295=>"110110111",
  15296=>"011101000",
  15297=>"011100110",
  15298=>"100100101",
  15299=>"011110010",
  15300=>"011110000",
  15301=>"001111010",
  15302=>"010000100",
  15303=>"011101111",
  15304=>"001011001",
  15305=>"100001110",
  15306=>"111011110",
  15307=>"101001000",
  15308=>"000110010",
  15309=>"111101001",
  15310=>"001011011",
  15311=>"011111110",
  15312=>"101100000",
  15313=>"011001010",
  15314=>"010001011",
  15315=>"110100011",
  15316=>"100101011",
  15317=>"000011001",
  15318=>"001100000",
  15319=>"110101001",
  15320=>"011110000",
  15321=>"010011110",
  15322=>"111111111",
  15323=>"001011110",
  15324=>"010011110",
  15325=>"111111000",
  15326=>"111100100",
  15327=>"001000110",
  15328=>"010101101",
  15329=>"011001011",
  15330=>"111110001",
  15331=>"100010001",
  15332=>"000111110",
  15333=>"001111000",
  15334=>"111010111",
  15335=>"000001000",
  15336=>"000000000",
  15337=>"101001010",
  15338=>"011011110",
  15339=>"000000101",
  15340=>"011001110",
  15341=>"011000010",
  15342=>"001011100",
  15343=>"010011101",
  15344=>"010000010",
  15345=>"101100111",
  15346=>"110101001",
  15347=>"101111001",
  15348=>"111100101",
  15349=>"000110100",
  15350=>"111101000",
  15351=>"001000111",
  15352=>"101100101",
  15353=>"101001011",
  15354=>"001110011",
  15355=>"110000010",
  15356=>"111110110",
  15357=>"110000011",
  15358=>"110101110",
  15359=>"000101111",
  15360=>"111100011",
  15361=>"000000011",
  15362=>"010011011",
  15363=>"000000000",
  15364=>"000111010",
  15365=>"111111001",
  15366=>"100101011",
  15367=>"000100100",
  15368=>"010000001",
  15369=>"100001110",
  15370=>"001010101",
  15371=>"110101110",
  15372=>"010111001",
  15373=>"101101110",
  15374=>"000100101",
  15375=>"111010010",
  15376=>"010110001",
  15377=>"100001101",
  15378=>"000101101",
  15379=>"011010101",
  15380=>"011111010",
  15381=>"001101010",
  15382=>"110101001",
  15383=>"111101110",
  15384=>"100000101",
  15385=>"101110011",
  15386=>"100010000",
  15387=>"111011010",
  15388=>"100000110",
  15389=>"011110001",
  15390=>"001001000",
  15391=>"101000000",
  15392=>"100100100",
  15393=>"100001010",
  15394=>"110011010",
  15395=>"010100111",
  15396=>"101100011",
  15397=>"110011110",
  15398=>"110101001",
  15399=>"110001001",
  15400=>"010011101",
  15401=>"110111110",
  15402=>"110001011",
  15403=>"111100100",
  15404=>"110000100",
  15405=>"001001101",
  15406=>"010010110",
  15407=>"000000110",
  15408=>"100011101",
  15409=>"000010101",
  15410=>"110101000",
  15411=>"011010000",
  15412=>"011000010",
  15413=>"100010010",
  15414=>"000000010",
  15415=>"101111111",
  15416=>"110001111",
  15417=>"101101010",
  15418=>"110000000",
  15419=>"110110111",
  15420=>"000000000",
  15421=>"110110100",
  15422=>"000111100",
  15423=>"111000100",
  15424=>"101000101",
  15425=>"000100000",
  15426=>"010110001",
  15427=>"010010101",
  15428=>"010000001",
  15429=>"101101000",
  15430=>"101001110",
  15431=>"110111100",
  15432=>"100100001",
  15433=>"011101110",
  15434=>"010001011",
  15435=>"111000001",
  15436=>"100111101",
  15437=>"011110101",
  15438=>"111000111",
  15439=>"101101110",
  15440=>"001000000",
  15441=>"111110001",
  15442=>"111010000",
  15443=>"100001111",
  15444=>"001011100",
  15445=>"101001000",
  15446=>"011011010",
  15447=>"100001110",
  15448=>"101000000",
  15449=>"111100011",
  15450=>"011110011",
  15451=>"010111110",
  15452=>"111110001",
  15453=>"111001011",
  15454=>"110110111",
  15455=>"000110010",
  15456=>"000110001",
  15457=>"010100010",
  15458=>"001111111",
  15459=>"000110010",
  15460=>"000000000",
  15461=>"101111111",
  15462=>"011010000",
  15463=>"110000000",
  15464=>"011110111",
  15465=>"000000010",
  15466=>"101000001",
  15467=>"010101001",
  15468=>"110000101",
  15469=>"100100001",
  15470=>"101000101",
  15471=>"001011001",
  15472=>"001100101",
  15473=>"101001001",
  15474=>"111111110",
  15475=>"001101100",
  15476=>"010101000",
  15477=>"100000011",
  15478=>"101011100",
  15479=>"001110101",
  15480=>"001010100",
  15481=>"110101110",
  15482=>"101110111",
  15483=>"011101010",
  15484=>"101101010",
  15485=>"111000001",
  15486=>"010110110",
  15487=>"011100000",
  15488=>"000001010",
  15489=>"010101011",
  15490=>"010101111",
  15491=>"100101000",
  15492=>"000010000",
  15493=>"011001000",
  15494=>"101111110",
  15495=>"111010010",
  15496=>"111101101",
  15497=>"110110100",
  15498=>"111100110",
  15499=>"111001101",
  15500=>"001001110",
  15501=>"100110111",
  15502=>"101101100",
  15503=>"011010000",
  15504=>"011010110",
  15505=>"000100100",
  15506=>"110010111",
  15507=>"100100100",
  15508=>"011000111",
  15509=>"111111010",
  15510=>"000000101",
  15511=>"100101111",
  15512=>"101000000",
  15513=>"001010000",
  15514=>"111111000",
  15515=>"011010100",
  15516=>"110101000",
  15517=>"000100000",
  15518=>"001011011",
  15519=>"010100010",
  15520=>"111001111",
  15521=>"101011110",
  15522=>"111001000",
  15523=>"001000101",
  15524=>"110110001",
  15525=>"111010001",
  15526=>"101100010",
  15527=>"110010010",
  15528=>"111110000",
  15529=>"010000111",
  15530=>"000000101",
  15531=>"011011001",
  15532=>"001010011",
  15533=>"001000110",
  15534=>"010110001",
  15535=>"001101100",
  15536=>"011000101",
  15537=>"011000110",
  15538=>"100011100",
  15539=>"111100100",
  15540=>"001101101",
  15541=>"110111011",
  15542=>"110000000",
  15543=>"100000100",
  15544=>"010100000",
  15545=>"000101101",
  15546=>"110110111",
  15547=>"001011001",
  15548=>"001100100",
  15549=>"110000001",
  15550=>"001000111",
  15551=>"111100011",
  15552=>"001100001",
  15553=>"001011001",
  15554=>"111101101",
  15555=>"011000000",
  15556=>"110001111",
  15557=>"010101011",
  15558=>"110110011",
  15559=>"111101010",
  15560=>"100011001",
  15561=>"011100010",
  15562=>"001110101",
  15563=>"000000100",
  15564=>"010010110",
  15565=>"111101110",
  15566=>"111010000",
  15567=>"111101110",
  15568=>"001110011",
  15569=>"111110101",
  15570=>"110101101",
  15571=>"000011101",
  15572=>"010100001",
  15573=>"011010011",
  15574=>"001000111",
  15575=>"000111000",
  15576=>"010000000",
  15577=>"111011000",
  15578=>"011111011",
  15579=>"001011111",
  15580=>"011011111",
  15581=>"111010111",
  15582=>"110001101",
  15583=>"010100100",
  15584=>"111111111",
  15585=>"101001111",
  15586=>"001011000",
  15587=>"100100001",
  15588=>"110011111",
  15589=>"111011001",
  15590=>"100111010",
  15591=>"001010010",
  15592=>"010000100",
  15593=>"000101101",
  15594=>"010111011",
  15595=>"101011111",
  15596=>"101111000",
  15597=>"001011111",
  15598=>"011010011",
  15599=>"110111110",
  15600=>"111010000",
  15601=>"001101100",
  15602=>"110000110",
  15603=>"110111101",
  15604=>"000100101",
  15605=>"010111000",
  15606=>"001111111",
  15607=>"100110111",
  15608=>"111001101",
  15609=>"101101101",
  15610=>"100011100",
  15611=>"011111111",
  15612=>"000001100",
  15613=>"110111110",
  15614=>"110110101",
  15615=>"010001010",
  15616=>"100100011",
  15617=>"010100011",
  15618=>"011111100",
  15619=>"101101000",
  15620=>"000111011",
  15621=>"011110100",
  15622=>"100101100",
  15623=>"000101100",
  15624=>"010001101",
  15625=>"000010111",
  15626=>"001110111",
  15627=>"100111111",
  15628=>"100010110",
  15629=>"011100010",
  15630=>"000011010",
  15631=>"011100010",
  15632=>"000001001",
  15633=>"010001101",
  15634=>"100100100",
  15635=>"000011010",
  15636=>"000101011",
  15637=>"010100000",
  15638=>"001111011",
  15639=>"110010111",
  15640=>"101001111",
  15641=>"010100001",
  15642=>"001100000",
  15643=>"111001001",
  15644=>"111111110",
  15645=>"000110110",
  15646=>"011011001",
  15647=>"101100110",
  15648=>"100111110",
  15649=>"001111010",
  15650=>"110011011",
  15651=>"100001110",
  15652=>"001100101",
  15653=>"110100111",
  15654=>"000001011",
  15655=>"000111010",
  15656=>"100111001",
  15657=>"000111010",
  15658=>"101110001",
  15659=>"110000000",
  15660=>"000111100",
  15661=>"110110000",
  15662=>"000000100",
  15663=>"110011000",
  15664=>"100010101",
  15665=>"111000100",
  15666=>"110111010",
  15667=>"101101011",
  15668=>"011110100",
  15669=>"111001000",
  15670=>"000010101",
  15671=>"110011001",
  15672=>"001101111",
  15673=>"110000000",
  15674=>"101000011",
  15675=>"000010101",
  15676=>"111011010",
  15677=>"111100010",
  15678=>"000010111",
  15679=>"100011001",
  15680=>"001011010",
  15681=>"011101100",
  15682=>"110110111",
  15683=>"101010100",
  15684=>"001001010",
  15685=>"010010101",
  15686=>"001110101",
  15687=>"101110111",
  15688=>"010010111",
  15689=>"010110111",
  15690=>"110110101",
  15691=>"111011100",
  15692=>"100001100",
  15693=>"110010100",
  15694=>"111000100",
  15695=>"111011001",
  15696=>"000101111",
  15697=>"001111000",
  15698=>"101100101",
  15699=>"110111100",
  15700=>"101000000",
  15701=>"000111111",
  15702=>"011010010",
  15703=>"111101110",
  15704=>"100110010",
  15705=>"111011001",
  15706=>"100101000",
  15707=>"001010011",
  15708=>"101111001",
  15709=>"100001000",
  15710=>"000010010",
  15711=>"010000000",
  15712=>"111000110",
  15713=>"100111110",
  15714=>"100110111",
  15715=>"101110111",
  15716=>"001101010",
  15717=>"101000001",
  15718=>"011101000",
  15719=>"110101001",
  15720=>"000111000",
  15721=>"001111111",
  15722=>"011111000",
  15723=>"100111101",
  15724=>"101100001",
  15725=>"101011000",
  15726=>"100001110",
  15727=>"011101100",
  15728=>"101011000",
  15729=>"100111011",
  15730=>"000011000",
  15731=>"100010110",
  15732=>"111111011",
  15733=>"110010101",
  15734=>"100100111",
  15735=>"101011110",
  15736=>"010101001",
  15737=>"110001001",
  15738=>"100111011",
  15739=>"000111110",
  15740=>"101010011",
  15741=>"101111001",
  15742=>"100111101",
  15743=>"110011110",
  15744=>"100101110",
  15745=>"000100011",
  15746=>"000110011",
  15747=>"101101011",
  15748=>"111100110",
  15749=>"111111111",
  15750=>"111100100",
  15751=>"101101011",
  15752=>"101101011",
  15753=>"011010101",
  15754=>"101010010",
  15755=>"111110100",
  15756=>"110000101",
  15757=>"100000000",
  15758=>"101101110",
  15759=>"100010000",
  15760=>"010000000",
  15761=>"000111011",
  15762=>"101110010",
  15763=>"000011011",
  15764=>"011100110",
  15765=>"011001101",
  15766=>"001001011",
  15767=>"000010100",
  15768=>"110101000",
  15769=>"111111110",
  15770=>"101001110",
  15771=>"011111100",
  15772=>"111110111",
  15773=>"001000100",
  15774=>"111001110",
  15775=>"111100000",
  15776=>"011110100",
  15777=>"010000100",
  15778=>"110001110",
  15779=>"010010110",
  15780=>"011010101",
  15781=>"100010010",
  15782=>"011011001",
  15783=>"000100010",
  15784=>"001001110",
  15785=>"000000010",
  15786=>"110011011",
  15787=>"100001110",
  15788=>"110010111",
  15789=>"110110111",
  15790=>"001111000",
  15791=>"001010011",
  15792=>"101011100",
  15793=>"000010110",
  15794=>"010011000",
  15795=>"101101111",
  15796=>"110011111",
  15797=>"110101011",
  15798=>"111101011",
  15799=>"010111001",
  15800=>"011101111",
  15801=>"101101111",
  15802=>"111110111",
  15803=>"111000111",
  15804=>"111101111",
  15805=>"111000010",
  15806=>"111011011",
  15807=>"011000111",
  15808=>"011000001",
  15809=>"111101101",
  15810=>"000010010",
  15811=>"001011111",
  15812=>"011110110",
  15813=>"001101011",
  15814=>"101001001",
  15815=>"000101001",
  15816=>"111100001",
  15817=>"001011100",
  15818=>"101111110",
  15819=>"010000010",
  15820=>"101011111",
  15821=>"001110001",
  15822=>"000000110",
  15823=>"100111000",
  15824=>"100010000",
  15825=>"011111101",
  15826=>"111001111",
  15827=>"001110101",
  15828=>"100001100",
  15829=>"100100010",
  15830=>"010010010",
  15831=>"000001010",
  15832=>"110010100",
  15833=>"011100000",
  15834=>"101110001",
  15835=>"111100111",
  15836=>"000011011",
  15837=>"100110101",
  15838=>"100110011",
  15839=>"110111100",
  15840=>"111101101",
  15841=>"010010100",
  15842=>"011110000",
  15843=>"101101111",
  15844=>"010000111",
  15845=>"110110111",
  15846=>"010100110",
  15847=>"010100111",
  15848=>"100111110",
  15849=>"011110111",
  15850=>"011001110",
  15851=>"111001001",
  15852=>"010101011",
  15853=>"111110100",
  15854=>"111101101",
  15855=>"001101011",
  15856=>"101000111",
  15857=>"100011010",
  15858=>"111000010",
  15859=>"000011101",
  15860=>"111111111",
  15861=>"101110000",
  15862=>"010110110",
  15863=>"010000100",
  15864=>"101000101",
  15865=>"110001010",
  15866=>"110001110",
  15867=>"110100110",
  15868=>"101110110",
  15869=>"100011000",
  15870=>"010110101",
  15871=>"000100101",
  15872=>"110010001",
  15873=>"011101100",
  15874=>"011101100",
  15875=>"010001111",
  15876=>"100110100",
  15877=>"001101011",
  15878=>"000010110",
  15879=>"001000100",
  15880=>"010000000",
  15881=>"101010101",
  15882=>"101011100",
  15883=>"010010001",
  15884=>"100101101",
  15885=>"011100000",
  15886=>"000111101",
  15887=>"010001001",
  15888=>"101000001",
  15889=>"010011100",
  15890=>"011011001",
  15891=>"100100111",
  15892=>"100111101",
  15893=>"000111110",
  15894=>"100111111",
  15895=>"110001111",
  15896=>"000011011",
  15897=>"111111100",
  15898=>"011000111",
  15899=>"000101010",
  15900=>"010110001",
  15901=>"110001100",
  15902=>"010100001",
  15903=>"010110100",
  15904=>"100100101",
  15905=>"001101100",
  15906=>"011110011",
  15907=>"000001011",
  15908=>"100010010",
  15909=>"110110000",
  15910=>"001011001",
  15911=>"111111111",
  15912=>"010100000",
  15913=>"101111111",
  15914=>"001011111",
  15915=>"111000001",
  15916=>"000111010",
  15917=>"010110110",
  15918=>"100100001",
  15919=>"010000010",
  15920=>"010001111",
  15921=>"101010000",
  15922=>"101001000",
  15923=>"101101111",
  15924=>"001101111",
  15925=>"010001011",
  15926=>"100111011",
  15927=>"000111100",
  15928=>"100010111",
  15929=>"101011101",
  15930=>"010110011",
  15931=>"100111001",
  15932=>"000110010",
  15933=>"110011111",
  15934=>"110110000",
  15935=>"111101110",
  15936=>"010010100",
  15937=>"111011000",
  15938=>"101000110",
  15939=>"010111010",
  15940=>"010010001",
  15941=>"110011100",
  15942=>"001111111",
  15943=>"010110000",
  15944=>"110110111",
  15945=>"010110010",
  15946=>"100010010",
  15947=>"000111100",
  15948=>"011010000",
  15949=>"100101000",
  15950=>"100000001",
  15951=>"101100000",
  15952=>"000011110",
  15953=>"001101000",
  15954=>"010001011",
  15955=>"100010110",
  15956=>"001100100",
  15957=>"100011111",
  15958=>"011100100",
  15959=>"001011111",
  15960=>"100001011",
  15961=>"110101110",
  15962=>"011111010",
  15963=>"111110010",
  15964=>"100000010",
  15965=>"010000111",
  15966=>"111110010",
  15967=>"010010110",
  15968=>"000001111",
  15969=>"100111001",
  15970=>"110000010",
  15971=>"001000100",
  15972=>"011010101",
  15973=>"000001110",
  15974=>"111100111",
  15975=>"001011000",
  15976=>"000110011",
  15977=>"110000100",
  15978=>"100101011",
  15979=>"100110001",
  15980=>"111011011",
  15981=>"100100011",
  15982=>"100011011",
  15983=>"100011000",
  15984=>"001100111",
  15985=>"000110000",
  15986=>"100010100",
  15987=>"000001010",
  15988=>"111110011",
  15989=>"111110001",
  15990=>"011100001",
  15991=>"010001000",
  15992=>"000111110",
  15993=>"111100100",
  15994=>"101101111",
  15995=>"111010000",
  15996=>"100001010",
  15997=>"000100111",
  15998=>"011000001",
  15999=>"001001011",
  16000=>"010001110",
  16001=>"011101101",
  16002=>"101110011",
  16003=>"011111011",
  16004=>"001001011",
  16005=>"111001101",
  16006=>"100001001",
  16007=>"110110010",
  16008=>"000100010",
  16009=>"100101110",
  16010=>"010110101",
  16011=>"011011100",
  16012=>"110010011",
  16013=>"000100001",
  16014=>"100100111",
  16015=>"000110101",
  16016=>"010011010",
  16017=>"111011111",
  16018=>"001011101",
  16019=>"100000000",
  16020=>"111001110",
  16021=>"000010101",
  16022=>"010110011",
  16023=>"000001000",
  16024=>"111101101",
  16025=>"011001010",
  16026=>"011000011",
  16027=>"111001001",
  16028=>"001101001",
  16029=>"111001001",
  16030=>"000001100",
  16031=>"100000011",
  16032=>"100011101",
  16033=>"000110110",
  16034=>"111101000",
  16035=>"110000110",
  16036=>"110011010",
  16037=>"110001100",
  16038=>"100011000",
  16039=>"011100110",
  16040=>"101101010",
  16041=>"110111011",
  16042=>"011001100",
  16043=>"110011011",
  16044=>"110100001",
  16045=>"110011000",
  16046=>"011000111",
  16047=>"010110010",
  16048=>"000111001",
  16049=>"011011101",
  16050=>"110010101",
  16051=>"101101101",
  16052=>"001000100",
  16053=>"100001111",
  16054=>"110110001",
  16055=>"010001000",
  16056=>"101010100",
  16057=>"010011111",
  16058=>"011100011",
  16059=>"100100100",
  16060=>"110100010",
  16061=>"101101101",
  16062=>"111011010",
  16063=>"100110011",
  16064=>"110111111",
  16065=>"110000100",
  16066=>"101110010",
  16067=>"110010111",
  16068=>"111011001",
  16069=>"100100110",
  16070=>"100111101",
  16071=>"010100000",
  16072=>"011000010",
  16073=>"100001000",
  16074=>"000101100",
  16075=>"010101100",
  16076=>"110101011",
  16077=>"101111001",
  16078=>"011011111",
  16079=>"010101101",
  16080=>"010001100",
  16081=>"000000011",
  16082=>"100110111",
  16083=>"001011111",
  16084=>"001100101",
  16085=>"100100000",
  16086=>"011100011",
  16087=>"101010000",
  16088=>"111010001",
  16089=>"001011000",
  16090=>"001000000",
  16091=>"001011100",
  16092=>"001110111",
  16093=>"111101110",
  16094=>"010011111",
  16095=>"101001101",
  16096=>"100111110",
  16097=>"011111101",
  16098=>"101010001",
  16099=>"111110111",
  16100=>"001111101",
  16101=>"101111101",
  16102=>"101001011",
  16103=>"000011110",
  16104=>"101010110",
  16105=>"110001011",
  16106=>"111100000",
  16107=>"101010010",
  16108=>"001101111",
  16109=>"010011101",
  16110=>"111011100",
  16111=>"000011101",
  16112=>"110000101",
  16113=>"000100101",
  16114=>"011100001",
  16115=>"100001111",
  16116=>"010110000",
  16117=>"001110111",
  16118=>"101101110",
  16119=>"110111110",
  16120=>"001111010",
  16121=>"101110010",
  16122=>"010101011",
  16123=>"110100111",
  16124=>"100110000",
  16125=>"011100111",
  16126=>"110010010",
  16127=>"101011011",
  16128=>"000010010",
  16129=>"110000101",
  16130=>"010010001",
  16131=>"000011110",
  16132=>"111110101",
  16133=>"100000000",
  16134=>"110111100",
  16135=>"001111011",
  16136=>"011101010",
  16137=>"000000110",
  16138=>"010111101",
  16139=>"100011010",
  16140=>"110100010",
  16141=>"111110110",
  16142=>"000001000",
  16143=>"010001000",
  16144=>"111000001",
  16145=>"100111001",
  16146=>"111010001",
  16147=>"010001010",
  16148=>"111011100",
  16149=>"011101110",
  16150=>"110110100",
  16151=>"100100001",
  16152=>"111001111",
  16153=>"000001111",
  16154=>"110101100",
  16155=>"110010010",
  16156=>"000000011",
  16157=>"010110000",
  16158=>"010011111",
  16159=>"010101101",
  16160=>"011111011",
  16161=>"001100011",
  16162=>"000000100",
  16163=>"011000000",
  16164=>"111001110",
  16165=>"010111000",
  16166=>"000100011",
  16167=>"011111111",
  16168=>"111111011",
  16169=>"011010101",
  16170=>"100110110",
  16171=>"001110110",
  16172=>"010101000",
  16173=>"101001111",
  16174=>"001011001",
  16175=>"110000010",
  16176=>"101011100",
  16177=>"101000100",
  16178=>"001111111",
  16179=>"000000100",
  16180=>"101101000",
  16181=>"111000111",
  16182=>"111111110",
  16183=>"110111000",
  16184=>"111100100",
  16185=>"100110010",
  16186=>"110011110",
  16187=>"100110101",
  16188=>"100010110",
  16189=>"011001100",
  16190=>"000001100",
  16191=>"111001011",
  16192=>"010011000",
  16193=>"110001100",
  16194=>"000110101",
  16195=>"110010101",
  16196=>"110110001",
  16197=>"011000001",
  16198=>"110001111",
  16199=>"100011111",
  16200=>"010100111",
  16201=>"111100101",
  16202=>"110100100",
  16203=>"101001100",
  16204=>"111000011",
  16205=>"010101001",
  16206=>"000111100",
  16207=>"110111101",
  16208=>"101111111",
  16209=>"110000111",
  16210=>"110101111",
  16211=>"001100100",
  16212=>"100101100",
  16213=>"100111011",
  16214=>"101110101",
  16215=>"110110011",
  16216=>"010010010",
  16217=>"111100001",
  16218=>"100100101",
  16219=>"101100101",
  16220=>"010011110",
  16221=>"101101010",
  16222=>"010010001",
  16223=>"000000011",
  16224=>"111111110",
  16225=>"001111100",
  16226=>"111011111",
  16227=>"101111010",
  16228=>"101010100",
  16229=>"010100000",
  16230=>"110100010",
  16231=>"111000101",
  16232=>"011001011",
  16233=>"001010110",
  16234=>"111001010",
  16235=>"011100101",
  16236=>"010001010",
  16237=>"100001001",
  16238=>"111010101",
  16239=>"001011000",
  16240=>"111000011",
  16241=>"000001100",
  16242=>"011000110",
  16243=>"110101000",
  16244=>"111111101",
  16245=>"011101011",
  16246=>"000111100",
  16247=>"110000011",
  16248=>"101000110",
  16249=>"001001100",
  16250=>"010111010",
  16251=>"001101110",
  16252=>"101111001",
  16253=>"101001000",
  16254=>"000000000",
  16255=>"110010101",
  16256=>"101011010",
  16257=>"101010001",
  16258=>"101101100",
  16259=>"100101110",
  16260=>"110111001",
  16261=>"111010001",
  16262=>"110110011",
  16263=>"100110001",
  16264=>"000111010",
  16265=>"000001011",
  16266=>"011111011",
  16267=>"000011000",
  16268=>"111101111",
  16269=>"111001000",
  16270=>"111110010",
  16271=>"111110010",
  16272=>"000101101",
  16273=>"011110001",
  16274=>"100110111",
  16275=>"100000101",
  16276=>"010101110",
  16277=>"000111111",
  16278=>"011001111",
  16279=>"110001000",
  16280=>"011001111",
  16281=>"010111011",
  16282=>"100110100",
  16283=>"110100110",
  16284=>"001111010",
  16285=>"000001111",
  16286=>"111100011",
  16287=>"000100100",
  16288=>"000100110",
  16289=>"110001000",
  16290=>"111110101",
  16291=>"100101111",
  16292=>"010100000",
  16293=>"010011001",
  16294=>"011011000",
  16295=>"010001100",
  16296=>"001000111",
  16297=>"011101111",
  16298=>"010000001",
  16299=>"001101000",
  16300=>"000000111",
  16301=>"000000000",
  16302=>"111011110",
  16303=>"011001111",
  16304=>"001111010",
  16305=>"010000010",
  16306=>"001011100",
  16307=>"001000000",
  16308=>"101000110",
  16309=>"101001001",
  16310=>"101001011",
  16311=>"000111111",
  16312=>"001000000",
  16313=>"011111000",
  16314=>"000010011",
  16315=>"101110111",
  16316=>"110100100",
  16317=>"010010001",
  16318=>"000001000",
  16319=>"111101001",
  16320=>"010111111",
  16321=>"101110011",
  16322=>"111010001",
  16323=>"001010000",
  16324=>"110110111",
  16325=>"000100010",
  16326=>"111111011",
  16327=>"111111011",
  16328=>"000001101",
  16329=>"101101011",
  16330=>"110000000",
  16331=>"000011011",
  16332=>"001100101",
  16333=>"100000101",
  16334=>"010101001",
  16335=>"111111101",
  16336=>"001110010",
  16337=>"011001101",
  16338=>"000011111",
  16339=>"001001001",
  16340=>"000110100",
  16341=>"010011101",
  16342=>"010010101",
  16343=>"100010110",
  16344=>"110001111",
  16345=>"111000010",
  16346=>"111001001",
  16347=>"110010110",
  16348=>"001101110",
  16349=>"001110001",
  16350=>"001101011",
  16351=>"011100110",
  16352=>"110110011",
  16353=>"111011011",
  16354=>"010000110",
  16355=>"000111101",
  16356=>"100101111",
  16357=>"000010010",
  16358=>"110010001",
  16359=>"001101011",
  16360=>"001110001",
  16361=>"000110110",
  16362=>"001101101",
  16363=>"001010011",
  16364=>"010100010",
  16365=>"110010011",
  16366=>"110101100",
  16367=>"101001001",
  16368=>"111111010",
  16369=>"010011011",
  16370=>"000100111",
  16371=>"000001100",
  16372=>"100110011",
  16373=>"101100111",
  16374=>"000111111",
  16375=>"110000001",
  16376=>"111001111",
  16377=>"011110110",
  16378=>"100101000",
  16379=>"111111000",
  16380=>"011101110",
  16381=>"000000010",
  16382=>"001001101",
  16383=>"001101101",
  16384=>"000001010",
  16385=>"110111101",
  16386=>"001110011",
  16387=>"000110001",
  16388=>"000010010",
  16389=>"100110110",
  16390=>"101100101",
  16391=>"101101111",
  16392=>"110110000",
  16393=>"111111100",
  16394=>"100000111",
  16395=>"111001001",
  16396=>"101111110",
  16397=>"100111010",
  16398=>"111010000",
  16399=>"101101001",
  16400=>"010101100",
  16401=>"100100101",
  16402=>"011100010",
  16403=>"011111001",
  16404=>"000011110",
  16405=>"110101110",
  16406=>"100010001",
  16407=>"110110101",
  16408=>"111111111",
  16409=>"100100100",
  16410=>"011000000",
  16411=>"000010010",
  16412=>"111000100",
  16413=>"001000110",
  16414=>"001010101",
  16415=>"000000000",
  16416=>"110100001",
  16417=>"101101101",
  16418=>"101100010",
  16419=>"011101111",
  16420=>"000011111",
  16421=>"110000101",
  16422=>"010110011",
  16423=>"110111111",
  16424=>"011100101",
  16425=>"001101000",
  16426=>"001101010",
  16427=>"010111110",
  16428=>"110111001",
  16429=>"111010011",
  16430=>"110010010",
  16431=>"001000110",
  16432=>"001000000",
  16433=>"000000001",
  16434=>"111100110",
  16435=>"001010010",
  16436=>"001110110",
  16437=>"101111111",
  16438=>"110100100",
  16439=>"111010111",
  16440=>"111111111",
  16441=>"001110110",
  16442=>"011010010",
  16443=>"000011110",
  16444=>"001110000",
  16445=>"110001000",
  16446=>"111101101",
  16447=>"110001000",
  16448=>"010110101",
  16449=>"101111111",
  16450=>"111001111",
  16451=>"011000110",
  16452=>"000111010",
  16453=>"101011011",
  16454=>"101011001",
  16455=>"111110000",
  16456=>"111111101",
  16457=>"000001010",
  16458=>"110100000",
  16459=>"101001000",
  16460=>"001111010",
  16461=>"101010101",
  16462=>"110011000",
  16463=>"101001100",
  16464=>"100110000",
  16465=>"110010110",
  16466=>"100111110",
  16467=>"010101000",
  16468=>"000010101",
  16469=>"011101001",
  16470=>"010000100",
  16471=>"100101000",
  16472=>"011101110",
  16473=>"110110101",
  16474=>"001100001",
  16475=>"101000101",
  16476=>"001010100",
  16477=>"111001111",
  16478=>"111100000",
  16479=>"101111010",
  16480=>"111100000",
  16481=>"100101110",
  16482=>"110011100",
  16483=>"000001101",
  16484=>"001001100",
  16485=>"011001100",
  16486=>"101100100",
  16487=>"000001010",
  16488=>"000001110",
  16489=>"011100111",
  16490=>"111001001",
  16491=>"111011010",
  16492=>"000110000",
  16493=>"100000100",
  16494=>"111100011",
  16495=>"000101011",
  16496=>"000100000",
  16497=>"000111010",
  16498=>"111101000",
  16499=>"110111111",
  16500=>"100001001",
  16501=>"110001010",
  16502=>"110011001",
  16503=>"001111010",
  16504=>"110011000",
  16505=>"000100101",
  16506=>"100100000",
  16507=>"110100010",
  16508=>"100010000",
  16509=>"010011000",
  16510=>"110010110",
  16511=>"111110111",
  16512=>"001001100",
  16513=>"111111010",
  16514=>"001111000",
  16515=>"000100111",
  16516=>"000111111",
  16517=>"111100111",
  16518=>"010101110",
  16519=>"111111101",
  16520=>"100010100",
  16521=>"001001001",
  16522=>"011010001",
  16523=>"000100110",
  16524=>"111001000",
  16525=>"110111001",
  16526=>"001011000",
  16527=>"001001100",
  16528=>"100100111",
  16529=>"011110101",
  16530=>"111010100",
  16531=>"011101000",
  16532=>"011100000",
  16533=>"100011011",
  16534=>"011011000",
  16535=>"110000101",
  16536=>"101001001",
  16537=>"101000011",
  16538=>"110011110",
  16539=>"110101011",
  16540=>"101110111",
  16541=>"010100010",
  16542=>"001001100",
  16543=>"011011101",
  16544=>"010100111",
  16545=>"000101111",
  16546=>"100011110",
  16547=>"110010110",
  16548=>"100000111",
  16549=>"010111010",
  16550=>"111100011",
  16551=>"001101110",
  16552=>"101111110",
  16553=>"011000101",
  16554=>"011011100",
  16555=>"101101110",
  16556=>"000011010",
  16557=>"011000100",
  16558=>"101111011",
  16559=>"000111000",
  16560=>"100011011",
  16561=>"110100110",
  16562=>"011000111",
  16563=>"011110001",
  16564=>"111100000",
  16565=>"110110000",
  16566=>"010000111",
  16567=>"110111110",
  16568=>"100011101",
  16569=>"111001001",
  16570=>"101111111",
  16571=>"001101111",
  16572=>"100101110",
  16573=>"010101111",
  16574=>"110011111",
  16575=>"100011001",
  16576=>"010011100",
  16577=>"001100000",
  16578=>"101011010",
  16579=>"100000101",
  16580=>"000100101",
  16581=>"011000011",
  16582=>"101001010",
  16583=>"101011111",
  16584=>"101000011",
  16585=>"011001111",
  16586=>"111001000",
  16587=>"011101001",
  16588=>"111110001",
  16589=>"001101001",
  16590=>"001101011",
  16591=>"000100001",
  16592=>"100010110",
  16593=>"011101100",
  16594=>"011010110",
  16595=>"100110111",
  16596=>"110011100",
  16597=>"000100110",
  16598=>"101010101",
  16599=>"101100001",
  16600=>"000010101",
  16601=>"001011001",
  16602=>"001001010",
  16603=>"010010100",
  16604=>"001001001",
  16605=>"100110110",
  16606=>"110100110",
  16607=>"000000001",
  16608=>"000011000",
  16609=>"000100011",
  16610=>"100101010",
  16611=>"101100101",
  16612=>"010110110",
  16613=>"000110011",
  16614=>"011001011",
  16615=>"000001010",
  16616=>"010111101",
  16617=>"010011101",
  16618=>"001011011",
  16619=>"111000011",
  16620=>"000011010",
  16621=>"001010111",
  16622=>"011000101",
  16623=>"110011001",
  16624=>"001110011",
  16625=>"000010000",
  16626=>"000111001",
  16627=>"001101000",
  16628=>"111010110",
  16629=>"110010000",
  16630=>"001001100",
  16631=>"110100100",
  16632=>"111110011",
  16633=>"001110011",
  16634=>"111000010",
  16635=>"001010010",
  16636=>"010000010",
  16637=>"000001100",
  16638=>"001111101",
  16639=>"011000001",
  16640=>"100010010",
  16641=>"011011011",
  16642=>"001101111",
  16643=>"111000101",
  16644=>"011100000",
  16645=>"001110111",
  16646=>"000101100",
  16647=>"101101011",
  16648=>"100101100",
  16649=>"100000000",
  16650=>"011011001",
  16651=>"111100101",
  16652=>"000100010",
  16653=>"000100111",
  16654=>"000001010",
  16655=>"010101110",
  16656=>"101010100",
  16657=>"010010010",
  16658=>"111100110",
  16659=>"110011011",
  16660=>"010101100",
  16661=>"110000110",
  16662=>"010111000",
  16663=>"100000110",
  16664=>"011100101",
  16665=>"101001001",
  16666=>"101001110",
  16667=>"001100111",
  16668=>"001110101",
  16669=>"100010111",
  16670=>"100110110",
  16671=>"001101101",
  16672=>"011110111",
  16673=>"011000001",
  16674=>"100001001",
  16675=>"001101100",
  16676=>"011100101",
  16677=>"000110001",
  16678=>"100101101",
  16679=>"000100001",
  16680=>"111111111",
  16681=>"001001110",
  16682=>"000010001",
  16683=>"011111100",
  16684=>"000011111",
  16685=>"100101001",
  16686=>"101000100",
  16687=>"000111110",
  16688=>"010100001",
  16689=>"011100101",
  16690=>"010011110",
  16691=>"000001100",
  16692=>"101000001",
  16693=>"001011111",
  16694=>"011110111",
  16695=>"101000101",
  16696=>"011101111",
  16697=>"001100100",
  16698=>"111100100",
  16699=>"101001001",
  16700=>"000100011",
  16701=>"110110100",
  16702=>"111011000",
  16703=>"111111111",
  16704=>"111100001",
  16705=>"110011110",
  16706=>"111111011",
  16707=>"110010110",
  16708=>"000000010",
  16709=>"010110101",
  16710=>"011000111",
  16711=>"101010101",
  16712=>"001010111",
  16713=>"100100011",
  16714=>"010001110",
  16715=>"000110000",
  16716=>"111011000",
  16717=>"110101110",
  16718=>"011011111",
  16719=>"111101111",
  16720=>"100001010",
  16721=>"011001100",
  16722=>"111011001",
  16723=>"101011011",
  16724=>"000100100",
  16725=>"111111101",
  16726=>"100100010",
  16727=>"101110010",
  16728=>"000110110",
  16729=>"110110010",
  16730=>"111110111",
  16731=>"110001101",
  16732=>"010011011",
  16733=>"100010010",
  16734=>"011010101",
  16735=>"010111001",
  16736=>"010101001",
  16737=>"100110111",
  16738=>"001001010",
  16739=>"001100000",
  16740=>"111000000",
  16741=>"110000001",
  16742=>"010111000",
  16743=>"101000001",
  16744=>"011001110",
  16745=>"100111100",
  16746=>"110100010",
  16747=>"010010001",
  16748=>"101111010",
  16749=>"100110111",
  16750=>"010100011",
  16751=>"110011101",
  16752=>"100100000",
  16753=>"010100101",
  16754=>"010101010",
  16755=>"111011000",
  16756=>"110010111",
  16757=>"010110111",
  16758=>"010110011",
  16759=>"101011010",
  16760=>"000111001",
  16761=>"100010101",
  16762=>"100001000",
  16763=>"100010011",
  16764=>"000110011",
  16765=>"000100000",
  16766=>"011110110",
  16767=>"101101101",
  16768=>"001001000",
  16769=>"011010100",
  16770=>"011110010",
  16771=>"000101010",
  16772=>"011100000",
  16773=>"111111000",
  16774=>"111100101",
  16775=>"011110000",
  16776=>"001100010",
  16777=>"101010010",
  16778=>"100111001",
  16779=>"000111101",
  16780=>"010011011",
  16781=>"100111000",
  16782=>"100111100",
  16783=>"100001100",
  16784=>"110010101",
  16785=>"000001110",
  16786=>"111101000",
  16787=>"100000011",
  16788=>"001010000",
  16789=>"110000100",
  16790=>"100001000",
  16791=>"111000010",
  16792=>"001101000",
  16793=>"000101101",
  16794=>"010100011",
  16795=>"010000111",
  16796=>"111000111",
  16797=>"001110001",
  16798=>"110010110",
  16799=>"010110110",
  16800=>"001001001",
  16801=>"110000111",
  16802=>"000001101",
  16803=>"110111001",
  16804=>"010001110",
  16805=>"111111000",
  16806=>"010100111",
  16807=>"110001100",
  16808=>"110111010",
  16809=>"110011001",
  16810=>"000000110",
  16811=>"111110101",
  16812=>"100100000",
  16813=>"111100001",
  16814=>"000111010",
  16815=>"011000101",
  16816=>"000101011",
  16817=>"110000100",
  16818=>"000111000",
  16819=>"101001000",
  16820=>"011011110",
  16821=>"010001110",
  16822=>"101111010",
  16823=>"000001000",
  16824=>"010011101",
  16825=>"011101000",
  16826=>"010001011",
  16827=>"010101111",
  16828=>"111111000",
  16829=>"010110001",
  16830=>"100000000",
  16831=>"011110001",
  16832=>"010010110",
  16833=>"010100110",
  16834=>"110011001",
  16835=>"011000000",
  16836=>"011111110",
  16837=>"000000000",
  16838=>"001110100",
  16839=>"111001011",
  16840=>"110000000",
  16841=>"011001110",
  16842=>"101101101",
  16843=>"001101111",
  16844=>"010111101",
  16845=>"100001101",
  16846=>"110100111",
  16847=>"010110010",
  16848=>"110111011",
  16849=>"010010000",
  16850=>"111010111",
  16851=>"111111100",
  16852=>"011010111",
  16853=>"001000110",
  16854=>"000010111",
  16855=>"110000111",
  16856=>"101011010",
  16857=>"010100000",
  16858=>"000010101",
  16859=>"100100010",
  16860=>"001101001",
  16861=>"100011011",
  16862=>"111010010",
  16863=>"000000001",
  16864=>"011010011",
  16865=>"011111011",
  16866=>"000100110",
  16867=>"001100100",
  16868=>"110001110",
  16869=>"100000101",
  16870=>"101101100",
  16871=>"111001011",
  16872=>"011101110",
  16873=>"001011100",
  16874=>"110111111",
  16875=>"010110111",
  16876=>"000111010",
  16877=>"000000011",
  16878=>"001100000",
  16879=>"011100011",
  16880=>"101000110",
  16881=>"111100101",
  16882=>"000110000",
  16883=>"100101111",
  16884=>"000010011",
  16885=>"101000010",
  16886=>"110001011",
  16887=>"100100110",
  16888=>"011101110",
  16889=>"100011010",
  16890=>"101101110",
  16891=>"011011010",
  16892=>"000000110",
  16893=>"001000010",
  16894=>"011100010",
  16895=>"011010011",
  16896=>"111111111",
  16897=>"101100110",
  16898=>"001000010",
  16899=>"110011110",
  16900=>"000110111",
  16901=>"110010001",
  16902=>"100111001",
  16903=>"001110011",
  16904=>"101000110",
  16905=>"000010010",
  16906=>"100010011",
  16907=>"011011110",
  16908=>"001001111",
  16909=>"001011100",
  16910=>"100111010",
  16911=>"000010001",
  16912=>"011110101",
  16913=>"100110111",
  16914=>"101001011",
  16915=>"111111010",
  16916=>"000010010",
  16917=>"110010111",
  16918=>"101110001",
  16919=>"001100000",
  16920=>"111001110",
  16921=>"100000111",
  16922=>"101100000",
  16923=>"111110111",
  16924=>"001110110",
  16925=>"100110110",
  16926=>"111000011",
  16927=>"010110100",
  16928=>"010011000",
  16929=>"111111001",
  16930=>"101000000",
  16931=>"101101010",
  16932=>"101111000",
  16933=>"111111110",
  16934=>"000100001",
  16935=>"110010111",
  16936=>"101110010",
  16937=>"111101010",
  16938=>"101001100",
  16939=>"100000000",
  16940=>"001101011",
  16941=>"010111011",
  16942=>"000010101",
  16943=>"001010000",
  16944=>"111001000",
  16945=>"110110100",
  16946=>"001101101",
  16947=>"100100110",
  16948=>"011101100",
  16949=>"101100010",
  16950=>"001100010",
  16951=>"000011100",
  16952=>"000110111",
  16953=>"101001100",
  16954=>"101011010",
  16955=>"011001101",
  16956=>"010111110",
  16957=>"000001110",
  16958=>"111000101",
  16959=>"101011110",
  16960=>"101110111",
  16961=>"111101011",
  16962=>"010101111",
  16963=>"010010001",
  16964=>"000111100",
  16965=>"110111110",
  16966=>"101001010",
  16967=>"000100000",
  16968=>"010110100",
  16969=>"000010011",
  16970=>"111101010",
  16971=>"001101010",
  16972=>"100010001",
  16973=>"101001011",
  16974=>"001111010",
  16975=>"111110110",
  16976=>"000111101",
  16977=>"011011101",
  16978=>"110110011",
  16979=>"111111001",
  16980=>"111100100",
  16981=>"111001000",
  16982=>"011000010",
  16983=>"011110111",
  16984=>"001001000",
  16985=>"110100111",
  16986=>"010000111",
  16987=>"010111101",
  16988=>"000010110",
  16989=>"110010110",
  16990=>"110111001",
  16991=>"110110101",
  16992=>"110001011",
  16993=>"001100110",
  16994=>"111010100",
  16995=>"001000101",
  16996=>"111000000",
  16997=>"111101100",
  16998=>"011011001",
  16999=>"100010000",
  17000=>"011011000",
  17001=>"110001101",
  17002=>"111001111",
  17003=>"110011001",
  17004=>"101101001",
  17005=>"000110001",
  17006=>"010100110",
  17007=>"111111110",
  17008=>"110010000",
  17009=>"010101010",
  17010=>"110100001",
  17011=>"010010100",
  17012=>"000110100",
  17013=>"000111111",
  17014=>"000101011",
  17015=>"111100111",
  17016=>"000000100",
  17017=>"100110101",
  17018=>"111010011",
  17019=>"001000011",
  17020=>"110101011",
  17021=>"000010000",
  17022=>"001110111",
  17023=>"111110101",
  17024=>"010101011",
  17025=>"100110110",
  17026=>"101001110",
  17027=>"001100000",
  17028=>"100101001",
  17029=>"010110000",
  17030=>"010010100",
  17031=>"111110000",
  17032=>"000010111",
  17033=>"110011001",
  17034=>"110111111",
  17035=>"100011111",
  17036=>"010001011",
  17037=>"101111011",
  17038=>"000100100",
  17039=>"010101001",
  17040=>"100101100",
  17041=>"100011011",
  17042=>"111001011",
  17043=>"110110011",
  17044=>"101000100",
  17045=>"010011110",
  17046=>"101111101",
  17047=>"001000110",
  17048=>"111001100",
  17049=>"100110010",
  17050=>"011000101",
  17051=>"001000010",
  17052=>"100110000",
  17053=>"110100110",
  17054=>"101101010",
  17055=>"011101101",
  17056=>"011100101",
  17057=>"010010001",
  17058=>"100000111",
  17059=>"110011011",
  17060=>"010111110",
  17061=>"010010101",
  17062=>"101110100",
  17063=>"100111110",
  17064=>"000100000",
  17065=>"110110000",
  17066=>"101000001",
  17067=>"110001011",
  17068=>"100011011",
  17069=>"010110011",
  17070=>"001010000",
  17071=>"011011111",
  17072=>"100000010",
  17073=>"001000011",
  17074=>"100001110",
  17075=>"111001101",
  17076=>"011001010",
  17077=>"011011010",
  17078=>"010110000",
  17079=>"111100001",
  17080=>"010100111",
  17081=>"101100011",
  17082=>"010011110",
  17083=>"000110001",
  17084=>"110000110",
  17085=>"000000011",
  17086=>"111011110",
  17087=>"001110110",
  17088=>"110000011",
  17089=>"010001011",
  17090=>"001110111",
  17091=>"101001001",
  17092=>"111001111",
  17093=>"110101111",
  17094=>"100100000",
  17095=>"001001111",
  17096=>"111001111",
  17097=>"111111101",
  17098=>"110001100",
  17099=>"000011001",
  17100=>"011110101",
  17101=>"011001011",
  17102=>"000001010",
  17103=>"010111110",
  17104=>"111010010",
  17105=>"100101101",
  17106=>"110110110",
  17107=>"011100100",
  17108=>"001101110",
  17109=>"010100101",
  17110=>"011010011",
  17111=>"001001010",
  17112=>"001011101",
  17113=>"101100100",
  17114=>"011000001",
  17115=>"011001010",
  17116=>"101001100",
  17117=>"111010100",
  17118=>"101011111",
  17119=>"110001101",
  17120=>"110101010",
  17121=>"001000101",
  17122=>"000011101",
  17123=>"001001010",
  17124=>"011100110",
  17125=>"111111001",
  17126=>"111000010",
  17127=>"100001110",
  17128=>"101010111",
  17129=>"010101110",
  17130=>"001000000",
  17131=>"010110011",
  17132=>"001010011",
  17133=>"011111100",
  17134=>"110100010",
  17135=>"001000111",
  17136=>"001110001",
  17137=>"010001001",
  17138=>"101111100",
  17139=>"111111011",
  17140=>"011011001",
  17141=>"000100110",
  17142=>"000000000",
  17143=>"011111001",
  17144=>"111110011",
  17145=>"101010100",
  17146=>"101010100",
  17147=>"110000001",
  17148=>"101101000",
  17149=>"011111011",
  17150=>"111101000",
  17151=>"010011101",
  17152=>"001101000",
  17153=>"001100110",
  17154=>"001011110",
  17155=>"000111110",
  17156=>"110101111",
  17157=>"110001000",
  17158=>"111001111",
  17159=>"011001101",
  17160=>"111011101",
  17161=>"101101111",
  17162=>"101011011",
  17163=>"101101111",
  17164=>"011100101",
  17165=>"110000001",
  17166=>"101000000",
  17167=>"010101010",
  17168=>"000000011",
  17169=>"110111010",
  17170=>"000110000",
  17171=>"110111110",
  17172=>"111101110",
  17173=>"010010100",
  17174=>"100100001",
  17175=>"101110100",
  17176=>"010000011",
  17177=>"101000000",
  17178=>"101101000",
  17179=>"011001011",
  17180=>"010011011",
  17181=>"011100010",
  17182=>"000111110",
  17183=>"010100010",
  17184=>"110101100",
  17185=>"110110011",
  17186=>"000000100",
  17187=>"001101001",
  17188=>"110001000",
  17189=>"001100000",
  17190=>"111100110",
  17191=>"111010010",
  17192=>"010000001",
  17193=>"101001111",
  17194=>"110000111",
  17195=>"001001110",
  17196=>"001111111",
  17197=>"001101010",
  17198=>"111010100",
  17199=>"011101000",
  17200=>"010001001",
  17201=>"100111110",
  17202=>"001111111",
  17203=>"110011101",
  17204=>"100110111",
  17205=>"101011110",
  17206=>"001001011",
  17207=>"001000010",
  17208=>"111111011",
  17209=>"100011000",
  17210=>"111111111",
  17211=>"111100011",
  17212=>"010001111",
  17213=>"010111000",
  17214=>"101111001",
  17215=>"001011110",
  17216=>"101010110",
  17217=>"011011000",
  17218=>"111101110",
  17219=>"001010000",
  17220=>"111110000",
  17221=>"111111110",
  17222=>"001101001",
  17223=>"111001111",
  17224=>"101110111",
  17225=>"001001001",
  17226=>"010110110",
  17227=>"010100100",
  17228=>"011011100",
  17229=>"010010011",
  17230=>"101001001",
  17231=>"101100011",
  17232=>"001001111",
  17233=>"101110111",
  17234=>"000010111",
  17235=>"001001000",
  17236=>"111110101",
  17237=>"101101101",
  17238=>"000011111",
  17239=>"110000001",
  17240=>"000000111",
  17241=>"111100000",
  17242=>"101001001",
  17243=>"011010000",
  17244=>"110011001",
  17245=>"100111101",
  17246=>"000100110",
  17247=>"111000010",
  17248=>"101111011",
  17249=>"111110111",
  17250=>"000100001",
  17251=>"101001100",
  17252=>"100011000",
  17253=>"010011011",
  17254=>"110001101",
  17255=>"100110100",
  17256=>"111110000",
  17257=>"100100101",
  17258=>"000100110",
  17259=>"110000000",
  17260=>"100101010",
  17261=>"011001111",
  17262=>"101101101",
  17263=>"010101011",
  17264=>"000010110",
  17265=>"101100000",
  17266=>"100110100",
  17267=>"010110011",
  17268=>"001010000",
  17269=>"011011100",
  17270=>"101010111",
  17271=>"110001001",
  17272=>"111111100",
  17273=>"010111110",
  17274=>"111101011",
  17275=>"100011011",
  17276=>"001111110",
  17277=>"110101001",
  17278=>"111001001",
  17279=>"110011001",
  17280=>"100011001",
  17281=>"011101111",
  17282=>"100011011",
  17283=>"011110011",
  17284=>"111010111",
  17285=>"111101100",
  17286=>"100110111",
  17287=>"000100010",
  17288=>"110011001",
  17289=>"000111011",
  17290=>"010001100",
  17291=>"010011100",
  17292=>"111111101",
  17293=>"111011000",
  17294=>"110011000",
  17295=>"000111000",
  17296=>"001010010",
  17297=>"110010111",
  17298=>"000001100",
  17299=>"101111110",
  17300=>"011011011",
  17301=>"110111100",
  17302=>"000110010",
  17303=>"101001010",
  17304=>"110101111",
  17305=>"110110111",
  17306=>"010001010",
  17307=>"110011111",
  17308=>"110101101",
  17309=>"111000111",
  17310=>"111110101",
  17311=>"011000001",
  17312=>"101101100",
  17313=>"011110000",
  17314=>"100110011",
  17315=>"111100000",
  17316=>"111101001",
  17317=>"010000100",
  17318=>"000001111",
  17319=>"010011110",
  17320=>"001000110",
  17321=>"000010111",
  17322=>"011010100",
  17323=>"000111110",
  17324=>"011011011",
  17325=>"000110110",
  17326=>"101011100",
  17327=>"110101000",
  17328=>"010111010",
  17329=>"110100111",
  17330=>"100111011",
  17331=>"100010110",
  17332=>"001010011",
  17333=>"100111111",
  17334=>"111110110",
  17335=>"101101110",
  17336=>"000110000",
  17337=>"111000011",
  17338=>"111101000",
  17339=>"100100100",
  17340=>"100010101",
  17341=>"011000101",
  17342=>"101101010",
  17343=>"000101000",
  17344=>"100000011",
  17345=>"011101100",
  17346=>"001110100",
  17347=>"011001100",
  17348=>"101010000",
  17349=>"101011101",
  17350=>"111010000",
  17351=>"011010001",
  17352=>"000101101",
  17353=>"001011101",
  17354=>"011111001",
  17355=>"001011010",
  17356=>"100110110",
  17357=>"000011111",
  17358=>"011100111",
  17359=>"111111110",
  17360=>"011100000",
  17361=>"001110111",
  17362=>"101111000",
  17363=>"100110101",
  17364=>"101100101",
  17365=>"010100001",
  17366=>"100111010",
  17367=>"000011010",
  17368=>"000000001",
  17369=>"111000110",
  17370=>"001011110",
  17371=>"101100011",
  17372=>"011100110",
  17373=>"000001111",
  17374=>"000100101",
  17375=>"100011100",
  17376=>"000101010",
  17377=>"101110100",
  17378=>"010100110",
  17379=>"111110000",
  17380=>"000010011",
  17381=>"011010100",
  17382=>"010111000",
  17383=>"010101101",
  17384=>"100011101",
  17385=>"000110111",
  17386=>"000001101",
  17387=>"110011100",
  17388=>"000001110",
  17389=>"110110101",
  17390=>"101111101",
  17391=>"011101000",
  17392=>"100111110",
  17393=>"101111000",
  17394=>"111000110",
  17395=>"001111101",
  17396=>"000101010",
  17397=>"111010111",
  17398=>"001010000",
  17399=>"011101010",
  17400=>"111011101",
  17401=>"100100010",
  17402=>"100000100",
  17403=>"101101100",
  17404=>"011011000",
  17405=>"111101111",
  17406=>"100100101",
  17407=>"101010111",
  17408=>"110101110",
  17409=>"001000000",
  17410=>"110000110",
  17411=>"111101100",
  17412=>"111110101",
  17413=>"011101110",
  17414=>"001001001",
  17415=>"111101101",
  17416=>"111101010",
  17417=>"011110001",
  17418=>"101111110",
  17419=>"011100100",
  17420=>"001010000",
  17421=>"001101101",
  17422=>"011000100",
  17423=>"110101100",
  17424=>"111110111",
  17425=>"000000011",
  17426=>"011101011",
  17427=>"010101001",
  17428=>"010101011",
  17429=>"110010010",
  17430=>"110111110",
  17431=>"010001110",
  17432=>"001100110",
  17433=>"010111101",
  17434=>"100110010",
  17435=>"011001111",
  17436=>"111110110",
  17437=>"101001101",
  17438=>"001100010",
  17439=>"010011011",
  17440=>"110101111",
  17441=>"010000000",
  17442=>"011100011",
  17443=>"110111100",
  17444=>"111001111",
  17445=>"010001000",
  17446=>"001101110",
  17447=>"011100011",
  17448=>"001011011",
  17449=>"111101101",
  17450=>"111110000",
  17451=>"110111011",
  17452=>"101101001",
  17453=>"011000101",
  17454=>"110011001",
  17455=>"101101001",
  17456=>"011011101",
  17457=>"111110111",
  17458=>"101010001",
  17459=>"101000000",
  17460=>"101110011",
  17461=>"001101111",
  17462=>"100111000",
  17463=>"111011101",
  17464=>"100010011",
  17465=>"010101110",
  17466=>"001000101",
  17467=>"000001011",
  17468=>"001100000",
  17469=>"100011111",
  17470=>"111100101",
  17471=>"101001101",
  17472=>"001100010",
  17473=>"100001100",
  17474=>"001011100",
  17475=>"000011000",
  17476=>"001001110",
  17477=>"111111011",
  17478=>"000110011",
  17479=>"110000000",
  17480=>"110101010",
  17481=>"000111100",
  17482=>"010100100",
  17483=>"001101001",
  17484=>"001101101",
  17485=>"111110111",
  17486=>"110011110",
  17487=>"010111000",
  17488=>"010111111",
  17489=>"011001010",
  17490=>"011011011",
  17491=>"000011011",
  17492=>"010001100",
  17493=>"011101110",
  17494=>"110110101",
  17495=>"100100100",
  17496=>"101000011",
  17497=>"111111101",
  17498=>"001000110",
  17499=>"101000110",
  17500=>"110001011",
  17501=>"010101101",
  17502=>"110011010",
  17503=>"101000000",
  17504=>"010110000",
  17505=>"101101011",
  17506=>"000011011",
  17507=>"010110010",
  17508=>"011110000",
  17509=>"110010100",
  17510=>"000111101",
  17511=>"101110000",
  17512=>"110011001",
  17513=>"111010011",
  17514=>"010001110",
  17515=>"011101100",
  17516=>"110001011",
  17517=>"111100100",
  17518=>"000101000",
  17519=>"100110001",
  17520=>"011001111",
  17521=>"101010001",
  17522=>"001001101",
  17523=>"011111111",
  17524=>"001000000",
  17525=>"111000111",
  17526=>"110011011",
  17527=>"101101011",
  17528=>"110101100",
  17529=>"100100111",
  17530=>"111111011",
  17531=>"101100001",
  17532=>"011000101",
  17533=>"100101011",
  17534=>"010011111",
  17535=>"011110101",
  17536=>"010010110",
  17537=>"101001100",
  17538=>"101001001",
  17539=>"001001011",
  17540=>"000101101",
  17541=>"010000001",
  17542=>"100010010",
  17543=>"001110001",
  17544=>"110100101",
  17545=>"010111100",
  17546=>"110011010",
  17547=>"000110000",
  17548=>"101101110",
  17549=>"010100010",
  17550=>"111101000",
  17551=>"000100010",
  17552=>"101011000",
  17553=>"100111010",
  17554=>"111011010",
  17555=>"001101100",
  17556=>"000001011",
  17557=>"000111001",
  17558=>"001011001",
  17559=>"001010101",
  17560=>"000011101",
  17561=>"111110011",
  17562=>"001110111",
  17563=>"011100111",
  17564=>"000011000",
  17565=>"011111110",
  17566=>"100110000",
  17567=>"100111101",
  17568=>"000110001",
  17569=>"001100010",
  17570=>"001100001",
  17571=>"110000010",
  17572=>"101110010",
  17573=>"110110011",
  17574=>"010001011",
  17575=>"101110001",
  17576=>"100010000",
  17577=>"111111101",
  17578=>"000010010",
  17579=>"000000101",
  17580=>"110011101",
  17581=>"111001111",
  17582=>"010101011",
  17583=>"000001000",
  17584=>"001101011",
  17585=>"101001110",
  17586=>"001000011",
  17587=>"000001001",
  17588=>"110100011",
  17589=>"000011111",
  17590=>"000001000",
  17591=>"111111001",
  17592=>"101001100",
  17593=>"000001010",
  17594=>"001010011",
  17595=>"100111001",
  17596=>"010100000",
  17597=>"011011111",
  17598=>"001001010",
  17599=>"000110000",
  17600=>"011110101",
  17601=>"001101001",
  17602=>"111010111",
  17603=>"101010111",
  17604=>"100100000",
  17605=>"110101001",
  17606=>"001001101",
  17607=>"100100111",
  17608=>"011110101",
  17609=>"100010000",
  17610=>"011111101",
  17611=>"001100101",
  17612=>"010110100",
  17613=>"000101000",
  17614=>"001001100",
  17615=>"000000001",
  17616=>"111100011",
  17617=>"001101000",
  17618=>"010000101",
  17619=>"000101111",
  17620=>"011101111",
  17621=>"110000010",
  17622=>"110011111",
  17623=>"111011011",
  17624=>"110100100",
  17625=>"100111000",
  17626=>"100001000",
  17627=>"100111100",
  17628=>"000100100",
  17629=>"100000110",
  17630=>"000100110",
  17631=>"111111110",
  17632=>"100101011",
  17633=>"101100000",
  17634=>"010011001",
  17635=>"101010011",
  17636=>"010010111",
  17637=>"011011001",
  17638=>"000000000",
  17639=>"111001101",
  17640=>"000101000",
  17641=>"001100100",
  17642=>"001011101",
  17643=>"111010000",
  17644=>"111101010",
  17645=>"110011010",
  17646=>"011010010",
  17647=>"001001011",
  17648=>"111001111",
  17649=>"110110111",
  17650=>"111011101",
  17651=>"101001001",
  17652=>"100111001",
  17653=>"000100100",
  17654=>"001011100",
  17655=>"000001000",
  17656=>"001011111",
  17657=>"100000100",
  17658=>"001110011",
  17659=>"101010001",
  17660=>"111101010",
  17661=>"101011100",
  17662=>"000001001",
  17663=>"011010111",
  17664=>"110100001",
  17665=>"011100101",
  17666=>"111010101",
  17667=>"000111011",
  17668=>"101111110",
  17669=>"000001101",
  17670=>"001000101",
  17671=>"000001110",
  17672=>"100111010",
  17673=>"010000011",
  17674=>"000001001",
  17675=>"001101100",
  17676=>"100100101",
  17677=>"010010001",
  17678=>"100001100",
  17679=>"111101000",
  17680=>"000000111",
  17681=>"010111001",
  17682=>"000000101",
  17683=>"111100011",
  17684=>"000000101",
  17685=>"011110000",
  17686=>"101010011",
  17687=>"010101011",
  17688=>"000011001",
  17689=>"010100110",
  17690=>"011111010",
  17691=>"111001000",
  17692=>"010010010",
  17693=>"001101100",
  17694=>"001010100",
  17695=>"000000100",
  17696=>"000000011",
  17697=>"100000110",
  17698=>"100001111",
  17699=>"010010101",
  17700=>"001110110",
  17701=>"000000011",
  17702=>"001011101",
  17703=>"110010010",
  17704=>"110011000",
  17705=>"110001010",
  17706=>"001101010",
  17707=>"000111111",
  17708=>"010001000",
  17709=>"111011110",
  17710=>"111101011",
  17711=>"010001000",
  17712=>"001011000",
  17713=>"010001101",
  17714=>"001100001",
  17715=>"011010111",
  17716=>"001001101",
  17717=>"001000000",
  17718=>"001100001",
  17719=>"101101011",
  17720=>"000011001",
  17721=>"000011000",
  17722=>"000011010",
  17723=>"011001001",
  17724=>"101100010",
  17725=>"111100010",
  17726=>"111111111",
  17727=>"101110111",
  17728=>"010000000",
  17729=>"001100000",
  17730=>"100110100",
  17731=>"101001110",
  17732=>"010101010",
  17733=>"110100001",
  17734=>"000010000",
  17735=>"111001110",
  17736=>"100101100",
  17737=>"001101111",
  17738=>"111010010",
  17739=>"010001011",
  17740=>"000000001",
  17741=>"111111010",
  17742=>"000001001",
  17743=>"011011000",
  17744=>"000000110",
  17745=>"011010010",
  17746=>"001000101",
  17747=>"100001101",
  17748=>"001000110",
  17749=>"101011111",
  17750=>"100100100",
  17751=>"001000101",
  17752=>"001001000",
  17753=>"110111101",
  17754=>"110000001",
  17755=>"101001110",
  17756=>"100010011",
  17757=>"010100010",
  17758=>"111001010",
  17759=>"010000010",
  17760=>"101001001",
  17761=>"010100110",
  17762=>"011111100",
  17763=>"001010000",
  17764=>"111100100",
  17765=>"110001101",
  17766=>"011110100",
  17767=>"111111101",
  17768=>"011110011",
  17769=>"011000101",
  17770=>"000111010",
  17771=>"101110000",
  17772=>"111011011",
  17773=>"010000010",
  17774=>"001011100",
  17775=>"010011010",
  17776=>"100001001",
  17777=>"111011000",
  17778=>"001101100",
  17779=>"000100100",
  17780=>"111111011",
  17781=>"100000010",
  17782=>"101100110",
  17783=>"110000011",
  17784=>"001011011",
  17785=>"010000101",
  17786=>"000000110",
  17787=>"110000000",
  17788=>"001000010",
  17789=>"111111011",
  17790=>"000100110",
  17791=>"000001100",
  17792=>"110011101",
  17793=>"011011110",
  17794=>"101000111",
  17795=>"001101010",
  17796=>"101110001",
  17797=>"010001001",
  17798=>"011100000",
  17799=>"000000010",
  17800=>"010001000",
  17801=>"000000110",
  17802=>"101001010",
  17803=>"110000000",
  17804=>"010001111",
  17805=>"001000100",
  17806=>"111111001",
  17807=>"010010100",
  17808=>"001001001",
  17809=>"010101000",
  17810=>"001001010",
  17811=>"000011011",
  17812=>"101100111",
  17813=>"100000101",
  17814=>"011111000",
  17815=>"011011001",
  17816=>"101100101",
  17817=>"000110011",
  17818=>"010101110",
  17819=>"001000110",
  17820=>"011111000",
  17821=>"010110010",
  17822=>"001000000",
  17823=>"000101000",
  17824=>"101100000",
  17825=>"101100011",
  17826=>"100001010",
  17827=>"000000011",
  17828=>"001111100",
  17829=>"110000011",
  17830=>"001011011",
  17831=>"101011100",
  17832=>"011101110",
  17833=>"000100001",
  17834=>"101101000",
  17835=>"110000110",
  17836=>"010010101",
  17837=>"101101101",
  17838=>"011101001",
  17839=>"001110100",
  17840=>"010111100",
  17841=>"000110100",
  17842=>"010000111",
  17843=>"010011100",
  17844=>"001101000",
  17845=>"011100100",
  17846=>"001110111",
  17847=>"111110100",
  17848=>"011100000",
  17849=>"111110011",
  17850=>"011000000",
  17851=>"111000111",
  17852=>"111101101",
  17853=>"110110001",
  17854=>"101101001",
  17855=>"101001001",
  17856=>"110011100",
  17857=>"110000001",
  17858=>"101111100",
  17859=>"100101111",
  17860=>"111111110",
  17861=>"010000100",
  17862=>"111110111",
  17863=>"100011010",
  17864=>"001011001",
  17865=>"110011101",
  17866=>"110011010",
  17867=>"001001001",
  17868=>"001001110",
  17869=>"111000010",
  17870=>"100110000",
  17871=>"101110001",
  17872=>"011110011",
  17873=>"101011011",
  17874=>"001001001",
  17875=>"011010000",
  17876=>"111011111",
  17877=>"111001000",
  17878=>"000101101",
  17879=>"010000011",
  17880=>"001000110",
  17881=>"100001101",
  17882=>"101011000",
  17883=>"111100101",
  17884=>"001110111",
  17885=>"001011000",
  17886=>"111110100",
  17887=>"011001011",
  17888=>"111010000",
  17889=>"000100011",
  17890=>"010100000",
  17891=>"111010100",
  17892=>"000001011",
  17893=>"111000010",
  17894=>"111110010",
  17895=>"110110001",
  17896=>"110000100",
  17897=>"011111001",
  17898=>"001001001",
  17899=>"101010110",
  17900=>"011110001",
  17901=>"111010001",
  17902=>"010100010",
  17903=>"100111001",
  17904=>"110101001",
  17905=>"010010001",
  17906=>"111111111",
  17907=>"101010011",
  17908=>"001000111",
  17909=>"010000111",
  17910=>"100110110",
  17911=>"001010001",
  17912=>"010000010",
  17913=>"101000011",
  17914=>"010010001",
  17915=>"000111000",
  17916=>"010011011",
  17917=>"000010110",
  17918=>"110100111",
  17919=>"110001000",
  17920=>"110000101",
  17921=>"001011011",
  17922=>"101001001",
  17923=>"000101011",
  17924=>"010010111",
  17925=>"001011100",
  17926=>"110001110",
  17927=>"011000000",
  17928=>"000010110",
  17929=>"110101010",
  17930=>"100110100",
  17931=>"011001100",
  17932=>"000001110",
  17933=>"000010010",
  17934=>"101110100",
  17935=>"100001011",
  17936=>"001111101",
  17937=>"010101111",
  17938=>"101111010",
  17939=>"011111111",
  17940=>"010010010",
  17941=>"011111011",
  17942=>"000001111",
  17943=>"110111010",
  17944=>"000101001",
  17945=>"000111011",
  17946=>"001110010",
  17947=>"110000011",
  17948=>"000010111",
  17949=>"010101001",
  17950=>"000000010",
  17951=>"110111100",
  17952=>"011011001",
  17953=>"001110000",
  17954=>"001100111",
  17955=>"010111010",
  17956=>"101110001",
  17957=>"111110000",
  17958=>"100000010",
  17959=>"011110101",
  17960=>"110000011",
  17961=>"100010111",
  17962=>"001101100",
  17963=>"001110000",
  17964=>"010000101",
  17965=>"011101010",
  17966=>"101001100",
  17967=>"110001011",
  17968=>"001000001",
  17969=>"011100101",
  17970=>"100000101",
  17971=>"000100111",
  17972=>"001000101",
  17973=>"010000010",
  17974=>"101100101",
  17975=>"010001011",
  17976=>"101010110",
  17977=>"001100010",
  17978=>"111110101",
  17979=>"100011000",
  17980=>"100101111",
  17981=>"001100010",
  17982=>"110001100",
  17983=>"111001111",
  17984=>"001010010",
  17985=>"101010101",
  17986=>"001101101",
  17987=>"001010000",
  17988=>"001101000",
  17989=>"001100000",
  17990=>"011100100",
  17991=>"110111110",
  17992=>"010010011",
  17993=>"000101100",
  17994=>"101100001",
  17995=>"111100000",
  17996=>"110110111",
  17997=>"101100000",
  17998=>"010001100",
  17999=>"011101010",
  18000=>"110111011",
  18001=>"011011100",
  18002=>"010101010",
  18003=>"000101111",
  18004=>"001111000",
  18005=>"010100010",
  18006=>"000001010",
  18007=>"101010011",
  18008=>"101011000",
  18009=>"110010010",
  18010=>"001001011",
  18011=>"010100110",
  18012=>"101100111",
  18013=>"101000000",
  18014=>"110000101",
  18015=>"111010011",
  18016=>"001000011",
  18017=>"010101010",
  18018=>"010100111",
  18019=>"100010001",
  18020=>"001110110",
  18021=>"111101100",
  18022=>"111111101",
  18023=>"111010010",
  18024=>"100100110",
  18025=>"110111001",
  18026=>"011100111",
  18027=>"010011110",
  18028=>"111101010",
  18029=>"000101010",
  18030=>"111011101",
  18031=>"110111111",
  18032=>"001010100",
  18033=>"000101100",
  18034=>"001100111",
  18035=>"110010001",
  18036=>"101111111",
  18037=>"000111001",
  18038=>"100000111",
  18039=>"100110110",
  18040=>"001100000",
  18041=>"111001010",
  18042=>"010001000",
  18043=>"111011111",
  18044=>"110011001",
  18045=>"101010111",
  18046=>"001111010",
  18047=>"111011001",
  18048=>"111111010",
  18049=>"101110000",
  18050=>"101101001",
  18051=>"001100110",
  18052=>"000000011",
  18053=>"011010101",
  18054=>"011111111",
  18055=>"101010000",
  18056=>"111001010",
  18057=>"001000000",
  18058=>"010001101",
  18059=>"111111101",
  18060=>"101011110",
  18061=>"011100100",
  18062=>"011000001",
  18063=>"001000101",
  18064=>"110100010",
  18065=>"010010101",
  18066=>"010011011",
  18067=>"000111111",
  18068=>"111111011",
  18069=>"010110010",
  18070=>"110000110",
  18071=>"000000100",
  18072=>"110011111",
  18073=>"111001001",
  18074=>"101000001",
  18075=>"101010000",
  18076=>"011001100",
  18077=>"110111001",
  18078=>"110001101",
  18079=>"011000001",
  18080=>"100100010",
  18081=>"000111110",
  18082=>"011110100",
  18083=>"011001101",
  18084=>"011111110",
  18085=>"101101001",
  18086=>"111100101",
  18087=>"101000010",
  18088=>"101001011",
  18089=>"010001000",
  18090=>"001011100",
  18091=>"000001000",
  18092=>"100010101",
  18093=>"000000001",
  18094=>"101010000",
  18095=>"000111111",
  18096=>"101011000",
  18097=>"001001001",
  18098=>"011101010",
  18099=>"110010011",
  18100=>"100111001",
  18101=>"000010000",
  18102=>"010010001",
  18103=>"000001110",
  18104=>"000011110",
  18105=>"100000101",
  18106=>"001110100",
  18107=>"000101011",
  18108=>"101100110",
  18109=>"000001001",
  18110=>"000100101",
  18111=>"000000010",
  18112=>"101110000",
  18113=>"011001000",
  18114=>"111011010",
  18115=>"101010111",
  18116=>"000111010",
  18117=>"010010111",
  18118=>"110010010",
  18119=>"011011010",
  18120=>"001001010",
  18121=>"110011001",
  18122=>"100100010",
  18123=>"011100101",
  18124=>"011100110",
  18125=>"110110101",
  18126=>"010010010",
  18127=>"001001100",
  18128=>"001001111",
  18129=>"011111100",
  18130=>"001011000",
  18131=>"111010000",
  18132=>"000100111",
  18133=>"110010100",
  18134=>"100110110",
  18135=>"111001111",
  18136=>"101101100",
  18137=>"010111111",
  18138=>"001001101",
  18139=>"100011001",
  18140=>"100100001",
  18141=>"000000101",
  18142=>"010100010",
  18143=>"110110100",
  18144=>"110011111",
  18145=>"000110100",
  18146=>"001001100",
  18147=>"101111000",
  18148=>"101101111",
  18149=>"011110101",
  18150=>"011101011",
  18151=>"000100111",
  18152=>"101000100",
  18153=>"011110000",
  18154=>"000100111",
  18155=>"010100110",
  18156=>"100001101",
  18157=>"110011101",
  18158=>"101010101",
  18159=>"000011100",
  18160=>"101000100",
  18161=>"010111000",
  18162=>"001011111",
  18163=>"110000101",
  18164=>"101001111",
  18165=>"000110011",
  18166=>"011111100",
  18167=>"011101100",
  18168=>"001010001",
  18169=>"111110000",
  18170=>"100110000",
  18171=>"010001000",
  18172=>"010010100",
  18173=>"010011010",
  18174=>"001000001",
  18175=>"110110001",
  18176=>"010011100",
  18177=>"100010100",
  18178=>"001101001",
  18179=>"101011101",
  18180=>"001101101",
  18181=>"110000001",
  18182=>"100111000",
  18183=>"111000110",
  18184=>"101101111",
  18185=>"100111111",
  18186=>"111110110",
  18187=>"000000101",
  18188=>"010100000",
  18189=>"101111011",
  18190=>"111111101",
  18191=>"110101011",
  18192=>"101101111",
  18193=>"011000101",
  18194=>"101001101",
  18195=>"111011111",
  18196=>"101110011",
  18197=>"001010011",
  18198=>"000010111",
  18199=>"110100001",
  18200=>"000111101",
  18201=>"010110000",
  18202=>"010011011",
  18203=>"111100001",
  18204=>"010111011",
  18205=>"111111100",
  18206=>"101010110",
  18207=>"010110010",
  18208=>"111001001",
  18209=>"101011001",
  18210=>"100000101",
  18211=>"100010000",
  18212=>"100000000",
  18213=>"100101001",
  18214=>"010110010",
  18215=>"001010101",
  18216=>"110101100",
  18217=>"000001001",
  18218=>"101101101",
  18219=>"110011101",
  18220=>"100110111",
  18221=>"101000011",
  18222=>"001101000",
  18223=>"101111101",
  18224=>"100011001",
  18225=>"001000000",
  18226=>"111001101",
  18227=>"101001011",
  18228=>"101111110",
  18229=>"110111110",
  18230=>"010101100",
  18231=>"000100111",
  18232=>"111101100",
  18233=>"101011000",
  18234=>"010000110",
  18235=>"010101110",
  18236=>"011001010",
  18237=>"100100100",
  18238=>"010011011",
  18239=>"001011000",
  18240=>"101100011",
  18241=>"010110101",
  18242=>"111111001",
  18243=>"101100100",
  18244=>"100000010",
  18245=>"110001111",
  18246=>"001110110",
  18247=>"100011001",
  18248=>"101101100",
  18249=>"111001011",
  18250=>"001000100",
  18251=>"100101011",
  18252=>"111001111",
  18253=>"101100110",
  18254=>"110101011",
  18255=>"101001100",
  18256=>"000000110",
  18257=>"100001011",
  18258=>"001011001",
  18259=>"111110110",
  18260=>"011110110",
  18261=>"010010101",
  18262=>"100101111",
  18263=>"010010001",
  18264=>"111000010",
  18265=>"100101111",
  18266=>"101010101",
  18267=>"110111010",
  18268=>"000111101",
  18269=>"100011100",
  18270=>"011110000",
  18271=>"110100010",
  18272=>"011011111",
  18273=>"010010100",
  18274=>"001000111",
  18275=>"011101000",
  18276=>"011111000",
  18277=>"011000110",
  18278=>"001101011",
  18279=>"001001001",
  18280=>"111011111",
  18281=>"110110011",
  18282=>"101000001",
  18283=>"011100000",
  18284=>"100111101",
  18285=>"000001011",
  18286=>"100001001",
  18287=>"100111000",
  18288=>"010101111",
  18289=>"101111111",
  18290=>"001010111",
  18291=>"011101100",
  18292=>"101101001",
  18293=>"111100110",
  18294=>"011111101",
  18295=>"101100000",
  18296=>"010111111",
  18297=>"001000000",
  18298=>"100111001",
  18299=>"101011101",
  18300=>"001010101",
  18301=>"100000111",
  18302=>"011000010",
  18303=>"011011011",
  18304=>"101001011",
  18305=>"111000001",
  18306=>"111110101",
  18307=>"000110000",
  18308=>"011001101",
  18309=>"000111000",
  18310=>"010001111",
  18311=>"000101111",
  18312=>"001000101",
  18313=>"010100010",
  18314=>"010010001",
  18315=>"101111100",
  18316=>"110100100",
  18317=>"000011011",
  18318=>"010010111",
  18319=>"100101010",
  18320=>"000111110",
  18321=>"101000011",
  18322=>"010000110",
  18323=>"100101010",
  18324=>"110100001",
  18325=>"110100110",
  18326=>"010100001",
  18327=>"101000000",
  18328=>"001000111",
  18329=>"111101001",
  18330=>"000110011",
  18331=>"001110011",
  18332=>"100100100",
  18333=>"000000000",
  18334=>"010000110",
  18335=>"000101011",
  18336=>"011101110",
  18337=>"001010010",
  18338=>"110110100",
  18339=>"000111100",
  18340=>"001100001",
  18341=>"000111110",
  18342=>"001000001",
  18343=>"010000010",
  18344=>"001010010",
  18345=>"101001110",
  18346=>"101111101",
  18347=>"001010011",
  18348=>"000011110",
  18349=>"110101110",
  18350=>"010011101",
  18351=>"000110010",
  18352=>"010101001",
  18353=>"111010010",
  18354=>"011111011",
  18355=>"000110111",
  18356=>"111111011",
  18357=>"100110000",
  18358=>"000011111",
  18359=>"110000010",
  18360=>"100010110",
  18361=>"000111011",
  18362=>"100011100",
  18363=>"100100100",
  18364=>"000011100",
  18365=>"101010100",
  18366=>"110111111",
  18367=>"010110101",
  18368=>"011000011",
  18369=>"000010101",
  18370=>"101010001",
  18371=>"100000010",
  18372=>"000001000",
  18373=>"111110010",
  18374=>"111011110",
  18375=>"101000010",
  18376=>"001001010",
  18377=>"101111000",
  18378=>"010000001",
  18379=>"011101011",
  18380=>"011011101",
  18381=>"111100000",
  18382=>"011011111",
  18383=>"101110110",
  18384=>"111010110",
  18385=>"011000010",
  18386=>"111110001",
  18387=>"100110010",
  18388=>"010111100",
  18389=>"101000001",
  18390=>"000110111",
  18391=>"001000100",
  18392=>"111110111",
  18393=>"111100110",
  18394=>"111111111",
  18395=>"001011010",
  18396=>"100000011",
  18397=>"011000000",
  18398=>"001101101",
  18399=>"111001111",
  18400=>"011101010",
  18401=>"101101100",
  18402=>"100011100",
  18403=>"111110010",
  18404=>"100011110",
  18405=>"101101011",
  18406=>"100101001",
  18407=>"111011101",
  18408=>"101110111",
  18409=>"000001011",
  18410=>"010000110",
  18411=>"110100110",
  18412=>"000110100",
  18413=>"010101000",
  18414=>"001010101",
  18415=>"000101111",
  18416=>"101111010",
  18417=>"101100111",
  18418=>"000110000",
  18419=>"010000000",
  18420=>"011110010",
  18421=>"010011011",
  18422=>"001001011",
  18423=>"110100101",
  18424=>"100011101",
  18425=>"010100101",
  18426=>"111000100",
  18427=>"101111101",
  18428=>"000011111",
  18429=>"010101010",
  18430=>"111101011",
  18431=>"011000000",
  18432=>"011111010",
  18433=>"100011110",
  18434=>"101000110",
  18435=>"010000000",
  18436=>"101101101",
  18437=>"100110011",
  18438=>"010000100",
  18439=>"100100101",
  18440=>"111001101",
  18441=>"110000101",
  18442=>"111000100",
  18443=>"000110101",
  18444=>"111010100",
  18445=>"010011101",
  18446=>"010100111",
  18447=>"110101111",
  18448=>"100000010",
  18449=>"010111101",
  18450=>"011011000",
  18451=>"111011100",
  18452=>"111101100",
  18453=>"110100101",
  18454=>"000100001",
  18455=>"011000000",
  18456=>"101000111",
  18457=>"111100011",
  18458=>"011110101",
  18459=>"001100000",
  18460=>"100001111",
  18461=>"011100010",
  18462=>"010011000",
  18463=>"001011111",
  18464=>"011011111",
  18465=>"011010101",
  18466=>"111111001",
  18467=>"111111000",
  18468=>"011110110",
  18469=>"111111111",
  18470=>"011010100",
  18471=>"010100111",
  18472=>"101001110",
  18473=>"011011110",
  18474=>"110010110",
  18475=>"111110111",
  18476=>"100001001",
  18477=>"001101100",
  18478=>"111111111",
  18479=>"101100111",
  18480=>"101101111",
  18481=>"100001110",
  18482=>"100011001",
  18483=>"111011001",
  18484=>"111110010",
  18485=>"111001000",
  18486=>"000001100",
  18487=>"001000001",
  18488=>"001000000",
  18489=>"010100000",
  18490=>"101010101",
  18491=>"100011101",
  18492=>"100000000",
  18493=>"101001011",
  18494=>"001100010",
  18495=>"010110001",
  18496=>"011000110",
  18497=>"001000100",
  18498=>"010000011",
  18499=>"101100001",
  18500=>"101111110",
  18501=>"100010100",
  18502=>"011011101",
  18503=>"011010111",
  18504=>"000111000",
  18505=>"110000110",
  18506=>"010111111",
  18507=>"110000010",
  18508=>"111011110",
  18509=>"001010000",
  18510=>"000011001",
  18511=>"111111010",
  18512=>"111010111",
  18513=>"000110100",
  18514=>"111110001",
  18515=>"101100001",
  18516=>"100101100",
  18517=>"010010100",
  18518=>"100101010",
  18519=>"010001100",
  18520=>"111100100",
  18521=>"001000100",
  18522=>"110111000",
  18523=>"010100000",
  18524=>"100001100",
  18525=>"110100010",
  18526=>"101011000",
  18527=>"110100001",
  18528=>"000111010",
  18529=>"110011110",
  18530=>"000110011",
  18531=>"000110110",
  18532=>"111111000",
  18533=>"111100001",
  18534=>"111011101",
  18535=>"100010111",
  18536=>"010110000",
  18537=>"111000101",
  18538=>"111001101",
  18539=>"101100101",
  18540=>"010000010",
  18541=>"000000110",
  18542=>"111110001",
  18543=>"011010101",
  18544=>"100110111",
  18545=>"000001100",
  18546=>"101010001",
  18547=>"101000101",
  18548=>"110010111",
  18549=>"010111001",
  18550=>"101101111",
  18551=>"100100011",
  18552=>"000000011",
  18553=>"101000010",
  18554=>"101100011",
  18555=>"010100011",
  18556=>"001101010",
  18557=>"111110100",
  18558=>"001101100",
  18559=>"000110000",
  18560=>"011010111",
  18561=>"000001000",
  18562=>"010101110",
  18563=>"000001001",
  18564=>"101001100",
  18565=>"011100110",
  18566=>"110111011",
  18567=>"001110000",
  18568=>"110101011",
  18569=>"111010001",
  18570=>"111011010",
  18571=>"001111110",
  18572=>"110100011",
  18573=>"100011101",
  18574=>"100001011",
  18575=>"010010101",
  18576=>"111001101",
  18577=>"101101100",
  18578=>"110011100",
  18579=>"101001011",
  18580=>"101011000",
  18581=>"101100101",
  18582=>"100111110",
  18583=>"001001111",
  18584=>"111100100",
  18585=>"111101101",
  18586=>"000101011",
  18587=>"011000100",
  18588=>"011011101",
  18589=>"000011000",
  18590=>"111111111",
  18591=>"110010101",
  18592=>"110000110",
  18593=>"111110000",
  18594=>"111111011",
  18595=>"110000111",
  18596=>"010110001",
  18597=>"010010001",
  18598=>"011000011",
  18599=>"000111001",
  18600=>"011011101",
  18601=>"000011110",
  18602=>"001101100",
  18603=>"001100100",
  18604=>"111000000",
  18605=>"010010001",
  18606=>"111001110",
  18607=>"011011001",
  18608=>"001000110",
  18609=>"001110010",
  18610=>"010011001",
  18611=>"000011100",
  18612=>"101000111",
  18613=>"101110100",
  18614=>"101111011",
  18615=>"000000000",
  18616=>"000000101",
  18617=>"001001000",
  18618=>"010110100",
  18619=>"000011010",
  18620=>"110110101",
  18621=>"101001000",
  18622=>"000101011",
  18623=>"010011001",
  18624=>"010000011",
  18625=>"111001110",
  18626=>"001000000",
  18627=>"010000011",
  18628=>"110001011",
  18629=>"001000101",
  18630=>"010000100",
  18631=>"011101110",
  18632=>"101110011",
  18633=>"101110001",
  18634=>"010011010",
  18635=>"011000010",
  18636=>"100001110",
  18637=>"011110100",
  18638=>"111100011",
  18639=>"101010010",
  18640=>"100011011",
  18641=>"000101110",
  18642=>"000000001",
  18643=>"011110100",
  18644=>"101010000",
  18645=>"011000010",
  18646=>"001000011",
  18647=>"001001010",
  18648=>"000000000",
  18649=>"011101010",
  18650=>"110001011",
  18651=>"010010010",
  18652=>"100101100",
  18653=>"000100100",
  18654=>"010010000",
  18655=>"110000001",
  18656=>"111100110",
  18657=>"001101000",
  18658=>"011110001",
  18659=>"111010000",
  18660=>"110010100",
  18661=>"111100111",
  18662=>"101000000",
  18663=>"101000000",
  18664=>"000100100",
  18665=>"111101110",
  18666=>"010000010",
  18667=>"101111000",
  18668=>"101000111",
  18669=>"010000111",
  18670=>"001111010",
  18671=>"000010100",
  18672=>"010101010",
  18673=>"101111000",
  18674=>"110000110",
  18675=>"000011100",
  18676=>"111110000",
  18677=>"111001111",
  18678=>"111110101",
  18679=>"110000010",
  18680=>"000111000",
  18681=>"111011010",
  18682=>"100101010",
  18683=>"110110001",
  18684=>"110100111",
  18685=>"000111100",
  18686=>"111011011",
  18687=>"010011110",
  18688=>"001010001",
  18689=>"100100110",
  18690=>"110111100",
  18691=>"110100100",
  18692=>"101101100",
  18693=>"011010110",
  18694=>"100000000",
  18695=>"010011000",
  18696=>"100101111",
  18697=>"100001101",
  18698=>"111101011",
  18699=>"011001000",
  18700=>"001100101",
  18701=>"011011011",
  18702=>"110010011",
  18703=>"000000000",
  18704=>"001011110",
  18705=>"010001011",
  18706=>"101001110",
  18707=>"001111110",
  18708=>"110011011",
  18709=>"100100010",
  18710=>"011111000",
  18711=>"000011011",
  18712=>"011111000",
  18713=>"101110101",
  18714=>"100000001",
  18715=>"100001100",
  18716=>"111100110",
  18717=>"100010000",
  18718=>"101001000",
  18719=>"010110010",
  18720=>"111000000",
  18721=>"010100000",
  18722=>"111011111",
  18723=>"111010010",
  18724=>"001010011",
  18725=>"101000000",
  18726=>"111101101",
  18727=>"001111000",
  18728=>"000000110",
  18729=>"011100111",
  18730=>"110000010",
  18731=>"100001000",
  18732=>"111000000",
  18733=>"101010000",
  18734=>"111101000",
  18735=>"111110110",
  18736=>"010000100",
  18737=>"111101100",
  18738=>"001000000",
  18739=>"001100010",
  18740=>"101100111",
  18741=>"110101110",
  18742=>"001111001",
  18743=>"101011010",
  18744=>"100011101",
  18745=>"100101000",
  18746=>"111111101",
  18747=>"111100110",
  18748=>"000000100",
  18749=>"011110000",
  18750=>"110101111",
  18751=>"111100001",
  18752=>"101100011",
  18753=>"111111001",
  18754=>"101010110",
  18755=>"001010010",
  18756=>"100000000",
  18757=>"111111011",
  18758=>"110011101",
  18759=>"011101111",
  18760=>"010001100",
  18761=>"110001001",
  18762=>"101001110",
  18763=>"111000101",
  18764=>"000101000",
  18765=>"011101101",
  18766=>"001011101",
  18767=>"000111011",
  18768=>"110111001",
  18769=>"110100110",
  18770=>"111111110",
  18771=>"001100100",
  18772=>"010110100",
  18773=>"001010101",
  18774=>"000101010",
  18775=>"110110011",
  18776=>"010011001",
  18777=>"011000010",
  18778=>"000001111",
  18779=>"111000000",
  18780=>"010110110",
  18781=>"110010001",
  18782=>"011100010",
  18783=>"100010001",
  18784=>"000100100",
  18785=>"000010110",
  18786=>"001101101",
  18787=>"100010111",
  18788=>"010001100",
  18789=>"100000110",
  18790=>"011110100",
  18791=>"011100100",
  18792=>"001101110",
  18793=>"011100001",
  18794=>"110101100",
  18795=>"000001101",
  18796=>"100100000",
  18797=>"001001001",
  18798=>"011001100",
  18799=>"011010100",
  18800=>"100001100",
  18801=>"100000110",
  18802=>"100010001",
  18803=>"010101011",
  18804=>"000001100",
  18805=>"101110001",
  18806=>"101110001",
  18807=>"110011001",
  18808=>"100000100",
  18809=>"100000011",
  18810=>"110011101",
  18811=>"001000100",
  18812=>"000000110",
  18813=>"010110011",
  18814=>"111111001",
  18815=>"100100011",
  18816=>"010110111",
  18817=>"011101011",
  18818=>"100101001",
  18819=>"100001111",
  18820=>"111010111",
  18821=>"101111011",
  18822=>"111010111",
  18823=>"101010001",
  18824=>"001001110",
  18825=>"010000010",
  18826=>"001101001",
  18827=>"000011101",
  18828=>"101010111",
  18829=>"011000000",
  18830=>"101010110",
  18831=>"110000101",
  18832=>"000001111",
  18833=>"111000111",
  18834=>"011000110",
  18835=>"001111011",
  18836=>"110101110",
  18837=>"100111011",
  18838=>"111100000",
  18839=>"101000110",
  18840=>"100000010",
  18841=>"101100001",
  18842=>"110111110",
  18843=>"110011010",
  18844=>"101110111",
  18845=>"011000001",
  18846=>"011100111",
  18847=>"101101111",
  18848=>"111011010",
  18849=>"100111001",
  18850=>"010000001",
  18851=>"110001010",
  18852=>"000011100",
  18853=>"110010001",
  18854=>"100101110",
  18855=>"110010100",
  18856=>"110110011",
  18857=>"100111101",
  18858=>"100100110",
  18859=>"001010110",
  18860=>"101111011",
  18861=>"100011111",
  18862=>"010010100",
  18863=>"010010110",
  18864=>"000111101",
  18865=>"011111100",
  18866=>"011101100",
  18867=>"110110000",
  18868=>"000010101",
  18869=>"001101011",
  18870=>"000100100",
  18871=>"011010110",
  18872=>"111101001",
  18873=>"011110000",
  18874=>"000100010",
  18875=>"100001100",
  18876=>"110011100",
  18877=>"111001111",
  18878=>"001101101",
  18879=>"111100101",
  18880=>"101100000",
  18881=>"110101111",
  18882=>"000101111",
  18883=>"110110010",
  18884=>"010000100",
  18885=>"000011001",
  18886=>"000101111",
  18887=>"011000000",
  18888=>"011110001",
  18889=>"000111111",
  18890=>"001000000",
  18891=>"100111010",
  18892=>"110110011",
  18893=>"010100101",
  18894=>"010001100",
  18895=>"110001101",
  18896=>"100110110",
  18897=>"100100011",
  18898=>"100001000",
  18899=>"000111000",
  18900=>"011111001",
  18901=>"100000000",
  18902=>"111111011",
  18903=>"111001011",
  18904=>"000111111",
  18905=>"101000100",
  18906=>"001001011",
  18907=>"111111110",
  18908=>"000000000",
  18909=>"101000000",
  18910=>"010011001",
  18911=>"000111111",
  18912=>"111011100",
  18913=>"000000111",
  18914=>"101101011",
  18915=>"010000000",
  18916=>"000100111",
  18917=>"101111001",
  18918=>"001001101",
  18919=>"111111101",
  18920=>"001000101",
  18921=>"100110000",
  18922=>"001111000",
  18923=>"111101101",
  18924=>"111000010",
  18925=>"111101000",
  18926=>"010000000",
  18927=>"111000011",
  18928=>"101101110",
  18929=>"100101011",
  18930=>"010111100",
  18931=>"001110000",
  18932=>"100000011",
  18933=>"010000001",
  18934=>"110101111",
  18935=>"000101101",
  18936=>"010110010",
  18937=>"111101101",
  18938=>"000101111",
  18939=>"010111010",
  18940=>"001111010",
  18941=>"001001100",
  18942=>"100101011",
  18943=>"001001011",
  18944=>"001011100",
  18945=>"100010011",
  18946=>"101101011",
  18947=>"011100011",
  18948=>"100000101",
  18949=>"100101010",
  18950=>"001001111",
  18951=>"100111111",
  18952=>"010111000",
  18953=>"010010010",
  18954=>"010010000",
  18955=>"000000000",
  18956=>"000011010",
  18957=>"000000000",
  18958=>"010001100",
  18959=>"000011000",
  18960=>"110110101",
  18961=>"110110000",
  18962=>"100110011",
  18963=>"010111110",
  18964=>"010000000",
  18965=>"010101010",
  18966=>"100001011",
  18967=>"110000100",
  18968=>"000010110",
  18969=>"000110011",
  18970=>"101000101",
  18971=>"111010100",
  18972=>"011000101",
  18973=>"000101111",
  18974=>"011111011",
  18975=>"111111100",
  18976=>"111101111",
  18977=>"110011000",
  18978=>"110000001",
  18979=>"000010100",
  18980=>"001111100",
  18981=>"101001111",
  18982=>"000011000",
  18983=>"010000010",
  18984=>"110010001",
  18985=>"101001111",
  18986=>"011101101",
  18987=>"011010110",
  18988=>"110011101",
  18989=>"110000010",
  18990=>"110000001",
  18991=>"101110000",
  18992=>"100000010",
  18993=>"110111001",
  18994=>"100000110",
  18995=>"011100011",
  18996=>"100000010",
  18997=>"010100010",
  18998=>"010101110",
  18999=>"000111001",
  19000=>"000100001",
  19001=>"000000100",
  19002=>"110110010",
  19003=>"110000010",
  19004=>"100100000",
  19005=>"111100000",
  19006=>"101011001",
  19007=>"111111011",
  19008=>"010000110",
  19009=>"000000000",
  19010=>"100000011",
  19011=>"010101011",
  19012=>"000000111",
  19013=>"101001011",
  19014=>"000000011",
  19015=>"110111001",
  19016=>"110011111",
  19017=>"101010110",
  19018=>"010111011",
  19019=>"111000100",
  19020=>"011001111",
  19021=>"010110110",
  19022=>"011000100",
  19023=>"001000001",
  19024=>"000010101",
  19025=>"010000101",
  19026=>"000100111",
  19027=>"010111100",
  19028=>"001000101",
  19029=>"001001100",
  19030=>"011110010",
  19031=>"110011100",
  19032=>"011111110",
  19033=>"100100101",
  19034=>"101100000",
  19035=>"010111011",
  19036=>"010011011",
  19037=>"010010011",
  19038=>"011001111",
  19039=>"010011010",
  19040=>"111001110",
  19041=>"010110000",
  19042=>"011011110",
  19043=>"001111010",
  19044=>"001001101",
  19045=>"001101110",
  19046=>"000000011",
  19047=>"001001011",
  19048=>"110110111",
  19049=>"000111111",
  19050=>"101101010",
  19051=>"011110110",
  19052=>"101100111",
  19053=>"001011110",
  19054=>"111010110",
  19055=>"001111100",
  19056=>"100100010",
  19057=>"111001100",
  19058=>"010101001",
  19059=>"111111100",
  19060=>"011000001",
  19061=>"101010000",
  19062=>"010100111",
  19063=>"010110101",
  19064=>"100101000",
  19065=>"111010010",
  19066=>"101110110",
  19067=>"100101001",
  19068=>"101100000",
  19069=>"110000110",
  19070=>"000000111",
  19071=>"010000000",
  19072=>"111011001",
  19073=>"101011001",
  19074=>"011100001",
  19075=>"000100100",
  19076=>"010001110",
  19077=>"100100000",
  19078=>"111100101",
  19079=>"111011100",
  19080=>"011111000",
  19081=>"111101101",
  19082=>"011110110",
  19083=>"110110111",
  19084=>"100011010",
  19085=>"100110100",
  19086=>"100011100",
  19087=>"110100011",
  19088=>"110011100",
  19089=>"000000011",
  19090=>"010111100",
  19091=>"101101110",
  19092=>"000001010",
  19093=>"100111100",
  19094=>"111010100",
  19095=>"111100101",
  19096=>"101110110",
  19097=>"101101000",
  19098=>"101010101",
  19099=>"000010110",
  19100=>"111000000",
  19101=>"110011110",
  19102=>"001111110",
  19103=>"100011100",
  19104=>"100011110",
  19105=>"111110001",
  19106=>"000110110",
  19107=>"110111010",
  19108=>"100001100",
  19109=>"110110110",
  19110=>"011000101",
  19111=>"001100110",
  19112=>"101100010",
  19113=>"010111000",
  19114=>"000010011",
  19115=>"011111110",
  19116=>"111011001",
  19117=>"101110000",
  19118=>"101100001",
  19119=>"100100101",
  19120=>"000001001",
  19121=>"001101100",
  19122=>"000001101",
  19123=>"100101001",
  19124=>"010100011",
  19125=>"111110000",
  19126=>"101111000",
  19127=>"100100100",
  19128=>"010001001",
  19129=>"101101001",
  19130=>"000001100",
  19131=>"001011011",
  19132=>"000110101",
  19133=>"100000101",
  19134=>"000100010",
  19135=>"101100011",
  19136=>"000000110",
  19137=>"001110000",
  19138=>"010010011",
  19139=>"110001110",
  19140=>"100001000",
  19141=>"100101101",
  19142=>"010001100",
  19143=>"011111000",
  19144=>"001111111",
  19145=>"101011001",
  19146=>"011001110",
  19147=>"100111010",
  19148=>"011100011",
  19149=>"111001001",
  19150=>"011110011",
  19151=>"111010110",
  19152=>"111111001",
  19153=>"011011000",
  19154=>"000001101",
  19155=>"110000101",
  19156=>"110010010",
  19157=>"101011010",
  19158=>"011000001",
  19159=>"100001111",
  19160=>"101111010",
  19161=>"000001110",
  19162=>"011010000",
  19163=>"010100000",
  19164=>"100100111",
  19165=>"110111000",
  19166=>"001100101",
  19167=>"001010011",
  19168=>"111001000",
  19169=>"011110001",
  19170=>"101001011",
  19171=>"001001000",
  19172=>"110000110",
  19173=>"010110101",
  19174=>"000011101",
  19175=>"000010000",
  19176=>"001001101",
  19177=>"111111101",
  19178=>"011001111",
  19179=>"101100100",
  19180=>"010010101",
  19181=>"100011100",
  19182=>"111111110",
  19183=>"100000100",
  19184=>"110111110",
  19185=>"110110111",
  19186=>"000111001",
  19187=>"110110011",
  19188=>"101110001",
  19189=>"011001101",
  19190=>"101000001",
  19191=>"011101000",
  19192=>"100000011",
  19193=>"111000100",
  19194=>"111110010",
  19195=>"000010100",
  19196=>"110000000",
  19197=>"001110000",
  19198=>"010001111",
  19199=>"111111110",
  19200=>"001001110",
  19201=>"111011011",
  19202=>"010111000",
  19203=>"100010100",
  19204=>"000101101",
  19205=>"000000000",
  19206=>"100001011",
  19207=>"000001111",
  19208=>"001010111",
  19209=>"000000101",
  19210=>"101111000",
  19211=>"010011000",
  19212=>"110011011",
  19213=>"101000101",
  19214=>"111010010",
  19215=>"110001000",
  19216=>"111100001",
  19217=>"001100101",
  19218=>"101010001",
  19219=>"111000011",
  19220=>"011100101",
  19221=>"110110010",
  19222=>"111011110",
  19223=>"010100100",
  19224=>"010011010",
  19225=>"001011110",
  19226=>"110011010",
  19227=>"110111001",
  19228=>"000000010",
  19229=>"111011001",
  19230=>"000001000",
  19231=>"000100011",
  19232=>"111110100",
  19233=>"000001110",
  19234=>"000100101",
  19235=>"011101101",
  19236=>"110000000",
  19237=>"011001010",
  19238=>"110111110",
  19239=>"100110101",
  19240=>"010010000",
  19241=>"000010010",
  19242=>"110111001",
  19243=>"001000011",
  19244=>"010110100",
  19245=>"000000111",
  19246=>"110010111",
  19247=>"100110011",
  19248=>"000100001",
  19249=>"001011010",
  19250=>"000110011",
  19251=>"010001000",
  19252=>"101111001",
  19253=>"000010001",
  19254=>"111010111",
  19255=>"101110100",
  19256=>"000010110",
  19257=>"100100100",
  19258=>"100110010",
  19259=>"100111010",
  19260=>"100101001",
  19261=>"110111000",
  19262=>"111100101",
  19263=>"101010100",
  19264=>"010000001",
  19265=>"111000100",
  19266=>"001101100",
  19267=>"110011110",
  19268=>"101001001",
  19269=>"000000101",
  19270=>"011000010",
  19271=>"101011000",
  19272=>"110001100",
  19273=>"010110111",
  19274=>"010010101",
  19275=>"100111010",
  19276=>"100100001",
  19277=>"001010101",
  19278=>"010000000",
  19279=>"001001000",
  19280=>"111011101",
  19281=>"010000001",
  19282=>"010110011",
  19283=>"100111001",
  19284=>"001101011",
  19285=>"110101111",
  19286=>"111011000",
  19287=>"010111110",
  19288=>"011010110",
  19289=>"000011100",
  19290=>"011110010",
  19291=>"000000111",
  19292=>"001111011",
  19293=>"111111110",
  19294=>"100100011",
  19295=>"011111001",
  19296=>"010100101",
  19297=>"001111111",
  19298=>"100101000",
  19299=>"011111010",
  19300=>"000011100",
  19301=>"011010100",
  19302=>"111100110",
  19303=>"001100011",
  19304=>"101110100",
  19305=>"010100000",
  19306=>"100100110",
  19307=>"011100110",
  19308=>"010010100",
  19309=>"111001000",
  19310=>"010010111",
  19311=>"100010010",
  19312=>"011100101",
  19313=>"001100101",
  19314=>"011010111",
  19315=>"101110110",
  19316=>"100110110",
  19317=>"010010010",
  19318=>"111010101",
  19319=>"110011011",
  19320=>"101100101",
  19321=>"111100111",
  19322=>"000000101",
  19323=>"110111011",
  19324=>"000000000",
  19325=>"110101101",
  19326=>"100101011",
  19327=>"100111011",
  19328=>"011111010",
  19329=>"101101101",
  19330=>"101000101",
  19331=>"000011101",
  19332=>"010101001",
  19333=>"000011100",
  19334=>"101001000",
  19335=>"100111101",
  19336=>"000000111",
  19337=>"000100001",
  19338=>"000110100",
  19339=>"000011010",
  19340=>"001010011",
  19341=>"101110100",
  19342=>"110101000",
  19343=>"110001000",
  19344=>"111010001",
  19345=>"100110110",
  19346=>"011010111",
  19347=>"010001011",
  19348=>"000011010",
  19349=>"010111101",
  19350=>"011101000",
  19351=>"011111101",
  19352=>"010110011",
  19353=>"111111011",
  19354=>"010011011",
  19355=>"110001111",
  19356=>"100011011",
  19357=>"100100000",
  19358=>"101100100",
  19359=>"000010000",
  19360=>"000110000",
  19361=>"001100001",
  19362=>"101010111",
  19363=>"001101101",
  19364=>"101010111",
  19365=>"111100011",
  19366=>"011111110",
  19367=>"100010000",
  19368=>"110010001",
  19369=>"011000000",
  19370=>"001001100",
  19371=>"110000110",
  19372=>"100101011",
  19373=>"110011001",
  19374=>"010110011",
  19375=>"000101110",
  19376=>"110110010",
  19377=>"100100111",
  19378=>"010001111",
  19379=>"101001010",
  19380=>"011111100",
  19381=>"110100000",
  19382=>"110010101",
  19383=>"100010101",
  19384=>"100100011",
  19385=>"011101110",
  19386=>"011110011",
  19387=>"010000000",
  19388=>"000111000",
  19389=>"111001111",
  19390=>"100111010",
  19391=>"111110111",
  19392=>"001001100",
  19393=>"011010111",
  19394=>"010100100",
  19395=>"101110100",
  19396=>"111110101",
  19397=>"010001000",
  19398=>"100110101",
  19399=>"000110001",
  19400=>"110001010",
  19401=>"010001000",
  19402=>"000010000",
  19403=>"010010011",
  19404=>"000000011",
  19405=>"100001000",
  19406=>"111100001",
  19407=>"101011100",
  19408=>"111000111",
  19409=>"010001100",
  19410=>"000011101",
  19411=>"101110101",
  19412=>"010111000",
  19413=>"001001001",
  19414=>"000100101",
  19415=>"010100011",
  19416=>"100000100",
  19417=>"011010010",
  19418=>"011000101",
  19419=>"100010101",
  19420=>"110101111",
  19421=>"111000110",
  19422=>"001001110",
  19423=>"011011100",
  19424=>"001000111",
  19425=>"000111001",
  19426=>"110000001",
  19427=>"111110110",
  19428=>"011010000",
  19429=>"010000110",
  19430=>"110110011",
  19431=>"101100001",
  19432=>"110011010",
  19433=>"101101010",
  19434=>"011001110",
  19435=>"001100001",
  19436=>"011001011",
  19437=>"100000101",
  19438=>"000101000",
  19439=>"101100011",
  19440=>"010001001",
  19441=>"100010110",
  19442=>"100101011",
  19443=>"101000000",
  19444=>"010010010",
  19445=>"011101011",
  19446=>"101110010",
  19447=>"110011011",
  19448=>"010000000",
  19449=>"000010011",
  19450=>"010101100",
  19451=>"111101111",
  19452=>"100000010",
  19453=>"011001011",
  19454=>"010001011",
  19455=>"010010011",
  19456=>"001010111",
  19457=>"000000011",
  19458=>"001001101",
  19459=>"111111110",
  19460=>"111110011",
  19461=>"000011011",
  19462=>"000100110",
  19463=>"111011010",
  19464=>"001100011",
  19465=>"000001110",
  19466=>"011011010",
  19467=>"000000011",
  19468=>"001011000",
  19469=>"011111101",
  19470=>"101111111",
  19471=>"010001000",
  19472=>"011000010",
  19473=>"010110000",
  19474=>"110101011",
  19475=>"111011101",
  19476=>"100100101",
  19477=>"001111111",
  19478=>"100001011",
  19479=>"101000100",
  19480=>"001001001",
  19481=>"010001011",
  19482=>"010111100",
  19483=>"000101101",
  19484=>"110110111",
  19485=>"000000101",
  19486=>"101100001",
  19487=>"111100010",
  19488=>"000110111",
  19489=>"101101100",
  19490=>"110000101",
  19491=>"100001111",
  19492=>"111100010",
  19493=>"000111011",
  19494=>"011111010",
  19495=>"000000000",
  19496=>"011000010",
  19497=>"010101000",
  19498=>"111110111",
  19499=>"011110110",
  19500=>"110010111",
  19501=>"010101001",
  19502=>"011100111",
  19503=>"011111110",
  19504=>"110010111",
  19505=>"111110010",
  19506=>"010111110",
  19507=>"101101101",
  19508=>"000011011",
  19509=>"011000100",
  19510=>"111101011",
  19511=>"110010100",
  19512=>"011011101",
  19513=>"110000110",
  19514=>"011000110",
  19515=>"000001100",
  19516=>"001001101",
  19517=>"010001010",
  19518=>"101100011",
  19519=>"010111000",
  19520=>"100000111",
  19521=>"000010011",
  19522=>"000100011",
  19523=>"101100010",
  19524=>"101010001",
  19525=>"111101000",
  19526=>"001000001",
  19527=>"000001001",
  19528=>"000001111",
  19529=>"010000000",
  19530=>"100001111",
  19531=>"001011010",
  19532=>"001011000",
  19533=>"111111010",
  19534=>"101111100",
  19535=>"011010010",
  19536=>"010000101",
  19537=>"111001101",
  19538=>"011101111",
  19539=>"010000111",
  19540=>"101000101",
  19541=>"110011110",
  19542=>"101011111",
  19543=>"010011000",
  19544=>"111110111",
  19545=>"001101001",
  19546=>"111100010",
  19547=>"100000111",
  19548=>"101101101",
  19549=>"000101110",
  19550=>"110010011",
  19551=>"110000111",
  19552=>"101110100",
  19553=>"011011011",
  19554=>"100010000",
  19555=>"001010000",
  19556=>"101101101",
  19557=>"000001111",
  19558=>"011010110",
  19559=>"000000010",
  19560=>"110001100",
  19561=>"110011001",
  19562=>"000001011",
  19563=>"001010100",
  19564=>"011000000",
  19565=>"110000111",
  19566=>"010010000",
  19567=>"110000111",
  19568=>"111000000",
  19569=>"100001111",
  19570=>"111001110",
  19571=>"110001010",
  19572=>"000111110",
  19573=>"011001111",
  19574=>"101110000",
  19575=>"101101000",
  19576=>"001010111",
  19577=>"000000101",
  19578=>"100001110",
  19579=>"101011110",
  19580=>"110001000",
  19581=>"000010011",
  19582=>"010000001",
  19583=>"011110100",
  19584=>"111001010",
  19585=>"001001110",
  19586=>"000000010",
  19587=>"010110011",
  19588=>"000101010",
  19589=>"010010010",
  19590=>"111010000",
  19591=>"111110111",
  19592=>"101110111",
  19593=>"001110010",
  19594=>"000000010",
  19595=>"111001100",
  19596=>"001101101",
  19597=>"101100011",
  19598=>"001110001",
  19599=>"001110011",
  19600=>"001000100",
  19601=>"101010100",
  19602=>"111111000",
  19603=>"111010101",
  19604=>"100011111",
  19605=>"001011101",
  19606=>"010111101",
  19607=>"101011010",
  19608=>"111011001",
  19609=>"010101100",
  19610=>"001001101",
  19611=>"111101111",
  19612=>"001100011",
  19613=>"010110000",
  19614=>"111110000",
  19615=>"000101001",
  19616=>"101110110",
  19617=>"010110011",
  19618=>"110001111",
  19619=>"010011000",
  19620=>"101101001",
  19621=>"000000110",
  19622=>"001001011",
  19623=>"101110101",
  19624=>"100011010",
  19625=>"110111011",
  19626=>"001111110",
  19627=>"111000101",
  19628=>"111101010",
  19629=>"100000000",
  19630=>"010111110",
  19631=>"011000001",
  19632=>"100000010",
  19633=>"111101000",
  19634=>"011000111",
  19635=>"001000100",
  19636=>"110000000",
  19637=>"001001011",
  19638=>"011110110",
  19639=>"001101111",
  19640=>"111100011",
  19641=>"011000110",
  19642=>"111011001",
  19643=>"110000000",
  19644=>"011101001",
  19645=>"101101111",
  19646=>"111001110",
  19647=>"110010011",
  19648=>"111100110",
  19649=>"010100000",
  19650=>"011000011",
  19651=>"000100110",
  19652=>"100111000",
  19653=>"010010000",
  19654=>"101110010",
  19655=>"010011100",
  19656=>"111001001",
  19657=>"101100100",
  19658=>"111010000",
  19659=>"100110110",
  19660=>"101101010",
  19661=>"000100111",
  19662=>"010000101",
  19663=>"011011001",
  19664=>"011010101",
  19665=>"000111001",
  19666=>"010000111",
  19667=>"010001100",
  19668=>"001000001",
  19669=>"000010010",
  19670=>"001001001",
  19671=>"000110111",
  19672=>"101110110",
  19673=>"101111111",
  19674=>"000000000",
  19675=>"111100101",
  19676=>"101100110",
  19677=>"010000001",
  19678=>"111111101",
  19679=>"110111100",
  19680=>"100010000",
  19681=>"001110011",
  19682=>"101000011",
  19683=>"000111111",
  19684=>"011010100",
  19685=>"011100111",
  19686=>"110101000",
  19687=>"100000010",
  19688=>"011111111",
  19689=>"100001010",
  19690=>"100101110",
  19691=>"000110111",
  19692=>"001011101",
  19693=>"001110110",
  19694=>"010100010",
  19695=>"000011100",
  19696=>"111110110",
  19697=>"001100001",
  19698=>"000010100",
  19699=>"100011100",
  19700=>"110001111",
  19701=>"001010110",
  19702=>"100101000",
  19703=>"101000000",
  19704=>"110101100",
  19705=>"110011110",
  19706=>"001101011",
  19707=>"111011000",
  19708=>"000100001",
  19709=>"011100010",
  19710=>"011001010",
  19711=>"101111000",
  19712=>"110110000",
  19713=>"011101100",
  19714=>"000100101",
  19715=>"001000110",
  19716=>"010000010",
  19717=>"101000010",
  19718=>"111010100",
  19719=>"011010001",
  19720=>"000100111",
  19721=>"110001111",
  19722=>"100010100",
  19723=>"111110000",
  19724=>"001110011",
  19725=>"110010110",
  19726=>"100011010",
  19727=>"001001001",
  19728=>"101000101",
  19729=>"111110001",
  19730=>"100110001",
  19731=>"100011101",
  19732=>"000101001",
  19733=>"101110011",
  19734=>"011110010",
  19735=>"010011110",
  19736=>"000011001",
  19737=>"111010011",
  19738=>"111011101",
  19739=>"110101100",
  19740=>"011000100",
  19741=>"101000110",
  19742=>"000011000",
  19743=>"100101011",
  19744=>"000001010",
  19745=>"101010011",
  19746=>"000010110",
  19747=>"011000100",
  19748=>"010110010",
  19749=>"010010100",
  19750=>"010000010",
  19751=>"010110110",
  19752=>"010000000",
  19753=>"100100110",
  19754=>"010001011",
  19755=>"110111101",
  19756=>"110001100",
  19757=>"111111100",
  19758=>"000001001",
  19759=>"010011110",
  19760=>"011000010",
  19761=>"010001000",
  19762=>"111100111",
  19763=>"011000111",
  19764=>"000110011",
  19765=>"100110000",
  19766=>"000000010",
  19767=>"110000011",
  19768=>"101110110",
  19769=>"110100010",
  19770=>"000111100",
  19771=>"100010000",
  19772=>"001011110",
  19773=>"000010001",
  19774=>"010011101",
  19775=>"010001110",
  19776=>"100010011",
  19777=>"001011000",
  19778=>"101101001",
  19779=>"100101000",
  19780=>"100001010",
  19781=>"110011011",
  19782=>"111000000",
  19783=>"000100111",
  19784=>"111111000",
  19785=>"100000000",
  19786=>"010001100",
  19787=>"010101101",
  19788=>"001110101",
  19789=>"101011100",
  19790=>"100000001",
  19791=>"011100110",
  19792=>"011111011",
  19793=>"010000001",
  19794=>"101110000",
  19795=>"000101010",
  19796=>"000110001",
  19797=>"010111100",
  19798=>"011111110",
  19799=>"111000001",
  19800=>"000001001",
  19801=>"100001010",
  19802=>"011001010",
  19803=>"000000011",
  19804=>"010010000",
  19805=>"000011010",
  19806=>"111001100",
  19807=>"011001000",
  19808=>"101001010",
  19809=>"011011001",
  19810=>"111011111",
  19811=>"001100011",
  19812=>"011011001",
  19813=>"100100000",
  19814=>"110010010",
  19815=>"101000100",
  19816=>"101001100",
  19817=>"001001011",
  19818=>"110000101",
  19819=>"010100111",
  19820=>"001000010",
  19821=>"000110111",
  19822=>"010101111",
  19823=>"100110011",
  19824=>"010010010",
  19825=>"100000100",
  19826=>"100010001",
  19827=>"000101010",
  19828=>"000110000",
  19829=>"000011010",
  19830=>"101000111",
  19831=>"010100000",
  19832=>"101100011",
  19833=>"101010001",
  19834=>"100011010",
  19835=>"110000001",
  19836=>"000010100",
  19837=>"100111110",
  19838=>"001010011",
  19839=>"110000100",
  19840=>"100111000",
  19841=>"011100111",
  19842=>"001111101",
  19843=>"010000100",
  19844=>"011100111",
  19845=>"100000000",
  19846=>"110101100",
  19847=>"101011001",
  19848=>"000100011",
  19849=>"111011101",
  19850=>"101001000",
  19851=>"110111010",
  19852=>"110101111",
  19853=>"010001001",
  19854=>"001001000",
  19855=>"100100000",
  19856=>"110101110",
  19857=>"000011010",
  19858=>"100001001",
  19859=>"100101010",
  19860=>"001010101",
  19861=>"100100000",
  19862=>"111100101",
  19863=>"101101011",
  19864=>"000001101",
  19865=>"000101010",
  19866=>"010100101",
  19867=>"110101000",
  19868=>"100111111",
  19869=>"101100011",
  19870=>"001001001",
  19871=>"000010110",
  19872=>"000100101",
  19873=>"000011110",
  19874=>"100111010",
  19875=>"101000001",
  19876=>"010101000",
  19877=>"100110101",
  19878=>"010111011",
  19879=>"111101110",
  19880=>"000110110",
  19881=>"010001111",
  19882=>"001101111",
  19883=>"111111101",
  19884=>"000010000",
  19885=>"011000000",
  19886=>"011011010",
  19887=>"001110011",
  19888=>"001101101",
  19889=>"111011101",
  19890=>"001110000",
  19891=>"010100000",
  19892=>"000111111",
  19893=>"111000011",
  19894=>"100110101",
  19895=>"011010011",
  19896=>"011101111",
  19897=>"000011111",
  19898=>"101000000",
  19899=>"010000010",
  19900=>"010110011",
  19901=>"100001111",
  19902=>"101111101",
  19903=>"011110011",
  19904=>"111010110",
  19905=>"011101001",
  19906=>"101110100",
  19907=>"001101111",
  19908=>"000100100",
  19909=>"111001010",
  19910=>"011001000",
  19911=>"011000111",
  19912=>"001110001",
  19913=>"100011101",
  19914=>"011000000",
  19915=>"111111000",
  19916=>"111001100",
  19917=>"111000000",
  19918=>"111100000",
  19919=>"001100000",
  19920=>"101011100",
  19921=>"001101011",
  19922=>"111100010",
  19923=>"001011001",
  19924=>"010000100",
  19925=>"000101010",
  19926=>"000010110",
  19927=>"100100101",
  19928=>"001101010",
  19929=>"101000011",
  19930=>"011000000",
  19931=>"111000111",
  19932=>"100111101",
  19933=>"001000011",
  19934=>"101111011",
  19935=>"001001111",
  19936=>"101111111",
  19937=>"100000000",
  19938=>"100111110",
  19939=>"101000010",
  19940=>"001101000",
  19941=>"000101011",
  19942=>"000000110",
  19943=>"100111001",
  19944=>"100110011",
  19945=>"110011011",
  19946=>"011111010",
  19947=>"100000100",
  19948=>"100000100",
  19949=>"000011000",
  19950=>"011011101",
  19951=>"001000100",
  19952=>"001011111",
  19953=>"000000010",
  19954=>"001100100",
  19955=>"011001000",
  19956=>"110101000",
  19957=>"011001010",
  19958=>"010110100",
  19959=>"011011000",
  19960=>"100010100",
  19961=>"100101011",
  19962=>"011101101",
  19963=>"011111111",
  19964=>"101001000",
  19965=>"000111111",
  19966=>"000101110",
  19967=>"011110010",
  19968=>"010000001",
  19969=>"110110011",
  19970=>"111110100",
  19971=>"010110100",
  19972=>"010001101",
  19973=>"001100010",
  19974=>"111000000",
  19975=>"010100001",
  19976=>"100100111",
  19977=>"101110111",
  19978=>"100000001",
  19979=>"000000000",
  19980=>"100101110",
  19981=>"010110111",
  19982=>"001010010",
  19983=>"001100110",
  19984=>"011010100",
  19985=>"100010011",
  19986=>"010101011",
  19987=>"110110001",
  19988=>"111000011",
  19989=>"010101000",
  19990=>"111100011",
  19991=>"010101100",
  19992=>"101000101",
  19993=>"001001011",
  19994=>"001000001",
  19995=>"011110001",
  19996=>"011100110",
  19997=>"010101011",
  19998=>"011001000",
  19999=>"001000100",
  20000=>"011101110",
  20001=>"111011011",
  20002=>"010101100",
  20003=>"001000001",
  20004=>"101101010",
  20005=>"110010000",
  20006=>"001000111",
  20007=>"000010110",
  20008=>"001111111",
  20009=>"110100111",
  20010=>"110010100",
  20011=>"111101011",
  20012=>"010101110",
  20013=>"010001011",
  20014=>"010001010",
  20015=>"100000010",
  20016=>"110000011",
  20017=>"111001011",
  20018=>"011001011",
  20019=>"100000101",
  20020=>"100000010",
  20021=>"100111010",
  20022=>"011011101",
  20023=>"110011101",
  20024=>"111001100",
  20025=>"001011001",
  20026=>"010000010",
  20027=>"010011101",
  20028=>"111001011",
  20029=>"111100011",
  20030=>"010010101",
  20031=>"111011110",
  20032=>"110001100",
  20033=>"001111001",
  20034=>"100000001",
  20035=>"000010000",
  20036=>"000000110",
  20037=>"011100000",
  20038=>"101111001",
  20039=>"100100011",
  20040=>"111101100",
  20041=>"000101011",
  20042=>"000001000",
  20043=>"000111100",
  20044=>"100101001",
  20045=>"101010111",
  20046=>"011100111",
  20047=>"110000100",
  20048=>"101000011",
  20049=>"001110101",
  20050=>"101110000",
  20051=>"000000001",
  20052=>"000011011",
  20053=>"011111001",
  20054=>"010100010",
  20055=>"011100010",
  20056=>"001000111",
  20057=>"101010001",
  20058=>"000000100",
  20059=>"000001101",
  20060=>"001010101",
  20061=>"110001100",
  20062=>"000100111",
  20063=>"011001100",
  20064=>"101100011",
  20065=>"100011011",
  20066=>"111100000",
  20067=>"101100010",
  20068=>"011011011",
  20069=>"010000100",
  20070=>"000100000",
  20071=>"010100100",
  20072=>"111011101",
  20073=>"101000100",
  20074=>"011111000",
  20075=>"001110011",
  20076=>"000110011",
  20077=>"011011001",
  20078=>"110110011",
  20079=>"011111011",
  20080=>"011000111",
  20081=>"100011101",
  20082=>"000101101",
  20083=>"001011111",
  20084=>"110100000",
  20085=>"001111100",
  20086=>"100001000",
  20087=>"100100000",
  20088=>"101000100",
  20089=>"000110010",
  20090=>"101011010",
  20091=>"111011010",
  20092=>"000001011",
  20093=>"100110010",
  20094=>"110101000",
  20095=>"000011101",
  20096=>"101101001",
  20097=>"111100100",
  20098=>"000001011",
  20099=>"010001101",
  20100=>"111001110",
  20101=>"100001100",
  20102=>"110001011",
  20103=>"110001000",
  20104=>"000011101",
  20105=>"000001101",
  20106=>"110001111",
  20107=>"010010000",
  20108=>"000011101",
  20109=>"110101011",
  20110=>"100101100",
  20111=>"000000001",
  20112=>"010110001",
  20113=>"000100010",
  20114=>"111010110",
  20115=>"100100101",
  20116=>"010100100",
  20117=>"010110010",
  20118=>"000010000",
  20119=>"101010001",
  20120=>"000011101",
  20121=>"010011111",
  20122=>"110001111",
  20123=>"010111100",
  20124=>"101110111",
  20125=>"101101100",
  20126=>"100011001",
  20127=>"001100011",
  20128=>"011101011",
  20129=>"010001110",
  20130=>"000000011",
  20131=>"010001110",
  20132=>"100110111",
  20133=>"100111000",
  20134=>"000010010",
  20135=>"001100010",
  20136=>"011100000",
  20137=>"101111010",
  20138=>"000010110",
  20139=>"010110101",
  20140=>"101000101",
  20141=>"001110010",
  20142=>"001100100",
  20143=>"010111011",
  20144=>"001010001",
  20145=>"010010111",
  20146=>"001001101",
  20147=>"011001111",
  20148=>"010111111",
  20149=>"010111111",
  20150=>"011111011",
  20151=>"000111000",
  20152=>"110011100",
  20153=>"101011110",
  20154=>"001100101",
  20155=>"101001011",
  20156=>"000100001",
  20157=>"010111011",
  20158=>"011000000",
  20159=>"101010100",
  20160=>"101000110",
  20161=>"001001011",
  20162=>"010001011",
  20163=>"111000010",
  20164=>"100011001",
  20165=>"100111100",
  20166=>"100101100",
  20167=>"010111011",
  20168=>"101111100",
  20169=>"110001001",
  20170=>"011101100",
  20171=>"000100010",
  20172=>"001010100",
  20173=>"001010011",
  20174=>"100011011",
  20175=>"010000010",
  20176=>"000111011",
  20177=>"110010111",
  20178=>"010110100",
  20179=>"001000101",
  20180=>"100110101",
  20181=>"100111101",
  20182=>"101000011",
  20183=>"011000011",
  20184=>"001010001",
  20185=>"010010001",
  20186=>"111110101",
  20187=>"110101110",
  20188=>"010101001",
  20189=>"111010110",
  20190=>"110001101",
  20191=>"110010110",
  20192=>"011000001",
  20193=>"101110000",
  20194=>"110110111",
  20195=>"011011000",
  20196=>"010001101",
  20197=>"001100011",
  20198=>"011110001",
  20199=>"110111010",
  20200=>"110011001",
  20201=>"001010100",
  20202=>"000010000",
  20203=>"001101011",
  20204=>"011100000",
  20205=>"100110011",
  20206=>"101100111",
  20207=>"000010011",
  20208=>"110111111",
  20209=>"111011000",
  20210=>"110100110",
  20211=>"101011111",
  20212=>"100010101",
  20213=>"110011010",
  20214=>"111110011",
  20215=>"000010110",
  20216=>"111011110",
  20217=>"001101100",
  20218=>"110110111",
  20219=>"001011000",
  20220=>"111101101",
  20221=>"101001011",
  20222=>"010000110",
  20223=>"010100010",
  20224=>"101101101",
  20225=>"000010110",
  20226=>"101011100",
  20227=>"011100010",
  20228=>"110000000",
  20229=>"100110100",
  20230=>"111110100",
  20231=>"110110000",
  20232=>"111001001",
  20233=>"101111010",
  20234=>"100010011",
  20235=>"000111010",
  20236=>"000001010",
  20237=>"100010010",
  20238=>"100000100",
  20239=>"001110010",
  20240=>"110010110",
  20241=>"000110111",
  20242=>"111101100",
  20243=>"100000101",
  20244=>"101001001",
  20245=>"110010000",
  20246=>"111010000",
  20247=>"011011100",
  20248=>"111011100",
  20249=>"011111011",
  20250=>"001101010",
  20251=>"001100110",
  20252=>"010110001",
  20253=>"111001010",
  20254=>"001100010",
  20255=>"100111011",
  20256=>"110001111",
  20257=>"111010101",
  20258=>"011001011",
  20259=>"011101001",
  20260=>"101101100",
  20261=>"101001111",
  20262=>"101010010",
  20263=>"110111001",
  20264=>"110000000",
  20265=>"000010110",
  20266=>"011100011",
  20267=>"010111010",
  20268=>"000111100",
  20269=>"001000001",
  20270=>"011010001",
  20271=>"110001010",
  20272=>"010111101",
  20273=>"000011111",
  20274=>"010111010",
  20275=>"101011001",
  20276=>"011110101",
  20277=>"110010001",
  20278=>"000001011",
  20279=>"011101100",
  20280=>"101010110",
  20281=>"110101001",
  20282=>"111111111",
  20283=>"000100111",
  20284=>"001001101",
  20285=>"000000000",
  20286=>"111110110",
  20287=>"101111011",
  20288=>"110010001",
  20289=>"100110001",
  20290=>"101100011",
  20291=>"011010110",
  20292=>"100010101",
  20293=>"010010100",
  20294=>"110110001",
  20295=>"010110101",
  20296=>"000001101",
  20297=>"000101011",
  20298=>"101111011",
  20299=>"011011101",
  20300=>"111010110",
  20301=>"101111101",
  20302=>"011101011",
  20303=>"101110100",
  20304=>"110110101",
  20305=>"010001010",
  20306=>"111000000",
  20307=>"000101100",
  20308=>"011100100",
  20309=>"110100111",
  20310=>"011011110",
  20311=>"000111111",
  20312=>"100001000",
  20313=>"100100100",
  20314=>"101111100",
  20315=>"011110100",
  20316=>"101001001",
  20317=>"010101100",
  20318=>"011111011",
  20319=>"000001100",
  20320=>"110110001",
  20321=>"111010100",
  20322=>"010101000",
  20323=>"001011000",
  20324=>"100001001",
  20325=>"000110110",
  20326=>"111000111",
  20327=>"000101110",
  20328=>"111101111",
  20329=>"000110010",
  20330=>"111010000",
  20331=>"011110001",
  20332=>"100100100",
  20333=>"110000011",
  20334=>"111111000",
  20335=>"101100111",
  20336=>"010110110",
  20337=>"111000001",
  20338=>"000100000",
  20339=>"000001010",
  20340=>"010011000",
  20341=>"111110110",
  20342=>"101111100",
  20343=>"100101100",
  20344=>"110010100",
  20345=>"101100010",
  20346=>"010000101",
  20347=>"111101001",
  20348=>"010100100",
  20349=>"010011010",
  20350=>"101111111",
  20351=>"111111010",
  20352=>"010111110",
  20353=>"100101110",
  20354=>"000101010",
  20355=>"111100011",
  20356=>"101110110",
  20357=>"001110010",
  20358=>"010010000",
  20359=>"000000000",
  20360=>"001100111",
  20361=>"100101010",
  20362=>"110111010",
  20363=>"010100011",
  20364=>"100010011",
  20365=>"100010010",
  20366=>"010001111",
  20367=>"000001100",
  20368=>"100110110",
  20369=>"111000010",
  20370=>"001110011",
  20371=>"110010000",
  20372=>"111111111",
  20373=>"100001001",
  20374=>"000100001",
  20375=>"011111011",
  20376=>"110010110",
  20377=>"000101011",
  20378=>"010011000",
  20379=>"001001000",
  20380=>"101000111",
  20381=>"110110100",
  20382=>"110111101",
  20383=>"010001111",
  20384=>"011001011",
  20385=>"111110010",
  20386=>"110100101",
  20387=>"111101111",
  20388=>"000101101",
  20389=>"000001101",
  20390=>"010001110",
  20391=>"001010111",
  20392=>"111010110",
  20393=>"001110111",
  20394=>"100011000",
  20395=>"101110001",
  20396=>"001110100",
  20397=>"110001011",
  20398=>"110000110",
  20399=>"001011100",
  20400=>"011010100",
  20401=>"001001100",
  20402=>"000110011",
  20403=>"111111001",
  20404=>"010101000",
  20405=>"001001010",
  20406=>"110011001",
  20407=>"101001100",
  20408=>"111011101",
  20409=>"111111100",
  20410=>"000001000",
  20411=>"100000100",
  20412=>"110001001",
  20413=>"111000110",
  20414=>"111110111",
  20415=>"011001111",
  20416=>"011011010",
  20417=>"001000010",
  20418=>"110001111",
  20419=>"111101100",
  20420=>"001101010",
  20421=>"100010010",
  20422=>"110100010",
  20423=>"111110100",
  20424=>"110110011",
  20425=>"010010111",
  20426=>"010110110",
  20427=>"101000100",
  20428=>"110110000",
  20429=>"111001111",
  20430=>"000011101",
  20431=>"001101011",
  20432=>"001111001",
  20433=>"101000000",
  20434=>"100011011",
  20435=>"011110110",
  20436=>"001001011",
  20437=>"000011000",
  20438=>"000100101",
  20439=>"111001000",
  20440=>"010110000",
  20441=>"000011010",
  20442=>"111110010",
  20443=>"111110010",
  20444=>"111111111",
  20445=>"110101010",
  20446=>"011101001",
  20447=>"100110000",
  20448=>"001011111",
  20449=>"010100011",
  20450=>"110111111",
  20451=>"010010000",
  20452=>"101011000",
  20453=>"010010001",
  20454=>"000100111",
  20455=>"010001010",
  20456=>"111010011",
  20457=>"011010111",
  20458=>"110111000",
  20459=>"100011110",
  20460=>"010101011",
  20461=>"000101111",
  20462=>"111100111",
  20463=>"101011101",
  20464=>"011111111",
  20465=>"101000000",
  20466=>"101100011",
  20467=>"111100000",
  20468=>"001110001",
  20469=>"100110000",
  20470=>"111111001",
  20471=>"111001011",
  20472=>"000000000",
  20473=>"000110001",
  20474=>"100100110",
  20475=>"111101100",
  20476=>"000101010",
  20477=>"001000101",
  20478=>"010110101",
  20479=>"111101101",
  20480=>"101010100",
  20481=>"111111000",
  20482=>"110101110",
  20483=>"010101101",
  20484=>"110010111",
  20485=>"010111110",
  20486=>"110111001",
  20487=>"010011010",
  20488=>"111110100",
  20489=>"001110111",
  20490=>"110110101",
  20491=>"101110101",
  20492=>"110000111",
  20493=>"011000100",
  20494=>"110100000",
  20495=>"110100000",
  20496=>"001010111",
  20497=>"111001001",
  20498=>"111100001",
  20499=>"000011110",
  20500=>"000000011",
  20501=>"010001010",
  20502=>"100010011",
  20503=>"101000000",
  20504=>"100111101",
  20505=>"001110100",
  20506=>"110011011",
  20507=>"011110001",
  20508=>"110101111",
  20509=>"001110001",
  20510=>"100110111",
  20511=>"110101100",
  20512=>"011101001",
  20513=>"100101011",
  20514=>"101100111",
  20515=>"001011011",
  20516=>"011110100",
  20517=>"111000100",
  20518=>"100101100",
  20519=>"001011101",
  20520=>"001010000",
  20521=>"011011010",
  20522=>"100011011",
  20523=>"111011001",
  20524=>"010100001",
  20525=>"000001101",
  20526=>"001100111",
  20527=>"110101100",
  20528=>"010111011",
  20529=>"011100011",
  20530=>"010000000",
  20531=>"011111100",
  20532=>"000011110",
  20533=>"011101111",
  20534=>"011001110",
  20535=>"001010011",
  20536=>"001010111",
  20537=>"110010001",
  20538=>"010110011",
  20539=>"001000010",
  20540=>"101000011",
  20541=>"001110100",
  20542=>"000001111",
  20543=>"101111001",
  20544=>"100011011",
  20545=>"111010000",
  20546=>"011010100",
  20547=>"010001101",
  20548=>"111000110",
  20549=>"000010011",
  20550=>"110101001",
  20551=>"011101000",
  20552=>"101110011",
  20553=>"000111011",
  20554=>"010110010",
  20555=>"000010011",
  20556=>"011001001",
  20557=>"100100110",
  20558=>"001100111",
  20559=>"000110111",
  20560=>"101000111",
  20561=>"110110101",
  20562=>"101100000",
  20563=>"110001011",
  20564=>"001111111",
  20565=>"000011000",
  20566=>"010110011",
  20567=>"000001011",
  20568=>"111100110",
  20569=>"011111101",
  20570=>"001001110",
  20571=>"011011111",
  20572=>"000011100",
  20573=>"000011010",
  20574=>"001011011",
  20575=>"110000110",
  20576=>"100111010",
  20577=>"010011100",
  20578=>"000000000",
  20579=>"101000010",
  20580=>"001101001",
  20581=>"101111001",
  20582=>"100101100",
  20583=>"010100000",
  20584=>"001110111",
  20585=>"010011011",
  20586=>"010100111",
  20587=>"110001011",
  20588=>"000000000",
  20589=>"111000110",
  20590=>"101001101",
  20591=>"000011111",
  20592=>"000011100",
  20593=>"011011011",
  20594=>"110101110",
  20595=>"000100001",
  20596=>"100000001",
  20597=>"111110101",
  20598=>"010110011",
  20599=>"011011111",
  20600=>"110100011",
  20601=>"110101101",
  20602=>"010000000",
  20603=>"000010100",
  20604=>"100000101",
  20605=>"000101101",
  20606=>"000000111",
  20607=>"101011100",
  20608=>"111010010",
  20609=>"000111000",
  20610=>"010010100",
  20611=>"111010010",
  20612=>"000111011",
  20613=>"000111110",
  20614=>"011110010",
  20615=>"100000000",
  20616=>"010110111",
  20617=>"000100001",
  20618=>"111101100",
  20619=>"010011111",
  20620=>"110000111",
  20621=>"000111101",
  20622=>"000001100",
  20623=>"000111100",
  20624=>"000001000",
  20625=>"011110000",
  20626=>"011111111",
  20627=>"011110010",
  20628=>"000100100",
  20629=>"100010100",
  20630=>"100010000",
  20631=>"010100001",
  20632=>"101110001",
  20633=>"110100110",
  20634=>"011110001",
  20635=>"110010011",
  20636=>"000001000",
  20637=>"110111011",
  20638=>"001110101",
  20639=>"000000010",
  20640=>"001110100",
  20641=>"111111011",
  20642=>"011010111",
  20643=>"101001010",
  20644=>"001000010",
  20645=>"000111101",
  20646=>"101111001",
  20647=>"101101010",
  20648=>"111001010",
  20649=>"001001100",
  20650=>"111100110",
  20651=>"110100110",
  20652=>"010001101",
  20653=>"110111001",
  20654=>"011111011",
  20655=>"000111101",
  20656=>"011011000",
  20657=>"010010110",
  20658=>"011110110",
  20659=>"100011001",
  20660=>"101010110",
  20661=>"001010010",
  20662=>"000001011",
  20663=>"010111110",
  20664=>"011110110",
  20665=>"011100100",
  20666=>"011111010",
  20667=>"010111111",
  20668=>"000000011",
  20669=>"110011010",
  20670=>"100101011",
  20671=>"000100111",
  20672=>"010000001",
  20673=>"011101101",
  20674=>"011010011",
  20675=>"100011110",
  20676=>"101111111",
  20677=>"011001001",
  20678=>"010110100",
  20679=>"101010110",
  20680=>"010111000",
  20681=>"001101110",
  20682=>"111101001",
  20683=>"000101101",
  20684=>"101001101",
  20685=>"101000110",
  20686=>"111000111",
  20687=>"100001000",
  20688=>"100101101",
  20689=>"101110101",
  20690=>"101110001",
  20691=>"110010111",
  20692=>"101111001",
  20693=>"101100010",
  20694=>"001110000",
  20695=>"111011001",
  20696=>"010111100",
  20697=>"100010110",
  20698=>"010010011",
  20699=>"000110001",
  20700=>"100001000",
  20701=>"010111000",
  20702=>"001110101",
  20703=>"100101101",
  20704=>"000110011",
  20705=>"000010000",
  20706=>"001000000",
  20707=>"100100001",
  20708=>"111010001",
  20709=>"000101110",
  20710=>"100110000",
  20711=>"010000111",
  20712=>"011000101",
  20713=>"011101000",
  20714=>"001011001",
  20715=>"001101101",
  20716=>"101010101",
  20717=>"001100111",
  20718=>"011011100",
  20719=>"000101101",
  20720=>"101110010",
  20721=>"000011010",
  20722=>"111011011",
  20723=>"001100111",
  20724=>"001111110",
  20725=>"010111111",
  20726=>"100111000",
  20727=>"000000001",
  20728=>"010100100",
  20729=>"001110001",
  20730=>"101111010",
  20731=>"000010101",
  20732=>"100110001",
  20733=>"000110011",
  20734=>"011100111",
  20735=>"110110101",
  20736=>"101101101",
  20737=>"111100010",
  20738=>"001000010",
  20739=>"110011000",
  20740=>"110101110",
  20741=>"110011011",
  20742=>"101100001",
  20743=>"110001011",
  20744=>"011010010",
  20745=>"100110010",
  20746=>"010011010",
  20747=>"000001100",
  20748=>"010001000",
  20749=>"100010010",
  20750=>"100000000",
  20751=>"000101000",
  20752=>"111011110",
  20753=>"000101101",
  20754=>"010011101",
  20755=>"110010101",
  20756=>"101100010",
  20757=>"111110000",
  20758=>"101010100",
  20759=>"010000101",
  20760=>"111000010",
  20761=>"101011011",
  20762=>"001110001",
  20763=>"100101111",
  20764=>"111011001",
  20765=>"000011111",
  20766=>"010000111",
  20767=>"011011010",
  20768=>"000011011",
  20769=>"100100110",
  20770=>"000001000",
  20771=>"010111001",
  20772=>"000110011",
  20773=>"001001011",
  20774=>"100101100",
  20775=>"100000100",
  20776=>"000001110",
  20777=>"001010111",
  20778=>"011101010",
  20779=>"010110011",
  20780=>"111101111",
  20781=>"100001010",
  20782=>"111000100",
  20783=>"010100110",
  20784=>"011101110",
  20785=>"111111101",
  20786=>"111000000",
  20787=>"000111110",
  20788=>"110001011",
  20789=>"001000001",
  20790=>"100011110",
  20791=>"011101001",
  20792=>"000100111",
  20793=>"000010101",
  20794=>"110100100",
  20795=>"000001100",
  20796=>"010101110",
  20797=>"111010100",
  20798=>"100100110",
  20799=>"000010101",
  20800=>"011110011",
  20801=>"000000111",
  20802=>"100001100",
  20803=>"100000000",
  20804=>"000011101",
  20805=>"111101111",
  20806=>"100100001",
  20807=>"010111010",
  20808=>"111101010",
  20809=>"111110100",
  20810=>"011010000",
  20811=>"000000111",
  20812=>"101011110",
  20813=>"011010101",
  20814=>"110111111",
  20815=>"011001101",
  20816=>"101001111",
  20817=>"111110101",
  20818=>"010000100",
  20819=>"101011100",
  20820=>"101101111",
  20821=>"101001111",
  20822=>"110000110",
  20823=>"000110010",
  20824=>"100000001",
  20825=>"101100101",
  20826=>"100111011",
  20827=>"011111111",
  20828=>"110111001",
  20829=>"010010110",
  20830=>"111111000",
  20831=>"011111000",
  20832=>"000000000",
  20833=>"101011000",
  20834=>"100100100",
  20835=>"000100010",
  20836=>"111011101",
  20837=>"000101000",
  20838=>"000110000",
  20839=>"111111111",
  20840=>"100110101",
  20841=>"000110011",
  20842=>"010101100",
  20843=>"101010011",
  20844=>"110101010",
  20845=>"001011000",
  20846=>"010000000",
  20847=>"110010101",
  20848=>"000110000",
  20849=>"000110001",
  20850=>"110101011",
  20851=>"110111000",
  20852=>"111111011",
  20853=>"001011011",
  20854=>"001110100",
  20855=>"101101001",
  20856=>"001111101",
  20857=>"100010000",
  20858=>"111110011",
  20859=>"101110110",
  20860=>"000000010",
  20861=>"100011001",
  20862=>"101010101",
  20863=>"001000001",
  20864=>"100101010",
  20865=>"000010010",
  20866=>"011110101",
  20867=>"100001100",
  20868=>"100110011",
  20869=>"101001111",
  20870=>"001010111",
  20871=>"111001101",
  20872=>"000010101",
  20873=>"111001110",
  20874=>"100100100",
  20875=>"110000000",
  20876=>"000110110",
  20877=>"001000110",
  20878=>"111111011",
  20879=>"100001101",
  20880=>"000101110",
  20881=>"110000100",
  20882=>"001001101",
  20883=>"001100011",
  20884=>"000000100",
  20885=>"101111010",
  20886=>"110111011",
  20887=>"111010101",
  20888=>"111010101",
  20889=>"111110010",
  20890=>"111101010",
  20891=>"101000101",
  20892=>"000011110",
  20893=>"101100111",
  20894=>"000110011",
  20895=>"111111111",
  20896=>"010101111",
  20897=>"111000101",
  20898=>"011101010",
  20899=>"000101100",
  20900=>"011000010",
  20901=>"100110110",
  20902=>"011000001",
  20903=>"000101110",
  20904=>"100011110",
  20905=>"110101110",
  20906=>"000001000",
  20907=>"011011000",
  20908=>"010100100",
  20909=>"111111110",
  20910=>"010010100",
  20911=>"110010000",
  20912=>"011100000",
  20913=>"010111110",
  20914=>"110101111",
  20915=>"001001000",
  20916=>"101101010",
  20917=>"000111001",
  20918=>"010100101",
  20919=>"001110100",
  20920=>"001000111",
  20921=>"100101010",
  20922=>"000000000",
  20923=>"011011000",
  20924=>"101111111",
  20925=>"001000110",
  20926=>"011111101",
  20927=>"110101011",
  20928=>"000111000",
  20929=>"101001101",
  20930=>"011100001",
  20931=>"000111110",
  20932=>"001010000",
  20933=>"001011000",
  20934=>"000011011",
  20935=>"000111101",
  20936=>"001000001",
  20937=>"110011101",
  20938=>"000011111",
  20939=>"001101110",
  20940=>"111000110",
  20941=>"000111001",
  20942=>"101001000",
  20943=>"001110011",
  20944=>"101000000",
  20945=>"000000111",
  20946=>"001110101",
  20947=>"100100001",
  20948=>"010011100",
  20949=>"010111110",
  20950=>"100101011",
  20951=>"100110100",
  20952=>"000000001",
  20953=>"101111011",
  20954=>"011100001",
  20955=>"110100011",
  20956=>"000000101",
  20957=>"100110011",
  20958=>"000011010",
  20959=>"110000000",
  20960=>"000011100",
  20961=>"010000000",
  20962=>"010101110",
  20963=>"111001111",
  20964=>"100111101",
  20965=>"000101011",
  20966=>"111100010",
  20967=>"111000000",
  20968=>"010001010",
  20969=>"110101010",
  20970=>"101011001",
  20971=>"001111010",
  20972=>"100101110",
  20973=>"100100101",
  20974=>"001000000",
  20975=>"110000000",
  20976=>"000011011",
  20977=>"000100110",
  20978=>"111010001",
  20979=>"000100100",
  20980=>"000110000",
  20981=>"100001101",
  20982=>"000110001",
  20983=>"100011111",
  20984=>"000000000",
  20985=>"000001000",
  20986=>"101100010",
  20987=>"000100110",
  20988=>"101011110",
  20989=>"110011110",
  20990=>"001101101",
  20991=>"110010011",
  20992=>"000010110",
  20993=>"111110001",
  20994=>"011001110",
  20995=>"000000100",
  20996=>"000111011",
  20997=>"011001100",
  20998=>"110110010",
  20999=>"011010101",
  21000=>"001110110",
  21001=>"000011110",
  21002=>"110011101",
  21003=>"010011010",
  21004=>"101010001",
  21005=>"101010100",
  21006=>"100000100",
  21007=>"110111110",
  21008=>"100100110",
  21009=>"100001101",
  21010=>"011110001",
  21011=>"000011111",
  21012=>"001101001",
  21013=>"100010101",
  21014=>"111011101",
  21015=>"110101010",
  21016=>"011011010",
  21017=>"000100110",
  21018=>"010100000",
  21019=>"000000101",
  21020=>"111111010",
  21021=>"000101010",
  21022=>"000101110",
  21023=>"111110110",
  21024=>"111000001",
  21025=>"001001110",
  21026=>"000001110",
  21027=>"010010111",
  21028=>"011111100",
  21029=>"000110111",
  21030=>"110110011",
  21031=>"110000110",
  21032=>"100011000",
  21033=>"100111011",
  21034=>"011000000",
  21035=>"100101001",
  21036=>"111001001",
  21037=>"100111110",
  21038=>"101001101",
  21039=>"111011011",
  21040=>"010111100",
  21041=>"111101010",
  21042=>"000011000",
  21043=>"101111110",
  21044=>"011100011",
  21045=>"100011011",
  21046=>"111000000",
  21047=>"110111010",
  21048=>"110010010",
  21049=>"111110111",
  21050=>"101010110",
  21051=>"000011011",
  21052=>"000100000",
  21053=>"010110001",
  21054=>"011111100",
  21055=>"101000111",
  21056=>"001001010",
  21057=>"000000111",
  21058=>"110100110",
  21059=>"100011110",
  21060=>"100001101",
  21061=>"110110111",
  21062=>"011100000",
  21063=>"111101110",
  21064=>"001001101",
  21065=>"011000101",
  21066=>"001000010",
  21067=>"011100100",
  21068=>"010100000",
  21069=>"101000100",
  21070=>"110001011",
  21071=>"011011111",
  21072=>"100110001",
  21073=>"010010101",
  21074=>"000011011",
  21075=>"001001011",
  21076=>"101000110",
  21077=>"001011101",
  21078=>"111111011",
  21079=>"101011100",
  21080=>"111110100",
  21081=>"000010001",
  21082=>"111001011",
  21083=>"111001100",
  21084=>"011001111",
  21085=>"111100011",
  21086=>"001110011",
  21087=>"011100011",
  21088=>"100000011",
  21089=>"000001011",
  21090=>"101111111",
  21091=>"110111111",
  21092=>"111100000",
  21093=>"110011000",
  21094=>"111010101",
  21095=>"101101011",
  21096=>"011111001",
  21097=>"110100011",
  21098=>"000000111",
  21099=>"010001000",
  21100=>"001110101",
  21101=>"001111010",
  21102=>"111101000",
  21103=>"110010011",
  21104=>"110111110",
  21105=>"001001000",
  21106=>"000010001",
  21107=>"111100011",
  21108=>"001100110",
  21109=>"001001110",
  21110=>"000001100",
  21111=>"101010001",
  21112=>"111010111",
  21113=>"011111110",
  21114=>"110101010",
  21115=>"001001101",
  21116=>"110000010",
  21117=>"101100001",
  21118=>"110101110",
  21119=>"101100011",
  21120=>"111110110",
  21121=>"001110011",
  21122=>"010110000",
  21123=>"110000111",
  21124=>"100101111",
  21125=>"000100011",
  21126=>"110001111",
  21127=>"101101101",
  21128=>"011011011",
  21129=>"010100100",
  21130=>"111110001",
  21131=>"110000110",
  21132=>"100010100",
  21133=>"101011010",
  21134=>"010110011",
  21135=>"110111110",
  21136=>"101011011",
  21137=>"010100001",
  21138=>"001111010",
  21139=>"111011110",
  21140=>"010011100",
  21141=>"000010110",
  21142=>"010001010",
  21143=>"100110101",
  21144=>"100111010",
  21145=>"011001010",
  21146=>"100000000",
  21147=>"101010111",
  21148=>"110000000",
  21149=>"100001001",
  21150=>"111101111",
  21151=>"110011111",
  21152=>"011110111",
  21153=>"011001001",
  21154=>"011101110",
  21155=>"010011000",
  21156=>"100011000",
  21157=>"101000001",
  21158=>"101110101",
  21159=>"000001001",
  21160=>"001010011",
  21161=>"100010110",
  21162=>"010101001",
  21163=>"010111101",
  21164=>"101101110",
  21165=>"001000000",
  21166=>"011011010",
  21167=>"000001101",
  21168=>"000101110",
  21169=>"001111111",
  21170=>"010001000",
  21171=>"101111100",
  21172=>"111111100",
  21173=>"000100000",
  21174=>"011111100",
  21175=>"000111111",
  21176=>"100010110",
  21177=>"100100101",
  21178=>"010100110",
  21179=>"111100000",
  21180=>"010111010",
  21181=>"000000011",
  21182=>"010100110",
  21183=>"000110101",
  21184=>"010110010",
  21185=>"100011010",
  21186=>"000111000",
  21187=>"001110100",
  21188=>"000001110",
  21189=>"111001100",
  21190=>"001111100",
  21191=>"100000010",
  21192=>"110000100",
  21193=>"001001010",
  21194=>"000101000",
  21195=>"011110111",
  21196=>"010110010",
  21197=>"010110000",
  21198=>"011011101",
  21199=>"001100110",
  21200=>"111000010",
  21201=>"101000100",
  21202=>"101000000",
  21203=>"010100110",
  21204=>"110000101",
  21205=>"001000001",
  21206=>"111100111",
  21207=>"110010011",
  21208=>"101110110",
  21209=>"111001101",
  21210=>"111110101",
  21211=>"001110110",
  21212=>"111001011",
  21213=>"110111101",
  21214=>"101100000",
  21215=>"011011111",
  21216=>"101100111",
  21217=>"000010001",
  21218=>"011010011",
  21219=>"111111001",
  21220=>"111111111",
  21221=>"111101011",
  21222=>"011011100",
  21223=>"000001110",
  21224=>"100000001",
  21225=>"100100001",
  21226=>"101100010",
  21227=>"010000011",
  21228=>"010011000",
  21229=>"000100111",
  21230=>"101001100",
  21231=>"110100000",
  21232=>"011001011",
  21233=>"101001001",
  21234=>"111000111",
  21235=>"000000100",
  21236=>"111100110",
  21237=>"101100001",
  21238=>"001001010",
  21239=>"011110000",
  21240=>"100000110",
  21241=>"010110111",
  21242=>"010101011",
  21243=>"001110100",
  21244=>"011001100",
  21245=>"011100011",
  21246=>"001101001",
  21247=>"000100110",
  21248=>"010000000",
  21249=>"001000011",
  21250=>"001011000",
  21251=>"010001111",
  21252=>"111100110",
  21253=>"111011011",
  21254=>"110010000",
  21255=>"011101101",
  21256=>"111011001",
  21257=>"100110100",
  21258=>"100000101",
  21259=>"111011000",
  21260=>"100000000",
  21261=>"110111011",
  21262=>"010101001",
  21263=>"110000001",
  21264=>"101111011",
  21265=>"100110100",
  21266=>"111111111",
  21267=>"001011010",
  21268=>"011110000",
  21269=>"100100111",
  21270=>"011000101",
  21271=>"011111011",
  21272=>"110001001",
  21273=>"101100110",
  21274=>"001000011",
  21275=>"100010001",
  21276=>"111011000",
  21277=>"011110001",
  21278=>"100000110",
  21279=>"111011001",
  21280=>"101001011",
  21281=>"001101000",
  21282=>"101100111",
  21283=>"010010001",
  21284=>"100101011",
  21285=>"011001100",
  21286=>"100110010",
  21287=>"010110100",
  21288=>"000000101",
  21289=>"001000111",
  21290=>"100110001",
  21291=>"011110001",
  21292=>"011101111",
  21293=>"101000100",
  21294=>"001111101",
  21295=>"011110110",
  21296=>"001000011",
  21297=>"001101001",
  21298=>"101000011",
  21299=>"100111101",
  21300=>"001110100",
  21301=>"111010101",
  21302=>"111111111",
  21303=>"011101110",
  21304=>"101000000",
  21305=>"110010110",
  21306=>"110110010",
  21307=>"100101011",
  21308=>"101111001",
  21309=>"010101001",
  21310=>"001001000",
  21311=>"111000100",
  21312=>"101011110",
  21313=>"000011111",
  21314=>"100101100",
  21315=>"100001101",
  21316=>"111011001",
  21317=>"110100101",
  21318=>"111111011",
  21319=>"001000110",
  21320=>"110010001",
  21321=>"110000001",
  21322=>"101011110",
  21323=>"001000000",
  21324=>"011010110",
  21325=>"100011000",
  21326=>"000001010",
  21327=>"010000011",
  21328=>"001111001",
  21329=>"000100010",
  21330=>"110101010",
  21331=>"011001011",
  21332=>"011110010",
  21333=>"010010110",
  21334=>"010101011",
  21335=>"111010110",
  21336=>"010100111",
  21337=>"100011011",
  21338=>"011001001",
  21339=>"100100101",
  21340=>"100110000",
  21341=>"001011111",
  21342=>"000111010",
  21343=>"010100000",
  21344=>"101110010",
  21345=>"011010010",
  21346=>"011101000",
  21347=>"001111100",
  21348=>"000001001",
  21349=>"011000011",
  21350=>"010000000",
  21351=>"011111111",
  21352=>"110101011",
  21353=>"110000011",
  21354=>"111110100",
  21355=>"000010001",
  21356=>"110000010",
  21357=>"001111011",
  21358=>"111001010",
  21359=>"101000010",
  21360=>"010100000",
  21361=>"010011011",
  21362=>"001111000",
  21363=>"100010000",
  21364=>"111000000",
  21365=>"100110100",
  21366=>"010001000",
  21367=>"111011111",
  21368=>"010011110",
  21369=>"100001111",
  21370=>"000111101",
  21371=>"000001001",
  21372=>"100000011",
  21373=>"101100110",
  21374=>"110000001",
  21375=>"011111010",
  21376=>"100101011",
  21377=>"011001011",
  21378=>"100101101",
  21379=>"000110100",
  21380=>"010001010",
  21381=>"111101110",
  21382=>"000010100",
  21383=>"000000011",
  21384=>"110001110",
  21385=>"100101110",
  21386=>"011000001",
  21387=>"101000101",
  21388=>"000010001",
  21389=>"000000111",
  21390=>"101010001",
  21391=>"011101111",
  21392=>"101110111",
  21393=>"110000010",
  21394=>"110100111",
  21395=>"011100110",
  21396=>"001001010",
  21397=>"001011111",
  21398=>"000110111",
  21399=>"011001000",
  21400=>"000000101",
  21401=>"101001100",
  21402=>"000100000",
  21403=>"010010101",
  21404=>"001011110",
  21405=>"001111101",
  21406=>"010010100",
  21407=>"010000000",
  21408=>"011010111",
  21409=>"000111001",
  21410=>"010101011",
  21411=>"111101011",
  21412=>"100010001",
  21413=>"011011001",
  21414=>"111101111",
  21415=>"000111110",
  21416=>"100001001",
  21417=>"000001011",
  21418=>"101001110",
  21419=>"011101100",
  21420=>"111111110",
  21421=>"111100111",
  21422=>"010011000",
  21423=>"000001110",
  21424=>"010000000",
  21425=>"110001110",
  21426=>"111001011",
  21427=>"000100001",
  21428=>"010000010",
  21429=>"001010001",
  21430=>"110101000",
  21431=>"011110101",
  21432=>"111100011",
  21433=>"100010111",
  21434=>"010111001",
  21435=>"001011110",
  21436=>"001010001",
  21437=>"111010001",
  21438=>"100000110",
  21439=>"110100110",
  21440=>"100000001",
  21441=>"011001101",
  21442=>"000011011",
  21443=>"110011100",
  21444=>"100111010",
  21445=>"011111111",
  21446=>"101010011",
  21447=>"100001000",
  21448=>"010000111",
  21449=>"101001100",
  21450=>"010110010",
  21451=>"010101110",
  21452=>"001100000",
  21453=>"000000011",
  21454=>"101000010",
  21455=>"000001011",
  21456=>"000101110",
  21457=>"001001100",
  21458=>"101111110",
  21459=>"011001000",
  21460=>"000001001",
  21461=>"000010010",
  21462=>"101111111",
  21463=>"001000010",
  21464=>"011110001",
  21465=>"100111110",
  21466=>"001010001",
  21467=>"000100100",
  21468=>"100100010",
  21469=>"001011010",
  21470=>"010000101",
  21471=>"100000010",
  21472=>"111111010",
  21473=>"100011100",
  21474=>"011111110",
  21475=>"000110001",
  21476=>"101000010",
  21477=>"011001100",
  21478=>"100110001",
  21479=>"010011011",
  21480=>"010101111",
  21481=>"001100101",
  21482=>"001110001",
  21483=>"000010000",
  21484=>"101111011",
  21485=>"101000001",
  21486=>"011010101",
  21487=>"010101110",
  21488=>"101100010",
  21489=>"111100101",
  21490=>"001001111",
  21491=>"001100110",
  21492=>"101001101",
  21493=>"000110101",
  21494=>"010001101",
  21495=>"111110110",
  21496=>"011011011",
  21497=>"101011110",
  21498=>"000011010",
  21499=>"001001010",
  21500=>"111101010",
  21501=>"000010010",
  21502=>"000010101",
  21503=>"110110111",
  21504=>"000000001",
  21505=>"110010001",
  21506=>"110111110",
  21507=>"101000000",
  21508=>"111110000",
  21509=>"010000110",
  21510=>"010011000",
  21511=>"111111000",
  21512=>"010011100",
  21513=>"010001000",
  21514=>"101110111",
  21515=>"100101011",
  21516=>"110101111",
  21517=>"110000100",
  21518=>"010011000",
  21519=>"000001001",
  21520=>"100111100",
  21521=>"011001100",
  21522=>"001110111",
  21523=>"011010100",
  21524=>"010100010",
  21525=>"000001000",
  21526=>"011100101",
  21527=>"010000011",
  21528=>"000100111",
  21529=>"011010010",
  21530=>"110110100",
  21531=>"100010101",
  21532=>"100110100",
  21533=>"010101001",
  21534=>"011010001",
  21535=>"000001110",
  21536=>"100000000",
  21537=>"101101010",
  21538=>"101101110",
  21539=>"101100100",
  21540=>"101000111",
  21541=>"101111101",
  21542=>"101010010",
  21543=>"001101100",
  21544=>"100100000",
  21545=>"110001001",
  21546=>"010111011",
  21547=>"000010001",
  21548=>"001001000",
  21549=>"001110000",
  21550=>"011101110",
  21551=>"010101111",
  21552=>"101000101",
  21553=>"101000000",
  21554=>"001100001",
  21555=>"001111100",
  21556=>"010111101",
  21557=>"000110110",
  21558=>"001000101",
  21559=>"111101111",
  21560=>"001011110",
  21561=>"100010011",
  21562=>"111001011",
  21563=>"010011110",
  21564=>"100011100",
  21565=>"000111000",
  21566=>"010111010",
  21567=>"011101101",
  21568=>"000110111",
  21569=>"011100001",
  21570=>"001010000",
  21571=>"111000011",
  21572=>"101011011",
  21573=>"001010101",
  21574=>"000110100",
  21575=>"111111000",
  21576=>"100111011",
  21577=>"111001111",
  21578=>"101000100",
  21579=>"111011001",
  21580=>"011100011",
  21581=>"000100100",
  21582=>"101011110",
  21583=>"001000101",
  21584=>"000101001",
  21585=>"010010111",
  21586=>"001010111",
  21587=>"010111010",
  21588=>"010000000",
  21589=>"100101000",
  21590=>"010111011",
  21591=>"000000001",
  21592=>"111000000",
  21593=>"000010011",
  21594=>"001101000",
  21595=>"001111100",
  21596=>"000010100",
  21597=>"110110010",
  21598=>"000010000",
  21599=>"100100101",
  21600=>"111110100",
  21601=>"110001010",
  21602=>"111010011",
  21603=>"011001010",
  21604=>"111110000",
  21605=>"110000001",
  21606=>"001010011",
  21607=>"111010111",
  21608=>"100000011",
  21609=>"010000000",
  21610=>"101001100",
  21611=>"011010001",
  21612=>"111110000",
  21613=>"101110100",
  21614=>"011101000",
  21615=>"010011100",
  21616=>"011111111",
  21617=>"101011000",
  21618=>"000110000",
  21619=>"111101010",
  21620=>"011110011",
  21621=>"010001101",
  21622=>"011111111",
  21623=>"011010011",
  21624=>"000100010",
  21625=>"101010101",
  21626=>"000110010",
  21627=>"001100010",
  21628=>"010111111",
  21629=>"001010111",
  21630=>"101011011",
  21631=>"011011111",
  21632=>"000110100",
  21633=>"011110101",
  21634=>"000001011",
  21635=>"001101011",
  21636=>"001011111",
  21637=>"100110110",
  21638=>"101101010",
  21639=>"010111100",
  21640=>"111110101",
  21641=>"101101110",
  21642=>"001101101",
  21643=>"111101011",
  21644=>"100000011",
  21645=>"111100111",
  21646=>"001010101",
  21647=>"001110110",
  21648=>"100010110",
  21649=>"011100000",
  21650=>"111101010",
  21651=>"111100010",
  21652=>"000001011",
  21653=>"110111101",
  21654=>"001011110",
  21655=>"001110100",
  21656=>"001001010",
  21657=>"001010010",
  21658=>"111110101",
  21659=>"100001011",
  21660=>"001011010",
  21661=>"011010001",
  21662=>"100000111",
  21663=>"001000011",
  21664=>"000110000",
  21665=>"100101111",
  21666=>"000000111",
  21667=>"010100001",
  21668=>"111101000",
  21669=>"111110000",
  21670=>"110001110",
  21671=>"001000111",
  21672=>"001101111",
  21673=>"101011001",
  21674=>"011010101",
  21675=>"010010011",
  21676=>"000111101",
  21677=>"101001011",
  21678=>"111111100",
  21679=>"110010110",
  21680=>"000101110",
  21681=>"011100110",
  21682=>"011110100",
  21683=>"011100100",
  21684=>"111110001",
  21685=>"011101010",
  21686=>"110110001",
  21687=>"101101010",
  21688=>"110110110",
  21689=>"011111000",
  21690=>"001010010",
  21691=>"100100111",
  21692=>"010000010",
  21693=>"111000001",
  21694=>"001101111",
  21695=>"011110010",
  21696=>"110110110",
  21697=>"111101010",
  21698=>"011100011",
  21699=>"100010011",
  21700=>"011100001",
  21701=>"010010111",
  21702=>"011111111",
  21703=>"010000101",
  21704=>"010111001",
  21705=>"100100010",
  21706=>"011111010",
  21707=>"110111111",
  21708=>"101111100",
  21709=>"011000000",
  21710=>"110101111",
  21711=>"110001010",
  21712=>"010000100",
  21713=>"011100011",
  21714=>"010110111",
  21715=>"001000000",
  21716=>"001100100",
  21717=>"100100001",
  21718=>"101000010",
  21719=>"111001010",
  21720=>"100000100",
  21721=>"101111111",
  21722=>"100001101",
  21723=>"111100001",
  21724=>"111000101",
  21725=>"000001101",
  21726=>"000000010",
  21727=>"111011010",
  21728=>"101010100",
  21729=>"001010000",
  21730=>"100010001",
  21731=>"100011101",
  21732=>"101011010",
  21733=>"110011000",
  21734=>"001100001",
  21735=>"110010101",
  21736=>"101111010",
  21737=>"010101000",
  21738=>"010000100",
  21739=>"110110100",
  21740=>"011011000",
  21741=>"010001100",
  21742=>"110001000",
  21743=>"111010000",
  21744=>"011011111",
  21745=>"111111110",
  21746=>"010110000",
  21747=>"111010000",
  21748=>"100111100",
  21749=>"001111010",
  21750=>"101001101",
  21751=>"000000001",
  21752=>"100011101",
  21753=>"111011011",
  21754=>"010111100",
  21755=>"000101001",
  21756=>"000000101",
  21757=>"001000000",
  21758=>"010001001",
  21759=>"010000000",
  21760=>"111101000",
  21761=>"101000110",
  21762=>"101111110",
  21763=>"000111001",
  21764=>"110010000",
  21765=>"011110111",
  21766=>"000101111",
  21767=>"110110001",
  21768=>"001111000",
  21769=>"111101110",
  21770=>"010010011",
  21771=>"110001010",
  21772=>"100000010",
  21773=>"001011110",
  21774=>"100111111",
  21775=>"011010100",
  21776=>"110111110",
  21777=>"100010001",
  21778=>"100100110",
  21779=>"100100110",
  21780=>"010101011",
  21781=>"010010111",
  21782=>"100111001",
  21783=>"111100001",
  21784=>"101011010",
  21785=>"101001001",
  21786=>"001110000",
  21787=>"101001001",
  21788=>"010101011",
  21789=>"101111000",
  21790=>"101111000",
  21791=>"000110000",
  21792=>"010110101",
  21793=>"000101001",
  21794=>"010010010",
  21795=>"100101001",
  21796=>"000001110",
  21797=>"100000100",
  21798=>"110000001",
  21799=>"001011110",
  21800=>"011000101",
  21801=>"010011111",
  21802=>"000001111",
  21803=>"100111001",
  21804=>"000000001",
  21805=>"001000011",
  21806=>"001101001",
  21807=>"001011011",
  21808=>"100000000",
  21809=>"001010100",
  21810=>"110010010",
  21811=>"100110001",
  21812=>"010101011",
  21813=>"000001110",
  21814=>"000001110",
  21815=>"100000011",
  21816=>"011100101",
  21817=>"001101011",
  21818=>"000101111",
  21819=>"100100000",
  21820=>"011000100",
  21821=>"110011111",
  21822=>"000010100",
  21823=>"110000001",
  21824=>"011100110",
  21825=>"001111111",
  21826=>"100000111",
  21827=>"101111010",
  21828=>"101001000",
  21829=>"010101010",
  21830=>"000100110",
  21831=>"001010001",
  21832=>"111010101",
  21833=>"010100101",
  21834=>"000011010",
  21835=>"001110110",
  21836=>"101101000",
  21837=>"100000011",
  21838=>"111011111",
  21839=>"010010011",
  21840=>"110110001",
  21841=>"110100011",
  21842=>"000100010",
  21843=>"001001100",
  21844=>"000111000",
  21845=>"011001110",
  21846=>"101101110",
  21847=>"101010101",
  21848=>"000000000",
  21849=>"110100100",
  21850=>"010011010",
  21851=>"110110101",
  21852=>"000000011",
  21853=>"111011100",
  21854=>"010011111",
  21855=>"100101111",
  21856=>"111110010",
  21857=>"100011011",
  21858=>"100100111",
  21859=>"000000011",
  21860=>"100100000",
  21861=>"110110110",
  21862=>"001110101",
  21863=>"101101000",
  21864=>"000000111",
  21865=>"101000000",
  21866=>"110110010",
  21867=>"010001101",
  21868=>"100101010",
  21869=>"111000110",
  21870=>"101011111",
  21871=>"110000111",
  21872=>"001101111",
  21873=>"011001011",
  21874=>"110111001",
  21875=>"111101110",
  21876=>"111010000",
  21877=>"001000100",
  21878=>"010011111",
  21879=>"110100111",
  21880=>"010011000",
  21881=>"001000010",
  21882=>"001100001",
  21883=>"011000000",
  21884=>"001111100",
  21885=>"111110110",
  21886=>"000100000",
  21887=>"111000000",
  21888=>"100010010",
  21889=>"000110111",
  21890=>"100000100",
  21891=>"011011111",
  21892=>"011100100",
  21893=>"110000001",
  21894=>"000111110",
  21895=>"111100110",
  21896=>"111101110",
  21897=>"011100011",
  21898=>"100110100",
  21899=>"111100000",
  21900=>"011000011",
  21901=>"010110100",
  21902=>"110101111",
  21903=>"000000110",
  21904=>"010110010",
  21905=>"100111010",
  21906=>"010110100",
  21907=>"011100000",
  21908=>"001111111",
  21909=>"111010000",
  21910=>"100110010",
  21911=>"101011000",
  21912=>"000101001",
  21913=>"100100101",
  21914=>"100001000",
  21915=>"000010000",
  21916=>"110101110",
  21917=>"000101001",
  21918=>"011010000",
  21919=>"000111010",
  21920=>"011010100",
  21921=>"110010001",
  21922=>"100100000",
  21923=>"001010010",
  21924=>"010100010",
  21925=>"000101111",
  21926=>"001010011",
  21927=>"111100011",
  21928=>"111101010",
  21929=>"110110001",
  21930=>"010000001",
  21931=>"101101011",
  21932=>"011011001",
  21933=>"101111110",
  21934=>"000010000",
  21935=>"110100011",
  21936=>"001100110",
  21937=>"111101000",
  21938=>"011111101",
  21939=>"000011000",
  21940=>"011000010",
  21941=>"101000101",
  21942=>"011101010",
  21943=>"011001000",
  21944=>"111001000",
  21945=>"000000010",
  21946=>"000001011",
  21947=>"100111110",
  21948=>"100110001",
  21949=>"110111101",
  21950=>"101011000",
  21951=>"000011000",
  21952=>"011101011",
  21953=>"100011010",
  21954=>"101100101",
  21955=>"000101010",
  21956=>"110101010",
  21957=>"101000000",
  21958=>"001010000",
  21959=>"000001110",
  21960=>"001011011",
  21961=>"100001000",
  21962=>"010111111",
  21963=>"111011111",
  21964=>"000011101",
  21965=>"010011101",
  21966=>"100011010",
  21967=>"000001100",
  21968=>"011011001",
  21969=>"111000111",
  21970=>"101001000",
  21971=>"000100000",
  21972=>"111100111",
  21973=>"100010111",
  21974=>"011011101",
  21975=>"010110010",
  21976=>"001100011",
  21977=>"111110101",
  21978=>"110001110",
  21979=>"110000010",
  21980=>"001000000",
  21981=>"110111110",
  21982=>"000001110",
  21983=>"100110101",
  21984=>"011101010",
  21985=>"001010001",
  21986=>"111111111",
  21987=>"111110000",
  21988=>"100000110",
  21989=>"000010001",
  21990=>"001100110",
  21991=>"110010010",
  21992=>"011100100",
  21993=>"010000101",
  21994=>"010000000",
  21995=>"010000010",
  21996=>"010000101",
  21997=>"001001110",
  21998=>"101100101",
  21999=>"101010101",
  22000=>"011001010",
  22001=>"111001001",
  22002=>"100101000",
  22003=>"101010011",
  22004=>"101110001",
  22005=>"001110000",
  22006=>"101001111",
  22007=>"000000010",
  22008=>"111011000",
  22009=>"000011000",
  22010=>"111001100",
  22011=>"011110001",
  22012=>"100000000",
  22013=>"101100011",
  22014=>"011001111",
  22015=>"101110110",
  22016=>"010000111",
  22017=>"001101101",
  22018=>"101111101",
  22019=>"111110100",
  22020=>"101011000",
  22021=>"100010100",
  22022=>"111001001",
  22023=>"001110101",
  22024=>"001100011",
  22025=>"101000101",
  22026=>"111010101",
  22027=>"011100000",
  22028=>"101010100",
  22029=>"010111111",
  22030=>"100001000",
  22031=>"000100110",
  22032=>"111110011",
  22033=>"000101110",
  22034=>"100011110",
  22035=>"001110110",
  22036=>"001000111",
  22037=>"000100110",
  22038=>"101101010",
  22039=>"110100100",
  22040=>"010101110",
  22041=>"111111010",
  22042=>"000101100",
  22043=>"111011011",
  22044=>"110110010",
  22045=>"000100100",
  22046=>"101000100",
  22047=>"101100000",
  22048=>"111001001",
  22049=>"101111001",
  22050=>"111110000",
  22051=>"110001100",
  22052=>"110110010",
  22053=>"000110111",
  22054=>"101001001",
  22055=>"110111111",
  22056=>"010000100",
  22057=>"111110110",
  22058=>"100000000",
  22059=>"000101111",
  22060=>"011101101",
  22061=>"110011001",
  22062=>"101100011",
  22063=>"011000101",
  22064=>"110011111",
  22065=>"101101010",
  22066=>"110101000",
  22067=>"100100001",
  22068=>"111010010",
  22069=>"010001000",
  22070=>"010011111",
  22071=>"010010000",
  22072=>"011111110",
  22073=>"111010000",
  22074=>"101101100",
  22075=>"111010001",
  22076=>"100000101",
  22077=>"000010001",
  22078=>"100101001",
  22079=>"000001011",
  22080=>"001001011",
  22081=>"110010100",
  22082=>"100111011",
  22083=>"100000001",
  22084=>"001010000",
  22085=>"000011110",
  22086=>"010011000",
  22087=>"101101011",
  22088=>"101100010",
  22089=>"011101000",
  22090=>"111110111",
  22091=>"111001000",
  22092=>"010101111",
  22093=>"000111110",
  22094=>"101110001",
  22095=>"110001011",
  22096=>"101110111",
  22097=>"111101111",
  22098=>"100010000",
  22099=>"100001010",
  22100=>"000000101",
  22101=>"100000100",
  22102=>"000111001",
  22103=>"000111011",
  22104=>"110111100",
  22105=>"100111101",
  22106=>"010111000",
  22107=>"111111010",
  22108=>"100100001",
  22109=>"000000001",
  22110=>"100100101",
  22111=>"001111111",
  22112=>"000001101",
  22113=>"100101011",
  22114=>"010110000",
  22115=>"100111001",
  22116=>"000011011",
  22117=>"011110111",
  22118=>"000001110",
  22119=>"010101100",
  22120=>"000000110",
  22121=>"101110000",
  22122=>"111011111",
  22123=>"011001101",
  22124=>"001101110",
  22125=>"101100100",
  22126=>"100111010",
  22127=>"100111001",
  22128=>"101101101",
  22129=>"110000000",
  22130=>"001011111",
  22131=>"010100000",
  22132=>"010010011",
  22133=>"100110010",
  22134=>"111010111",
  22135=>"111011100",
  22136=>"100100010",
  22137=>"000111011",
  22138=>"101010010",
  22139=>"000001000",
  22140=>"001011001",
  22141=>"010000111",
  22142=>"001000000",
  22143=>"111110001",
  22144=>"100001010",
  22145=>"111011111",
  22146=>"000001011",
  22147=>"011000011",
  22148=>"111010111",
  22149=>"101001100",
  22150=>"000000101",
  22151=>"011011111",
  22152=>"110100011",
  22153=>"001010011",
  22154=>"110000101",
  22155=>"101111011",
  22156=>"011110101",
  22157=>"111101101",
  22158=>"110100100",
  22159=>"001000100",
  22160=>"001000110",
  22161=>"110110111",
  22162=>"001100111",
  22163=>"100001001",
  22164=>"011100011",
  22165=>"010100111",
  22166=>"100101100",
  22167=>"001010100",
  22168=>"111111101",
  22169=>"011111101",
  22170=>"100110110",
  22171=>"011100011",
  22172=>"000011101",
  22173=>"101100000",
  22174=>"001010001",
  22175=>"001000000",
  22176=>"011101111",
  22177=>"101110100",
  22178=>"001010011",
  22179=>"110111011",
  22180=>"101111110",
  22181=>"010001011",
  22182=>"110010000",
  22183=>"001100010",
  22184=>"001100011",
  22185=>"000110000",
  22186=>"110011010",
  22187=>"000000001",
  22188=>"100101011",
  22189=>"000011101",
  22190=>"110110101",
  22191=>"001000111",
  22192=>"110000110",
  22193=>"011000001",
  22194=>"100110111",
  22195=>"110110001",
  22196=>"011100111",
  22197=>"110010100",
  22198=>"111010100",
  22199=>"000110010",
  22200=>"100010101",
  22201=>"010110000",
  22202=>"101100010",
  22203=>"001110000",
  22204=>"001010111",
  22205=>"110000100",
  22206=>"000001000",
  22207=>"111000000",
  22208=>"111110110",
  22209=>"100000111",
  22210=>"001011011",
  22211=>"100011101",
  22212=>"001000100",
  22213=>"110100011",
  22214=>"100110110",
  22215=>"110110000",
  22216=>"011001101",
  22217=>"110100100",
  22218=>"010011101",
  22219=>"101001000",
  22220=>"100110011",
  22221=>"101011010",
  22222=>"001001010",
  22223=>"110110010",
  22224=>"001000101",
  22225=>"111001100",
  22226=>"101101001",
  22227=>"100010111",
  22228=>"010100010",
  22229=>"111000100",
  22230=>"011011011",
  22231=>"111010011",
  22232=>"111010010",
  22233=>"001010110",
  22234=>"001001111",
  22235=>"010001101",
  22236=>"101110101",
  22237=>"011000011",
  22238=>"000111111",
  22239=>"110111001",
  22240=>"001010001",
  22241=>"000110101",
  22242=>"101100110",
  22243=>"111010011",
  22244=>"010001101",
  22245=>"110111101",
  22246=>"101110100",
  22247=>"111111100",
  22248=>"000010011",
  22249=>"011100011",
  22250=>"100101100",
  22251=>"011000010",
  22252=>"000000001",
  22253=>"010001110",
  22254=>"100010011",
  22255=>"001010100",
  22256=>"101110111",
  22257=>"100100101",
  22258=>"001000110",
  22259=>"011111110",
  22260=>"101010000",
  22261=>"011000000",
  22262=>"100111001",
  22263=>"111011110",
  22264=>"000010101",
  22265=>"011101101",
  22266=>"100001101",
  22267=>"000101000",
  22268=>"100011000",
  22269=>"000010001",
  22270=>"010000001",
  22271=>"000100000",
  22272=>"001011111",
  22273=>"001001111",
  22274=>"111101101",
  22275=>"101010101",
  22276=>"111101011",
  22277=>"110110001",
  22278=>"101110110",
  22279=>"110100011",
  22280=>"000010111",
  22281=>"011101000",
  22282=>"011011111",
  22283=>"001001011",
  22284=>"000000000",
  22285=>"100000011",
  22286=>"100110001",
  22287=>"110101100",
  22288=>"011011110",
  22289=>"101010100",
  22290=>"001110010",
  22291=>"111000110",
  22292=>"100010010",
  22293=>"000001100",
  22294=>"101101001",
  22295=>"111111101",
  22296=>"110111110",
  22297=>"110000001",
  22298=>"100100111",
  22299=>"100101111",
  22300=>"000100101",
  22301=>"100101111",
  22302=>"100101111",
  22303=>"001011011",
  22304=>"000000000",
  22305=>"100100010",
  22306=>"101111000",
  22307=>"010011010",
  22308=>"100101011",
  22309=>"011110100",
  22310=>"010101101",
  22311=>"111111011",
  22312=>"010100110",
  22313=>"000111101",
  22314=>"001000010",
  22315=>"010100010",
  22316=>"100111011",
  22317=>"011100101",
  22318=>"000110100",
  22319=>"111001001",
  22320=>"010110011",
  22321=>"110000111",
  22322=>"110111110",
  22323=>"100000000",
  22324=>"110001110",
  22325=>"010101000",
  22326=>"000010101",
  22327=>"011011001",
  22328=>"011010010",
  22329=>"011110000",
  22330=>"101001010",
  22331=>"100000111",
  22332=>"000101001",
  22333=>"001010000",
  22334=>"001000111",
  22335=>"111110000",
  22336=>"110010010",
  22337=>"100000011",
  22338=>"110101111",
  22339=>"101111101",
  22340=>"000101101",
  22341=>"111110100",
  22342=>"110010001",
  22343=>"000111001",
  22344=>"111111010",
  22345=>"001101110",
  22346=>"000100001",
  22347=>"101111001",
  22348=>"010001010",
  22349=>"111011110",
  22350=>"100011011",
  22351=>"100101110",
  22352=>"000001001",
  22353=>"001001111",
  22354=>"100010001",
  22355=>"010001010",
  22356=>"010001011",
  22357=>"111111111",
  22358=>"011101011",
  22359=>"100100010",
  22360=>"011000101",
  22361=>"100010001",
  22362=>"110000101",
  22363=>"100110100",
  22364=>"101101111",
  22365=>"010111000",
  22366=>"111010110",
  22367=>"010011000",
  22368=>"000000101",
  22369=>"101111010",
  22370=>"011100010",
  22371=>"101010101",
  22372=>"111010010",
  22373=>"011001000",
  22374=>"100000001",
  22375=>"001111000",
  22376=>"001000100",
  22377=>"010101111",
  22378=>"110001010",
  22379=>"011010010",
  22380=>"000111100",
  22381=>"011001111",
  22382=>"101000000",
  22383=>"111000111",
  22384=>"010001010",
  22385=>"010000110",
  22386=>"110101111",
  22387=>"111111101",
  22388=>"000100001",
  22389=>"001101101",
  22390=>"011010011",
  22391=>"100101000",
  22392=>"101111100",
  22393=>"000110100",
  22394=>"101110110",
  22395=>"000001010",
  22396=>"011010111",
  22397=>"001000010",
  22398=>"111101011",
  22399=>"011110101",
  22400=>"001001001",
  22401=>"011010010",
  22402=>"111101111",
  22403=>"100100010",
  22404=>"001000110",
  22405=>"011111011",
  22406=>"111001000",
  22407=>"011111000",
  22408=>"101001011",
  22409=>"000110111",
  22410=>"010010000",
  22411=>"101001001",
  22412=>"110011001",
  22413=>"110101101",
  22414=>"100000000",
  22415=>"000101000",
  22416=>"111001011",
  22417=>"001100000",
  22418=>"010011010",
  22419=>"001010011",
  22420=>"000011000",
  22421=>"011001001",
  22422=>"000000100",
  22423=>"101011110",
  22424=>"111011011",
  22425=>"111110111",
  22426=>"111000100",
  22427=>"001000010",
  22428=>"010011100",
  22429=>"000111111",
  22430=>"010000010",
  22431=>"111111111",
  22432=>"001110010",
  22433=>"101101111",
  22434=>"011010001",
  22435=>"011111110",
  22436=>"111010100",
  22437=>"110101010",
  22438=>"110011111",
  22439=>"001100101",
  22440=>"101011011",
  22441=>"111101111",
  22442=>"001011010",
  22443=>"001010101",
  22444=>"100111001",
  22445=>"010001110",
  22446=>"111100001",
  22447=>"100010000",
  22448=>"100101010",
  22449=>"101011101",
  22450=>"101101101",
  22451=>"000001100",
  22452=>"111101001",
  22453=>"110110011",
  22454=>"000010011",
  22455=>"001010001",
  22456=>"110011100",
  22457=>"111000101",
  22458=>"011110111",
  22459=>"010011101",
  22460=>"111101001",
  22461=>"110100000",
  22462=>"111001101",
  22463=>"011110110",
  22464=>"100000010",
  22465=>"000000000",
  22466=>"111000000",
  22467=>"001011001",
  22468=>"111010110",
  22469=>"001001011",
  22470=>"010000100",
  22471=>"101010000",
  22472=>"000100000",
  22473=>"011111001",
  22474=>"110110100",
  22475=>"111111101",
  22476=>"011110011",
  22477=>"111111111",
  22478=>"101110011",
  22479=>"011110000",
  22480=>"001011001",
  22481=>"001100101",
  22482=>"111111110",
  22483=>"000000111",
  22484=>"000010000",
  22485=>"111110010",
  22486=>"111001100",
  22487=>"101100101",
  22488=>"010100010",
  22489=>"100110110",
  22490=>"111100111",
  22491=>"000011011",
  22492=>"101101001",
  22493=>"110101011",
  22494=>"111100100",
  22495=>"001010010",
  22496=>"100010110",
  22497=>"110101111",
  22498=>"111010000",
  22499=>"001100011",
  22500=>"001010110",
  22501=>"000000001",
  22502=>"000111111",
  22503=>"110111110",
  22504=>"100011111",
  22505=>"101010100",
  22506=>"000011101",
  22507=>"010010111",
  22508=>"001101111",
  22509=>"000100001",
  22510=>"100010110",
  22511=>"101100000",
  22512=>"010011001",
  22513=>"010000101",
  22514=>"001010011",
  22515=>"000101100",
  22516=>"011000000",
  22517=>"000010010",
  22518=>"101101101",
  22519=>"000111110",
  22520=>"011110101",
  22521=>"101111100",
  22522=>"010101010",
  22523=>"001011100",
  22524=>"100101011",
  22525=>"011101101",
  22526=>"001101100",
  22527=>"000100010",
  22528=>"001100000",
  22529=>"110011001",
  22530=>"110000101",
  22531=>"011100011",
  22532=>"111101010",
  22533=>"011010001",
  22534=>"100101011",
  22535=>"011001100",
  22536=>"111100001",
  22537=>"110111111",
  22538=>"101010011",
  22539=>"011010011",
  22540=>"100110000",
  22541=>"000010111",
  22542=>"001101111",
  22543=>"100110001",
  22544=>"111101001",
  22545=>"000000010",
  22546=>"011101101",
  22547=>"110101101",
  22548=>"000111011",
  22549=>"101100011",
  22550=>"010010010",
  22551=>"011001110",
  22552=>"000110111",
  22553=>"101111110",
  22554=>"001001111",
  22555=>"111011111",
  22556=>"000011111",
  22557=>"001111010",
  22558=>"110111000",
  22559=>"101010011",
  22560=>"111101010",
  22561=>"100010011",
  22562=>"100000001",
  22563=>"011011101",
  22564=>"001101001",
  22565=>"010010111",
  22566=>"101101000",
  22567=>"010101000",
  22568=>"101000001",
  22569=>"010100101",
  22570=>"110100010",
  22571=>"101011101",
  22572=>"100110011",
  22573=>"100011010",
  22574=>"111100001",
  22575=>"000000010",
  22576=>"111101111",
  22577=>"110100001",
  22578=>"000011001",
  22579=>"110101010",
  22580=>"111111001",
  22581=>"001011001",
  22582=>"111001100",
  22583=>"111110110",
  22584=>"000010111",
  22585=>"100101010",
  22586=>"000001011",
  22587=>"010010110",
  22588=>"011010000",
  22589=>"110110010",
  22590=>"110100111",
  22591=>"011111010",
  22592=>"111010011",
  22593=>"111010101",
  22594=>"100110101",
  22595=>"011101000",
  22596=>"010000110",
  22597=>"111011111",
  22598=>"101010001",
  22599=>"110010001",
  22600=>"000101011",
  22601=>"110101010",
  22602=>"001110010",
  22603=>"101111000",
  22604=>"001100111",
  22605=>"111111110",
  22606=>"110000100",
  22607=>"000001011",
  22608=>"001010110",
  22609=>"101001111",
  22610=>"110100010",
  22611=>"111100100",
  22612=>"001011000",
  22613=>"101100110",
  22614=>"111010111",
  22615=>"011010000",
  22616=>"000111011",
  22617=>"000000001",
  22618=>"100010100",
  22619=>"100110100",
  22620=>"010011001",
  22621=>"110110010",
  22622=>"010011111",
  22623=>"111111000",
  22624=>"100000111",
  22625=>"010011101",
  22626=>"000111100",
  22627=>"000000000",
  22628=>"100011011",
  22629=>"010110010",
  22630=>"100110010",
  22631=>"111000010",
  22632=>"110101100",
  22633=>"001010110",
  22634=>"101100100",
  22635=>"011011100",
  22636=>"110001000",
  22637=>"110110001",
  22638=>"100010011",
  22639=>"010001110",
  22640=>"110100010",
  22641=>"100000110",
  22642=>"001100101",
  22643=>"100111010",
  22644=>"010001000",
  22645=>"111101100",
  22646=>"111111010",
  22647=>"000001110",
  22648=>"100000000",
  22649=>"100100100",
  22650=>"001110011",
  22651=>"000011101",
  22652=>"000000100",
  22653=>"101000010",
  22654=>"010110000",
  22655=>"000101100",
  22656=>"001111100",
  22657=>"101000011",
  22658=>"100000000",
  22659=>"100001101",
  22660=>"111001001",
  22661=>"001000001",
  22662=>"011100000",
  22663=>"000010110",
  22664=>"010001001",
  22665=>"011000110",
  22666=>"111001111",
  22667=>"011001110",
  22668=>"010010010",
  22669=>"111011110",
  22670=>"111110101",
  22671=>"010001100",
  22672=>"100000001",
  22673=>"101010110",
  22674=>"011100101",
  22675=>"000011001",
  22676=>"100100000",
  22677=>"101001111",
  22678=>"000100000",
  22679=>"101111101",
  22680=>"110010110",
  22681=>"110111111",
  22682=>"011101101",
  22683=>"110111110",
  22684=>"010111101",
  22685=>"000011000",
  22686=>"100110110",
  22687=>"000101111",
  22688=>"111000111",
  22689=>"101100011",
  22690=>"110111110",
  22691=>"110001111",
  22692=>"010101110",
  22693=>"111011110",
  22694=>"000101100",
  22695=>"011001011",
  22696=>"011001011",
  22697=>"110001010",
  22698=>"000010010",
  22699=>"101010111",
  22700=>"101101000",
  22701=>"010011000",
  22702=>"000001000",
  22703=>"100011001",
  22704=>"000111111",
  22705=>"011100111",
  22706=>"011001110",
  22707=>"011100011",
  22708=>"000110100",
  22709=>"000111010",
  22710=>"100010110",
  22711=>"011110111",
  22712=>"011001111",
  22713=>"000010001",
  22714=>"000101001",
  22715=>"111001011",
  22716=>"000111110",
  22717=>"101011000",
  22718=>"100010011",
  22719=>"001000000",
  22720=>"110000010",
  22721=>"001001100",
  22722=>"100011001",
  22723=>"011000001",
  22724=>"101000111",
  22725=>"001110000",
  22726=>"100111101",
  22727=>"111111111",
  22728=>"001011010",
  22729=>"111111001",
  22730=>"011111010",
  22731=>"100101011",
  22732=>"100010010",
  22733=>"011100110",
  22734=>"000010111",
  22735=>"100000010",
  22736=>"110100010",
  22737=>"100110010",
  22738=>"001110001",
  22739=>"011111111",
  22740=>"010011000",
  22741=>"011100101",
  22742=>"100001100",
  22743=>"011101100",
  22744=>"011100111",
  22745=>"000101100",
  22746=>"000100110",
  22747=>"001111001",
  22748=>"111011101",
  22749=>"110111101",
  22750=>"100011100",
  22751=>"010000110",
  22752=>"100110011",
  22753=>"100011011",
  22754=>"011001110",
  22755=>"101110110",
  22756=>"011111001",
  22757=>"010110110",
  22758=>"110100010",
  22759=>"110110011",
  22760=>"010101000",
  22761=>"000010100",
  22762=>"010101111",
  22763=>"000010011",
  22764=>"111011110",
  22765=>"110010000",
  22766=>"010111010",
  22767=>"001001000",
  22768=>"101001110",
  22769=>"101100001",
  22770=>"101111111",
  22771=>"110010111",
  22772=>"000110011",
  22773=>"011000101",
  22774=>"101110111",
  22775=>"110000100",
  22776=>"111010101",
  22777=>"011010110",
  22778=>"100000111",
  22779=>"001010000",
  22780=>"110100101",
  22781=>"010101110",
  22782=>"110011101",
  22783=>"000000000",
  22784=>"001010101",
  22785=>"110101001",
  22786=>"101010111",
  22787=>"000100000",
  22788=>"111010110",
  22789=>"001100111",
  22790=>"001010011",
  22791=>"011010110",
  22792=>"111011010",
  22793=>"001000010",
  22794=>"001101010",
  22795=>"000001111",
  22796=>"010001000",
  22797=>"101111100",
  22798=>"111111000",
  22799=>"010100011",
  22800=>"001010010",
  22801=>"011111011",
  22802=>"000000101",
  22803=>"001101110",
  22804=>"111010100",
  22805=>"010100010",
  22806=>"011011100",
  22807=>"111110110",
  22808=>"010001010",
  22809=>"010111111",
  22810=>"011100000",
  22811=>"100001111",
  22812=>"110000001",
  22813=>"011111000",
  22814=>"100100111",
  22815=>"110100111",
  22816=>"010010110",
  22817=>"000010110",
  22818=>"010101000",
  22819=>"110000000",
  22820=>"101010101",
  22821=>"101000100",
  22822=>"000100011",
  22823=>"011100101",
  22824=>"010010010",
  22825=>"101010000",
  22826=>"111011001",
  22827=>"010100001",
  22828=>"011110011",
  22829=>"010101010",
  22830=>"010001010",
  22831=>"111000011",
  22832=>"010100001",
  22833=>"011101101",
  22834=>"111101001",
  22835=>"110010011",
  22836=>"101101101",
  22837=>"101011111",
  22838=>"000010111",
  22839=>"011111000",
  22840=>"100110110",
  22841=>"011011010",
  22842=>"110101100",
  22843=>"011111110",
  22844=>"110101100",
  22845=>"011101110",
  22846=>"100011101",
  22847=>"111010011",
  22848=>"101100111",
  22849=>"110100001",
  22850=>"101101000",
  22851=>"111011001",
  22852=>"001000101",
  22853=>"101100011",
  22854=>"110001110",
  22855=>"111100111",
  22856=>"000111101",
  22857=>"010111010",
  22858=>"111001010",
  22859=>"001111011",
  22860=>"010111010",
  22861=>"010111001",
  22862=>"001110011",
  22863=>"000101111",
  22864=>"100110100",
  22865=>"011000011",
  22866=>"000001111",
  22867=>"011000111",
  22868=>"000011000",
  22869=>"011011111",
  22870=>"001110101",
  22871=>"010001011",
  22872=>"000001101",
  22873=>"110101111",
  22874=>"011111101",
  22875=>"100010111",
  22876=>"110010100",
  22877=>"100000010",
  22878=>"111000111",
  22879=>"000100001",
  22880=>"000010000",
  22881=>"110011101",
  22882=>"111001100",
  22883=>"001101011",
  22884=>"011111010",
  22885=>"100010100",
  22886=>"101101010",
  22887=>"101011010",
  22888=>"011000110",
  22889=>"100000110",
  22890=>"101101110",
  22891=>"011011001",
  22892=>"010000110",
  22893=>"000101100",
  22894=>"010001011",
  22895=>"101111100",
  22896=>"000101000",
  22897=>"110000011",
  22898=>"000101110",
  22899=>"111011010",
  22900=>"001011101",
  22901=>"111011110",
  22902=>"011110010",
  22903=>"010100000",
  22904=>"110110011",
  22905=>"011011110",
  22906=>"101111001",
  22907=>"101101000",
  22908=>"000111011",
  22909=>"110101010",
  22910=>"100011010",
  22911=>"100010001",
  22912=>"111001101",
  22913=>"001000110",
  22914=>"001000011",
  22915=>"110100011",
  22916=>"001000111",
  22917=>"000011010",
  22918=>"101000111",
  22919=>"110111010",
  22920=>"111000001",
  22921=>"011000010",
  22922=>"001101001",
  22923=>"100111011",
  22924=>"100110001",
  22925=>"001010000",
  22926=>"011110111",
  22927=>"101110011",
  22928=>"111000010",
  22929=>"001100111",
  22930=>"101100010",
  22931=>"101010011",
  22932=>"011000001",
  22933=>"110010010",
  22934=>"010000111",
  22935=>"011001111",
  22936=>"101111100",
  22937=>"101001010",
  22938=>"011101001",
  22939=>"011111111",
  22940=>"001111010",
  22941=>"011001001",
  22942=>"001001100",
  22943=>"001101101",
  22944=>"011100001",
  22945=>"011110100",
  22946=>"000101000",
  22947=>"110101011",
  22948=>"101111001",
  22949=>"110010100",
  22950=>"001011000",
  22951=>"111110100",
  22952=>"010001011",
  22953=>"000100100",
  22954=>"111100111",
  22955=>"101110000",
  22956=>"101000001",
  22957=>"101011100",
  22958=>"101010011",
  22959=>"010000001",
  22960=>"010111110",
  22961=>"101100111",
  22962=>"110110100",
  22963=>"011011001",
  22964=>"111011001",
  22965=>"000101001",
  22966=>"011100101",
  22967=>"010010111",
  22968=>"001000000",
  22969=>"010110110",
  22970=>"101111110",
  22971=>"110100001",
  22972=>"110111001",
  22973=>"010111001",
  22974=>"110010000",
  22975=>"100010011",
  22976=>"011110101",
  22977=>"111000010",
  22978=>"100110001",
  22979=>"111110101",
  22980=>"011101110",
  22981=>"011111001",
  22982=>"001010100",
  22983=>"111101010",
  22984=>"100110110",
  22985=>"111011001",
  22986=>"001000110",
  22987=>"110001110",
  22988=>"011000010",
  22989=>"111001111",
  22990=>"000101100",
  22991=>"011011000",
  22992=>"001101001",
  22993=>"100000101",
  22994=>"111111110",
  22995=>"010001011",
  22996=>"110000100",
  22997=>"000100111",
  22998=>"010100010",
  22999=>"011111101",
  23000=>"111011101",
  23001=>"001011100",
  23002=>"101011001",
  23003=>"101111110",
  23004=>"001011010",
  23005=>"101100000",
  23006=>"111011110",
  23007=>"001100001",
  23008=>"010111001",
  23009=>"110100001",
  23010=>"000011111",
  23011=>"100111100",
  23012=>"000100011",
  23013=>"000010111",
  23014=>"011001110",
  23015=>"111111000",
  23016=>"110010001",
  23017=>"011100000",
  23018=>"010100010",
  23019=>"000000001",
  23020=>"100111011",
  23021=>"001000000",
  23022=>"000001101",
  23023=>"110000011",
  23024=>"001001100",
  23025=>"100000000",
  23026=>"011000111",
  23027=>"101111011",
  23028=>"111111101",
  23029=>"001010100",
  23030=>"010100001",
  23031=>"010111001",
  23032=>"001000110",
  23033=>"011110100",
  23034=>"011111000",
  23035=>"111100001",
  23036=>"101011100",
  23037=>"101000001",
  23038=>"101100010",
  23039=>"011100010",
  23040=>"011111001",
  23041=>"000110111",
  23042=>"010100001",
  23043=>"111010111",
  23044=>"011010110",
  23045=>"100010111",
  23046=>"010100001",
  23047=>"100100000",
  23048=>"111100111",
  23049=>"111111010",
  23050=>"011011110",
  23051=>"100110111",
  23052=>"000100111",
  23053=>"010010101",
  23054=>"010100011",
  23055=>"000111111",
  23056=>"101110110",
  23057=>"010000011",
  23058=>"100010001",
  23059=>"110101110",
  23060=>"111000000",
  23061=>"010010010",
  23062=>"000110001",
  23063=>"101101101",
  23064=>"100011111",
  23065=>"000110110",
  23066=>"011011101",
  23067=>"011010010",
  23068=>"010110001",
  23069=>"110101000",
  23070=>"110101100",
  23071=>"010011011",
  23072=>"101011111",
  23073=>"101001011",
  23074=>"010110010",
  23075=>"101110001",
  23076=>"011011110",
  23077=>"111100100",
  23078=>"101100111",
  23079=>"101111111",
  23080=>"110100110",
  23081=>"010001001",
  23082=>"111001000",
  23083=>"001010010",
  23084=>"110111010",
  23085=>"110001010",
  23086=>"110011100",
  23087=>"011100100",
  23088=>"011011110",
  23089=>"011101000",
  23090=>"101000111",
  23091=>"100100110",
  23092=>"010000100",
  23093=>"111101000",
  23094=>"111100000",
  23095=>"011001100",
  23096=>"000010000",
  23097=>"011011000",
  23098=>"010110000",
  23099=>"011010011",
  23100=>"111000000",
  23101=>"011100111",
  23102=>"000001101",
  23103=>"110110000",
  23104=>"101111111",
  23105=>"101110110",
  23106=>"110101001",
  23107=>"100100100",
  23108=>"011010101",
  23109=>"000101110",
  23110=>"111100110",
  23111=>"100101100",
  23112=>"111010110",
  23113=>"001111000",
  23114=>"001011010",
  23115=>"001000100",
  23116=>"011001011",
  23117=>"010110000",
  23118=>"011001101",
  23119=>"000001001",
  23120=>"111110110",
  23121=>"110010010",
  23122=>"111000111",
  23123=>"010000110",
  23124=>"011010111",
  23125=>"111101101",
  23126=>"111010111",
  23127=>"111110111",
  23128=>"101011010",
  23129=>"100101011",
  23130=>"110000001",
  23131=>"101010101",
  23132=>"100101011",
  23133=>"101110101",
  23134=>"000011101",
  23135=>"000101001",
  23136=>"101101111",
  23137=>"110010100",
  23138=>"101101100",
  23139=>"000101111",
  23140=>"011100110",
  23141=>"101001111",
  23142=>"111111110",
  23143=>"110011000",
  23144=>"000100000",
  23145=>"110101010",
  23146=>"010000110",
  23147=>"011001101",
  23148=>"110001010",
  23149=>"110001010",
  23150=>"100111111",
  23151=>"001001001",
  23152=>"000010001",
  23153=>"010000110",
  23154=>"000010011",
  23155=>"101101011",
  23156=>"110101011",
  23157=>"101000111",
  23158=>"001011010",
  23159=>"100101100",
  23160=>"001010100",
  23161=>"101001001",
  23162=>"001111110",
  23163=>"100110110",
  23164=>"001001110",
  23165=>"001111001",
  23166=>"111111011",
  23167=>"000111010",
  23168=>"100101011",
  23169=>"010110011",
  23170=>"110000100",
  23171=>"101100100",
  23172=>"000010011",
  23173=>"000000000",
  23174=>"001010000",
  23175=>"001000100",
  23176=>"010111111",
  23177=>"000000010",
  23178=>"101100000",
  23179=>"100000010",
  23180=>"100001110",
  23181=>"000100001",
  23182=>"010000001",
  23183=>"110100110",
  23184=>"100110001",
  23185=>"110001110",
  23186=>"111100111",
  23187=>"100011011",
  23188=>"010100111",
  23189=>"101101001",
  23190=>"101000100",
  23191=>"110110111",
  23192=>"110000011",
  23193=>"001110101",
  23194=>"000001010",
  23195=>"110001110",
  23196=>"101000000",
  23197=>"110101110",
  23198=>"001011110",
  23199=>"010000010",
  23200=>"000110101",
  23201=>"110100111",
  23202=>"011101101",
  23203=>"001010001",
  23204=>"101001010",
  23205=>"111110000",
  23206=>"101100011",
  23207=>"010001011",
  23208=>"110010110",
  23209=>"101011101",
  23210=>"111101001",
  23211=>"100100001",
  23212=>"011010110",
  23213=>"111110010",
  23214=>"110111001",
  23215=>"110100111",
  23216=>"001001110",
  23217=>"100100001",
  23218=>"111100000",
  23219=>"001000010",
  23220=>"111000010",
  23221=>"101010111",
  23222=>"110101000",
  23223=>"111100110",
  23224=>"000000100",
  23225=>"110111110",
  23226=>"000010110",
  23227=>"010110001",
  23228=>"001001011",
  23229=>"001000101",
  23230=>"101010101",
  23231=>"010000000",
  23232=>"101001000",
  23233=>"000101110",
  23234=>"101101111",
  23235=>"111010111",
  23236=>"111111010",
  23237=>"101001110",
  23238=>"100001000",
  23239=>"100001101",
  23240=>"101101111",
  23241=>"111101010",
  23242=>"101000001",
  23243=>"011110001",
  23244=>"011101000",
  23245=>"000100000",
  23246=>"111110001",
  23247=>"110010110",
  23248=>"111101111",
  23249=>"100111000",
  23250=>"111101111",
  23251=>"101011111",
  23252=>"111101111",
  23253=>"100111000",
  23254=>"101010001",
  23255=>"011000101",
  23256=>"111011001",
  23257=>"010110010",
  23258=>"000000101",
  23259=>"101010110",
  23260=>"001101100",
  23261=>"000011010",
  23262=>"011100001",
  23263=>"110111110",
  23264=>"010011000",
  23265=>"001100101",
  23266=>"111010110",
  23267=>"000101001",
  23268=>"101101110",
  23269=>"010100111",
  23270=>"010100111",
  23271=>"110110100",
  23272=>"100100011",
  23273=>"100001101",
  23274=>"110000011",
  23275=>"110010101",
  23276=>"110000101",
  23277=>"101011000",
  23278=>"010010111",
  23279=>"010011110",
  23280=>"100100000",
  23281=>"011011100",
  23282=>"101000011",
  23283=>"101110010",
  23284=>"101010110",
  23285=>"111100011",
  23286=>"100001011",
  23287=>"010000000",
  23288=>"101111100",
  23289=>"100101111",
  23290=>"010001000",
  23291=>"111001100",
  23292=>"101000011",
  23293=>"110101101",
  23294=>"110100110",
  23295=>"101001101",
  23296=>"000101111",
  23297=>"100000000",
  23298=>"110101000",
  23299=>"011000010",
  23300=>"011010110",
  23301=>"011110000",
  23302=>"110010100",
  23303=>"100000011",
  23304=>"011100011",
  23305=>"110101111",
  23306=>"111011001",
  23307=>"000110000",
  23308=>"000000101",
  23309=>"101000000",
  23310=>"110000111",
  23311=>"010101111",
  23312=>"111001010",
  23313=>"110010101",
  23314=>"000000010",
  23315=>"000011101",
  23316=>"100111011",
  23317=>"001001110",
  23318=>"101001011",
  23319=>"111111011",
  23320=>"010110000",
  23321=>"001110001",
  23322=>"111010100",
  23323=>"111110011",
  23324=>"100010010",
  23325=>"001000001",
  23326=>"101110010",
  23327=>"001111101",
  23328=>"000100011",
  23329=>"101101010",
  23330=>"100110000",
  23331=>"110000011",
  23332=>"100100000",
  23333=>"111111111",
  23334=>"101000010",
  23335=>"100100011",
  23336=>"100000000",
  23337=>"000000101",
  23338=>"011101101",
  23339=>"011000010",
  23340=>"000111011",
  23341=>"011010111",
  23342=>"001000010",
  23343=>"010001000",
  23344=>"100100101",
  23345=>"000111000",
  23346=>"100011000",
  23347=>"100000101",
  23348=>"110110010",
  23349=>"100011100",
  23350=>"100101101",
  23351=>"011011010",
  23352=>"110010001",
  23353=>"100110101",
  23354=>"111101000",
  23355=>"010110101",
  23356=>"110111110",
  23357=>"010110100",
  23358=>"010000011",
  23359=>"110111101",
  23360=>"000001001",
  23361=>"110110000",
  23362=>"110001000",
  23363=>"000100111",
  23364=>"111110100",
  23365=>"111010010",
  23366=>"110001011",
  23367=>"111101011",
  23368=>"000100001",
  23369=>"011011111",
  23370=>"000011100",
  23371=>"000011111",
  23372=>"010010101",
  23373=>"011101110",
  23374=>"101110000",
  23375=>"110001001",
  23376=>"011011100",
  23377=>"001100110",
  23378=>"010110101",
  23379=>"001010010",
  23380=>"011000000",
  23381=>"110000111",
  23382=>"000100100",
  23383=>"011011011",
  23384=>"111111001",
  23385=>"011010010",
  23386=>"101100111",
  23387=>"000101110",
  23388=>"011000100",
  23389=>"001111100",
  23390=>"100001101",
  23391=>"111000101",
  23392=>"101100111",
  23393=>"010100001",
  23394=>"111111011",
  23395=>"100000010",
  23396=>"100011110",
  23397=>"010011001",
  23398=>"100101011",
  23399=>"000010001",
  23400=>"001110010",
  23401=>"100101101",
  23402=>"000000111",
  23403=>"100111110",
  23404=>"010000010",
  23405=>"111001001",
  23406=>"000001111",
  23407=>"010011010",
  23408=>"101010100",
  23409=>"110110000",
  23410=>"000101011",
  23411=>"101111001",
  23412=>"001010110",
  23413=>"010100010",
  23414=>"110110010",
  23415=>"100001001",
  23416=>"011001111",
  23417=>"111011101",
  23418=>"100000101",
  23419=>"101011011",
  23420=>"100111101",
  23421=>"010111011",
  23422=>"011000101",
  23423=>"011010000",
  23424=>"011101101",
  23425=>"000111110",
  23426=>"011000101",
  23427=>"000100000",
  23428=>"001011111",
  23429=>"011111011",
  23430=>"001010001",
  23431=>"110111101",
  23432=>"010001010",
  23433=>"011010000",
  23434=>"010000000",
  23435=>"011100000",
  23436=>"111111011",
  23437=>"111100011",
  23438=>"101100000",
  23439=>"100101110",
  23440=>"000000011",
  23441=>"110100101",
  23442=>"100000111",
  23443=>"000110101",
  23444=>"101110111",
  23445=>"100001101",
  23446=>"011111110",
  23447=>"000010101",
  23448=>"110000101",
  23449=>"110111011",
  23450=>"110100000",
  23451=>"010011110",
  23452=>"010101111",
  23453=>"101100110",
  23454=>"001011111",
  23455=>"010111110",
  23456=>"101101011",
  23457=>"101011101",
  23458=>"010001101",
  23459=>"110101111",
  23460=>"001000001",
  23461=>"010101011",
  23462=>"111001101",
  23463=>"111000011",
  23464=>"000010000",
  23465=>"000101010",
  23466=>"111101111",
  23467=>"010101011",
  23468=>"001100101",
  23469=>"100000000",
  23470=>"110101010",
  23471=>"101111000",
  23472=>"110100110",
  23473=>"010100111",
  23474=>"011011000",
  23475=>"001011001",
  23476=>"101100010",
  23477=>"100010000",
  23478=>"101111011",
  23479=>"010000110",
  23480=>"100011001",
  23481=>"000100001",
  23482=>"010011010",
  23483=>"001101101",
  23484=>"010101101",
  23485=>"111111111",
  23486=>"010001011",
  23487=>"010010010",
  23488=>"010101101",
  23489=>"010000110",
  23490=>"000011101",
  23491=>"100001101",
  23492=>"000001101",
  23493=>"110001010",
  23494=>"011110110",
  23495=>"111111111",
  23496=>"101011110",
  23497=>"000001010",
  23498=>"100001010",
  23499=>"010110010",
  23500=>"100010010",
  23501=>"111100101",
  23502=>"001110101",
  23503=>"001000101",
  23504=>"111100111",
  23505=>"011110011",
  23506=>"111100111",
  23507=>"100100101",
  23508=>"011000001",
  23509=>"111000000",
  23510=>"100001001",
  23511=>"101101001",
  23512=>"011000110",
  23513=>"001110000",
  23514=>"111111001",
  23515=>"100001010",
  23516=>"101111011",
  23517=>"100101110",
  23518=>"011111000",
  23519=>"001010000",
  23520=>"011001001",
  23521=>"110010010",
  23522=>"100000010",
  23523=>"101101110",
  23524=>"010110010",
  23525=>"010110101",
  23526=>"000010000",
  23527=>"001110011",
  23528=>"010100110",
  23529=>"110011001",
  23530=>"110110101",
  23531=>"101001010",
  23532=>"101001110",
  23533=>"010101000",
  23534=>"011010100",
  23535=>"011100010",
  23536=>"001011010",
  23537=>"110000101",
  23538=>"100001000",
  23539=>"011110111",
  23540=>"100110010",
  23541=>"011011010",
  23542=>"011010011",
  23543=>"011001101",
  23544=>"001000000",
  23545=>"110011101",
  23546=>"100110101",
  23547=>"111100111",
  23548=>"110010111",
  23549=>"001010000",
  23550=>"100000000",
  23551=>"111110011",
  23552=>"011111111",
  23553=>"000001000",
  23554=>"111101000",
  23555=>"101100011",
  23556=>"101100000",
  23557=>"111001011",
  23558=>"100110101",
  23559=>"100101000",
  23560=>"001100011",
  23561=>"010001001",
  23562=>"110111000",
  23563=>"111111000",
  23564=>"111000101",
  23565=>"010101110",
  23566=>"111110000",
  23567=>"011000101",
  23568=>"001000001",
  23569=>"000110000",
  23570=>"000110011",
  23571=>"110000001",
  23572=>"111011101",
  23573=>"001010101",
  23574=>"111100110",
  23575=>"111000011",
  23576=>"110101110",
  23577=>"111100001",
  23578=>"000100001",
  23579=>"011011011",
  23580=>"100001010",
  23581=>"111000100",
  23582=>"101010111",
  23583=>"001010100",
  23584=>"100001000",
  23585=>"111111111",
  23586=>"110100000",
  23587=>"011110010",
  23588=>"001111111",
  23589=>"001110100",
  23590=>"010110000",
  23591=>"011101000",
  23592=>"010010100",
  23593=>"001000010",
  23594=>"101111001",
  23595=>"100001010",
  23596=>"111111101",
  23597=>"101010101",
  23598=>"011100111",
  23599=>"000111011",
  23600=>"101100101",
  23601=>"100101100",
  23602=>"100001101",
  23603=>"110011000",
  23604=>"000000000",
  23605=>"111111010",
  23606=>"111010111",
  23607=>"101111100",
  23608=>"011100001",
  23609=>"001001010",
  23610=>"110001110",
  23611=>"110000010",
  23612=>"011010000",
  23613=>"100011011",
  23614=>"001000000",
  23615=>"000001101",
  23616=>"101010101",
  23617=>"001000011",
  23618=>"000100000",
  23619=>"010011001",
  23620=>"011000101",
  23621=>"000110010",
  23622=>"000110110",
  23623=>"010111111",
  23624=>"110101010",
  23625=>"000110011",
  23626=>"000110001",
  23627=>"001101111",
  23628=>"101111101",
  23629=>"000101010",
  23630=>"101011100",
  23631=>"000110101",
  23632=>"100001101",
  23633=>"001111000",
  23634=>"011010011",
  23635=>"100100111",
  23636=>"101110001",
  23637=>"100101111",
  23638=>"100111101",
  23639=>"000001100",
  23640=>"100111010",
  23641=>"100011111",
  23642=>"000011111",
  23643=>"011010110",
  23644=>"111011001",
  23645=>"010101101",
  23646=>"010000011",
  23647=>"011000000",
  23648=>"010111010",
  23649=>"100111001",
  23650=>"101000111",
  23651=>"001001001",
  23652=>"000101111",
  23653=>"001101010",
  23654=>"111110101",
  23655=>"001000100",
  23656=>"110100101",
  23657=>"000111000",
  23658=>"101010001",
  23659=>"011111101",
  23660=>"101000101",
  23661=>"100011001",
  23662=>"001011100",
  23663=>"001000011",
  23664=>"001001011",
  23665=>"110101101",
  23666=>"000110000",
  23667=>"100011011",
  23668=>"101101100",
  23669=>"110110111",
  23670=>"010001010",
  23671=>"011010101",
  23672=>"101100110",
  23673=>"011010000",
  23674=>"111010110",
  23675=>"010101110",
  23676=>"111000100",
  23677=>"100001100",
  23678=>"110001101",
  23679=>"111111010",
  23680=>"011010100",
  23681=>"010100110",
  23682=>"011000000",
  23683=>"110010010",
  23684=>"000110100",
  23685=>"100010100",
  23686=>"000010101",
  23687=>"001010001",
  23688=>"110110000",
  23689=>"010100011",
  23690=>"001000011",
  23691=>"010100101",
  23692=>"011001110",
  23693=>"101010011",
  23694=>"010000011",
  23695=>"010000110",
  23696=>"110100111",
  23697=>"110010111",
  23698=>"000101001",
  23699=>"010001101",
  23700=>"110001111",
  23701=>"010110001",
  23702=>"010101111",
  23703=>"001010011",
  23704=>"111001110",
  23705=>"101011101",
  23706=>"001011010",
  23707=>"100110100",
  23708=>"000000011",
  23709=>"100000100",
  23710=>"011100111",
  23711=>"010000011",
  23712=>"010000011",
  23713=>"110111111",
  23714=>"001110111",
  23715=>"111001011",
  23716=>"110001001",
  23717=>"111000001",
  23718=>"001000001",
  23719=>"010100001",
  23720=>"010001111",
  23721=>"001101011",
  23722=>"110111000",
  23723=>"001000111",
  23724=>"011011110",
  23725=>"001001111",
  23726=>"111111101",
  23727=>"011000010",
  23728=>"100000100",
  23729=>"000011111",
  23730=>"001011000",
  23731=>"000101101",
  23732=>"010000001",
  23733=>"101110111",
  23734=>"111101101",
  23735=>"111001000",
  23736=>"001011010",
  23737=>"010001100",
  23738=>"100110110",
  23739=>"100110001",
  23740=>"001100100",
  23741=>"101101101",
  23742=>"011011111",
  23743=>"101110101",
  23744=>"010001001",
  23745=>"001001111",
  23746=>"000100101",
  23747=>"111011100",
  23748=>"011001101",
  23749=>"101010110",
  23750=>"100000010",
  23751=>"001001100",
  23752=>"000101010",
  23753=>"101010100",
  23754=>"100010011",
  23755=>"100110101",
  23756=>"010001000",
  23757=>"111011000",
  23758=>"000001000",
  23759=>"011011101",
  23760=>"010100111",
  23761=>"100101001",
  23762=>"100001111",
  23763=>"001101011",
  23764=>"010001001",
  23765=>"100100110",
  23766=>"100010001",
  23767=>"111110110",
  23768=>"001000011",
  23769=>"010101110",
  23770=>"001100010",
  23771=>"111000000",
  23772=>"110010011",
  23773=>"111011111",
  23774=>"000010000",
  23775=>"011110000",
  23776=>"001010110",
  23777=>"011001101",
  23778=>"110101100",
  23779=>"110101100",
  23780=>"010000110",
  23781=>"000110111",
  23782=>"100111011",
  23783=>"110010110",
  23784=>"111011100",
  23785=>"000010010",
  23786=>"010111000",
  23787=>"010010011",
  23788=>"000110110",
  23789=>"111111110",
  23790=>"101100110",
  23791=>"111110101",
  23792=>"010110010",
  23793=>"010100000",
  23794=>"111111011",
  23795=>"011011100",
  23796=>"111001011",
  23797=>"101111000",
  23798=>"010001001",
  23799=>"100011011",
  23800=>"101111000",
  23801=>"011101010",
  23802=>"011111111",
  23803=>"110101000",
  23804=>"011111111",
  23805=>"110111110",
  23806=>"111000100",
  23807=>"000111011",
  23808=>"111001001",
  23809=>"010101110",
  23810=>"010011011",
  23811=>"101010110",
  23812=>"001100011",
  23813=>"110111001",
  23814=>"010100000",
  23815=>"100111111",
  23816=>"110110111",
  23817=>"000101111",
  23818=>"001100001",
  23819=>"111001110",
  23820=>"000000010",
  23821=>"010101101",
  23822=>"100110010",
  23823=>"000010100",
  23824=>"111000011",
  23825=>"100000011",
  23826=>"001100110",
  23827=>"101101001",
  23828=>"100101100",
  23829=>"111111100",
  23830=>"111011100",
  23831=>"000111011",
  23832=>"001100001",
  23833=>"110111111",
  23834=>"000010110",
  23835=>"011110000",
  23836=>"111000000",
  23837=>"110001000",
  23838=>"100101111",
  23839=>"010001110",
  23840=>"001010110",
  23841=>"111001000",
  23842=>"001101111",
  23843=>"110001110",
  23844=>"111001100",
  23845=>"111011000",
  23846=>"101111011",
  23847=>"101100010",
  23848=>"111000111",
  23849=>"010100111",
  23850=>"001010101",
  23851=>"100111010",
  23852=>"100111100",
  23853=>"110100101",
  23854=>"010101000",
  23855=>"011001000",
  23856=>"010010011",
  23857=>"011010001",
  23858=>"110010111",
  23859=>"101001100",
  23860=>"010101110",
  23861=>"001010001",
  23862=>"111111010",
  23863=>"001111001",
  23864=>"011100000",
  23865=>"011001110",
  23866=>"111010111",
  23867=>"010110000",
  23868=>"000101001",
  23869=>"101111100",
  23870=>"110111110",
  23871=>"101100000",
  23872=>"100101001",
  23873=>"110010001",
  23874=>"111011110",
  23875=>"110101001",
  23876=>"011101000",
  23877=>"011000100",
  23878=>"100000010",
  23879=>"110001001",
  23880=>"100011100",
  23881=>"100011101",
  23882=>"101100000",
  23883=>"011000000",
  23884=>"010011111",
  23885=>"111001001",
  23886=>"000101000",
  23887=>"111111001",
  23888=>"101010000",
  23889=>"100111010",
  23890=>"101001010",
  23891=>"001101111",
  23892=>"111011101",
  23893=>"010101011",
  23894=>"111010110",
  23895=>"101011110",
  23896=>"100001110",
  23897=>"001101101",
  23898=>"100100100",
  23899=>"000110001",
  23900=>"011001000",
  23901=>"011100010",
  23902=>"001111101",
  23903=>"000100010",
  23904=>"011010110",
  23905=>"111001101",
  23906=>"100101110",
  23907=>"101001111",
  23908=>"000000011",
  23909=>"011111001",
  23910=>"101011000",
  23911=>"101111000",
  23912=>"001101010",
  23913=>"011001011",
  23914=>"001000011",
  23915=>"111111110",
  23916=>"101111010",
  23917=>"100000000",
  23918=>"101011100",
  23919=>"000100010",
  23920=>"110010000",
  23921=>"010101101",
  23922=>"010000001",
  23923=>"100000000",
  23924=>"011000110",
  23925=>"111001100",
  23926=>"110111111",
  23927=>"010111001",
  23928=>"001110100",
  23929=>"010011000",
  23930=>"101011000",
  23931=>"101110011",
  23932=>"100011111",
  23933=>"101111111",
  23934=>"001100111",
  23935=>"101110011",
  23936=>"111111010",
  23937=>"010110010",
  23938=>"100001001",
  23939=>"001100111",
  23940=>"001000101",
  23941=>"000111010",
  23942=>"110111011",
  23943=>"000000111",
  23944=>"110111100",
  23945=>"111110110",
  23946=>"011011100",
  23947=>"111000101",
  23948=>"110010001",
  23949=>"000010010",
  23950=>"010000001",
  23951=>"011011100",
  23952=>"001101110",
  23953=>"110101000",
  23954=>"001110000",
  23955=>"100000111",
  23956=>"110110001",
  23957=>"110010100",
  23958=>"011010111",
  23959=>"100000110",
  23960=>"101101010",
  23961=>"000000001",
  23962=>"001100010",
  23963=>"000000100",
  23964=>"001110000",
  23965=>"111000010",
  23966=>"101110011",
  23967=>"100111000",
  23968=>"111001011",
  23969=>"001011000",
  23970=>"001001010",
  23971=>"100011001",
  23972=>"100100110",
  23973=>"011000010",
  23974=>"111011001",
  23975=>"100101011",
  23976=>"001001111",
  23977=>"111010100",
  23978=>"110100101",
  23979=>"010010101",
  23980=>"011011111",
  23981=>"110110101",
  23982=>"001101001",
  23983=>"101000010",
  23984=>"100001110",
  23985=>"111101010",
  23986=>"001111000",
  23987=>"001000001",
  23988=>"011110001",
  23989=>"011011011",
  23990=>"001000011",
  23991=>"111111110",
  23992=>"010101011",
  23993=>"110010011",
  23994=>"001101101",
  23995=>"010010100",
  23996=>"111110111",
  23997=>"011001100",
  23998=>"110000110",
  23999=>"011011001",
  24000=>"111001001",
  24001=>"001011101",
  24002=>"011010001",
  24003=>"100001010",
  24004=>"111111100",
  24005=>"010010100",
  24006=>"001000000",
  24007=>"011000100",
  24008=>"010010101",
  24009=>"100110011",
  24010=>"110110011",
  24011=>"010111101",
  24012=>"111110111",
  24013=>"111000011",
  24014=>"111000010",
  24015=>"111110110",
  24016=>"111101001",
  24017=>"111001101",
  24018=>"001001111",
  24019=>"000100000",
  24020=>"011000101",
  24021=>"101001100",
  24022=>"110001110",
  24023=>"100001101",
  24024=>"010101101",
  24025=>"101110100",
  24026=>"011001011",
  24027=>"010000110",
  24028=>"101110000",
  24029=>"000000111",
  24030=>"101110110",
  24031=>"100001110",
  24032=>"100111010",
  24033=>"011110011",
  24034=>"111101001",
  24035=>"001111010",
  24036=>"110110110",
  24037=>"000111110",
  24038=>"111101110",
  24039=>"110111001",
  24040=>"000100000",
  24041=>"001000100",
  24042=>"010100101",
  24043=>"000011000",
  24044=>"000001010",
  24045=>"010100010",
  24046=>"011001001",
  24047=>"011110111",
  24048=>"111100101",
  24049=>"101010010",
  24050=>"000110101",
  24051=>"101111010",
  24052=>"100111010",
  24053=>"000010110",
  24054=>"101101010",
  24055=>"000000010",
  24056=>"000111110",
  24057=>"010010100",
  24058=>"111101100",
  24059=>"010000011",
  24060=>"100000011",
  24061=>"111000000",
  24062=>"100001000",
  24063=>"111011100",
  24064=>"010110111",
  24065=>"110010011",
  24066=>"000000011",
  24067=>"011010111",
  24068=>"001101110",
  24069=>"110101011",
  24070=>"011010100",
  24071=>"011011110",
  24072=>"001100110",
  24073=>"100100011",
  24074=>"111111011",
  24075=>"000011111",
  24076=>"011101010",
  24077=>"001110101",
  24078=>"111000110",
  24079=>"011011011",
  24080=>"100000000",
  24081=>"100111010",
  24082=>"010111111",
  24083=>"011111000",
  24084=>"100000001",
  24085=>"011101000",
  24086=>"010100100",
  24087=>"000001100",
  24088=>"011001111",
  24089=>"010110110",
  24090=>"100111000",
  24091=>"011010010",
  24092=>"100100110",
  24093=>"101000101",
  24094=>"010001000",
  24095=>"110111000",
  24096=>"011010000",
  24097=>"011000010",
  24098=>"010110111",
  24099=>"111011101",
  24100=>"101010110",
  24101=>"100001110",
  24102=>"011110110",
  24103=>"000000100",
  24104=>"011110110",
  24105=>"110010111",
  24106=>"011000111",
  24107=>"011011000",
  24108=>"001110110",
  24109=>"011111000",
  24110=>"110001110",
  24111=>"111001110",
  24112=>"110010010",
  24113=>"111100111",
  24114=>"110001100",
  24115=>"001101001",
  24116=>"101100001",
  24117=>"010100100",
  24118=>"101110100",
  24119=>"110101011",
  24120=>"111000001",
  24121=>"100101010",
  24122=>"111100111",
  24123=>"001011111",
  24124=>"000000111",
  24125=>"100111100",
  24126=>"001001100",
  24127=>"001011010",
  24128=>"001111111",
  24129=>"101111110",
  24130=>"001010111",
  24131=>"010001101",
  24132=>"001110101",
  24133=>"111000101",
  24134=>"001110101",
  24135=>"011001100",
  24136=>"011011110",
  24137=>"011100001",
  24138=>"111110001",
  24139=>"101001001",
  24140=>"100000110",
  24141=>"100100010",
  24142=>"110011011",
  24143=>"111111110",
  24144=>"111100010",
  24145=>"100011100",
  24146=>"000101111",
  24147=>"100100101",
  24148=>"001111111",
  24149=>"001100101",
  24150=>"100000000",
  24151=>"001001010",
  24152=>"010100111",
  24153=>"110001001",
  24154=>"100000011",
  24155=>"110010000",
  24156=>"101001001",
  24157=>"000001010",
  24158=>"111010100",
  24159=>"001001000",
  24160=>"001101010",
  24161=>"011000110",
  24162=>"000011011",
  24163=>"000000001",
  24164=>"000000111",
  24165=>"111111001",
  24166=>"101101111",
  24167=>"011000101",
  24168=>"101110011",
  24169=>"011110010",
  24170=>"110111101",
  24171=>"110001000",
  24172=>"100000001",
  24173=>"101100111",
  24174=>"110111100",
  24175=>"100010001",
  24176=>"001011110",
  24177=>"001001011",
  24178=>"111100101",
  24179=>"010101011",
  24180=>"010010110",
  24181=>"110111000",
  24182=>"100100101",
  24183=>"101011001",
  24184=>"100010111",
  24185=>"000011100",
  24186=>"011010100",
  24187=>"000100010",
  24188=>"001011101",
  24189=>"010101000",
  24190=>"001000000",
  24191=>"100110010",
  24192=>"000110100",
  24193=>"011011000",
  24194=>"111101110",
  24195=>"000001001",
  24196=>"100011111",
  24197=>"101101001",
  24198=>"011100011",
  24199=>"000111110",
  24200=>"110001001",
  24201=>"011111110",
  24202=>"111111110",
  24203=>"010110100",
  24204=>"101110110",
  24205=>"001011111",
  24206=>"100001000",
  24207=>"000110001",
  24208=>"110100110",
  24209=>"001010011",
  24210=>"000110001",
  24211=>"010110010",
  24212=>"001101011",
  24213=>"101000001",
  24214=>"100110101",
  24215=>"100011100",
  24216=>"110000011",
  24217=>"000010000",
  24218=>"101000101",
  24219=>"110000111",
  24220=>"000110110",
  24221=>"000010100",
  24222=>"001110001",
  24223=>"011110011",
  24224=>"001011101",
  24225=>"100001100",
  24226=>"000110111",
  24227=>"010001001",
  24228=>"011110000",
  24229=>"010111011",
  24230=>"010101001",
  24231=>"010110100",
  24232=>"010000100",
  24233=>"101010000",
  24234=>"111101110",
  24235=>"010010100",
  24236=>"111101111",
  24237=>"011111001",
  24238=>"001101111",
  24239=>"001111000",
  24240=>"001000001",
  24241=>"000001011",
  24242=>"111011000",
  24243=>"011011001",
  24244=>"011001010",
  24245=>"111101010",
  24246=>"111000111",
  24247=>"110110001",
  24248=>"010001101",
  24249=>"011101111",
  24250=>"100001110",
  24251=>"001100101",
  24252=>"011000101",
  24253=>"110001110",
  24254=>"001111000",
  24255=>"000100011",
  24256=>"001010001",
  24257=>"011011010",
  24258=>"011000100",
  24259=>"111000100",
  24260=>"010000111",
  24261=>"000100111",
  24262=>"011000000",
  24263=>"101101001",
  24264=>"001111011",
  24265=>"111010000",
  24266=>"000000011",
  24267=>"110110011",
  24268=>"001000101",
  24269=>"110000010",
  24270=>"110010110",
  24271=>"001000100",
  24272=>"101100101",
  24273=>"011110100",
  24274=>"111110110",
  24275=>"000001001",
  24276=>"100111001",
  24277=>"101000100",
  24278=>"110000110",
  24279=>"001010011",
  24280=>"011010100",
  24281=>"110110010",
  24282=>"010100111",
  24283=>"110010000",
  24284=>"101110111",
  24285=>"111000010",
  24286=>"010001101",
  24287=>"100011111",
  24288=>"000000100",
  24289=>"001111111",
  24290=>"111111010",
  24291=>"101000000",
  24292=>"000101100",
  24293=>"000101110",
  24294=>"011111110",
  24295=>"100111000",
  24296=>"100010111",
  24297=>"011000010",
  24298=>"000000101",
  24299=>"100101001",
  24300=>"110001110",
  24301=>"011110111",
  24302=>"111101011",
  24303=>"010101011",
  24304=>"011000111",
  24305=>"011110010",
  24306=>"010010010",
  24307=>"010010100",
  24308=>"110101001",
  24309=>"110010111",
  24310=>"111010010",
  24311=>"010100111",
  24312=>"101010101",
  24313=>"111101111",
  24314=>"110001111",
  24315=>"101101011",
  24316=>"101101010",
  24317=>"101000100",
  24318=>"111110011",
  24319=>"000011010",
  24320=>"110110101",
  24321=>"110010000",
  24322=>"101010110",
  24323=>"111010011",
  24324=>"101001110",
  24325=>"111100101",
  24326=>"001111001",
  24327=>"000001011",
  24328=>"010100001",
  24329=>"001011001",
  24330=>"100011101",
  24331=>"011110001",
  24332=>"111000011",
  24333=>"010111101",
  24334=>"111011010",
  24335=>"111001101",
  24336=>"110001011",
  24337=>"101010000",
  24338=>"111000110",
  24339=>"101010010",
  24340=>"011110011",
  24341=>"000111011",
  24342=>"010101000",
  24343=>"010110001",
  24344=>"111101111",
  24345=>"100110111",
  24346=>"000001001",
  24347=>"010110100",
  24348=>"000010100",
  24349=>"111001001",
  24350=>"010011111",
  24351=>"111000100",
  24352=>"110110000",
  24353=>"111111111",
  24354=>"111000000",
  24355=>"010110011",
  24356=>"001000110",
  24357=>"100010001",
  24358=>"000111101",
  24359=>"000111101",
  24360=>"100110110",
  24361=>"111001110",
  24362=>"010101000",
  24363=>"111001011",
  24364=>"111001101",
  24365=>"011001101",
  24366=>"000000100",
  24367=>"110111001",
  24368=>"110100111",
  24369=>"001010010",
  24370=>"011111100",
  24371=>"100100011",
  24372=>"000111101",
  24373=>"001011010",
  24374=>"100001110",
  24375=>"001111010",
  24376=>"000101111",
  24377=>"010011100",
  24378=>"000100001",
  24379=>"100110011",
  24380=>"100000110",
  24381=>"100110101",
  24382=>"111000100",
  24383=>"111000111",
  24384=>"111100011",
  24385=>"110011000",
  24386=>"111111100",
  24387=>"011100011",
  24388=>"011000010",
  24389=>"010001001",
  24390=>"001000011",
  24391=>"101110001",
  24392=>"010001110",
  24393=>"111011101",
  24394=>"001011101",
  24395=>"101010100",
  24396=>"111101010",
  24397=>"100111010",
  24398=>"001101011",
  24399=>"101111010",
  24400=>"001110000",
  24401=>"100001101",
  24402=>"111000100",
  24403=>"111101011",
  24404=>"001011000",
  24405=>"010000111",
  24406=>"011001010",
  24407=>"100100011",
  24408=>"011000101",
  24409=>"000101101",
  24410=>"111111001",
  24411=>"010010100",
  24412=>"111011001",
  24413=>"000101000",
  24414=>"101100110",
  24415=>"010111001",
  24416=>"110111010",
  24417=>"000110000",
  24418=>"100100001",
  24419=>"101100010",
  24420=>"100010000",
  24421=>"010111010",
  24422=>"010111111",
  24423=>"011010011",
  24424=>"000110010",
  24425=>"101000100",
  24426=>"011110101",
  24427=>"101000110",
  24428=>"011010100",
  24429=>"011100000",
  24430=>"110111011",
  24431=>"000110110",
  24432=>"110110001",
  24433=>"111101101",
  24434=>"001101000",
  24435=>"010101000",
  24436=>"001011110",
  24437=>"000000100",
  24438=>"100110100",
  24439=>"110001001",
  24440=>"110101001",
  24441=>"101111001",
  24442=>"001110000",
  24443=>"001111011",
  24444=>"110110011",
  24445=>"010100110",
  24446=>"001101011",
  24447=>"100110101",
  24448=>"010101011",
  24449=>"111001110",
  24450=>"100010010",
  24451=>"111010010",
  24452=>"100010000",
  24453=>"101011011",
  24454=>"011110001",
  24455=>"001101101",
  24456=>"101100100",
  24457=>"000010100",
  24458=>"101100000",
  24459=>"000101010",
  24460=>"111100001",
  24461=>"100100111",
  24462=>"100110000",
  24463=>"000101010",
  24464=>"110111101",
  24465=>"011001001",
  24466=>"011100111",
  24467=>"100100010",
  24468=>"111010101",
  24469=>"100011011",
  24470=>"011000100",
  24471=>"111010010",
  24472=>"111011111",
  24473=>"100110001",
  24474=>"000011001",
  24475=>"101010101",
  24476=>"001000011",
  24477=>"110110000",
  24478=>"100000111",
  24479=>"001111111",
  24480=>"101110010",
  24481=>"110111000",
  24482=>"011011111",
  24483=>"000000000",
  24484=>"010001000",
  24485=>"001011111",
  24486=>"110011110",
  24487=>"101001100",
  24488=>"101000111",
  24489=>"010101001",
  24490=>"101001011",
  24491=>"111000101",
  24492=>"000111001",
  24493=>"011100011",
  24494=>"001000101",
  24495=>"001100011",
  24496=>"000101101",
  24497=>"010101100",
  24498=>"001101100",
  24499=>"110110101",
  24500=>"101001001",
  24501=>"000100001",
  24502=>"000001110",
  24503=>"111001110",
  24504=>"101001000",
  24505=>"100010000",
  24506=>"110011100",
  24507=>"111000111",
  24508=>"111000110",
  24509=>"111011010",
  24510=>"011010011",
  24511=>"011100010",
  24512=>"101001111",
  24513=>"000100101",
  24514=>"000011110",
  24515=>"000001100",
  24516=>"101110000",
  24517=>"011100100",
  24518=>"010111010",
  24519=>"111001000",
  24520=>"000010010",
  24521=>"110100010",
  24522=>"111111010",
  24523=>"010011101",
  24524=>"001111010",
  24525=>"111101000",
  24526=>"010011001",
  24527=>"010100000",
  24528=>"001010001",
  24529=>"111010000",
  24530=>"011101111",
  24531=>"000111011",
  24532=>"000110110",
  24533=>"000100000",
  24534=>"101011010",
  24535=>"100010101",
  24536=>"111110010",
  24537=>"001001101",
  24538=>"110111111",
  24539=>"001001101",
  24540=>"100001011",
  24541=>"110100101",
  24542=>"100000001",
  24543=>"101101110",
  24544=>"010111001",
  24545=>"000110011",
  24546=>"111110100",
  24547=>"011100110",
  24548=>"000000001",
  24549=>"111001011",
  24550=>"001111101",
  24551=>"001111110",
  24552=>"000001101",
  24553=>"011100101",
  24554=>"110001110",
  24555=>"100110111",
  24556=>"001011011",
  24557=>"011001110",
  24558=>"011101110",
  24559=>"010101111",
  24560=>"010000000",
  24561=>"101000110",
  24562=>"101101001",
  24563=>"100010010",
  24564=>"111111110",
  24565=>"011100001",
  24566=>"101011000",
  24567=>"010100010",
  24568=>"011011000",
  24569=>"011001011",
  24570=>"101000000",
  24571=>"111110000",
  24572=>"010011100",
  24573=>"100000101",
  24574=>"111110100",
  24575=>"011010000",
  24576=>"001010010",
  24577=>"001101101",
  24578=>"010001111",
  24579=>"000100010",
  24580=>"011100101",
  24581=>"000001000",
  24582=>"101111111",
  24583=>"101110101",
  24584=>"001100010",
  24585=>"101100011",
  24586=>"100010010",
  24587=>"111011011",
  24588=>"110000011",
  24589=>"010010110",
  24590=>"010001001",
  24591=>"001110100",
  24592=>"101111101",
  24593=>"011000000",
  24594=>"111110010",
  24595=>"010011010",
  24596=>"011110001",
  24597=>"110011001",
  24598=>"000011011",
  24599=>"010110001",
  24600=>"010101110",
  24601=>"110111100",
  24602=>"111001111",
  24603=>"110101100",
  24604=>"011111110",
  24605=>"101001111",
  24606=>"111100110",
  24607=>"110110001",
  24608=>"101001001",
  24609=>"100111001",
  24610=>"001000111",
  24611=>"001001110",
  24612=>"100000110",
  24613=>"011111000",
  24614=>"100100001",
  24615=>"001011110",
  24616=>"011001111",
  24617=>"001100111",
  24618=>"011010001",
  24619=>"001001111",
  24620=>"000010010",
  24621=>"110011000",
  24622=>"001101000",
  24623=>"000011001",
  24624=>"000011001",
  24625=>"101001010",
  24626=>"010001010",
  24627=>"010001001",
  24628=>"011001011",
  24629=>"011011010",
  24630=>"100011110",
  24631=>"000011110",
  24632=>"101001110",
  24633=>"010011000",
  24634=>"010000101",
  24635=>"101011011",
  24636=>"110000000",
  24637=>"010101100",
  24638=>"111101000",
  24639=>"101100000",
  24640=>"000000001",
  24641=>"000001010",
  24642=>"001001010",
  24643=>"000101011",
  24644=>"101001111",
  24645=>"001001111",
  24646=>"101101010",
  24647=>"001111000",
  24648=>"110100000",
  24649=>"010110111",
  24650=>"111111101",
  24651=>"011010111",
  24652=>"111100111",
  24653=>"110011100",
  24654=>"111000010",
  24655=>"111101111",
  24656=>"011010001",
  24657=>"100011100",
  24658=>"001010011",
  24659=>"100110001",
  24660=>"110100111",
  24661=>"100010110",
  24662=>"011111010",
  24663=>"001000011",
  24664=>"111110111",
  24665=>"010000000",
  24666=>"101110110",
  24667=>"100110001",
  24668=>"001011011",
  24669=>"111101111",
  24670=>"111011011",
  24671=>"011000101",
  24672=>"010000101",
  24673=>"100000101",
  24674=>"001101011",
  24675=>"011000001",
  24676=>"111110010",
  24677=>"000000111",
  24678=>"000010110",
  24679=>"000000001",
  24680=>"000000001",
  24681=>"101111110",
  24682=>"101000111",
  24683=>"101101010",
  24684=>"011010111",
  24685=>"011110011",
  24686=>"111101000",
  24687=>"110101100",
  24688=>"101100010",
  24689=>"110101011",
  24690=>"110010011",
  24691=>"010000000",
  24692=>"110010100",
  24693=>"100000010",
  24694=>"101001001",
  24695=>"101001110",
  24696=>"100010111",
  24697=>"100110101",
  24698=>"011000001",
  24699=>"110111110",
  24700=>"010000000",
  24701=>"100000001",
  24702=>"011101110",
  24703=>"011101000",
  24704=>"110001011",
  24705=>"110011110",
  24706=>"110111000",
  24707=>"100010010",
  24708=>"000000000",
  24709=>"001110100",
  24710=>"011111011",
  24711=>"101000110",
  24712=>"010000010",
  24713=>"101110110",
  24714=>"111000101",
  24715=>"111001010",
  24716=>"110101101",
  24717=>"110101100",
  24718=>"101001000",
  24719=>"011011110",
  24720=>"100000001",
  24721=>"000111110",
  24722=>"011000010",
  24723=>"110000100",
  24724=>"011111011",
  24725=>"110100010",
  24726=>"110010011",
  24727=>"000000001",
  24728=>"000100101",
  24729=>"010111110",
  24730=>"010101110",
  24731=>"111010000",
  24732=>"101000011",
  24733=>"110011000",
  24734=>"101110011",
  24735=>"110001111",
  24736=>"011110110",
  24737=>"101101110",
  24738=>"000000001",
  24739=>"100100011",
  24740=>"011001101",
  24741=>"011100000",
  24742=>"100101011",
  24743=>"011101010",
  24744=>"010100000",
  24745=>"100001011",
  24746=>"011010011",
  24747=>"110111110",
  24748=>"000011111",
  24749=>"010010101",
  24750=>"001110000",
  24751=>"001010011",
  24752=>"101111111",
  24753=>"110111111",
  24754=>"011010001",
  24755=>"001001011",
  24756=>"100000010",
  24757=>"010100100",
  24758=>"000001100",
  24759=>"101110011",
  24760=>"101010101",
  24761=>"110111000",
  24762=>"101111001",
  24763=>"111000111",
  24764=>"010110000",
  24765=>"111101010",
  24766=>"001000011",
  24767=>"110110011",
  24768=>"100001101",
  24769=>"111010100",
  24770=>"001110100",
  24771=>"011011110",
  24772=>"011000000",
  24773=>"000001101",
  24774=>"001000111",
  24775=>"011100111",
  24776=>"011110100",
  24777=>"101101001",
  24778=>"101101101",
  24779=>"111101011",
  24780=>"111010110",
  24781=>"001001111",
  24782=>"001001011",
  24783=>"101000000",
  24784=>"011110000",
  24785=>"010000011",
  24786=>"110110000",
  24787=>"100110100",
  24788=>"110111000",
  24789=>"111001100",
  24790=>"101010001",
  24791=>"010100101",
  24792=>"010101100",
  24793=>"000011010",
  24794=>"001010001",
  24795=>"010001001",
  24796=>"010000010",
  24797=>"010000100",
  24798=>"010110001",
  24799=>"111111011",
  24800=>"000110110",
  24801=>"111010110",
  24802=>"110111010",
  24803=>"110101110",
  24804=>"000101001",
  24805=>"111110111",
  24806=>"110110100",
  24807=>"000101111",
  24808=>"100010111",
  24809=>"100111000",
  24810=>"111001010",
  24811=>"110000111",
  24812=>"110111100",
  24813=>"110000101",
  24814=>"101110001",
  24815=>"001000111",
  24816=>"110011111",
  24817=>"011110010",
  24818=>"011000100",
  24819=>"000000001",
  24820=>"011001011",
  24821=>"011101001",
  24822=>"100110110",
  24823=>"000100011",
  24824=>"010000110",
  24825=>"111010001",
  24826=>"000101001",
  24827=>"110000100",
  24828=>"100000110",
  24829=>"110100011",
  24830=>"000101001",
  24831=>"110111011",
  24832=>"101000101",
  24833=>"101111101",
  24834=>"001001010",
  24835=>"001010001",
  24836=>"010011100",
  24837=>"000001110",
  24838=>"101011101",
  24839=>"011101000",
  24840=>"111001100",
  24841=>"100000000",
  24842=>"101000010",
  24843=>"110110010",
  24844=>"001000100",
  24845=>"100000010",
  24846=>"000100001",
  24847=>"111110100",
  24848=>"111110001",
  24849=>"101101100",
  24850=>"100010010",
  24851=>"111100100",
  24852=>"010110101",
  24853=>"111110100",
  24854=>"011000101",
  24855=>"011010011",
  24856=>"001001010",
  24857=>"000001010",
  24858=>"111110010",
  24859=>"001011010",
  24860=>"000101000",
  24861=>"110011111",
  24862=>"100010000",
  24863=>"001110000",
  24864=>"010010111",
  24865=>"011111011",
  24866=>"111101101",
  24867=>"111010101",
  24868=>"111101010",
  24869=>"011111011",
  24870=>"000110010",
  24871=>"000001111",
  24872=>"000000011",
  24873=>"000100111",
  24874=>"010001001",
  24875=>"011101110",
  24876=>"000100100",
  24877=>"001011010",
  24878=>"000100000",
  24879=>"100101011",
  24880=>"110010111",
  24881=>"100001000",
  24882=>"111011101",
  24883=>"011010010",
  24884=>"011100011",
  24885=>"110110111",
  24886=>"000111110",
  24887=>"110111111",
  24888=>"010100001",
  24889=>"011111111",
  24890=>"100111101",
  24891=>"001000001",
  24892=>"100001110",
  24893=>"111001011",
  24894=>"110100110",
  24895=>"001001000",
  24896=>"100011011",
  24897=>"001111110",
  24898=>"111000010",
  24899=>"111111101",
  24900=>"101101100",
  24901=>"010110100",
  24902=>"100000011",
  24903=>"010010101",
  24904=>"111101010",
  24905=>"000101100",
  24906=>"001111110",
  24907=>"000010011",
  24908=>"101000101",
  24909=>"000100100",
  24910=>"001010110",
  24911=>"011111111",
  24912=>"101110111",
  24913=>"001000001",
  24914=>"101101100",
  24915=>"110011011",
  24916=>"010110101",
  24917=>"100100001",
  24918=>"111010111",
  24919=>"011101010",
  24920=>"001000011",
  24921=>"001010100",
  24922=>"010000000",
  24923=>"100011110",
  24924=>"010100000",
  24925=>"010010001",
  24926=>"101110111",
  24927=>"100110010",
  24928=>"011010100",
  24929=>"000110100",
  24930=>"000001100",
  24931=>"100000110",
  24932=>"000011111",
  24933=>"000110001",
  24934=>"111001110",
  24935=>"110111001",
  24936=>"000100000",
  24937=>"101000010",
  24938=>"011100100",
  24939=>"001001111",
  24940=>"000101111",
  24941=>"000111010",
  24942=>"100110101",
  24943=>"110101100",
  24944=>"001010111",
  24945=>"010001100",
  24946=>"101101011",
  24947=>"011011001",
  24948=>"001110001",
  24949=>"001000000",
  24950=>"011000010",
  24951=>"101000001",
  24952=>"111111010",
  24953=>"000100111",
  24954=>"001101001",
  24955=>"010000011",
  24956=>"101111000",
  24957=>"000101011",
  24958=>"100111111",
  24959=>"010001001",
  24960=>"001100001",
  24961=>"100000001",
  24962=>"001100011",
  24963=>"101001000",
  24964=>"010101110",
  24965=>"001000101",
  24966=>"001011100",
  24967=>"100010101",
  24968=>"010000111",
  24969=>"111110110",
  24970=>"010011010",
  24971=>"100100111",
  24972=>"010111111",
  24973=>"001001000",
  24974=>"011010000",
  24975=>"110000000",
  24976=>"110010001",
  24977=>"101010000",
  24978=>"010000110",
  24979=>"010101111",
  24980=>"010101101",
  24981=>"000010010",
  24982=>"011001010",
  24983=>"111110101",
  24984=>"000101001",
  24985=>"111001111",
  24986=>"100111100",
  24987=>"100001111",
  24988=>"100010110",
  24989=>"010110110",
  24990=>"100101110",
  24991=>"111000111",
  24992=>"111111111",
  24993=>"110100010",
  24994=>"010010000",
  24995=>"000001001",
  24996=>"100011011",
  24997=>"001000000",
  24998=>"011111111",
  24999=>"100010000",
  25000=>"000110111",
  25001=>"101011100",
  25002=>"000010110",
  25003=>"100000000",
  25004=>"111100111",
  25005=>"001110011",
  25006=>"001110111",
  25007=>"001011000",
  25008=>"110111110",
  25009=>"110100110",
  25010=>"000110101",
  25011=>"000111111",
  25012=>"010110110",
  25013=>"011011010",
  25014=>"100111100",
  25015=>"100101010",
  25016=>"110111011",
  25017=>"101011000",
  25018=>"111001010",
  25019=>"100001001",
  25020=>"111011111",
  25021=>"110011011",
  25022=>"001111100",
  25023=>"100001110",
  25024=>"111101000",
  25025=>"111011000",
  25026=>"111011011",
  25027=>"110011000",
  25028=>"111101011",
  25029=>"111001001",
  25030=>"110000111",
  25031=>"000001110",
  25032=>"100000001",
  25033=>"010111100",
  25034=>"011111011",
  25035=>"111010010",
  25036=>"101000011",
  25037=>"111111110",
  25038=>"000010011",
  25039=>"011001011",
  25040=>"011001100",
  25041=>"110011100",
  25042=>"100101010",
  25043=>"111100101",
  25044=>"011110110",
  25045=>"111011000",
  25046=>"100101001",
  25047=>"110000111",
  25048=>"111100101",
  25049=>"111100001",
  25050=>"110100010",
  25051=>"010100011",
  25052=>"110000001",
  25053=>"100111110",
  25054=>"110101101",
  25055=>"011000110",
  25056=>"110110100",
  25057=>"110010000",
  25058=>"100111000",
  25059=>"111111000",
  25060=>"000110000",
  25061=>"000000101",
  25062=>"100111100",
  25063=>"111101111",
  25064=>"010001010",
  25065=>"011011011",
  25066=>"000001001",
  25067=>"101010101",
  25068=>"100101001",
  25069=>"111110100",
  25070=>"001010101",
  25071=>"011101011",
  25072=>"010111101",
  25073=>"110100101",
  25074=>"101011010",
  25075=>"110100011",
  25076=>"111011011",
  25077=>"000000011",
  25078=>"011011011",
  25079=>"001001010",
  25080=>"001010011",
  25081=>"100100001",
  25082=>"011110111",
  25083=>"001111110",
  25084=>"100010111",
  25085=>"111110010",
  25086=>"110010111",
  25087=>"011110000",
  25088=>"111011101",
  25089=>"000011001",
  25090=>"110000000",
  25091=>"000000101",
  25092=>"101000010",
  25093=>"100010101",
  25094=>"110111011",
  25095=>"011100001",
  25096=>"110101000",
  25097=>"011111110",
  25098=>"110010010",
  25099=>"000110000",
  25100=>"101011110",
  25101=>"111001001",
  25102=>"000110010",
  25103=>"111110111",
  25104=>"011000010",
  25105=>"001010000",
  25106=>"100010111",
  25107=>"001000101",
  25108=>"011011011",
  25109=>"100101010",
  25110=>"010111110",
  25111=>"010111001",
  25112=>"100110011",
  25113=>"110011010",
  25114=>"100001000",
  25115=>"110010010",
  25116=>"100101001",
  25117=>"111010010",
  25118=>"001011101",
  25119=>"010001101",
  25120=>"100100111",
  25121=>"111010000",
  25122=>"010011000",
  25123=>"011001000",
  25124=>"011000010",
  25125=>"010000010",
  25126=>"000100011",
  25127=>"010001100",
  25128=>"001000001",
  25129=>"110111111",
  25130=>"010010000",
  25131=>"111111000",
  25132=>"111111101",
  25133=>"000011110",
  25134=>"101110110",
  25135=>"101111001",
  25136=>"100111111",
  25137=>"000101000",
  25138=>"100110000",
  25139=>"011010101",
  25140=>"101101011",
  25141=>"101010010",
  25142=>"001101011",
  25143=>"010110010",
  25144=>"111111010",
  25145=>"111001100",
  25146=>"100011011",
  25147=>"000000111",
  25148=>"000010001",
  25149=>"110000001",
  25150=>"100011001",
  25151=>"101001111",
  25152=>"111111100",
  25153=>"111100111",
  25154=>"000010101",
  25155=>"110000011",
  25156=>"011010000",
  25157=>"011001000",
  25158=>"100000111",
  25159=>"100101000",
  25160=>"011101011",
  25161=>"001100001",
  25162=>"001101001",
  25163=>"110011000",
  25164=>"011010010",
  25165=>"111100010",
  25166=>"111010000",
  25167=>"001010000",
  25168=>"000010001",
  25169=>"011011100",
  25170=>"100100010",
  25171=>"110110001",
  25172=>"100100010",
  25173=>"000110011",
  25174=>"101110100",
  25175=>"000000110",
  25176=>"001000000",
  25177=>"001001010",
  25178=>"111011011",
  25179=>"000100100",
  25180=>"010010001",
  25181=>"111011111",
  25182=>"111101001",
  25183=>"000001101",
  25184=>"001001010",
  25185=>"110101000",
  25186=>"010001001",
  25187=>"100110101",
  25188=>"000100110",
  25189=>"101101001",
  25190=>"100000010",
  25191=>"110010110",
  25192=>"101010001",
  25193=>"001000000",
  25194=>"110110010",
  25195=>"101000101",
  25196=>"000111100",
  25197=>"001101000",
  25198=>"001100011",
  25199=>"001010111",
  25200=>"010100011",
  25201=>"011000011",
  25202=>"000111011",
  25203=>"111010010",
  25204=>"100101100",
  25205=>"000110010",
  25206=>"011110010",
  25207=>"101100110",
  25208=>"100011000",
  25209=>"111011000",
  25210=>"000111011",
  25211=>"001100001",
  25212=>"110011010",
  25213=>"010001111",
  25214=>"101111000",
  25215=>"111001110",
  25216=>"010000110",
  25217=>"110001110",
  25218=>"110110110",
  25219=>"010100110",
  25220=>"010111111",
  25221=>"010000101",
  25222=>"111000111",
  25223=>"101011001",
  25224=>"011110010",
  25225=>"010000010",
  25226=>"001101110",
  25227=>"000010101",
  25228=>"011000101",
  25229=>"011110111",
  25230=>"000111111",
  25231=>"010111110",
  25232=>"001010011",
  25233=>"000111110",
  25234=>"010010111",
  25235=>"110101011",
  25236=>"011000011",
  25237=>"011101100",
  25238=>"000011010",
  25239=>"111001001",
  25240=>"001000110",
  25241=>"011111010",
  25242=>"000010000",
  25243=>"101111010",
  25244=>"000000010",
  25245=>"100100101",
  25246=>"001100111",
  25247=>"110101111",
  25248=>"011000010",
  25249=>"100011100",
  25250=>"101011110",
  25251=>"001000101",
  25252=>"111101100",
  25253=>"101101111",
  25254=>"110000011",
  25255=>"101000000",
  25256=>"101011001",
  25257=>"101010100",
  25258=>"111001010",
  25259=>"100001100",
  25260=>"101111001",
  25261=>"010010001",
  25262=>"100011101",
  25263=>"110010100",
  25264=>"110100010",
  25265=>"010110100",
  25266=>"010000011",
  25267=>"100100010",
  25268=>"111110011",
  25269=>"001101100",
  25270=>"111110110",
  25271=>"100111111",
  25272=>"010001111",
  25273=>"110001100",
  25274=>"010010100",
  25275=>"001100001",
  25276=>"100001101",
  25277=>"100000110",
  25278=>"101110110",
  25279=>"011101010",
  25280=>"100000111",
  25281=>"000101100",
  25282=>"110010111",
  25283=>"111110100",
  25284=>"000001101",
  25285=>"001101001",
  25286=>"011011100",
  25287=>"111011100",
  25288=>"001100110",
  25289=>"110000000",
  25290=>"001110001",
  25291=>"011011010",
  25292=>"010100010",
  25293=>"111101001",
  25294=>"111011000",
  25295=>"010111110",
  25296=>"010010000",
  25297=>"011101111",
  25298=>"101101010",
  25299=>"110110000",
  25300=>"011111010",
  25301=>"111001000",
  25302=>"100100111",
  25303=>"110001111",
  25304=>"110111100",
  25305=>"010101111",
  25306=>"101111011",
  25307=>"110000101",
  25308=>"100101011",
  25309=>"011010110",
  25310=>"111101110",
  25311=>"010001011",
  25312=>"001111010",
  25313=>"001001110",
  25314=>"111110110",
  25315=>"100111000",
  25316=>"111011001",
  25317=>"111101110",
  25318=>"110010001",
  25319=>"000000011",
  25320=>"101100101",
  25321=>"011101110",
  25322=>"111101100",
  25323=>"111000001",
  25324=>"111111100",
  25325=>"010111101",
  25326=>"101110101",
  25327=>"000000000",
  25328=>"111100000",
  25329=>"001111111",
  25330=>"011001001",
  25331=>"001001111",
  25332=>"010101011",
  25333=>"010010010",
  25334=>"101110101",
  25335=>"100011001",
  25336=>"011110001",
  25337=>"011111000",
  25338=>"001001010",
  25339=>"001011100",
  25340=>"111110111",
  25341=>"100010111",
  25342=>"101100101",
  25343=>"110010110",
  25344=>"000000001",
  25345=>"100100011",
  25346=>"111011001",
  25347=>"000101100",
  25348=>"000000111",
  25349=>"001001010",
  25350=>"100100001",
  25351=>"001001101",
  25352=>"101101110",
  25353=>"011100001",
  25354=>"101001110",
  25355=>"000001101",
  25356=>"110100110",
  25357=>"111110000",
  25358=>"000110011",
  25359=>"111100000",
  25360=>"011011101",
  25361=>"100101110",
  25362=>"101001110",
  25363=>"000011011",
  25364=>"011101111",
  25365=>"100000110",
  25366=>"011011101",
  25367=>"110010110",
  25368=>"000011010",
  25369=>"000010100",
  25370=>"110001101",
  25371=>"001000101",
  25372=>"111010000",
  25373=>"110100101",
  25374=>"110000011",
  25375=>"010000110",
  25376=>"010000111",
  25377=>"101001011",
  25378=>"010101100",
  25379=>"101101010",
  25380=>"001111101",
  25381=>"010010111",
  25382=>"011110001",
  25383=>"010110110",
  25384=>"010100000",
  25385=>"101000000",
  25386=>"100111111",
  25387=>"001100001",
  25388=>"011100101",
  25389=>"010110101",
  25390=>"100010010",
  25391=>"010101110",
  25392=>"100110100",
  25393=>"101100110",
  25394=>"010100001",
  25395=>"000101011",
  25396=>"100101011",
  25397=>"100110010",
  25398=>"001111001",
  25399=>"000111101",
  25400=>"000111000",
  25401=>"000110011",
  25402=>"110010111",
  25403=>"001000001",
  25404=>"010111110",
  25405=>"010111101",
  25406=>"000111110",
  25407=>"010011001",
  25408=>"110001011",
  25409=>"010100000",
  25410=>"111011010",
  25411=>"000110000",
  25412=>"000100100",
  25413=>"010010111",
  25414=>"101111111",
  25415=>"111110001",
  25416=>"010011000",
  25417=>"110000000",
  25418=>"001101101",
  25419=>"000100110",
  25420=>"110101010",
  25421=>"111101001",
  25422=>"010010111",
  25423=>"101111111",
  25424=>"101111111",
  25425=>"010000010",
  25426=>"001010000",
  25427=>"010001001",
  25428=>"010101000",
  25429=>"111101100",
  25430=>"011001110",
  25431=>"111000110",
  25432=>"100000100",
  25433=>"110000100",
  25434=>"101111011",
  25435=>"001001100",
  25436=>"110110010",
  25437=>"011000000",
  25438=>"000100010",
  25439=>"000000000",
  25440=>"110011000",
  25441=>"110110010",
  25442=>"111010101",
  25443=>"101100000",
  25444=>"010111110",
  25445=>"100111000",
  25446=>"101100111",
  25447=>"101110001",
  25448=>"110001001",
  25449=>"001110011",
  25450=>"000001000",
  25451=>"000000111",
  25452=>"111010000",
  25453=>"000011100",
  25454=>"100101100",
  25455=>"001011001",
  25456=>"111110001",
  25457=>"000010100",
  25458=>"110110010",
  25459=>"010000000",
  25460=>"000011100",
  25461=>"000001000",
  25462=>"010010100",
  25463=>"001010100",
  25464=>"010111010",
  25465=>"100011001",
  25466=>"000111111",
  25467=>"001011110",
  25468=>"000100100",
  25469=>"111001100",
  25470=>"110100100",
  25471=>"100100001",
  25472=>"101010100",
  25473=>"111001001",
  25474=>"010010011",
  25475=>"111111111",
  25476=>"011111011",
  25477=>"100011100",
  25478=>"111101010",
  25479=>"111010000",
  25480=>"010110000",
  25481=>"100001010",
  25482=>"000111111",
  25483=>"000100100",
  25484=>"100100011",
  25485=>"010110101",
  25486=>"001011100",
  25487=>"110100000",
  25488=>"111001111",
  25489=>"100111101",
  25490=>"000011111",
  25491=>"011111000",
  25492=>"001100000",
  25493=>"110001011",
  25494=>"110111001",
  25495=>"001011100",
  25496=>"011000011",
  25497=>"010110101",
  25498=>"100000011",
  25499=>"100001110",
  25500=>"001001101",
  25501=>"011000011",
  25502=>"100101001",
  25503=>"011001001",
  25504=>"000111110",
  25505=>"001100110",
  25506=>"010010000",
  25507=>"101100101",
  25508=>"001100000",
  25509=>"001111111",
  25510=>"000011010",
  25511=>"000111101",
  25512=>"100110100",
  25513=>"000000010",
  25514=>"110001101",
  25515=>"010000000",
  25516=>"010100011",
  25517=>"100001001",
  25518=>"111001000",
  25519=>"110100001",
  25520=>"100000011",
  25521=>"100011000",
  25522=>"001000101",
  25523=>"001110001",
  25524=>"100110100",
  25525=>"110001000",
  25526=>"110010110",
  25527=>"010000010",
  25528=>"111001111",
  25529=>"111101011",
  25530=>"101110111",
  25531=>"001100100",
  25532=>"000011010",
  25533=>"101010000",
  25534=>"101110000",
  25535=>"100000110",
  25536=>"010110011",
  25537=>"100010111",
  25538=>"001110101",
  25539=>"001111110",
  25540=>"000000001",
  25541=>"101011001",
  25542=>"001110000",
  25543=>"101000010",
  25544=>"011001000",
  25545=>"011111010",
  25546=>"101101100",
  25547=>"011111111",
  25548=>"010110010",
  25549=>"111100000",
  25550=>"011011100",
  25551=>"011000110",
  25552=>"101111111",
  25553=>"111110011",
  25554=>"111000110",
  25555=>"000000010",
  25556=>"110000101",
  25557=>"011110011",
  25558=>"111011010",
  25559=>"101011101",
  25560=>"110111111",
  25561=>"110111110",
  25562=>"000000000",
  25563=>"110110100",
  25564=>"111011010",
  25565=>"100010001",
  25566=>"001011111",
  25567=>"001001010",
  25568=>"110011011",
  25569=>"100000100",
  25570=>"101001010",
  25571=>"101010100",
  25572=>"000110000",
  25573=>"110101111",
  25574=>"010011101",
  25575=>"111110000",
  25576=>"000011111",
  25577=>"000000110",
  25578=>"110000000",
  25579=>"000011111",
  25580=>"000100001",
  25581=>"000010100",
  25582=>"100101000",
  25583=>"011111110",
  25584=>"011110001",
  25585=>"001101100",
  25586=>"000110110",
  25587=>"111011001",
  25588=>"010100110",
  25589=>"100101011",
  25590=>"110011010",
  25591=>"111011011",
  25592=>"110101011",
  25593=>"101110100",
  25594=>"101111001",
  25595=>"011111110",
  25596=>"110110111",
  25597=>"100111100",
  25598=>"011001101",
  25599=>"010101110",
  25600=>"111111000",
  25601=>"101011011",
  25602=>"011100110",
  25603=>"111011101",
  25604=>"110100111",
  25605=>"101001000",
  25606=>"011011110",
  25607=>"001010011",
  25608=>"111001110",
  25609=>"110110101",
  25610=>"000001110",
  25611=>"110001011",
  25612=>"111111011",
  25613=>"011001100",
  25614=>"000100110",
  25615=>"011110000",
  25616=>"101011011",
  25617=>"000111100",
  25618=>"101011000",
  25619=>"000001011",
  25620=>"100100001",
  25621=>"100110101",
  25622=>"001000100",
  25623=>"100100011",
  25624=>"000100110",
  25625=>"011111000",
  25626=>"100101111",
  25627=>"011111010",
  25628=>"011111011",
  25629=>"001100110",
  25630=>"101100000",
  25631=>"111110111",
  25632=>"001101111",
  25633=>"110111101",
  25634=>"011100011",
  25635=>"001001100",
  25636=>"011001110",
  25637=>"000111100",
  25638=>"001000000",
  25639=>"111001110",
  25640=>"101101110",
  25641=>"101111100",
  25642=>"111001011",
  25643=>"111101011",
  25644=>"011110110",
  25645=>"101101000",
  25646=>"011000111",
  25647=>"001010010",
  25648=>"111100111",
  25649=>"001001001",
  25650=>"100000011",
  25651=>"111000000",
  25652=>"010101101",
  25653=>"000000111",
  25654=>"110110001",
  25655=>"100011011",
  25656=>"100101101",
  25657=>"001110000",
  25658=>"110111110",
  25659=>"010001001",
  25660=>"000100100",
  25661=>"101001000",
  25662=>"111001001",
  25663=>"101111010",
  25664=>"000100101",
  25665=>"010001000",
  25666=>"000100100",
  25667=>"101110111",
  25668=>"101000011",
  25669=>"000001101",
  25670=>"100110100",
  25671=>"000110010",
  25672=>"100100111",
  25673=>"001001000",
  25674=>"111011011",
  25675=>"000110111",
  25676=>"001110010",
  25677=>"000010010",
  25678=>"101001001",
  25679=>"100000010",
  25680=>"001100101",
  25681=>"001001110",
  25682=>"101000100",
  25683=>"010110110",
  25684=>"111000011",
  25685=>"000111101",
  25686=>"101011000",
  25687=>"011100111",
  25688=>"101100100",
  25689=>"011001010",
  25690=>"111100100",
  25691=>"110010001",
  25692=>"001101011",
  25693=>"111000101",
  25694=>"111000010",
  25695=>"011101010",
  25696=>"100111100",
  25697=>"110010011",
  25698=>"101000100",
  25699=>"001101100",
  25700=>"110100011",
  25701=>"111111110",
  25702=>"110001010",
  25703=>"110001000",
  25704=>"011011000",
  25705=>"000111101",
  25706=>"101100001",
  25707=>"111001110",
  25708=>"101111101",
  25709=>"101110111",
  25710=>"111111010",
  25711=>"010100011",
  25712=>"010010111",
  25713=>"001100010",
  25714=>"000001111",
  25715=>"111111110",
  25716=>"010111111",
  25717=>"001101110",
  25718=>"110111000",
  25719=>"000001100",
  25720=>"011011010",
  25721=>"101000100",
  25722=>"010110110",
  25723=>"001100101",
  25724=>"000111011",
  25725=>"110111100",
  25726=>"000011001",
  25727=>"110001110",
  25728=>"010000010",
  25729=>"011001100",
  25730=>"111101010",
  25731=>"100010011",
  25732=>"000100011",
  25733=>"010101100",
  25734=>"001100100",
  25735=>"101000111",
  25736=>"101101101",
  25737=>"010100101",
  25738=>"001000000",
  25739=>"011011100",
  25740=>"000010000",
  25741=>"101101111",
  25742=>"111111101",
  25743=>"110110011",
  25744=>"000110011",
  25745=>"101100110",
  25746=>"010001001",
  25747=>"111001111",
  25748=>"001000110",
  25749=>"100101010",
  25750=>"101000000",
  25751=>"010100101",
  25752=>"110110001",
  25753=>"011011100",
  25754=>"000100100",
  25755=>"010100001",
  25756=>"111110011",
  25757=>"111011110",
  25758=>"000101000",
  25759=>"001010111",
  25760=>"101010110",
  25761=>"101100110",
  25762=>"100010110",
  25763=>"100000011",
  25764=>"111111101",
  25765=>"010011010",
  25766=>"110101110",
  25767=>"010100100",
  25768=>"011101000",
  25769=>"110011010",
  25770=>"101001011",
  25771=>"001111010",
  25772=>"100000101",
  25773=>"000001000",
  25774=>"101110100",
  25775=>"110101111",
  25776=>"000011000",
  25777=>"000001000",
  25778=>"000110011",
  25779=>"100110111",
  25780=>"100100100",
  25781=>"010101001",
  25782=>"100000110",
  25783=>"001001101",
  25784=>"001010111",
  25785=>"101010010",
  25786=>"101101111",
  25787=>"110010111",
  25788=>"011101001",
  25789=>"000100000",
  25790=>"110101111",
  25791=>"110110000",
  25792=>"000111011",
  25793=>"001011111",
  25794=>"000000000",
  25795=>"101101000",
  25796=>"111111111",
  25797=>"010001100",
  25798=>"010100001",
  25799=>"000101011",
  25800=>"011111001",
  25801=>"111111010",
  25802=>"110001101",
  25803=>"111110000",
  25804=>"100000010",
  25805=>"111101011",
  25806=>"100110001",
  25807=>"111000010",
  25808=>"100101101",
  25809=>"000000010",
  25810=>"111011010",
  25811=>"000011001",
  25812=>"010100101",
  25813=>"000110001",
  25814=>"001011101",
  25815=>"000010000",
  25816=>"100011100",
  25817=>"111110001",
  25818=>"011100101",
  25819=>"110001000",
  25820=>"000011001",
  25821=>"011111111",
  25822=>"100101000",
  25823=>"111111001",
  25824=>"001100100",
  25825=>"001010110",
  25826=>"011100001",
  25827=>"001110101",
  25828=>"010000000",
  25829=>"110101010",
  25830=>"100011000",
  25831=>"011001111",
  25832=>"110001000",
  25833=>"101010001",
  25834=>"001011001",
  25835=>"110101110",
  25836=>"100111101",
  25837=>"101100000",
  25838=>"000100011",
  25839=>"010000010",
  25840=>"010111100",
  25841=>"011000111",
  25842=>"100000110",
  25843=>"000010111",
  25844=>"100001111",
  25845=>"001010010",
  25846=>"110111000",
  25847=>"011100000",
  25848=>"101111100",
  25849=>"110001111",
  25850=>"001001000",
  25851=>"001100001",
  25852=>"011111101",
  25853=>"111001011",
  25854=>"100111101",
  25855=>"111111101",
  25856=>"001101010",
  25857=>"010010010",
  25858=>"101100110",
  25859=>"000011000",
  25860=>"010010011",
  25861=>"100111011",
  25862=>"000101111",
  25863=>"011111111",
  25864=>"101001101",
  25865=>"010100001",
  25866=>"100011000",
  25867=>"100111001",
  25868=>"001010001",
  25869=>"111110110",
  25870=>"011111001",
  25871=>"010010011",
  25872=>"100011000",
  25873=>"010001111",
  25874=>"011011000",
  25875=>"101111100",
  25876=>"101011011",
  25877=>"011101100",
  25878=>"000001111",
  25879=>"000101010",
  25880=>"111100001",
  25881=>"001111001",
  25882=>"100110001",
  25883=>"010010101",
  25884=>"111100011",
  25885=>"111010000",
  25886=>"011110011",
  25887=>"110111111",
  25888=>"101000000",
  25889=>"110010111",
  25890=>"101101110",
  25891=>"100111011",
  25892=>"110001111",
  25893=>"101100100",
  25894=>"011101010",
  25895=>"110001010",
  25896=>"001000010",
  25897=>"011000011",
  25898=>"011111011",
  25899=>"010001001",
  25900=>"001000111",
  25901=>"001110011",
  25902=>"111110000",
  25903=>"001100101",
  25904=>"011101011",
  25905=>"000001110",
  25906=>"001101101",
  25907=>"101111001",
  25908=>"010101110",
  25909=>"110010011",
  25910=>"001101000",
  25911=>"011110000",
  25912=>"000001101",
  25913=>"110000000",
  25914=>"001001000",
  25915=>"110011011",
  25916=>"001100111",
  25917=>"010000011",
  25918=>"111000100",
  25919=>"011011100",
  25920=>"001100010",
  25921=>"111011101",
  25922=>"010100100",
  25923=>"111101010",
  25924=>"001011011",
  25925=>"110101010",
  25926=>"000000010",
  25927=>"100010100",
  25928=>"101001101",
  25929=>"000010100",
  25930=>"101001001",
  25931=>"111111000",
  25932=>"110101011",
  25933=>"000101001",
  25934=>"101001000",
  25935=>"000011110",
  25936=>"011100110",
  25937=>"101010000",
  25938=>"101001111",
  25939=>"000100010",
  25940=>"010100010",
  25941=>"011111010",
  25942=>"100010100",
  25943=>"111010001",
  25944=>"111110001",
  25945=>"011101110",
  25946=>"101101101",
  25947=>"011100000",
  25948=>"101110000",
  25949=>"010111100",
  25950=>"100000000",
  25951=>"100001011",
  25952=>"100000011",
  25953=>"011010110",
  25954=>"101000110",
  25955=>"011000000",
  25956=>"011010001",
  25957=>"011010010",
  25958=>"001010001",
  25959=>"001010011",
  25960=>"001001010",
  25961=>"110110000",
  25962=>"000111101",
  25963=>"000100111",
  25964=>"001010100",
  25965=>"000001101",
  25966=>"111011101",
  25967=>"011101010",
  25968=>"111010111",
  25969=>"001110000",
  25970=>"010000111",
  25971=>"000101100",
  25972=>"100110110",
  25973=>"100000110",
  25974=>"100111101",
  25975=>"001100110",
  25976=>"100110010",
  25977=>"011010111",
  25978=>"110100010",
  25979=>"111000001",
  25980=>"111011101",
  25981=>"011111001",
  25982=>"010110111",
  25983=>"101101101",
  25984=>"010010011",
  25985=>"110110101",
  25986=>"011110110",
  25987=>"000100100",
  25988=>"100111000",
  25989=>"001010001",
  25990=>"010111111",
  25991=>"001000000",
  25992=>"111100001",
  25993=>"000000101",
  25994=>"001000111",
  25995=>"000010100",
  25996=>"110100100",
  25997=>"100100101",
  25998=>"000000010",
  25999=>"011011101",
  26000=>"011010011",
  26001=>"111110011",
  26002=>"001100100",
  26003=>"010000000",
  26004=>"010101001",
  26005=>"111101000",
  26006=>"111000011",
  26007=>"111011100",
  26008=>"011100000",
  26009=>"010110111",
  26010=>"000011011",
  26011=>"101001100",
  26012=>"110111000",
  26013=>"001011111",
  26014=>"111011110",
  26015=>"001001110",
  26016=>"100111110",
  26017=>"100101000",
  26018=>"001110000",
  26019=>"100110011",
  26020=>"011010000",
  26021=>"011111001",
  26022=>"111111100",
  26023=>"110111100",
  26024=>"111010100",
  26025=>"111001110",
  26026=>"110000101",
  26027=>"110111101",
  26028=>"011000011",
  26029=>"010001110",
  26030=>"000010010",
  26031=>"110010111",
  26032=>"000111111",
  26033=>"100101011",
  26034=>"011110111",
  26035=>"011001011",
  26036=>"000011110",
  26037=>"111000011",
  26038=>"011110000",
  26039=>"100101001",
  26040=>"100010100",
  26041=>"000010110",
  26042=>"010111101",
  26043=>"110111110",
  26044=>"110010011",
  26045=>"000100000",
  26046=>"111110011",
  26047=>"110111110",
  26048=>"101011100",
  26049=>"011000101",
  26050=>"001110100",
  26051=>"011000011",
  26052=>"010011100",
  26053=>"000100011",
  26054=>"001010101",
  26055=>"001110010",
  26056=>"111011000",
  26057=>"100001001",
  26058=>"100100001",
  26059=>"001101000",
  26060=>"011000100",
  26061=>"111001000",
  26062=>"100111110",
  26063=>"000101111",
  26064=>"111000101",
  26065=>"001110110",
  26066=>"101100001",
  26067=>"010001100",
  26068=>"101011001",
  26069=>"000111110",
  26070=>"100100000",
  26071=>"000010001",
  26072=>"000110000",
  26073=>"111111010",
  26074=>"001001011",
  26075=>"101000001",
  26076=>"101100100",
  26077=>"100110111",
  26078=>"101011100",
  26079=>"011001101",
  26080=>"011100000",
  26081=>"100000010",
  26082=>"010111110",
  26083=>"110000001",
  26084=>"000100111",
  26085=>"001000001",
  26086=>"011111101",
  26087=>"101111101",
  26088=>"010111100",
  26089=>"110110001",
  26090=>"100001010",
  26091=>"111111111",
  26092=>"001110100",
  26093=>"110000010",
  26094=>"100001011",
  26095=>"010101111",
  26096=>"101111100",
  26097=>"001100110",
  26098=>"101000111",
  26099=>"000110110",
  26100=>"111110011",
  26101=>"110101111",
  26102=>"000111001",
  26103=>"100011000",
  26104=>"011101000",
  26105=>"111000011",
  26106=>"000111001",
  26107=>"000111010",
  26108=>"000110110",
  26109=>"100000101",
  26110=>"110110110",
  26111=>"101011101",
  26112=>"110001010",
  26113=>"011011000",
  26114=>"100110010",
  26115=>"000001100",
  26116=>"101111100",
  26117=>"000110000",
  26118=>"110111100",
  26119=>"100111000",
  26120=>"000111111",
  26121=>"110111001",
  26122=>"000000110",
  26123=>"000011000",
  26124=>"000110111",
  26125=>"110111111",
  26126=>"001010100",
  26127=>"110001110",
  26128=>"111010000",
  26129=>"100011101",
  26130=>"000010100",
  26131=>"011111010",
  26132=>"111110111",
  26133=>"110010010",
  26134=>"100110111",
  26135=>"110100101",
  26136=>"011010010",
  26137=>"000111000",
  26138=>"000010111",
  26139=>"111011010",
  26140=>"011100111",
  26141=>"111111000",
  26142=>"100011100",
  26143=>"110111000",
  26144=>"001011110",
  26145=>"111101111",
  26146=>"101010010",
  26147=>"001010000",
  26148=>"001001000",
  26149=>"101010000",
  26150=>"101010011",
  26151=>"000000001",
  26152=>"101000100",
  26153=>"110101110",
  26154=>"110100110",
  26155=>"010111110",
  26156=>"100101100",
  26157=>"110111101",
  26158=>"000001000",
  26159=>"010111010",
  26160=>"110000000",
  26161=>"000001001",
  26162=>"001011000",
  26163=>"000001101",
  26164=>"000010110",
  26165=>"001111110",
  26166=>"111000010",
  26167=>"001010001",
  26168=>"001001100",
  26169=>"101011101",
  26170=>"100001011",
  26171=>"011011000",
  26172=>"101011010",
  26173=>"010011110",
  26174=>"101001111",
  26175=>"110110000",
  26176=>"110011101",
  26177=>"001111110",
  26178=>"011101111",
  26179=>"001101101",
  26180=>"101111101",
  26181=>"110100111",
  26182=>"010111110",
  26183=>"011010011",
  26184=>"011111000",
  26185=>"011110110",
  26186=>"101100101",
  26187=>"101001000",
  26188=>"001000000",
  26189=>"011000000",
  26190=>"111110101",
  26191=>"101011100",
  26192=>"010110001",
  26193=>"111011000",
  26194=>"101110010",
  26195=>"000000011",
  26196=>"110010001",
  26197=>"110000001",
  26198=>"011000111",
  26199=>"101101000",
  26200=>"000001111",
  26201=>"000000101",
  26202=>"100101011",
  26203=>"100000101",
  26204=>"001001110",
  26205=>"111010100",
  26206=>"000001011",
  26207=>"100000011",
  26208=>"011010101",
  26209=>"011011100",
  26210=>"001111000",
  26211=>"010011011",
  26212=>"011010000",
  26213=>"000101000",
  26214=>"011100111",
  26215=>"011011001",
  26216=>"001101111",
  26217=>"100101011",
  26218=>"100111000",
  26219=>"001111100",
  26220=>"000010001",
  26221=>"001111001",
  26222=>"110011110",
  26223=>"011100011",
  26224=>"110110010",
  26225=>"111110011",
  26226=>"000110101",
  26227=>"101101110",
  26228=>"100001010",
  26229=>"110100000",
  26230=>"001010110",
  26231=>"001000000",
  26232=>"011111100",
  26233=>"001111001",
  26234=>"011001011",
  26235=>"100111110",
  26236=>"000111100",
  26237=>"100010000",
  26238=>"110101110",
  26239=>"001110010",
  26240=>"100101100",
  26241=>"100001011",
  26242=>"000101111",
  26243=>"110010100",
  26244=>"010111111",
  26245=>"010000100",
  26246=>"100110111",
  26247=>"011001001",
  26248=>"100000111",
  26249=>"001000110",
  26250=>"011010011",
  26251=>"011101011",
  26252=>"000001010",
  26253=>"010101001",
  26254=>"100001010",
  26255=>"101010010",
  26256=>"111000010",
  26257=>"001011000",
  26258=>"000100011",
  26259=>"001101011",
  26260=>"000110010",
  26261=>"001000010",
  26262=>"000101000",
  26263=>"101100101",
  26264=>"001101010",
  26265=>"110000011",
  26266=>"101111100",
  26267=>"101111000",
  26268=>"111001100",
  26269=>"100100010",
  26270=>"010100000",
  26271=>"000101110",
  26272=>"000111111",
  26273=>"101010101",
  26274=>"010011101",
  26275=>"100100001",
  26276=>"100100111",
  26277=>"011000110",
  26278=>"100111000",
  26279=>"100000001",
  26280=>"001000110",
  26281=>"101111011",
  26282=>"011000111",
  26283=>"110110000",
  26284=>"110010110",
  26285=>"100000011",
  26286=>"100000110",
  26287=>"101001000",
  26288=>"000100011",
  26289=>"100110100",
  26290=>"010110010",
  26291=>"001110100",
  26292=>"001101111",
  26293=>"101001011",
  26294=>"000001110",
  26295=>"111010100",
  26296=>"101101000",
  26297=>"010100001",
  26298=>"111010011",
  26299=>"010101111",
  26300=>"000001001",
  26301=>"111001111",
  26302=>"010000111",
  26303=>"010101010",
  26304=>"101100100",
  26305=>"000000110",
  26306=>"101101111",
  26307=>"110111001",
  26308=>"010001010",
  26309=>"001001101",
  26310=>"001001100",
  26311=>"111101100",
  26312=>"011111011",
  26313=>"101110001",
  26314=>"101010100",
  26315=>"001010000",
  26316=>"100101011",
  26317=>"111111111",
  26318=>"110000010",
  26319=>"011010100",
  26320=>"110001101",
  26321=>"110011001",
  26322=>"100001110",
  26323=>"011101101",
  26324=>"100011101",
  26325=>"011000011",
  26326=>"011110111",
  26327=>"100110100",
  26328=>"110000000",
  26329=>"111100000",
  26330=>"101001101",
  26331=>"100010001",
  26332=>"011001110",
  26333=>"000110000",
  26334=>"010010110",
  26335=>"101000010",
  26336=>"111111111",
  26337=>"010100010",
  26338=>"101110100",
  26339=>"101110010",
  26340=>"011001101",
  26341=>"101111101",
  26342=>"101011001",
  26343=>"111100011",
  26344=>"011010101",
  26345=>"000000000",
  26346=>"111101010",
  26347=>"101000011",
  26348=>"000011001",
  26349=>"100000111",
  26350=>"000011000",
  26351=>"101110000",
  26352=>"100100010",
  26353=>"000100011",
  26354=>"001111110",
  26355=>"111111100",
  26356=>"001001100",
  26357=>"100000010",
  26358=>"101110011",
  26359=>"011110000",
  26360=>"011111111",
  26361=>"010000000",
  26362=>"111000000",
  26363=>"111010111",
  26364=>"100010001",
  26365=>"000101110",
  26366=>"101010110",
  26367=>"011010000",
  26368=>"110101101",
  26369=>"100100011",
  26370=>"101010011",
  26371=>"000001110",
  26372=>"110011010",
  26373=>"101111110",
  26374=>"011100010",
  26375=>"110011001",
  26376=>"010000010",
  26377=>"110010110",
  26378=>"111011001",
  26379=>"010111000",
  26380=>"011011111",
  26381=>"110010010",
  26382=>"000101101",
  26383=>"111111101",
  26384=>"001111010",
  26385=>"010010011",
  26386=>"010111111",
  26387=>"100110000",
  26388=>"001111101",
  26389=>"111001110",
  26390=>"111011100",
  26391=>"011010100",
  26392=>"100001001",
  26393=>"101011100",
  26394=>"101000000",
  26395=>"101110010",
  26396=>"001000100",
  26397=>"110000110",
  26398=>"011101100",
  26399=>"100000000",
  26400=>"101000101",
  26401=>"001111000",
  26402=>"000111000",
  26403=>"011101000",
  26404=>"100101010",
  26405=>"100100010",
  26406=>"001010100",
  26407=>"001101100",
  26408=>"111100000",
  26409=>"100000111",
  26410=>"110001110",
  26411=>"110101100",
  26412=>"101010100",
  26413=>"010111100",
  26414=>"100101000",
  26415=>"101011101",
  26416=>"111011010",
  26417=>"111100101",
  26418=>"101111101",
  26419=>"110111111",
  26420=>"010100000",
  26421=>"100110100",
  26422=>"100111111",
  26423=>"100011100",
  26424=>"111011001",
  26425=>"111000010",
  26426=>"001111101",
  26427=>"111011110",
  26428=>"000110110",
  26429=>"100010110",
  26430=>"000000101",
  26431=>"110111000",
  26432=>"100001010",
  26433=>"101110001",
  26434=>"001111111",
  26435=>"000111110",
  26436=>"111000100",
  26437=>"010110110",
  26438=>"100001010",
  26439=>"010000101",
  26440=>"000011111",
  26441=>"000011100",
  26442=>"111011111",
  26443=>"010100010",
  26444=>"001100000",
  26445=>"101111101",
  26446=>"010010010",
  26447=>"111000011",
  26448=>"110110110",
  26449=>"110110111",
  26450=>"001101101",
  26451=>"110110100",
  26452=>"101100010",
  26453=>"011001110",
  26454=>"000001111",
  26455=>"110001000",
  26456=>"100101000",
  26457=>"011100110",
  26458=>"100101000",
  26459=>"000010101",
  26460=>"111111000",
  26461=>"001101011",
  26462=>"111111011",
  26463=>"000011101",
  26464=>"110100110",
  26465=>"000011011",
  26466=>"000010110",
  26467=>"110110100",
  26468=>"100010000",
  26469=>"011010101",
  26470=>"011010101",
  26471=>"110110100",
  26472=>"000001000",
  26473=>"001101000",
  26474=>"101011000",
  26475=>"011010010",
  26476=>"111011001",
  26477=>"110000010",
  26478=>"000100111",
  26479=>"101000111",
  26480=>"110110101",
  26481=>"000110011",
  26482=>"101001001",
  26483=>"001010101",
  26484=>"110100010",
  26485=>"101010101",
  26486=>"101111111",
  26487=>"001000101",
  26488=>"101111111",
  26489=>"111011100",
  26490=>"100000101",
  26491=>"011100001",
  26492=>"010110011",
  26493=>"010110110",
  26494=>"101100001",
  26495=>"011011111",
  26496=>"010010011",
  26497=>"010100001",
  26498=>"111110010",
  26499=>"110010110",
  26500=>"111000010",
  26501=>"111000010",
  26502=>"100101001",
  26503=>"000110000",
  26504=>"110000011",
  26505=>"001111110",
  26506=>"111101110",
  26507=>"000101100",
  26508=>"110101010",
  26509=>"010010001",
  26510=>"000101100",
  26511=>"010110100",
  26512=>"000111111",
  26513=>"011111010",
  26514=>"100000100",
  26515=>"111000011",
  26516=>"011110000",
  26517=>"001001000",
  26518=>"010010110",
  26519=>"000111100",
  26520=>"100111110",
  26521=>"000110000",
  26522=>"010100111",
  26523=>"001100011",
  26524=>"110100001",
  26525=>"111101011",
  26526=>"011000111",
  26527=>"000111010",
  26528=>"001011010",
  26529=>"111101101",
  26530=>"001001111",
  26531=>"111101001",
  26532=>"010011010",
  26533=>"100101011",
  26534=>"001101001",
  26535=>"110010001",
  26536=>"000001111",
  26537=>"001000111",
  26538=>"001011111",
  26539=>"101001110",
  26540=>"001011110",
  26541=>"001111011",
  26542=>"000101011",
  26543=>"001111010",
  26544=>"011010001",
  26545=>"011100010",
  26546=>"100111000",
  26547=>"000111111",
  26548=>"001101001",
  26549=>"001100101",
  26550=>"011101110",
  26551=>"110010011",
  26552=>"111100100",
  26553=>"011000010",
  26554=>"010100101",
  26555=>"010100000",
  26556=>"011101001",
  26557=>"101111111",
  26558=>"100001100",
  26559=>"110011111",
  26560=>"000100100",
  26561=>"100011100",
  26562=>"000010101",
  26563=>"111011011",
  26564=>"000101010",
  26565=>"001010101",
  26566=>"111101001",
  26567=>"000011001",
  26568=>"110011001",
  26569=>"011011011",
  26570=>"101000100",
  26571=>"011110110",
  26572=>"000000111",
  26573=>"000111110",
  26574=>"011010010",
  26575=>"000000001",
  26576=>"101100000",
  26577=>"001100010",
  26578=>"111001010",
  26579=>"000101110",
  26580=>"001001000",
  26581=>"111101001",
  26582=>"101001111",
  26583=>"011101110",
  26584=>"000111111",
  26585=>"000111111",
  26586=>"100110001",
  26587=>"111011000",
  26588=>"101101100",
  26589=>"011100011",
  26590=>"101101001",
  26591=>"100000100",
  26592=>"000110111",
  26593=>"100010010",
  26594=>"100001010",
  26595=>"000100011",
  26596=>"011101111",
  26597=>"010011110",
  26598=>"100010100",
  26599=>"101110000",
  26600=>"000101000",
  26601=>"111011111",
  26602=>"110101100",
  26603=>"000111101",
  26604=>"111110111",
  26605=>"101101111",
  26606=>"011110010",
  26607=>"100110101",
  26608=>"100101111",
  26609=>"100110100",
  26610=>"011011111",
  26611=>"111110110",
  26612=>"101010110",
  26613=>"101100001",
  26614=>"000110111",
  26615=>"001001001",
  26616=>"000101100",
  26617=>"110110010",
  26618=>"010011101",
  26619=>"011100011",
  26620=>"110101101",
  26621=>"001011110",
  26622=>"000111010",
  26623=>"101100101",
  26624=>"001000111",
  26625=>"000111001",
  26626=>"010001001",
  26627=>"110101111",
  26628=>"111000110",
  26629=>"100000001",
  26630=>"000011000",
  26631=>"110111111",
  26632=>"000011101",
  26633=>"010110100",
  26634=>"101001011",
  26635=>"100101010",
  26636=>"111010000",
  26637=>"010111011",
  26638=>"001000111",
  26639=>"101111001",
  26640=>"000000111",
  26641=>"110001111",
  26642=>"100110110",
  26643=>"101101110",
  26644=>"001110100",
  26645=>"100000110",
  26646=>"000100011",
  26647=>"011011110",
  26648=>"011111101",
  26649=>"010011000",
  26650=>"111011111",
  26651=>"010010101",
  26652=>"001001101",
  26653=>"110100010",
  26654=>"010000000",
  26655=>"000011011",
  26656=>"111001000",
  26657=>"010001000",
  26658=>"100110011",
  26659=>"001111100",
  26660=>"010111101",
  26661=>"110110010",
  26662=>"100100010",
  26663=>"010011010",
  26664=>"000010011",
  26665=>"111001111",
  26666=>"101100110",
  26667=>"111000100",
  26668=>"110110011",
  26669=>"010101111",
  26670=>"100000100",
  26671=>"111000000",
  26672=>"001110111",
  26673=>"100000100",
  26674=>"110110110",
  26675=>"011010101",
  26676=>"100110011",
  26677=>"001111110",
  26678=>"000001010",
  26679=>"111110110",
  26680=>"010100011",
  26681=>"110011000",
  26682=>"001111100",
  26683=>"111001011",
  26684=>"101110101",
  26685=>"001010010",
  26686=>"110110100",
  26687=>"110010100",
  26688=>"100111100",
  26689=>"111101001",
  26690=>"010000101",
  26691=>"001001110",
  26692=>"001100001",
  26693=>"101100011",
  26694=>"010110100",
  26695=>"010100100",
  26696=>"100001111",
  26697=>"000100000",
  26698=>"111011111",
  26699=>"101111011",
  26700=>"111011110",
  26701=>"010101001",
  26702=>"000001110",
  26703=>"100111110",
  26704=>"110101111",
  26705=>"011001011",
  26706=>"101001110",
  26707=>"001011001",
  26708=>"010001100",
  26709=>"000101010",
  26710=>"100001011",
  26711=>"111111111",
  26712=>"111110011",
  26713=>"111001000",
  26714=>"101000001",
  26715=>"000100100",
  26716=>"000011101",
  26717=>"110000010",
  26718=>"101000100",
  26719=>"011000001",
  26720=>"111100101",
  26721=>"111011010",
  26722=>"110010010",
  26723=>"000101111",
  26724=>"100100010",
  26725=>"100011000",
  26726=>"000011111",
  26727=>"111010011",
  26728=>"110010010",
  26729=>"001101010",
  26730=>"011111011",
  26731=>"000110010",
  26732=>"101101100",
  26733=>"101110101",
  26734=>"001110010",
  26735=>"011000011",
  26736=>"010001011",
  26737=>"111101111",
  26738=>"011000111",
  26739=>"000110101",
  26740=>"001111000",
  26741=>"010110000",
  26742=>"111010011",
  26743=>"000100100",
  26744=>"000101101",
  26745=>"101110110",
  26746=>"110110111",
  26747=>"001011000",
  26748=>"010111010",
  26749=>"100101001",
  26750=>"000001110",
  26751=>"101001010",
  26752=>"001000010",
  26753=>"110001100",
  26754=>"110100011",
  26755=>"110001011",
  26756=>"000000001",
  26757=>"001111111",
  26758=>"100000000",
  26759=>"000101011",
  26760=>"000111001",
  26761=>"110100110",
  26762=>"101100100",
  26763=>"111110111",
  26764=>"000111110",
  26765=>"101000100",
  26766=>"000100100",
  26767=>"101111011",
  26768=>"101010000",
  26769=>"001100001",
  26770=>"011010110",
  26771=>"111110010",
  26772=>"000000011",
  26773=>"011100100",
  26774=>"001010001",
  26775=>"000011100",
  26776=>"100111001",
  26777=>"000001011",
  26778=>"001011100",
  26779=>"110100110",
  26780=>"101111000",
  26781=>"000011000",
  26782=>"010011000",
  26783=>"010001110",
  26784=>"010001011",
  26785=>"111011000",
  26786=>"011010000",
  26787=>"010110011",
  26788=>"100101000",
  26789=>"001101111",
  26790=>"011110000",
  26791=>"011111100",
  26792=>"101010011",
  26793=>"100111000",
  26794=>"101010101",
  26795=>"000000000",
  26796=>"001101011",
  26797=>"101101101",
  26798=>"110100001",
  26799=>"010110111",
  26800=>"101010110",
  26801=>"010001000",
  26802=>"101110100",
  26803=>"001110110",
  26804=>"001110101",
  26805=>"111011101",
  26806=>"011010011",
  26807=>"000000000",
  26808=>"100010001",
  26809=>"110011111",
  26810=>"111010000",
  26811=>"000111101",
  26812=>"101101110",
  26813=>"111001111",
  26814=>"001111101",
  26815=>"101010100",
  26816=>"001000111",
  26817=>"110010111",
  26818=>"110010101",
  26819=>"111111011",
  26820=>"111001100",
  26821=>"110000011",
  26822=>"101110101",
  26823=>"011000011",
  26824=>"110101111",
  26825=>"010100111",
  26826=>"000011000",
  26827=>"110100110",
  26828=>"101000100",
  26829=>"100101011",
  26830=>"111000000",
  26831=>"001010100",
  26832=>"010001101",
  26833=>"010010110",
  26834=>"111001011",
  26835=>"001001100",
  26836=>"010000101",
  26837=>"101001101",
  26838=>"110111000",
  26839=>"110000000",
  26840=>"101011111",
  26841=>"010101010",
  26842=>"100100001",
  26843=>"010100000",
  26844=>"101111100",
  26845=>"010000100",
  26846=>"001111111",
  26847=>"111110101",
  26848=>"000011000",
  26849=>"011110000",
  26850=>"100010001",
  26851=>"001101010",
  26852=>"100010111",
  26853=>"111001111",
  26854=>"111001111",
  26855=>"011011111",
  26856=>"111110111",
  26857=>"100110000",
  26858=>"100110010",
  26859=>"010101011",
  26860=>"110101010",
  26861=>"111101000",
  26862=>"101100100",
  26863=>"111001111",
  26864=>"110100001",
  26865=>"001111000",
  26866=>"011110000",
  26867=>"011111001",
  26868=>"001010100",
  26869=>"001011111",
  26870=>"100011000",
  26871=>"111100101",
  26872=>"100010110",
  26873=>"110000011",
  26874=>"011011011",
  26875=>"000110101",
  26876=>"001010111",
  26877=>"100000010",
  26878=>"111111111",
  26879=>"111111101",
  26880=>"110000100",
  26881=>"000000111",
  26882=>"001011111",
  26883=>"101010001",
  26884=>"001100000",
  26885=>"011001001",
  26886=>"101011001",
  26887=>"110010100",
  26888=>"011010110",
  26889=>"111101011",
  26890=>"101110100",
  26891=>"110010100",
  26892=>"011000001",
  26893=>"001101111",
  26894=>"101111011",
  26895=>"111011000",
  26896=>"010011111",
  26897=>"001101010",
  26898=>"100111011",
  26899=>"100101111",
  26900=>"100000110",
  26901=>"000001011",
  26902=>"010100001",
  26903=>"101010110",
  26904=>"110000110",
  26905=>"011101100",
  26906=>"000000010",
  26907=>"001101001",
  26908=>"110100110",
  26909=>"011100110",
  26910=>"010000000",
  26911=>"101111001",
  26912=>"000010101",
  26913=>"001111110",
  26914=>"101011111",
  26915=>"100111011",
  26916=>"010110101",
  26917=>"111011111",
  26918=>"000011001",
  26919=>"111010010",
  26920=>"110001000",
  26921=>"111000000",
  26922=>"111110000",
  26923=>"111111001",
  26924=>"100010111",
  26925=>"000000101",
  26926=>"110000101",
  26927=>"001000111",
  26928=>"001110010",
  26929=>"000000001",
  26930=>"100010000",
  26931=>"100101111",
  26932=>"111000001",
  26933=>"011000000",
  26934=>"001101101",
  26935=>"101001100",
  26936=>"110111110",
  26937=>"111101100",
  26938=>"001111111",
  26939=>"000101011",
  26940=>"000010111",
  26941=>"001000001",
  26942=>"011001011",
  26943=>"101001101",
  26944=>"111000011",
  26945=>"110101010",
  26946=>"011011001",
  26947=>"110111011",
  26948=>"010100110",
  26949=>"101111111",
  26950=>"110110011",
  26951=>"110100001",
  26952=>"001001000",
  26953=>"000000010",
  26954=>"111011100",
  26955=>"110111001",
  26956=>"111000000",
  26957=>"110100101",
  26958=>"000101011",
  26959=>"110111101",
  26960=>"111101001",
  26961=>"001110010",
  26962=>"011111101",
  26963=>"111011010",
  26964=>"111011011",
  26965=>"110110111",
  26966=>"110001011",
  26967=>"100101100",
  26968=>"010100110",
  26969=>"010101111",
  26970=>"111011111",
  26971=>"010000010",
  26972=>"110111110",
  26973=>"101100001",
  26974=>"110110000",
  26975=>"000110101",
  26976=>"101111001",
  26977=>"100000101",
  26978=>"101000111",
  26979=>"110100111",
  26980=>"100110111",
  26981=>"011111100",
  26982=>"011100110",
  26983=>"011001010",
  26984=>"011011111",
  26985=>"001101111",
  26986=>"101010110",
  26987=>"101110111",
  26988=>"111001010",
  26989=>"010011111",
  26990=>"111001100",
  26991=>"110101111",
  26992=>"101100011",
  26993=>"011110000",
  26994=>"110000011",
  26995=>"000011111",
  26996=>"010000111",
  26997=>"001001111",
  26998=>"011100001",
  26999=>"111101101",
  27000=>"101100110",
  27001=>"011001011",
  27002=>"001001100",
  27003=>"011011110",
  27004=>"110010000",
  27005=>"100111111",
  27006=>"011101011",
  27007=>"000011011",
  27008=>"110111000",
  27009=>"000010011",
  27010=>"110011110",
  27011=>"001011111",
  27012=>"011001100",
  27013=>"001100101",
  27014=>"001111111",
  27015=>"000010000",
  27016=>"101001111",
  27017=>"000110100",
  27018=>"011011011",
  27019=>"010000011",
  27020=>"110001011",
  27021=>"010111011",
  27022=>"000100001",
  27023=>"100001111",
  27024=>"111010011",
  27025=>"101101000",
  27026=>"011110101",
  27027=>"011100100",
  27028=>"101101010",
  27029=>"101100100",
  27030=>"010011011",
  27031=>"100000100",
  27032=>"100010100",
  27033=>"011010010",
  27034=>"000111101",
  27035=>"000010010",
  27036=>"010010001",
  27037=>"111000011",
  27038=>"010100111",
  27039=>"011001001",
  27040=>"111111011",
  27041=>"111000000",
  27042=>"111110010",
  27043=>"000010001",
  27044=>"011000100",
  27045=>"001111110",
  27046=>"100000110",
  27047=>"001001101",
  27048=>"000100100",
  27049=>"011001010",
  27050=>"111001111",
  27051=>"110011100",
  27052=>"111111101",
  27053=>"110111011",
  27054=>"010001111",
  27055=>"011111100",
  27056=>"101011000",
  27057=>"001111010",
  27058=>"001100110",
  27059=>"111110111",
  27060=>"001010001",
  27061=>"011010001",
  27062=>"100101101",
  27063=>"110001000",
  27064=>"111010100",
  27065=>"001111111",
  27066=>"101011110",
  27067=>"010010010",
  27068=>"010010100",
  27069=>"010000010",
  27070=>"000011111",
  27071=>"111100100",
  27072=>"100001000",
  27073=>"111010101",
  27074=>"011010011",
  27075=>"101000010",
  27076=>"001000010",
  27077=>"100010101",
  27078=>"100110111",
  27079=>"100000000",
  27080=>"110101111",
  27081=>"101011111",
  27082=>"101000000",
  27083=>"001110011",
  27084=>"111010001",
  27085=>"110011101",
  27086=>"100101000",
  27087=>"000101101",
  27088=>"010011101",
  27089=>"011000011",
  27090=>"111110010",
  27091=>"001101100",
  27092=>"110000000",
  27093=>"010111011",
  27094=>"000001001",
  27095=>"010010010",
  27096=>"101100011",
  27097=>"101110100",
  27098=>"010010111",
  27099=>"001011010",
  27100=>"011010001",
  27101=>"001111100",
  27102=>"110110000",
  27103=>"010010011",
  27104=>"100001010",
  27105=>"110100100",
  27106=>"000110011",
  27107=>"111101100",
  27108=>"111100001",
  27109=>"111100010",
  27110=>"011011000",
  27111=>"101011000",
  27112=>"100010000",
  27113=>"111001011",
  27114=>"110101010",
  27115=>"010100100",
  27116=>"101011101",
  27117=>"001001000",
  27118=>"010101011",
  27119=>"100100111",
  27120=>"001010110",
  27121=>"111000010",
  27122=>"011110000",
  27123=>"001000111",
  27124=>"100010110",
  27125=>"000111001",
  27126=>"100110111",
  27127=>"001000111",
  27128=>"101001110",
  27129=>"101001010",
  27130=>"011010101",
  27131=>"010101111",
  27132=>"111100111",
  27133=>"010001001",
  27134=>"001111110",
  27135=>"101110000",
  27136=>"011011000",
  27137=>"001000011",
  27138=>"110101110",
  27139=>"001001111",
  27140=>"101111011",
  27141=>"000000100",
  27142=>"010110000",
  27143=>"001111110",
  27144=>"100011111",
  27145=>"111111101",
  27146=>"100110110",
  27147=>"101011111",
  27148=>"100110000",
  27149=>"011100101",
  27150=>"000010111",
  27151=>"000101011",
  27152=>"000100001",
  27153=>"100010010",
  27154=>"000001111",
  27155=>"111011110",
  27156=>"110101000",
  27157=>"110000001",
  27158=>"010100010",
  27159=>"001101111",
  27160=>"101000000",
  27161=>"110000001",
  27162=>"110101001",
  27163=>"001011001",
  27164=>"100100011",
  27165=>"001110010",
  27166=>"111101001",
  27167=>"011100001",
  27168=>"000010011",
  27169=>"111110011",
  27170=>"110110110",
  27171=>"110111000",
  27172=>"111100010",
  27173=>"101011111",
  27174=>"100000110",
  27175=>"011111101",
  27176=>"001101111",
  27177=>"000000001",
  27178=>"000011000",
  27179=>"101011110",
  27180=>"001111111",
  27181=>"000100011",
  27182=>"100000110",
  27183=>"111110101",
  27184=>"000001110",
  27185=>"010010001",
  27186=>"011111011",
  27187=>"101110110",
  27188=>"101111000",
  27189=>"010010100",
  27190=>"111001011",
  27191=>"010011011",
  27192=>"111001100",
  27193=>"111100010",
  27194=>"110000110",
  27195=>"111101101",
  27196=>"000101001",
  27197=>"010000000",
  27198=>"010000000",
  27199=>"000001000",
  27200=>"011100100",
  27201=>"101111001",
  27202=>"010100001",
  27203=>"001101111",
  27204=>"000101001",
  27205=>"110100010",
  27206=>"010010101",
  27207=>"001000111",
  27208=>"011110011",
  27209=>"000010111",
  27210=>"010001111",
  27211=>"000111011",
  27212=>"011000110",
  27213=>"100111010",
  27214=>"011010001",
  27215=>"111111000",
  27216=>"100011010",
  27217=>"110100100",
  27218=>"000001011",
  27219=>"100100100",
  27220=>"001101001",
  27221=>"110100001",
  27222=>"111110100",
  27223=>"110100101",
  27224=>"000000011",
  27225=>"111110001",
  27226=>"111110011",
  27227=>"111010001",
  27228=>"010111000",
  27229=>"010100001",
  27230=>"000101101",
  27231=>"111110001",
  27232=>"110010111",
  27233=>"000001101",
  27234=>"101010010",
  27235=>"110011001",
  27236=>"010100011",
  27237=>"100100010",
  27238=>"111101100",
  27239=>"110010111",
  27240=>"110110111",
  27241=>"000101110",
  27242=>"011010100",
  27243=>"000100110",
  27244=>"011100110",
  27245=>"110010101",
  27246=>"011110010",
  27247=>"000010101",
  27248=>"111010011",
  27249=>"111001111",
  27250=>"010101011",
  27251=>"100000101",
  27252=>"111111110",
  27253=>"010000110",
  27254=>"001100010",
  27255=>"000101010",
  27256=>"100010100",
  27257=>"110110111",
  27258=>"101010000",
  27259=>"100001101",
  27260=>"111100101",
  27261=>"000101000",
  27262=>"001001001",
  27263=>"000010110",
  27264=>"011110000",
  27265=>"101010011",
  27266=>"000011111",
  27267=>"100110110",
  27268=>"111011110",
  27269=>"110110101",
  27270=>"111010111",
  27271=>"101110110",
  27272=>"011100110",
  27273=>"000101101",
  27274=>"110010011",
  27275=>"110011100",
  27276=>"101100010",
  27277=>"100000110",
  27278=>"000000100",
  27279=>"010010111",
  27280=>"011111101",
  27281=>"011111101",
  27282=>"111111101",
  27283=>"101110011",
  27284=>"010000111",
  27285=>"100001001",
  27286=>"010001111",
  27287=>"101101101",
  27288=>"010110000",
  27289=>"010011000",
  27290=>"100100000",
  27291=>"101101100",
  27292=>"000110011",
  27293=>"000001110",
  27294=>"010110000",
  27295=>"100000101",
  27296=>"011111101",
  27297=>"100101011",
  27298=>"011001000",
  27299=>"011110111",
  27300=>"000100111",
  27301=>"111000001",
  27302=>"001100010",
  27303=>"001110010",
  27304=>"000001011",
  27305=>"010100111",
  27306=>"110001100",
  27307=>"101000010",
  27308=>"011001111",
  27309=>"011111101",
  27310=>"000000011",
  27311=>"010111101",
  27312=>"011010001",
  27313=>"100110111",
  27314=>"110001111",
  27315=>"011011101",
  27316=>"101110110",
  27317=>"001101010",
  27318=>"000011011",
  27319=>"001101011",
  27320=>"010111010",
  27321=>"001100101",
  27322=>"001000100",
  27323=>"100110010",
  27324=>"011000011",
  27325=>"011001111",
  27326=>"101000101",
  27327=>"000000000",
  27328=>"000110111",
  27329=>"010011100",
  27330=>"100101101",
  27331=>"010111111",
  27332=>"111110010",
  27333=>"000100001",
  27334=>"111000110",
  27335=>"001100011",
  27336=>"100100101",
  27337=>"001111101",
  27338=>"010001001",
  27339=>"010100101",
  27340=>"001110101",
  27341=>"000000110",
  27342=>"011110001",
  27343=>"001101111",
  27344=>"101101010",
  27345=>"000100000",
  27346=>"010011110",
  27347=>"111011011",
  27348=>"100000101",
  27349=>"101101001",
  27350=>"001100011",
  27351=>"011110011",
  27352=>"001001100",
  27353=>"110111111",
  27354=>"011000001",
  27355=>"000001110",
  27356=>"110011101",
  27357=>"100110000",
  27358=>"111001100",
  27359=>"100111001",
  27360=>"100101001",
  27361=>"110000110",
  27362=>"111101001",
  27363=>"001101011",
  27364=>"110000110",
  27365=>"111001000",
  27366=>"000110100",
  27367=>"000000111",
  27368=>"110111110",
  27369=>"001000001",
  27370=>"010000101",
  27371=>"111001100",
  27372=>"000100111",
  27373=>"110100110",
  27374=>"011101111",
  27375=>"111111111",
  27376=>"100001111",
  27377=>"101000100",
  27378=>"011000110",
  27379=>"100100101",
  27380=>"100110100",
  27381=>"110100100",
  27382=>"110010001",
  27383=>"101000011",
  27384=>"111011111",
  27385=>"100000010",
  27386=>"110001001",
  27387=>"001010010",
  27388=>"101110000",
  27389=>"010001110",
  27390=>"101111111",
  27391=>"111011111",
  27392=>"011100101",
  27393=>"101111110",
  27394=>"000000101",
  27395=>"101111000",
  27396=>"111000100",
  27397=>"101110010",
  27398=>"011001110",
  27399=>"010100001",
  27400=>"100110110",
  27401=>"100001101",
  27402=>"100010001",
  27403=>"010111100",
  27404=>"000000001",
  27405=>"110100101",
  27406=>"010110111",
  27407=>"010010101",
  27408=>"110111100",
  27409=>"101101111",
  27410=>"110110100",
  27411=>"010110001",
  27412=>"111111010",
  27413=>"010111000",
  27414=>"000001100",
  27415=>"101101000",
  27416=>"111101001",
  27417=>"001110011",
  27418=>"101100100",
  27419=>"010101000",
  27420=>"010111100",
  27421=>"100001110",
  27422=>"000011110",
  27423=>"111101111",
  27424=>"010000111",
  27425=>"110101100",
  27426=>"101011111",
  27427=>"001000001",
  27428=>"101010100",
  27429=>"001110100",
  27430=>"110111010",
  27431=>"000011000",
  27432=>"000010000",
  27433=>"100001010",
  27434=>"011001111",
  27435=>"010010110",
  27436=>"111111110",
  27437=>"001000001",
  27438=>"101110011",
  27439=>"101101011",
  27440=>"010001110",
  27441=>"011010111",
  27442=>"101010001",
  27443=>"100010111",
  27444=>"011001000",
  27445=>"010010100",
  27446=>"000001100",
  27447=>"000110100",
  27448=>"000110110",
  27449=>"000001111",
  27450=>"110011110",
  27451=>"000011000",
  27452=>"001000111",
  27453=>"011010110",
  27454=>"010000101",
  27455=>"101000011",
  27456=>"100010111",
  27457=>"001011100",
  27458=>"001100101",
  27459=>"000101010",
  27460=>"000101010",
  27461=>"110010110",
  27462=>"101001101",
  27463=>"101001101",
  27464=>"000111110",
  27465=>"011000111",
  27466=>"111001110",
  27467=>"000100010",
  27468=>"110111100",
  27469=>"011100111",
  27470=>"000010111",
  27471=>"110010001",
  27472=>"000000000",
  27473=>"010101110",
  27474=>"010110011",
  27475=>"010000001",
  27476=>"010110111",
  27477=>"110011010",
  27478=>"111111110",
  27479=>"000100011",
  27480=>"011110010",
  27481=>"011100010",
  27482=>"010010111",
  27483=>"011001010",
  27484=>"001111010",
  27485=>"100001111",
  27486=>"000010101",
  27487=>"101111001",
  27488=>"111000010",
  27489=>"000000100",
  27490=>"101001101",
  27491=>"001101110",
  27492=>"100000010",
  27493=>"111101010",
  27494=>"000001000",
  27495=>"100111000",
  27496=>"011000000",
  27497=>"110111001",
  27498=>"110100001",
  27499=>"010010111",
  27500=>"100000011",
  27501=>"101111111",
  27502=>"100111110",
  27503=>"101100100",
  27504=>"110100100",
  27505=>"010110011",
  27506=>"111011110",
  27507=>"111010001",
  27508=>"110100111",
  27509=>"001000111",
  27510=>"011001000",
  27511=>"111101010",
  27512=>"111111111",
  27513=>"010111110",
  27514=>"011010001",
  27515=>"100101010",
  27516=>"010111011",
  27517=>"100000101",
  27518=>"010000110",
  27519=>"110000011",
  27520=>"111111111",
  27521=>"010101000",
  27522=>"110101011",
  27523=>"101000101",
  27524=>"001010100",
  27525=>"111101100",
  27526=>"111100000",
  27527=>"101110001",
  27528=>"000111010",
  27529=>"101000000",
  27530=>"011000000",
  27531=>"011111010",
  27532=>"011010100",
  27533=>"001001011",
  27534=>"111010110",
  27535=>"101001111",
  27536=>"011101110",
  27537=>"100011111",
  27538=>"000001111",
  27539=>"000110000",
  27540=>"001101101",
  27541=>"101000000",
  27542=>"001101001",
  27543=>"001111011",
  27544=>"000000011",
  27545=>"001000001",
  27546=>"111110001",
  27547=>"010010011",
  27548=>"010000000",
  27549=>"011100101",
  27550=>"000001011",
  27551=>"111100101",
  27552=>"010110100",
  27553=>"010101000",
  27554=>"101101010",
  27555=>"111011111",
  27556=>"000100000",
  27557=>"010110100",
  27558=>"101110011",
  27559=>"100000101",
  27560=>"100001111",
  27561=>"110101000",
  27562=>"101111011",
  27563=>"100010101",
  27564=>"001111010",
  27565=>"100100111",
  27566=>"101010011",
  27567=>"011100100",
  27568=>"111100101",
  27569=>"110100101",
  27570=>"100101001",
  27571=>"111100101",
  27572=>"111000000",
  27573=>"001111010",
  27574=>"101101100",
  27575=>"011110010",
  27576=>"111111001",
  27577=>"000101001",
  27578=>"011010111",
  27579=>"000000110",
  27580=>"000101111",
  27581=>"001101010",
  27582=>"000111111",
  27583=>"011001000",
  27584=>"011111000",
  27585=>"001110101",
  27586=>"101100010",
  27587=>"000000011",
  27588=>"100101101",
  27589=>"101011100",
  27590=>"001100011",
  27591=>"011000101",
  27592=>"011001000",
  27593=>"001000010",
  27594=>"010101110",
  27595=>"001000001",
  27596=>"001101010",
  27597=>"011001000",
  27598=>"111001100",
  27599=>"010010101",
  27600=>"111100101",
  27601=>"101101110",
  27602=>"011110100",
  27603=>"010011110",
  27604=>"100010001",
  27605=>"110101010",
  27606=>"000100100",
  27607=>"101100100",
  27608=>"101011001",
  27609=>"001110101",
  27610=>"001100110",
  27611=>"010001100",
  27612=>"000101110",
  27613=>"001000000",
  27614=>"000000111",
  27615=>"110000011",
  27616=>"111010000",
  27617=>"101111110",
  27618=>"010101001",
  27619=>"111011101",
  27620=>"000011000",
  27621=>"101101001",
  27622=>"101110011",
  27623=>"010001000",
  27624=>"111111110",
  27625=>"000001001",
  27626=>"110011100",
  27627=>"000000111",
  27628=>"010111110",
  27629=>"100011011",
  27630=>"001100111",
  27631=>"011001110",
  27632=>"010001101",
  27633=>"010100111",
  27634=>"110011000",
  27635=>"111100000",
  27636=>"101100101",
  27637=>"100101111",
  27638=>"110101100",
  27639=>"011000000",
  27640=>"111110100",
  27641=>"101000000",
  27642=>"111110111",
  27643=>"111011010",
  27644=>"001011111",
  27645=>"110110000",
  27646=>"110000101",
  27647=>"011111011",
  27648=>"010010101",
  27649=>"101110111",
  27650=>"010101000",
  27651=>"100100101",
  27652=>"011101011",
  27653=>"111110111",
  27654=>"111010011",
  27655=>"110011000",
  27656=>"010100111",
  27657=>"111001101",
  27658=>"111000011",
  27659=>"010111010",
  27660=>"011001001",
  27661=>"100010000",
  27662=>"110111111",
  27663=>"000110001",
  27664=>"011010011",
  27665=>"010101111",
  27666=>"101110000",
  27667=>"111010011",
  27668=>"001011001",
  27669=>"100001001",
  27670=>"110001001",
  27671=>"001010011",
  27672=>"111010100",
  27673=>"111110111",
  27674=>"001010011",
  27675=>"000110110",
  27676=>"111001110",
  27677=>"101001010",
  27678=>"010010100",
  27679=>"011000011",
  27680=>"111101010",
  27681=>"011101000",
  27682=>"011011000",
  27683=>"000111000",
  27684=>"011001011",
  27685=>"101011111",
  27686=>"100001000",
  27687=>"111111101",
  27688=>"011101000",
  27689=>"000110111",
  27690=>"000111111",
  27691=>"110011111",
  27692=>"100101101",
  27693=>"000010010",
  27694=>"011000100",
  27695=>"000010011",
  27696=>"111000101",
  27697=>"110001000",
  27698=>"010101101",
  27699=>"110001001",
  27700=>"100011101",
  27701=>"110110100",
  27702=>"010110001",
  27703=>"110100010",
  27704=>"110111000",
  27705=>"001100000",
  27706=>"001000100",
  27707=>"101000010",
  27708=>"011100010",
  27709=>"100011101",
  27710=>"011111111",
  27711=>"111101111",
  27712=>"111111010",
  27713=>"111010010",
  27714=>"100100000",
  27715=>"111101000",
  27716=>"100101111",
  27717=>"001111111",
  27718=>"111111001",
  27719=>"101010011",
  27720=>"000001000",
  27721=>"111001000",
  27722=>"101001011",
  27723=>"111100001",
  27724=>"111010001",
  27725=>"101010101",
  27726=>"100110111",
  27727=>"111110100",
  27728=>"000100110",
  27729=>"000100000",
  27730=>"111011001",
  27731=>"011010111",
  27732=>"010111011",
  27733=>"011010010",
  27734=>"000100110",
  27735=>"010001010",
  27736=>"111001010",
  27737=>"010110011",
  27738=>"101010000",
  27739=>"100001100",
  27740=>"001110011",
  27741=>"011111010",
  27742=>"010111100",
  27743=>"110101000",
  27744=>"000000101",
  27745=>"011100100",
  27746=>"000001101",
  27747=>"000000011",
  27748=>"010101110",
  27749=>"001011111",
  27750=>"010000011",
  27751=>"111110110",
  27752=>"110010100",
  27753=>"000001010",
  27754=>"011100000",
  27755=>"100010100",
  27756=>"011001010",
  27757=>"001001000",
  27758=>"110010010",
  27759=>"101111010",
  27760=>"111000111",
  27761=>"111100010",
  27762=>"101010111",
  27763=>"000110010",
  27764=>"110001011",
  27765=>"111001111",
  27766=>"010000110",
  27767=>"000100110",
  27768=>"010011110",
  27769=>"110001101",
  27770=>"111110000",
  27771=>"101101110",
  27772=>"011111101",
  27773=>"101110000",
  27774=>"011111011",
  27775=>"000110011",
  27776=>"110100111",
  27777=>"110011101",
  27778=>"100011001",
  27779=>"001001001",
  27780=>"000001111",
  27781=>"110111110",
  27782=>"110101000",
  27783=>"000111000",
  27784=>"000001010",
  27785=>"100100000",
  27786=>"001001111",
  27787=>"010111100",
  27788=>"100111010",
  27789=>"010101010",
  27790=>"011100110",
  27791=>"010100110",
  27792=>"101111101",
  27793=>"111110011",
  27794=>"100001000",
  27795=>"010111111",
  27796=>"011000100",
  27797=>"011111010",
  27798=>"000000011",
  27799=>"101111011",
  27800=>"100100101",
  27801=>"101000011",
  27802=>"101110000",
  27803=>"001000100",
  27804=>"011111111",
  27805=>"100111010",
  27806=>"010101111",
  27807=>"111011110",
  27808=>"100000111",
  27809=>"010000000",
  27810=>"110010001",
  27811=>"100111001",
  27812=>"110010101",
  27813=>"111101111",
  27814=>"111101000",
  27815=>"101101111",
  27816=>"001100100",
  27817=>"000101010",
  27818=>"000010000",
  27819=>"011100100",
  27820=>"110000000",
  27821=>"110111001",
  27822=>"001101101",
  27823=>"101001001",
  27824=>"100001000",
  27825=>"000111001",
  27826=>"001011001",
  27827=>"110100101",
  27828=>"010111110",
  27829=>"101101111",
  27830=>"011010010",
  27831=>"101111111",
  27832=>"110101101",
  27833=>"111000100",
  27834=>"011101111",
  27835=>"000111011",
  27836=>"110101011",
  27837=>"000111001",
  27838=>"101001101",
  27839=>"000001010",
  27840=>"001011110",
  27841=>"001101000",
  27842=>"100001110",
  27843=>"000100110",
  27844=>"000100001",
  27845=>"011001110",
  27846=>"111011010",
  27847=>"101011000",
  27848=>"010000011",
  27849=>"011111010",
  27850=>"100111010",
  27851=>"011110000",
  27852=>"010101010",
  27853=>"110100011",
  27854=>"101011101",
  27855=>"100001001",
  27856=>"000000000",
  27857=>"100101000",
  27858=>"010110101",
  27859=>"111111101",
  27860=>"100001111",
  27861=>"010110011",
  27862=>"110011010",
  27863=>"101110000",
  27864=>"100000100",
  27865=>"000011010",
  27866=>"110000000",
  27867=>"001001111",
  27868=>"010110110",
  27869=>"001001100",
  27870=>"101001001",
  27871=>"000010000",
  27872=>"110110010",
  27873=>"111111110",
  27874=>"101100010",
  27875=>"010110001",
  27876=>"010100110",
  27877=>"010000011",
  27878=>"000110110",
  27879=>"101011001",
  27880=>"010111010",
  27881=>"000000110",
  27882=>"111111011",
  27883=>"110011000",
  27884=>"111001010",
  27885=>"110011111",
  27886=>"011001011",
  27887=>"000100000",
  27888=>"111000000",
  27889=>"101100111",
  27890=>"101001101",
  27891=>"101100111",
  27892=>"010000001",
  27893=>"110100011",
  27894=>"101110110",
  27895=>"011110101",
  27896=>"001101001",
  27897=>"000001001",
  27898=>"111110000",
  27899=>"000000000",
  27900=>"100011000",
  27901=>"000111101",
  27902=>"111000011",
  27903=>"110011100",
  27904=>"000000000",
  27905=>"011010010",
  27906=>"011011110",
  27907=>"000111111",
  27908=>"010101000",
  27909=>"000100011",
  27910=>"000001111",
  27911=>"110101111",
  27912=>"110001111",
  27913=>"000110001",
  27914=>"001111101",
  27915=>"101111111",
  27916=>"010101110",
  27917=>"001001110",
  27918=>"111010111",
  27919=>"011111101",
  27920=>"001100000",
  27921=>"010100001",
  27922=>"000001010",
  27923=>"101111110",
  27924=>"111010000",
  27925=>"111111011",
  27926=>"010111001",
  27927=>"000110110",
  27928=>"001001101",
  27929=>"101011010",
  27930=>"001101011",
  27931=>"110110110",
  27932=>"001010110",
  27933=>"010110010",
  27934=>"011100001",
  27935=>"011110100",
  27936=>"001000001",
  27937=>"111101110",
  27938=>"011000100",
  27939=>"110100011",
  27940=>"000011011",
  27941=>"111011011",
  27942=>"111001001",
  27943=>"110000010",
  27944=>"011010010",
  27945=>"101101100",
  27946=>"100100010",
  27947=>"101111000",
  27948=>"101100000",
  27949=>"010011101",
  27950=>"000100100",
  27951=>"010001001",
  27952=>"000001111",
  27953=>"001100111",
  27954=>"001101011",
  27955=>"000110100",
  27956=>"001000100",
  27957=>"001111101",
  27958=>"000111100",
  27959=>"101010111",
  27960=>"111110100",
  27961=>"001100101",
  27962=>"111010111",
  27963=>"111000000",
  27964=>"101001000",
  27965=>"000010010",
  27966=>"110111100",
  27967=>"000010101",
  27968=>"100000100",
  27969=>"010011110",
  27970=>"001100101",
  27971=>"001010000",
  27972=>"111111001",
  27973=>"110100101",
  27974=>"011000000",
  27975=>"010111101",
  27976=>"110010110",
  27977=>"000100001",
  27978=>"111111100",
  27979=>"101111101",
  27980=>"111011011",
  27981=>"011100100",
  27982=>"011111000",
  27983=>"001000000",
  27984=>"100010110",
  27985=>"000010100",
  27986=>"000101001",
  27987=>"111100000",
  27988=>"001100111",
  27989=>"110000001",
  27990=>"100100001",
  27991=>"011110010",
  27992=>"110001100",
  27993=>"010111100",
  27994=>"110001011",
  27995=>"001110100",
  27996=>"101111111",
  27997=>"110101000",
  27998=>"001100100",
  27999=>"111111011",
  28000=>"000101100",
  28001=>"100101110",
  28002=>"110100111",
  28003=>"011010010",
  28004=>"111111110",
  28005=>"001110011",
  28006=>"001111110",
  28007=>"100010110",
  28008=>"011001001",
  28009=>"111001111",
  28010=>"001100111",
  28011=>"001110001",
  28012=>"000000011",
  28013=>"001000000",
  28014=>"101000111",
  28015=>"000010110",
  28016=>"011000110",
  28017=>"100010011",
  28018=>"010001101",
  28019=>"011001001",
  28020=>"100111001",
  28021=>"100011110",
  28022=>"100001010",
  28023=>"000000110",
  28024=>"000000011",
  28025=>"111101100",
  28026=>"110101101",
  28027=>"011101010",
  28028=>"110101010",
  28029=>"101110111",
  28030=>"011001110",
  28031=>"111110000",
  28032=>"000000110",
  28033=>"001110001",
  28034=>"011000000",
  28035=>"100100111",
  28036=>"001100110",
  28037=>"000100010",
  28038=>"001000000",
  28039=>"001010101",
  28040=>"001011110",
  28041=>"000100000",
  28042=>"111101101",
  28043=>"101111110",
  28044=>"001101011",
  28045=>"101110011",
  28046=>"111001000",
  28047=>"110110011",
  28048=>"010101000",
  28049=>"010111111",
  28050=>"000111110",
  28051=>"100100011",
  28052=>"000111101",
  28053=>"101001101",
  28054=>"010111111",
  28055=>"000101110",
  28056=>"000001101",
  28057=>"111000110",
  28058=>"011011111",
  28059=>"001000111",
  28060=>"101000100",
  28061=>"001010111",
  28062=>"111100000",
  28063=>"111000010",
  28064=>"100001111",
  28065=>"111110000",
  28066=>"011111000",
  28067=>"001110101",
  28068=>"111000001",
  28069=>"001111000",
  28070=>"000111111",
  28071=>"111110001",
  28072=>"001010010",
  28073=>"101011110",
  28074=>"000000111",
  28075=>"010100100",
  28076=>"111000110",
  28077=>"101010010",
  28078=>"110011110",
  28079=>"101001010",
  28080=>"101100101",
  28081=>"101010000",
  28082=>"011110111",
  28083=>"110111111",
  28084=>"101111111",
  28085=>"100001010",
  28086=>"000010011",
  28087=>"100000110",
  28088=>"100000000",
  28089=>"000010010",
  28090=>"101100100",
  28091=>"010001011",
  28092=>"110000000",
  28093=>"010011001",
  28094=>"000101111",
  28095=>"010000000",
  28096=>"111101110",
  28097=>"010011000",
  28098=>"101101000",
  28099=>"111011111",
  28100=>"000010111",
  28101=>"001010000",
  28102=>"111100111",
  28103=>"111110110",
  28104=>"110100110",
  28105=>"111111110",
  28106=>"001010001",
  28107=>"101000001",
  28108=>"111101100",
  28109=>"011001111",
  28110=>"000110000",
  28111=>"101110010",
  28112=>"101100010",
  28113=>"110010111",
  28114=>"111010100",
  28115=>"010110001",
  28116=>"011100110",
  28117=>"101111101",
  28118=>"111000000",
  28119=>"111101010",
  28120=>"101001011",
  28121=>"111111011",
  28122=>"000010111",
  28123=>"010011111",
  28124=>"111110100",
  28125=>"011011111",
  28126=>"000110111",
  28127=>"110110100",
  28128=>"001010011",
  28129=>"010100011",
  28130=>"010110100",
  28131=>"111001100",
  28132=>"100101000",
  28133=>"010111010",
  28134=>"101101001",
  28135=>"010011000",
  28136=>"011000000",
  28137=>"011100100",
  28138=>"010010010",
  28139=>"101001101",
  28140=>"001000001",
  28141=>"000000011",
  28142=>"101100000",
  28143=>"000101000",
  28144=>"011011010",
  28145=>"110100001",
  28146=>"011111001",
  28147=>"110001001",
  28148=>"010101110",
  28149=>"000111000",
  28150=>"001001011",
  28151=>"000011101",
  28152=>"101111000",
  28153=>"111101000",
  28154=>"011011000",
  28155=>"110100001",
  28156=>"001111001",
  28157=>"010011001",
  28158=>"011011010",
  28159=>"100110000",
  28160=>"010010001",
  28161=>"010011111",
  28162=>"100101110",
  28163=>"101010110",
  28164=>"110100101",
  28165=>"101111110",
  28166=>"101100001",
  28167=>"100110001",
  28168=>"000010110",
  28169=>"100110110",
  28170=>"101101001",
  28171=>"110100010",
  28172=>"101111010",
  28173=>"001000000",
  28174=>"001111001",
  28175=>"110101011",
  28176=>"100111110",
  28177=>"110001011",
  28178=>"101111101",
  28179=>"001001010",
  28180=>"010000010",
  28181=>"010100110",
  28182=>"000001101",
  28183=>"100001010",
  28184=>"000110011",
  28185=>"101110110",
  28186=>"110011110",
  28187=>"100010010",
  28188=>"111111000",
  28189=>"010100011",
  28190=>"101001001",
  28191=>"101101010",
  28192=>"010000111",
  28193=>"100111000",
  28194=>"010100001",
  28195=>"000100100",
  28196=>"010110110",
  28197=>"110010000",
  28198=>"111000100",
  28199=>"101001011",
  28200=>"010100011",
  28201=>"011010101",
  28202=>"110111011",
  28203=>"101010101",
  28204=>"111111000",
  28205=>"000010100",
  28206=>"000101110",
  28207=>"101111010",
  28208=>"110001111",
  28209=>"111000110",
  28210=>"011000001",
  28211=>"111110011",
  28212=>"111101011",
  28213=>"001110111",
  28214=>"111111000",
  28215=>"110001101",
  28216=>"100111010",
  28217=>"000100101",
  28218=>"010101110",
  28219=>"000001010",
  28220=>"101011110",
  28221=>"001010101",
  28222=>"000101001",
  28223=>"111011100",
  28224=>"111011100",
  28225=>"100011100",
  28226=>"001001111",
  28227=>"100101011",
  28228=>"011111000",
  28229=>"011000100",
  28230=>"001110011",
  28231=>"001001001",
  28232=>"001110011",
  28233=>"111101101",
  28234=>"100111111",
  28235=>"011100101",
  28236=>"011110101",
  28237=>"011010011",
  28238=>"111110011",
  28239=>"001001110",
  28240=>"101111111",
  28241=>"000011001",
  28242=>"100111111",
  28243=>"001100010",
  28244=>"100001000",
  28245=>"011110001",
  28246=>"010101110",
  28247=>"111101110",
  28248=>"001001101",
  28249=>"101111011",
  28250=>"110100111",
  28251=>"110110111",
  28252=>"010111100",
  28253=>"011101011",
  28254=>"011101010",
  28255=>"111111101",
  28256=>"000100001",
  28257=>"101110100",
  28258=>"010001000",
  28259=>"111000011",
  28260=>"000100010",
  28261=>"101110011",
  28262=>"101111101",
  28263=>"111111110",
  28264=>"000011111",
  28265=>"011111101",
  28266=>"001001111",
  28267=>"101101111",
  28268=>"110011110",
  28269=>"101010000",
  28270=>"100010011",
  28271=>"010101011",
  28272=>"011000001",
  28273=>"000000010",
  28274=>"111111111",
  28275=>"111010000",
  28276=>"011011010",
  28277=>"110010001",
  28278=>"000001011",
  28279=>"010011101",
  28280=>"101011001",
  28281=>"000111011",
  28282=>"111100110",
  28283=>"110110110",
  28284=>"110010000",
  28285=>"011010001",
  28286=>"101111101",
  28287=>"101011001",
  28288=>"100010010",
  28289=>"000011100",
  28290=>"111111110",
  28291=>"000010100",
  28292=>"101100001",
  28293=>"000110011",
  28294=>"001110100",
  28295=>"000010010",
  28296=>"001001010",
  28297=>"011010010",
  28298=>"010011010",
  28299=>"110100100",
  28300=>"000000010",
  28301=>"101110111",
  28302=>"101011011",
  28303=>"111111000",
  28304=>"010000111",
  28305=>"111101001",
  28306=>"110101101",
  28307=>"001000011",
  28308=>"010011000",
  28309=>"000100000",
  28310=>"001110011",
  28311=>"101010100",
  28312=>"110110010",
  28313=>"011110011",
  28314=>"000001100",
  28315=>"001011000",
  28316=>"000110110",
  28317=>"011001101",
  28318=>"111101100",
  28319=>"011100100",
  28320=>"000010101",
  28321=>"110000000",
  28322=>"111011111",
  28323=>"001000111",
  28324=>"000101100",
  28325=>"111111101",
  28326=>"011100000",
  28327=>"000000000",
  28328=>"011101011",
  28329=>"111111101",
  28330=>"110100110",
  28331=>"010100101",
  28332=>"100001001",
  28333=>"100011001",
  28334=>"000110001",
  28335=>"100111000",
  28336=>"010110100",
  28337=>"111001101",
  28338=>"001001001",
  28339=>"100100000",
  28340=>"111101011",
  28341=>"001011010",
  28342=>"000100110",
  28343=>"000101011",
  28344=>"100001010",
  28345=>"110010110",
  28346=>"111111110",
  28347=>"010110011",
  28348=>"110011111",
  28349=>"001100001",
  28350=>"100110101",
  28351=>"001100110",
  28352=>"100010101",
  28353=>"111111101",
  28354=>"110101110",
  28355=>"100000000",
  28356=>"011011111",
  28357=>"111101101",
  28358=>"100101011",
  28359=>"100010010",
  28360=>"101101101",
  28361=>"101111011",
  28362=>"110111110",
  28363=>"011110100",
  28364=>"011001010",
  28365=>"110011111",
  28366=>"000111011",
  28367=>"101011100",
  28368=>"011101111",
  28369=>"100100010",
  28370=>"101110001",
  28371=>"110111110",
  28372=>"101011010",
  28373=>"111110110",
  28374=>"110111111",
  28375=>"100011010",
  28376=>"100010111",
  28377=>"010001010",
  28378=>"001100011",
  28379=>"111011111",
  28380=>"111110111",
  28381=>"101101101",
  28382=>"100001010",
  28383=>"000001010",
  28384=>"110100101",
  28385=>"011111110",
  28386=>"101010011",
  28387=>"100010111",
  28388=>"101000010",
  28389=>"110000001",
  28390=>"010010100",
  28391=>"010100100",
  28392=>"001010000",
  28393=>"100011111",
  28394=>"011010010",
  28395=>"100000100",
  28396=>"110000000",
  28397=>"001000100",
  28398=>"011001001",
  28399=>"101111101",
  28400=>"010010010",
  28401=>"111100001",
  28402=>"000010000",
  28403=>"100100010",
  28404=>"011001000",
  28405=>"111001101",
  28406=>"101001110",
  28407=>"101100110",
  28408=>"100100010",
  28409=>"000001100",
  28410=>"110110000",
  28411=>"100011101",
  28412=>"010111011",
  28413=>"011011000",
  28414=>"011111110",
  28415=>"111010111",
  28416=>"011111110",
  28417=>"111010000",
  28418=>"101010000",
  28419=>"101100000",
  28420=>"011001001",
  28421=>"110111101",
  28422=>"000010001",
  28423=>"010110001",
  28424=>"000100010",
  28425=>"110000010",
  28426=>"110100111",
  28427=>"000000000",
  28428=>"100101111",
  28429=>"001110011",
  28430=>"000010011",
  28431=>"001110000",
  28432=>"100110010",
  28433=>"111001101",
  28434=>"011101100",
  28435=>"001111100",
  28436=>"010000100",
  28437=>"100110000",
  28438=>"110010101",
  28439=>"100001001",
  28440=>"010000000",
  28441=>"000001000",
  28442=>"101100100",
  28443=>"111111001",
  28444=>"001100100",
  28445=>"011100111",
  28446=>"101011000",
  28447=>"000001111",
  28448=>"111100100",
  28449=>"101010001",
  28450=>"100000011",
  28451=>"000000101",
  28452=>"001100000",
  28453=>"101110110",
  28454=>"011001100",
  28455=>"010111011",
  28456=>"100001010",
  28457=>"111101000",
  28458=>"101101110",
  28459=>"011010110",
  28460=>"011110001",
  28461=>"100010100",
  28462=>"111011110",
  28463=>"001111001",
  28464=>"001001001",
  28465=>"000101101",
  28466=>"000101000",
  28467=>"101011010",
  28468=>"011101011",
  28469=>"111010110",
  28470=>"110110100",
  28471=>"000111000",
  28472=>"000101111",
  28473=>"100000100",
  28474=>"010001000",
  28475=>"101100101",
  28476=>"100000100",
  28477=>"101011010",
  28478=>"000011110",
  28479=>"110000111",
  28480=>"011110010",
  28481=>"000001000",
  28482=>"110110000",
  28483=>"000000010",
  28484=>"001100001",
  28485=>"100110110",
  28486=>"100000111",
  28487=>"111001001",
  28488=>"100001010",
  28489=>"101101011",
  28490=>"110000111",
  28491=>"111101101",
  28492=>"011010111",
  28493=>"110011011",
  28494=>"010010100",
  28495=>"101111001",
  28496=>"010100111",
  28497=>"011100001",
  28498=>"111001000",
  28499=>"100111111",
  28500=>"001000110",
  28501=>"000110111",
  28502=>"011000001",
  28503=>"100100001",
  28504=>"000000101",
  28505=>"101111100",
  28506=>"101101011",
  28507=>"010100000",
  28508=>"101100010",
  28509=>"111001100",
  28510=>"001111011",
  28511=>"000110000",
  28512=>"010111010",
  28513=>"110001011",
  28514=>"100110001",
  28515=>"110111010",
  28516=>"110111001",
  28517=>"101011011",
  28518=>"001001001",
  28519=>"011111000",
  28520=>"001001100",
  28521=>"100000101",
  28522=>"111100010",
  28523=>"101000110",
  28524=>"110101111",
  28525=>"110100011",
  28526=>"010111010",
  28527=>"110100111",
  28528=>"100001001",
  28529=>"011100010",
  28530=>"100111101",
  28531=>"111110110",
  28532=>"111101001",
  28533=>"100111000",
  28534=>"100000011",
  28535=>"000000111",
  28536=>"101101000",
  28537=>"001010000",
  28538=>"101110000",
  28539=>"100000000",
  28540=>"000100100",
  28541=>"101010110",
  28542=>"010111011",
  28543=>"001100011",
  28544=>"011010011",
  28545=>"000110110",
  28546=>"001010010",
  28547=>"000001111",
  28548=>"110101011",
  28549=>"101110110",
  28550=>"110001001",
  28551=>"100111011",
  28552=>"101001000",
  28553=>"001111111",
  28554=>"001111101",
  28555=>"001100110",
  28556=>"001011011",
  28557=>"000100100",
  28558=>"101101000",
  28559=>"011111000",
  28560=>"111010111",
  28561=>"001011100",
  28562=>"110001011",
  28563=>"100001001",
  28564=>"010100111",
  28565=>"011101111",
  28566=>"110111101",
  28567=>"001101011",
  28568=>"000101001",
  28569=>"000000110",
  28570=>"110100100",
  28571=>"101110101",
  28572=>"011000010",
  28573=>"010011010",
  28574=>"110000010",
  28575=>"010100110",
  28576=>"110011011",
  28577=>"001011110",
  28578=>"010101111",
  28579=>"110001011",
  28580=>"000000010",
  28581=>"111110110",
  28582=>"010000111",
  28583=>"100010111",
  28584=>"101110001",
  28585=>"010000100",
  28586=>"110111110",
  28587=>"000110111",
  28588=>"110010100",
  28589=>"000100110",
  28590=>"001010110",
  28591=>"101110000",
  28592=>"001100110",
  28593=>"111000011",
  28594=>"000011010",
  28595=>"111111100",
  28596=>"110110100",
  28597=>"101111000",
  28598=>"100011011",
  28599=>"000000110",
  28600=>"111101001",
  28601=>"100001111",
  28602=>"111010000",
  28603=>"110101100",
  28604=>"000101010",
  28605=>"101011101",
  28606=>"100000010",
  28607=>"111010000",
  28608=>"010100000",
  28609=>"000100100",
  28610=>"110100001",
  28611=>"000101100",
  28612=>"010010111",
  28613=>"101000101",
  28614=>"100110111",
  28615=>"111110100",
  28616=>"101111101",
  28617=>"110010001",
  28618=>"101110001",
  28619=>"000100100",
  28620=>"100010000",
  28621=>"011001110",
  28622=>"111111111",
  28623=>"101000010",
  28624=>"111100101",
  28625=>"001100001",
  28626=>"101110111",
  28627=>"000100101",
  28628=>"011101010",
  28629=>"110110110",
  28630=>"100001001",
  28631=>"111010100",
  28632=>"110010011",
  28633=>"111111010",
  28634=>"101000010",
  28635=>"100000000",
  28636=>"110101100",
  28637=>"110111100",
  28638=>"111100001",
  28639=>"111000100",
  28640=>"101000111",
  28641=>"000101111",
  28642=>"100000111",
  28643=>"011111110",
  28644=>"001110100",
  28645=>"110101001",
  28646=>"101010111",
  28647=>"000111001",
  28648=>"001110001",
  28649=>"100010010",
  28650=>"001010110",
  28651=>"000010111",
  28652=>"110001000",
  28653=>"100111010",
  28654=>"111111000",
  28655=>"000100101",
  28656=>"111111111",
  28657=>"000111101",
  28658=>"111110100",
  28659=>"101111000",
  28660=>"000110110",
  28661=>"111100111",
  28662=>"100001001",
  28663=>"100000001",
  28664=>"000110001",
  28665=>"101100001",
  28666=>"111110101",
  28667=>"110100001",
  28668=>"100000000",
  28669=>"011101100",
  28670=>"111110111",
  28671=>"111110000",
  28672=>"101010001",
  28673=>"100010110",
  28674=>"101011000",
  28675=>"010000000",
  28676=>"110111110",
  28677=>"000001111",
  28678=>"011011101",
  28679=>"100111010",
  28680=>"110011011",
  28681=>"010111101",
  28682=>"000011100",
  28683=>"000011001",
  28684=>"101110001",
  28685=>"000100001",
  28686=>"111010010",
  28687=>"110111011",
  28688=>"110111111",
  28689=>"010010111",
  28690=>"000010000",
  28691=>"111001110",
  28692=>"001111010",
  28693=>"010110010",
  28694=>"101110100",
  28695=>"111011000",
  28696=>"110010010",
  28697=>"010010100",
  28698=>"100000111",
  28699=>"011111010",
  28700=>"010010001",
  28701=>"101000101",
  28702=>"111101001",
  28703=>"100000111",
  28704=>"100010110",
  28705=>"001001111",
  28706=>"001000110",
  28707=>"100110110",
  28708=>"011101001",
  28709=>"100101100",
  28710=>"101011001",
  28711=>"010010000",
  28712=>"111111010",
  28713=>"101011110",
  28714=>"111000110",
  28715=>"001100011",
  28716=>"010010000",
  28717=>"111011101",
  28718=>"101100100",
  28719=>"110100010",
  28720=>"000100101",
  28721=>"110110011",
  28722=>"101110010",
  28723=>"001011111",
  28724=>"000111001",
  28725=>"000110010",
  28726=>"111100111",
  28727=>"000000000",
  28728=>"010111110",
  28729=>"011010001",
  28730=>"100011001",
  28731=>"111111000",
  28732=>"110110001",
  28733=>"010101011",
  28734=>"001110110",
  28735=>"011110001",
  28736=>"010001100",
  28737=>"010010000",
  28738=>"011001011",
  28739=>"010101001",
  28740=>"011000101",
  28741=>"101011001",
  28742=>"011111111",
  28743=>"110111011",
  28744=>"100000011",
  28745=>"011110110",
  28746=>"001100011",
  28747=>"101110101",
  28748=>"011110110",
  28749=>"100001001",
  28750=>"001111010",
  28751=>"110111010",
  28752=>"100100110",
  28753=>"000010110",
  28754=>"100001111",
  28755=>"010100101",
  28756=>"100011101",
  28757=>"000010010",
  28758=>"000110101",
  28759=>"000000010",
  28760=>"001001101",
  28761=>"101101000",
  28762=>"000011011",
  28763=>"110100111",
  28764=>"001110010",
  28765=>"011000101",
  28766=>"011100000",
  28767=>"010010110",
  28768=>"010110011",
  28769=>"100000100",
  28770=>"001001111",
  28771=>"011010110",
  28772=>"001110010",
  28773=>"010111100",
  28774=>"011010001",
  28775=>"111111111",
  28776=>"001110011",
  28777=>"100010110",
  28778=>"100111001",
  28779=>"010111010",
  28780=>"111110011",
  28781=>"011011101",
  28782=>"101010010",
  28783=>"100000111",
  28784=>"011110110",
  28785=>"010000110",
  28786=>"011110110",
  28787=>"110111110",
  28788=>"001111001",
  28789=>"001000000",
  28790=>"110111111",
  28791=>"101110100",
  28792=>"000010101",
  28793=>"011001000",
  28794=>"010011100",
  28795=>"010001000",
  28796=>"000101100",
  28797=>"000010011",
  28798=>"101001010",
  28799=>"000100101",
  28800=>"111010100",
  28801=>"110111111",
  28802=>"100100000",
  28803=>"110011011",
  28804=>"110100001",
  28805=>"111001110",
  28806=>"001010111",
  28807=>"101010111",
  28808=>"111111011",
  28809=>"001101111",
  28810=>"101111100",
  28811=>"111100101",
  28812=>"000001010",
  28813=>"000110010",
  28814=>"100000101",
  28815=>"011000111",
  28816=>"100100100",
  28817=>"010100101",
  28818=>"101011000",
  28819=>"011101000",
  28820=>"101101100",
  28821=>"001110000",
  28822=>"000010110",
  28823=>"111001111",
  28824=>"010101010",
  28825=>"101101111",
  28826=>"101000111",
  28827=>"100010100",
  28828=>"010100011",
  28829=>"010010101",
  28830=>"100011000",
  28831=>"111111110",
  28832=>"010101101",
  28833=>"010010111",
  28834=>"001110010",
  28835=>"011011011",
  28836=>"111011000",
  28837=>"000010010",
  28838=>"011101010",
  28839=>"011100100",
  28840=>"111101101",
  28841=>"010000110",
  28842=>"001101111",
  28843=>"010100110",
  28844=>"111010110",
  28845=>"111010000",
  28846=>"100111000",
  28847=>"010101011",
  28848=>"001000010",
  28849=>"010111000",
  28850=>"001011010",
  28851=>"001111000",
  28852=>"110100011",
  28853=>"110011101",
  28854=>"100101001",
  28855=>"000001101",
  28856=>"101101101",
  28857=>"101010001",
  28858=>"011110110",
  28859=>"100001010",
  28860=>"110001010",
  28861=>"001101100",
  28862=>"100111101",
  28863=>"101000001",
  28864=>"111101111",
  28865=>"011000110",
  28866=>"010101110",
  28867=>"001111011",
  28868=>"101110101",
  28869=>"110110011",
  28870=>"000001101",
  28871=>"010001000",
  28872=>"101001110",
  28873=>"101110011",
  28874=>"111101001",
  28875=>"111000010",
  28876=>"100000001",
  28877=>"000110100",
  28878=>"100001010",
  28879=>"011110110",
  28880=>"001110001",
  28881=>"010000100",
  28882=>"110101000",
  28883=>"100000100",
  28884=>"010000010",
  28885=>"100011110",
  28886=>"100001000",
  28887=>"110000000",
  28888=>"011010010",
  28889=>"010000100",
  28890=>"101111101",
  28891=>"010001000",
  28892=>"000101111",
  28893=>"010100110",
  28894=>"010010110",
  28895=>"000101110",
  28896=>"110101101",
  28897=>"000100010",
  28898=>"000001011",
  28899=>"011011001",
  28900=>"000110001",
  28901=>"110110101",
  28902=>"111010101",
  28903=>"010011110",
  28904=>"110100101",
  28905=>"000111011",
  28906=>"001000100",
  28907=>"001000001",
  28908=>"101001000",
  28909=>"110000010",
  28910=>"110111101",
  28911=>"110000001",
  28912=>"010101100",
  28913=>"001011011",
  28914=>"101110011",
  28915=>"011001001",
  28916=>"010000000",
  28917=>"110000010",
  28918=>"111111010",
  28919=>"000001011",
  28920=>"110110100",
  28921=>"100010111",
  28922=>"101100111",
  28923=>"110110011",
  28924=>"101000001",
  28925=>"000011010",
  28926=>"011011010",
  28927=>"110000101",
  28928=>"111111000",
  28929=>"000011110",
  28930=>"001101110",
  28931=>"110000100",
  28932=>"110011011",
  28933=>"010100000",
  28934=>"001010110",
  28935=>"001001100",
  28936=>"101010011",
  28937=>"110100101",
  28938=>"101010010",
  28939=>"010100000",
  28940=>"010001101",
  28941=>"110110011",
  28942=>"001001101",
  28943=>"100010000",
  28944=>"001010111",
  28945=>"011000100",
  28946=>"000011111",
  28947=>"001111010",
  28948=>"110110110",
  28949=>"010000110",
  28950=>"110101010",
  28951=>"100011000",
  28952=>"111101111",
  28953=>"001011011",
  28954=>"111101100",
  28955=>"010000010",
  28956=>"111111011",
  28957=>"100001100",
  28958=>"111100010",
  28959=>"010000000",
  28960=>"000000010",
  28961=>"111101011",
  28962=>"100110101",
  28963=>"111110010",
  28964=>"101010000",
  28965=>"111111110",
  28966=>"001010100",
  28967=>"010101010",
  28968=>"111010100",
  28969=>"001100001",
  28970=>"001101000",
  28971=>"110111110",
  28972=>"101110101",
  28973=>"100001010",
  28974=>"011110111",
  28975=>"101110111",
  28976=>"100011001",
  28977=>"111011100",
  28978=>"101010001",
  28979=>"111111101",
  28980=>"000001100",
  28981=>"011000001",
  28982=>"010001100",
  28983=>"010101100",
  28984=>"111000101",
  28985=>"110010000",
  28986=>"111010111",
  28987=>"011101101",
  28988=>"011011000",
  28989=>"000110011",
  28990=>"010110000",
  28991=>"100010011",
  28992=>"100000100",
  28993=>"100101011",
  28994=>"000001010",
  28995=>"100110101",
  28996=>"011010100",
  28997=>"000001110",
  28998=>"101001011",
  28999=>"100011001",
  29000=>"110000101",
  29001=>"010101001",
  29002=>"011000001",
  29003=>"010001010",
  29004=>"011000011",
  29005=>"010010000",
  29006=>"111111110",
  29007=>"100001111",
  29008=>"101000111",
  29009=>"001110110",
  29010=>"010110110",
  29011=>"010000010",
  29012=>"001011011",
  29013=>"000011100",
  29014=>"100000011",
  29015=>"000100011",
  29016=>"011100010",
  29017=>"101001100",
  29018=>"010101111",
  29019=>"001100100",
  29020=>"100100011",
  29021=>"000011100",
  29022=>"011010111",
  29023=>"000100111",
  29024=>"000001010",
  29025=>"000010000",
  29026=>"100001001",
  29027=>"111110001",
  29028=>"111110010",
  29029=>"010000101",
  29030=>"011011010",
  29031=>"001011111",
  29032=>"110010010",
  29033=>"101110100",
  29034=>"000010011",
  29035=>"100001111",
  29036=>"110111110",
  29037=>"100111011",
  29038=>"000111010",
  29039=>"001111011",
  29040=>"110100001",
  29041=>"000110101",
  29042=>"000101101",
  29043=>"001100001",
  29044=>"001011100",
  29045=>"111000101",
  29046=>"111100110",
  29047=>"111010100",
  29048=>"001010101",
  29049=>"100010011",
  29050=>"100111000",
  29051=>"011101000",
  29052=>"001011001",
  29053=>"100011011",
  29054=>"110000101",
  29055=>"110010100",
  29056=>"000001000",
  29057=>"011111011",
  29058=>"110001111",
  29059=>"001110000",
  29060=>"110111101",
  29061=>"111010001",
  29062=>"100100101",
  29063=>"001111110",
  29064=>"101111110",
  29065=>"000000011",
  29066=>"000010000",
  29067=>"001011000",
  29068=>"000101100",
  29069=>"010101111",
  29070=>"000000110",
  29071=>"111101111",
  29072=>"011111110",
  29073=>"001010010",
  29074=>"000101011",
  29075=>"101110100",
  29076=>"111110111",
  29077=>"010101110",
  29078=>"100101010",
  29079=>"110100010",
  29080=>"111001001",
  29081=>"010001011",
  29082=>"111110101",
  29083=>"000010000",
  29084=>"000110010",
  29085=>"110000000",
  29086=>"001100110",
  29087=>"100001111",
  29088=>"100010011",
  29089=>"001000000",
  29090=>"010110000",
  29091=>"000000110",
  29092=>"100011000",
  29093=>"000111111",
  29094=>"110010001",
  29095=>"101010100",
  29096=>"010100011",
  29097=>"111100000",
  29098=>"101011101",
  29099=>"111100011",
  29100=>"111101001",
  29101=>"010001110",
  29102=>"000000100",
  29103=>"100010111",
  29104=>"001000001",
  29105=>"001000011",
  29106=>"011101111",
  29107=>"000010011",
  29108=>"101100111",
  29109=>"001100000",
  29110=>"001001100",
  29111=>"100001010",
  29112=>"111011111",
  29113=>"110011100",
  29114=>"100000110",
  29115=>"100111011",
  29116=>"000101001",
  29117=>"110111000",
  29118=>"000010100",
  29119=>"111000110",
  29120=>"000000011",
  29121=>"000000001",
  29122=>"110101110",
  29123=>"100110001",
  29124=>"000011010",
  29125=>"000110001",
  29126=>"110011010",
  29127=>"010010010",
  29128=>"111000101",
  29129=>"101010001",
  29130=>"001001111",
  29131=>"010000010",
  29132=>"001001101",
  29133=>"110101000",
  29134=>"011110000",
  29135=>"001110000",
  29136=>"111111001",
  29137=>"111011111",
  29138=>"001000010",
  29139=>"101100010",
  29140=>"111010001",
  29141=>"110000111",
  29142=>"000001111",
  29143=>"011010110",
  29144=>"110110011",
  29145=>"111011100",
  29146=>"001101111",
  29147=>"100101011",
  29148=>"000011111",
  29149=>"001011010",
  29150=>"001101101",
  29151=>"101010011",
  29152=>"111110111",
  29153=>"001001111",
  29154=>"111100011",
  29155=>"010011100",
  29156=>"010110000",
  29157=>"000010100",
  29158=>"111100110",
  29159=>"010111101",
  29160=>"010100001",
  29161=>"000100000",
  29162=>"110101000",
  29163=>"011101110",
  29164=>"111101011",
  29165=>"000110110",
  29166=>"111110111",
  29167=>"100110110",
  29168=>"111110001",
  29169=>"001110010",
  29170=>"000001000",
  29171=>"101100111",
  29172=>"010100111",
  29173=>"010101100",
  29174=>"010101100",
  29175=>"100100100",
  29176=>"011110001",
  29177=>"001010101",
  29178=>"001001110",
  29179=>"110010111",
  29180=>"000100011",
  29181=>"000010100",
  29182=>"101001000",
  29183=>"110010001",
  29184=>"100011010",
  29185=>"110100001",
  29186=>"111001000",
  29187=>"110001000",
  29188=>"101001011",
  29189=>"110110111",
  29190=>"111100010",
  29191=>"111111110",
  29192=>"010000110",
  29193=>"110000111",
  29194=>"100000001",
  29195=>"000110111",
  29196=>"111100101",
  29197=>"110011010",
  29198=>"000011101",
  29199=>"000100011",
  29200=>"101001110",
  29201=>"111111000",
  29202=>"010110011",
  29203=>"110100100",
  29204=>"011101010",
  29205=>"001110000",
  29206=>"111011011",
  29207=>"111110110",
  29208=>"000111010",
  29209=>"110000000",
  29210=>"111000110",
  29211=>"010111010",
  29212=>"101100001",
  29213=>"000110010",
  29214=>"111010010",
  29215=>"011100000",
  29216=>"000011001",
  29217=>"111100110",
  29218=>"100001011",
  29219=>"000001101",
  29220=>"111101010",
  29221=>"111011000",
  29222=>"001011000",
  29223=>"100111001",
  29224=>"100000110",
  29225=>"100101000",
  29226=>"011011011",
  29227=>"000001001",
  29228=>"110100101",
  29229=>"011111101",
  29230=>"011011010",
  29231=>"010001000",
  29232=>"111101011",
  29233=>"101110011",
  29234=>"111111110",
  29235=>"001110101",
  29236=>"001000111",
  29237=>"000110010",
  29238=>"001011011",
  29239=>"001110111",
  29240=>"101010110",
  29241=>"100001000",
  29242=>"111100101",
  29243=>"110111000",
  29244=>"000000100",
  29245=>"000100111",
  29246=>"101010001",
  29247=>"000110110",
  29248=>"111000110",
  29249=>"111001111",
  29250=>"000010100",
  29251=>"011111111",
  29252=>"111000101",
  29253=>"100100111",
  29254=>"001011010",
  29255=>"100101001",
  29256=>"100011110",
  29257=>"001010001",
  29258=>"100101101",
  29259=>"111100110",
  29260=>"111110111",
  29261=>"001000101",
  29262=>"000000011",
  29263=>"010001000",
  29264=>"011001010",
  29265=>"001110101",
  29266=>"111011101",
  29267=>"100011111",
  29268=>"010001001",
  29269=>"011010100",
  29270=>"000011100",
  29271=>"001100011",
  29272=>"101001010",
  29273=>"001010101",
  29274=>"111110011",
  29275=>"110001010",
  29276=>"011101101",
  29277=>"010001101",
  29278=>"101010000",
  29279=>"010111101",
  29280=>"100010000",
  29281=>"010001001",
  29282=>"011111100",
  29283=>"100101110",
  29284=>"111111100",
  29285=>"110011001",
  29286=>"001110111",
  29287=>"010111000",
  29288=>"110100000",
  29289=>"100010000",
  29290=>"101100010",
  29291=>"100100000",
  29292=>"101110010",
  29293=>"000101101",
  29294=>"001011000",
  29295=>"110100100",
  29296=>"101100000",
  29297=>"110000000",
  29298=>"001010101",
  29299=>"101011110",
  29300=>"101011011",
  29301=>"100100011",
  29302=>"111111010",
  29303=>"110011010",
  29304=>"100010111",
  29305=>"101110001",
  29306=>"101000110",
  29307=>"001000100",
  29308=>"101001011",
  29309=>"011010100",
  29310=>"010011001",
  29311=>"010011001",
  29312=>"001110110",
  29313=>"110101101",
  29314=>"010011101",
  29315=>"001000011",
  29316=>"111000100",
  29317=>"011000000",
  29318=>"000100100",
  29319=>"110011000",
  29320=>"111111101",
  29321=>"001011000",
  29322=>"111111001",
  29323=>"000010011",
  29324=>"110010011",
  29325=>"100010101",
  29326=>"000100010",
  29327=>"000011001",
  29328=>"101101011",
  29329=>"000011010",
  29330=>"100010000",
  29331=>"010110010",
  29332=>"111110000",
  29333=>"100110110",
  29334=>"001001000",
  29335=>"111001100",
  29336=>"000001011",
  29337=>"111001100",
  29338=>"010010011",
  29339=>"101010110",
  29340=>"000110010",
  29341=>"011011000",
  29342=>"010011110",
  29343=>"000010000",
  29344=>"010011001",
  29345=>"011001100",
  29346=>"000000011",
  29347=>"101000010",
  29348=>"100100010",
  29349=>"011100001",
  29350=>"110111011",
  29351=>"010110001",
  29352=>"000010010",
  29353=>"100111000",
  29354=>"100110011",
  29355=>"010011110",
  29356=>"011001101",
  29357=>"001000110",
  29358=>"011100100",
  29359=>"011001100",
  29360=>"010001100",
  29361=>"011110011",
  29362=>"010000111",
  29363=>"111101001",
  29364=>"100100011",
  29365=>"111110010",
  29366=>"010100100",
  29367=>"001101010",
  29368=>"000000101",
  29369=>"100111010",
  29370=>"000001100",
  29371=>"100010011",
  29372=>"001101010",
  29373=>"111011110",
  29374=>"110101101",
  29375=>"001111000",
  29376=>"000101100",
  29377=>"100111011",
  29378=>"100011100",
  29379=>"110101110",
  29380=>"111000111",
  29381=>"010001010",
  29382=>"111010000",
  29383=>"000101111",
  29384=>"001000100",
  29385=>"110011111",
  29386=>"101010001",
  29387=>"110100011",
  29388=>"111101101",
  29389=>"010111111",
  29390=>"001100011",
  29391=>"010001000",
  29392=>"111000100",
  29393=>"000100000",
  29394=>"101011000",
  29395=>"000000100",
  29396=>"011001011",
  29397=>"100101110",
  29398=>"101000011",
  29399=>"011100000",
  29400=>"000011010",
  29401=>"111101100",
  29402=>"111000000",
  29403=>"011001100",
  29404=>"100101010",
  29405=>"011100001",
  29406=>"000000100",
  29407=>"101011001",
  29408=>"101010000",
  29409=>"011110000",
  29410=>"010011110",
  29411=>"111110110",
  29412=>"111001100",
  29413=>"000100111",
  29414=>"110100001",
  29415=>"111101101",
  29416=>"100010111",
  29417=>"110001100",
  29418=>"110001101",
  29419=>"011011010",
  29420=>"001011100",
  29421=>"010010010",
  29422=>"100110011",
  29423=>"001001001",
  29424=>"010000001",
  29425=>"110111110",
  29426=>"110001101",
  29427=>"110111001",
  29428=>"011100011",
  29429=>"111010000",
  29430=>"001101111",
  29431=>"101000110",
  29432=>"110100110",
  29433=>"000100001",
  29434=>"011111001",
  29435=>"101100111",
  29436=>"011011100",
  29437=>"010110001",
  29438=>"111101010",
  29439=>"011010010",
  29440=>"111110010",
  29441=>"001110100",
  29442=>"110101111",
  29443=>"010000100",
  29444=>"001010111",
  29445=>"000000110",
  29446=>"111010110",
  29447=>"111000001",
  29448=>"000001011",
  29449=>"111101110",
  29450=>"100001011",
  29451=>"001001100",
  29452=>"011010001",
  29453=>"110111111",
  29454=>"110101011",
  29455=>"101110111",
  29456=>"100010111",
  29457=>"111001000",
  29458=>"000001000",
  29459=>"110101011",
  29460=>"110101110",
  29461=>"000001011",
  29462=>"100000100",
  29463=>"010001111",
  29464=>"111011000",
  29465=>"001001111",
  29466=>"011110100",
  29467=>"100001001",
  29468=>"010010101",
  29469=>"101111001",
  29470=>"001110010",
  29471=>"110011101",
  29472=>"011000001",
  29473=>"111010000",
  29474=>"001001111",
  29475=>"101001010",
  29476=>"000100100",
  29477=>"000001010",
  29478=>"001100111",
  29479=>"111011011",
  29480=>"010111001",
  29481=>"110111010",
  29482=>"101000100",
  29483=>"100111111",
  29484=>"101110111",
  29485=>"100111001",
  29486=>"101010000",
  29487=>"111001110",
  29488=>"110110010",
  29489=>"101111110",
  29490=>"001001110",
  29491=>"001101101",
  29492=>"101010101",
  29493=>"011101000",
  29494=>"101100110",
  29495=>"000101111",
  29496=>"101111101",
  29497=>"000100000",
  29498=>"000010010",
  29499=>"001000001",
  29500=>"010001001",
  29501=>"001011111",
  29502=>"010011001",
  29503=>"010001110",
  29504=>"100011101",
  29505=>"110000010",
  29506=>"111110111",
  29507=>"000010110",
  29508=>"110111100",
  29509=>"000001110",
  29510=>"101000001",
  29511=>"101101111",
  29512=>"001110111",
  29513=>"010001011",
  29514=>"110101111",
  29515=>"000011000",
  29516=>"010101110",
  29517=>"001111000",
  29518=>"011100001",
  29519=>"001000010",
  29520=>"010100000",
  29521=>"011111111",
  29522=>"011010101",
  29523=>"011101111",
  29524=>"111100000",
  29525=>"111000100",
  29526=>"100100010",
  29527=>"101101101",
  29528=>"011010110",
  29529=>"001011100",
  29530=>"011110101",
  29531=>"001001000",
  29532=>"001100000",
  29533=>"000000101",
  29534=>"010110000",
  29535=>"001001010",
  29536=>"000001100",
  29537=>"100100010",
  29538=>"000010110",
  29539=>"101010110",
  29540=>"010110001",
  29541=>"100111000",
  29542=>"001011011",
  29543=>"001010111",
  29544=>"000001101",
  29545=>"111001001",
  29546=>"011000110",
  29547=>"001001000",
  29548=>"000011101",
  29549=>"111010010",
  29550=>"110101100",
  29551=>"110010100",
  29552=>"010011111",
  29553=>"010110110",
  29554=>"000110100",
  29555=>"110110101",
  29556=>"010010001",
  29557=>"110111101",
  29558=>"011010011",
  29559=>"000001101",
  29560=>"111001010",
  29561=>"101010110",
  29562=>"101110101",
  29563=>"011000111",
  29564=>"010111010",
  29565=>"100111111",
  29566=>"001101111",
  29567=>"010110011",
  29568=>"011011111",
  29569=>"110010011",
  29570=>"101010111",
  29571=>"000011100",
  29572=>"110111111",
  29573=>"000111001",
  29574=>"001000000",
  29575=>"101110010",
  29576=>"100010100",
  29577=>"001100011",
  29578=>"010000001",
  29579=>"111101100",
  29580=>"011000111",
  29581=>"000010001",
  29582=>"000111111",
  29583=>"101001111",
  29584=>"110111101",
  29585=>"100001110",
  29586=>"100001100",
  29587=>"111011101",
  29588=>"010111000",
  29589=>"110011101",
  29590=>"010001001",
  29591=>"110000111",
  29592=>"100010001",
  29593=>"110100111",
  29594=>"111100101",
  29595=>"111101101",
  29596=>"011011010",
  29597=>"000001101",
  29598=>"000111011",
  29599=>"111011010",
  29600=>"011000001",
  29601=>"001101101",
  29602=>"010101000",
  29603=>"111001110",
  29604=>"111101000",
  29605=>"011101110",
  29606=>"001000010",
  29607=>"101100001",
  29608=>"011111111",
  29609=>"111111101",
  29610=>"101010100",
  29611=>"011100000",
  29612=>"100001000",
  29613=>"000001000",
  29614=>"110010110",
  29615=>"011101010",
  29616=>"000101111",
  29617=>"001100000",
  29618=>"001011100",
  29619=>"000010100",
  29620=>"010101001",
  29621=>"101001111",
  29622=>"111111110",
  29623=>"100000000",
  29624=>"100000001",
  29625=>"001111111",
  29626=>"100101000",
  29627=>"110100000",
  29628=>"110011001",
  29629=>"011001111",
  29630=>"110001101",
  29631=>"010101110",
  29632=>"110110001",
  29633=>"000001010",
  29634=>"111000110",
  29635=>"011000110",
  29636=>"001111010",
  29637=>"100011101",
  29638=>"101111101",
  29639=>"110011111",
  29640=>"010111001",
  29641=>"010010011",
  29642=>"101001101",
  29643=>"111101000",
  29644=>"100000111",
  29645=>"111111110",
  29646=>"011000110",
  29647=>"001100111",
  29648=>"010110101",
  29649=>"110110110",
  29650=>"111001111",
  29651=>"100001100",
  29652=>"100110001",
  29653=>"000110000",
  29654=>"101000111",
  29655=>"111000000",
  29656=>"101011101",
  29657=>"101110110",
  29658=>"101110000",
  29659=>"100011100",
  29660=>"111011000",
  29661=>"010011000",
  29662=>"110111011",
  29663=>"110001100",
  29664=>"000000110",
  29665=>"101100110",
  29666=>"001000000",
  29667=>"010011000",
  29668=>"000101011",
  29669=>"101111001",
  29670=>"101011101",
  29671=>"100011011",
  29672=>"001111111",
  29673=>"101000000",
  29674=>"111001001",
  29675=>"111101001",
  29676=>"010101111",
  29677=>"010011100",
  29678=>"110110000",
  29679=>"011110011",
  29680=>"100100110",
  29681=>"000111001",
  29682=>"011110010",
  29683=>"011000000",
  29684=>"001010100",
  29685=>"101011010",
  29686=>"111000110",
  29687=>"111001001",
  29688=>"110111001",
  29689=>"110100101",
  29690=>"000000011",
  29691=>"000011100",
  29692=>"001110011",
  29693=>"100001110",
  29694=>"101011110",
  29695=>"011101001",
  29696=>"010000011",
  29697=>"100000101",
  29698=>"100010000",
  29699=>"011100001",
  29700=>"000001001",
  29701=>"101011111",
  29702=>"100011011",
  29703=>"011100001",
  29704=>"101110001",
  29705=>"111110100",
  29706=>"001001100",
  29707=>"000100000",
  29708=>"100001011",
  29709=>"100111110",
  29710=>"000100000",
  29711=>"010001111",
  29712=>"000101010",
  29713=>"011000011",
  29714=>"001000101",
  29715=>"011100000",
  29716=>"000101000",
  29717=>"100100010",
  29718=>"111111101",
  29719=>"111100010",
  29720=>"100000011",
  29721=>"000001010",
  29722=>"101110110",
  29723=>"110111011",
  29724=>"101011101",
  29725=>"001101011",
  29726=>"101100000",
  29727=>"100111011",
  29728=>"100110000",
  29729=>"010011001",
  29730=>"011100011",
  29731=>"101100111",
  29732=>"100010101",
  29733=>"100010111",
  29734=>"111101011",
  29735=>"101001110",
  29736=>"011001110",
  29737=>"000010100",
  29738=>"000010000",
  29739=>"010101001",
  29740=>"010000110",
  29741=>"000011011",
  29742=>"101001001",
  29743=>"111111011",
  29744=>"111111001",
  29745=>"110000011",
  29746=>"100001111",
  29747=>"010000100",
  29748=>"101000001",
  29749=>"111101101",
  29750=>"101010111",
  29751=>"010111111",
  29752=>"100101010",
  29753=>"010100000",
  29754=>"000101000",
  29755=>"000001101",
  29756=>"001000100",
  29757=>"010110110",
  29758=>"101010010",
  29759=>"000011111",
  29760=>"011110100",
  29761=>"001010011",
  29762=>"000001110",
  29763=>"110110100",
  29764=>"111011101",
  29765=>"010110001",
  29766=>"101010011",
  29767=>"100001101",
  29768=>"101001010",
  29769=>"011010001",
  29770=>"000001001",
  29771=>"110100001",
  29772=>"000000000",
  29773=>"110110010",
  29774=>"111110101",
  29775=>"000111001",
  29776=>"010100111",
  29777=>"011110111",
  29778=>"000011001",
  29779=>"001010111",
  29780=>"101000100",
  29781=>"111010111",
  29782=>"010111011",
  29783=>"110001010",
  29784=>"110101000",
  29785=>"110111110",
  29786=>"101000110",
  29787=>"010001011",
  29788=>"000001111",
  29789=>"110001111",
  29790=>"000100110",
  29791=>"100101111",
  29792=>"001011101",
  29793=>"111001100",
  29794=>"011111100",
  29795=>"001010110",
  29796=>"010001001",
  29797=>"111001010",
  29798=>"011001111",
  29799=>"000000011",
  29800=>"100001010",
  29801=>"010100110",
  29802=>"001100000",
  29803=>"111001011",
  29804=>"001001111",
  29805=>"101000000",
  29806=>"011000100",
  29807=>"010010101",
  29808=>"000010000",
  29809=>"001110010",
  29810=>"111101000",
  29811=>"101111011",
  29812=>"111001111",
  29813=>"100011111",
  29814=>"010100001",
  29815=>"101001001",
  29816=>"010100110",
  29817=>"111011011",
  29818=>"000110010",
  29819=>"101001110",
  29820=>"011001010",
  29821=>"110100111",
  29822=>"001111100",
  29823=>"010011000",
  29824=>"110001000",
  29825=>"100100100",
  29826=>"110110100",
  29827=>"101010000",
  29828=>"001001010",
  29829=>"000111011",
  29830=>"000001001",
  29831=>"011111000",
  29832=>"101110100",
  29833=>"101010100",
  29834=>"000100011",
  29835=>"011010001",
  29836=>"110001100",
  29837=>"010101000",
  29838=>"011001111",
  29839=>"100101001",
  29840=>"100011100",
  29841=>"000100100",
  29842=>"001100100",
  29843=>"001101110",
  29844=>"100010101",
  29845=>"110100110",
  29846=>"001111001",
  29847=>"000100000",
  29848=>"110010101",
  29849=>"011111001",
  29850=>"010001011",
  29851=>"100000111",
  29852=>"011111111",
  29853=>"100001001",
  29854=>"111110010",
  29855=>"010011111",
  29856=>"100010001",
  29857=>"000000000",
  29858=>"000101111",
  29859=>"001010001",
  29860=>"000000011",
  29861=>"101011010",
  29862=>"001100101",
  29863=>"111110111",
  29864=>"000101001",
  29865=>"010110111",
  29866=>"101101111",
  29867=>"111011110",
  29868=>"001010000",
  29869=>"000110111",
  29870=>"011100001",
  29871=>"110101000",
  29872=>"100110110",
  29873=>"000111000",
  29874=>"110001110",
  29875=>"001100010",
  29876=>"111001000",
  29877=>"110100000",
  29878=>"100011101",
  29879=>"101111010",
  29880=>"000100010",
  29881=>"100010100",
  29882=>"110111111",
  29883=>"000001101",
  29884=>"001101001",
  29885=>"011001111",
  29886=>"000100011",
  29887=>"010110011",
  29888=>"000101100",
  29889=>"010001000",
  29890=>"010010011",
  29891=>"101111101",
  29892=>"100000000",
  29893=>"001011011",
  29894=>"010011100",
  29895=>"100111101",
  29896=>"111110010",
  29897=>"101101110",
  29898=>"011111001",
  29899=>"111011000",
  29900=>"110110001",
  29901=>"111001110",
  29902=>"000000001",
  29903=>"101000110",
  29904=>"100000000",
  29905=>"110010010",
  29906=>"010010011",
  29907=>"101001111",
  29908=>"110011011",
  29909=>"100011010",
  29910=>"010001111",
  29911=>"100100100",
  29912=>"010011110",
  29913=>"111000011",
  29914=>"100000110",
  29915=>"101010000",
  29916=>"101111110",
  29917=>"101010101",
  29918=>"110011101",
  29919=>"001001000",
  29920=>"010010000",
  29921=>"101001111",
  29922=>"001100111",
  29923=>"011110100",
  29924=>"000100000",
  29925=>"011001110",
  29926=>"101001101",
  29927=>"011000110",
  29928=>"110000001",
  29929=>"010111010",
  29930=>"000100010",
  29931=>"001000111",
  29932=>"001101010",
  29933=>"101100111",
  29934=>"110101110",
  29935=>"010011111",
  29936=>"110100010",
  29937=>"010001000",
  29938=>"001100100",
  29939=>"001111010",
  29940=>"000111110",
  29941=>"111111110",
  29942=>"011010010",
  29943=>"001010011",
  29944=>"101000100",
  29945=>"111100110",
  29946=>"101001101",
  29947=>"110101011",
  29948=>"000001001",
  29949=>"101101101",
  29950=>"000101010",
  29951=>"001010001",
  29952=>"000011111",
  29953=>"001111101",
  29954=>"111101100",
  29955=>"110011111",
  29956=>"110011011",
  29957=>"111000011",
  29958=>"100011100",
  29959=>"000110001",
  29960=>"001110000",
  29961=>"111110110",
  29962=>"000111001",
  29963=>"011011000",
  29964=>"011010100",
  29965=>"111100011",
  29966=>"000100011",
  29967=>"100010111",
  29968=>"010111011",
  29969=>"111101110",
  29970=>"010110011",
  29971=>"011100001",
  29972=>"010000000",
  29973=>"111001011",
  29974=>"100110010",
  29975=>"001010101",
  29976=>"101101101",
  29977=>"111001100",
  29978=>"100110001",
  29979=>"010010010",
  29980=>"011000111",
  29981=>"100010110",
  29982=>"111100110",
  29983=>"000101100",
  29984=>"001001001",
  29985=>"000101000",
  29986=>"100000001",
  29987=>"111010110",
  29988=>"111100101",
  29989=>"101100011",
  29990=>"011000010",
  29991=>"110000001",
  29992=>"011000011",
  29993=>"000100001",
  29994=>"001100101",
  29995=>"011001100",
  29996=>"001000000",
  29997=>"000000110",
  29998=>"011000000",
  29999=>"101111110",
  30000=>"011000000",
  30001=>"010110110",
  30002=>"011010001",
  30003=>"001100101",
  30004=>"110011010",
  30005=>"101000010",
  30006=>"001001100",
  30007=>"111011110",
  30008=>"011100011",
  30009=>"010000001",
  30010=>"001000011",
  30011=>"010100111",
  30012=>"010001111",
  30013=>"100100001",
  30014=>"100110010",
  30015=>"010110100",
  30016=>"000010010",
  30017=>"111010000",
  30018=>"000110110",
  30019=>"100011101",
  30020=>"100011001",
  30021=>"000111110",
  30022=>"001000011",
  30023=>"101000000",
  30024=>"110000010",
  30025=>"111010111",
  30026=>"000101111",
  30027=>"000000010",
  30028=>"111001000",
  30029=>"010010101",
  30030=>"000011110",
  30031=>"100101100",
  30032=>"000100100",
  30033=>"010001101",
  30034=>"001111010",
  30035=>"001010000",
  30036=>"001011110",
  30037=>"101010111",
  30038=>"111011101",
  30039=>"110000100",
  30040=>"011000011",
  30041=>"110000101",
  30042=>"110010000",
  30043=>"100100111",
  30044=>"100111001",
  30045=>"010000110",
  30046=>"100000101",
  30047=>"110010100",
  30048=>"000011101",
  30049=>"110111010",
  30050=>"000000011",
  30051=>"110110000",
  30052=>"000000001",
  30053=>"101010001",
  30054=>"101000100",
  30055=>"000111010",
  30056=>"000010100",
  30057=>"001000001",
  30058=>"101100011",
  30059=>"011001001",
  30060=>"001010000",
  30061=>"011101100",
  30062=>"000110100",
  30063=>"010011100",
  30064=>"100011110",
  30065=>"110111110",
  30066=>"100011111",
  30067=>"011110111",
  30068=>"100110011",
  30069=>"100000000",
  30070=>"010111100",
  30071=>"001000000",
  30072=>"001010110",
  30073=>"000111111",
  30074=>"010111001",
  30075=>"101111000",
  30076=>"011001111",
  30077=>"100011100",
  30078=>"001111000",
  30079=>"110100000",
  30080=>"101000111",
  30081=>"001000111",
  30082=>"000101010",
  30083=>"011011001",
  30084=>"011111101",
  30085=>"111101101",
  30086=>"100100110",
  30087=>"110010110",
  30088=>"100101010",
  30089=>"010010111",
  30090=>"100111000",
  30091=>"000000011",
  30092=>"100100000",
  30093=>"011010000",
  30094=>"010001001",
  30095=>"111111101",
  30096=>"101011010",
  30097=>"001000010",
  30098=>"001101110",
  30099=>"101101101",
  30100=>"001110000",
  30101=>"110010011",
  30102=>"000000110",
  30103=>"101111001",
  30104=>"110101000",
  30105=>"000000011",
  30106=>"111111010",
  30107=>"010101101",
  30108=>"100001111",
  30109=>"110000100",
  30110=>"111110111",
  30111=>"001000000",
  30112=>"011110001",
  30113=>"111101010",
  30114=>"111100000",
  30115=>"111100001",
  30116=>"110100100",
  30117=>"010010000",
  30118=>"011100011",
  30119=>"101000111",
  30120=>"101000011",
  30121=>"001010000",
  30122=>"010000000",
  30123=>"010101101",
  30124=>"111100011",
  30125=>"010101101",
  30126=>"000110110",
  30127=>"001001001",
  30128=>"011101011",
  30129=>"110110100",
  30130=>"011110000",
  30131=>"001000101",
  30132=>"001110110",
  30133=>"011010010",
  30134=>"010110011",
  30135=>"111010110",
  30136=>"101001100",
  30137=>"001010000",
  30138=>"100100101",
  30139=>"100011000",
  30140=>"010001001",
  30141=>"111110001",
  30142=>"001001101",
  30143=>"111111000",
  30144=>"100010011",
  30145=>"100010001",
  30146=>"101110100",
  30147=>"110111010",
  30148=>"000010000",
  30149=>"100100001",
  30150=>"010000100",
  30151=>"001011001",
  30152=>"111100000",
  30153=>"100100011",
  30154=>"010101001",
  30155=>"111100001",
  30156=>"011101010",
  30157=>"110100110",
  30158=>"110010010",
  30159=>"111010001",
  30160=>"010000100",
  30161=>"111001011",
  30162=>"000110011",
  30163=>"010010000",
  30164=>"101110111",
  30165=>"101111111",
  30166=>"000110010",
  30167=>"001111001",
  30168=>"101110010",
  30169=>"001110011",
  30170=>"110101010",
  30171=>"011010100",
  30172=>"001011000",
  30173=>"011101011",
  30174=>"101011010",
  30175=>"010111010",
  30176=>"010111110",
  30177=>"011110010",
  30178=>"111100110",
  30179=>"011011100",
  30180=>"110101111",
  30181=>"000000001",
  30182=>"100111101",
  30183=>"001111111",
  30184=>"110001100",
  30185=>"110011010",
  30186=>"000000000",
  30187=>"100001101",
  30188=>"100110100",
  30189=>"010110101",
  30190=>"010000011",
  30191=>"001011001",
  30192=>"100110011",
  30193=>"010010101",
  30194=>"110001001",
  30195=>"001010010",
  30196=>"111000100",
  30197=>"011100010",
  30198=>"001101111",
  30199=>"100011000",
  30200=>"100100101",
  30201=>"111011000",
  30202=>"110010010",
  30203=>"000011111",
  30204=>"111111001",
  30205=>"000001101",
  30206=>"110100010",
  30207=>"110000010",
  30208=>"111101110",
  30209=>"101100011",
  30210=>"100011110",
  30211=>"101011001",
  30212=>"010001101",
  30213=>"010011110",
  30214=>"100100100",
  30215=>"110101000",
  30216=>"100010101",
  30217=>"111101010",
  30218=>"000010110",
  30219=>"110100000",
  30220=>"101010110",
  30221=>"111100010",
  30222=>"011100111",
  30223=>"010101001",
  30224=>"000011010",
  30225=>"010001010",
  30226=>"111011101",
  30227=>"011111111",
  30228=>"110001011",
  30229=>"011100110",
  30230=>"001000110",
  30231=>"011001011",
  30232=>"010001000",
  30233=>"011100101",
  30234=>"100111110",
  30235=>"001001010",
  30236=>"010001011",
  30237=>"000110011",
  30238=>"011111100",
  30239=>"101110110",
  30240=>"100110100",
  30241=>"010011101",
  30242=>"111101000",
  30243=>"000011011",
  30244=>"010111110",
  30245=>"011100010",
  30246=>"001110010",
  30247=>"110000010",
  30248=>"100001100",
  30249=>"101011101",
  30250=>"100110101",
  30251=>"111110111",
  30252=>"110111110",
  30253=>"001001101",
  30254=>"010011000",
  30255=>"100001100",
  30256=>"110001110",
  30257=>"001011010",
  30258=>"101101101",
  30259=>"111101001",
  30260=>"101101000",
  30261=>"111100000",
  30262=>"100110011",
  30263=>"110100010",
  30264=>"001010001",
  30265=>"011111100",
  30266=>"110111110",
  30267=>"100000011",
  30268=>"110000100",
  30269=>"001100100",
  30270=>"101111100",
  30271=>"011100010",
  30272=>"111010110",
  30273=>"011001001",
  30274=>"100101000",
  30275=>"101010000",
  30276=>"010011001",
  30277=>"000000011",
  30278=>"001100101",
  30279=>"101011001",
  30280=>"101111110",
  30281=>"010000011",
  30282=>"001000000",
  30283=>"110001000",
  30284=>"001000011",
  30285=>"101010001",
  30286=>"100101000",
  30287=>"111011100",
  30288=>"010000000",
  30289=>"110010011",
  30290=>"011111011",
  30291=>"001011001",
  30292=>"100000001",
  30293=>"110000011",
  30294=>"100001111",
  30295=>"101100001",
  30296=>"001000000",
  30297=>"110100011",
  30298=>"100100001",
  30299=>"101010111",
  30300=>"000101010",
  30301=>"010010101",
  30302=>"011010101",
  30303=>"011100001",
  30304=>"100100111",
  30305=>"010010111",
  30306=>"011001110",
  30307=>"100011110",
  30308=>"111110111",
  30309=>"001010111",
  30310=>"110010010",
  30311=>"101100101",
  30312=>"110100001",
  30313=>"000010101",
  30314=>"111111101",
  30315=>"011011111",
  30316=>"001101111",
  30317=>"110101011",
  30318=>"100010001",
  30319=>"001101101",
  30320=>"111100101",
  30321=>"000011000",
  30322=>"011011110",
  30323=>"000001000",
  30324=>"100001001",
  30325=>"010011001",
  30326=>"011000011",
  30327=>"011001100",
  30328=>"110010000",
  30329=>"010111110",
  30330=>"001100010",
  30331=>"010101111",
  30332=>"010010011",
  30333=>"001011110",
  30334=>"000001010",
  30335=>"011011001",
  30336=>"000000110",
  30337=>"111101010",
  30338=>"010010010",
  30339=>"110001110",
  30340=>"000000100",
  30341=>"101101111",
  30342=>"110001010",
  30343=>"111010000",
  30344=>"011111001",
  30345=>"001110000",
  30346=>"100101110",
  30347=>"110000110",
  30348=>"111001110",
  30349=>"101000110",
  30350=>"011000111",
  30351=>"110000111",
  30352=>"000001111",
  30353=>"101000011",
  30354=>"101011111",
  30355=>"110001100",
  30356=>"001100101",
  30357=>"100110000",
  30358=>"011111011",
  30359=>"101111101",
  30360=>"110000100",
  30361=>"010011010",
  30362=>"110000001",
  30363=>"110110101",
  30364=>"011011101",
  30365=>"001100101",
  30366=>"001011000",
  30367=>"101010100",
  30368=>"111101001",
  30369=>"100011010",
  30370=>"011110001",
  30371=>"110001101",
  30372=>"111111011",
  30373=>"000111101",
  30374=>"110111100",
  30375=>"101010011",
  30376=>"011100011",
  30377=>"000001001",
  30378=>"001100000",
  30379=>"001101001",
  30380=>"001000011",
  30381=>"010101101",
  30382=>"111010111",
  30383=>"111100001",
  30384=>"100110000",
  30385=>"101000000",
  30386=>"101000011",
  30387=>"000001111",
  30388=>"000011000",
  30389=>"111101110",
  30390=>"011101001",
  30391=>"001100010",
  30392=>"110011111",
  30393=>"100101001",
  30394=>"010010110",
  30395=>"011011111",
  30396=>"010100011",
  30397=>"100100101",
  30398=>"101101000",
  30399=>"011101100",
  30400=>"101001111",
  30401=>"100111011",
  30402=>"000100011",
  30403=>"011000110",
  30404=>"111110100",
  30405=>"001000110",
  30406=>"000100100",
  30407=>"101011000",
  30408=>"000000011",
  30409=>"111011010",
  30410=>"100100100",
  30411=>"000111111",
  30412=>"011000100",
  30413=>"111100001",
  30414=>"001000111",
  30415=>"000000000",
  30416=>"000000001",
  30417=>"101010100",
  30418=>"000010101",
  30419=>"001001010",
  30420=>"000110110",
  30421=>"110011001",
  30422=>"101100000",
  30423=>"100001000",
  30424=>"010001010",
  30425=>"111100000",
  30426=>"100001100",
  30427=>"000110101",
  30428=>"101001100",
  30429=>"010000000",
  30430=>"000011101",
  30431=>"100111110",
  30432=>"110111100",
  30433=>"011110001",
  30434=>"011100011",
  30435=>"111100010",
  30436=>"110010100",
  30437=>"100101100",
  30438=>"000011110",
  30439=>"011010101",
  30440=>"111110000",
  30441=>"000011111",
  30442=>"011110010",
  30443=>"110110000",
  30444=>"000110000",
  30445=>"111001110",
  30446=>"010101110",
  30447=>"101010100",
  30448=>"010000010",
  30449=>"111100011",
  30450=>"111011100",
  30451=>"001010011",
  30452=>"001110010",
  30453=>"110011010",
  30454=>"000000101",
  30455=>"011101110",
  30456=>"110010111",
  30457=>"010111110",
  30458=>"010111010",
  30459=>"111011100",
  30460=>"010000100",
  30461=>"101001001",
  30462=>"000000011",
  30463=>"111001011",
  30464=>"001011010",
  30465=>"000101100",
  30466=>"101100001",
  30467=>"100010010",
  30468=>"010010100",
  30469=>"111001011",
  30470=>"001010010",
  30471=>"101001011",
  30472=>"100110001",
  30473=>"001111110",
  30474=>"000100100",
  30475=>"010000000",
  30476=>"010011110",
  30477=>"010000110",
  30478=>"111010011",
  30479=>"101110111",
  30480=>"101100110",
  30481=>"000001100",
  30482=>"100001110",
  30483=>"001000110",
  30484=>"110010101",
  30485=>"011010100",
  30486=>"000101100",
  30487=>"110011001",
  30488=>"111001011",
  30489=>"101011000",
  30490=>"000010010",
  30491=>"000010111",
  30492=>"100110111",
  30493=>"000110110",
  30494=>"001010111",
  30495=>"011101111",
  30496=>"100110001",
  30497=>"101110101",
  30498=>"111000011",
  30499=>"111011001",
  30500=>"101110001",
  30501=>"001000111",
  30502=>"111010111",
  30503=>"100101011",
  30504=>"011001011",
  30505=>"000000110",
  30506=>"110101110",
  30507=>"000111101",
  30508=>"000111110",
  30509=>"101000000",
  30510=>"100000011",
  30511=>"001111110",
  30512=>"011111010",
  30513=>"100011110",
  30514=>"100101110",
  30515=>"011001110",
  30516=>"100110001",
  30517=>"011001100",
  30518=>"110111010",
  30519=>"101000011",
  30520=>"101000011",
  30521=>"101101100",
  30522=>"000101001",
  30523=>"111011000",
  30524=>"100100101",
  30525=>"000101000",
  30526=>"001011100",
  30527=>"010100100",
  30528=>"000100000",
  30529=>"000111110",
  30530=>"011100001",
  30531=>"001000100",
  30532=>"000010001",
  30533=>"111000011",
  30534=>"111001110",
  30535=>"100011000",
  30536=>"010010101",
  30537=>"000100110",
  30538=>"010111110",
  30539=>"011010111",
  30540=>"011011010",
  30541=>"110101110",
  30542=>"111111101",
  30543=>"100101011",
  30544=>"101110101",
  30545=>"100101111",
  30546=>"000100010",
  30547=>"111100101",
  30548=>"100011011",
  30549=>"001010010",
  30550=>"010111110",
  30551=>"110010010",
  30552=>"101101011",
  30553=>"011101110",
  30554=>"111011111",
  30555=>"100100011",
  30556=>"111000111",
  30557=>"010100100",
  30558=>"110011101",
  30559=>"110000000",
  30560=>"100011010",
  30561=>"101001110",
  30562=>"001010000",
  30563=>"111010011",
  30564=>"110001010",
  30565=>"111101001",
  30566=>"010101001",
  30567=>"011010010",
  30568=>"010000000",
  30569=>"010111000",
  30570=>"110101000",
  30571=>"011110001",
  30572=>"001111100",
  30573=>"111111001",
  30574=>"000111011",
  30575=>"111000011",
  30576=>"110010001",
  30577=>"110101100",
  30578=>"111001110",
  30579=>"011111010",
  30580=>"011011001",
  30581=>"110001100",
  30582=>"101100001",
  30583=>"001010000",
  30584=>"010100101",
  30585=>"000111000",
  30586=>"110101111",
  30587=>"001000101",
  30588=>"010100000",
  30589=>"110110011",
  30590=>"101101110",
  30591=>"111110110",
  30592=>"011010111",
  30593=>"110110001",
  30594=>"010010100",
  30595=>"001001000",
  30596=>"011110001",
  30597=>"000101011",
  30598=>"110110000",
  30599=>"011000100",
  30600=>"001000001",
  30601=>"110100100",
  30602=>"111011111",
  30603=>"011101100",
  30604=>"100001110",
  30605=>"101010001",
  30606=>"101010111",
  30607=>"101111111",
  30608=>"101001101",
  30609=>"101110001",
  30610=>"000110111",
  30611=>"011001011",
  30612=>"110100111",
  30613=>"011000100",
  30614=>"011000001",
  30615=>"010011000",
  30616=>"111000011",
  30617=>"010011110",
  30618=>"011110011",
  30619=>"100001110",
  30620=>"111000001",
  30621=>"001010101",
  30622=>"001010010",
  30623=>"010101010",
  30624=>"001001110",
  30625=>"010110110",
  30626=>"000100111",
  30627=>"110101000",
  30628=>"000001101",
  30629=>"001101010",
  30630=>"111001101",
  30631=>"010111100",
  30632=>"001011000",
  30633=>"110111100",
  30634=>"111000100",
  30635=>"000111110",
  30636=>"011010110",
  30637=>"110000100",
  30638=>"101111000",
  30639=>"010100011",
  30640=>"101100100",
  30641=>"111111111",
  30642=>"110111001",
  30643=>"010101001",
  30644=>"110100101",
  30645=>"110000000",
  30646=>"000010111",
  30647=>"100110111",
  30648=>"001011110",
  30649=>"100011010",
  30650=>"101111001",
  30651=>"100010001",
  30652=>"111011110",
  30653=>"000010010",
  30654=>"111010111",
  30655=>"111101011",
  30656=>"001110101",
  30657=>"000001010",
  30658=>"001100111",
  30659=>"101010111",
  30660=>"101100001",
  30661=>"101100100",
  30662=>"110101110",
  30663=>"101000001",
  30664=>"111110110",
  30665=>"101000001",
  30666=>"110001010",
  30667=>"101000010",
  30668=>"111010111",
  30669=>"101111100",
  30670=>"100010100",
  30671=>"010001000",
  30672=>"011111111",
  30673=>"010000110",
  30674=>"101011011",
  30675=>"000000000",
  30676=>"011011001",
  30677=>"010111100",
  30678=>"010010101",
  30679=>"001001001",
  30680=>"000000111",
  30681=>"111010000",
  30682=>"110010001",
  30683=>"110100111",
  30684=>"100000000",
  30685=>"110100110",
  30686=>"010111110",
  30687=>"101000110",
  30688=>"010100100",
  30689=>"000010110",
  30690=>"001011011",
  30691=>"011110011",
  30692=>"000101000",
  30693=>"000011101",
  30694=>"111100110",
  30695=>"111100000",
  30696=>"100100011",
  30697=>"010010100",
  30698=>"111011111",
  30699=>"100000001",
  30700=>"110110111",
  30701=>"010010111",
  30702=>"101100101",
  30703=>"010101011",
  30704=>"010110101",
  30705=>"010110100",
  30706=>"111010111",
  30707=>"011111111",
  30708=>"111011010",
  30709=>"000100011",
  30710=>"101010010",
  30711=>"100111011",
  30712=>"110001111",
  30713=>"010011100",
  30714=>"011001100",
  30715=>"000001111",
  30716=>"011101011",
  30717=>"101001110",
  30718=>"110000001",
  30719=>"010011010",
  30720=>"000110010",
  30721=>"010100010",
  30722=>"000110000",
  30723=>"101001101",
  30724=>"111001110",
  30725=>"100010000",
  30726=>"010010011",
  30727=>"010010100",
  30728=>"110111010",
  30729=>"100111101",
  30730=>"000110011",
  30731=>"110101101",
  30732=>"000011100",
  30733=>"110000100",
  30734=>"111100100",
  30735=>"100011100",
  30736=>"101110011",
  30737=>"110101110",
  30738=>"111111011",
  30739=>"111011111",
  30740=>"010101001",
  30741=>"011001000",
  30742=>"111001100",
  30743=>"101000101",
  30744=>"000001010",
  30745=>"100011011",
  30746=>"110000111",
  30747=>"001100101",
  30748=>"111111000",
  30749=>"110101000",
  30750=>"001001110",
  30751=>"000100011",
  30752=>"010111110",
  30753=>"110011101",
  30754=>"101100000",
  30755=>"011110110",
  30756=>"111100010",
  30757=>"100000111",
  30758=>"011010111",
  30759=>"010011110",
  30760=>"101100000",
  30761=>"000101111",
  30762=>"010111111",
  30763=>"010101011",
  30764=>"110000011",
  30765=>"011110011",
  30766=>"111111100",
  30767=>"111000000",
  30768=>"110111000",
  30769=>"010001000",
  30770=>"111000110",
  30771=>"000001010",
  30772=>"011000001",
  30773=>"011011010",
  30774=>"111000010",
  30775=>"110110110",
  30776=>"101000110",
  30777=>"111110110",
  30778=>"110011010",
  30779=>"100011110",
  30780=>"001011010",
  30781=>"000100101",
  30782=>"101011010",
  30783=>"011000001",
  30784=>"000001001",
  30785=>"000010001",
  30786=>"111111101",
  30787=>"110111010",
  30788=>"101111101",
  30789=>"000000100",
  30790=>"111010001",
  30791=>"011011101",
  30792=>"000101000",
  30793=>"000010100",
  30794=>"101000110",
  30795=>"101110100",
  30796=>"101000111",
  30797=>"001100111",
  30798=>"000101010",
  30799=>"110101010",
  30800=>"101110111",
  30801=>"111110100",
  30802=>"011000101",
  30803=>"110101111",
  30804=>"100010000",
  30805=>"111000011",
  30806=>"111000101",
  30807=>"011111001",
  30808=>"110100000",
  30809=>"100011000",
  30810=>"011101110",
  30811=>"000011010",
  30812=>"010010100",
  30813=>"101000100",
  30814=>"010000100",
  30815=>"101111100",
  30816=>"100000001",
  30817=>"100010000",
  30818=>"110111000",
  30819=>"100001001",
  30820=>"100010011",
  30821=>"100111011",
  30822=>"110100000",
  30823=>"011101111",
  30824=>"011010011",
  30825=>"110001100",
  30826=>"011011011",
  30827=>"011010110",
  30828=>"111111100",
  30829=>"100110100",
  30830=>"011111110",
  30831=>"110010010",
  30832=>"101101000",
  30833=>"011011011",
  30834=>"111000110",
  30835=>"111000110",
  30836=>"000000110",
  30837=>"101100011",
  30838=>"111111111",
  30839=>"011101011",
  30840=>"011000010",
  30841=>"101110000",
  30842=>"111000111",
  30843=>"000100011",
  30844=>"011111000",
  30845=>"101110110",
  30846=>"010100011",
  30847=>"011101010",
  30848=>"100010110",
  30849=>"100000100",
  30850=>"011011110",
  30851=>"011111111",
  30852=>"010001111",
  30853=>"110010011",
  30854=>"110001110",
  30855=>"110001100",
  30856=>"010001001",
  30857=>"100100100",
  30858=>"100000100",
  30859=>"101000010",
  30860=>"001010100",
  30861=>"101000100",
  30862=>"111100011",
  30863=>"100110010",
  30864=>"001110000",
  30865=>"110000111",
  30866=>"101000101",
  30867=>"000001110",
  30868=>"000001100",
  30869=>"000100011",
  30870=>"101110010",
  30871=>"010111001",
  30872=>"010111111",
  30873=>"101100011",
  30874=>"011000100",
  30875=>"111011111",
  30876=>"100101011",
  30877=>"100000001",
  30878=>"000111110",
  30879=>"000001101",
  30880=>"010101010",
  30881=>"110000001",
  30882=>"011010100",
  30883=>"001000100",
  30884=>"001010110",
  30885=>"000000111",
  30886=>"001000000",
  30887=>"000011000",
  30888=>"111111011",
  30889=>"011111110",
  30890=>"100001110",
  30891=>"111100010",
  30892=>"100101100",
  30893=>"001001100",
  30894=>"101111111",
  30895=>"111010010",
  30896=>"101001110",
  30897=>"010101110",
  30898=>"111111001",
  30899=>"000101110",
  30900=>"110101000",
  30901=>"100011000",
  30902=>"000111010",
  30903=>"101100000",
  30904=>"100000010",
  30905=>"010011110",
  30906=>"011111011",
  30907=>"001101110",
  30908=>"011010000",
  30909=>"010011000",
  30910=>"011100010",
  30911=>"001011101",
  30912=>"111111100",
  30913=>"001110011",
  30914=>"000101110",
  30915=>"110001010",
  30916=>"111001101",
  30917=>"111001010",
  30918=>"001000110",
  30919=>"110010010",
  30920=>"111010010",
  30921=>"100001011",
  30922=>"111101000",
  30923=>"001101100",
  30924=>"111100110",
  30925=>"110101001",
  30926=>"001000110",
  30927=>"011000001",
  30928=>"000110100",
  30929=>"101010110",
  30930=>"000101011",
  30931=>"101010111",
  30932=>"110001100",
  30933=>"100110011",
  30934=>"101111101",
  30935=>"111010111",
  30936=>"011100100",
  30937=>"100011001",
  30938=>"001111001",
  30939=>"111000001",
  30940=>"011110000",
  30941=>"001001000",
  30942=>"011111011",
  30943=>"001101001",
  30944=>"011000110",
  30945=>"111110001",
  30946=>"011111100",
  30947=>"111000000",
  30948=>"011100011",
  30949=>"110101000",
  30950=>"001001001",
  30951=>"100111000",
  30952=>"011100101",
  30953=>"110010100",
  30954=>"001010101",
  30955=>"100111111",
  30956=>"000101101",
  30957=>"011101111",
  30958=>"111110111",
  30959=>"000111000",
  30960=>"010110011",
  30961=>"001111000",
  30962=>"100101000",
  30963=>"001000100",
  30964=>"111011001",
  30965=>"101101000",
  30966=>"111000011",
  30967=>"001110011",
  30968=>"001110111",
  30969=>"000110001",
  30970=>"001100110",
  30971=>"101000000",
  30972=>"000010110",
  30973=>"110011011",
  30974=>"001000000",
  30975=>"011010001",
  30976=>"011010110",
  30977=>"111100000",
  30978=>"011110000",
  30979=>"000010101",
  30980=>"111000110",
  30981=>"000001111",
  30982=>"101100101",
  30983=>"111110001",
  30984=>"010100101",
  30985=>"101001101",
  30986=>"110110000",
  30987=>"100010100",
  30988=>"000011110",
  30989=>"111111100",
  30990=>"110000011",
  30991=>"000011100",
  30992=>"000110001",
  30993=>"101100100",
  30994=>"010011100",
  30995=>"011101100",
  30996=>"100110111",
  30997=>"101010011",
  30998=>"011011100",
  30999=>"101011011",
  31000=>"010110000",
  31001=>"110111000",
  31002=>"001110000",
  31003=>"000110100",
  31004=>"001110110",
  31005=>"101011011",
  31006=>"001001110",
  31007=>"011101011",
  31008=>"111001111",
  31009=>"101001010",
  31010=>"011111001",
  31011=>"011001100",
  31012=>"100110001",
  31013=>"001001011",
  31014=>"100101111",
  31015=>"000000010",
  31016=>"100000101",
  31017=>"111010000",
  31018=>"001010111",
  31019=>"100111100",
  31020=>"001010000",
  31021=>"111111000",
  31022=>"111000001",
  31023=>"100010110",
  31024=>"001011111",
  31025=>"001000101",
  31026=>"001000001",
  31027=>"100001100",
  31028=>"110011101",
  31029=>"011110000",
  31030=>"111101110",
  31031=>"111010000",
  31032=>"010100010",
  31033=>"110000011",
  31034=>"010011111",
  31035=>"011110011",
  31036=>"000001000",
  31037=>"100100111",
  31038=>"000011101",
  31039=>"001100000",
  31040=>"010011100",
  31041=>"101010011",
  31042=>"011110111",
  31043=>"111111000",
  31044=>"011111011",
  31045=>"010011011",
  31046=>"100110111",
  31047=>"101000101",
  31048=>"110001110",
  31049=>"110000100",
  31050=>"100110010",
  31051=>"111000001",
  31052=>"000110101",
  31053=>"000010000",
  31054=>"110101110",
  31055=>"001001011",
  31056=>"100110101",
  31057=>"010101100",
  31058=>"100000100",
  31059=>"110111111",
  31060=>"000000000",
  31061=>"001001000",
  31062=>"110010000",
  31063=>"001101000",
  31064=>"011110000",
  31065=>"110100111",
  31066=>"110110111",
  31067=>"111010101",
  31068=>"001010011",
  31069=>"101011011",
  31070=>"111001101",
  31071=>"101101001",
  31072=>"111001000",
  31073=>"110001111",
  31074=>"000000110",
  31075=>"101110001",
  31076=>"011111000",
  31077=>"001111011",
  31078=>"011110010",
  31079=>"001101100",
  31080=>"101101000",
  31081=>"100101011",
  31082=>"110111010",
  31083=>"110011101",
  31084=>"000001010",
  31085=>"000010000",
  31086=>"010110110",
  31087=>"000001101",
  31088=>"011001101",
  31089=>"010111100",
  31090=>"000000001",
  31091=>"100100000",
  31092=>"000101101",
  31093=>"010110001",
  31094=>"100000110",
  31095=>"101001000",
  31096=>"001000000",
  31097=>"000101110",
  31098=>"111010010",
  31099=>"010100000",
  31100=>"000111000",
  31101=>"001001000",
  31102=>"000001010",
  31103=>"000001101",
  31104=>"001110010",
  31105=>"011110111",
  31106=>"101111000",
  31107=>"000110110",
  31108=>"101011101",
  31109=>"110111011",
  31110=>"110000110",
  31111=>"010010011",
  31112=>"010010001",
  31113=>"000100100",
  31114=>"110101101",
  31115=>"000011000",
  31116=>"111110100",
  31117=>"001001001",
  31118=>"011111101",
  31119=>"111101110",
  31120=>"100001111",
  31121=>"100001011",
  31122=>"001110111",
  31123=>"001010101",
  31124=>"111111100",
  31125=>"101100101",
  31126=>"010101101",
  31127=>"101101011",
  31128=>"010001101",
  31129=>"010100010",
  31130=>"000001101",
  31131=>"110111101",
  31132=>"001001001",
  31133=>"001101100",
  31134=>"100011010",
  31135=>"101110000",
  31136=>"011000110",
  31137=>"111001010",
  31138=>"010111101",
  31139=>"111100011",
  31140=>"110001100",
  31141=>"010000011",
  31142=>"000001110",
  31143=>"001000000",
  31144=>"001111111",
  31145=>"111110111",
  31146=>"111000100",
  31147=>"111000011",
  31148=>"111010000",
  31149=>"001001100",
  31150=>"101000100",
  31151=>"111100011",
  31152=>"000110101",
  31153=>"111110000",
  31154=>"101000110",
  31155=>"101110100",
  31156=>"000011010",
  31157=>"011011111",
  31158=>"101111000",
  31159=>"001110011",
  31160=>"010010011",
  31161=>"101101111",
  31162=>"000011000",
  31163=>"010001000",
  31164=>"100001001",
  31165=>"111111001",
  31166=>"100000001",
  31167=>"011111100",
  31168=>"100001010",
  31169=>"101001101",
  31170=>"111011010",
  31171=>"000000011",
  31172=>"000101011",
  31173=>"110100110",
  31174=>"011000100",
  31175=>"011110011",
  31176=>"010110000",
  31177=>"110100110",
  31178=>"011100000",
  31179=>"101111111",
  31180=>"110000010",
  31181=>"000010010",
  31182=>"100000011",
  31183=>"100100110",
  31184=>"110001111",
  31185=>"010001101",
  31186=>"000001110",
  31187=>"111000011",
  31188=>"100001101",
  31189=>"010001110",
  31190=>"001101000",
  31191=>"101001110",
  31192=>"011010001",
  31193=>"111111100",
  31194=>"111110100",
  31195=>"010111011",
  31196=>"101001100",
  31197=>"110101000",
  31198=>"010001001",
  31199=>"111001010",
  31200=>"100111000",
  31201=>"101011010",
  31202=>"111011111",
  31203=>"100100100",
  31204=>"101001100",
  31205=>"010100001",
  31206=>"000011011",
  31207=>"101100001",
  31208=>"100100100",
  31209=>"100101111",
  31210=>"010111101",
  31211=>"010000001",
  31212=>"011011100",
  31213=>"100001000",
  31214=>"001000001",
  31215=>"111000010",
  31216=>"111000001",
  31217=>"011110010",
  31218=>"100011100",
  31219=>"001110100",
  31220=>"111100110",
  31221=>"111010111",
  31222=>"011011011",
  31223=>"000101010",
  31224=>"101101110",
  31225=>"101011010",
  31226=>"111100111",
  31227=>"100111110",
  31228=>"001111101",
  31229=>"100000010",
  31230=>"011111001",
  31231=>"010011001",
  31232=>"011011110",
  31233=>"111000101",
  31234=>"011111001",
  31235=>"101001010",
  31236=>"111011111",
  31237=>"001110111",
  31238=>"110011001",
  31239=>"101100100",
  31240=>"110000100",
  31241=>"101110010",
  31242=>"010011111",
  31243=>"111111110",
  31244=>"000000101",
  31245=>"001101010",
  31246=>"101010111",
  31247=>"110110010",
  31248=>"110000011",
  31249=>"111000111",
  31250=>"111000000",
  31251=>"111001011",
  31252=>"000101100",
  31253=>"111110001",
  31254=>"110110111",
  31255=>"001101101",
  31256=>"111111000",
  31257=>"101101110",
  31258=>"000101011",
  31259=>"010100111",
  31260=>"101010100",
  31261=>"000000010",
  31262=>"100101101",
  31263=>"001111110",
  31264=>"011111100",
  31265=>"010010001",
  31266=>"000000101",
  31267=>"011100011",
  31268=>"010011010",
  31269=>"111011001",
  31270=>"010011010",
  31271=>"001000011",
  31272=>"101010110",
  31273=>"000010000",
  31274=>"001000000",
  31275=>"010100110",
  31276=>"000000110",
  31277=>"010001100",
  31278=>"001110011",
  31279=>"000011101",
  31280=>"101001101",
  31281=>"000101010",
  31282=>"110001110",
  31283=>"100100010",
  31284=>"100010101",
  31285=>"000000001",
  31286=>"011000111",
  31287=>"000010101",
  31288=>"100011100",
  31289=>"000000011",
  31290=>"001111110",
  31291=>"011000001",
  31292=>"001110101",
  31293=>"000101100",
  31294=>"001001011",
  31295=>"010001011",
  31296=>"101001100",
  31297=>"000101110",
  31298=>"001001000",
  31299=>"010111001",
  31300=>"111101010",
  31301=>"110110111",
  31302=>"000100110",
  31303=>"010110101",
  31304=>"111110111",
  31305=>"101100100",
  31306=>"010101010",
  31307=>"010000110",
  31308=>"101111100",
  31309=>"110010010",
  31310=>"010000100",
  31311=>"000101000",
  31312=>"001100100",
  31313=>"011011100",
  31314=>"101000111",
  31315=>"101110000",
  31316=>"111010101",
  31317=>"110100010",
  31318=>"100011110",
  31319=>"001000101",
  31320=>"001010010",
  31321=>"001110110",
  31322=>"011110010",
  31323=>"011011111",
  31324=>"000011000",
  31325=>"101101100",
  31326=>"101010110",
  31327=>"110100001",
  31328=>"110100111",
  31329=>"001001001",
  31330=>"100000010",
  31331=>"101110110",
  31332=>"010110110",
  31333=>"001111010",
  31334=>"001010011",
  31335=>"101010111",
  31336=>"111111111",
  31337=>"010111100",
  31338=>"110111010",
  31339=>"011000000",
  31340=>"001111001",
  31341=>"111001011",
  31342=>"111100100",
  31343=>"101001000",
  31344=>"111000011",
  31345=>"110110000",
  31346=>"101100101",
  31347=>"000101110",
  31348=>"111000100",
  31349=>"011101001",
  31350=>"110111101",
  31351=>"010111000",
  31352=>"111100011",
  31353=>"001011010",
  31354=>"100100111",
  31355=>"101011110",
  31356=>"001100011",
  31357=>"000010011",
  31358=>"001000000",
  31359=>"001010001",
  31360=>"000000010",
  31361=>"101110111",
  31362=>"100100111",
  31363=>"111110111",
  31364=>"100100100",
  31365=>"011110110",
  31366=>"110101111",
  31367=>"101110011",
  31368=>"111111101",
  31369=>"110011101",
  31370=>"000100110",
  31371=>"111011000",
  31372=>"110010101",
  31373=>"000010111",
  31374=>"000000000",
  31375=>"100000111",
  31376=>"000011100",
  31377=>"000001111",
  31378=>"011010110",
  31379=>"101100100",
  31380=>"100010000",
  31381=>"010111111",
  31382=>"011000100",
  31383=>"101110011",
  31384=>"101001010",
  31385=>"010111000",
  31386=>"110111010",
  31387=>"111101110",
  31388=>"011111110",
  31389=>"101010111",
  31390=>"001010101",
  31391=>"110111100",
  31392=>"010110010",
  31393=>"100111010",
  31394=>"010111111",
  31395=>"101111100",
  31396=>"010111101",
  31397=>"100000001",
  31398=>"111011100",
  31399=>"011100001",
  31400=>"001101000",
  31401=>"010000100",
  31402=>"001100001",
  31403=>"110101111",
  31404=>"100110000",
  31405=>"011111010",
  31406=>"111110110",
  31407=>"100111110",
  31408=>"100010010",
  31409=>"110010111",
  31410=>"000001111",
  31411=>"101001111",
  31412=>"110110011",
  31413=>"110111101",
  31414=>"100011100",
  31415=>"111001000",
  31416=>"000010101",
  31417=>"000101011",
  31418=>"011001101",
  31419=>"110000000",
  31420=>"111101101",
  31421=>"100001001",
  31422=>"110011000",
  31423=>"100010100",
  31424=>"100011010",
  31425=>"011000010",
  31426=>"000010100",
  31427=>"110111100",
  31428=>"010110001",
  31429=>"110010100",
  31430=>"010010110",
  31431=>"010101100",
  31432=>"111100111",
  31433=>"011011110",
  31434=>"010010011",
  31435=>"101001100",
  31436=>"010101100",
  31437=>"000001001",
  31438=>"110001100",
  31439=>"110100000",
  31440=>"111000001",
  31441=>"000111011",
  31442=>"010011100",
  31443=>"111011111",
  31444=>"010110010",
  31445=>"100101010",
  31446=>"001110011",
  31447=>"110100100",
  31448=>"101100110",
  31449=>"010111101",
  31450=>"100100000",
  31451=>"000011001",
  31452=>"001111011",
  31453=>"111010000",
  31454=>"101100011",
  31455=>"100111001",
  31456=>"101111111",
  31457=>"100010111",
  31458=>"111111011",
  31459=>"111001001",
  31460=>"101101001",
  31461=>"100000000",
  31462=>"111101010",
  31463=>"011100110",
  31464=>"001000010",
  31465=>"111010000",
  31466=>"100000001",
  31467=>"010101001",
  31468=>"111111110",
  31469=>"100001010",
  31470=>"011110000",
  31471=>"010110011",
  31472=>"101010110",
  31473=>"111011110",
  31474=>"011110000",
  31475=>"011111101",
  31476=>"101010001",
  31477=>"110101111",
  31478=>"110101110",
  31479=>"000010000",
  31480=>"000110111",
  31481=>"100001000",
  31482=>"111010001",
  31483=>"100100001",
  31484=>"001101100",
  31485=>"110100011",
  31486=>"100110111",
  31487=>"110100011",
  31488=>"011000000",
  31489=>"111111101",
  31490=>"010010000",
  31491=>"110000011",
  31492=>"101101110",
  31493=>"101011111",
  31494=>"000001111",
  31495=>"101010011",
  31496=>"010101001",
  31497=>"001000010",
  31498=>"001101101",
  31499=>"101010111",
  31500=>"100111110",
  31501=>"110111111",
  31502=>"101000000",
  31503=>"100001110",
  31504=>"101101001",
  31505=>"101011001",
  31506=>"110101011",
  31507=>"110000101",
  31508=>"100100011",
  31509=>"110101000",
  31510=>"111000001",
  31511=>"101100110",
  31512=>"111111110",
  31513=>"010001010",
  31514=>"110111001",
  31515=>"111111100",
  31516=>"001000100",
  31517=>"110001010",
  31518=>"100110011",
  31519=>"110111000",
  31520=>"010110011",
  31521=>"101011000",
  31522=>"010001111",
  31523=>"010001101",
  31524=>"000100000",
  31525=>"111011101",
  31526=>"111111101",
  31527=>"111010100",
  31528=>"011110101",
  31529=>"011111000",
  31530=>"111110111",
  31531=>"101000001",
  31532=>"011011110",
  31533=>"111110111",
  31534=>"100110001",
  31535=>"001001000",
  31536=>"111001111",
  31537=>"100000000",
  31538=>"010001010",
  31539=>"111110110",
  31540=>"100000000",
  31541=>"010001110",
  31542=>"011011110",
  31543=>"100110101",
  31544=>"001111110",
  31545=>"101111111",
  31546=>"111000000",
  31547=>"000010000",
  31548=>"111000100",
  31549=>"101001000",
  31550=>"111111110",
  31551=>"011010011",
  31552=>"011000011",
  31553=>"001010100",
  31554=>"110010001",
  31555=>"101110011",
  31556=>"101011010",
  31557=>"110011001",
  31558=>"000010101",
  31559=>"111110101",
  31560=>"000000101",
  31561=>"001010010",
  31562=>"110000000",
  31563=>"010011011",
  31564=>"100011001",
  31565=>"000001110",
  31566=>"000011010",
  31567=>"011000001",
  31568=>"111010101",
  31569=>"111111010",
  31570=>"100100101",
  31571=>"110111101",
  31572=>"011000100",
  31573=>"000100011",
  31574=>"110000101",
  31575=>"101001010",
  31576=>"100011001",
  31577=>"101101010",
  31578=>"001001110",
  31579=>"100011100",
  31580=>"111110010",
  31581=>"111000101",
  31582=>"100010010",
  31583=>"100010011",
  31584=>"010010010",
  31585=>"010110010",
  31586=>"000100011",
  31587=>"011111000",
  31588=>"000011110",
  31589=>"110000001",
  31590=>"100011001",
  31591=>"110110110",
  31592=>"100000000",
  31593=>"111111110",
  31594=>"101110111",
  31595=>"111001100",
  31596=>"111001010",
  31597=>"010000110",
  31598=>"101101000",
  31599=>"001001011",
  31600=>"111010001",
  31601=>"001011010",
  31602=>"011111001",
  31603=>"111101100",
  31604=>"001011111",
  31605=>"010100011",
  31606=>"110110001",
  31607=>"010010000",
  31608=>"011101001",
  31609=>"000000011",
  31610=>"111111101",
  31611=>"001110101",
  31612=>"011000000",
  31613=>"110101110",
  31614=>"000111000",
  31615=>"001111101",
  31616=>"110010001",
  31617=>"000011110",
  31618=>"101000001",
  31619=>"110110101",
  31620=>"011110000",
  31621=>"101011001",
  31622=>"000100111",
  31623=>"111000010",
  31624=>"101101001",
  31625=>"001100000",
  31626=>"000111100",
  31627=>"010100000",
  31628=>"100101100",
  31629=>"101111010",
  31630=>"000010001",
  31631=>"001100100",
  31632=>"111000101",
  31633=>"000101000",
  31634=>"101010001",
  31635=>"000101001",
  31636=>"001000011",
  31637=>"101011001",
  31638=>"001010001",
  31639=>"010110110",
  31640=>"100010000",
  31641=>"001110110",
  31642=>"100101101",
  31643=>"111011001",
  31644=>"111001100",
  31645=>"011011110",
  31646=>"000010111",
  31647=>"100011010",
  31648=>"111010101",
  31649=>"000010110",
  31650=>"111111111",
  31651=>"010110000",
  31652=>"110101011",
  31653=>"101111111",
  31654=>"101011001",
  31655=>"101011111",
  31656=>"000110000",
  31657=>"011001000",
  31658=>"000100101",
  31659=>"000001000",
  31660=>"011001111",
  31661=>"100010001",
  31662=>"001011110",
  31663=>"011101110",
  31664=>"001100001",
  31665=>"110010000",
  31666=>"111101011",
  31667=>"000101100",
  31668=>"010001011",
  31669=>"110001100",
  31670=>"111010101",
  31671=>"100101000",
  31672=>"111110111",
  31673=>"110101110",
  31674=>"010101001",
  31675=>"100000110",
  31676=>"010011010",
  31677=>"100101000",
  31678=>"100100000",
  31679=>"000011011",
  31680=>"010010001",
  31681=>"010011010",
  31682=>"010111000",
  31683=>"100000011",
  31684=>"100001101",
  31685=>"110111001",
  31686=>"001100011",
  31687=>"111010001",
  31688=>"000000111",
  31689=>"000001111",
  31690=>"011001100",
  31691=>"011101001",
  31692=>"011001100",
  31693=>"001110010",
  31694=>"111110101",
  31695=>"010000100",
  31696=>"111100111",
  31697=>"000001101",
  31698=>"010001001",
  31699=>"000110010",
  31700=>"010101011",
  31701=>"110101101",
  31702=>"001000110",
  31703=>"000101010",
  31704=>"110110110",
  31705=>"101011100",
  31706=>"000000011",
  31707=>"101011011",
  31708=>"000010010",
  31709=>"111011101",
  31710=>"001001111",
  31711=>"010010000",
  31712=>"110101011",
  31713=>"010100100",
  31714=>"001000010",
  31715=>"011110111",
  31716=>"001000010",
  31717=>"011001100",
  31718=>"011101011",
  31719=>"100000000",
  31720=>"000100010",
  31721=>"001111101",
  31722=>"010001011",
  31723=>"111101100",
  31724=>"111100011",
  31725=>"000111010",
  31726=>"010010000",
  31727=>"011000110",
  31728=>"000100000",
  31729=>"101011010",
  31730=>"001111011",
  31731=>"111000111",
  31732=>"000011000",
  31733=>"111010101",
  31734=>"111101011",
  31735=>"101001101",
  31736=>"011100111",
  31737=>"111110100",
  31738=>"011011000",
  31739=>"010101110",
  31740=>"101101111",
  31741=>"111000010",
  31742=>"010010011",
  31743=>"000001111",
  31744=>"101100011",
  31745=>"010011111",
  31746=>"010111011",
  31747=>"110110100",
  31748=>"111111101",
  31749=>"001000011",
  31750=>"101110010",
  31751=>"101100110",
  31752=>"101111011",
  31753=>"001101010",
  31754=>"110000000",
  31755=>"011100010",
  31756=>"110110000",
  31757=>"110110111",
  31758=>"101011000",
  31759=>"001101110",
  31760=>"111011001",
  31761=>"010010111",
  31762=>"000110001",
  31763=>"111001010",
  31764=>"011110000",
  31765=>"000010101",
  31766=>"101011001",
  31767=>"101001100",
  31768=>"101111111",
  31769=>"001011001",
  31770=>"100110001",
  31771=>"101100001",
  31772=>"001100010",
  31773=>"010010100",
  31774=>"101101111",
  31775=>"100100001",
  31776=>"110100111",
  31777=>"001000011",
  31778=>"100110110",
  31779=>"111000111",
  31780=>"100001000",
  31781=>"001111001",
  31782=>"100000010",
  31783=>"100000110",
  31784=>"110100100",
  31785=>"000001110",
  31786=>"101010111",
  31787=>"100101110",
  31788=>"011000111",
  31789=>"111001011",
  31790=>"100010011",
  31791=>"010110000",
  31792=>"000011110",
  31793=>"111001001",
  31794=>"010000110",
  31795=>"110100100",
  31796=>"001101010",
  31797=>"101010010",
  31798=>"100111010",
  31799=>"010000000",
  31800=>"000010011",
  31801=>"001101111",
  31802=>"011000011",
  31803=>"101010001",
  31804=>"101001001",
  31805=>"111101000",
  31806=>"100000000",
  31807=>"110101000",
  31808=>"011010101",
  31809=>"110010001",
  31810=>"111010000",
  31811=>"111000011",
  31812=>"000000001",
  31813=>"101000000",
  31814=>"011110111",
  31815=>"000100011",
  31816=>"101110101",
  31817=>"000111011",
  31818=>"101001100",
  31819=>"110010110",
  31820=>"000000000",
  31821=>"010110011",
  31822=>"111000001",
  31823=>"101110011",
  31824=>"111100101",
  31825=>"111000111",
  31826=>"011100001",
  31827=>"000001111",
  31828=>"001010101",
  31829=>"100101110",
  31830=>"000110111",
  31831=>"000110110",
  31832=>"110000000",
  31833=>"000000101",
  31834=>"011000110",
  31835=>"010000000",
  31836=>"111011000",
  31837=>"100110011",
  31838=>"101100101",
  31839=>"110111001",
  31840=>"100001101",
  31841=>"011111010",
  31842=>"000110101",
  31843=>"101110101",
  31844=>"111110100",
  31845=>"001100000",
  31846=>"001011111",
  31847=>"110000011",
  31848=>"111110101",
  31849=>"011110010",
  31850=>"011100011",
  31851=>"101011000",
  31852=>"001010000",
  31853=>"000010011",
  31854=>"010000111",
  31855=>"010101000",
  31856=>"101111000",
  31857=>"000100101",
  31858=>"001010110",
  31859=>"011010110",
  31860=>"110010111",
  31861=>"100100100",
  31862=>"011100000",
  31863=>"100011001",
  31864=>"110010001",
  31865=>"110110110",
  31866=>"111111101",
  31867=>"001010000",
  31868=>"110010001",
  31869=>"100100010",
  31870=>"100011011",
  31871=>"110111010",
  31872=>"001010101",
  31873=>"000101100",
  31874=>"010000010",
  31875=>"000010010",
  31876=>"011111101",
  31877=>"000111000",
  31878=>"000011100",
  31879=>"101110011",
  31880=>"100100111",
  31881=>"111100111",
  31882=>"111000110",
  31883=>"111110110",
  31884=>"100000000",
  31885=>"001000001",
  31886=>"000100011",
  31887=>"010110101",
  31888=>"110001111",
  31889=>"000110100",
  31890=>"110101011",
  31891=>"110011111",
  31892=>"000011001",
  31893=>"000011111",
  31894=>"111001000",
  31895=>"101111011",
  31896=>"111101111",
  31897=>"000000000",
  31898=>"111100101",
  31899=>"001100010",
  31900=>"001111110",
  31901=>"111101111",
  31902=>"111010100",
  31903=>"011010001",
  31904=>"101001111",
  31905=>"011000010",
  31906=>"011110011",
  31907=>"010110111",
  31908=>"110100101",
  31909=>"100110101",
  31910=>"000010110",
  31911=>"000001011",
  31912=>"110001100",
  31913=>"110101011",
  31914=>"111111011",
  31915=>"100010100",
  31916=>"111010001",
  31917=>"100001111",
  31918=>"010000110",
  31919=>"111001101",
  31920=>"010011100",
  31921=>"011000101",
  31922=>"010111010",
  31923=>"011100101",
  31924=>"001100100",
  31925=>"011100011",
  31926=>"001001001",
  31927=>"011001001",
  31928=>"100000000",
  31929=>"110011000",
  31930=>"100110101",
  31931=>"000011001",
  31932=>"000111001",
  31933=>"101010110",
  31934=>"111101001",
  31935=>"101010111",
  31936=>"111010010",
  31937=>"101100001",
  31938=>"101110111",
  31939=>"001010010",
  31940=>"000011010",
  31941=>"101001110",
  31942=>"100110001",
  31943=>"111000011",
  31944=>"111011010",
  31945=>"011110001",
  31946=>"110011001",
  31947=>"011010111",
  31948=>"101001100",
  31949=>"111111100",
  31950=>"101001010",
  31951=>"111110010",
  31952=>"011110010",
  31953=>"100111110",
  31954=>"000001111",
  31955=>"011110100",
  31956=>"001001110",
  31957=>"010111101",
  31958=>"010111111",
  31959=>"101101010",
  31960=>"001100010",
  31961=>"100111111",
  31962=>"000110011",
  31963=>"111101101",
  31964=>"011101111",
  31965=>"110010111",
  31966=>"001011101",
  31967=>"101100001",
  31968=>"000110100",
  31969=>"110101111",
  31970=>"110010001",
  31971=>"010110000",
  31972=>"101000000",
  31973=>"001000111",
  31974=>"111100000",
  31975=>"110001111",
  31976=>"001100011",
  31977=>"110110111",
  31978=>"010111110",
  31979=>"001011001",
  31980=>"111111110",
  31981=>"001101110",
  31982=>"111000011",
  31983=>"110110100",
  31984=>"101001010",
  31985=>"100010001",
  31986=>"100000100",
  31987=>"110010101",
  31988=>"101011011",
  31989=>"100111111",
  31990=>"010010110",
  31991=>"111101000",
  31992=>"000010011",
  31993=>"100110001",
  31994=>"000101001",
  31995=>"111101001",
  31996=>"010001101",
  31997=>"110110111",
  31998=>"010100000",
  31999=>"001000101",
  32000=>"100001111",
  32001=>"110010110",
  32002=>"101100110",
  32003=>"100011110",
  32004=>"001000111",
  32005=>"000110001",
  32006=>"110110000",
  32007=>"000000111",
  32008=>"000110010",
  32009=>"100100010",
  32010=>"011001100",
  32011=>"111110110",
  32012=>"001000110",
  32013=>"010000110",
  32014=>"100100111",
  32015=>"110110101",
  32016=>"011010101",
  32017=>"100011000",
  32018=>"000001101",
  32019=>"011000110",
  32020=>"001101001",
  32021=>"001010011",
  32022=>"000110101",
  32023=>"110000101",
  32024=>"111010110",
  32025=>"001110110",
  32026=>"100000100",
  32027=>"000101100",
  32028=>"011011011",
  32029=>"010010100",
  32030=>"011110010",
  32031=>"101000110",
  32032=>"111001000",
  32033=>"011010010",
  32034=>"011110100",
  32035=>"010000000",
  32036=>"110010000",
  32037=>"011110000",
  32038=>"000000000",
  32039=>"000000110",
  32040=>"010000111",
  32041=>"010000111",
  32042=>"111110000",
  32043=>"010011100",
  32044=>"011101011",
  32045=>"101000101",
  32046=>"000100010",
  32047=>"010010110",
  32048=>"111001001",
  32049=>"110001110",
  32050=>"001100101",
  32051=>"110101100",
  32052=>"011000100",
  32053=>"000110100",
  32054=>"011000100",
  32055=>"011101101",
  32056=>"101001011",
  32057=>"010000010",
  32058=>"000100111",
  32059=>"110110011",
  32060=>"111000111",
  32061=>"100100011",
  32062=>"111110001",
  32063=>"011011111",
  32064=>"001101000",
  32065=>"101111011",
  32066=>"111001000",
  32067=>"111110011",
  32068=>"001010011",
  32069=>"111000010",
  32070=>"110110101",
  32071=>"010111010",
  32072=>"011000111",
  32073=>"110100000",
  32074=>"001000110",
  32075=>"001111101",
  32076=>"010010111",
  32077=>"010100000",
  32078=>"110101000",
  32079=>"001100000",
  32080=>"011001111",
  32081=>"100110110",
  32082=>"101011100",
  32083=>"011010100",
  32084=>"000011001",
  32085=>"010011010",
  32086=>"111011011",
  32087=>"111001100",
  32088=>"010010100",
  32089=>"001000101",
  32090=>"111001100",
  32091=>"011010000",
  32092=>"000101010",
  32093=>"000010001",
  32094=>"011011000",
  32095=>"100110011",
  32096=>"010000110",
  32097=>"000000001",
  32098=>"010110101",
  32099=>"000111100",
  32100=>"011010110",
  32101=>"101001110",
  32102=>"011111110",
  32103=>"110110100",
  32104=>"111001111",
  32105=>"111110000",
  32106=>"111010110",
  32107=>"100000101",
  32108=>"101100000",
  32109=>"110001111",
  32110=>"001110001",
  32111=>"010000101",
  32112=>"011000000",
  32113=>"001111001",
  32114=>"111111100",
  32115=>"000101100",
  32116=>"110011000",
  32117=>"011010100",
  32118=>"100000000",
  32119=>"001000000",
  32120=>"000010010",
  32121=>"011010111",
  32122=>"110000000",
  32123=>"101001110",
  32124=>"010111001",
  32125=>"110010000",
  32126=>"101001001",
  32127=>"111100011",
  32128=>"100001000",
  32129=>"010000000",
  32130=>"111101001",
  32131=>"101100110",
  32132=>"101010101",
  32133=>"010011000",
  32134=>"100110111",
  32135=>"100000101",
  32136=>"110000001",
  32137=>"011010100",
  32138=>"011010110",
  32139=>"101111001",
  32140=>"010111100",
  32141=>"111010001",
  32142=>"101101001",
  32143=>"101110100",
  32144=>"110111011",
  32145=>"010100011",
  32146=>"011111100",
  32147=>"110100100",
  32148=>"100001001",
  32149=>"110000111",
  32150=>"111101101",
  32151=>"001011000",
  32152=>"010000010",
  32153=>"110101000",
  32154=>"010110001",
  32155=>"110001110",
  32156=>"111100101",
  32157=>"111110100",
  32158=>"101100100",
  32159=>"010111101",
  32160=>"000100101",
  32161=>"100000111",
  32162=>"111011000",
  32163=>"001000100",
  32164=>"100101111",
  32165=>"001001110",
  32166=>"101101010",
  32167=>"100101110",
  32168=>"111100001",
  32169=>"101011110",
  32170=>"100111111",
  32171=>"111100010",
  32172=>"101101001",
  32173=>"110011000",
  32174=>"000111001",
  32175=>"111000000",
  32176=>"100100001",
  32177=>"111111010",
  32178=>"100100100",
  32179=>"111111000",
  32180=>"001011010",
  32181=>"110010100",
  32182=>"110101001",
  32183=>"000010110",
  32184=>"001001101",
  32185=>"010011101",
  32186=>"011010010",
  32187=>"000110101",
  32188=>"011101000",
  32189=>"100011011",
  32190=>"011100010",
  32191=>"010011011",
  32192=>"010100010",
  32193=>"001110101",
  32194=>"111110001",
  32195=>"000100111",
  32196=>"000010001",
  32197=>"000001001",
  32198=>"001011010",
  32199=>"010110001",
  32200=>"100011001",
  32201=>"101010011",
  32202=>"100011000",
  32203=>"111100100",
  32204=>"100101110",
  32205=>"010011110",
  32206=>"011010001",
  32207=>"001010101",
  32208=>"110000011",
  32209=>"101011001",
  32210=>"000100111",
  32211=>"010101010",
  32212=>"011110110",
  32213=>"010100001",
  32214=>"001101011",
  32215=>"010000011",
  32216=>"111111010",
  32217=>"111111110",
  32218=>"010101000",
  32219=>"011101100",
  32220=>"011000011",
  32221=>"101100100",
  32222=>"100101100",
  32223=>"001000011",
  32224=>"010011010",
  32225=>"100001000",
  32226=>"001111110",
  32227=>"101001010",
  32228=>"110011111",
  32229=>"010101010",
  32230=>"001011011",
  32231=>"011100101",
  32232=>"010010000",
  32233=>"111111101",
  32234=>"010011100",
  32235=>"110110110",
  32236=>"000010000",
  32237=>"110111101",
  32238=>"111100000",
  32239=>"000001101",
  32240=>"010110000",
  32241=>"000111010",
  32242=>"111101001",
  32243=>"000010001",
  32244=>"110110100",
  32245=>"111101011",
  32246=>"001011111",
  32247=>"101110110",
  32248=>"111100101",
  32249=>"110111010",
  32250=>"101000111",
  32251=>"101110010",
  32252=>"000000110",
  32253=>"011110100",
  32254=>"100100001",
  32255=>"001110001",
  32256=>"100110100",
  32257=>"101010010",
  32258=>"001010101",
  32259=>"010000100",
  32260=>"011001111",
  32261=>"101011100",
  32262=>"111111110",
  32263=>"000100111",
  32264=>"101101000",
  32265=>"100000000",
  32266=>"101110000",
  32267=>"011010010",
  32268=>"000111100",
  32269=>"100010011",
  32270=>"101100001",
  32271=>"101001000",
  32272=>"011011001",
  32273=>"110111110",
  32274=>"001101110",
  32275=>"000100000",
  32276=>"011100010",
  32277=>"011011110",
  32278=>"111011110",
  32279=>"001010010",
  32280=>"000000100",
  32281=>"101110000",
  32282=>"100110000",
  32283=>"001001100",
  32284=>"101000001",
  32285=>"010100101",
  32286=>"000100000",
  32287=>"011010011",
  32288=>"011101101",
  32289=>"001010001",
  32290=>"000101110",
  32291=>"011100011",
  32292=>"111010001",
  32293=>"101010111",
  32294=>"101001111",
  32295=>"100011001",
  32296=>"010100110",
  32297=>"111001100",
  32298=>"110010111",
  32299=>"000011110",
  32300=>"001011101",
  32301=>"110100011",
  32302=>"011111000",
  32303=>"101100100",
  32304=>"000101001",
  32305=>"000100000",
  32306=>"100001111",
  32307=>"010011111",
  32308=>"010010101",
  32309=>"110111111",
  32310=>"111100111",
  32311=>"010000000",
  32312=>"011110111",
  32313=>"011111001",
  32314=>"101010100",
  32315=>"110110110",
  32316=>"011111010",
  32317=>"101111011",
  32318=>"111111000",
  32319=>"101100100",
  32320=>"101001010",
  32321=>"100010000",
  32322=>"000101110",
  32323=>"010110000",
  32324=>"010100111",
  32325=>"000000100",
  32326=>"111100101",
  32327=>"010101000",
  32328=>"001000011",
  32329=>"101111111",
  32330=>"110110010",
  32331=>"011000010",
  32332=>"000010100",
  32333=>"110111011",
  32334=>"110100101",
  32335=>"001011001",
  32336=>"011101101",
  32337=>"000010000",
  32338=>"110111011",
  32339=>"011011111",
  32340=>"101010111",
  32341=>"001111101",
  32342=>"011000001",
  32343=>"100111000",
  32344=>"111111000",
  32345=>"000111011",
  32346=>"000000110",
  32347=>"110001101",
  32348=>"101011101",
  32349=>"111111101",
  32350=>"011010011",
  32351=>"111100110",
  32352=>"011000010",
  32353=>"011010111",
  32354=>"001101111",
  32355=>"101100011",
  32356=>"101000010",
  32357=>"101111001",
  32358=>"101101010",
  32359=>"001001110",
  32360=>"001010011",
  32361=>"011011101",
  32362=>"001110011",
  32363=>"110110100",
  32364=>"101100000",
  32365=>"100011110",
  32366=>"110001000",
  32367=>"101100110",
  32368=>"001011010",
  32369=>"101101100",
  32370=>"111000100",
  32371=>"110010011",
  32372=>"101010100",
  32373=>"101111101",
  32374=>"100111001",
  32375=>"000001100",
  32376=>"101010011",
  32377=>"100110110",
  32378=>"110011100",
  32379=>"011111001",
  32380=>"000011001",
  32381=>"010001101",
  32382=>"111101101",
  32383=>"111000100",
  32384=>"010100010",
  32385=>"011111100",
  32386=>"100111100",
  32387=>"110100111",
  32388=>"010011111",
  32389=>"010111101",
  32390=>"111100001",
  32391=>"110000100",
  32392=>"100101000",
  32393=>"100010000",
  32394=>"111100011",
  32395=>"011111000",
  32396=>"011111000",
  32397=>"101110111",
  32398=>"101110010",
  32399=>"011111000",
  32400=>"100011010",
  32401=>"110000111",
  32402=>"110100111",
  32403=>"001010000",
  32404=>"100010011",
  32405=>"000000101",
  32406=>"110010010",
  32407=>"100100100",
  32408=>"011101000",
  32409=>"010101010",
  32410=>"100111011",
  32411=>"100111011",
  32412=>"111100101",
  32413=>"111100011",
  32414=>"100111111",
  32415=>"101111000",
  32416=>"111000101",
  32417=>"001011100",
  32418=>"101011110",
  32419=>"001111001",
  32420=>"000110010",
  32421=>"100010000",
  32422=>"100010000",
  32423=>"111110101",
  32424=>"010011000",
  32425=>"101011001",
  32426=>"010100000",
  32427=>"001101101",
  32428=>"011111111",
  32429=>"010111010",
  32430=>"111111001",
  32431=>"111111000",
  32432=>"110000001",
  32433=>"001100100",
  32434=>"001001010",
  32435=>"111111110",
  32436=>"011011000",
  32437=>"010101111",
  32438=>"010100110",
  32439=>"110101100",
  32440=>"110110010",
  32441=>"101111001",
  32442=>"111101111",
  32443=>"111101110",
  32444=>"110000011",
  32445=>"001010000",
  32446=>"111110000",
  32447=>"001000000",
  32448=>"100010010",
  32449=>"010111001",
  32450=>"000000011",
  32451=>"110001010",
  32452=>"010001000",
  32453=>"000111000",
  32454=>"100011110",
  32455=>"001011100",
  32456=>"000100000",
  32457=>"001111100",
  32458=>"110110001",
  32459=>"010000001",
  32460=>"001110110",
  32461=>"010100010",
  32462=>"001000111",
  32463=>"110001010",
  32464=>"000101011",
  32465=>"101111011",
  32466=>"100000110",
  32467=>"000011011",
  32468=>"010110100",
  32469=>"000000000",
  32470=>"000100000",
  32471=>"011011010",
  32472=>"001000100",
  32473=>"110010110",
  32474=>"011000010",
  32475=>"000100100",
  32476=>"010111101",
  32477=>"111011101",
  32478=>"000101111",
  32479=>"000100001",
  32480=>"011000100",
  32481=>"001110001",
  32482=>"100001110",
  32483=>"100001010",
  32484=>"000100000",
  32485=>"011101110",
  32486=>"110010101",
  32487=>"000110000",
  32488=>"101000011",
  32489=>"011000010",
  32490=>"100010000",
  32491=>"101011111",
  32492=>"101000001",
  32493=>"110110110",
  32494=>"001000100",
  32495=>"100110010",
  32496=>"011001101",
  32497=>"010011100",
  32498=>"101011001",
  32499=>"100110111",
  32500=>"100110110",
  32501=>"101111110",
  32502=>"000111010",
  32503=>"011100111",
  32504=>"010011100",
  32505=>"010010110",
  32506=>"000001010",
  32507=>"010001010",
  32508=>"001010100",
  32509=>"000100111",
  32510=>"011100101",
  32511=>"110011100",
  32512=>"001100111",
  32513=>"010000100",
  32514=>"111110010",
  32515=>"110010011",
  32516=>"001110001",
  32517=>"111101100",
  32518=>"100111011",
  32519=>"100101001",
  32520=>"110011010",
  32521=>"100000100",
  32522=>"000000111",
  32523=>"101110100",
  32524=>"100100101",
  32525=>"011100111",
  32526=>"101001010",
  32527=>"001101111",
  32528=>"010101110",
  32529=>"001100010",
  32530=>"010101011",
  32531=>"011010010",
  32532=>"010011011",
  32533=>"101000111",
  32534=>"011000001",
  32535=>"111000110",
  32536=>"011100101",
  32537=>"110001111",
  32538=>"010100111",
  32539=>"100000101",
  32540=>"010000000",
  32541=>"000001010",
  32542=>"101010100",
  32543=>"100101101",
  32544=>"110011000",
  32545=>"011111001",
  32546=>"011111111",
  32547=>"110101101",
  32548=>"011101110",
  32549=>"000000111",
  32550=>"100000110",
  32551=>"101101110",
  32552=>"111101000",
  32553=>"000000110",
  32554=>"101001100",
  32555=>"001110111",
  32556=>"111110110",
  32557=>"000000000",
  32558=>"111111000",
  32559=>"101111110",
  32560=>"110001110",
  32561=>"011111001",
  32562=>"000010010",
  32563=>"101000000",
  32564=>"001001101",
  32565=>"110010100",
  32566=>"101100111",
  32567=>"010010011",
  32568=>"010011011",
  32569=>"111110100",
  32570=>"000101111",
  32571=>"001011110",
  32572=>"111001111",
  32573=>"010110101",
  32574=>"100101110",
  32575=>"101010011",
  32576=>"111010110",
  32577=>"000101010",
  32578=>"100001000",
  32579=>"100011100",
  32580=>"001000110",
  32581=>"100001101",
  32582=>"001111111",
  32583=>"010110110",
  32584=>"100010000",
  32585=>"111110000",
  32586=>"011101110",
  32587=>"101000010",
  32588=>"100001011",
  32589=>"111111011",
  32590=>"111101110",
  32591=>"101011101",
  32592=>"111110101",
  32593=>"110001000",
  32594=>"000100010",
  32595=>"111101001",
  32596=>"100111111",
  32597=>"110000001",
  32598=>"010010101",
  32599=>"110101111",
  32600=>"100100100",
  32601=>"101111100",
  32602=>"101010110",
  32603=>"111000110",
  32604=>"100011011",
  32605=>"101110000",
  32606=>"001110101",
  32607=>"111010001",
  32608=>"001011001",
  32609=>"000010000",
  32610=>"000000100",
  32611=>"110101100",
  32612=>"001011011",
  32613=>"010100100",
  32614=>"001110111",
  32615=>"000111110",
  32616=>"101111101",
  32617=>"100100000",
  32618=>"111100001",
  32619=>"110000100",
  32620=>"110101101",
  32621=>"011111111",
  32622=>"100001101",
  32623=>"101010010",
  32624=>"101110100",
  32625=>"011000001",
  32626=>"110010110",
  32627=>"101110101",
  32628=>"000001000",
  32629=>"111011010",
  32630=>"100110110",
  32631=>"110110011",
  32632=>"001011001",
  32633=>"001010110",
  32634=>"100001000",
  32635=>"110111000",
  32636=>"000011101",
  32637=>"011110111",
  32638=>"011101000",
  32639=>"100101000",
  32640=>"100010001",
  32641=>"011100111",
  32642=>"110001000",
  32643=>"001100111",
  32644=>"011011101",
  32645=>"010110010",
  32646=>"011110000",
  32647=>"110001001",
  32648=>"101000100",
  32649=>"110011010",
  32650=>"000111101",
  32651=>"110100101",
  32652=>"011011100",
  32653=>"000110100",
  32654=>"010001000",
  32655=>"010000010",
  32656=>"100111110",
  32657=>"100110010",
  32658=>"011100011",
  32659=>"010000000",
  32660=>"010111110",
  32661=>"111001010",
  32662=>"111010100",
  32663=>"010111101",
  32664=>"011011011",
  32665=>"100100000",
  32666=>"100010010",
  32667=>"010010001",
  32668=>"000001101",
  32669=>"110100001",
  32670=>"010010101",
  32671=>"110010111",
  32672=>"111010000",
  32673=>"110001111",
  32674=>"101010100",
  32675=>"100101111",
  32676=>"111001111",
  32677=>"000110000",
  32678=>"101110001",
  32679=>"100000000",
  32680=>"111101001",
  32681=>"110000000",
  32682=>"000100011",
  32683=>"010111010",
  32684=>"010111100",
  32685=>"000011011",
  32686=>"110000001",
  32687=>"010100101",
  32688=>"000101100",
  32689=>"000001010",
  32690=>"001011001",
  32691=>"111101111",
  32692=>"011100111",
  32693=>"101100001",
  32694=>"000110100",
  32695=>"000010000",
  32696=>"110110001",
  32697=>"100000010",
  32698=>"000011010",
  32699=>"010100011",
  32700=>"010000111",
  32701=>"000001100",
  32702=>"111011111",
  32703=>"111100111",
  32704=>"001100000",
  32705=>"100100110",
  32706=>"000111000",
  32707=>"111010010",
  32708=>"011010010",
  32709=>"110010010",
  32710=>"000011101",
  32711=>"100000000",
  32712=>"101110100",
  32713=>"000100101",
  32714=>"001111011",
  32715=>"100100000",
  32716=>"111111110",
  32717=>"111110111",
  32718=>"101011110",
  32719=>"101010010",
  32720=>"000010100",
  32721=>"011101110",
  32722=>"000111010",
  32723=>"101110011",
  32724=>"110111000",
  32725=>"011100011",
  32726=>"101010001",
  32727=>"110001101",
  32728=>"110100100",
  32729=>"101100101",
  32730=>"111110101",
  32731=>"101111101",
  32732=>"101001011",
  32733=>"010010000",
  32734=>"101001110",
  32735=>"001101001",
  32736=>"001011010",
  32737=>"101111001",
  32738=>"100101101",
  32739=>"110011000",
  32740=>"000110000",
  32741=>"111101001",
  32742=>"111101111",
  32743=>"001100010",
  32744=>"111110001",
  32745=>"000001010",
  32746=>"110110010",
  32747=>"110101000",
  32748=>"001010011",
  32749=>"000101111",
  32750=>"111000001",
  32751=>"001111000",
  32752=>"100001111",
  32753=>"111111111",
  32754=>"001010101",
  32755=>"110001010",
  32756=>"111000101",
  32757=>"011011010",
  32758=>"011000001",
  32759=>"101110010",
  32760=>"011110000",
  32761=>"000101011",
  32762=>"110110001",
  32763=>"011110010",
  32764=>"101101101",
  32765=>"011011101",
  32766=>"010011010",
  32767=>"101001110",
  32768=>"111100111",
  32769=>"110001000",
  32770=>"110000100",
  32771=>"100000100",
  32772=>"000110101",
  32773=>"111101101",
  32774=>"000000100",
  32775=>"111011011",
  32776=>"111000000",
  32777=>"101101111",
  32778=>"000010110",
  32779=>"101001000",
  32780=>"101111111",
  32781=>"010011001",
  32782=>"000011001",
  32783=>"101000100",
  32784=>"010110110",
  32785=>"000100000",
  32786=>"100000001",
  32787=>"110001001",
  32788=>"111111101",
  32789=>"000111101",
  32790=>"110100000",
  32791=>"110101000",
  32792=>"011111001",
  32793=>"111010110",
  32794=>"010110100",
  32795=>"110010111",
  32796=>"110110101",
  32797=>"001010000",
  32798=>"000000000",
  32799=>"000001001",
  32800=>"000001010",
  32801=>"011001010",
  32802=>"010001111",
  32803=>"100110101",
  32804=>"001111001",
  32805=>"000011101",
  32806=>"010001110",
  32807=>"101101000",
  32808=>"110010101",
  32809=>"001001110",
  32810=>"001100001",
  32811=>"011001110",
  32812=>"100110011",
  32813=>"111111011",
  32814=>"010111101",
  32815=>"010011101",
  32816=>"011000110",
  32817=>"011001101",
  32818=>"011101110",
  32819=>"000110111",
  32820=>"111110101",
  32821=>"011110011",
  32822=>"100100001",
  32823=>"111010110",
  32824=>"010100110",
  32825=>"101100100",
  32826=>"000110101",
  32827=>"110110011",
  32828=>"010110101",
  32829=>"111010001",
  32830=>"010011111",
  32831=>"110100101",
  32832=>"110111111",
  32833=>"001101110",
  32834=>"001111100",
  32835=>"100110101",
  32836=>"111001010",
  32837=>"111011011",
  32838=>"110111111",
  32839=>"001100001",
  32840=>"011110010",
  32841=>"001000100",
  32842=>"011100110",
  32843=>"001000011",
  32844=>"101110111",
  32845=>"011111011",
  32846=>"001011011",
  32847=>"110000011",
  32848=>"011010101",
  32849=>"100011000",
  32850=>"100010101",
  32851=>"000010111",
  32852=>"110100010",
  32853=>"000000100",
  32854=>"100010111",
  32855=>"101000001",
  32856=>"000000011",
  32857=>"011010100",
  32858=>"001010111",
  32859=>"011111010",
  32860=>"000111111",
  32861=>"111101101",
  32862=>"000101100",
  32863=>"001101111",
  32864=>"110011111",
  32865=>"001011000",
  32866=>"110001101",
  32867=>"110001111",
  32868=>"100010110",
  32869=>"100110001",
  32870=>"011111100",
  32871=>"111000111",
  32872=>"011001101",
  32873=>"001011011",
  32874=>"000000101",
  32875=>"110110010",
  32876=>"011011111",
  32877=>"100011111",
  32878=>"011000101",
  32879=>"111010110",
  32880=>"110010100",
  32881=>"011001110",
  32882=>"110111011",
  32883=>"111001001",
  32884=>"111001001",
  32885=>"110110001",
  32886=>"111011010",
  32887=>"100001110",
  32888=>"110110010",
  32889=>"111000110",
  32890=>"110110011",
  32891=>"100000101",
  32892=>"001110001",
  32893=>"100110100",
  32894=>"011110110",
  32895=>"101110101",
  32896=>"110000101",
  32897=>"100101110",
  32898=>"111100001",
  32899=>"110101111",
  32900=>"011111011",
  32901=>"101000101",
  32902=>"011111011",
  32903=>"100100101",
  32904=>"001001001",
  32905=>"100101101",
  32906=>"111001000",
  32907=>"010101111",
  32908=>"010000001",
  32909=>"110011111",
  32910=>"010111011",
  32911=>"101101101",
  32912=>"111001000",
  32913=>"001010000",
  32914=>"110100101",
  32915=>"001010100",
  32916=>"110010111",
  32917=>"101100001",
  32918=>"011011000",
  32919=>"101010011",
  32920=>"111011101",
  32921=>"011001001",
  32922=>"111111111",
  32923=>"000000101",
  32924=>"010001001",
  32925=>"110000111",
  32926=>"111011101",
  32927=>"111100000",
  32928=>"100100100",
  32929=>"001111111",
  32930=>"110100000",
  32931=>"101000010",
  32932=>"011010001",
  32933=>"101010011",
  32934=>"010100011",
  32935=>"100000111",
  32936=>"100101110",
  32937=>"111101010",
  32938=>"001010111",
  32939=>"011111011",
  32940=>"101001001",
  32941=>"100010000",
  32942=>"000000101",
  32943=>"111110010",
  32944=>"111011010",
  32945=>"000101110",
  32946=>"011000101",
  32947=>"100010001",
  32948=>"001111111",
  32949=>"111010111",
  32950=>"001000000",
  32951=>"010010010",
  32952=>"001000100",
  32953=>"010001111",
  32954=>"011001011",
  32955=>"000100101",
  32956=>"100100000",
  32957=>"101001111",
  32958=>"011101001",
  32959=>"010000001",
  32960=>"000100011",
  32961=>"000000100",
  32962=>"101111100",
  32963=>"000101110",
  32964=>"101110010",
  32965=>"010111001",
  32966=>"111100010",
  32967=>"010001011",
  32968=>"001101000",
  32969=>"001101101",
  32970=>"100010111",
  32971=>"100100011",
  32972=>"111100010",
  32973=>"010011000",
  32974=>"010110001",
  32975=>"001001011",
  32976=>"001010010",
  32977=>"000000101",
  32978=>"010001111",
  32979=>"110110010",
  32980=>"110110001",
  32981=>"100011011",
  32982=>"000001010",
  32983=>"111010101",
  32984=>"100110111",
  32985=>"100010110",
  32986=>"101001100",
  32987=>"111001010",
  32988=>"100101010",
  32989=>"010001001",
  32990=>"101000101",
  32991=>"110011101",
  32992=>"101000101",
  32993=>"010010110",
  32994=>"111001000",
  32995=>"011101010",
  32996=>"111011110",
  32997=>"001110100",
  32998=>"111000101",
  32999=>"111100101",
  33000=>"001000001",
  33001=>"111000001",
  33002=>"000011011",
  33003=>"001000110",
  33004=>"111100111",
  33005=>"011000010",
  33006=>"111100001",
  33007=>"001110010",
  33008=>"111011000",
  33009=>"011011011",
  33010=>"111101101",
  33011=>"001100100",
  33012=>"000011101",
  33013=>"000110100",
  33014=>"100101001",
  33015=>"110001010",
  33016=>"000111010",
  33017=>"011111010",
  33018=>"100111000",
  33019=>"101000101",
  33020=>"010000011",
  33021=>"010011011",
  33022=>"111010011",
  33023=>"110010110",
  33024=>"101101001",
  33025=>"110110011",
  33026=>"011001000",
  33027=>"010010001",
  33028=>"110010101",
  33029=>"010110110",
  33030=>"001011000",
  33031=>"101100010",
  33032=>"001100000",
  33033=>"000111000",
  33034=>"100101111",
  33035=>"010011010",
  33036=>"101001001",
  33037=>"011110110",
  33038=>"100001111",
  33039=>"001100001",
  33040=>"011001110",
  33041=>"011101100",
  33042=>"110100111",
  33043=>"101011011",
  33044=>"100110100",
  33045=>"000110110",
  33046=>"100011010",
  33047=>"101010111",
  33048=>"000100010",
  33049=>"111101011",
  33050=>"111001111",
  33051=>"101111100",
  33052=>"010001001",
  33053=>"000100001",
  33054=>"111011111",
  33055=>"000101111",
  33056=>"011010110",
  33057=>"001011100",
  33058=>"111000111",
  33059=>"000101111",
  33060=>"101011001",
  33061=>"101011001",
  33062=>"000101100",
  33063=>"111110101",
  33064=>"100000000",
  33065=>"110111010",
  33066=>"100000110",
  33067=>"110101110",
  33068=>"111010000",
  33069=>"101000111",
  33070=>"100001011",
  33071=>"111110011",
  33072=>"110110111",
  33073=>"000001001",
  33074=>"001001110",
  33075=>"000010010",
  33076=>"001110100",
  33077=>"000011000",
  33078=>"110010010",
  33079=>"111110000",
  33080=>"110011111",
  33081=>"001101110",
  33082=>"100110111",
  33083=>"001010101",
  33084=>"101000011",
  33085=>"100001000",
  33086=>"010000010",
  33087=>"000111100",
  33088=>"111010101",
  33089=>"111111100",
  33090=>"001001101",
  33091=>"110111000",
  33092=>"101000001",
  33093=>"000010101",
  33094=>"110001101",
  33095=>"000101010",
  33096=>"101101101",
  33097=>"010010010",
  33098=>"101010011",
  33099=>"100000110",
  33100=>"001100011",
  33101=>"011110000",
  33102=>"100001101",
  33103=>"010101010",
  33104=>"001000100",
  33105=>"010000010",
  33106=>"100000111",
  33107=>"010100001",
  33108=>"101100011",
  33109=>"110110001",
  33110=>"110000101",
  33111=>"011010001",
  33112=>"000010000",
  33113=>"100110001",
  33114=>"101110011",
  33115=>"010001110",
  33116=>"111011101",
  33117=>"110100111",
  33118=>"100110110",
  33119=>"101111110",
  33120=>"111111101",
  33121=>"001000101",
  33122=>"001001001",
  33123=>"111000101",
  33124=>"111100011",
  33125=>"001001110",
  33126=>"001101011",
  33127=>"111110111",
  33128=>"010101100",
  33129=>"100100101",
  33130=>"010111001",
  33131=>"011101101",
  33132=>"100110111",
  33133=>"000010101",
  33134=>"000100110",
  33135=>"111001110",
  33136=>"110100011",
  33137=>"001101000",
  33138=>"000001111",
  33139=>"101101100",
  33140=>"001101100",
  33141=>"101101110",
  33142=>"010000001",
  33143=>"111100000",
  33144=>"011001100",
  33145=>"011101101",
  33146=>"111101110",
  33147=>"100000101",
  33148=>"101111101",
  33149=>"110010001",
  33150=>"101011010",
  33151=>"110000111",
  33152=>"100000001",
  33153=>"001001110",
  33154=>"111101011",
  33155=>"110100110",
  33156=>"111011111",
  33157=>"110100110",
  33158=>"110111110",
  33159=>"110001111",
  33160=>"011010111",
  33161=>"000110111",
  33162=>"000100100",
  33163=>"110000001",
  33164=>"010100010",
  33165=>"010100111",
  33166=>"000000011",
  33167=>"001100011",
  33168=>"101111111",
  33169=>"010000000",
  33170=>"101010111",
  33171=>"111001110",
  33172=>"011110011",
  33173=>"001001000",
  33174=>"001011011",
  33175=>"011010100",
  33176=>"010000101",
  33177=>"100011001",
  33178=>"111011001",
  33179=>"010011000",
  33180=>"001100100",
  33181=>"010001000",
  33182=>"001010000",
  33183=>"011001011",
  33184=>"010000101",
  33185=>"001100001",
  33186=>"000110010",
  33187=>"100000000",
  33188=>"011100110",
  33189=>"100100000",
  33190=>"010110111",
  33191=>"001110111",
  33192=>"000101010",
  33193=>"111000011",
  33194=>"000001111",
  33195=>"000100101",
  33196=>"001101011",
  33197=>"101010000",
  33198=>"010010101",
  33199=>"000110111",
  33200=>"010000110",
  33201=>"011110100",
  33202=>"011000000",
  33203=>"000010011",
  33204=>"011110011",
  33205=>"100010110",
  33206=>"000011101",
  33207=>"001111100",
  33208=>"010000010",
  33209=>"010110110",
  33210=>"100001001",
  33211=>"000100100",
  33212=>"011010000",
  33213=>"111100000",
  33214=>"000000001",
  33215=>"111000000",
  33216=>"011000101",
  33217=>"100001110",
  33218=>"111111101",
  33219=>"010010110",
  33220=>"010011101",
  33221=>"111101100",
  33222=>"010000111",
  33223=>"001010111",
  33224=>"110010000",
  33225=>"101100101",
  33226=>"111111111",
  33227=>"100001000",
  33228=>"101001110",
  33229=>"111011110",
  33230=>"111010100",
  33231=>"010001001",
  33232=>"011010100",
  33233=>"110110010",
  33234=>"001000111",
  33235=>"111111110",
  33236=>"110100010",
  33237=>"110000100",
  33238=>"100001111",
  33239=>"000000000",
  33240=>"100001000",
  33241=>"101011110",
  33242=>"111010101",
  33243=>"111001100",
  33244=>"000000000",
  33245=>"110111111",
  33246=>"011110010",
  33247=>"000011111",
  33248=>"000101011",
  33249=>"011110001",
  33250=>"111010110",
  33251=>"011000011",
  33252=>"000001010",
  33253=>"000000001",
  33254=>"101000110",
  33255=>"011101011",
  33256=>"111000100",
  33257=>"011001000",
  33258=>"001111001",
  33259=>"111011000",
  33260=>"000010001",
  33261=>"000111111",
  33262=>"000001101",
  33263=>"100110000",
  33264=>"000111010",
  33265=>"011111111",
  33266=>"110111100",
  33267=>"011000100",
  33268=>"001011100",
  33269=>"100100111",
  33270=>"101000100",
  33271=>"110101111",
  33272=>"101011110",
  33273=>"111101100",
  33274=>"000110011",
  33275=>"010100110",
  33276=>"010001001",
  33277=>"100010100",
  33278=>"100011011",
  33279=>"110010100",
  33280=>"110101111",
  33281=>"101101110",
  33282=>"100100100",
  33283=>"101110001",
  33284=>"100000000",
  33285=>"100010001",
  33286=>"100010110",
  33287=>"011110000",
  33288=>"001101111",
  33289=>"011111001",
  33290=>"111111100",
  33291=>"000111000",
  33292=>"011111101",
  33293=>"111000011",
  33294=>"010010100",
  33295=>"111100111",
  33296=>"000101111",
  33297=>"111000010",
  33298=>"110010110",
  33299=>"110111111",
  33300=>"001010101",
  33301=>"000100100",
  33302=>"001001011",
  33303=>"100110001",
  33304=>"010001101",
  33305=>"101001101",
  33306=>"010111000",
  33307=>"011001011",
  33308=>"101101000",
  33309=>"111001100",
  33310=>"000100010",
  33311=>"111010000",
  33312=>"000000100",
  33313=>"010011111",
  33314=>"110000011",
  33315=>"000101011",
  33316=>"110001101",
  33317=>"000001110",
  33318=>"110100111",
  33319=>"111111100",
  33320=>"101101101",
  33321=>"110010000",
  33322=>"100111010",
  33323=>"111001100",
  33324=>"110110110",
  33325=>"000001001",
  33326=>"010101000",
  33327=>"000011100",
  33328=>"110011111",
  33329=>"110001111",
  33330=>"000100001",
  33331=>"110011010",
  33332=>"111001011",
  33333=>"000111010",
  33334=>"000100001",
  33335=>"101001110",
  33336=>"101000100",
  33337=>"000100001",
  33338=>"001000001",
  33339=>"000010000",
  33340=>"111001101",
  33341=>"011100110",
  33342=>"001111000",
  33343=>"101001111",
  33344=>"100101011",
  33345=>"111010101",
  33346=>"111010011",
  33347=>"110100110",
  33348=>"110111111",
  33349=>"010000010",
  33350=>"110001000",
  33351=>"010111000",
  33352=>"111010101",
  33353=>"100000011",
  33354=>"001111110",
  33355=>"110101011",
  33356=>"010101010",
  33357=>"001110111",
  33358=>"111110001",
  33359=>"001110011",
  33360=>"010101001",
  33361=>"111001101",
  33362=>"010111001",
  33363=>"111010101",
  33364=>"010000101",
  33365=>"001000010",
  33366=>"011001111",
  33367=>"001010011",
  33368=>"000100111",
  33369=>"101001100",
  33370=>"001000001",
  33371=>"111111111",
  33372=>"100100000",
  33373=>"000010010",
  33374=>"001010100",
  33375=>"011111010",
  33376=>"001101011",
  33377=>"101001000",
  33378=>"101101000",
  33379=>"100110001",
  33380=>"111101100",
  33381=>"111111010",
  33382=>"101010001",
  33383=>"000001010",
  33384=>"110100011",
  33385=>"100011011",
  33386=>"110011100",
  33387=>"101101101",
  33388=>"100101011",
  33389=>"100110011",
  33390=>"011010011",
  33391=>"110100001",
  33392=>"100000011",
  33393=>"101000001",
  33394=>"110010101",
  33395=>"001100100",
  33396=>"110100011",
  33397=>"000001100",
  33398=>"011110100",
  33399=>"001101101",
  33400=>"010110101",
  33401=>"110010110",
  33402=>"011111011",
  33403=>"101111000",
  33404=>"000001001",
  33405=>"001000100",
  33406=>"100100000",
  33407=>"111111101",
  33408=>"110101110",
  33409=>"100101110",
  33410=>"000000111",
  33411=>"100100110",
  33412=>"011111111",
  33413=>"101100010",
  33414=>"111001000",
  33415=>"111111000",
  33416=>"011001100",
  33417=>"100010000",
  33418=>"110000000",
  33419=>"101110010",
  33420=>"000001000",
  33421=>"101000011",
  33422=>"111110100",
  33423=>"100000011",
  33424=>"100001110",
  33425=>"101110010",
  33426=>"111100101",
  33427=>"111111110",
  33428=>"000101111",
  33429=>"110101000",
  33430=>"010111101",
  33431=>"001010000",
  33432=>"101010100",
  33433=>"111110010",
  33434=>"000011110",
  33435=>"111000011",
  33436=>"010101000",
  33437=>"000001111",
  33438=>"000101010",
  33439=>"110101110",
  33440=>"111001010",
  33441=>"010100100",
  33442=>"111001000",
  33443=>"111100001",
  33444=>"111001011",
  33445=>"101101001",
  33446=>"110101010",
  33447=>"100111101",
  33448=>"000000000",
  33449=>"111101111",
  33450=>"100001001",
  33451=>"011000100",
  33452=>"011100010",
  33453=>"011101110",
  33454=>"100000000",
  33455=>"001100110",
  33456=>"100000101",
  33457=>"110100011",
  33458=>"010110111",
  33459=>"100001111",
  33460=>"111001111",
  33461=>"000010010",
  33462=>"101011100",
  33463=>"011010100",
  33464=>"110000100",
  33465=>"010001011",
  33466=>"001010110",
  33467=>"010110110",
  33468=>"011001100",
  33469=>"010011110",
  33470=>"010010001",
  33471=>"001011101",
  33472=>"110001010",
  33473=>"100101011",
  33474=>"000001100",
  33475=>"010100101",
  33476=>"100011011",
  33477=>"000111010",
  33478=>"100100000",
  33479=>"001010010",
  33480=>"100100001",
  33481=>"001011110",
  33482=>"110001101",
  33483=>"111011011",
  33484=>"101000101",
  33485=>"010000001",
  33486=>"111111011",
  33487=>"111100110",
  33488=>"100110010",
  33489=>"110010000",
  33490=>"111001000",
  33491=>"001000101",
  33492=>"001111100",
  33493=>"101101110",
  33494=>"110100011",
  33495=>"111110000",
  33496=>"000111000",
  33497=>"101111111",
  33498=>"101101010",
  33499=>"111111111",
  33500=>"010100000",
  33501=>"111110000",
  33502=>"001111100",
  33503=>"001010000",
  33504=>"010111110",
  33505=>"101111101",
  33506=>"010101000",
  33507=>"001100000",
  33508=>"101111111",
  33509=>"100110000",
  33510=>"100111110",
  33511=>"000111000",
  33512=>"001110011",
  33513=>"011100100",
  33514=>"001001111",
  33515=>"111111111",
  33516=>"111011001",
  33517=>"000000011",
  33518=>"000010000",
  33519=>"111100111",
  33520=>"110010011",
  33521=>"101000001",
  33522=>"001010111",
  33523=>"110001110",
  33524=>"100110010",
  33525=>"011100010",
  33526=>"101011100",
  33527=>"001100111",
  33528=>"101101101",
  33529=>"110110001",
  33530=>"010100111",
  33531=>"110100000",
  33532=>"000100011",
  33533=>"100011100",
  33534=>"011101011",
  33535=>"100100001",
  33536=>"010111000",
  33537=>"100110100",
  33538=>"100100100",
  33539=>"000001100",
  33540=>"001000100",
  33541=>"111110001",
  33542=>"000101011",
  33543=>"010010100",
  33544=>"011011111",
  33545=>"000011000",
  33546=>"011111101",
  33547=>"001101010",
  33548=>"100001101",
  33549=>"110111011",
  33550=>"101010100",
  33551=>"010010111",
  33552=>"101001111",
  33553=>"001010110",
  33554=>"100010001",
  33555=>"011110101",
  33556=>"011101000",
  33557=>"100101001",
  33558=>"110110111",
  33559=>"100111000",
  33560=>"111001101",
  33561=>"110000010",
  33562=>"110110101",
  33563=>"001100000",
  33564=>"011110100",
  33565=>"010001111",
  33566=>"101010010",
  33567=>"011011010",
  33568=>"100011010",
  33569=>"001100110",
  33570=>"011110001",
  33571=>"100010101",
  33572=>"001001011",
  33573=>"100100011",
  33574=>"010010000",
  33575=>"011101110",
  33576=>"000011011",
  33577=>"111000100",
  33578=>"000111000",
  33579=>"101011111",
  33580=>"011011011",
  33581=>"101010001",
  33582=>"010010110",
  33583=>"111110111",
  33584=>"100101001",
  33585=>"110101111",
  33586=>"000010011",
  33587=>"011110011",
  33588=>"000110100",
  33589=>"111110001",
  33590=>"000100100",
  33591=>"100001101",
  33592=>"011011001",
  33593=>"000001000",
  33594=>"101111110",
  33595=>"110010001",
  33596=>"100111011",
  33597=>"100000000",
  33598=>"100101101",
  33599=>"001110000",
  33600=>"100001000",
  33601=>"011101101",
  33602=>"001101101",
  33603=>"000110111",
  33604=>"001010001",
  33605=>"111001000",
  33606=>"000110000",
  33607=>"010010001",
  33608=>"011011001",
  33609=>"101001000",
  33610=>"100001010",
  33611=>"011000001",
  33612=>"101100000",
  33613=>"011100000",
  33614=>"001110010",
  33615=>"101110110",
  33616=>"000001110",
  33617=>"111011001",
  33618=>"111000100",
  33619=>"001001100",
  33620=>"100100011",
  33621=>"011000110",
  33622=>"001001110",
  33623=>"000101101",
  33624=>"101000001",
  33625=>"111100111",
  33626=>"111001111",
  33627=>"111110101",
  33628=>"111011100",
  33629=>"010001101",
  33630=>"001010000",
  33631=>"000001010",
  33632=>"010000000",
  33633=>"101010010",
  33634=>"100111000",
  33635=>"100001001",
  33636=>"110100111",
  33637=>"011001011",
  33638=>"001010011",
  33639=>"001011011",
  33640=>"011010111",
  33641=>"001101100",
  33642=>"110001100",
  33643=>"001010111",
  33644=>"001111000",
  33645=>"001110001",
  33646=>"111000111",
  33647=>"011100111",
  33648=>"100100000",
  33649=>"010100010",
  33650=>"000001011",
  33651=>"011010001",
  33652=>"010000100",
  33653=>"001000101",
  33654=>"011111000",
  33655=>"111101010",
  33656=>"110010000",
  33657=>"010011011",
  33658=>"000011001",
  33659=>"101000100",
  33660=>"010010111",
  33661=>"100001011",
  33662=>"010011101",
  33663=>"001110111",
  33664=>"111101101",
  33665=>"010010110",
  33666=>"000001100",
  33667=>"010001100",
  33668=>"110000110",
  33669=>"011001111",
  33670=>"011000111",
  33671=>"001011100",
  33672=>"011000000",
  33673=>"110010001",
  33674=>"000010101",
  33675=>"101101101",
  33676=>"010100100",
  33677=>"100011011",
  33678=>"111110000",
  33679=>"001100010",
  33680=>"010001100",
  33681=>"111011010",
  33682=>"000101100",
  33683=>"011011101",
  33684=>"011101001",
  33685=>"101110010",
  33686=>"001010010",
  33687=>"110110110",
  33688=>"001010110",
  33689=>"001010000",
  33690=>"111101111",
  33691=>"010010010",
  33692=>"010011000",
  33693=>"100101111",
  33694=>"011111101",
  33695=>"011111100",
  33696=>"101100011",
  33697=>"000010100",
  33698=>"101011101",
  33699=>"111010110",
  33700=>"000100000",
  33701=>"101111011",
  33702=>"000100000",
  33703=>"100101111",
  33704=>"101100001",
  33705=>"111110111",
  33706=>"111100010",
  33707=>"110000011",
  33708=>"111001000",
  33709=>"010101101",
  33710=>"110100011",
  33711=>"100010100",
  33712=>"110010011",
  33713=>"100001011",
  33714=>"101011001",
  33715=>"001110110",
  33716=>"000011000",
  33717=>"111111011",
  33718=>"001111101",
  33719=>"000010010",
  33720=>"111000110",
  33721=>"100000100",
  33722=>"010111000",
  33723=>"110011100",
  33724=>"000010111",
  33725=>"110110011",
  33726=>"111001001",
  33727=>"001001100",
  33728=>"000011011",
  33729=>"000001111",
  33730=>"111100100",
  33731=>"000101101",
  33732=>"000001110",
  33733=>"011001101",
  33734=>"001101111",
  33735=>"110011110",
  33736=>"000100000",
  33737=>"010010101",
  33738=>"011101011",
  33739=>"001000111",
  33740=>"111101110",
  33741=>"101100100",
  33742=>"000001101",
  33743=>"011100101",
  33744=>"010110001",
  33745=>"010101010",
  33746=>"110101000",
  33747=>"101001011",
  33748=>"001101000",
  33749=>"001000110",
  33750=>"110000101",
  33751=>"101001111",
  33752=>"010011100",
  33753=>"001111110",
  33754=>"010110010",
  33755=>"101101011",
  33756=>"110110101",
  33757=>"101101000",
  33758=>"000100011",
  33759=>"100011010",
  33760=>"100101001",
  33761=>"101100111",
  33762=>"011111101",
  33763=>"010001110",
  33764=>"110010000",
  33765=>"111110101",
  33766=>"001001011",
  33767=>"011011100",
  33768=>"001000101",
  33769=>"000111110",
  33770=>"110011001",
  33771=>"011011001",
  33772=>"000001110",
  33773=>"100111101",
  33774=>"110110011",
  33775=>"010101011",
  33776=>"000101011",
  33777=>"011100100",
  33778=>"010100001",
  33779=>"100111110",
  33780=>"111010101",
  33781=>"000001101",
  33782=>"010100010",
  33783=>"111000000",
  33784=>"101011110",
  33785=>"101000001",
  33786=>"101000101",
  33787=>"011000010",
  33788=>"110001100",
  33789=>"010110011",
  33790=>"110101001",
  33791=>"001110010",
  33792=>"111011010",
  33793=>"101110101",
  33794=>"011011011",
  33795=>"011110010",
  33796=>"000000110",
  33797=>"001100010",
  33798=>"011100110",
  33799=>"100010011",
  33800=>"000100001",
  33801=>"111111011",
  33802=>"101000000",
  33803=>"100111011",
  33804=>"111000010",
  33805=>"101111011",
  33806=>"010100000",
  33807=>"101001101",
  33808=>"001001010",
  33809=>"101110101",
  33810=>"010101011",
  33811=>"000111100",
  33812=>"011101000",
  33813=>"111111111",
  33814=>"110011100",
  33815=>"101101111",
  33816=>"000011100",
  33817=>"001110000",
  33818=>"101000101",
  33819=>"101011110",
  33820=>"011111011",
  33821=>"110110111",
  33822=>"011101111",
  33823=>"010000111",
  33824=>"101111110",
  33825=>"010011011",
  33826=>"100100010",
  33827=>"010000100",
  33828=>"011000100",
  33829=>"001100110",
  33830=>"101001010",
  33831=>"100110000",
  33832=>"100101101",
  33833=>"110011000",
  33834=>"101110001",
  33835=>"010111111",
  33836=>"001101001",
  33837=>"011010100",
  33838=>"101111010",
  33839=>"001000101",
  33840=>"010110111",
  33841=>"110111101",
  33842=>"011011010",
  33843=>"111010111",
  33844=>"101000101",
  33845=>"110011000",
  33846=>"110001111",
  33847=>"101110001",
  33848=>"111101101",
  33849=>"111110110",
  33850=>"001001011",
  33851=>"000011101",
  33852=>"001111010",
  33853=>"100100111",
  33854=>"010000000",
  33855=>"000111101",
  33856=>"110000101",
  33857=>"011000111",
  33858=>"000010111",
  33859=>"010001000",
  33860=>"110110010",
  33861=>"110111100",
  33862=>"110101100",
  33863=>"111101101",
  33864=>"100001011",
  33865=>"000100001",
  33866=>"010001000",
  33867=>"100101111",
  33868=>"000011001",
  33869=>"011101110",
  33870=>"001101111",
  33871=>"100011010",
  33872=>"101111100",
  33873=>"000110000",
  33874=>"101110011",
  33875=>"111011010",
  33876=>"100000001",
  33877=>"000010011",
  33878=>"010011010",
  33879=>"011011110",
  33880=>"000100110",
  33881=>"001101000",
  33882=>"101000110",
  33883=>"100100101",
  33884=>"000001001",
  33885=>"010010010",
  33886=>"111100101",
  33887=>"001100011",
  33888=>"110110001",
  33889=>"001011010",
  33890=>"010110101",
  33891=>"110110001",
  33892=>"110100010",
  33893=>"011010000",
  33894=>"000110111",
  33895=>"100101111",
  33896=>"001000100",
  33897=>"001001101",
  33898=>"110011011",
  33899=>"011011110",
  33900=>"011010100",
  33901=>"101111100",
  33902=>"011000101",
  33903=>"011100100",
  33904=>"101011100",
  33905=>"101001101",
  33906=>"000010010",
  33907=>"000110000",
  33908=>"111011010",
  33909=>"111101101",
  33910=>"110110110",
  33911=>"010101001",
  33912=>"000000011",
  33913=>"011100110",
  33914=>"001010011",
  33915=>"010111110",
  33916=>"111010011",
  33917=>"100000100",
  33918=>"011101010",
  33919=>"101100100",
  33920=>"011001000",
  33921=>"001110000",
  33922=>"100001010",
  33923=>"001110001",
  33924=>"110000011",
  33925=>"000011110",
  33926=>"111100010",
  33927=>"000100100",
  33928=>"010010100",
  33929=>"100010000",
  33930=>"010111011",
  33931=>"011100100",
  33932=>"010010010",
  33933=>"000100010",
  33934=>"100011101",
  33935=>"000000011",
  33936=>"110101011",
  33937=>"111110111",
  33938=>"110010101",
  33939=>"011111011",
  33940=>"000110101",
  33941=>"101111110",
  33942=>"000000101",
  33943=>"010110101",
  33944=>"001001000",
  33945=>"000100011",
  33946=>"000101101",
  33947=>"010001001",
  33948=>"000111100",
  33949=>"010110100",
  33950=>"000011111",
  33951=>"110011101",
  33952=>"100001001",
  33953=>"000111000",
  33954=>"111101011",
  33955=>"000110101",
  33956=>"101011111",
  33957=>"111110111",
  33958=>"110000011",
  33959=>"100001001",
  33960=>"100001000",
  33961=>"100010110",
  33962=>"001010000",
  33963=>"001101100",
  33964=>"111011001",
  33965=>"010011010",
  33966=>"011111001",
  33967=>"000011111",
  33968=>"101011010",
  33969=>"000100000",
  33970=>"011001001",
  33971=>"000001000",
  33972=>"010101100",
  33973=>"000011011",
  33974=>"010101110",
  33975=>"101001111",
  33976=>"000011100",
  33977=>"001001010",
  33978=>"001110010",
  33979=>"100110010",
  33980=>"100101110",
  33981=>"101111101",
  33982=>"101001001",
  33983=>"100111110",
  33984=>"000000011",
  33985=>"101000001",
  33986=>"101000011",
  33987=>"110011000",
  33988=>"100000011",
  33989=>"111110111",
  33990=>"111110010",
  33991=>"000011110",
  33992=>"010110001",
  33993=>"101101111",
  33994=>"000010100",
  33995=>"011111101",
  33996=>"110110000",
  33997=>"000101110",
  33998=>"001110101",
  33999=>"110010101",
  34000=>"010111101",
  34001=>"101111010",
  34002=>"000010111",
  34003=>"100101111",
  34004=>"111100001",
  34005=>"100111100",
  34006=>"010101010",
  34007=>"010100110",
  34008=>"111110000",
  34009=>"100011100",
  34010=>"110111100",
  34011=>"110010111",
  34012=>"010011001",
  34013=>"110001011",
  34014=>"101000001",
  34015=>"100100111",
  34016=>"010011111",
  34017=>"011110000",
  34018=>"111101010",
  34019=>"001011111",
  34020=>"010101111",
  34021=>"101100011",
  34022=>"010001011",
  34023=>"111100100",
  34024=>"000000001",
  34025=>"110010101",
  34026=>"000001011",
  34027=>"111110010",
  34028=>"111000110",
  34029=>"000011111",
  34030=>"101000101",
  34031=>"101010001",
  34032=>"100101000",
  34033=>"010110111",
  34034=>"111110000",
  34035=>"000010110",
  34036=>"011111110",
  34037=>"000110101",
  34038=>"100001011",
  34039=>"011110100",
  34040=>"001100100",
  34041=>"110110010",
  34042=>"101110100",
  34043=>"010010011",
  34044=>"001100010",
  34045=>"100111111",
  34046=>"101111011",
  34047=>"100010000",
  34048=>"110001000",
  34049=>"001110111",
  34050=>"010000010",
  34051=>"101001101",
  34052=>"010111010",
  34053=>"110001010",
  34054=>"110011110",
  34055=>"001011001",
  34056=>"100000000",
  34057=>"011111010",
  34058=>"110001100",
  34059=>"101001111",
  34060=>"101001000",
  34061=>"101011011",
  34062=>"011100011",
  34063=>"000110111",
  34064=>"001101101",
  34065=>"000110001",
  34066=>"010001010",
  34067=>"110011110",
  34068=>"110100011",
  34069=>"010000100",
  34070=>"010101001",
  34071=>"000010110",
  34072=>"101111010",
  34073=>"011100111",
  34074=>"111001101",
  34075=>"100111111",
  34076=>"011010000",
  34077=>"110001111",
  34078=>"100110010",
  34079=>"000010100",
  34080=>"011100111",
  34081=>"110110100",
  34082=>"011000001",
  34083=>"000111100",
  34084=>"011110001",
  34085=>"000110100",
  34086=>"100111100",
  34087=>"100100101",
  34088=>"000011000",
  34089=>"010110100",
  34090=>"001010110",
  34091=>"100101000",
  34092=>"111001000",
  34093=>"100011100",
  34094=>"100000111",
  34095=>"001101001",
  34096=>"000100010",
  34097=>"101001001",
  34098=>"101011011",
  34099=>"100101110",
  34100=>"001000100",
  34101=>"111111010",
  34102=>"000000011",
  34103=>"111001101",
  34104=>"110110001",
  34105=>"101011011",
  34106=>"100000000",
  34107=>"101110100",
  34108=>"100111001",
  34109=>"100100001",
  34110=>"011100011",
  34111=>"111111100",
  34112=>"111101001",
  34113=>"100010000",
  34114=>"010001011",
  34115=>"001110011",
  34116=>"011000000",
  34117=>"110100100",
  34118=>"111010010",
  34119=>"111101010",
  34120=>"111101001",
  34121=>"010001010",
  34122=>"100010100",
  34123=>"011000001",
  34124=>"001111100",
  34125=>"111000001",
  34126=>"000100010",
  34127=>"101101101",
  34128=>"011010011",
  34129=>"000011001",
  34130=>"000001100",
  34131=>"010010001",
  34132=>"011001100",
  34133=>"010000110",
  34134=>"101100100",
  34135=>"100010000",
  34136=>"101000111",
  34137=>"110001101",
  34138=>"111111010",
  34139=>"001101010",
  34140=>"101011111",
  34141=>"011101101",
  34142=>"011100001",
  34143=>"011010001",
  34144=>"111111000",
  34145=>"010100010",
  34146=>"010011001",
  34147=>"001110111",
  34148=>"010100010",
  34149=>"001110110",
  34150=>"100001100",
  34151=>"011001011",
  34152=>"001101010",
  34153=>"110010010",
  34154=>"000010111",
  34155=>"100111000",
  34156=>"110001010",
  34157=>"010101010",
  34158=>"101011111",
  34159=>"011000001",
  34160=>"010100101",
  34161=>"010000000",
  34162=>"011100111",
  34163=>"100101001",
  34164=>"010101000",
  34165=>"011101110",
  34166=>"001101100",
  34167=>"000110110",
  34168=>"011100100",
  34169=>"110011110",
  34170=>"111101010",
  34171=>"000011100",
  34172=>"101100000",
  34173=>"111110000",
  34174=>"100010010",
  34175=>"010101111",
  34176=>"010110001",
  34177=>"100101100",
  34178=>"111111001",
  34179=>"101111100",
  34180=>"100011111",
  34181=>"110001110",
  34182=>"110010100",
  34183=>"000001111",
  34184=>"101100101",
  34185=>"101010000",
  34186=>"101110001",
  34187=>"100011011",
  34188=>"010000111",
  34189=>"001110011",
  34190=>"011111001",
  34191=>"101110010",
  34192=>"100010001",
  34193=>"000000110",
  34194=>"100111010",
  34195=>"111110010",
  34196=>"010001100",
  34197=>"001001111",
  34198=>"000110010",
  34199=>"011001000",
  34200=>"100111001",
  34201=>"001000000",
  34202=>"101101101",
  34203=>"100100110",
  34204=>"010000101",
  34205=>"010000001",
  34206=>"111110110",
  34207=>"000001001",
  34208=>"100111010",
  34209=>"011101000",
  34210=>"110000000",
  34211=>"010000001",
  34212=>"001110001",
  34213=>"001011011",
  34214=>"010010011",
  34215=>"101000011",
  34216=>"110110100",
  34217=>"000000000",
  34218=>"100011000",
  34219=>"100100100",
  34220=>"000111101",
  34221=>"111011100",
  34222=>"011010100",
  34223=>"101100000",
  34224=>"101000000",
  34225=>"001100001",
  34226=>"101100011",
  34227=>"001010100",
  34228=>"111111000",
  34229=>"011000010",
  34230=>"000100101",
  34231=>"001010111",
  34232=>"101000110",
  34233=>"110011011",
  34234=>"010110100",
  34235=>"001011010",
  34236=>"111110110",
  34237=>"110100111",
  34238=>"010110101",
  34239=>"111111011",
  34240=>"000110111",
  34241=>"101111111",
  34242=>"011101100",
  34243=>"101010110",
  34244=>"001100010",
  34245=>"000101000",
  34246=>"000000000",
  34247=>"001010011",
  34248=>"010100111",
  34249=>"000000010",
  34250=>"111000110",
  34251=>"011001001",
  34252=>"000111000",
  34253=>"111001001",
  34254=>"100100000",
  34255=>"111011110",
  34256=>"101111110",
  34257=>"001101100",
  34258=>"100000000",
  34259=>"100010110",
  34260=>"110100010",
  34261=>"001011101",
  34262=>"001101111",
  34263=>"000000000",
  34264=>"111001110",
  34265=>"000010101",
  34266=>"100000011",
  34267=>"010111110",
  34268=>"111110001",
  34269=>"101010111",
  34270=>"100101110",
  34271=>"000010111",
  34272=>"111111011",
  34273=>"111001010",
  34274=>"000000101",
  34275=>"111111111",
  34276=>"100011011",
  34277=>"100000010",
  34278=>"000000000",
  34279=>"110111001",
  34280=>"101001000",
  34281=>"011100100",
  34282=>"100000111",
  34283=>"101110010",
  34284=>"001010000",
  34285=>"000011100",
  34286=>"001010011",
  34287=>"001011110",
  34288=>"101100010",
  34289=>"000010010",
  34290=>"011110101",
  34291=>"111000100",
  34292=>"001010000",
  34293=>"110011011",
  34294=>"101111110",
  34295=>"010110111",
  34296=>"000000110",
  34297=>"011001111",
  34298=>"001110010",
  34299=>"000001010",
  34300=>"001011010",
  34301=>"010001101",
  34302=>"000001110",
  34303=>"110100111",
  34304=>"101100011",
  34305=>"101101110",
  34306=>"110101100",
  34307=>"000000001",
  34308=>"100000110",
  34309=>"110010011",
  34310=>"001011110",
  34311=>"101110111",
  34312=>"110000100",
  34313=>"111011001",
  34314=>"011110101",
  34315=>"101000111",
  34316=>"010001110",
  34317=>"111001010",
  34318=>"011000111",
  34319=>"010011000",
  34320=>"001010110",
  34321=>"000100100",
  34322=>"000111011",
  34323=>"001001111",
  34324=>"010100111",
  34325=>"110111111",
  34326=>"011110100",
  34327=>"100001101",
  34328=>"011010011",
  34329=>"100100100",
  34330=>"100010011",
  34331=>"110100011",
  34332=>"101110111",
  34333=>"000100101",
  34334=>"011111000",
  34335=>"001000110",
  34336=>"101010000",
  34337=>"111110111",
  34338=>"010001001",
  34339=>"010010010",
  34340=>"000110001",
  34341=>"101001111",
  34342=>"001101011",
  34343=>"110100110",
  34344=>"110101110",
  34345=>"101001100",
  34346=>"110111111",
  34347=>"101100001",
  34348=>"010001000",
  34349=>"000000010",
  34350=>"000000101",
  34351=>"001101010",
  34352=>"101101010",
  34353=>"101110000",
  34354=>"101111001",
  34355=>"101001111",
  34356=>"101101101",
  34357=>"100010100",
  34358=>"000101111",
  34359=>"001010100",
  34360=>"100100000",
  34361=>"111111010",
  34362=>"001111111",
  34363=>"100101001",
  34364=>"111000100",
  34365=>"110111000",
  34366=>"000011111",
  34367=>"100000001",
  34368=>"100011011",
  34369=>"000101011",
  34370=>"101101101",
  34371=>"000100110",
  34372=>"111000000",
  34373=>"101010000",
  34374=>"001000001",
  34375=>"100110111",
  34376=>"111011101",
  34377=>"001110011",
  34378=>"101110110",
  34379=>"001100001",
  34380=>"100001010",
  34381=>"010011001",
  34382=>"010010011",
  34383=>"111011110",
  34384=>"101111010",
  34385=>"100000000",
  34386=>"101011000",
  34387=>"111101111",
  34388=>"010000010",
  34389=>"110111100",
  34390=>"101000111",
  34391=>"110010101",
  34392=>"000000100",
  34393=>"010111111",
  34394=>"101000111",
  34395=>"111101011",
  34396=>"000010000",
  34397=>"101010001",
  34398=>"101000010",
  34399=>"111100110",
  34400=>"111111101",
  34401=>"000100110",
  34402=>"101001010",
  34403=>"011001011",
  34404=>"101011111",
  34405=>"100101101",
  34406=>"111111111",
  34407=>"000000101",
  34408=>"110010101",
  34409=>"100011001",
  34410=>"100011110",
  34411=>"001100010",
  34412=>"101010000",
  34413=>"111011100",
  34414=>"001100011",
  34415=>"100111111",
  34416=>"101110110",
  34417=>"001011001",
  34418=>"101101001",
  34419=>"111010111",
  34420=>"011111001",
  34421=>"101010110",
  34422=>"111001100",
  34423=>"110111000",
  34424=>"000001010",
  34425=>"001111010",
  34426=>"110010001",
  34427=>"110011101",
  34428=>"101000001",
  34429=>"001001100",
  34430=>"111000000",
  34431=>"001100100",
  34432=>"111110110",
  34433=>"011110001",
  34434=>"010000110",
  34435=>"101001010",
  34436=>"010011100",
  34437=>"001110100",
  34438=>"001100011",
  34439=>"011101111",
  34440=>"001011101",
  34441=>"001000000",
  34442=>"001100000",
  34443=>"000001100",
  34444=>"111001000",
  34445=>"011011110",
  34446=>"011101111",
  34447=>"010110010",
  34448=>"100110011",
  34449=>"010010101",
  34450=>"100110011",
  34451=>"011111100",
  34452=>"100101001",
  34453=>"100111011",
  34454=>"010001110",
  34455=>"011011100",
  34456=>"010111001",
  34457=>"110101101",
  34458=>"001100011",
  34459=>"000010101",
  34460=>"010001111",
  34461=>"000110100",
  34462=>"100111010",
  34463=>"000101100",
  34464=>"100000011",
  34465=>"101101000",
  34466=>"111010011",
  34467=>"011001011",
  34468=>"101110011",
  34469=>"101100010",
  34470=>"101101011",
  34471=>"101110100",
  34472=>"111000000",
  34473=>"101100111",
  34474=>"000110000",
  34475=>"001100111",
  34476=>"111111101",
  34477=>"101001100",
  34478=>"010111000",
  34479=>"111111010",
  34480=>"111001000",
  34481=>"110011111",
  34482=>"000111111",
  34483=>"010111100",
  34484=>"000011101",
  34485=>"000000010",
  34486=>"001011010",
  34487=>"100110000",
  34488=>"111101001",
  34489=>"111110100",
  34490=>"011001001",
  34491=>"111010101",
  34492=>"000011111",
  34493=>"101110111",
  34494=>"000001100",
  34495=>"010100100",
  34496=>"001111110",
  34497=>"110100100",
  34498=>"100100110",
  34499=>"000011111",
  34500=>"100011000",
  34501=>"100111001",
  34502=>"001010110",
  34503=>"010111010",
  34504=>"100010111",
  34505=>"010011100",
  34506=>"000100101",
  34507=>"001001100",
  34508=>"110111001",
  34509=>"111100011",
  34510=>"001010110",
  34511=>"111011101",
  34512=>"011001001",
  34513=>"000111100",
  34514=>"100001011",
  34515=>"101010101",
  34516=>"111110111",
  34517=>"011110011",
  34518=>"110110000",
  34519=>"100001010",
  34520=>"001101110",
  34521=>"110110101",
  34522=>"001101110",
  34523=>"110001111",
  34524=>"001101110",
  34525=>"001100110",
  34526=>"111011111",
  34527=>"100111000",
  34528=>"100100101",
  34529=>"111011010",
  34530=>"001100001",
  34531=>"011110100",
  34532=>"010010100",
  34533=>"000111011",
  34534=>"010100110",
  34535=>"110010010",
  34536=>"010111111",
  34537=>"001011101",
  34538=>"000001101",
  34539=>"011100100",
  34540=>"111010101",
  34541=>"010111000",
  34542=>"001100010",
  34543=>"111001011",
  34544=>"001010000",
  34545=>"101001000",
  34546=>"010111000",
  34547=>"001010111",
  34548=>"000111111",
  34549=>"010000100",
  34550=>"110011101",
  34551=>"010100111",
  34552=>"001010100",
  34553=>"100101001",
  34554=>"101101101",
  34555=>"011100111",
  34556=>"100011001",
  34557=>"001000010",
  34558=>"101101101",
  34559=>"100100000",
  34560=>"111100100",
  34561=>"100000111",
  34562=>"001000111",
  34563=>"011011011",
  34564=>"001100000",
  34565=>"101010010",
  34566=>"111011001",
  34567=>"100011011",
  34568=>"001111010",
  34569=>"110101111",
  34570=>"011000110",
  34571=>"000010000",
  34572=>"010010101",
  34573=>"101110111",
  34574=>"100011001",
  34575=>"001101010",
  34576=>"011000110",
  34577=>"110001101",
  34578=>"101010001",
  34579=>"000110100",
  34580=>"010011010",
  34581=>"011110101",
  34582=>"110011111",
  34583=>"111101010",
  34584=>"010010011",
  34585=>"001010011",
  34586=>"100001100",
  34587=>"001100110",
  34588=>"101101001",
  34589=>"011000111",
  34590=>"011100010",
  34591=>"110110111",
  34592=>"010000111",
  34593=>"101011101",
  34594=>"101010010",
  34595=>"000000111",
  34596=>"110011001",
  34597=>"011100011",
  34598=>"001011010",
  34599=>"110001100",
  34600=>"111010011",
  34601=>"111011100",
  34602=>"000111100",
  34603=>"001010100",
  34604=>"000010110",
  34605=>"001111000",
  34606=>"111001001",
  34607=>"000100000",
  34608=>"000011100",
  34609=>"111100111",
  34610=>"011000011",
  34611=>"010011110",
  34612=>"111101010",
  34613=>"101101111",
  34614=>"001001100",
  34615=>"000001001",
  34616=>"011001000",
  34617=>"101111100",
  34618=>"111001010",
  34619=>"111110001",
  34620=>"110001001",
  34621=>"010011101",
  34622=>"001001000",
  34623=>"111111111",
  34624=>"110110101",
  34625=>"010001010",
  34626=>"100011111",
  34627=>"000000000",
  34628=>"010100101",
  34629=>"000100100",
  34630=>"110001101",
  34631=>"001101000",
  34632=>"001110011",
  34633=>"111001001",
  34634=>"101110011",
  34635=>"010100001",
  34636=>"000011011",
  34637=>"110100110",
  34638=>"000101110",
  34639=>"000010111",
  34640=>"010010110",
  34641=>"100011001",
  34642=>"011011110",
  34643=>"100011111",
  34644=>"100101000",
  34645=>"000000010",
  34646=>"111000011",
  34647=>"000101011",
  34648=>"100011000",
  34649=>"000001000",
  34650=>"011110011",
  34651=>"101101011",
  34652=>"101100100",
  34653=>"011110100",
  34654=>"111110011",
  34655=>"010010001",
  34656=>"110101110",
  34657=>"000011001",
  34658=>"010100010",
  34659=>"000010000",
  34660=>"100000000",
  34661=>"011101001",
  34662=>"000000101",
  34663=>"111000011",
  34664=>"011000001",
  34665=>"000001111",
  34666=>"101110001",
  34667=>"000111101",
  34668=>"001010001",
  34669=>"010110100",
  34670=>"011101000",
  34671=>"101101001",
  34672=>"001100110",
  34673=>"011011111",
  34674=>"111011100",
  34675=>"000001101",
  34676=>"010001010",
  34677=>"111100000",
  34678=>"111100101",
  34679=>"000100111",
  34680=>"100001110",
  34681=>"000010000",
  34682=>"011001100",
  34683=>"000000110",
  34684=>"000010111",
  34685=>"111001001",
  34686=>"101100011",
  34687=>"001101011",
  34688=>"101000011",
  34689=>"111110100",
  34690=>"000010110",
  34691=>"110000101",
  34692=>"011111100",
  34693=>"101010000",
  34694=>"110000100",
  34695=>"000011100",
  34696=>"000110110",
  34697=>"011011101",
  34698=>"100111111",
  34699=>"000111010",
  34700=>"111011100",
  34701=>"110011111",
  34702=>"111010110",
  34703=>"110001000",
  34704=>"100111010",
  34705=>"001001011",
  34706=>"101011011",
  34707=>"111010001",
  34708=>"011010001",
  34709=>"000000101",
  34710=>"000100101",
  34711=>"110101010",
  34712=>"101110110",
  34713=>"101000000",
  34714=>"101001011",
  34715=>"111001100",
  34716=>"110011110",
  34717=>"001111111",
  34718=>"011000111",
  34719=>"011111010",
  34720=>"110110011",
  34721=>"001011111",
  34722=>"001011011",
  34723=>"110011011",
  34724=>"010011100",
  34725=>"101100001",
  34726=>"100000111",
  34727=>"100010100",
  34728=>"110110110",
  34729=>"101111001",
  34730=>"010001011",
  34731=>"111101000",
  34732=>"110101110",
  34733=>"010100101",
  34734=>"111001110",
  34735=>"000011110",
  34736=>"100100000",
  34737=>"111101001",
  34738=>"001011100",
  34739=>"001000001",
  34740=>"011110001",
  34741=>"001110011",
  34742=>"100010011",
  34743=>"101110101",
  34744=>"011111110",
  34745=>"100101100",
  34746=>"100010011",
  34747=>"100001101",
  34748=>"000100000",
  34749=>"111110001",
  34750=>"010000010",
  34751=>"011100010",
  34752=>"101011010",
  34753=>"011101001",
  34754=>"110010100",
  34755=>"010110110",
  34756=>"010101101",
  34757=>"000001100",
  34758=>"101011101",
  34759=>"100010010",
  34760=>"000011001",
  34761=>"000101000",
  34762=>"010000110",
  34763=>"000100000",
  34764=>"101100110",
  34765=>"111110000",
  34766=>"000010101",
  34767=>"101100111",
  34768=>"111100101",
  34769=>"000001010",
  34770=>"111111001",
  34771=>"010100000",
  34772=>"000001110",
  34773=>"000001111",
  34774=>"010001101",
  34775=>"010000101",
  34776=>"010101110",
  34777=>"001111110",
  34778=>"111100100",
  34779=>"101001111",
  34780=>"000010010",
  34781=>"111101111",
  34782=>"010010011",
  34783=>"011000011",
  34784=>"110101110",
  34785=>"000101011",
  34786=>"001110010",
  34787=>"001001001",
  34788=>"010000100",
  34789=>"111011111",
  34790=>"010000000",
  34791=>"000110100",
  34792=>"011001010",
  34793=>"011011101",
  34794=>"110110001",
  34795=>"100010111",
  34796=>"100001011",
  34797=>"111110100",
  34798=>"111111110",
  34799=>"111101101",
  34800=>"000000101",
  34801=>"010110111",
  34802=>"111100010",
  34803=>"001110010",
  34804=>"111101110",
  34805=>"110101011",
  34806=>"001101001",
  34807=>"110101000",
  34808=>"101000011",
  34809=>"100101101",
  34810=>"001100000",
  34811=>"001000100",
  34812=>"000100001",
  34813=>"100010010",
  34814=>"111001001",
  34815=>"001100100",
  34816=>"010000000",
  34817=>"001001001",
  34818=>"000110101",
  34819=>"100000111",
  34820=>"011001011",
  34821=>"000000001",
  34822=>"110000010",
  34823=>"001101000",
  34824=>"011000000",
  34825=>"111111100",
  34826=>"001000001",
  34827=>"011101011",
  34828=>"010111100",
  34829=>"000101000",
  34830=>"111111101",
  34831=>"010100110",
  34832=>"100011100",
  34833=>"001010000",
  34834=>"110110110",
  34835=>"110111101",
  34836=>"010010011",
  34837=>"110100001",
  34838=>"101111110",
  34839=>"000110100",
  34840=>"010001010",
  34841=>"000011001",
  34842=>"110101001",
  34843=>"000001101",
  34844=>"111100001",
  34845=>"111001101",
  34846=>"100010011",
  34847=>"101001001",
  34848=>"100001011",
  34849=>"101110111",
  34850=>"010111110",
  34851=>"000110010",
  34852=>"110110000",
  34853=>"101001100",
  34854=>"010111110",
  34855=>"011101010",
  34856=>"101011100",
  34857=>"110101111",
  34858=>"110011000",
  34859=>"010000010",
  34860=>"100000000",
  34861=>"000000000",
  34862=>"000111100",
  34863=>"000101110",
  34864=>"100000001",
  34865=>"111100111",
  34866=>"000010001",
  34867=>"100010001",
  34868=>"000110000",
  34869=>"110001000",
  34870=>"110000110",
  34871=>"011011011",
  34872=>"100011001",
  34873=>"110011100",
  34874=>"011101001",
  34875=>"010101100",
  34876=>"001001001",
  34877=>"001111110",
  34878=>"010111001",
  34879=>"101010000",
  34880=>"010000110",
  34881=>"000001100",
  34882=>"111011000",
  34883=>"010100110",
  34884=>"001100010",
  34885=>"100000000",
  34886=>"011110110",
  34887=>"101101110",
  34888=>"010011111",
  34889=>"110111001",
  34890=>"100100100",
  34891=>"001101101",
  34892=>"110000111",
  34893=>"100000011",
  34894=>"111101110",
  34895=>"001001111",
  34896=>"101110110",
  34897=>"000001011",
  34898=>"000010000",
  34899=>"111110010",
  34900=>"000110100",
  34901=>"100001111",
  34902=>"111011001",
  34903=>"010101010",
  34904=>"110001111",
  34905=>"111000011",
  34906=>"010010000",
  34907=>"010110000",
  34908=>"000111000",
  34909=>"110101101",
  34910=>"110010110",
  34911=>"011111011",
  34912=>"000111100",
  34913=>"100010101",
  34914=>"111100000",
  34915=>"001101001",
  34916=>"001001101",
  34917=>"101101001",
  34918=>"101100100",
  34919=>"100010110",
  34920=>"000001101",
  34921=>"111000001",
  34922=>"111110011",
  34923=>"010001101",
  34924=>"000111101",
  34925=>"101000010",
  34926=>"011100011",
  34927=>"101100100",
  34928=>"010111001",
  34929=>"011011110",
  34930=>"011000010",
  34931=>"010010100",
  34932=>"011010001",
  34933=>"101110111",
  34934=>"111000111",
  34935=>"100110010",
  34936=>"101111010",
  34937=>"110001110",
  34938=>"011011011",
  34939=>"101011111",
  34940=>"010101110",
  34941=>"101101000",
  34942=>"010110000",
  34943=>"111100110",
  34944=>"101010101",
  34945=>"110010001",
  34946=>"111101111",
  34947=>"111011010",
  34948=>"000000111",
  34949=>"110101010",
  34950=>"101110001",
  34951=>"101010110",
  34952=>"100001010",
  34953=>"111110000",
  34954=>"000001100",
  34955=>"110100011",
  34956=>"000010000",
  34957=>"000110000",
  34958=>"111010011",
  34959=>"111111101",
  34960=>"000001100",
  34961=>"100010101",
  34962=>"011010100",
  34963=>"000100111",
  34964=>"011011111",
  34965=>"011001100",
  34966=>"010010111",
  34967=>"000110101",
  34968=>"011001111",
  34969=>"101001010",
  34970=>"110010101",
  34971=>"101111000",
  34972=>"000100001",
  34973=>"110001000",
  34974=>"101001011",
  34975=>"001001111",
  34976=>"000100001",
  34977=>"110010000",
  34978=>"110110011",
  34979=>"101110000",
  34980=>"101001000",
  34981=>"110101110",
  34982=>"000001100",
  34983=>"100111101",
  34984=>"010001100",
  34985=>"000000000",
  34986=>"000001100",
  34987=>"010100010",
  34988=>"100011000",
  34989=>"111110010",
  34990=>"100111010",
  34991=>"111010111",
  34992=>"001111001",
  34993=>"011001100",
  34994=>"111001000",
  34995=>"000000001",
  34996=>"100011100",
  34997=>"100010001",
  34998=>"100000001",
  34999=>"010111011",
  35000=>"110100011",
  35001=>"010110111",
  35002=>"011010010",
  35003=>"111011010",
  35004=>"111000010",
  35005=>"011111110",
  35006=>"010010001",
  35007=>"100110000",
  35008=>"111010100",
  35009=>"000110111",
  35010=>"101110111",
  35011=>"000001001",
  35012=>"100100101",
  35013=>"101101110",
  35014=>"011000100",
  35015=>"000010001",
  35016=>"100000110",
  35017=>"000101110",
  35018=>"110000000",
  35019=>"111100100",
  35020=>"001011110",
  35021=>"010111110",
  35022=>"000111101",
  35023=>"100101111",
  35024=>"100111011",
  35025=>"011001110",
  35026=>"001000111",
  35027=>"110000010",
  35028=>"000000101",
  35029=>"001111111",
  35030=>"101000100",
  35031=>"010000101",
  35032=>"000000101",
  35033=>"110111001",
  35034=>"010101101",
  35035=>"000110011",
  35036=>"001001000",
  35037=>"111111111",
  35038=>"101110101",
  35039=>"011110110",
  35040=>"111000110",
  35041=>"011101100",
  35042=>"101000100",
  35043=>"010000111",
  35044=>"001010000",
  35045=>"111000111",
  35046=>"010110111",
  35047=>"010000101",
  35048=>"010111010",
  35049=>"100111101",
  35050=>"111011001",
  35051=>"110101010",
  35052=>"010001110",
  35053=>"000000110",
  35054=>"100011000",
  35055=>"111110101",
  35056=>"001110101",
  35057=>"010010011",
  35058=>"000011111",
  35059=>"000110000",
  35060=>"110010010",
  35061=>"011000001",
  35062=>"001100001",
  35063=>"000101100",
  35064=>"001011001",
  35065=>"110110011",
  35066=>"011000010",
  35067=>"011110110",
  35068=>"010011001",
  35069=>"000110110",
  35070=>"110000110",
  35071=>"101100000",
  35072=>"110111110",
  35073=>"111001001",
  35074=>"100101001",
  35075=>"110101010",
  35076=>"011011010",
  35077=>"101001100",
  35078=>"110001001",
  35079=>"111011100",
  35080=>"110101011",
  35081=>"100111010",
  35082=>"101110010",
  35083=>"110001010",
  35084=>"111100001",
  35085=>"111101011",
  35086=>"101100001",
  35087=>"010111010",
  35088=>"011010001",
  35089=>"110101010",
  35090=>"101110110",
  35091=>"101101110",
  35092=>"111000101",
  35093=>"110101010",
  35094=>"010100100",
  35095=>"011100011",
  35096=>"011000010",
  35097=>"100111100",
  35098=>"110001110",
  35099=>"011100100",
  35100=>"000010011",
  35101=>"010000011",
  35102=>"000000101",
  35103=>"000010100",
  35104=>"011010101",
  35105=>"111010110",
  35106=>"011011000",
  35107=>"010111011",
  35108=>"100011100",
  35109=>"111110010",
  35110=>"010001111",
  35111=>"011000010",
  35112=>"000000011",
  35113=>"111111110",
  35114=>"101111100",
  35115=>"011010000",
  35116=>"010001000",
  35117=>"001000101",
  35118=>"011111001",
  35119=>"001111000",
  35120=>"101011111",
  35121=>"100101101",
  35122=>"001010010",
  35123=>"110110110",
  35124=>"000000000",
  35125=>"000001011",
  35126=>"111111110",
  35127=>"011101111",
  35128=>"010000001",
  35129=>"001010101",
  35130=>"001101010",
  35131=>"111100110",
  35132=>"001000110",
  35133=>"101001010",
  35134=>"000010100",
  35135=>"101011011",
  35136=>"010011111",
  35137=>"101111111",
  35138=>"100101010",
  35139=>"110111000",
  35140=>"100111110",
  35141=>"001010010",
  35142=>"111011000",
  35143=>"111101000",
  35144=>"111100110",
  35145=>"111111110",
  35146=>"111011111",
  35147=>"010101100",
  35148=>"011000000",
  35149=>"001010010",
  35150=>"111100101",
  35151=>"110111001",
  35152=>"110110101",
  35153=>"101110101",
  35154=>"001110000",
  35155=>"111100110",
  35156=>"110100000",
  35157=>"111011110",
  35158=>"010011000",
  35159=>"011110110",
  35160=>"010010011",
  35161=>"101100010",
  35162=>"110100101",
  35163=>"100000011",
  35164=>"010001101",
  35165=>"001001101",
  35166=>"110110011",
  35167=>"111000101",
  35168=>"001001110",
  35169=>"000001110",
  35170=>"110001110",
  35171=>"001100001",
  35172=>"111101111",
  35173=>"001101110",
  35174=>"101001000",
  35175=>"010111000",
  35176=>"011000101",
  35177=>"001100001",
  35178=>"011111110",
  35179=>"101100101",
  35180=>"000011011",
  35181=>"000001110",
  35182=>"110010110",
  35183=>"001001001",
  35184=>"111111011",
  35185=>"111000000",
  35186=>"100001101",
  35187=>"110110001",
  35188=>"111000011",
  35189=>"100110000",
  35190=>"111110001",
  35191=>"001100001",
  35192=>"100001010",
  35193=>"010000000",
  35194=>"001100100",
  35195=>"111111110",
  35196=>"001101101",
  35197=>"001100001",
  35198=>"011110000",
  35199=>"000010110",
  35200=>"101001011",
  35201=>"011101010",
  35202=>"110111110",
  35203=>"111001110",
  35204=>"011011011",
  35205=>"001010100",
  35206=>"001111001",
  35207=>"010001011",
  35208=>"101101000",
  35209=>"100110101",
  35210=>"100011100",
  35211=>"101001001",
  35212=>"110000000",
  35213=>"100101100",
  35214=>"101110110",
  35215=>"110100001",
  35216=>"000100101",
  35217=>"110000000",
  35218=>"001010010",
  35219=>"010101000",
  35220=>"110111101",
  35221=>"100100100",
  35222=>"001011010",
  35223=>"010000011",
  35224=>"000110110",
  35225=>"010111101",
  35226=>"010010001",
  35227=>"101111111",
  35228=>"111010000",
  35229=>"010101011",
  35230=>"001000010",
  35231=>"011101010",
  35232=>"100100110",
  35233=>"111000010",
  35234=>"010001001",
  35235=>"100001011",
  35236=>"010100110",
  35237=>"111001011",
  35238=>"111100011",
  35239=>"100110001",
  35240=>"000100000",
  35241=>"001101111",
  35242=>"000101110",
  35243=>"000011101",
  35244=>"110011111",
  35245=>"001001111",
  35246=>"010110010",
  35247=>"110100101",
  35248=>"000111010",
  35249=>"000101010",
  35250=>"010011100",
  35251=>"101100011",
  35252=>"110110011",
  35253=>"110000101",
  35254=>"101111010",
  35255=>"001100000",
  35256=>"101001001",
  35257=>"010100010",
  35258=>"011000000",
  35259=>"101100110",
  35260=>"111010111",
  35261=>"100000111",
  35262=>"011011000",
  35263=>"110101001",
  35264=>"011011101",
  35265=>"111011010",
  35266=>"111000000",
  35267=>"001001101",
  35268=>"001000000",
  35269=>"110001010",
  35270=>"001000000",
  35271=>"101011001",
  35272=>"101001011",
  35273=>"000010001",
  35274=>"010000100",
  35275=>"100111011",
  35276=>"000001110",
  35277=>"011100001",
  35278=>"001110001",
  35279=>"011110000",
  35280=>"100000000",
  35281=>"101111111",
  35282=>"111111011",
  35283=>"101111001",
  35284=>"010000000",
  35285=>"111100010",
  35286=>"010100100",
  35287=>"001000011",
  35288=>"111110000",
  35289=>"111111010",
  35290=>"010000000",
  35291=>"000011001",
  35292=>"110101100",
  35293=>"100110100",
  35294=>"000111101",
  35295=>"100011111",
  35296=>"110111000",
  35297=>"000001110",
  35298=>"010101011",
  35299=>"101111010",
  35300=>"111111010",
  35301=>"100011010",
  35302=>"010110100",
  35303=>"010101001",
  35304=>"001000010",
  35305=>"011011010",
  35306=>"100010001",
  35307=>"011100100",
  35308=>"110111001",
  35309=>"000101101",
  35310=>"010010011",
  35311=>"000101101",
  35312=>"110101101",
  35313=>"110101011",
  35314=>"000100001",
  35315=>"001101100",
  35316=>"000000000",
  35317=>"110010111",
  35318=>"011110010",
  35319=>"111110010",
  35320=>"000100111",
  35321=>"011000110",
  35322=>"001001011",
  35323=>"000101011",
  35324=>"010001100",
  35325=>"000000010",
  35326=>"110110111",
  35327=>"010010110",
  35328=>"100001011",
  35329=>"011100100",
  35330=>"001010110",
  35331=>"101000101",
  35332=>"100110001",
  35333=>"000110001",
  35334=>"111111101",
  35335=>"010110000",
  35336=>"100011000",
  35337=>"100110010",
  35338=>"010011010",
  35339=>"111100010",
  35340=>"101011001",
  35341=>"111100001",
  35342=>"000110001",
  35343=>"101101011",
  35344=>"000000111",
  35345=>"001001010",
  35346=>"101010001",
  35347=>"010001011",
  35348=>"110011010",
  35349=>"101000111",
  35350=>"110100000",
  35351=>"100001011",
  35352=>"111111110",
  35353=>"111110100",
  35354=>"111000000",
  35355=>"001100000",
  35356=>"000110011",
  35357=>"000110001",
  35358=>"000111110",
  35359=>"010001111",
  35360=>"111010000",
  35361=>"010101010",
  35362=>"100100010",
  35363=>"100000000",
  35364=>"011001111",
  35365=>"011010111",
  35366=>"110011110",
  35367=>"100010001",
  35368=>"110000000",
  35369=>"001101010",
  35370=>"000010100",
  35371=>"000100010",
  35372=>"110111001",
  35373=>"110010010",
  35374=>"111111101",
  35375=>"110100001",
  35376=>"110011111",
  35377=>"111100001",
  35378=>"010010010",
  35379=>"100000110",
  35380=>"001001010",
  35381=>"100010111",
  35382=>"011011111",
  35383=>"111011111",
  35384=>"101110100",
  35385=>"011011010",
  35386=>"100111111",
  35387=>"001011101",
  35388=>"001101010",
  35389=>"010001000",
  35390=>"000100010",
  35391=>"011001100",
  35392=>"000111000",
  35393=>"111101110",
  35394=>"001001000",
  35395=>"011111111",
  35396=>"000101101",
  35397=>"001101010",
  35398=>"001100010",
  35399=>"010100111",
  35400=>"100110001",
  35401=>"011111101",
  35402=>"001001111",
  35403=>"010001111",
  35404=>"100011100",
  35405=>"111001001",
  35406=>"101000000",
  35407=>"110000111",
  35408=>"010100010",
  35409=>"101011101",
  35410=>"001011111",
  35411=>"101110100",
  35412=>"110100010",
  35413=>"100001010",
  35414=>"101101011",
  35415=>"111110010",
  35416=>"010111110",
  35417=>"100101011",
  35418=>"100111011",
  35419=>"110110011",
  35420=>"010101001",
  35421=>"100001100",
  35422=>"001111111",
  35423=>"111001100",
  35424=>"101011100",
  35425=>"000110100",
  35426=>"100010001",
  35427=>"101010100",
  35428=>"000010111",
  35429=>"010000010",
  35430=>"110011010",
  35431=>"001000010",
  35432=>"101001101",
  35433=>"101010000",
  35434=>"011111000",
  35435=>"100100001",
  35436=>"010110111",
  35437=>"110000110",
  35438=>"100111000",
  35439=>"111010110",
  35440=>"101101111",
  35441=>"010001100",
  35442=>"101110111",
  35443=>"010110101",
  35444=>"000110101",
  35445=>"101011111",
  35446=>"000010111",
  35447=>"100011111",
  35448=>"010100110",
  35449=>"101001111",
  35450=>"100100011",
  35451=>"111101000",
  35452=>"111111111",
  35453=>"010101100",
  35454=>"001011111",
  35455=>"101111100",
  35456=>"010001000",
  35457=>"100011110",
  35458=>"010000001",
  35459=>"001000101",
  35460=>"110011110",
  35461=>"011000111",
  35462=>"111101010",
  35463=>"111110111",
  35464=>"001001111",
  35465=>"101001011",
  35466=>"010011110",
  35467=>"001001110",
  35468=>"101100010",
  35469=>"101001110",
  35470=>"100101111",
  35471=>"110001111",
  35472=>"111001110",
  35473=>"111010111",
  35474=>"110000010",
  35475=>"000000100",
  35476=>"100100101",
  35477=>"110010111",
  35478=>"100000001",
  35479=>"100000010",
  35480=>"011101010",
  35481=>"000010111",
  35482=>"001000000",
  35483=>"110111010",
  35484=>"001010111",
  35485=>"101010010",
  35486=>"101011101",
  35487=>"011111010",
  35488=>"111000011",
  35489=>"101001101",
  35490=>"111001100",
  35491=>"010011000",
  35492=>"001000101",
  35493=>"101010001",
  35494=>"101111010",
  35495=>"110101101",
  35496=>"001011001",
  35497=>"001110110",
  35498=>"010101100",
  35499=>"111011001",
  35500=>"111100011",
  35501=>"111000011",
  35502=>"010000100",
  35503=>"101100110",
  35504=>"010001001",
  35505=>"111110010",
  35506=>"011010001",
  35507=>"011110100",
  35508=>"011000101",
  35509=>"001011000",
  35510=>"101000100",
  35511=>"011100101",
  35512=>"101100111",
  35513=>"001011000",
  35514=>"100100000",
  35515=>"001100000",
  35516=>"110011101",
  35517=>"000110011",
  35518=>"001100101",
  35519=>"001000000",
  35520=>"010111101",
  35521=>"010010011",
  35522=>"101010011",
  35523=>"101111010",
  35524=>"110001011",
  35525=>"111011000",
  35526=>"010101100",
  35527=>"000001000",
  35528=>"111000110",
  35529=>"010011110",
  35530=>"000011111",
  35531=>"011000101",
  35532=>"010011101",
  35533=>"011100111",
  35534=>"000101110",
  35535=>"010100010",
  35536=>"000100111",
  35537=>"110101100",
  35538=>"011001101",
  35539=>"001000100",
  35540=>"000111001",
  35541=>"010001001",
  35542=>"000000111",
  35543=>"111110101",
  35544=>"110100100",
  35545=>"111100101",
  35546=>"011011111",
  35547=>"100001100",
  35548=>"110011111",
  35549=>"000100010",
  35550=>"000110100",
  35551=>"101111110",
  35552=>"011010011",
  35553=>"010011111",
  35554=>"110000100",
  35555=>"010001001",
  35556=>"010101100",
  35557=>"100011010",
  35558=>"000110110",
  35559=>"001101110",
  35560=>"111010011",
  35561=>"001110011",
  35562=>"001001001",
  35563=>"011001000",
  35564=>"010001101",
  35565=>"000100111",
  35566=>"010101100",
  35567=>"010110010",
  35568=>"011111111",
  35569=>"001000000",
  35570=>"011100000",
  35571=>"011010100",
  35572=>"101011110",
  35573=>"000110101",
  35574=>"100111111",
  35575=>"010011100",
  35576=>"101100011",
  35577=>"111010001",
  35578=>"111000000",
  35579=>"101010111",
  35580=>"111100111",
  35581=>"100110110",
  35582=>"010010110",
  35583=>"001001000",
  35584=>"010010011",
  35585=>"000110110",
  35586=>"011000011",
  35587=>"011101111",
  35588=>"000011110",
  35589=>"000000100",
  35590=>"100110111",
  35591=>"000011101",
  35592=>"110111000",
  35593=>"111110111",
  35594=>"101010000",
  35595=>"010100000",
  35596=>"010000011",
  35597=>"011011101",
  35598=>"101101000",
  35599=>"001100000",
  35600=>"000001110",
  35601=>"001001111",
  35602=>"101110101",
  35603=>"001000101",
  35604=>"110100101",
  35605=>"000110110",
  35606=>"000101110",
  35607=>"111001101",
  35608=>"111010111",
  35609=>"001100000",
  35610=>"010000111",
  35611=>"001000110",
  35612=>"001101010",
  35613=>"100000000",
  35614=>"000000111",
  35615=>"000000100",
  35616=>"110100010",
  35617=>"111001010",
  35618=>"100001010",
  35619=>"111000101",
  35620=>"010100001",
  35621=>"101000111",
  35622=>"110101010",
  35623=>"100000110",
  35624=>"101000000",
  35625=>"111000111",
  35626=>"000111000",
  35627=>"010110010",
  35628=>"100111011",
  35629=>"001001011",
  35630=>"001010000",
  35631=>"011000111",
  35632=>"010011011",
  35633=>"001101010",
  35634=>"011100110",
  35635=>"110000100",
  35636=>"010110101",
  35637=>"000111000",
  35638=>"010101111",
  35639=>"100001101",
  35640=>"111000011",
  35641=>"000001000",
  35642=>"001101000",
  35643=>"010110011",
  35644=>"111011000",
  35645=>"011101001",
  35646=>"000000001",
  35647=>"010000111",
  35648=>"000001100",
  35649=>"110010000",
  35650=>"111000101",
  35651=>"010000011",
  35652=>"010001010",
  35653=>"001000100",
  35654=>"001000101",
  35655=>"111110101",
  35656=>"001101001",
  35657=>"100001110",
  35658=>"001001101",
  35659=>"011100010",
  35660=>"100100001",
  35661=>"100011000",
  35662=>"000000010",
  35663=>"000100011",
  35664=>"111010000",
  35665=>"000010001",
  35666=>"001111101",
  35667=>"001101100",
  35668=>"110000100",
  35669=>"010100100",
  35670=>"111011000",
  35671=>"100000000",
  35672=>"111101001",
  35673=>"111101011",
  35674=>"000010110",
  35675=>"000010010",
  35676=>"110100000",
  35677=>"010001010",
  35678=>"000110110",
  35679=>"101001111",
  35680=>"010111010",
  35681=>"001110101",
  35682=>"111111101",
  35683=>"001100011",
  35684=>"111001100",
  35685=>"010001011",
  35686=>"000110111",
  35687=>"111010011",
  35688=>"001100100",
  35689=>"111111111",
  35690=>"010111101",
  35691=>"100111011",
  35692=>"111000100",
  35693=>"100101100",
  35694=>"110011000",
  35695=>"000001100",
  35696=>"001011100",
  35697=>"001111101",
  35698=>"010100000",
  35699=>"001011110",
  35700=>"011101111",
  35701=>"001000001",
  35702=>"100001110",
  35703=>"000000100",
  35704=>"111101001",
  35705=>"010000111",
  35706=>"101111011",
  35707=>"011011101",
  35708=>"010001100",
  35709=>"011000101",
  35710=>"011011010",
  35711=>"011100111",
  35712=>"111011010",
  35713=>"001010011",
  35714=>"111010111",
  35715=>"001110101",
  35716=>"000100100",
  35717=>"110100000",
  35718=>"110110110",
  35719=>"000011110",
  35720=>"001000010",
  35721=>"101111010",
  35722=>"111000101",
  35723=>"011110000",
  35724=>"010100101",
  35725=>"101100101",
  35726=>"111111111",
  35727=>"101101110",
  35728=>"110001101",
  35729=>"100110010",
  35730=>"000111111",
  35731=>"011001100",
  35732=>"010010100",
  35733=>"110000110",
  35734=>"110011001",
  35735=>"010000101",
  35736=>"111111011",
  35737=>"000101111",
  35738=>"111111100",
  35739=>"100111111",
  35740=>"110001010",
  35741=>"011101101",
  35742=>"011011010",
  35743=>"000111011",
  35744=>"101100111",
  35745=>"101001011",
  35746=>"010100101",
  35747=>"001001100",
  35748=>"101111000",
  35749=>"111111111",
  35750=>"100101101",
  35751=>"111110001",
  35752=>"010011000",
  35753=>"110110110",
  35754=>"001111111",
  35755=>"110111000",
  35756=>"101001010",
  35757=>"000000100",
  35758=>"101001111",
  35759=>"001110010",
  35760=>"110011010",
  35761=>"111101111",
  35762=>"001111100",
  35763=>"110001010",
  35764=>"110001001",
  35765=>"011101110",
  35766=>"011111110",
  35767=>"101001001",
  35768=>"110100110",
  35769=>"110011010",
  35770=>"100101110",
  35771=>"010010110",
  35772=>"100011000",
  35773=>"000110011",
  35774=>"100111001",
  35775=>"010101000",
  35776=>"111111001",
  35777=>"110101101",
  35778=>"101010011",
  35779=>"001110100",
  35780=>"011010001",
  35781=>"000100111",
  35782=>"111011011",
  35783=>"010000000",
  35784=>"010100000",
  35785=>"111111111",
  35786=>"000000001",
  35787=>"100111000",
  35788=>"110111111",
  35789=>"000011010",
  35790=>"110100111",
  35791=>"100110110",
  35792=>"100011110",
  35793=>"101110111",
  35794=>"001111000",
  35795=>"000101111",
  35796=>"000010100",
  35797=>"001101001",
  35798=>"000010110",
  35799=>"110011111",
  35800=>"111111110",
  35801=>"000001011",
  35802=>"111001000",
  35803=>"101001111",
  35804=>"100110010",
  35805=>"111000010",
  35806=>"001000000",
  35807=>"001100101",
  35808=>"101011110",
  35809=>"010001011",
  35810=>"010001001",
  35811=>"011010111",
  35812=>"111010000",
  35813=>"101001110",
  35814=>"110100100",
  35815=>"101000000",
  35816=>"101101111",
  35817=>"010001111",
  35818=>"110000110",
  35819=>"110111111",
  35820=>"101110001",
  35821=>"111010110",
  35822=>"010101000",
  35823=>"110111110",
  35824=>"010101111",
  35825=>"100010001",
  35826=>"001001100",
  35827=>"011110110",
  35828=>"100101111",
  35829=>"010001000",
  35830=>"100110001",
  35831=>"101001010",
  35832=>"011110100",
  35833=>"101100011",
  35834=>"100100001",
  35835=>"110111001",
  35836=>"101100110",
  35837=>"100011011",
  35838=>"110011010",
  35839=>"001111101",
  35840=>"001110110",
  35841=>"101111110",
  35842=>"100100000",
  35843=>"001001010",
  35844=>"010101011",
  35845=>"100011010",
  35846=>"100111001",
  35847=>"001010000",
  35848=>"010111110",
  35849=>"100111010",
  35850=>"100000111",
  35851=>"100000011",
  35852=>"111110101",
  35853=>"001001110",
  35854=>"011010110",
  35855=>"100100011",
  35856=>"010010000",
  35857=>"100011101",
  35858=>"111001000",
  35859=>"000011001",
  35860=>"000101000",
  35861=>"011110001",
  35862=>"011110111",
  35863=>"000000100",
  35864=>"101111000",
  35865=>"100110000",
  35866=>"000010000",
  35867=>"100101000",
  35868=>"110001110",
  35869=>"011000110",
  35870=>"011001100",
  35871=>"010000110",
  35872=>"000000010",
  35873=>"000000100",
  35874=>"111111001",
  35875=>"011011111",
  35876=>"100111101",
  35877=>"100011101",
  35878=>"001000001",
  35879=>"110111000",
  35880=>"111001000",
  35881=>"001100000",
  35882=>"111010100",
  35883=>"101101110",
  35884=>"011001010",
  35885=>"011101001",
  35886=>"101011111",
  35887=>"001101011",
  35888=>"001000010",
  35889=>"001011000",
  35890=>"010000011",
  35891=>"101001011",
  35892=>"011011001",
  35893=>"100100101",
  35894=>"110100010",
  35895=>"110011001",
  35896=>"000000000",
  35897=>"001110011",
  35898=>"010011000",
  35899=>"011100000",
  35900=>"111011011",
  35901=>"110000100",
  35902=>"010100000",
  35903=>"000100100",
  35904=>"001001000",
  35905=>"000101000",
  35906=>"011100001",
  35907=>"000111101",
  35908=>"100110100",
  35909=>"110110100",
  35910=>"011010011",
  35911=>"000101010",
  35912=>"111100001",
  35913=>"100001111",
  35914=>"000110011",
  35915=>"111000111",
  35916=>"010100001",
  35917=>"111111110",
  35918=>"011100101",
  35919=>"000100101",
  35920=>"000101010",
  35921=>"101000101",
  35922=>"000000101",
  35923=>"101100111",
  35924=>"100001110",
  35925=>"001010010",
  35926=>"111000001",
  35927=>"000011010",
  35928=>"011101111",
  35929=>"001010001",
  35930=>"011000100",
  35931=>"111101010",
  35932=>"011100011",
  35933=>"000010000",
  35934=>"001000001",
  35935=>"001010001",
  35936=>"011000100",
  35937=>"101011110",
  35938=>"001000111",
  35939=>"000011000",
  35940=>"010001101",
  35941=>"100010111",
  35942=>"110010010",
  35943=>"000011100",
  35944=>"110010110",
  35945=>"111000110",
  35946=>"000011100",
  35947=>"101101000",
  35948=>"101110011",
  35949=>"101110000",
  35950=>"101010100",
  35951=>"000111010",
  35952=>"100111110",
  35953=>"111011110",
  35954=>"110001011",
  35955=>"000101100",
  35956=>"010100011",
  35957=>"111000001",
  35958=>"011101010",
  35959=>"110001010",
  35960=>"001000001",
  35961=>"110110111",
  35962=>"110100100",
  35963=>"110100100",
  35964=>"011000110",
  35965=>"111110101",
  35966=>"101010011",
  35967=>"110101100",
  35968=>"011011110",
  35969=>"010111011",
  35970=>"100000000",
  35971=>"000010011",
  35972=>"111111010",
  35973=>"101001111",
  35974=>"000001111",
  35975=>"010001101",
  35976=>"100101001",
  35977=>"001001010",
  35978=>"111111011",
  35979=>"011000110",
  35980=>"011001100",
  35981=>"111100101",
  35982=>"001100110",
  35983=>"110100011",
  35984=>"011000110",
  35985=>"110111010",
  35986=>"100001110",
  35987=>"101000000",
  35988=>"000100001",
  35989=>"010001111",
  35990=>"101100100",
  35991=>"001110010",
  35992=>"011101010",
  35993=>"000110110",
  35994=>"011110100",
  35995=>"101101001",
  35996=>"000100110",
  35997=>"110001001",
  35998=>"011101110",
  35999=>"000111100",
  36000=>"111100011",
  36001=>"011111001",
  36002=>"001000001",
  36003=>"101010011",
  36004=>"110011101",
  36005=>"000010001",
  36006=>"101101000",
  36007=>"111111010",
  36008=>"000101110",
  36009=>"011101010",
  36010=>"111110101",
  36011=>"111110011",
  36012=>"000111000",
  36013=>"011001110",
  36014=>"011100101",
  36015=>"100001110",
  36016=>"001100001",
  36017=>"111011101",
  36018=>"101011100",
  36019=>"111111100",
  36020=>"101000000",
  36021=>"100000110",
  36022=>"110100111",
  36023=>"100101010",
  36024=>"111000001",
  36025=>"000100010",
  36026=>"111000100",
  36027=>"100111101",
  36028=>"100111001",
  36029=>"111100110",
  36030=>"111011010",
  36031=>"101101011",
  36032=>"100111000",
  36033=>"110111011",
  36034=>"100010010",
  36035=>"000000011",
  36036=>"110001001",
  36037=>"100000000",
  36038=>"110010000",
  36039=>"101100110",
  36040=>"110011101",
  36041=>"101000001",
  36042=>"111111111",
  36043=>"110110111",
  36044=>"110101011",
  36045=>"010000100",
  36046=>"001111000",
  36047=>"110101110",
  36048=>"011101000",
  36049=>"111101101",
  36050=>"000111101",
  36051=>"111011111",
  36052=>"111100010",
  36053=>"010111100",
  36054=>"101100000",
  36055=>"001001101",
  36056=>"001100000",
  36057=>"111010000",
  36058=>"000000001",
  36059=>"101100000",
  36060=>"111111110",
  36061=>"100101011",
  36062=>"110100101",
  36063=>"100011110",
  36064=>"011110111",
  36065=>"100001110",
  36066=>"011110011",
  36067=>"101000010",
  36068=>"111000110",
  36069=>"100111000",
  36070=>"100100000",
  36071=>"010111001",
  36072=>"011100011",
  36073=>"100001110",
  36074=>"000011100",
  36075=>"010000100",
  36076=>"000100101",
  36077=>"001001010",
  36078=>"110110010",
  36079=>"010111010",
  36080=>"001110101",
  36081=>"101010110",
  36082=>"100111011",
  36083=>"010001001",
  36084=>"110100000",
  36085=>"010000001",
  36086=>"110000100",
  36087=>"110000010",
  36088=>"111001010",
  36089=>"000010110",
  36090=>"111101011",
  36091=>"101101100",
  36092=>"011010101",
  36093=>"001101001",
  36094=>"011101100",
  36095=>"010000001",
  36096=>"000000001",
  36097=>"100111011",
  36098=>"000010100",
  36099=>"101111100",
  36100=>"000111000",
  36101=>"101101110",
  36102=>"100001100",
  36103=>"111001101",
  36104=>"000111110",
  36105=>"010001001",
  36106=>"100010100",
  36107=>"110000010",
  36108=>"100011010",
  36109=>"111101101",
  36110=>"100001001",
  36111=>"110000110",
  36112=>"010011001",
  36113=>"000001001",
  36114=>"100101110",
  36115=>"110100010",
  36116=>"111100010",
  36117=>"110011011",
  36118=>"001110010",
  36119=>"011011000",
  36120=>"011010111",
  36121=>"100000110",
  36122=>"110000010",
  36123=>"101000111",
  36124=>"100100001",
  36125=>"101011100",
  36126=>"101100100",
  36127=>"100000100",
  36128=>"100100001",
  36129=>"100101111",
  36130=>"101000110",
  36131=>"010001111",
  36132=>"010110001",
  36133=>"011100100",
  36134=>"110101110",
  36135=>"001001100",
  36136=>"001010111",
  36137=>"110001111",
  36138=>"001101110",
  36139=>"010100001",
  36140=>"001110100",
  36141=>"111101010",
  36142=>"000011100",
  36143=>"000101011",
  36144=>"011001111",
  36145=>"100101001",
  36146=>"001000100",
  36147=>"000110000",
  36148=>"001110110",
  36149=>"110000001",
  36150=>"001000101",
  36151=>"111010101",
  36152=>"000000000",
  36153=>"111011110",
  36154=>"101100110",
  36155=>"111110000",
  36156=>"110111111",
  36157=>"000000100",
  36158=>"101110101",
  36159=>"101011110",
  36160=>"011101010",
  36161=>"001111000",
  36162=>"101110000",
  36163=>"001000001",
  36164=>"100010100",
  36165=>"001111101",
  36166=>"110110001",
  36167=>"000101110",
  36168=>"011110011",
  36169=>"000101001",
  36170=>"011011001",
  36171=>"011101111",
  36172=>"100000111",
  36173=>"011100111",
  36174=>"010111110",
  36175=>"001111101",
  36176=>"011011010",
  36177=>"001000000",
  36178=>"011011001",
  36179=>"001010000",
  36180=>"101010111",
  36181=>"001001000",
  36182=>"010111100",
  36183=>"000011000",
  36184=>"011111100",
  36185=>"011101001",
  36186=>"111111001",
  36187=>"101011101",
  36188=>"100001000",
  36189=>"100100000",
  36190=>"010001100",
  36191=>"001001010",
  36192=>"000000100",
  36193=>"111010111",
  36194=>"010100000",
  36195=>"100110001",
  36196=>"111100111",
  36197=>"100100110",
  36198=>"010011110",
  36199=>"001110001",
  36200=>"000011101",
  36201=>"111101010",
  36202=>"100000001",
  36203=>"100011101",
  36204=>"011001001",
  36205=>"000101100",
  36206=>"011010101",
  36207=>"010001100",
  36208=>"010011101",
  36209=>"110110001",
  36210=>"111011001",
  36211=>"000010101",
  36212=>"111000111",
  36213=>"101111100",
  36214=>"111011110",
  36215=>"110100010",
  36216=>"010011000",
  36217=>"111001110",
  36218=>"100000101",
  36219=>"100010101",
  36220=>"000100000",
  36221=>"011000100",
  36222=>"101100000",
  36223=>"101111111",
  36224=>"111010000",
  36225=>"101001110",
  36226=>"110101010",
  36227=>"011110000",
  36228=>"100010011",
  36229=>"010000101",
  36230=>"001110001",
  36231=>"011110100",
  36232=>"110011001",
  36233=>"110001100",
  36234=>"101111111",
  36235=>"111000000",
  36236=>"110110110",
  36237=>"110001101",
  36238=>"111010011",
  36239=>"010010101",
  36240=>"101010011",
  36241=>"111011000",
  36242=>"111111000",
  36243=>"011001011",
  36244=>"000111010",
  36245=>"001000001",
  36246=>"111111010",
  36247=>"101101001",
  36248=>"010111010",
  36249=>"000001010",
  36250=>"000000000",
  36251=>"101100001",
  36252=>"111001010",
  36253=>"101000010",
  36254=>"011110001",
  36255=>"000101101",
  36256=>"110101110",
  36257=>"111001010",
  36258=>"000001000",
  36259=>"111000001",
  36260=>"111110101",
  36261=>"101111010",
  36262=>"000010111",
  36263=>"111101011",
  36264=>"101000101",
  36265=>"100110010",
  36266=>"011010000",
  36267=>"011101000",
  36268=>"100001110",
  36269=>"010001000",
  36270=>"111010100",
  36271=>"111100100",
  36272=>"010011100",
  36273=>"100011101",
  36274=>"011101111",
  36275=>"000011001",
  36276=>"010001101",
  36277=>"101010100",
  36278=>"000101101",
  36279=>"101101011",
  36280=>"100011011",
  36281=>"000010100",
  36282=>"001110110",
  36283=>"011010101",
  36284=>"101011111",
  36285=>"101010100",
  36286=>"101111010",
  36287=>"110001100",
  36288=>"010100101",
  36289=>"100100101",
  36290=>"011000101",
  36291=>"010101100",
  36292=>"101111110",
  36293=>"000110000",
  36294=>"001001100",
  36295=>"110010100",
  36296=>"100001001",
  36297=>"111001110",
  36298=>"011011110",
  36299=>"011110010",
  36300=>"001101001",
  36301=>"101111110",
  36302=>"010100110",
  36303=>"101100010",
  36304=>"101110011",
  36305=>"001010000",
  36306=>"101101110",
  36307=>"011010110",
  36308=>"001000010",
  36309=>"101000000",
  36310=>"000000010",
  36311=>"110110001",
  36312=>"100000011",
  36313=>"000100011",
  36314=>"110101111",
  36315=>"001100010",
  36316=>"110000011",
  36317=>"101010011",
  36318=>"011110111",
  36319=>"000110000",
  36320=>"100110010",
  36321=>"101110110",
  36322=>"000100000",
  36323=>"000111110",
  36324=>"100110100",
  36325=>"001000000",
  36326=>"111111111",
  36327=>"100010010",
  36328=>"010010011",
  36329=>"001100010",
  36330=>"011101010",
  36331=>"100000011",
  36332=>"111001011",
  36333=>"100101010",
  36334=>"101000101",
  36335=>"110100100",
  36336=>"000110100",
  36337=>"100110101",
  36338=>"111010100",
  36339=>"110111110",
  36340=>"011000010",
  36341=>"100001111",
  36342=>"101001011",
  36343=>"010101101",
  36344=>"111100010",
  36345=>"010111111",
  36346=>"001110111",
  36347=>"101111010",
  36348=>"011110000",
  36349=>"101001111",
  36350=>"011111011",
  36351=>"101110100",
  36352=>"011001101",
  36353=>"111011001",
  36354=>"011010101",
  36355=>"100101100",
  36356=>"000000010",
  36357=>"100110100",
  36358=>"100100101",
  36359=>"111100001",
  36360=>"011001100",
  36361=>"000110111",
  36362=>"111000000",
  36363=>"011010100",
  36364=>"100000000",
  36365=>"111011100",
  36366=>"111010000",
  36367=>"110111010",
  36368=>"000110101",
  36369=>"000101011",
  36370=>"001101000",
  36371=>"111001010",
  36372=>"111001000",
  36373=>"101010101",
  36374=>"001000010",
  36375=>"111001111",
  36376=>"000010100",
  36377=>"100111011",
  36378=>"010010010",
  36379=>"111100111",
  36380=>"000000001",
  36381=>"001000110",
  36382=>"100011011",
  36383=>"001010010",
  36384=>"101100010",
  36385=>"100110100",
  36386=>"001001001",
  36387=>"111101110",
  36388=>"011101111",
  36389=>"011100111",
  36390=>"111110000",
  36391=>"110001111",
  36392=>"111100101",
  36393=>"111011100",
  36394=>"000101101",
  36395=>"011011111",
  36396=>"000101101",
  36397=>"101101011",
  36398=>"110110101",
  36399=>"000101111",
  36400=>"100010100",
  36401=>"101100100",
  36402=>"100100000",
  36403=>"001011000",
  36404=>"001010111",
  36405=>"111101000",
  36406=>"010010100",
  36407=>"101001001",
  36408=>"010100101",
  36409=>"100011101",
  36410=>"011010010",
  36411=>"111100000",
  36412=>"010100100",
  36413=>"110010001",
  36414=>"111011101",
  36415=>"111011110",
  36416=>"110000000",
  36417=>"111000000",
  36418=>"101101001",
  36419=>"101101010",
  36420=>"111010001",
  36421=>"100010100",
  36422=>"011011000",
  36423=>"100010100",
  36424=>"111010110",
  36425=>"001110011",
  36426=>"111010010",
  36427=>"101100010",
  36428=>"011111000",
  36429=>"100101001",
  36430=>"111010101",
  36431=>"101110011",
  36432=>"011000010",
  36433=>"011000110",
  36434=>"110100110",
  36435=>"011110101",
  36436=>"010000001",
  36437=>"000111001",
  36438=>"000100000",
  36439=>"100001001",
  36440=>"010111111",
  36441=>"101011111",
  36442=>"110100010",
  36443=>"111101110",
  36444=>"111000011",
  36445=>"011101000",
  36446=>"001001001",
  36447=>"101011110",
  36448=>"111111011",
  36449=>"111010100",
  36450=>"010010110",
  36451=>"010000001",
  36452=>"101000000",
  36453=>"001111110",
  36454=>"011010101",
  36455=>"101000100",
  36456=>"110010100",
  36457=>"000101011",
  36458=>"111010000",
  36459=>"111111110",
  36460=>"000100110",
  36461=>"101111100",
  36462=>"110010011",
  36463=>"010100010",
  36464=>"011011100",
  36465=>"001010100",
  36466=>"010110010",
  36467=>"000000100",
  36468=>"111001011",
  36469=>"111110000",
  36470=>"001111000",
  36471=>"110110010",
  36472=>"111000000",
  36473=>"110101110",
  36474=>"101111000",
  36475=>"001001010",
  36476=>"111100001",
  36477=>"111011110",
  36478=>"111111100",
  36479=>"001000011",
  36480=>"101011101",
  36481=>"000111011",
  36482=>"101000110",
  36483=>"000000011",
  36484=>"100111100",
  36485=>"100000001",
  36486=>"011001000",
  36487=>"100001110",
  36488=>"111100111",
  36489=>"010010110",
  36490=>"110110001",
  36491=>"101010001",
  36492=>"100110010",
  36493=>"011011001",
  36494=>"011101011",
  36495=>"100111100",
  36496=>"000000111",
  36497=>"100101101",
  36498=>"011111101",
  36499=>"010100101",
  36500=>"100011100",
  36501=>"010010111",
  36502=>"111010001",
  36503=>"101101111",
  36504=>"000001001",
  36505=>"110001011",
  36506=>"101011011",
  36507=>"000100010",
  36508=>"101010110",
  36509=>"101110110",
  36510=>"111010110",
  36511=>"011110001",
  36512=>"101111100",
  36513=>"101110101",
  36514=>"110000011",
  36515=>"010110001",
  36516=>"100111111",
  36517=>"001001111",
  36518=>"111110110",
  36519=>"001111011",
  36520=>"111000010",
  36521=>"010101000",
  36522=>"100000100",
  36523=>"110100010",
  36524=>"000000001",
  36525=>"110010111",
  36526=>"111000001",
  36527=>"001111010",
  36528=>"110101111",
  36529=>"000000000",
  36530=>"101000111",
  36531=>"101111000",
  36532=>"001100010",
  36533=>"000111001",
  36534=>"001010111",
  36535=>"110100111",
  36536=>"111001111",
  36537=>"101011011",
  36538=>"010010100",
  36539=>"000100000",
  36540=>"000010100",
  36541=>"100011000",
  36542=>"101100000",
  36543=>"011001000",
  36544=>"101111111",
  36545=>"101000001",
  36546=>"100100110",
  36547=>"010000100",
  36548=>"000011001",
  36549=>"001000110",
  36550=>"111101010",
  36551=>"101111111",
  36552=>"111000011",
  36553=>"011000001",
  36554=>"101011111",
  36555=>"010000011",
  36556=>"010010110",
  36557=>"111111111",
  36558=>"000010111",
  36559=>"010111010",
  36560=>"000000111",
  36561=>"111010110",
  36562=>"001111110",
  36563=>"110110101",
  36564=>"110100000",
  36565=>"001000001",
  36566=>"000110100",
  36567=>"000010010",
  36568=>"111110101",
  36569=>"011010111",
  36570=>"010010110",
  36571=>"101011100",
  36572=>"110001011",
  36573=>"110111111",
  36574=>"010111110",
  36575=>"110100011",
  36576=>"001100011",
  36577=>"001111010",
  36578=>"100011111",
  36579=>"011001001",
  36580=>"101001000",
  36581=>"101000110",
  36582=>"101111111",
  36583=>"111000111",
  36584=>"010111101",
  36585=>"101101111",
  36586=>"001000000",
  36587=>"011001011",
  36588=>"111110001",
  36589=>"000101111",
  36590=>"110010000",
  36591=>"100100111",
  36592=>"100000000",
  36593=>"011001100",
  36594=>"101000100",
  36595=>"111010011",
  36596=>"001110101",
  36597=>"000101100",
  36598=>"010101010",
  36599=>"100110000",
  36600=>"100111011",
  36601=>"100010101",
  36602=>"100100111",
  36603=>"000010111",
  36604=>"010011010",
  36605=>"010101000",
  36606=>"111000100",
  36607=>"001001000",
  36608=>"011111010",
  36609=>"010010000",
  36610=>"011001000",
  36611=>"111100111",
  36612=>"011111010",
  36613=>"000000011",
  36614=>"001011111",
  36615=>"100110101",
  36616=>"001111000",
  36617=>"110010000",
  36618=>"111010111",
  36619=>"100100010",
  36620=>"000110001",
  36621=>"000111101",
  36622=>"100010100",
  36623=>"011001100",
  36624=>"100110110",
  36625=>"101101111",
  36626=>"110010100",
  36627=>"000101001",
  36628=>"110011100",
  36629=>"110101011",
  36630=>"000111011",
  36631=>"111001110",
  36632=>"000110011",
  36633=>"010010000",
  36634=>"000000100",
  36635=>"100010011",
  36636=>"011110000",
  36637=>"100011111",
  36638=>"011100100",
  36639=>"011000000",
  36640=>"100101001",
  36641=>"010010011",
  36642=>"111011111",
  36643=>"101001100",
  36644=>"110010110",
  36645=>"110111001",
  36646=>"101101110",
  36647=>"000111101",
  36648=>"111110101",
  36649=>"000000111",
  36650=>"110110001",
  36651=>"101011000",
  36652=>"001111100",
  36653=>"000101010",
  36654=>"010011000",
  36655=>"101001101",
  36656=>"100000000",
  36657=>"100001110",
  36658=>"011010001",
  36659=>"011001000",
  36660=>"111101111",
  36661=>"110000010",
  36662=>"001110110",
  36663=>"001110011",
  36664=>"011110111",
  36665=>"010100111",
  36666=>"010011001",
  36667=>"000001100",
  36668=>"111011000",
  36669=>"101100111",
  36670=>"110000001",
  36671=>"011111111",
  36672=>"100100111",
  36673=>"011000011",
  36674=>"101111010",
  36675=>"010111100",
  36676=>"001101001",
  36677=>"111101101",
  36678=>"010110000",
  36679=>"100111110",
  36680=>"010011100",
  36681=>"100000011",
  36682=>"010011011",
  36683=>"100111101",
  36684=>"101001110",
  36685=>"010000010",
  36686=>"011110100",
  36687=>"111001011",
  36688=>"110110110",
  36689=>"001000101",
  36690=>"000010100",
  36691=>"110011001",
  36692=>"001001000",
  36693=>"000001000",
  36694=>"001110000",
  36695=>"010110001",
  36696=>"101010110",
  36697=>"001111110",
  36698=>"110001011",
  36699=>"111010011",
  36700=>"001010110",
  36701=>"001001001",
  36702=>"111101000",
  36703=>"010000100",
  36704=>"101011100",
  36705=>"100001110",
  36706=>"000111111",
  36707=>"110110010",
  36708=>"111100011",
  36709=>"110011110",
  36710=>"110011010",
  36711=>"011100101",
  36712=>"101101101",
  36713=>"000111110",
  36714=>"001111010",
  36715=>"110001001",
  36716=>"100100000",
  36717=>"010101110",
  36718=>"101010101",
  36719=>"001110010",
  36720=>"111100101",
  36721=>"010011011",
  36722=>"001110111",
  36723=>"111010111",
  36724=>"011101010",
  36725=>"000001010",
  36726=>"010000100",
  36727=>"011101101",
  36728=>"110011000",
  36729=>"000001101",
  36730=>"101111110",
  36731=>"000111001",
  36732=>"100100000",
  36733=>"110011000",
  36734=>"101000100",
  36735=>"000111011",
  36736=>"111110000",
  36737=>"001011010",
  36738=>"000000010",
  36739=>"000010111",
  36740=>"011110000",
  36741=>"110111011",
  36742=>"001001111",
  36743=>"111111100",
  36744=>"001001110",
  36745=>"101101110",
  36746=>"001000100",
  36747=>"000100110",
  36748=>"001101111",
  36749=>"001111100",
  36750=>"001011100",
  36751=>"001110000",
  36752=>"111100100",
  36753=>"010001000",
  36754=>"111001000",
  36755=>"110101110",
  36756=>"111111001",
  36757=>"100110101",
  36758=>"111000010",
  36759=>"000011101",
  36760=>"001100111",
  36761=>"110101000",
  36762=>"111010000",
  36763=>"001000100",
  36764=>"010011000",
  36765=>"011010011",
  36766=>"110000000",
  36767=>"000100000",
  36768=>"011001110",
  36769=>"101111111",
  36770=>"011000100",
  36771=>"000001110",
  36772=>"101001000",
  36773=>"100001100",
  36774=>"000000000",
  36775=>"010010001",
  36776=>"001001001",
  36777=>"110111001",
  36778=>"010000010",
  36779=>"100100111",
  36780=>"011000100",
  36781=>"000110001",
  36782=>"101101010",
  36783=>"101011011",
  36784=>"000001100",
  36785=>"011100100",
  36786=>"000110100",
  36787=>"001010000",
  36788=>"111000011",
  36789=>"011000110",
  36790=>"100101111",
  36791=>"111010101",
  36792=>"001000010",
  36793=>"001000101",
  36794=>"100010101",
  36795=>"000110011",
  36796=>"010111100",
  36797=>"100110100",
  36798=>"111101110",
  36799=>"110111111",
  36800=>"101010100",
  36801=>"000111010",
  36802=>"101010000",
  36803=>"110111110",
  36804=>"100100100",
  36805=>"110100110",
  36806=>"000011111",
  36807=>"001010100",
  36808=>"101001010",
  36809=>"111110001",
  36810=>"010011000",
  36811=>"111111011",
  36812=>"101010010",
  36813=>"011000100",
  36814=>"010000111",
  36815=>"101101101",
  36816=>"000111011",
  36817=>"100011011",
  36818=>"111011101",
  36819=>"100000000",
  36820=>"101000001",
  36821=>"000110111",
  36822=>"010010001",
  36823=>"101100101",
  36824=>"100010110",
  36825=>"100001011",
  36826=>"100011111",
  36827=>"011000010",
  36828=>"101111110",
  36829=>"100110110",
  36830=>"010111110",
  36831=>"000001100",
  36832=>"000111100",
  36833=>"001110101",
  36834=>"001000100",
  36835=>"100010100",
  36836=>"110110100",
  36837=>"110110101",
  36838=>"100010101",
  36839=>"000110100",
  36840=>"000001111",
  36841=>"000100110",
  36842=>"000100100",
  36843=>"011001000",
  36844=>"011000011",
  36845=>"010011111",
  36846=>"000100010",
  36847=>"011000000",
  36848=>"000010000",
  36849=>"111110100",
  36850=>"011011100",
  36851=>"100111010",
  36852=>"100110110",
  36853=>"000010000",
  36854=>"000011100",
  36855=>"010100000",
  36856=>"011011110",
  36857=>"000000101",
  36858=>"100000011",
  36859=>"111001011",
  36860=>"110011001",
  36861=>"100110001",
  36862=>"000000011",
  36863=>"100110010",
  36864=>"101001111",
  36865=>"101110010",
  36866=>"111111100",
  36867=>"001001011",
  36868=>"111110111",
  36869=>"101101111",
  36870=>"001000110",
  36871=>"011011000",
  36872=>"001000000",
  36873=>"111001000",
  36874=>"101011011",
  36875=>"010100100",
  36876=>"111101011",
  36877=>"000010111",
  36878=>"110010000",
  36879=>"010011000",
  36880=>"111111101",
  36881=>"010000111",
  36882=>"100100001",
  36883=>"010010001",
  36884=>"010101000",
  36885=>"101100100",
  36886=>"001001010",
  36887=>"011001010",
  36888=>"001100111",
  36889=>"111011101",
  36890=>"000100010",
  36891=>"110011100",
  36892=>"010111111",
  36893=>"001110111",
  36894=>"110100111",
  36895=>"011110111",
  36896=>"110111101",
  36897=>"100000111",
  36898=>"111100110",
  36899=>"010101100",
  36900=>"011111001",
  36901=>"011001010",
  36902=>"110001000",
  36903=>"000111011",
  36904=>"111100111",
  36905=>"000110100",
  36906=>"111110011",
  36907=>"000101001",
  36908=>"111111101",
  36909=>"001010111",
  36910=>"111100100",
  36911=>"110101010",
  36912=>"010001100",
  36913=>"011010011",
  36914=>"000011001",
  36915=>"111110000",
  36916=>"011101000",
  36917=>"111110110",
  36918=>"010000100",
  36919=>"010000010",
  36920=>"010001001",
  36921=>"010110111",
  36922=>"011011001",
  36923=>"100000011",
  36924=>"001011001",
  36925=>"001000100",
  36926=>"111000110",
  36927=>"001100101",
  36928=>"000011001",
  36929=>"110110001",
  36930=>"010111011",
  36931=>"010001001",
  36932=>"111101000",
  36933=>"100100111",
  36934=>"011001001",
  36935=>"101100001",
  36936=>"011001101",
  36937=>"111110010",
  36938=>"101001110",
  36939=>"001100110",
  36940=>"010000111",
  36941=>"101111001",
  36942=>"111101111",
  36943=>"011010000",
  36944=>"110101001",
  36945=>"011000010",
  36946=>"101110110",
  36947=>"100001010",
  36948=>"001100011",
  36949=>"001101000",
  36950=>"110100011",
  36951=>"010011011",
  36952=>"100001101",
  36953=>"110101000",
  36954=>"001101000",
  36955=>"000100000",
  36956=>"000110111",
  36957=>"000000100",
  36958=>"000001100",
  36959=>"001101111",
  36960=>"011011001",
  36961=>"111010011",
  36962=>"111111001",
  36963=>"111011010",
  36964=>"101100000",
  36965=>"001001101",
  36966=>"111101000",
  36967=>"100100100",
  36968=>"011001000",
  36969=>"000110011",
  36970=>"000111110",
  36971=>"011110100",
  36972=>"001000101",
  36973=>"011011000",
  36974=>"000111011",
  36975=>"111110001",
  36976=>"101111011",
  36977=>"100001000",
  36978=>"000010011",
  36979=>"000011000",
  36980=>"110000100",
  36981=>"010101111",
  36982=>"010001000",
  36983=>"110001011",
  36984=>"000101010",
  36985=>"111101101",
  36986=>"111000011",
  36987=>"111011011",
  36988=>"010110100",
  36989=>"111110101",
  36990=>"000010100",
  36991=>"001110000",
  36992=>"100101100",
  36993=>"100111011",
  36994=>"110110011",
  36995=>"100100001",
  36996=>"010110011",
  36997=>"110001011",
  36998=>"001011010",
  36999=>"011101101",
  37000=>"010100011",
  37001=>"100110010",
  37002=>"111001110",
  37003=>"010111010",
  37004=>"011111001",
  37005=>"100000000",
  37006=>"100100010",
  37007=>"111001100",
  37008=>"111100100",
  37009=>"001001111",
  37010=>"111011010",
  37011=>"110011001",
  37012=>"001101010",
  37013=>"000001101",
  37014=>"111100011",
  37015=>"110010000",
  37016=>"011110110",
  37017=>"111110000",
  37018=>"010001010",
  37019=>"011111101",
  37020=>"101010001",
  37021=>"000010001",
  37022=>"100110001",
  37023=>"011110111",
  37024=>"010101001",
  37025=>"111010001",
  37026=>"010011101",
  37027=>"100100101",
  37028=>"010001100",
  37029=>"110101101",
  37030=>"101001000",
  37031=>"110101101",
  37032=>"110110100",
  37033=>"111000100",
  37034=>"111100100",
  37035=>"110000001",
  37036=>"101001101",
  37037=>"101001111",
  37038=>"011100011",
  37039=>"011001001",
  37040=>"110010001",
  37041=>"111100110",
  37042=>"010100010",
  37043=>"001100000",
  37044=>"111001011",
  37045=>"111111101",
  37046=>"010111011",
  37047=>"001010010",
  37048=>"001011110",
  37049=>"001011011",
  37050=>"001001110",
  37051=>"110000110",
  37052=>"001110101",
  37053=>"011011100",
  37054=>"111111000",
  37055=>"111100001",
  37056=>"001000110",
  37057=>"111011010",
  37058=>"110000101",
  37059=>"110110111",
  37060=>"110011111",
  37061=>"110100001",
  37062=>"001000011",
  37063=>"000000111",
  37064=>"101010111",
  37065=>"000111110",
  37066=>"011000011",
  37067=>"100110000",
  37068=>"010010110",
  37069=>"110110001",
  37070=>"110001110",
  37071=>"001001101",
  37072=>"101001011",
  37073=>"101001011",
  37074=>"011011000",
  37075=>"001111100",
  37076=>"111010100",
  37077=>"001000100",
  37078=>"111011101",
  37079=>"001010010",
  37080=>"000010010",
  37081=>"110101100",
  37082=>"000011000",
  37083=>"011000111",
  37084=>"011110101",
  37085=>"100010111",
  37086=>"011001011",
  37087=>"000010111",
  37088=>"000010011",
  37089=>"011010000",
  37090=>"100111111",
  37091=>"001001110",
  37092=>"100111001",
  37093=>"001110001",
  37094=>"000101011",
  37095=>"111011111",
  37096=>"100010111",
  37097=>"001101001",
  37098=>"101101001",
  37099=>"111001100",
  37100=>"100100010",
  37101=>"000111101",
  37102=>"011101111",
  37103=>"010000001",
  37104=>"111111011",
  37105=>"100111111",
  37106=>"011011010",
  37107=>"100011110",
  37108=>"110011110",
  37109=>"000000110",
  37110=>"000000100",
  37111=>"010000100",
  37112=>"011010011",
  37113=>"111101101",
  37114=>"001011001",
  37115=>"100111010",
  37116=>"111000100",
  37117=>"111110001",
  37118=>"101111111",
  37119=>"010000111",
  37120=>"101001010",
  37121=>"011110101",
  37122=>"100010100",
  37123=>"111010010",
  37124=>"101001000",
  37125=>"011001011",
  37126=>"001100100",
  37127=>"100100100",
  37128=>"000110111",
  37129=>"111000011",
  37130=>"100101101",
  37131=>"100101000",
  37132=>"100110000",
  37133=>"100011101",
  37134=>"110110101",
  37135=>"000001001",
  37136=>"111101000",
  37137=>"011100111",
  37138=>"000101000",
  37139=>"010100000",
  37140=>"100000001",
  37141=>"001000001",
  37142=>"111010000",
  37143=>"111110000",
  37144=>"101110111",
  37145=>"111111111",
  37146=>"000100101",
  37147=>"101101110",
  37148=>"111000110",
  37149=>"010000001",
  37150=>"111000010",
  37151=>"011101000",
  37152=>"100111100",
  37153=>"001110100",
  37154=>"000110100",
  37155=>"101000100",
  37156=>"110101101",
  37157=>"010111000",
  37158=>"011111000",
  37159=>"110100100",
  37160=>"111001001",
  37161=>"000110110",
  37162=>"010000010",
  37163=>"010110001",
  37164=>"111110101",
  37165=>"001000100",
  37166=>"111001110",
  37167=>"010000110",
  37168=>"011011000",
  37169=>"111011101",
  37170=>"000011011",
  37171=>"000000111",
  37172=>"000110000",
  37173=>"001011111",
  37174=>"001000001",
  37175=>"001001001",
  37176=>"101100000",
  37177=>"100110001",
  37178=>"001101010",
  37179=>"001111111",
  37180=>"111011100",
  37181=>"100010011",
  37182=>"111001100",
  37183=>"110111000",
  37184=>"111010101",
  37185=>"000110100",
  37186=>"101010011",
  37187=>"111011001",
  37188=>"111011011",
  37189=>"100111111",
  37190=>"100111101",
  37191=>"011100010",
  37192=>"101010011",
  37193=>"111011011",
  37194=>"001111001",
  37195=>"111101011",
  37196=>"011011110",
  37197=>"111110111",
  37198=>"111111110",
  37199=>"011001000",
  37200=>"101101100",
  37201=>"111011000",
  37202=>"111000111",
  37203=>"010001101",
  37204=>"000111000",
  37205=>"110110010",
  37206=>"110100111",
  37207=>"000010010",
  37208=>"100100001",
  37209=>"000100011",
  37210=>"001110101",
  37211=>"100001111",
  37212=>"100110000",
  37213=>"000010100",
  37214=>"101100100",
  37215=>"000010011",
  37216=>"100011011",
  37217=>"111010100",
  37218=>"100011001",
  37219=>"110100010",
  37220=>"110011000",
  37221=>"011110001",
  37222=>"000101010",
  37223=>"111011000",
  37224=>"110000010",
  37225=>"010011011",
  37226=>"101111010",
  37227=>"100001111",
  37228=>"111110010",
  37229=>"111100001",
  37230=>"011110010",
  37231=>"101100010",
  37232=>"101011000",
  37233=>"010001100",
  37234=>"000011111",
  37235=>"001001001",
  37236=>"000100111",
  37237=>"001001000",
  37238=>"010010000",
  37239=>"010011110",
  37240=>"001000101",
  37241=>"011000000",
  37242=>"100000010",
  37243=>"001110110",
  37244=>"110000000",
  37245=>"111100101",
  37246=>"111101010",
  37247=>"001110110",
  37248=>"011001001",
  37249=>"010011100",
  37250=>"001011111",
  37251=>"101110011",
  37252=>"110101101",
  37253=>"001111101",
  37254=>"010111010",
  37255=>"110011000",
  37256=>"100111100",
  37257=>"110100100",
  37258=>"111101010",
  37259=>"011010010",
  37260=>"001010110",
  37261=>"010000100",
  37262=>"000000101",
  37263=>"011111100",
  37264=>"000000111",
  37265=>"111011000",
  37266=>"111011000",
  37267=>"101001011",
  37268=>"000101001",
  37269=>"011001011",
  37270=>"110000100",
  37271=>"111100010",
  37272=>"001110000",
  37273=>"001001000",
  37274=>"001111101",
  37275=>"111001000",
  37276=>"111000000",
  37277=>"101101000",
  37278=>"011010111",
  37279=>"101001101",
  37280=>"101001100",
  37281=>"111001000",
  37282=>"010111111",
  37283=>"111010110",
  37284=>"110001111",
  37285=>"010110011",
  37286=>"000010110",
  37287=>"110111110",
  37288=>"111100100",
  37289=>"101000010",
  37290=>"010011000",
  37291=>"000111111",
  37292=>"101000111",
  37293=>"011001010",
  37294=>"000001011",
  37295=>"011011010",
  37296=>"010111011",
  37297=>"000001001",
  37298=>"111100001",
  37299=>"100000000",
  37300=>"101101110",
  37301=>"111111101",
  37302=>"000001011",
  37303=>"111100111",
  37304=>"110100000",
  37305=>"101011110",
  37306=>"001011010",
  37307=>"110001101",
  37308=>"110110011",
  37309=>"011000010",
  37310=>"001010101",
  37311=>"100010001",
  37312=>"111110000",
  37313=>"100101001",
  37314=>"110000010",
  37315=>"101100110",
  37316=>"111010001",
  37317=>"000011010",
  37318=>"010011101",
  37319=>"111111001",
  37320=>"110100101",
  37321=>"000110101",
  37322=>"011101000",
  37323=>"111011011",
  37324=>"000010100",
  37325=>"100111101",
  37326=>"000101101",
  37327=>"110100100",
  37328=>"001000011",
  37329=>"010011011",
  37330=>"000100110",
  37331=>"010000011",
  37332=>"000010111",
  37333=>"011000110",
  37334=>"110000110",
  37335=>"111001011",
  37336=>"111110001",
  37337=>"010110110",
  37338=>"011001000",
  37339=>"010111001",
  37340=>"110110010",
  37341=>"011011011",
  37342=>"010110111",
  37343=>"011000100",
  37344=>"011011000",
  37345=>"111101111",
  37346=>"101001010",
  37347=>"010100101",
  37348=>"001000000",
  37349=>"011010000",
  37350=>"010000100",
  37351=>"111101010",
  37352=>"110100110",
  37353=>"000000011",
  37354=>"111001100",
  37355=>"001111111",
  37356=>"000010110",
  37357=>"011111111",
  37358=>"001010000",
  37359=>"001101000",
  37360=>"110101110",
  37361=>"010100111",
  37362=>"001001101",
  37363=>"010100000",
  37364=>"000001000",
  37365=>"000001000",
  37366=>"010000011",
  37367=>"010110100",
  37368=>"111111011",
  37369=>"101011110",
  37370=>"101111101",
  37371=>"110000111",
  37372=>"011110110",
  37373=>"111100110",
  37374=>"000010001",
  37375=>"110110001",
  37376=>"001111110",
  37377=>"101111011",
  37378=>"011111010",
  37379=>"001011000",
  37380=>"100110011",
  37381=>"111000111",
  37382=>"001100001",
  37383=>"100001000",
  37384=>"010011111",
  37385=>"011001010",
  37386=>"000010101",
  37387=>"001110111",
  37388=>"011000011",
  37389=>"010101111",
  37390=>"011001000",
  37391=>"110100110",
  37392=>"111111011",
  37393=>"101001110",
  37394=>"001110101",
  37395=>"010000001",
  37396=>"000111011",
  37397=>"111111111",
  37398=>"001111110",
  37399=>"100100100",
  37400=>"010100000",
  37401=>"011010111",
  37402=>"111010001",
  37403=>"111011010",
  37404=>"101011010",
  37405=>"110001010",
  37406=>"000110100",
  37407=>"101100000",
  37408=>"111011001",
  37409=>"100110000",
  37410=>"100111111",
  37411=>"111110110",
  37412=>"000111010",
  37413=>"001011101",
  37414=>"000110111",
  37415=>"011000110",
  37416=>"101101111",
  37417=>"101011011",
  37418=>"001000000",
  37419=>"100110111",
  37420=>"100011111",
  37421=>"100010000",
  37422=>"000010001",
  37423=>"101111011",
  37424=>"011011101",
  37425=>"001010110",
  37426=>"111101111",
  37427=>"001000010",
  37428=>"100000111",
  37429=>"011001000",
  37430=>"110000000",
  37431=>"100110101",
  37432=>"101100110",
  37433=>"011111100",
  37434=>"001101111",
  37435=>"001100100",
  37436=>"010000100",
  37437=>"110101010",
  37438=>"001101100",
  37439=>"110000101",
  37440=>"111001001",
  37441=>"010111000",
  37442=>"111101010",
  37443=>"101000001",
  37444=>"110100111",
  37445=>"011111011",
  37446=>"010001010",
  37447=>"010110010",
  37448=>"101000000",
  37449=>"001011111",
  37450=>"010110010",
  37451=>"000000001",
  37452=>"000100100",
  37453=>"011111000",
  37454=>"101101011",
  37455=>"010001001",
  37456=>"110100001",
  37457=>"011100001",
  37458=>"000110010",
  37459=>"001010000",
  37460=>"101110100",
  37461=>"010110001",
  37462=>"011111100",
  37463=>"000001000",
  37464=>"011000110",
  37465=>"100101011",
  37466=>"011010100",
  37467=>"101011111",
  37468=>"011101101",
  37469=>"000001000",
  37470=>"101010111",
  37471=>"010010100",
  37472=>"101010101",
  37473=>"111000101",
  37474=>"101010100",
  37475=>"110010010",
  37476=>"110000001",
  37477=>"010011111",
  37478=>"111110101",
  37479=>"101000001",
  37480=>"111111110",
  37481=>"110101000",
  37482=>"010010010",
  37483=>"101101111",
  37484=>"000000111",
  37485=>"110001111",
  37486=>"101100010",
  37487=>"000011101",
  37488=>"101010001",
  37489=>"001111111",
  37490=>"100111101",
  37491=>"110000010",
  37492=>"001001001",
  37493=>"010110000",
  37494=>"111001110",
  37495=>"111001001",
  37496=>"010100101",
  37497=>"001110000",
  37498=>"111100100",
  37499=>"111111111",
  37500=>"101001101",
  37501=>"111001100",
  37502=>"111000101",
  37503=>"011001011",
  37504=>"010010000",
  37505=>"110010100",
  37506=>"111011011",
  37507=>"111101000",
  37508=>"000100100",
  37509=>"110110111",
  37510=>"100110110",
  37511=>"000110001",
  37512=>"001111100",
  37513=>"110000100",
  37514=>"000100101",
  37515=>"001111010",
  37516=>"001111110",
  37517=>"011010001",
  37518=>"101101010",
  37519=>"111011100",
  37520=>"011100110",
  37521=>"001111111",
  37522=>"011111110",
  37523=>"110000001",
  37524=>"000000010",
  37525=>"001011100",
  37526=>"000111010",
  37527=>"110111111",
  37528=>"101010111",
  37529=>"100010010",
  37530=>"000000110",
  37531=>"000000001",
  37532=>"111000000",
  37533=>"111010001",
  37534=>"100100010",
  37535=>"111000000",
  37536=>"001001001",
  37537=>"010100111",
  37538=>"011110111",
  37539=>"101000010",
  37540=>"011001011",
  37541=>"010000010",
  37542=>"000100101",
  37543=>"110101111",
  37544=>"111111001",
  37545=>"011000101",
  37546=>"010111010",
  37547=>"111111001",
  37548=>"000101010",
  37549=>"110111110",
  37550=>"111110101",
  37551=>"110000011",
  37552=>"000001011",
  37553=>"000100011",
  37554=>"010110100",
  37555=>"010111001",
  37556=>"010101001",
  37557=>"111110110",
  37558=>"010010011",
  37559=>"110101100",
  37560=>"110001001",
  37561=>"000100011",
  37562=>"001011101",
  37563=>"001110100",
  37564=>"101010000",
  37565=>"011101000",
  37566=>"010000010",
  37567=>"010111100",
  37568=>"011000000",
  37569=>"111011110",
  37570=>"000011101",
  37571=>"011100011",
  37572=>"100000000",
  37573=>"101101100",
  37574=>"111110101",
  37575=>"110001101",
  37576=>"111111100",
  37577=>"000110001",
  37578=>"100001000",
  37579=>"100011111",
  37580=>"001011101",
  37581=>"101100010",
  37582=>"011011001",
  37583=>"001111101",
  37584=>"110011001",
  37585=>"110110110",
  37586=>"000000001",
  37587=>"001011000",
  37588=>"101111110",
  37589=>"000001010",
  37590=>"100101001",
  37591=>"011000010",
  37592=>"011110111",
  37593=>"101111111",
  37594=>"010101000",
  37595=>"101000010",
  37596=>"010100000",
  37597=>"110100110",
  37598=>"100101100",
  37599=>"000010011",
  37600=>"010000000",
  37601=>"101011100",
  37602=>"110111100",
  37603=>"111101110",
  37604=>"110001110",
  37605=>"111101001",
  37606=>"111010100",
  37607=>"001000101",
  37608=>"001011100",
  37609=>"010100011",
  37610=>"100111101",
  37611=>"110100101",
  37612=>"100110101",
  37613=>"110101000",
  37614=>"011011001",
  37615=>"001000101",
  37616=>"010111110",
  37617=>"101001100",
  37618=>"011100100",
  37619=>"110000100",
  37620=>"100010110",
  37621=>"111110111",
  37622=>"110011100",
  37623=>"101011011",
  37624=>"000010011",
  37625=>"101010001",
  37626=>"100000111",
  37627=>"111000001",
  37628=>"100110001",
  37629=>"011000001",
  37630=>"100111011",
  37631=>"010111010",
  37632=>"110101110",
  37633=>"000111110",
  37634=>"000010010",
  37635=>"111011001",
  37636=>"101101100",
  37637=>"001100011",
  37638=>"000100110",
  37639=>"000010101",
  37640=>"110110001",
  37641=>"101100101",
  37642=>"110100001",
  37643=>"111111000",
  37644=>"011000100",
  37645=>"111100110",
  37646=>"101110101",
  37647=>"011101100",
  37648=>"110010000",
  37649=>"111011000",
  37650=>"110101111",
  37651=>"000000100",
  37652=>"110001110",
  37653=>"011000110",
  37654=>"110101111",
  37655=>"011000011",
  37656=>"111001111",
  37657=>"011000101",
  37658=>"000000000",
  37659=>"010001111",
  37660=>"100101010",
  37661=>"100010100",
  37662=>"101011010",
  37663=>"011111001",
  37664=>"000011100",
  37665=>"011111011",
  37666=>"111000101",
  37667=>"011000010",
  37668=>"100000001",
  37669=>"011100001",
  37670=>"101001101",
  37671=>"110111010",
  37672=>"101001010",
  37673=>"101011001",
  37674=>"110111111",
  37675=>"000110110",
  37676=>"100111101",
  37677=>"000000001",
  37678=>"101010001",
  37679=>"111011101",
  37680=>"110011000",
  37681=>"101000111",
  37682=>"100111000",
  37683=>"001010000",
  37684=>"111101111",
  37685=>"111011101",
  37686=>"001100111",
  37687=>"001100110",
  37688=>"101111111",
  37689=>"011100001",
  37690=>"110100011",
  37691=>"110010001",
  37692=>"100000000",
  37693=>"111000001",
  37694=>"101011100",
  37695=>"000000111",
  37696=>"110000111",
  37697=>"010100111",
  37698=>"000110001",
  37699=>"100000000",
  37700=>"001111000",
  37701=>"001110010",
  37702=>"110001100",
  37703=>"101000001",
  37704=>"010000010",
  37705=>"001011100",
  37706=>"000100011",
  37707=>"010111001",
  37708=>"101011010",
  37709=>"011001011",
  37710=>"101000000",
  37711=>"000101010",
  37712=>"111000100",
  37713=>"100010101",
  37714=>"111010001",
  37715=>"010000000",
  37716=>"001111000",
  37717=>"000001100",
  37718=>"010111101",
  37719=>"100110000",
  37720=>"000111111",
  37721=>"111110011",
  37722=>"101100100",
  37723=>"110001011",
  37724=>"011101111",
  37725=>"001000011",
  37726=>"111011011",
  37727=>"101001001",
  37728=>"111011000",
  37729=>"111111100",
  37730=>"001000101",
  37731=>"101100110",
  37732=>"101011001",
  37733=>"010101010",
  37734=>"110000111",
  37735=>"000010100",
  37736=>"111110110",
  37737=>"001010110",
  37738=>"010010000",
  37739=>"110111010",
  37740=>"100100111",
  37741=>"010011001",
  37742=>"111100001",
  37743=>"111001100",
  37744=>"100001101",
  37745=>"101100101",
  37746=>"101101111",
  37747=>"111110110",
  37748=>"110001101",
  37749=>"011000010",
  37750=>"111101100",
  37751=>"110011011",
  37752=>"001010001",
  37753=>"010100101",
  37754=>"001101100",
  37755=>"111001011",
  37756=>"010001000",
  37757=>"110101011",
  37758=>"111100110",
  37759=>"011001001",
  37760=>"110111110",
  37761=>"001001000",
  37762=>"000100100",
  37763=>"000000011",
  37764=>"011001000",
  37765=>"111101111",
  37766=>"010000101",
  37767=>"011001111",
  37768=>"011010100",
  37769=>"010110101",
  37770=>"011000100",
  37771=>"010111011",
  37772=>"101011000",
  37773=>"001111111",
  37774=>"011110110",
  37775=>"101100101",
  37776=>"000100010",
  37777=>"110011011",
  37778=>"111001000",
  37779=>"110101101",
  37780=>"011000010",
  37781=>"000100111",
  37782=>"001001011",
  37783=>"000101111",
  37784=>"111101101",
  37785=>"111101001",
  37786=>"000101100",
  37787=>"011011011",
  37788=>"111000101",
  37789=>"110110010",
  37790=>"011001010",
  37791=>"101111100",
  37792=>"000110110",
  37793=>"011011111",
  37794=>"011101000",
  37795=>"111100010",
  37796=>"010011001",
  37797=>"000010001",
  37798=>"100100010",
  37799=>"100011001",
  37800=>"000100101",
  37801=>"011000100",
  37802=>"100100110",
  37803=>"110111111",
  37804=>"010011011",
  37805=>"011100100",
  37806=>"001101111",
  37807=>"011000001",
  37808=>"111111111",
  37809=>"110000010",
  37810=>"110101001",
  37811=>"110111101",
  37812=>"010001000",
  37813=>"101101111",
  37814=>"100111110",
  37815=>"100001001",
  37816=>"110111101",
  37817=>"100000110",
  37818=>"010010011",
  37819=>"111101110",
  37820=>"001111001",
  37821=>"101001000",
  37822=>"110111110",
  37823=>"001001011",
  37824=>"010011011",
  37825=>"100000101",
  37826=>"110110111",
  37827=>"110000000",
  37828=>"000001111",
  37829=>"010101001",
  37830=>"100010100",
  37831=>"000000010",
  37832=>"111100100",
  37833=>"111101111",
  37834=>"100101010",
  37835=>"011110001",
  37836=>"000110111",
  37837=>"101001100",
  37838=>"111101010",
  37839=>"100100001",
  37840=>"010000010",
  37841=>"011000110",
  37842=>"000001011",
  37843=>"011001100",
  37844=>"110101010",
  37845=>"110001101",
  37846=>"000110110",
  37847=>"000110111",
  37848=>"101100001",
  37849=>"101000000",
  37850=>"101011111",
  37851=>"100101101",
  37852=>"000101100",
  37853=>"010011111",
  37854=>"100001100",
  37855=>"111000110",
  37856=>"011110000",
  37857=>"101110101",
  37858=>"101011101",
  37859=>"011111011",
  37860=>"011011001",
  37861=>"001110010",
  37862=>"010001001",
  37863=>"110110011",
  37864=>"001111100",
  37865=>"101111000",
  37866=>"010101000",
  37867=>"000010001",
  37868=>"000100100",
  37869=>"000111100",
  37870=>"111011110",
  37871=>"111101100",
  37872=>"110101010",
  37873=>"111000001",
  37874=>"010100000",
  37875=>"011110111",
  37876=>"010011010",
  37877=>"011111000",
  37878=>"000000100",
  37879=>"010100011",
  37880=>"011000000",
  37881=>"101001100",
  37882=>"000011110",
  37883=>"011001110",
  37884=>"010000001",
  37885=>"000000101",
  37886=>"001000101",
  37887=>"010000001",
  37888=>"111100011",
  37889=>"000010100",
  37890=>"001110110",
  37891=>"001001111",
  37892=>"010110111",
  37893=>"011011110",
  37894=>"011110000",
  37895=>"111111111",
  37896=>"111110101",
  37897=>"111100101",
  37898=>"100001111",
  37899=>"000000111",
  37900=>"111111010",
  37901=>"000101001",
  37902=>"001101011",
  37903=>"000010001",
  37904=>"000000000",
  37905=>"001001100",
  37906=>"111101001",
  37907=>"010011101",
  37908=>"000011000",
  37909=>"111111101",
  37910=>"100010000",
  37911=>"110111101",
  37912=>"101001110",
  37913=>"001001111",
  37914=>"111010010",
  37915=>"011111101",
  37916=>"001000010",
  37917=>"001111111",
  37918=>"110000101",
  37919=>"111001100",
  37920=>"000111011",
  37921=>"100110100",
  37922=>"110000100",
  37923=>"101001111",
  37924=>"001001001",
  37925=>"111111011",
  37926=>"010010000",
  37927=>"010101111",
  37928=>"010000000",
  37929=>"101011011",
  37930=>"101001011",
  37931=>"000110010",
  37932=>"010000001",
  37933=>"011000110",
  37934=>"100000111",
  37935=>"110000011",
  37936=>"101100101",
  37937=>"100010001",
  37938=>"000110000",
  37939=>"011011100",
  37940=>"001101000",
  37941=>"101011000",
  37942=>"111100000",
  37943=>"000001101",
  37944=>"100001111",
  37945=>"000001010",
  37946=>"101110000",
  37947=>"001010110",
  37948=>"111000010",
  37949=>"000001010",
  37950=>"101001101",
  37951=>"001111011",
  37952=>"111101011",
  37953=>"001001000",
  37954=>"001000110",
  37955=>"000010111",
  37956=>"100101001",
  37957=>"011000000",
  37958=>"000101101",
  37959=>"010001100",
  37960=>"110001010",
  37961=>"010110011",
  37962=>"001101010",
  37963=>"000100010",
  37964=>"001000010",
  37965=>"001100101",
  37966=>"010100010",
  37967=>"001001000",
  37968=>"100010110",
  37969=>"011110001",
  37970=>"001011001",
  37971=>"001100101",
  37972=>"101110001",
  37973=>"110110010",
  37974=>"100001011",
  37975=>"011000100",
  37976=>"111111100",
  37977=>"100011001",
  37978=>"101000001",
  37979=>"101001110",
  37980=>"101001101",
  37981=>"111101011",
  37982=>"000101101",
  37983=>"110001111",
  37984=>"000000111",
  37985=>"011000100",
  37986=>"011110000",
  37987=>"000000011",
  37988=>"010100110",
  37989=>"100010111",
  37990=>"000010101",
  37991=>"100000100",
  37992=>"100001011",
  37993=>"001001010",
  37994=>"111000111",
  37995=>"110000111",
  37996=>"100111010",
  37997=>"101011111",
  37998=>"100100111",
  37999=>"000100011",
  38000=>"111111010",
  38001=>"100101010",
  38002=>"011110011",
  38003=>"110100000",
  38004=>"011000101",
  38005=>"000111111",
  38006=>"010110000",
  38007=>"110110101",
  38008=>"001110001",
  38009=>"110110011",
  38010=>"110111010",
  38011=>"111010011",
  38012=>"000001001",
  38013=>"111100100",
  38014=>"011100100",
  38015=>"010101111",
  38016=>"110111111",
  38017=>"000111010",
  38018=>"111010011",
  38019=>"111000011",
  38020=>"111111100",
  38021=>"100101101",
  38022=>"100010110",
  38023=>"010010010",
  38024=>"110000001",
  38025=>"011011110",
  38026=>"110100100",
  38027=>"010010011",
  38028=>"001111101",
  38029=>"010110100",
  38030=>"000000110",
  38031=>"111000110",
  38032=>"100000011",
  38033=>"110110001",
  38034=>"100100110",
  38035=>"011010001",
  38036=>"010100100",
  38037=>"000000001",
  38038=>"110111101",
  38039=>"111001000",
  38040=>"111100011",
  38041=>"011011101",
  38042=>"011010011",
  38043=>"000001110",
  38044=>"000110110",
  38045=>"010100101",
  38046=>"011010000",
  38047=>"000000011",
  38048=>"101100011",
  38049=>"001001110",
  38050=>"110010011",
  38051=>"111010011",
  38052=>"110100111",
  38053=>"000000101",
  38054=>"010000110",
  38055=>"111111100",
  38056=>"001100110",
  38057=>"101111001",
  38058=>"100100101",
  38059=>"010010011",
  38060=>"000000000",
  38061=>"111100101",
  38062=>"011001011",
  38063=>"111011001",
  38064=>"000101110",
  38065=>"010110100",
  38066=>"000110101",
  38067=>"000010011",
  38068=>"000001101",
  38069=>"111100000",
  38070=>"110101101",
  38071=>"011110001",
  38072=>"111100101",
  38073=>"010110100",
  38074=>"011100110",
  38075=>"110111010",
  38076=>"111111000",
  38077=>"001011001",
  38078=>"001101111",
  38079=>"100100100",
  38080=>"100001011",
  38081=>"110100011",
  38082=>"010110110",
  38083=>"110101011",
  38084=>"001111111",
  38085=>"001100110",
  38086=>"000001100",
  38087=>"000110011",
  38088=>"001011100",
  38089=>"101010010",
  38090=>"000001110",
  38091=>"010001110",
  38092=>"000001001",
  38093=>"011111000",
  38094=>"010100110",
  38095=>"011000100",
  38096=>"111100010",
  38097=>"110000011",
  38098=>"011111110",
  38099=>"001011001",
  38100=>"111100000",
  38101=>"000111101",
  38102=>"011100001",
  38103=>"100001100",
  38104=>"101011001",
  38105=>"111000011",
  38106=>"000011101",
  38107=>"111000111",
  38108=>"110111010",
  38109=>"101010101",
  38110=>"011101110",
  38111=>"011100101",
  38112=>"100000001",
  38113=>"011011111",
  38114=>"100100000",
  38115=>"001000000",
  38116=>"001111110",
  38117=>"000101110",
  38118=>"011000000",
  38119=>"111011110",
  38120=>"001000101",
  38121=>"110000011",
  38122=>"010011011",
  38123=>"000111110",
  38124=>"000110010",
  38125=>"001101110",
  38126=>"000101011",
  38127=>"000000100",
  38128=>"100001100",
  38129=>"100110000",
  38130=>"110111010",
  38131=>"010101011",
  38132=>"110010011",
  38133=>"110011011",
  38134=>"010000111",
  38135=>"100101111",
  38136=>"111011010",
  38137=>"100000001",
  38138=>"110011101",
  38139=>"000001010",
  38140=>"101011101",
  38141=>"110010101",
  38142=>"010101100",
  38143=>"011111101",
  38144=>"011001110",
  38145=>"100111000",
  38146=>"000010110",
  38147=>"100001000",
  38148=>"011110111",
  38149=>"111100000",
  38150=>"101000101",
  38151=>"000101000",
  38152=>"001111100",
  38153=>"100011101",
  38154=>"000101101",
  38155=>"110010011",
  38156=>"101000001",
  38157=>"000000101",
  38158=>"111000010",
  38159=>"101010111",
  38160=>"110101001",
  38161=>"111111000",
  38162=>"100010110",
  38163=>"011011001",
  38164=>"111101101",
  38165=>"010110110",
  38166=>"101110111",
  38167=>"000110111",
  38168=>"101100101",
  38169=>"010011000",
  38170=>"000011011",
  38171=>"010100111",
  38172=>"110111101",
  38173=>"000111010",
  38174=>"111000100",
  38175=>"110111101",
  38176=>"001100101",
  38177=>"000100000",
  38178=>"010110001",
  38179=>"110100101",
  38180=>"101010001",
  38181=>"000111011",
  38182=>"011011100",
  38183=>"011000011",
  38184=>"101010000",
  38185=>"110100111",
  38186=>"100010101",
  38187=>"101001100",
  38188=>"111011010",
  38189=>"111000100",
  38190=>"101110000",
  38191=>"001100101",
  38192=>"010101011",
  38193=>"100100100",
  38194=>"111011101",
  38195=>"110101011",
  38196=>"111111000",
  38197=>"010110000",
  38198=>"001100011",
  38199=>"110110011",
  38200=>"010010000",
  38201=>"110111011",
  38202=>"000000100",
  38203=>"100100000",
  38204=>"111011000",
  38205=>"000010010",
  38206=>"110001010",
  38207=>"010100001",
  38208=>"001110000",
  38209=>"000111111",
  38210=>"101011000",
  38211=>"010010010",
  38212=>"000101111",
  38213=>"101011010",
  38214=>"101110010",
  38215=>"011000001",
  38216=>"101000010",
  38217=>"010110010",
  38218=>"111101110",
  38219=>"110010101",
  38220=>"111111111",
  38221=>"010001001",
  38222=>"010011110",
  38223=>"001000110",
  38224=>"111001001",
  38225=>"010011010",
  38226=>"010111011",
  38227=>"000101011",
  38228=>"100100100",
  38229=>"111100111",
  38230=>"010001010",
  38231=>"110010011",
  38232=>"011101111",
  38233=>"000111001",
  38234=>"111010000",
  38235=>"100100001",
  38236=>"111001110",
  38237=>"011010100",
  38238=>"000010110",
  38239=>"110010100",
  38240=>"111001101",
  38241=>"101100011",
  38242=>"111110000",
  38243=>"000011100",
  38244=>"001001101",
  38245=>"101010010",
  38246=>"000101011",
  38247=>"001011111",
  38248=>"001000110",
  38249=>"001110010",
  38250=>"110010010",
  38251=>"100110111",
  38252=>"110001000",
  38253=>"000001100",
  38254=>"001100101",
  38255=>"001101001",
  38256=>"001100110",
  38257=>"011010011",
  38258=>"100100000",
  38259=>"111011001",
  38260=>"011110001",
  38261=>"000010001",
  38262=>"010100011",
  38263=>"100111000",
  38264=>"111011111",
  38265=>"000001011",
  38266=>"001010011",
  38267=>"101111000",
  38268=>"100101111",
  38269=>"011001001",
  38270=>"000111101",
  38271=>"000110000",
  38272=>"000000011",
  38273=>"110000010",
  38274=>"110100110",
  38275=>"000111100",
  38276=>"001100011",
  38277=>"110110100",
  38278=>"000010100",
  38279=>"010000000",
  38280=>"000110010",
  38281=>"100110011",
  38282=>"110111000",
  38283=>"100010010",
  38284=>"001010000",
  38285=>"110101111",
  38286=>"111110010",
  38287=>"101001001",
  38288=>"010111011",
  38289=>"111100000",
  38290=>"100010101",
  38291=>"100001111",
  38292=>"010110111",
  38293=>"001001001",
  38294=>"101101111",
  38295=>"111001001",
  38296=>"110111111",
  38297=>"000010111",
  38298=>"001011001",
  38299=>"011111001",
  38300=>"110100100",
  38301=>"101111101",
  38302=>"100110101",
  38303=>"001100111",
  38304=>"110101100",
  38305=>"100001100",
  38306=>"101100101",
  38307=>"110010111",
  38308=>"101111001",
  38309=>"111011010",
  38310=>"010100001",
  38311=>"000111110",
  38312=>"010100111",
  38313=>"010000110",
  38314=>"011101010",
  38315=>"101000010",
  38316=>"000000110",
  38317=>"110010010",
  38318=>"000100101",
  38319=>"011000010",
  38320=>"000101111",
  38321=>"110000011",
  38322=>"110110000",
  38323=>"110110011",
  38324=>"101011111",
  38325=>"001010000",
  38326=>"110011000",
  38327=>"001101111",
  38328=>"000010010",
  38329=>"100100100",
  38330=>"101100100",
  38331=>"011010011",
  38332=>"111100010",
  38333=>"010100101",
  38334=>"110000100",
  38335=>"111111001",
  38336=>"111111010",
  38337=>"000000111",
  38338=>"100001000",
  38339=>"101101111",
  38340=>"010101010",
  38341=>"111001000",
  38342=>"110011001",
  38343=>"011100100",
  38344=>"100101000",
  38345=>"001001101",
  38346=>"000010101",
  38347=>"101110111",
  38348=>"010110001",
  38349=>"010101011",
  38350=>"110100111",
  38351=>"011000010",
  38352=>"001110111",
  38353=>"010011011",
  38354=>"001110100",
  38355=>"011010101",
  38356=>"100010101",
  38357=>"000111010",
  38358=>"100111111",
  38359=>"111111011",
  38360=>"000111001",
  38361=>"011001100",
  38362=>"100001010",
  38363=>"111100001",
  38364=>"100101010",
  38365=>"011101111",
  38366=>"011000001",
  38367=>"000101110",
  38368=>"001100111",
  38369=>"000011100",
  38370=>"010000110",
  38371=>"001111111",
  38372=>"001110110",
  38373=>"111110101",
  38374=>"001110010",
  38375=>"010011000",
  38376=>"111100011",
  38377=>"000010010",
  38378=>"101100000",
  38379=>"111011110",
  38380=>"000000000",
  38381=>"111001000",
  38382=>"000100000",
  38383=>"000010010",
  38384=>"000001000",
  38385=>"100100001",
  38386=>"110000101",
  38387=>"111111000",
  38388=>"010010001",
  38389=>"010101011",
  38390=>"000011111",
  38391=>"110011000",
  38392=>"101111110",
  38393=>"111101010",
  38394=>"101000000",
  38395=>"001100101",
  38396=>"010111110",
  38397=>"111101111",
  38398=>"000111001",
  38399=>"011001111",
  38400=>"000001100",
  38401=>"110000110",
  38402=>"000010010",
  38403=>"110101001",
  38404=>"000010100",
  38405=>"000000101",
  38406=>"100100110",
  38407=>"010001111",
  38408=>"110110110",
  38409=>"101100111",
  38410=>"111000111",
  38411=>"100111110",
  38412=>"111010101",
  38413=>"111111011",
  38414=>"110001010",
  38415=>"100101110",
  38416=>"010011101",
  38417=>"111001101",
  38418=>"111001010",
  38419=>"111110110",
  38420=>"111000000",
  38421=>"100011011",
  38422=>"010010010",
  38423=>"100000110",
  38424=>"001011101",
  38425=>"110010000",
  38426=>"101110001",
  38427=>"011011001",
  38428=>"111000110",
  38429=>"110100101",
  38430=>"000101111",
  38431=>"011111100",
  38432=>"111111111",
  38433=>"001001010",
  38434=>"101000000",
  38435=>"010111011",
  38436=>"101000000",
  38437=>"010001000",
  38438=>"111110011",
  38439=>"110011000",
  38440=>"001100000",
  38441=>"100000100",
  38442=>"100100011",
  38443=>"101010110",
  38444=>"111010111",
  38445=>"101100011",
  38446=>"100100111",
  38447=>"101000101",
  38448=>"001111110",
  38449=>"100010010",
  38450=>"101101001",
  38451=>"111011100",
  38452=>"110110110",
  38453=>"010101001",
  38454=>"000011010",
  38455=>"111011010",
  38456=>"101111100",
  38457=>"110010100",
  38458=>"100001001",
  38459=>"111100100",
  38460=>"000110001",
  38461=>"111110111",
  38462=>"110011010",
  38463=>"100110010",
  38464=>"010100101",
  38465=>"001101101",
  38466=>"100110110",
  38467=>"011010111",
  38468=>"100000000",
  38469=>"110001001",
  38470=>"110000101",
  38471=>"011101110",
  38472=>"010010000",
  38473=>"000110110",
  38474=>"101100000",
  38475=>"000101000",
  38476=>"101000001",
  38477=>"010101001",
  38478=>"110111100",
  38479=>"110010111",
  38480=>"011100001",
  38481=>"101110011",
  38482=>"110101000",
  38483=>"001100001",
  38484=>"001100000",
  38485=>"000010011",
  38486=>"111000101",
  38487=>"001001101",
  38488=>"010000100",
  38489=>"011101110",
  38490=>"100011010",
  38491=>"000101111",
  38492=>"110011000",
  38493=>"011010111",
  38494=>"000000110",
  38495=>"001001110",
  38496=>"010110010",
  38497=>"110010011",
  38498=>"000111010",
  38499=>"101111000",
  38500=>"100111110",
  38501=>"011101111",
  38502=>"101100111",
  38503=>"001100100",
  38504=>"111001110",
  38505=>"111001101",
  38506=>"111000010",
  38507=>"010000001",
  38508=>"000011110",
  38509=>"010010100",
  38510=>"111011101",
  38511=>"000110001",
  38512=>"001011010",
  38513=>"011110101",
  38514=>"010101011",
  38515=>"001000001",
  38516=>"111001110",
  38517=>"100101000",
  38518=>"111101110",
  38519=>"111000010",
  38520=>"110110111",
  38521=>"110110100",
  38522=>"111100011",
  38523=>"110101100",
  38524=>"000001101",
  38525=>"111110011",
  38526=>"101110011",
  38527=>"010000100",
  38528=>"000110011",
  38529=>"101001111",
  38530=>"111111111",
  38531=>"000001101",
  38532=>"100101101",
  38533=>"011010010",
  38534=>"001001110",
  38535=>"000101101",
  38536=>"011001101",
  38537=>"010101000",
  38538=>"000011110",
  38539=>"000111111",
  38540=>"110111101",
  38541=>"110011000",
  38542=>"011001000",
  38543=>"000011000",
  38544=>"101010000",
  38545=>"111110000",
  38546=>"111001100",
  38547=>"001001101",
  38548=>"000001101",
  38549=>"111001111",
  38550=>"011110100",
  38551=>"000001001",
  38552=>"100111101",
  38553=>"001110111",
  38554=>"101010010",
  38555=>"011011001",
  38556=>"111101000",
  38557=>"010110111",
  38558=>"100000011",
  38559=>"110111011",
  38560=>"010111110",
  38561=>"010111000",
  38562=>"001101010",
  38563=>"100101101",
  38564=>"101011101",
  38565=>"011111001",
  38566=>"101001000",
  38567=>"000110101",
  38568=>"000000011",
  38569=>"010001010",
  38570=>"110001100",
  38571=>"011101100",
  38572=>"000001001",
  38573=>"000100100",
  38574=>"101100111",
  38575=>"111111110",
  38576=>"100011111",
  38577=>"011000101",
  38578=>"010000001",
  38579=>"011110001",
  38580=>"101000011",
  38581=>"111010001",
  38582=>"111101011",
  38583=>"001101110",
  38584=>"101011100",
  38585=>"010100000",
  38586=>"000111011",
  38587=>"000111101",
  38588=>"101000111",
  38589=>"101010101",
  38590=>"110010101",
  38591=>"011110010",
  38592=>"110000111",
  38593=>"010111001",
  38594=>"010111101",
  38595=>"100111000",
  38596=>"000001101",
  38597=>"001010000",
  38598=>"111011001",
  38599=>"010100110",
  38600=>"111111110",
  38601=>"010010101",
  38602=>"110111001",
  38603=>"110100001",
  38604=>"011001101",
  38605=>"001110000",
  38606=>"100110110",
  38607=>"000001011",
  38608=>"111110011",
  38609=>"000000100",
  38610=>"110000101",
  38611=>"110110110",
  38612=>"101110010",
  38613=>"111110000",
  38614=>"001110111",
  38615=>"001001100",
  38616=>"110000101",
  38617=>"001100011",
  38618=>"000000010",
  38619=>"101010000",
  38620=>"110000001",
  38621=>"010111110",
  38622=>"010111111",
  38623=>"101101001",
  38624=>"110100010",
  38625=>"111101101",
  38626=>"010010000",
  38627=>"101110001",
  38628=>"100100111",
  38629=>"101011110",
  38630=>"111010101",
  38631=>"010100001",
  38632=>"111000001",
  38633=>"101101001",
  38634=>"000011000",
  38635=>"111100011",
  38636=>"010011011",
  38637=>"000101110",
  38638=>"101000111",
  38639=>"001111010",
  38640=>"111111000",
  38641=>"101111011",
  38642=>"100000000",
  38643=>"001000010",
  38644=>"010110000",
  38645=>"110111000",
  38646=>"110111001",
  38647=>"111111010",
  38648=>"111011100",
  38649=>"011000110",
  38650=>"100011111",
  38651=>"110100101",
  38652=>"011001011",
  38653=>"001010111",
  38654=>"110000000",
  38655=>"001011101",
  38656=>"000010101",
  38657=>"111110011",
  38658=>"001110011",
  38659=>"010100101",
  38660=>"011111000",
  38661=>"111101110",
  38662=>"001101101",
  38663=>"001101101",
  38664=>"100000100",
  38665=>"011010010",
  38666=>"111110010",
  38667=>"110100110",
  38668=>"110010010",
  38669=>"000101101",
  38670=>"100011101",
  38671=>"101001010",
  38672=>"110111110",
  38673=>"110011011",
  38674=>"011110011",
  38675=>"101001101",
  38676=>"110111110",
  38677=>"000100001",
  38678=>"011101010",
  38679=>"010100101",
  38680=>"110001100",
  38681=>"101010111",
  38682=>"101110100",
  38683=>"100100000",
  38684=>"011100000",
  38685=>"100101011",
  38686=>"011010000",
  38687=>"110011000",
  38688=>"000111001",
  38689=>"111001100",
  38690=>"111001000",
  38691=>"001011101",
  38692=>"000000100",
  38693=>"010010000",
  38694=>"110011101",
  38695=>"010000101",
  38696=>"000101010",
  38697=>"111000101",
  38698=>"100010000",
  38699=>"001011101",
  38700=>"000110001",
  38701=>"100000100",
  38702=>"011101001",
  38703=>"111000010",
  38704=>"101111101",
  38705=>"000000010",
  38706=>"101000000",
  38707=>"110100111",
  38708=>"000101011",
  38709=>"111111101",
  38710=>"110101100",
  38711=>"011111010",
  38712=>"101011010",
  38713=>"000011110",
  38714=>"111110110",
  38715=>"010010011",
  38716=>"100101011",
  38717=>"111100010",
  38718=>"101001010",
  38719=>"100110011",
  38720=>"100100000",
  38721=>"111100111",
  38722=>"010100111",
  38723=>"111011110",
  38724=>"100111110",
  38725=>"111010111",
  38726=>"110110000",
  38727=>"011111111",
  38728=>"101000000",
  38729=>"011010000",
  38730=>"010110001",
  38731=>"000000100",
  38732=>"011000101",
  38733=>"011000110",
  38734=>"111001000",
  38735=>"000101010",
  38736=>"100000010",
  38737=>"001011100",
  38738=>"110101001",
  38739=>"011101110",
  38740=>"001100110",
  38741=>"110101100",
  38742=>"000011101",
  38743=>"101100011",
  38744=>"000011100",
  38745=>"100111000",
  38746=>"100101001",
  38747=>"010111100",
  38748=>"111110011",
  38749=>"100100101",
  38750=>"111011011",
  38751=>"011101000",
  38752=>"111100111",
  38753=>"111000100",
  38754=>"111011010",
  38755=>"000001110",
  38756=>"000100000",
  38757=>"000100111",
  38758=>"101101001",
  38759=>"000000100",
  38760=>"101110010",
  38761=>"100110111",
  38762=>"011110110",
  38763=>"101101101",
  38764=>"011011111",
  38765=>"111100000",
  38766=>"011100001",
  38767=>"001001111",
  38768=>"011111110",
  38769=>"010000000",
  38770=>"101011010",
  38771=>"101110010",
  38772=>"100110011",
  38773=>"001010111",
  38774=>"010110000",
  38775=>"101000110",
  38776=>"001010011",
  38777=>"011001100",
  38778=>"001100010",
  38779=>"100110111",
  38780=>"111100000",
  38781=>"110000010",
  38782=>"010000000",
  38783=>"101101011",
  38784=>"000100010",
  38785=>"010100101",
  38786=>"010000100",
  38787=>"100011010",
  38788=>"001011111",
  38789=>"000011000",
  38790=>"110001000",
  38791=>"010110100",
  38792=>"001000001",
  38793=>"000001100",
  38794=>"000000010",
  38795=>"100110011",
  38796=>"101100111",
  38797=>"001111111",
  38798=>"111010100",
  38799=>"010100100",
  38800=>"010111000",
  38801=>"110110011",
  38802=>"100100100",
  38803=>"110000111",
  38804=>"101110101",
  38805=>"010111000",
  38806=>"110010110",
  38807=>"010110000",
  38808=>"101100011",
  38809=>"101100000",
  38810=>"000110111",
  38811=>"100100010",
  38812=>"110111011",
  38813=>"111100010",
  38814=>"010001001",
  38815=>"000110100",
  38816=>"001101100",
  38817=>"000011111",
  38818=>"001110000",
  38819=>"000110100",
  38820=>"100100110",
  38821=>"101100101",
  38822=>"100100101",
  38823=>"010101101",
  38824=>"001011000",
  38825=>"010000111",
  38826=>"001011100",
  38827=>"010100100",
  38828=>"000010001",
  38829=>"111001011",
  38830=>"001111101",
  38831=>"110110000",
  38832=>"010000111",
  38833=>"100111100",
  38834=>"011010000",
  38835=>"100011100",
  38836=>"100101011",
  38837=>"101100011",
  38838=>"000011111",
  38839=>"001100110",
  38840=>"011011100",
  38841=>"010110000",
  38842=>"110001110",
  38843=>"110101111",
  38844=>"110011110",
  38845=>"111101001",
  38846=>"111110111",
  38847=>"111101100",
  38848=>"001100010",
  38849=>"100100111",
  38850=>"010010000",
  38851=>"010101011",
  38852=>"010111001",
  38853=>"001001111",
  38854=>"111011100",
  38855=>"011111110",
  38856=>"111101101",
  38857=>"000100101",
  38858=>"110111100",
  38859=>"000001110",
  38860=>"000000100",
  38861=>"010010000",
  38862=>"000111111",
  38863=>"110110001",
  38864=>"111000110",
  38865=>"111110001",
  38866=>"101000100",
  38867=>"011100101",
  38868=>"001100111",
  38869=>"110111001",
  38870=>"101100000",
  38871=>"011101110",
  38872=>"000001011",
  38873=>"101111010",
  38874=>"011100001",
  38875=>"011100110",
  38876=>"110010000",
  38877=>"011001100",
  38878=>"010000110",
  38879=>"101001000",
  38880=>"011111100",
  38881=>"000001000",
  38882=>"101000110",
  38883=>"011100110",
  38884=>"101101100",
  38885=>"101110100",
  38886=>"111000101",
  38887=>"001011100",
  38888=>"001000100",
  38889=>"110011110",
  38890=>"110011010",
  38891=>"110011011",
  38892=>"110110111",
  38893=>"011100010",
  38894=>"010011011",
  38895=>"100100111",
  38896=>"110100110",
  38897=>"001111100",
  38898=>"000001111",
  38899=>"100000101",
  38900=>"111011001",
  38901=>"110000100",
  38902=>"010111011",
  38903=>"011100110",
  38904=>"010100110",
  38905=>"001111110",
  38906=>"010001000",
  38907=>"001110011",
  38908=>"000111011",
  38909=>"010000100",
  38910=>"111000000",
  38911=>"001000110",
  38912=>"111101111",
  38913=>"100011010",
  38914=>"100110110",
  38915=>"110110111",
  38916=>"011001101",
  38917=>"000100100",
  38918=>"011111101",
  38919=>"001011001",
  38920=>"110100011",
  38921=>"110110100",
  38922=>"101110011",
  38923=>"010011100",
  38924=>"000101001",
  38925=>"000111100",
  38926=>"001011001",
  38927=>"010011111",
  38928=>"010000000",
  38929=>"110111110",
  38930=>"100000011",
  38931=>"001101011",
  38932=>"111111011",
  38933=>"101111100",
  38934=>"111011100",
  38935=>"010001001",
  38936=>"000110111",
  38937=>"101110011",
  38938=>"010101110",
  38939=>"110010011",
  38940=>"001011000",
  38941=>"111011101",
  38942=>"101100100",
  38943=>"111101010",
  38944=>"001010000",
  38945=>"011001010",
  38946=>"110100101",
  38947=>"111001001",
  38948=>"110111010",
  38949=>"010011100",
  38950=>"011110010",
  38951=>"011000010",
  38952=>"000001110",
  38953=>"101111110",
  38954=>"111001001",
  38955=>"111011100",
  38956=>"101110111",
  38957=>"010010000",
  38958=>"001011100",
  38959=>"111101100",
  38960=>"111011001",
  38961=>"111110101",
  38962=>"111001101",
  38963=>"111011010",
  38964=>"100010010",
  38965=>"010010011",
  38966=>"111111011",
  38967=>"111010110",
  38968=>"101101000",
  38969=>"010111000",
  38970=>"101000001",
  38971=>"111000001",
  38972=>"010110000",
  38973=>"111100010",
  38974=>"100110111",
  38975=>"000001110",
  38976=>"111100000",
  38977=>"010110000",
  38978=>"011110111",
  38979=>"111100010",
  38980=>"001111010",
  38981=>"111111111",
  38982=>"110000100",
  38983=>"010111010",
  38984=>"010111101",
  38985=>"111010110",
  38986=>"101010100",
  38987=>"011111100",
  38988=>"100011110",
  38989=>"111100001",
  38990=>"010001011",
  38991=>"110100010",
  38992=>"000001011",
  38993=>"010010000",
  38994=>"000111110",
  38995=>"001000011",
  38996=>"011011101",
  38997=>"011111101",
  38998=>"001011010",
  38999=>"111011110",
  39000=>"001110000",
  39001=>"011100101",
  39002=>"011100111",
  39003=>"011101110",
  39004=>"100100100",
  39005=>"111000010",
  39006=>"011101000",
  39007=>"010011111",
  39008=>"101110000",
  39009=>"000001001",
  39010=>"011101001",
  39011=>"110111000",
  39012=>"000011000",
  39013=>"011011011",
  39014=>"110000011",
  39015=>"110101101",
  39016=>"001100000",
  39017=>"010001000",
  39018=>"010000110",
  39019=>"001011110",
  39020=>"001110011",
  39021=>"111000100",
  39022=>"100011111",
  39023=>"100110010",
  39024=>"010110100",
  39025=>"010010111",
  39026=>"011100110",
  39027=>"001100111",
  39028=>"001001111",
  39029=>"001010110",
  39030=>"100111100",
  39031=>"001000000",
  39032=>"111101000",
  39033=>"110111000",
  39034=>"000101111",
  39035=>"010010000",
  39036=>"110000001",
  39037=>"000010111",
  39038=>"000011110",
  39039=>"101010100",
  39040=>"001001011",
  39041=>"110101100",
  39042=>"100100100",
  39043=>"000100000",
  39044=>"011011001",
  39045=>"001110100",
  39046=>"101101001",
  39047=>"110111001",
  39048=>"101011001",
  39049=>"111110011",
  39050=>"111000110",
  39051=>"100001100",
  39052=>"111101111",
  39053=>"110000101",
  39054=>"000111001",
  39055=>"001011001",
  39056=>"100011110",
  39057=>"111010110",
  39058=>"010110100",
  39059=>"101001100",
  39060=>"010111011",
  39061=>"101110111",
  39062=>"010001010",
  39063=>"101010011",
  39064=>"001110001",
  39065=>"001001111",
  39066=>"111110111",
  39067=>"000001100",
  39068=>"111101100",
  39069=>"001110111",
  39070=>"110100001",
  39071=>"111010111",
  39072=>"111111101",
  39073=>"100010110",
  39074=>"001110110",
  39075=>"110001011",
  39076=>"011101111",
  39077=>"000110010",
  39078=>"100011001",
  39079=>"000101011",
  39080=>"110011100",
  39081=>"000100100",
  39082=>"000000111",
  39083=>"000001000",
  39084=>"001010100",
  39085=>"011101111",
  39086=>"000000110",
  39087=>"100000101",
  39088=>"000011110",
  39089=>"111010101",
  39090=>"001111111",
  39091=>"000101110",
  39092=>"110011100",
  39093=>"011111001",
  39094=>"100100000",
  39095=>"100000001",
  39096=>"000101001",
  39097=>"000110111",
  39098=>"110110111",
  39099=>"111110110",
  39100=>"000001001",
  39101=>"010001010",
  39102=>"001100000",
  39103=>"110110111",
  39104=>"111010011",
  39105=>"001010010",
  39106=>"100000010",
  39107=>"010100001",
  39108=>"101011110",
  39109=>"011110110",
  39110=>"010011111",
  39111=>"110001100",
  39112=>"001101110",
  39113=>"110011101",
  39114=>"111101111",
  39115=>"010101011",
  39116=>"001100101",
  39117=>"101010001",
  39118=>"111100110",
  39119=>"011000010",
  39120=>"011001110",
  39121=>"001000010",
  39122=>"110011100",
  39123=>"000001000",
  39124=>"000110011",
  39125=>"100001001",
  39126=>"001011110",
  39127=>"001110101",
  39128=>"011110010",
  39129=>"100010011",
  39130=>"111010101",
  39131=>"000001100",
  39132=>"100000011",
  39133=>"011010110",
  39134=>"011011010",
  39135=>"001000111",
  39136=>"001100100",
  39137=>"000001111",
  39138=>"110010101",
  39139=>"100010100",
  39140=>"010100100",
  39141=>"001110010",
  39142=>"011111101",
  39143=>"111101011",
  39144=>"000100101",
  39145=>"001110010",
  39146=>"000100100",
  39147=>"101100101",
  39148=>"011110000",
  39149=>"011110110",
  39150=>"111011000",
  39151=>"010100100",
  39152=>"010010000",
  39153=>"111011111",
  39154=>"111011101",
  39155=>"001001110",
  39156=>"001010110",
  39157=>"000011101",
  39158=>"100101100",
  39159=>"101100111",
  39160=>"110011010",
  39161=>"110110000",
  39162=>"101010100",
  39163=>"010110010",
  39164=>"111111000",
  39165=>"011110111",
  39166=>"011111110",
  39167=>"010011001",
  39168=>"110001001",
  39169=>"010010001",
  39170=>"100100000",
  39171=>"001100110",
  39172=>"100010101",
  39173=>"111111011",
  39174=>"010011010",
  39175=>"111001111",
  39176=>"101001111",
  39177=>"101100010",
  39178=>"100111100",
  39179=>"011010111",
  39180=>"010010011",
  39181=>"110001001",
  39182=>"101111110",
  39183=>"101011100",
  39184=>"011101101",
  39185=>"000000100",
  39186=>"101111101",
  39187=>"000010000",
  39188=>"111100100",
  39189=>"000010101",
  39190=>"111110100",
  39191=>"011111100",
  39192=>"000110110",
  39193=>"110100111",
  39194=>"011100100",
  39195=>"111110100",
  39196=>"000011111",
  39197=>"101001000",
  39198=>"111000110",
  39199=>"100001000",
  39200=>"100110100",
  39201=>"010110010",
  39202=>"010100111",
  39203=>"100000010",
  39204=>"101101000",
  39205=>"101011001",
  39206=>"000011011",
  39207=>"101011010",
  39208=>"100111110",
  39209=>"010110001",
  39210=>"010101010",
  39211=>"000110110",
  39212=>"111110111",
  39213=>"101100011",
  39214=>"101000111",
  39215=>"011000111",
  39216=>"010100000",
  39217=>"100110100",
  39218=>"110111000",
  39219=>"110011010",
  39220=>"110100000",
  39221=>"011100100",
  39222=>"100110110",
  39223=>"100110101",
  39224=>"110011110",
  39225=>"100001100",
  39226=>"101111001",
  39227=>"010001111",
  39228=>"001110100",
  39229=>"001101010",
  39230=>"011101110",
  39231=>"100010000",
  39232=>"000111001",
  39233=>"001110111",
  39234=>"000111110",
  39235=>"011100101",
  39236=>"111111010",
  39237=>"001100010",
  39238=>"101011000",
  39239=>"000111001",
  39240=>"111101101",
  39241=>"011000111",
  39242=>"100100000",
  39243=>"011110011",
  39244=>"110111010",
  39245=>"111101100",
  39246=>"000001001",
  39247=>"111000101",
  39248=>"010000010",
  39249=>"011000101",
  39250=>"110101000",
  39251=>"110101000",
  39252=>"010111100",
  39253=>"111110101",
  39254=>"111000100",
  39255=>"111110110",
  39256=>"100100011",
  39257=>"011110011",
  39258=>"100011101",
  39259=>"100110000",
  39260=>"110011001",
  39261=>"110000011",
  39262=>"100000011",
  39263=>"000111110",
  39264=>"101010111",
  39265=>"110111111",
  39266=>"011001000",
  39267=>"110001001",
  39268=>"010010101",
  39269=>"001101101",
  39270=>"111111010",
  39271=>"000110111",
  39272=>"001010000",
  39273=>"101110110",
  39274=>"101001111",
  39275=>"111001100",
  39276=>"111001010",
  39277=>"111100100",
  39278=>"111001101",
  39279=>"000101111",
  39280=>"111010011",
  39281=>"001010001",
  39282=>"110100101",
  39283=>"111011010",
  39284=>"011101101",
  39285=>"111111111",
  39286=>"111101000",
  39287=>"110100000",
  39288=>"011111000",
  39289=>"011110101",
  39290=>"100001010",
  39291=>"000100101",
  39292=>"010111111",
  39293=>"101110111",
  39294=>"100110110",
  39295=>"000111101",
  39296=>"110111100",
  39297=>"100011100",
  39298=>"001000101",
  39299=>"101000110",
  39300=>"011111000",
  39301=>"101111000",
  39302=>"000011101",
  39303=>"010100010",
  39304=>"011011000",
  39305=>"111011111",
  39306=>"000011011",
  39307=>"101101111",
  39308=>"110011111",
  39309=>"101010010",
  39310=>"101011110",
  39311=>"111010000",
  39312=>"001110101",
  39313=>"001011100",
  39314=>"101110010",
  39315=>"001011000",
  39316=>"000000000",
  39317=>"001101010",
  39318=>"010111010",
  39319=>"111101111",
  39320=>"011010010",
  39321=>"101001011",
  39322=>"010000000",
  39323=>"010001001",
  39324=>"111001010",
  39325=>"000100011",
  39326=>"100000000",
  39327=>"011000001",
  39328=>"111101000",
  39329=>"000000000",
  39330=>"110011010",
  39331=>"101010110",
  39332=>"111001010",
  39333=>"100101001",
  39334=>"111010110",
  39335=>"001111010",
  39336=>"001001010",
  39337=>"010011111",
  39338=>"100010000",
  39339=>"101000100",
  39340=>"111101000",
  39341=>"000001000",
  39342=>"001011000",
  39343=>"001101001",
  39344=>"000110010",
  39345=>"011001101",
  39346=>"111101111",
  39347=>"011010011",
  39348=>"110110000",
  39349=>"101001101",
  39350=>"011000100",
  39351=>"011101010",
  39352=>"001110100",
  39353=>"100010110",
  39354=>"111010001",
  39355=>"110011110",
  39356=>"010000100",
  39357=>"101110110",
  39358=>"000110111",
  39359=>"010100000",
  39360=>"111110011",
  39361=>"001011100",
  39362=>"100110110",
  39363=>"010110000",
  39364=>"111000101",
  39365=>"110101111",
  39366=>"110100011",
  39367=>"101111101",
  39368=>"000111000",
  39369=>"110100110",
  39370=>"010110000",
  39371=>"110110000",
  39372=>"001011101",
  39373=>"111011010",
  39374=>"000111100",
  39375=>"111110101",
  39376=>"011011111",
  39377=>"110111110",
  39378=>"110101111",
  39379=>"000010101",
  39380=>"101010110",
  39381=>"110101001",
  39382=>"111101101",
  39383=>"101110001",
  39384=>"101110010",
  39385=>"111110001",
  39386=>"000110100",
  39387=>"100100000",
  39388=>"001000110",
  39389=>"010000100",
  39390=>"011110110",
  39391=>"010010110",
  39392=>"010010100",
  39393=>"010000110",
  39394=>"011000101",
  39395=>"001111010",
  39396=>"010111100",
  39397=>"001000001",
  39398=>"000011001",
  39399=>"000010001",
  39400=>"001011010",
  39401=>"000111010",
  39402=>"011101011",
  39403=>"000101110",
  39404=>"110100101",
  39405=>"010011101",
  39406=>"101101100",
  39407=>"101111010",
  39408=>"000101110",
  39409=>"101111000",
  39410=>"100100100",
  39411=>"111111001",
  39412=>"000010000",
  39413=>"110101000",
  39414=>"000111010",
  39415=>"111011101",
  39416=>"101000011",
  39417=>"011001100",
  39418=>"101001010",
  39419=>"101011011",
  39420=>"100100111",
  39421=>"001001000",
  39422=>"110000110",
  39423=>"100010011",
  39424=>"100111100",
  39425=>"100010000",
  39426=>"110000100",
  39427=>"010011100",
  39428=>"010000001",
  39429=>"011111111",
  39430=>"011100101",
  39431=>"001110001",
  39432=>"100101010",
  39433=>"111001010",
  39434=>"100010101",
  39435=>"000000010",
  39436=>"010111011",
  39437=>"011100111",
  39438=>"000000010",
  39439=>"001101000",
  39440=>"100111101",
  39441=>"101101101",
  39442=>"110101101",
  39443=>"001000101",
  39444=>"010000111",
  39445=>"100001110",
  39446=>"100100010",
  39447=>"101100110",
  39448=>"101000010",
  39449=>"100100011",
  39450=>"100011101",
  39451=>"111000110",
  39452=>"011101111",
  39453=>"110001001",
  39454=>"101101100",
  39455=>"101100010",
  39456=>"001010101",
  39457=>"010111111",
  39458=>"101111110",
  39459=>"001111111",
  39460=>"111110110",
  39461=>"011111111",
  39462=>"000011000",
  39463=>"100101011",
  39464=>"111101111",
  39465=>"010101010",
  39466=>"010111101",
  39467=>"111011111",
  39468=>"000000000",
  39469=>"111010001",
  39470=>"000011110",
  39471=>"011111000",
  39472=>"110100111",
  39473=>"110010111",
  39474=>"011100100",
  39475=>"000101011",
  39476=>"010111111",
  39477=>"001101011",
  39478=>"101110000",
  39479=>"111101101",
  39480=>"100100101",
  39481=>"000101100",
  39482=>"001110011",
  39483=>"110111100",
  39484=>"110111111",
  39485=>"101001000",
  39486=>"100001010",
  39487=>"101100110",
  39488=>"010101010",
  39489=>"010011101",
  39490=>"001101011",
  39491=>"111110011",
  39492=>"110110000",
  39493=>"100110001",
  39494=>"111101001",
  39495=>"101100110",
  39496=>"000001110",
  39497=>"011110011",
  39498=>"000000111",
  39499=>"010010000",
  39500=>"110000101",
  39501=>"000010001",
  39502=>"100001111",
  39503=>"101001001",
  39504=>"101011010",
  39505=>"001111000",
  39506=>"010110100",
  39507=>"011000011",
  39508=>"111011111",
  39509=>"011010011",
  39510=>"001111111",
  39511=>"111000011",
  39512=>"000000101",
  39513=>"000011010",
  39514=>"101010001",
  39515=>"011011110",
  39516=>"010101001",
  39517=>"101100110",
  39518=>"011010110",
  39519=>"100110010",
  39520=>"010011110",
  39521=>"100000000",
  39522=>"110000101",
  39523=>"111110011",
  39524=>"011011011",
  39525=>"110100111",
  39526=>"001010101",
  39527=>"100100001",
  39528=>"011001000",
  39529=>"001111110",
  39530=>"111110000",
  39531=>"110010101",
  39532=>"101011110",
  39533=>"111001111",
  39534=>"110001101",
  39535=>"101010010",
  39536=>"011101001",
  39537=>"111111011",
  39538=>"001001011",
  39539=>"010111100",
  39540=>"000100111",
  39541=>"010100100",
  39542=>"111010110",
  39543=>"100101101",
  39544=>"000100000",
  39545=>"110111111",
  39546=>"100111010",
  39547=>"111111101",
  39548=>"111001000",
  39549=>"011011110",
  39550=>"011110001",
  39551=>"110111110",
  39552=>"100110010",
  39553=>"011011010",
  39554=>"111010010",
  39555=>"001001011",
  39556=>"100101111",
  39557=>"110000110",
  39558=>"011000101",
  39559=>"111011011",
  39560=>"001111010",
  39561=>"011011001",
  39562=>"110111011",
  39563=>"010001111",
  39564=>"001000010",
  39565=>"000000011",
  39566=>"111010111",
  39567=>"111111001",
  39568=>"111011011",
  39569=>"100000111",
  39570=>"011100000",
  39571=>"000011111",
  39572=>"100010101",
  39573=>"001101110",
  39574=>"100100010",
  39575=>"110101111",
  39576=>"011011111",
  39577=>"001001000",
  39578=>"100101010",
  39579=>"111010010",
  39580=>"101110100",
  39581=>"101000001",
  39582=>"000001111",
  39583=>"010111011",
  39584=>"100001011",
  39585=>"010001100",
  39586=>"101111000",
  39587=>"010111110",
  39588=>"101000010",
  39589=>"011011111",
  39590=>"101011100",
  39591=>"100110001",
  39592=>"110100111",
  39593=>"000111000",
  39594=>"011000110",
  39595=>"001110010",
  39596=>"011001100",
  39597=>"111111101",
  39598=>"000000110",
  39599=>"100001100",
  39600=>"101011000",
  39601=>"000101000",
  39602=>"000000111",
  39603=>"111000111",
  39604=>"000010111",
  39605=>"110100100",
  39606=>"001010010",
  39607=>"111010100",
  39608=>"001101011",
  39609=>"010111111",
  39610=>"110000010",
  39611=>"000111111",
  39612=>"010000110",
  39613=>"010110001",
  39614=>"001001100",
  39615=>"100011111",
  39616=>"111100010",
  39617=>"100000100",
  39618=>"111111000",
  39619=>"000101101",
  39620=>"011001010",
  39621=>"000100000",
  39622=>"110110111",
  39623=>"101000100",
  39624=>"111001111",
  39625=>"110011101",
  39626=>"000110010",
  39627=>"011110010",
  39628=>"100110101",
  39629=>"110101111",
  39630=>"111100010",
  39631=>"011100000",
  39632=>"001010000",
  39633=>"011001110",
  39634=>"011011000",
  39635=>"010010111",
  39636=>"101011011",
  39637=>"101101110",
  39638=>"011011011",
  39639=>"101101100",
  39640=>"010011110",
  39641=>"101100001",
  39642=>"001010110",
  39643=>"001010111",
  39644=>"111101001",
  39645=>"100110010",
  39646=>"001110001",
  39647=>"001011010",
  39648=>"111000101",
  39649=>"111110101",
  39650=>"101110111",
  39651=>"010110111",
  39652=>"110110001",
  39653=>"011100111",
  39654=>"101100011",
  39655=>"001100110",
  39656=>"101110111",
  39657=>"000101001",
  39658=>"011110111",
  39659=>"101101010",
  39660=>"111011110",
  39661=>"010001111",
  39662=>"100010110",
  39663=>"000010000",
  39664=>"011111101",
  39665=>"000101101",
  39666=>"000010101",
  39667=>"001000011",
  39668=>"101101001",
  39669=>"101001100",
  39670=>"111000001",
  39671=>"111101010",
  39672=>"000001011",
  39673=>"000100011",
  39674=>"101000100",
  39675=>"110011111",
  39676=>"000000010",
  39677=>"100010000",
  39678=>"001000000",
  39679=>"010100101",
  39680=>"011100010",
  39681=>"110111000",
  39682=>"110110000",
  39683=>"000000011",
  39684=>"000010111",
  39685=>"110111011",
  39686=>"010100111",
  39687=>"011100000",
  39688=>"001001000",
  39689=>"001001001",
  39690=>"111011101",
  39691=>"110101101",
  39692=>"010001001",
  39693=>"111101110",
  39694=>"011001101",
  39695=>"000000010",
  39696=>"001110011",
  39697=>"100011110",
  39698=>"001010001",
  39699=>"110001011",
  39700=>"100001000",
  39701=>"100110010",
  39702=>"000100110",
  39703=>"011101001",
  39704=>"100010001",
  39705=>"111000010",
  39706=>"001000001",
  39707=>"001011001",
  39708=>"001000100",
  39709=>"110001111",
  39710=>"011000100",
  39711=>"000000111",
  39712=>"001101111",
  39713=>"000010011",
  39714=>"011001010",
  39715=>"111110000",
  39716=>"001010001",
  39717=>"001010011",
  39718=>"100001100",
  39719=>"011100101",
  39720=>"111110001",
  39721=>"101000000",
  39722=>"100000000",
  39723=>"110111101",
  39724=>"110100101",
  39725=>"111011100",
  39726=>"100101010",
  39727=>"101000111",
  39728=>"000101001",
  39729=>"001010110",
  39730=>"110110101",
  39731=>"011111010",
  39732=>"001101011",
  39733=>"000110111",
  39734=>"011111011",
  39735=>"000000011",
  39736=>"011100110",
  39737=>"010011001",
  39738=>"100000110",
  39739=>"100111000",
  39740=>"110101111",
  39741=>"010110001",
  39742=>"001110001",
  39743=>"000000010",
  39744=>"110110111",
  39745=>"010001101",
  39746=>"010101111",
  39747=>"101111111",
  39748=>"000110001",
  39749=>"000101110",
  39750=>"110000100",
  39751=>"011010010",
  39752=>"100010000",
  39753=>"000110110",
  39754=>"010000100",
  39755=>"100011100",
  39756=>"000101010",
  39757=>"010111001",
  39758=>"111000010",
  39759=>"110011000",
  39760=>"100001001",
  39761=>"111101000",
  39762=>"111110111",
  39763=>"100101001",
  39764=>"111001101",
  39765=>"010001100",
  39766=>"000010010",
  39767=>"011001010",
  39768=>"111101000",
  39769=>"100101010",
  39770=>"100111111",
  39771=>"100101000",
  39772=>"000011000",
  39773=>"111000101",
  39774=>"000110000",
  39775=>"110001100",
  39776=>"010000010",
  39777=>"000110100",
  39778=>"011011111",
  39779=>"011010101",
  39780=>"001101000",
  39781=>"101101110",
  39782=>"101010010",
  39783=>"111111100",
  39784=>"000001001",
  39785=>"111001011",
  39786=>"010111001",
  39787=>"100101001",
  39788=>"101101010",
  39789=>"011001110",
  39790=>"110000101",
  39791=>"010001001",
  39792=>"100000010",
  39793=>"011111000",
  39794=>"010000011",
  39795=>"011110111",
  39796=>"110110011",
  39797=>"011011111",
  39798=>"001101000",
  39799=>"001101000",
  39800=>"111111100",
  39801=>"000000010",
  39802=>"000111111",
  39803=>"001100110",
  39804=>"000010111",
  39805=>"111000101",
  39806=>"111111000",
  39807=>"111011000",
  39808=>"111111010",
  39809=>"010011101",
  39810=>"101101101",
  39811=>"110111101",
  39812=>"010110101",
  39813=>"010000001",
  39814=>"000001001",
  39815=>"000111111",
  39816=>"011111110",
  39817=>"101011000",
  39818=>"001011000",
  39819=>"100101000",
  39820=>"111100010",
  39821=>"000010110",
  39822=>"110110110",
  39823=>"011010001",
  39824=>"111111100",
  39825=>"011001001",
  39826=>"111110001",
  39827=>"100011111",
  39828=>"001011000",
  39829=>"010101001",
  39830=>"000110001",
  39831=>"001100111",
  39832=>"001000010",
  39833=>"100001101",
  39834=>"100100101",
  39835=>"111011011",
  39836=>"110110011",
  39837=>"001001101",
  39838=>"110001000",
  39839=>"010000110",
  39840=>"111101100",
  39841=>"110100011",
  39842=>"010111101",
  39843=>"000001101",
  39844=>"101111011",
  39845=>"001101110",
  39846=>"110010111",
  39847=>"010100101",
  39848=>"001011110",
  39849=>"101111000",
  39850=>"010001000",
  39851=>"010001010",
  39852=>"101100110",
  39853=>"110100001",
  39854=>"101010011",
  39855=>"110011011",
  39856=>"000010110",
  39857=>"011111010",
  39858=>"100000001",
  39859=>"000000011",
  39860=>"011110010",
  39861=>"110000000",
  39862=>"101010010",
  39863=>"000011100",
  39864=>"000111100",
  39865=>"100001111",
  39866=>"011111111",
  39867=>"011101111",
  39868=>"101110000",
  39869=>"111101010",
  39870=>"000111011",
  39871=>"011101101",
  39872=>"001101011",
  39873=>"111100010",
  39874=>"110111110",
  39875=>"010010101",
  39876=>"000010010",
  39877=>"111010010",
  39878=>"010111110",
  39879=>"010110000",
  39880=>"010000100",
  39881=>"011110100",
  39882=>"101111110",
  39883=>"010111000",
  39884=>"000010000",
  39885=>"001111111",
  39886=>"010110011",
  39887=>"010011100",
  39888=>"101010101",
  39889=>"100010101",
  39890=>"101110110",
  39891=>"010001011",
  39892=>"000001100",
  39893=>"111110000",
  39894=>"111100111",
  39895=>"011010110",
  39896=>"001010100",
  39897=>"100000000",
  39898=>"001000010",
  39899=>"001000011",
  39900=>"100101011",
  39901=>"011100010",
  39902=>"101111001",
  39903=>"100001010",
  39904=>"000101011",
  39905=>"100010101",
  39906=>"110001111",
  39907=>"000101100",
  39908=>"110110010",
  39909=>"001001000",
  39910=>"101000000",
  39911=>"101000011",
  39912=>"101100000",
  39913=>"011011000",
  39914=>"111101000",
  39915=>"001001000",
  39916=>"011011101",
  39917=>"101100011",
  39918=>"010100110",
  39919=>"110101111",
  39920=>"000111111",
  39921=>"001011111",
  39922=>"101111011",
  39923=>"001110000",
  39924=>"000001111",
  39925=>"000010110",
  39926=>"011101110",
  39927=>"111001001",
  39928=>"110001100",
  39929=>"110000100",
  39930=>"111001111",
  39931=>"111111001",
  39932=>"111011010",
  39933=>"010001110",
  39934=>"010000111",
  39935=>"010000110",
  39936=>"110111000",
  39937=>"111001000",
  39938=>"101111111",
  39939=>"010110101",
  39940=>"111111111",
  39941=>"110100111",
  39942=>"010000011",
  39943=>"010000000",
  39944=>"110111101",
  39945=>"001101101",
  39946=>"000010010",
  39947=>"101110111",
  39948=>"000000000",
  39949=>"010000111",
  39950=>"011101011",
  39951=>"100111110",
  39952=>"001111000",
  39953=>"000001110",
  39954=>"111110100",
  39955=>"011111011",
  39956=>"001001111",
  39957=>"101100111",
  39958=>"111111111",
  39959=>"100000001",
  39960=>"110101000",
  39961=>"111110110",
  39962=>"010100110",
  39963=>"110010110",
  39964=>"000100110",
  39965=>"101000011",
  39966=>"101001111",
  39967=>"010001111",
  39968=>"001000110",
  39969=>"010011110",
  39970=>"011111001",
  39971=>"000100100",
  39972=>"101001000",
  39973=>"100111111",
  39974=>"011111110",
  39975=>"010100101",
  39976=>"001100111",
  39977=>"011010100",
  39978=>"100101011",
  39979=>"000101111",
  39980=>"010011111",
  39981=>"111011010",
  39982=>"101111110",
  39983=>"001100100",
  39984=>"110010101",
  39985=>"110111100",
  39986=>"111100010",
  39987=>"111111001",
  39988=>"011110111",
  39989=>"011101001",
  39990=>"010101001",
  39991=>"000111001",
  39992=>"100010000",
  39993=>"011000110",
  39994=>"101010111",
  39995=>"100010100",
  39996=>"000001110",
  39997=>"101110000",
  39998=>"001010001",
  39999=>"010001000",
  40000=>"001110100",
  40001=>"001001111",
  40002=>"001001100",
  40003=>"001010001",
  40004=>"010000111",
  40005=>"110000010",
  40006=>"111011101",
  40007=>"001001001",
  40008=>"100010100",
  40009=>"011110011",
  40010=>"010110110",
  40011=>"000010000",
  40012=>"101000110",
  40013=>"101101100",
  40014=>"010100000",
  40015=>"110101001",
  40016=>"000011111",
  40017=>"001100101",
  40018=>"011111111",
  40019=>"001011111",
  40020=>"000110111",
  40021=>"000101001",
  40022=>"001010011",
  40023=>"000110000",
  40024=>"001000101",
  40025=>"011011111",
  40026=>"100111001",
  40027=>"001001000",
  40028=>"010101000",
  40029=>"000101110",
  40030=>"101111001",
  40031=>"100000001",
  40032=>"000110001",
  40033=>"000000100",
  40034=>"000001101",
  40035=>"011100100",
  40036=>"001000111",
  40037=>"011001101",
  40038=>"001011001",
  40039=>"101100111",
  40040=>"111100011",
  40041=>"110111111",
  40042=>"000110111",
  40043=>"111100110",
  40044=>"101000001",
  40045=>"101101001",
  40046=>"010011000",
  40047=>"110011111",
  40048=>"010010111",
  40049=>"111001100",
  40050=>"111011010",
  40051=>"111011001",
  40052=>"010010100",
  40053=>"111001000",
  40054=>"100000110",
  40055=>"110000110",
  40056=>"101101100",
  40057=>"000101101",
  40058=>"010110111",
  40059=>"101010110",
  40060=>"011111101",
  40061=>"101111110",
  40062=>"100000001",
  40063=>"111000100",
  40064=>"011001010",
  40065=>"001000010",
  40066=>"000010011",
  40067=>"011101001",
  40068=>"011110001",
  40069=>"110000110",
  40070=>"011000110",
  40071=>"100010011",
  40072=>"110101000",
  40073=>"001101111",
  40074=>"001110100",
  40075=>"101001101",
  40076=>"100110000",
  40077=>"001000111",
  40078=>"010000101",
  40079=>"100110100",
  40080=>"010100100",
  40081=>"100101010",
  40082=>"110000000",
  40083=>"010010110",
  40084=>"100000001",
  40085=>"001000010",
  40086=>"100100010",
  40087=>"111100010",
  40088=>"001001010",
  40089=>"000101001",
  40090=>"001010011",
  40091=>"011111100",
  40092=>"101010110",
  40093=>"010011011",
  40094=>"110110010",
  40095=>"110011110",
  40096=>"001001100",
  40097=>"111000110",
  40098=>"111001001",
  40099=>"000000011",
  40100=>"110101001",
  40101=>"000100001",
  40102=>"100101010",
  40103=>"010111001",
  40104=>"110010000",
  40105=>"101101011",
  40106=>"110000001",
  40107=>"101110111",
  40108=>"101010010",
  40109=>"111101001",
  40110=>"010000011",
  40111=>"001000000",
  40112=>"001101110",
  40113=>"001010011",
  40114=>"000011011",
  40115=>"000000011",
  40116=>"100110111",
  40117=>"111010101",
  40118=>"001001010",
  40119=>"010100001",
  40120=>"101100100",
  40121=>"010000000",
  40122=>"101010011",
  40123=>"001010100",
  40124=>"011101111",
  40125=>"110110010",
  40126=>"110000000",
  40127=>"111110101",
  40128=>"000010000",
  40129=>"111001111",
  40130=>"110100011",
  40131=>"000011010",
  40132=>"110011100",
  40133=>"010010100",
  40134=>"010101010",
  40135=>"101001001",
  40136=>"111101000",
  40137=>"001001100",
  40138=>"101101111",
  40139=>"000111111",
  40140=>"010101000",
  40141=>"100010001",
  40142=>"000011111",
  40143=>"001011001",
  40144=>"001000111",
  40145=>"110111001",
  40146=>"100100000",
  40147=>"010111100",
  40148=>"101001110",
  40149=>"110010111",
  40150=>"010011111",
  40151=>"100110100",
  40152=>"111011000",
  40153=>"111011001",
  40154=>"000000000",
  40155=>"100110101",
  40156=>"000101001",
  40157=>"010100101",
  40158=>"010000100",
  40159=>"110101010",
  40160=>"101001100",
  40161=>"110100111",
  40162=>"000110000",
  40163=>"000000011",
  40164=>"011011110",
  40165=>"001110011",
  40166=>"000000101",
  40167=>"011111100",
  40168=>"011000000",
  40169=>"101001111",
  40170=>"000000000",
  40171=>"110000100",
  40172=>"010000111",
  40173=>"100000111",
  40174=>"101101001",
  40175=>"001010011",
  40176=>"111001110",
  40177=>"011100101",
  40178=>"110010010",
  40179=>"101001100",
  40180=>"101100101",
  40181=>"100011100",
  40182=>"010001001",
  40183=>"010011111",
  40184=>"100100110",
  40185=>"110101010",
  40186=>"001101101",
  40187=>"010010000",
  40188=>"100110110",
  40189=>"111110010",
  40190=>"010010110",
  40191=>"101010000",
  40192=>"111101101",
  40193=>"111010001",
  40194=>"111010111",
  40195=>"000001000",
  40196=>"010011011",
  40197=>"001011010",
  40198=>"010000010",
  40199=>"100010100",
  40200=>"000000010",
  40201=>"100010010",
  40202=>"110011100",
  40203=>"011001010",
  40204=>"100110001",
  40205=>"001110010",
  40206=>"011111011",
  40207=>"001111111",
  40208=>"001100001",
  40209=>"111110000",
  40210=>"101000010",
  40211=>"010110111",
  40212=>"100100100",
  40213=>"000011001",
  40214=>"011010100",
  40215=>"000111011",
  40216=>"001000001",
  40217=>"100111000",
  40218=>"001100100",
  40219=>"011001010",
  40220=>"010011001",
  40221=>"011000101",
  40222=>"100110010",
  40223=>"000000110",
  40224=>"101001011",
  40225=>"000110000",
  40226=>"010010100",
  40227=>"110000100",
  40228=>"000001011",
  40229=>"000101111",
  40230=>"111010111",
  40231=>"001111110",
  40232=>"110010101",
  40233=>"111010011",
  40234=>"001000101",
  40235=>"101011000",
  40236=>"110100011",
  40237=>"011001000",
  40238=>"000010110",
  40239=>"000100110",
  40240=>"011111101",
  40241=>"000110100",
  40242=>"010001110",
  40243=>"001110111",
  40244=>"101110100",
  40245=>"000100110",
  40246=>"000011011",
  40247=>"110000011",
  40248=>"000000111",
  40249=>"100000000",
  40250=>"111111101",
  40251=>"100110100",
  40252=>"001111001",
  40253=>"111111100",
  40254=>"110111110",
  40255=>"001001001",
  40256=>"001010111",
  40257=>"000001101",
  40258=>"111110100",
  40259=>"001101101",
  40260=>"000100011",
  40261=>"110101000",
  40262=>"011000101",
  40263=>"110011110",
  40264=>"010111100",
  40265=>"000000000",
  40266=>"100010000",
  40267=>"001010010",
  40268=>"111100111",
  40269=>"101001111",
  40270=>"110111111",
  40271=>"010110010",
  40272=>"011100100",
  40273=>"100010011",
  40274=>"000000011",
  40275=>"000100101",
  40276=>"010110100",
  40277=>"111000100",
  40278=>"110110101",
  40279=>"000100011",
  40280=>"101010000",
  40281=>"001101010",
  40282=>"100110101",
  40283=>"110000010",
  40284=>"111001101",
  40285=>"111100011",
  40286=>"111001011",
  40287=>"110000011",
  40288=>"001010000",
  40289=>"110001001",
  40290=>"000100011",
  40291=>"010111011",
  40292=>"110001000",
  40293=>"101110011",
  40294=>"010001001",
  40295=>"011100010",
  40296=>"111011001",
  40297=>"001111011",
  40298=>"000101000",
  40299=>"001100000",
  40300=>"111101101",
  40301=>"100101100",
  40302=>"010100001",
  40303=>"111101101",
  40304=>"100011100",
  40305=>"100110000",
  40306=>"111011011",
  40307=>"110100010",
  40308=>"101011110",
  40309=>"111100010",
  40310=>"111010010",
  40311=>"111110110",
  40312=>"001101011",
  40313=>"101110000",
  40314=>"011111111",
  40315=>"100111100",
  40316=>"010100001",
  40317=>"100010111",
  40318=>"100000111",
  40319=>"000001000",
  40320=>"110011111",
  40321=>"110011111",
  40322=>"101110101",
  40323=>"001101011",
  40324=>"000110001",
  40325=>"110000000",
  40326=>"000111111",
  40327=>"111011111",
  40328=>"011000000",
  40329=>"001011110",
  40330=>"111101111",
  40331=>"101010010",
  40332=>"100000110",
  40333=>"000010001",
  40334=>"000001100",
  40335=>"110011110",
  40336=>"000111011",
  40337=>"001110000",
  40338=>"111001110",
  40339=>"000001101",
  40340=>"000110010",
  40341=>"110010100",
  40342=>"111110100",
  40343=>"111011011",
  40344=>"001111111",
  40345=>"101000011",
  40346=>"000111011",
  40347=>"101011001",
  40348=>"100110100",
  40349=>"101111100",
  40350=>"100001010",
  40351=>"011101001",
  40352=>"111111111",
  40353=>"001111100",
  40354=>"001101001",
  40355=>"101001010",
  40356=>"101000000",
  40357=>"100010101",
  40358=>"011010001",
  40359=>"100001010",
  40360=>"010010111",
  40361=>"000011011",
  40362=>"111011001",
  40363=>"101110011",
  40364=>"110011010",
  40365=>"011101001",
  40366=>"010011110",
  40367=>"110101101",
  40368=>"000100100",
  40369=>"110011110",
  40370=>"100000101",
  40371=>"001010001",
  40372=>"010001000",
  40373=>"100100000",
  40374=>"111101000",
  40375=>"000000011",
  40376=>"000110001",
  40377=>"010110010",
  40378=>"010001110",
  40379=>"010100111",
  40380=>"011110100",
  40381=>"011111001",
  40382=>"000000000",
  40383=>"110110111",
  40384=>"010010000",
  40385=>"010011111",
  40386=>"000011001",
  40387=>"001000110",
  40388=>"110001110",
  40389=>"010001001",
  40390=>"001011110",
  40391=>"001001100",
  40392=>"111001101",
  40393=>"001110110",
  40394=>"010111001",
  40395=>"010010010",
  40396=>"110011000",
  40397=>"110111100",
  40398=>"011000001",
  40399=>"001010101",
  40400=>"000100010",
  40401=>"000000001",
  40402=>"000010000",
  40403=>"011000000",
  40404=>"100010000",
  40405=>"000010100",
  40406=>"100110011",
  40407=>"011010101",
  40408=>"100001100",
  40409=>"111111011",
  40410=>"011100010",
  40411=>"100000101",
  40412=>"010011110",
  40413=>"010000110",
  40414=>"000011001",
  40415=>"111101111",
  40416=>"110000111",
  40417=>"010110000",
  40418=>"110000010",
  40419=>"010001001",
  40420=>"000101011",
  40421=>"101110001",
  40422=>"100010010",
  40423=>"001101001",
  40424=>"001111011",
  40425=>"111000101",
  40426=>"110011111",
  40427=>"000000010",
  40428=>"001111000",
  40429=>"111010001",
  40430=>"101100111",
  40431=>"010010000",
  40432=>"110000000",
  40433=>"110010101",
  40434=>"111000101",
  40435=>"110010010",
  40436=>"001000011",
  40437=>"111001111",
  40438=>"010111011",
  40439=>"000011010",
  40440=>"000011000",
  40441=>"101011111",
  40442=>"111111100",
  40443=>"001010010",
  40444=>"011001010",
  40445=>"101000110",
  40446=>"101100111",
  40447=>"111100011",
  40448=>"111000110",
  40449=>"110100111",
  40450=>"100100101",
  40451=>"000001110",
  40452=>"001111111",
  40453=>"001100111",
  40454=>"111110111",
  40455=>"010111100",
  40456=>"010010010",
  40457=>"000011100",
  40458=>"001110110",
  40459=>"000110110",
  40460=>"001101001",
  40461=>"000000001",
  40462=>"100100000",
  40463=>"010000000",
  40464=>"011110011",
  40465=>"001100010",
  40466=>"011001011",
  40467=>"110111110",
  40468=>"110000000",
  40469=>"000100000",
  40470=>"110100100",
  40471=>"011001110",
  40472=>"110011100",
  40473=>"010111111",
  40474=>"000011001",
  40475=>"100000110",
  40476=>"011011100",
  40477=>"001100101",
  40478=>"111010011",
  40479=>"101110101",
  40480=>"000100111",
  40481=>"111100101",
  40482=>"010000100",
  40483=>"111001110",
  40484=>"110111101",
  40485=>"100000100",
  40486=>"011111001",
  40487=>"001110111",
  40488=>"000000011",
  40489=>"011101111",
  40490=>"101100010",
  40491=>"111100000",
  40492=>"110010010",
  40493=>"010101111",
  40494=>"001001111",
  40495=>"101010100",
  40496=>"000001100",
  40497=>"011010100",
  40498=>"001100101",
  40499=>"000000011",
  40500=>"010010000",
  40501=>"011001011",
  40502=>"000011010",
  40503=>"100110100",
  40504=>"000000100",
  40505=>"110101100",
  40506=>"000101010",
  40507=>"010100111",
  40508=>"100110100",
  40509=>"010100000",
  40510=>"100110000",
  40511=>"111110110",
  40512=>"110100000",
  40513=>"001110110",
  40514=>"001011010",
  40515=>"001010111",
  40516=>"101010001",
  40517=>"001001011",
  40518=>"010100110",
  40519=>"010010110",
  40520=>"010000111",
  40521=>"111101101",
  40522=>"011000101",
  40523=>"000000100",
  40524=>"000111000",
  40525=>"100100010",
  40526=>"111011110",
  40527=>"101001101",
  40528=>"101000110",
  40529=>"101010111",
  40530=>"100100011",
  40531=>"101000000",
  40532=>"010000001",
  40533=>"100010000",
  40534=>"010110100",
  40535=>"000001100",
  40536=>"100110100",
  40537=>"011111010",
  40538=>"001101010",
  40539=>"010001001",
  40540=>"001001100",
  40541=>"100011111",
  40542=>"001000101",
  40543=>"100100101",
  40544=>"000011010",
  40545=>"100110010",
  40546=>"101101101",
  40547=>"110110100",
  40548=>"010110101",
  40549=>"011010000",
  40550=>"011011010",
  40551=>"100010001",
  40552=>"000000110",
  40553=>"010010110",
  40554=>"000011100",
  40555=>"001110000",
  40556=>"000001111",
  40557=>"011000110",
  40558=>"100110100",
  40559=>"111000010",
  40560=>"010010000",
  40561=>"011000000",
  40562=>"101011100",
  40563=>"101111111",
  40564=>"111101100",
  40565=>"111011011",
  40566=>"111110101",
  40567=>"101011011",
  40568=>"001101000",
  40569=>"100100010",
  40570=>"111101011",
  40571=>"100001000",
  40572=>"000011101",
  40573=>"011000101",
  40574=>"101001110",
  40575=>"010111101",
  40576=>"000111100",
  40577=>"000011111",
  40578=>"110100110",
  40579=>"101000011",
  40580=>"101001000",
  40581=>"101111010",
  40582=>"111100111",
  40583=>"111011011",
  40584=>"100010110",
  40585=>"100111111",
  40586=>"100111001",
  40587=>"000100100",
  40588=>"000110100",
  40589=>"111110100",
  40590=>"111011110",
  40591=>"010100010",
  40592=>"011101110",
  40593=>"100010101",
  40594=>"101100001",
  40595=>"001110011",
  40596=>"100100001",
  40597=>"001000000",
  40598=>"111011101",
  40599=>"000100001",
  40600=>"111111100",
  40601=>"100000100",
  40602=>"000001000",
  40603=>"000001011",
  40604=>"010100000",
  40605=>"101100110",
  40606=>"101101000",
  40607=>"110101100",
  40608=>"101011000",
  40609=>"001110011",
  40610=>"110110010",
  40611=>"111101001",
  40612=>"001010000",
  40613=>"001100000",
  40614=>"001110010",
  40615=>"000101110",
  40616=>"111101001",
  40617=>"001001001",
  40618=>"101000001",
  40619=>"101101001",
  40620=>"010010101",
  40621=>"100101101",
  40622=>"010001101",
  40623=>"011001000",
  40624=>"000000110",
  40625=>"110010011",
  40626=>"001101111",
  40627=>"000100000",
  40628=>"000010101",
  40629=>"010100010",
  40630=>"010010010",
  40631=>"100011100",
  40632=>"111101111",
  40633=>"101000010",
  40634=>"111110110",
  40635=>"000100010",
  40636=>"011110011",
  40637=>"100010011",
  40638=>"101101001",
  40639=>"011110111",
  40640=>"100010000",
  40641=>"101110111",
  40642=>"001011100",
  40643=>"110110011",
  40644=>"100000110",
  40645=>"011100101",
  40646=>"010110111",
  40647=>"110111111",
  40648=>"111000100",
  40649=>"011000000",
  40650=>"011011000",
  40651=>"001110011",
  40652=>"011111010",
  40653=>"100010001",
  40654=>"110110010",
  40655=>"011001011",
  40656=>"011010101",
  40657=>"100101110",
  40658=>"001011011",
  40659=>"110010000",
  40660=>"010000011",
  40661=>"110011100",
  40662=>"100001011",
  40663=>"111110111",
  40664=>"001010110",
  40665=>"010101101",
  40666=>"110101011",
  40667=>"110100000",
  40668=>"100101010",
  40669=>"010100110",
  40670=>"110101001",
  40671=>"100100010",
  40672=>"110001101",
  40673=>"100110101",
  40674=>"111000100",
  40675=>"100100100",
  40676=>"011001100",
  40677=>"011111111",
  40678=>"100010010",
  40679=>"011101000",
  40680=>"100100101",
  40681=>"101100101",
  40682=>"011100010",
  40683=>"000011110",
  40684=>"100000100",
  40685=>"101100110",
  40686=>"100010110",
  40687=>"100110101",
  40688=>"000100000",
  40689=>"100000001",
  40690=>"101111101",
  40691=>"101011100",
  40692=>"110001000",
  40693=>"011001101",
  40694=>"001110101",
  40695=>"111100111",
  40696=>"010011000",
  40697=>"010100101",
  40698=>"001010101",
  40699=>"010001011",
  40700=>"110010011",
  40701=>"101110011",
  40702=>"111111000",
  40703=>"101101001",
  40704=>"000110100",
  40705=>"111101011",
  40706=>"011011011",
  40707=>"010101000",
  40708=>"111110001",
  40709=>"110000010",
  40710=>"101111101",
  40711=>"001111111",
  40712=>"011110001",
  40713=>"100101011",
  40714=>"010011011",
  40715=>"010011011",
  40716=>"101010100",
  40717=>"111010000",
  40718=>"110011101",
  40719=>"100011010",
  40720=>"010001001",
  40721=>"100100110",
  40722=>"110011100",
  40723=>"001100110",
  40724=>"111111100",
  40725=>"110100000",
  40726=>"100110001",
  40727=>"100000111",
  40728=>"010110000",
  40729=>"001100010",
  40730=>"000001111",
  40731=>"111100000",
  40732=>"001110100",
  40733=>"100011100",
  40734=>"000001110",
  40735=>"110001010",
  40736=>"001000100",
  40737=>"110001001",
  40738=>"000110011",
  40739=>"100011001",
  40740=>"000011110",
  40741=>"100010111",
  40742=>"001100011",
  40743=>"100110111",
  40744=>"111110011",
  40745=>"010101010",
  40746=>"101110100",
  40747=>"001110101",
  40748=>"101101101",
  40749=>"000101101",
  40750=>"101000001",
  40751=>"010011010",
  40752=>"110001000",
  40753=>"010111101",
  40754=>"001011001",
  40755=>"010111100",
  40756=>"110110100",
  40757=>"111110100",
  40758=>"011000110",
  40759=>"000101000",
  40760=>"100001111",
  40761=>"101100101",
  40762=>"101010011",
  40763=>"101010011",
  40764=>"011101000",
  40765=>"100100100",
  40766=>"100000000",
  40767=>"110011110",
  40768=>"101110010",
  40769=>"101011011",
  40770=>"100110100",
  40771=>"001101111",
  40772=>"100000100",
  40773=>"111001001",
  40774=>"010000100",
  40775=>"010011111",
  40776=>"110001010",
  40777=>"011111001",
  40778=>"001011110",
  40779=>"000001111",
  40780=>"010010011",
  40781=>"110010010",
  40782=>"100110111",
  40783=>"000011001",
  40784=>"111110100",
  40785=>"000011000",
  40786=>"101010010",
  40787=>"000111001",
  40788=>"001001111",
  40789=>"000100100",
  40790=>"101100000",
  40791=>"001100110",
  40792=>"100011001",
  40793=>"100100100",
  40794=>"110011110",
  40795=>"101010101",
  40796=>"000110111",
  40797=>"100010001",
  40798=>"010011011",
  40799=>"001100000",
  40800=>"111001111",
  40801=>"111110010",
  40802=>"000101100",
  40803=>"100100101",
  40804=>"001001110",
  40805=>"100100100",
  40806=>"110101000",
  40807=>"011101011",
  40808=>"011011110",
  40809=>"010001000",
  40810=>"101101001",
  40811=>"010011101",
  40812=>"111000001",
  40813=>"001001000",
  40814=>"010011111",
  40815=>"011011111",
  40816=>"000101110",
  40817=>"001000100",
  40818=>"110000101",
  40819=>"101000010",
  40820=>"000011000",
  40821=>"001111001",
  40822=>"010000010",
  40823=>"000101110",
  40824=>"111100001",
  40825=>"001111110",
  40826=>"001100111",
  40827=>"110000101",
  40828=>"000000000",
  40829=>"000100100",
  40830=>"110111111",
  40831=>"010001100",
  40832=>"011011001",
  40833=>"101011000",
  40834=>"001000011",
  40835=>"101101010",
  40836=>"000110000",
  40837=>"111110011",
  40838=>"011111100",
  40839=>"110110000",
  40840=>"111001111",
  40841=>"000110001",
  40842=>"000101101",
  40843=>"101000100",
  40844=>"000100010",
  40845=>"000111000",
  40846=>"100011011",
  40847=>"001110100",
  40848=>"110111110",
  40849=>"111111011",
  40850=>"110001010",
  40851=>"110100010",
  40852=>"110000111",
  40853=>"110010110",
  40854=>"100000101",
  40855=>"101100001",
  40856=>"010100010",
  40857=>"101000100",
  40858=>"010111001",
  40859=>"111001010",
  40860=>"100010110",
  40861=>"011011100",
  40862=>"011000000",
  40863=>"110000010",
  40864=>"110011000",
  40865=>"111000101",
  40866=>"100000011",
  40867=>"100001001",
  40868=>"001000000",
  40869=>"101101001",
  40870=>"011011011",
  40871=>"010111000",
  40872=>"111010111",
  40873=>"011101000",
  40874=>"001010010",
  40875=>"000011001",
  40876=>"010000000",
  40877=>"100100110",
  40878=>"010110100",
  40879=>"001010111",
  40880=>"111100000",
  40881=>"110100111",
  40882=>"000011110",
  40883=>"100100001",
  40884=>"000110000",
  40885=>"011011001",
  40886=>"110011110",
  40887=>"110000010",
  40888=>"111010110",
  40889=>"101010101",
  40890=>"110110000",
  40891=>"110111011",
  40892=>"111100011",
  40893=>"010000100",
  40894=>"111100110",
  40895=>"111100111",
  40896=>"011000100",
  40897=>"111000100",
  40898=>"001001001",
  40899=>"000010000",
  40900=>"011100111",
  40901=>"001010001",
  40902=>"001110010",
  40903=>"000010100",
  40904=>"100000000",
  40905=>"010001000",
  40906=>"101101010",
  40907=>"011111101",
  40908=>"001010100",
  40909=>"111101010",
  40910=>"111000110",
  40911=>"110110100",
  40912=>"000110100",
  40913=>"001001001",
  40914=>"101111000",
  40915=>"001011110",
  40916=>"010000011",
  40917=>"110000100",
  40918=>"110011100",
  40919=>"001101101",
  40920=>"100100101",
  40921=>"000000100",
  40922=>"010101010",
  40923=>"000001011",
  40924=>"110111011",
  40925=>"001011100",
  40926=>"011100000",
  40927=>"110110100",
  40928=>"000011101",
  40929=>"101111111",
  40930=>"111011110",
  40931=>"001010000",
  40932=>"110010100",
  40933=>"111011001",
  40934=>"111010100",
  40935=>"000010010",
  40936=>"110000000",
  40937=>"111011010",
  40938=>"110111010",
  40939=>"000100001",
  40940=>"110001100",
  40941=>"010101000",
  40942=>"100010100",
  40943=>"011100100",
  40944=>"111010000",
  40945=>"111011011",
  40946=>"100001100",
  40947=>"100001001",
  40948=>"110001100",
  40949=>"110100001",
  40950=>"000000001",
  40951=>"011010011",
  40952=>"010101100",
  40953=>"001000100",
  40954=>"011111100",
  40955=>"011010110",
  40956=>"110011000",
  40957=>"001100100",
  40958=>"010011001",
  40959=>"100101001",
  40960=>"010100101",
  40961=>"101110011",
  40962=>"100011110",
  40963=>"100000111",
  40964=>"101000101",
  40965=>"000001010",
  40966=>"000010101",
  40967=>"010111100",
  40968=>"111111010",
  40969=>"000011011",
  40970=>"010100000",
  40971=>"110111011",
  40972=>"101100101",
  40973=>"101111111",
  40974=>"101100100",
  40975=>"101100110",
  40976=>"111111110",
  40977=>"001100000",
  40978=>"100000011",
  40979=>"101100101",
  40980=>"111110000",
  40981=>"010111001",
  40982=>"100111010",
  40983=>"011010111",
  40984=>"010000100",
  40985=>"010011101",
  40986=>"111111011",
  40987=>"010010000",
  40988=>"101000010",
  40989=>"010000001",
  40990=>"010000001",
  40991=>"011110001",
  40992=>"011000001",
  40993=>"111010110",
  40994=>"111111111",
  40995=>"001000101",
  40996=>"000001000",
  40997=>"001101010",
  40998=>"101001110",
  40999=>"010111111",
  41000=>"110010000",
  41001=>"110001011",
  41002=>"000011111",
  41003=>"011010111",
  41004=>"000011100",
  41005=>"101000000",
  41006=>"011100101",
  41007=>"111110010",
  41008=>"010110111",
  41009=>"110110110",
  41010=>"100100000",
  41011=>"011110110",
  41012=>"100001101",
  41013=>"100011100",
  41014=>"000110100",
  41015=>"001100100",
  41016=>"110011100",
  41017=>"111101010",
  41018=>"111011110",
  41019=>"010000010",
  41020=>"000110011",
  41021=>"100000101",
  41022=>"101101000",
  41023=>"111100010",
  41024=>"101010100",
  41025=>"010010011",
  41026=>"001011010",
  41027=>"100110110",
  41028=>"100010101",
  41029=>"011101111",
  41030=>"001011011",
  41031=>"000000110",
  41032=>"101111001",
  41033=>"010111101",
  41034=>"010100101",
  41035=>"001010000",
  41036=>"101000100",
  41037=>"100001111",
  41038=>"101101000",
  41039=>"000111110",
  41040=>"100010011",
  41041=>"010011100",
  41042=>"010000100",
  41043=>"011001110",
  41044=>"110011010",
  41045=>"111110000",
  41046=>"000001111",
  41047=>"100110111",
  41048=>"101001100",
  41049=>"001001110",
  41050=>"011001010",
  41051=>"111110100",
  41052=>"010110101",
  41053=>"011000110",
  41054=>"111101110",
  41055=>"111100010",
  41056=>"000000011",
  41057=>"100100011",
  41058=>"110101000",
  41059=>"110110101",
  41060=>"010011101",
  41061=>"101010111",
  41062=>"110101111",
  41063=>"011101000",
  41064=>"110100001",
  41065=>"000011010",
  41066=>"110111001",
  41067=>"100101111",
  41068=>"010110001",
  41069=>"101010010",
  41070=>"000111100",
  41071=>"111100100",
  41072=>"000101100",
  41073=>"010000000",
  41074=>"001001110",
  41075=>"011000001",
  41076=>"101000001",
  41077=>"110111101",
  41078=>"101101101",
  41079=>"010100101",
  41080=>"011110010",
  41081=>"111101011",
  41082=>"111110111",
  41083=>"101011100",
  41084=>"011101000",
  41085=>"111001010",
  41086=>"000001111",
  41087=>"101111110",
  41088=>"111100011",
  41089=>"111001100",
  41090=>"001110111",
  41091=>"000010100",
  41092=>"100001101",
  41093=>"110000100",
  41094=>"111100010",
  41095=>"000100011",
  41096=>"110111011",
  41097=>"001001011",
  41098=>"100001000",
  41099=>"110010111",
  41100=>"010111101",
  41101=>"011011111",
  41102=>"001101010",
  41103=>"011100010",
  41104=>"110100110",
  41105=>"000111111",
  41106=>"010001110",
  41107=>"100111010",
  41108=>"111001011",
  41109=>"100000110",
  41110=>"100000001",
  41111=>"011000111",
  41112=>"110011110",
  41113=>"101111100",
  41114=>"110111101",
  41115=>"100110111",
  41116=>"101011111",
  41117=>"001011101",
  41118=>"001101000",
  41119=>"000000100",
  41120=>"001010111",
  41121=>"011100001",
  41122=>"010011110",
  41123=>"101011010",
  41124=>"000011001",
  41125=>"110011100",
  41126=>"011010111",
  41127=>"111100111",
  41128=>"011001001",
  41129=>"011111000",
  41130=>"010000110",
  41131=>"000101010",
  41132=>"001110100",
  41133=>"011100100",
  41134=>"100100101",
  41135=>"100110000",
  41136=>"001110000",
  41137=>"010010001",
  41138=>"000110110",
  41139=>"111000101",
  41140=>"101101001",
  41141=>"100000000",
  41142=>"011010001",
  41143=>"010110001",
  41144=>"010010001",
  41145=>"100100110",
  41146=>"010010011",
  41147=>"100000000",
  41148=>"100111010",
  41149=>"011010110",
  41150=>"001110000",
  41151=>"111111001",
  41152=>"111010101",
  41153=>"001101111",
  41154=>"010110101",
  41155=>"110001101",
  41156=>"111111100",
  41157=>"100100110",
  41158=>"100111110",
  41159=>"111000101",
  41160=>"100110001",
  41161=>"000001110",
  41162=>"111111011",
  41163=>"111011011",
  41164=>"111011100",
  41165=>"011001110",
  41166=>"100011110",
  41167=>"000000011",
  41168=>"001001101",
  41169=>"001110101",
  41170=>"110110011",
  41171=>"001110101",
  41172=>"110000110",
  41173=>"111010000",
  41174=>"111100101",
  41175=>"100100111",
  41176=>"001100010",
  41177=>"000011011",
  41178=>"101101111",
  41179=>"100110001",
  41180=>"110110000",
  41181=>"010100100",
  41182=>"100001010",
  41183=>"111001110",
  41184=>"101001011",
  41185=>"000100100",
  41186=>"001101100",
  41187=>"000100111",
  41188=>"000000000",
  41189=>"101010110",
  41190=>"110000001",
  41191=>"110100001",
  41192=>"110101111",
  41193=>"100100000",
  41194=>"000010110",
  41195=>"111101100",
  41196=>"001100000",
  41197=>"101010010",
  41198=>"101001000",
  41199=>"110011111",
  41200=>"010011010",
  41201=>"100110101",
  41202=>"000101100",
  41203=>"100100111",
  41204=>"000001010",
  41205=>"111101100",
  41206=>"101011000",
  41207=>"011100000",
  41208=>"110010111",
  41209=>"110100000",
  41210=>"011011011",
  41211=>"110110110",
  41212=>"111100101",
  41213=>"011110000",
  41214=>"101011100",
  41215=>"011010011",
  41216=>"101010010",
  41217=>"111101111",
  41218=>"101000111",
  41219=>"110000010",
  41220=>"011000100",
  41221=>"100111010",
  41222=>"000101111",
  41223=>"011000011",
  41224=>"110000011",
  41225=>"101010111",
  41226=>"000010010",
  41227=>"101110101",
  41228=>"101001110",
  41229=>"001110101",
  41230=>"001011001",
  41231=>"001010001",
  41232=>"000110100",
  41233=>"101101111",
  41234=>"011110110",
  41235=>"101011000",
  41236=>"111011111",
  41237=>"001000101",
  41238=>"000110001",
  41239=>"110001110",
  41240=>"101110110",
  41241=>"101011011",
  41242=>"010011000",
  41243=>"010100011",
  41244=>"110101111",
  41245=>"010010000",
  41246=>"010111100",
  41247=>"111111001",
  41248=>"111000000",
  41249=>"000110111",
  41250=>"000011000",
  41251=>"111000011",
  41252=>"111100010",
  41253=>"001011000",
  41254=>"010000100",
  41255=>"011100101",
  41256=>"011111001",
  41257=>"010011000",
  41258=>"101010100",
  41259=>"001000110",
  41260=>"110011010",
  41261=>"011001101",
  41262=>"011101000",
  41263=>"010101011",
  41264=>"100011011",
  41265=>"111001011",
  41266=>"000111100",
  41267=>"001000011",
  41268=>"011101111",
  41269=>"000001110",
  41270=>"001110110",
  41271=>"101100001",
  41272=>"010000111",
  41273=>"000111100",
  41274=>"000001011",
  41275=>"101001100",
  41276=>"000000100",
  41277=>"001100110",
  41278=>"001010000",
  41279=>"001001010",
  41280=>"001110110",
  41281=>"000110100",
  41282=>"100000111",
  41283=>"111110100",
  41284=>"111010100",
  41285=>"110010011",
  41286=>"111100001",
  41287=>"101111000",
  41288=>"111011011",
  41289=>"100111100",
  41290=>"110010010",
  41291=>"101000101",
  41292=>"111011000",
  41293=>"011001100",
  41294=>"000101001",
  41295=>"100111000",
  41296=>"100001110",
  41297=>"010101111",
  41298=>"001010000",
  41299=>"101101100",
  41300=>"011000001",
  41301=>"001111111",
  41302=>"101000000",
  41303=>"001000111",
  41304=>"001000001",
  41305=>"001101100",
  41306=>"000101001",
  41307=>"101000011",
  41308=>"101000111",
  41309=>"100100110",
  41310=>"101011010",
  41311=>"000010100",
  41312=>"001010011",
  41313=>"111001100",
  41314=>"110101111",
  41315=>"011011011",
  41316=>"000000000",
  41317=>"001110000",
  41318=>"101110011",
  41319=>"000111001",
  41320=>"111000110",
  41321=>"010110001",
  41322=>"101001101",
  41323=>"110000010",
  41324=>"001111000",
  41325=>"011011110",
  41326=>"000000101",
  41327=>"101010101",
  41328=>"100111010",
  41329=>"000001111",
  41330=>"000000101",
  41331=>"100110111",
  41332=>"101100000",
  41333=>"001000010",
  41334=>"110101110",
  41335=>"001010110",
  41336=>"101111101",
  41337=>"101100011",
  41338=>"110111111",
  41339=>"100001101",
  41340=>"111001110",
  41341=>"001110000",
  41342=>"111000111",
  41343=>"001101001",
  41344=>"011001100",
  41345=>"000010011",
  41346=>"101011001",
  41347=>"110001000",
  41348=>"100001110",
  41349=>"000011110",
  41350=>"011010000",
  41351=>"001110110",
  41352=>"000100111",
  41353=>"000001000",
  41354=>"101011101",
  41355=>"101010001",
  41356=>"100010010",
  41357=>"010100111",
  41358=>"010110100",
  41359=>"101011110",
  41360=>"111101001",
  41361=>"110001001",
  41362=>"111100010",
  41363=>"000000100",
  41364=>"000111110",
  41365=>"110011100",
  41366=>"011111111",
  41367=>"111110111",
  41368=>"100110111",
  41369=>"010001010",
  41370=>"010001011",
  41371=>"010100011",
  41372=>"111111101",
  41373=>"011111101",
  41374=>"101110111",
  41375=>"101100110",
  41376=>"101101001",
  41377=>"101101010",
  41378=>"110100100",
  41379=>"110111111",
  41380=>"001101011",
  41381=>"001000101",
  41382=>"001101000",
  41383=>"110010110",
  41384=>"100100011",
  41385=>"101101110",
  41386=>"001000000",
  41387=>"000101110",
  41388=>"011101110",
  41389=>"001100110",
  41390=>"110101011",
  41391=>"111111111",
  41392=>"101110111",
  41393=>"010001101",
  41394=>"001010001",
  41395=>"111101110",
  41396=>"010101010",
  41397=>"111101011",
  41398=>"100111100",
  41399=>"111101000",
  41400=>"101001010",
  41401=>"000110100",
  41402=>"000100101",
  41403=>"000011001",
  41404=>"100001011",
  41405=>"000011011",
  41406=>"111001101",
  41407=>"100010111",
  41408=>"001110100",
  41409=>"000000011",
  41410=>"001010001",
  41411=>"110011111",
  41412=>"001001111",
  41413=>"010100110",
  41414=>"010100011",
  41415=>"110010000",
  41416=>"110000000",
  41417=>"111001100",
  41418=>"100111001",
  41419=>"001111101",
  41420=>"111001101",
  41421=>"000110110",
  41422=>"010001011",
  41423=>"111110111",
  41424=>"010000011",
  41425=>"101110010",
  41426=>"101000111",
  41427=>"000101101",
  41428=>"111101000",
  41429=>"000010110",
  41430=>"110000101",
  41431=>"110111011",
  41432=>"101001001",
  41433=>"101010001",
  41434=>"100100110",
  41435=>"001000100",
  41436=>"111101111",
  41437=>"001010010",
  41438=>"000010010",
  41439=>"100101110",
  41440=>"101011011",
  41441=>"000000110",
  41442=>"101010010",
  41443=>"110100001",
  41444=>"111111110",
  41445=>"100100000",
  41446=>"111000011",
  41447=>"101110000",
  41448=>"000010000",
  41449=>"111100110",
  41450=>"010100110",
  41451=>"001111111",
  41452=>"011110001",
  41453=>"000101110",
  41454=>"100000100",
  41455=>"100010101",
  41456=>"010110100",
  41457=>"010011110",
  41458=>"111000000",
  41459=>"100011101",
  41460=>"110100111",
  41461=>"001100101",
  41462=>"010001100",
  41463=>"111000000",
  41464=>"101011010",
  41465=>"110111100",
  41466=>"011110001",
  41467=>"110000110",
  41468=>"111000010",
  41469=>"001011100",
  41470=>"111110110",
  41471=>"011001010",
  41472=>"111001101",
  41473=>"010111110",
  41474=>"100001010",
  41475=>"011011111",
  41476=>"111111101",
  41477=>"000101001",
  41478=>"111010111",
  41479=>"111011011",
  41480=>"111000110",
  41481=>"010011101",
  41482=>"110101010",
  41483=>"110111101",
  41484=>"110100000",
  41485=>"010110101",
  41486=>"110110111",
  41487=>"101001101",
  41488=>"000011101",
  41489=>"000110011",
  41490=>"011010010",
  41491=>"110111100",
  41492=>"101101111",
  41493=>"110000000",
  41494=>"001001111",
  41495=>"111001011",
  41496=>"111001001",
  41497=>"110110111",
  41498=>"001101111",
  41499=>"111100010",
  41500=>"000001011",
  41501=>"110010011",
  41502=>"000000010",
  41503=>"100000001",
  41504=>"111100110",
  41505=>"100000100",
  41506=>"110011110",
  41507=>"011111001",
  41508=>"000101000",
  41509=>"101000110",
  41510=>"101101110",
  41511=>"001100010",
  41512=>"001011110",
  41513=>"011001110",
  41514=>"001111010",
  41515=>"011110011",
  41516=>"001110011",
  41517=>"000010111",
  41518=>"110101100",
  41519=>"100111000",
  41520=>"100001001",
  41521=>"100100100",
  41522=>"110010101",
  41523=>"000101000",
  41524=>"111110000",
  41525=>"010110111",
  41526=>"110011011",
  41527=>"110010111",
  41528=>"111101001",
  41529=>"010001011",
  41530=>"001001011",
  41531=>"110010001",
  41532=>"011111100",
  41533=>"110110111",
  41534=>"000110011",
  41535=>"100101111",
  41536=>"001111101",
  41537=>"010001011",
  41538=>"001101111",
  41539=>"110010010",
  41540=>"111111111",
  41541=>"110001110",
  41542=>"011001111",
  41543=>"111010000",
  41544=>"001011110",
  41545=>"111111011",
  41546=>"000010000",
  41547=>"100110100",
  41548=>"000101101",
  41549=>"001101001",
  41550=>"000010000",
  41551=>"100011010",
  41552=>"100000011",
  41553=>"010000000",
  41554=>"011111011",
  41555=>"110110101",
  41556=>"010010110",
  41557=>"000000100",
  41558=>"101111011",
  41559=>"100011111",
  41560=>"111011111",
  41561=>"010010010",
  41562=>"011110011",
  41563=>"001100010",
  41564=>"101111111",
  41565=>"000110001",
  41566=>"001110001",
  41567=>"110011100",
  41568=>"100000111",
  41569=>"110101111",
  41570=>"000101011",
  41571=>"101001111",
  41572=>"000110000",
  41573=>"100101010",
  41574=>"011110001",
  41575=>"111111001",
  41576=>"001101111",
  41577=>"101100000",
  41578=>"000111010",
  41579=>"111000010",
  41580=>"011001100",
  41581=>"000101111",
  41582=>"101011101",
  41583=>"111011010",
  41584=>"011011101",
  41585=>"101000101",
  41586=>"110011000",
  41587=>"100111111",
  41588=>"010000011",
  41589=>"011000010",
  41590=>"110011110",
  41591=>"100011110",
  41592=>"011101001",
  41593=>"001000110",
  41594=>"110110101",
  41595=>"111010111",
  41596=>"001000100",
  41597=>"100111100",
  41598=>"001000101",
  41599=>"000100011",
  41600=>"010101100",
  41601=>"001100000",
  41602=>"001100111",
  41603=>"101011110",
  41604=>"100111111",
  41605=>"000010100",
  41606=>"000100101",
  41607=>"100101101",
  41608=>"100100001",
  41609=>"001101100",
  41610=>"011010111",
  41611=>"011110110",
  41612=>"011011011",
  41613=>"010101101",
  41614=>"101001000",
  41615=>"011101001",
  41616=>"000100010",
  41617=>"101011011",
  41618=>"101011001",
  41619=>"100000111",
  41620=>"000000111",
  41621=>"101110101",
  41622=>"001000011",
  41623=>"110110010",
  41624=>"011001010",
  41625=>"000110000",
  41626=>"001010111",
  41627=>"111001100",
  41628=>"000111010",
  41629=>"010110010",
  41630=>"000011001",
  41631=>"111000011",
  41632=>"110100001",
  41633=>"011111101",
  41634=>"001001100",
  41635=>"010101101",
  41636=>"000100010",
  41637=>"101011100",
  41638=>"001010000",
  41639=>"000100001",
  41640=>"001010000",
  41641=>"100011010",
  41642=>"011010111",
  41643=>"010001111",
  41644=>"011110001",
  41645=>"000100110",
  41646=>"101001001",
  41647=>"101110110",
  41648=>"110010111",
  41649=>"100100111",
  41650=>"011010101",
  41651=>"011000010",
  41652=>"101001010",
  41653=>"001110110",
  41654=>"000010110",
  41655=>"001011111",
  41656=>"011100110",
  41657=>"000111110",
  41658=>"011010011",
  41659=>"000010111",
  41660=>"001110111",
  41661=>"011110000",
  41662=>"010011010",
  41663=>"110010001",
  41664=>"111001010",
  41665=>"100100111",
  41666=>"000111101",
  41667=>"011101111",
  41668=>"001111011",
  41669=>"001111001",
  41670=>"001101100",
  41671=>"110110101",
  41672=>"111111111",
  41673=>"011111110",
  41674=>"110100110",
  41675=>"011000001",
  41676=>"000100010",
  41677=>"001000101",
  41678=>"001111100",
  41679=>"011111011",
  41680=>"110101111",
  41681=>"000000111",
  41682=>"111010110",
  41683=>"010100011",
  41684=>"101000000",
  41685=>"101000101",
  41686=>"001110111",
  41687=>"010111100",
  41688=>"111111010",
  41689=>"010000101",
  41690=>"000110000",
  41691=>"111011100",
  41692=>"110110011",
  41693=>"001000001",
  41694=>"000001101",
  41695=>"101011010",
  41696=>"111100011",
  41697=>"100000001",
  41698=>"000110000",
  41699=>"001111100",
  41700=>"000010000",
  41701=>"010000010",
  41702=>"110001000",
  41703=>"110111111",
  41704=>"111001111",
  41705=>"101010000",
  41706=>"000000101",
  41707=>"010110101",
  41708=>"010010010",
  41709=>"000100011",
  41710=>"100010001",
  41711=>"010001000",
  41712=>"010100111",
  41713=>"011100111",
  41714=>"011101101",
  41715=>"110000100",
  41716=>"011001000",
  41717=>"001101100",
  41718=>"001011100",
  41719=>"000110010",
  41720=>"011110000",
  41721=>"000010000",
  41722=>"001100001",
  41723=>"011110001",
  41724=>"110110001",
  41725=>"000110111",
  41726=>"110100101",
  41727=>"000101011",
  41728=>"001001001",
  41729=>"101100101",
  41730=>"111111011",
  41731=>"010001000",
  41732=>"000000011",
  41733=>"101111111",
  41734=>"001100101",
  41735=>"110000000",
  41736=>"000101100",
  41737=>"010110010",
  41738=>"110101011",
  41739=>"110000011",
  41740=>"011100100",
  41741=>"100101100",
  41742=>"000010101",
  41743=>"101000100",
  41744=>"000101110",
  41745=>"000010100",
  41746=>"100100011",
  41747=>"110110001",
  41748=>"010001011",
  41749=>"010000001",
  41750=>"111101101",
  41751=>"010111010",
  41752=>"011110001",
  41753=>"101100001",
  41754=>"000100111",
  41755=>"111011011",
  41756=>"101010011",
  41757=>"110110100",
  41758=>"000000101",
  41759=>"111111011",
  41760=>"100010011",
  41761=>"100010010",
  41762=>"011011110",
  41763=>"110000111",
  41764=>"001010111",
  41765=>"101011001",
  41766=>"010011010",
  41767=>"111101010",
  41768=>"010101110",
  41769=>"010100001",
  41770=>"111100011",
  41771=>"110010000",
  41772=>"010001111",
  41773=>"111111101",
  41774=>"110110111",
  41775=>"111101111",
  41776=>"001001001",
  41777=>"010010100",
  41778=>"100010001",
  41779=>"000100010",
  41780=>"001000010",
  41781=>"100000000",
  41782=>"111111111",
  41783=>"010100001",
  41784=>"110100011",
  41785=>"000101110",
  41786=>"101101011",
  41787=>"001111000",
  41788=>"000011011",
  41789=>"000011000",
  41790=>"010111110",
  41791=>"111001100",
  41792=>"100101010",
  41793=>"111011011",
  41794=>"100100010",
  41795=>"110110110",
  41796=>"001101101",
  41797=>"010001100",
  41798=>"101000011",
  41799=>"011111010",
  41800=>"000101110",
  41801=>"000101101",
  41802=>"001110100",
  41803=>"001100000",
  41804=>"100110000",
  41805=>"111011011",
  41806=>"011111010",
  41807=>"000100100",
  41808=>"000111001",
  41809=>"000111101",
  41810=>"011000011",
  41811=>"111110011",
  41812=>"000010010",
  41813=>"000101101",
  41814=>"011100101",
  41815=>"110110110",
  41816=>"011001010",
  41817=>"111111111",
  41818=>"000011100",
  41819=>"111111111",
  41820=>"101110100",
  41821=>"001001000",
  41822=>"001110010",
  41823=>"101001011",
  41824=>"110111011",
  41825=>"100001111",
  41826=>"100010000",
  41827=>"010000000",
  41828=>"111000010",
  41829=>"000010010",
  41830=>"101010001",
  41831=>"100101110",
  41832=>"111001001",
  41833=>"101011001",
  41834=>"011100000",
  41835=>"101001100",
  41836=>"111111011",
  41837=>"011011011",
  41838=>"010011011",
  41839=>"011001100",
  41840=>"110001010",
  41841=>"101111111",
  41842=>"010110111",
  41843=>"111001011",
  41844=>"001111011",
  41845=>"000010111",
  41846=>"101011010",
  41847=>"000010010",
  41848=>"001001011",
  41849=>"100110101",
  41850=>"011111010",
  41851=>"000000011",
  41852=>"000101011",
  41853=>"011001000",
  41854=>"011011110",
  41855=>"010001101",
  41856=>"100110000",
  41857=>"101000101",
  41858=>"111111001",
  41859=>"101010101",
  41860=>"110000100",
  41861=>"100111010",
  41862=>"111001001",
  41863=>"111110111",
  41864=>"100000010",
  41865=>"100111000",
  41866=>"010110000",
  41867=>"111111111",
  41868=>"001000010",
  41869=>"010001011",
  41870=>"101101110",
  41871=>"010001101",
  41872=>"111101010",
  41873=>"100000011",
  41874=>"010000000",
  41875=>"101111110",
  41876=>"011111110",
  41877=>"001110010",
  41878=>"000100010",
  41879=>"110000111",
  41880=>"111111111",
  41881=>"011101110",
  41882=>"000111100",
  41883=>"100011011",
  41884=>"100011100",
  41885=>"101000010",
  41886=>"000000000",
  41887=>"110011110",
  41888=>"010010011",
  41889=>"110110000",
  41890=>"001000010",
  41891=>"010001011",
  41892=>"000000110",
  41893=>"111000110",
  41894=>"000000010",
  41895=>"100011111",
  41896=>"000110001",
  41897=>"100101000",
  41898=>"011100011",
  41899=>"100010110",
  41900=>"100010111",
  41901=>"011111001",
  41902=>"000101100",
  41903=>"110010001",
  41904=>"110000000",
  41905=>"011111011",
  41906=>"110000001",
  41907=>"010101011",
  41908=>"000111001",
  41909=>"000101001",
  41910=>"000001000",
  41911=>"000011000",
  41912=>"001100000",
  41913=>"100111111",
  41914=>"100111010",
  41915=>"110001001",
  41916=>"110101110",
  41917=>"001000000",
  41918=>"101001010",
  41919=>"111110111",
  41920=>"100111110",
  41921=>"100101101",
  41922=>"100101000",
  41923=>"111100011",
  41924=>"001011010",
  41925=>"000101000",
  41926=>"110100000",
  41927=>"001001110",
  41928=>"001000111",
  41929=>"101111001",
  41930=>"010001000",
  41931=>"111000010",
  41932=>"110000110",
  41933=>"001100111",
  41934=>"111111111",
  41935=>"100000000",
  41936=>"101001100",
  41937=>"100011011",
  41938=>"000010100",
  41939=>"000001100",
  41940=>"000011000",
  41941=>"100000111",
  41942=>"000011001",
  41943=>"111111011",
  41944=>"011110100",
  41945=>"001110101",
  41946=>"000010111",
  41947=>"001011010",
  41948=>"011011001",
  41949=>"011001000",
  41950=>"000011101",
  41951=>"000011000",
  41952=>"111111111",
  41953=>"110010110",
  41954=>"101110101",
  41955=>"000101010",
  41956=>"000000010",
  41957=>"000011000",
  41958=>"111100000",
  41959=>"101111001",
  41960=>"000101000",
  41961=>"111111001",
  41962=>"000100010",
  41963=>"110011101",
  41964=>"111001110",
  41965=>"010000010",
  41966=>"001101000",
  41967=>"001010110",
  41968=>"111110101",
  41969=>"100110010",
  41970=>"000100100",
  41971=>"101011110",
  41972=>"100111110",
  41973=>"000110011",
  41974=>"000011001",
  41975=>"110011111",
  41976=>"100001110",
  41977=>"000110000",
  41978=>"110011111",
  41979=>"011000001",
  41980=>"010110111",
  41981=>"110011100",
  41982=>"000000001",
  41983=>"011011101",
  41984=>"110110101",
  41985=>"110111001",
  41986=>"110111111",
  41987=>"001011101",
  41988=>"001001001",
  41989=>"110100010",
  41990=>"000100010",
  41991=>"011010011",
  41992=>"111010111",
  41993=>"110011111",
  41994=>"110001001",
  41995=>"000000111",
  41996=>"000100011",
  41997=>"100010100",
  41998=>"001100010",
  41999=>"001010110",
  42000=>"110100010",
  42001=>"000110011",
  42002=>"010111100",
  42003=>"010110111",
  42004=>"010010000",
  42005=>"100010110",
  42006=>"110010011",
  42007=>"010010010",
  42008=>"101101011",
  42009=>"110101001",
  42010=>"011000100",
  42011=>"110000000",
  42012=>"011101001",
  42013=>"000000111",
  42014=>"001001000",
  42015=>"111010011",
  42016=>"111110110",
  42017=>"011110100",
  42018=>"011110010",
  42019=>"011010000",
  42020=>"001101010",
  42021=>"001110011",
  42022=>"111101010",
  42023=>"110101111",
  42024=>"000011000",
  42025=>"110110101",
  42026=>"010100110",
  42027=>"110010101",
  42028=>"010100101",
  42029=>"001110001",
  42030=>"001110101",
  42031=>"010001010",
  42032=>"011100111",
  42033=>"100111010",
  42034=>"111010110",
  42035=>"100101101",
  42036=>"111110111",
  42037=>"010100110",
  42038=>"000110111",
  42039=>"101111110",
  42040=>"001010111",
  42041=>"000010010",
  42042=>"100000110",
  42043=>"001000000",
  42044=>"011101010",
  42045=>"001100110",
  42046=>"000110011",
  42047=>"000101000",
  42048=>"001111111",
  42049=>"111110000",
  42050=>"111001110",
  42051=>"000001010",
  42052=>"101010011",
  42053=>"000010000",
  42054=>"010000101",
  42055=>"001001111",
  42056=>"111101011",
  42057=>"000000000",
  42058=>"110011010",
  42059=>"011011110",
  42060=>"110110100",
  42061=>"110010001",
  42062=>"001011010",
  42063=>"111010000",
  42064=>"001010100",
  42065=>"110111000",
  42066=>"001000011",
  42067=>"010110000",
  42068=>"110111100",
  42069=>"111100111",
  42070=>"010000001",
  42071=>"000001010",
  42072=>"111111000",
  42073=>"001100101",
  42074=>"110111111",
  42075=>"101001110",
  42076=>"101111001",
  42077=>"100100100",
  42078=>"100110011",
  42079=>"010001010",
  42080=>"001101001",
  42081=>"101110101",
  42082=>"111010101",
  42083=>"001001100",
  42084=>"000110101",
  42085=>"100101111",
  42086=>"011100001",
  42087=>"011100001",
  42088=>"100000111",
  42089=>"010111011",
  42090=>"011101110",
  42091=>"100110001",
  42092=>"111010111",
  42093=>"010100101",
  42094=>"100110000",
  42095=>"110110010",
  42096=>"001001101",
  42097=>"110000100",
  42098=>"011010101",
  42099=>"100101111",
  42100=>"001001010",
  42101=>"111111101",
  42102=>"001110011",
  42103=>"001001010",
  42104=>"001111011",
  42105=>"001111101",
  42106=>"110001000",
  42107=>"111011000",
  42108=>"110011000",
  42109=>"011100111",
  42110=>"000010111",
  42111=>"000101001",
  42112=>"101110011",
  42113=>"100100100",
  42114=>"100100000",
  42115=>"110001101",
  42116=>"101101110",
  42117=>"111110011",
  42118=>"110101011",
  42119=>"001000111",
  42120=>"011000100",
  42121=>"011000100",
  42122=>"010011100",
  42123=>"010110000",
  42124=>"001110011",
  42125=>"100011010",
  42126=>"111100110",
  42127=>"111001010",
  42128=>"100000001",
  42129=>"001001101",
  42130=>"110110001",
  42131=>"011101000",
  42132=>"000001101",
  42133=>"001101001",
  42134=>"010010100",
  42135=>"110100000",
  42136=>"011100110",
  42137=>"111100001",
  42138=>"010000100",
  42139=>"111011011",
  42140=>"011110001",
  42141=>"101011101",
  42142=>"111111010",
  42143=>"111101010",
  42144=>"101010011",
  42145=>"000100111",
  42146=>"001001011",
  42147=>"001010101",
  42148=>"010111001",
  42149=>"011111110",
  42150=>"110010001",
  42151=>"000101000",
  42152=>"101000100",
  42153=>"111001010",
  42154=>"111101111",
  42155=>"011110010",
  42156=>"111111101",
  42157=>"000111001",
  42158=>"001001010",
  42159=>"000011001",
  42160=>"011100010",
  42161=>"100111010",
  42162=>"000110101",
  42163=>"100011100",
  42164=>"111000011",
  42165=>"010010101",
  42166=>"011110111",
  42167=>"110111110",
  42168=>"001011000",
  42169=>"111111010",
  42170=>"001001100",
  42171=>"000000001",
  42172=>"010101111",
  42173=>"001110100",
  42174=>"011101110",
  42175=>"000010011",
  42176=>"001011100",
  42177=>"111000010",
  42178=>"010011110",
  42179=>"111100001",
  42180=>"101011111",
  42181=>"100000111",
  42182=>"000100111",
  42183=>"101011001",
  42184=>"110111000",
  42185=>"000111001",
  42186=>"111101010",
  42187=>"001000010",
  42188=>"111011010",
  42189=>"101110001",
  42190=>"001010110",
  42191=>"111111001",
  42192=>"010000100",
  42193=>"000011010",
  42194=>"001001011",
  42195=>"100001110",
  42196=>"111010011",
  42197=>"111000001",
  42198=>"000101000",
  42199=>"011010110",
  42200=>"001111111",
  42201=>"110010110",
  42202=>"101101110",
  42203=>"100000110",
  42204=>"101001101",
  42205=>"001111001",
  42206=>"001000101",
  42207=>"000010110",
  42208=>"111110011",
  42209=>"000110000",
  42210=>"101001101",
  42211=>"000011000",
  42212=>"011011100",
  42213=>"010101011",
  42214=>"011110100",
  42215=>"000110101",
  42216=>"110010001",
  42217=>"010110101",
  42218=>"111110011",
  42219=>"101001110",
  42220=>"101100000",
  42221=>"000101101",
  42222=>"111001000",
  42223=>"101001110",
  42224=>"001000110",
  42225=>"000011101",
  42226=>"110001110",
  42227=>"111011100",
  42228=>"111000011",
  42229=>"100100001",
  42230=>"101110101",
  42231=>"111111111",
  42232=>"100101111",
  42233=>"000010010",
  42234=>"110001001",
  42235=>"011011100",
  42236=>"101000010",
  42237=>"001010001",
  42238=>"001001100",
  42239=>"000111110",
  42240=>"111101011",
  42241=>"111100100",
  42242=>"011101110",
  42243=>"000111010",
  42244=>"011111101",
  42245=>"011001110",
  42246=>"100011001",
  42247=>"000011011",
  42248=>"111111011",
  42249=>"001101111",
  42250=>"111100010",
  42251=>"111110110",
  42252=>"001110110",
  42253=>"011101100",
  42254=>"001001110",
  42255=>"000100001",
  42256=>"111000010",
  42257=>"111111111",
  42258=>"011011001",
  42259=>"111011111",
  42260=>"001110010",
  42261=>"001011001",
  42262=>"110100111",
  42263=>"001111011",
  42264=>"101110101",
  42265=>"100010101",
  42266=>"100101101",
  42267=>"110111100",
  42268=>"101011001",
  42269=>"010100001",
  42270=>"110011110",
  42271=>"101110101",
  42272=>"010001001",
  42273=>"101101111",
  42274=>"000110110",
  42275=>"111111001",
  42276=>"111101001",
  42277=>"111010101",
  42278=>"101010000",
  42279=>"100001110",
  42280=>"101111000",
  42281=>"010000100",
  42282=>"011101101",
  42283=>"011101111",
  42284=>"110010010",
  42285=>"011000000",
  42286=>"100110011",
  42287=>"000100100",
  42288=>"010001101",
  42289=>"011011101",
  42290=>"010101111",
  42291=>"111110100",
  42292=>"110101000",
  42293=>"101001101",
  42294=>"111110000",
  42295=>"100001010",
  42296=>"010011100",
  42297=>"111111000",
  42298=>"001000010",
  42299=>"101101101",
  42300=>"111011101",
  42301=>"110001110",
  42302=>"100100100",
  42303=>"100011011",
  42304=>"010110010",
  42305=>"011011010",
  42306=>"000100000",
  42307=>"011110011",
  42308=>"011010001",
  42309=>"111000010",
  42310=>"100001001",
  42311=>"010011101",
  42312=>"010101000",
  42313=>"100100001",
  42314=>"011100101",
  42315=>"100100100",
  42316=>"010001100",
  42317=>"001100010",
  42318=>"111111101",
  42319=>"000111011",
  42320=>"000000000",
  42321=>"010110000",
  42322=>"001001001",
  42323=>"010011000",
  42324=>"000100001",
  42325=>"010100001",
  42326=>"101010110",
  42327=>"110000111",
  42328=>"010111011",
  42329=>"000000011",
  42330=>"011101101",
  42331=>"011011010",
  42332=>"110100010",
  42333=>"001010000",
  42334=>"001011111",
  42335=>"000100101",
  42336=>"110101110",
  42337=>"101000101",
  42338=>"100111100",
  42339=>"011111100",
  42340=>"001100100",
  42341=>"011111100",
  42342=>"101110100",
  42343=>"001011001",
  42344=>"000101001",
  42345=>"001110011",
  42346=>"110000101",
  42347=>"010001110",
  42348=>"100011011",
  42349=>"101000101",
  42350=>"011101111",
  42351=>"111000110",
  42352=>"111011000",
  42353=>"010110011",
  42354=>"110110000",
  42355=>"110100011",
  42356=>"001000110",
  42357=>"001101011",
  42358=>"001011110",
  42359=>"101100000",
  42360=>"110100110",
  42361=>"110010100",
  42362=>"100100011",
  42363=>"111011111",
  42364=>"101010110",
  42365=>"001001011",
  42366=>"000010101",
  42367=>"010010101",
  42368=>"100110100",
  42369=>"010000111",
  42370=>"010100001",
  42371=>"010001101",
  42372=>"111001010",
  42373=>"010011011",
  42374=>"010001000",
  42375=>"001110100",
  42376=>"100001011",
  42377=>"000010000",
  42378=>"011011011",
  42379=>"111100011",
  42380=>"110000000",
  42381=>"100011010",
  42382=>"101111111",
  42383=>"110000100",
  42384=>"011000011",
  42385=>"111011001",
  42386=>"100111001",
  42387=>"111000101",
  42388=>"010011111",
  42389=>"110000000",
  42390=>"000010000",
  42391=>"101000111",
  42392=>"110011011",
  42393=>"101000100",
  42394=>"011100011",
  42395=>"001100001",
  42396=>"011101010",
  42397=>"011101110",
  42398=>"011101000",
  42399=>"100010101",
  42400=>"100100100",
  42401=>"001011011",
  42402=>"011000111",
  42403=>"110111011",
  42404=>"101101110",
  42405=>"001001001",
  42406=>"001000010",
  42407=>"110100000",
  42408=>"010000001",
  42409=>"101111010",
  42410=>"111011001",
  42411=>"001100010",
  42412=>"101100101",
  42413=>"000000011",
  42414=>"110011110",
  42415=>"101100110",
  42416=>"100111100",
  42417=>"011000000",
  42418=>"100010111",
  42419=>"000001110",
  42420=>"101010110",
  42421=>"001101000",
  42422=>"101010110",
  42423=>"011100010",
  42424=>"100111011",
  42425=>"010110001",
  42426=>"011101010",
  42427=>"101110010",
  42428=>"101001110",
  42429=>"001110100",
  42430=>"110110111",
  42431=>"111101111",
  42432=>"001110101",
  42433=>"100010011",
  42434=>"000000101",
  42435=>"110001000",
  42436=>"011001001",
  42437=>"110001100",
  42438=>"100110101",
  42439=>"111101111",
  42440=>"011001111",
  42441=>"110101111",
  42442=>"001101101",
  42443=>"110110100",
  42444=>"010101111",
  42445=>"010101010",
  42446=>"000001111",
  42447=>"111010111",
  42448=>"011110000",
  42449=>"000101111",
  42450=>"101001011",
  42451=>"100001001",
  42452=>"010100001",
  42453=>"010001011",
  42454=>"101000111",
  42455=>"010001001",
  42456=>"000001110",
  42457=>"010001111",
  42458=>"111000011",
  42459=>"011000001",
  42460=>"010101100",
  42461=>"011111001",
  42462=>"010110110",
  42463=>"101111101",
  42464=>"111101110",
  42465=>"001000101",
  42466=>"100001110",
  42467=>"101011001",
  42468=>"001111011",
  42469=>"011000000",
  42470=>"001111000",
  42471=>"001001100",
  42472=>"111011100",
  42473=>"000001111",
  42474=>"101111100",
  42475=>"001111010",
  42476=>"111111000",
  42477=>"110101100",
  42478=>"110000111",
  42479=>"111111110",
  42480=>"110010000",
  42481=>"101101111",
  42482=>"011001110",
  42483=>"010111011",
  42484=>"011100101",
  42485=>"001101001",
  42486=>"011101110",
  42487=>"101101010",
  42488=>"100000100",
  42489=>"111101011",
  42490=>"111011100",
  42491=>"111100111",
  42492=>"011101010",
  42493=>"100100101",
  42494=>"000011000",
  42495=>"000011000",
  42496=>"100000110",
  42497=>"101110111",
  42498=>"100011000",
  42499=>"101011000",
  42500=>"011110101",
  42501=>"101110110",
  42502=>"100100000",
  42503=>"000010011",
  42504=>"000000010",
  42505=>"110110000",
  42506=>"000101011",
  42507=>"111100110",
  42508=>"110101100",
  42509=>"101000101",
  42510=>"110001001",
  42511=>"100010011",
  42512=>"011110010",
  42513=>"000111100",
  42514=>"111111111",
  42515=>"010111000",
  42516=>"111010111",
  42517=>"011001000",
  42518=>"101001011",
  42519=>"010011111",
  42520=>"110110111",
  42521=>"111101110",
  42522=>"111011011",
  42523=>"001000100",
  42524=>"011100101",
  42525=>"101111111",
  42526=>"100100011",
  42527=>"010011010",
  42528=>"111001110",
  42529=>"101100001",
  42530=>"111010000",
  42531=>"101110011",
  42532=>"101111110",
  42533=>"110111001",
  42534=>"110101100",
  42535=>"101011111",
  42536=>"101100000",
  42537=>"110100101",
  42538=>"011111001",
  42539=>"110010101",
  42540=>"001000111",
  42541=>"111111011",
  42542=>"010111000",
  42543=>"111000001",
  42544=>"010111001",
  42545=>"110111111",
  42546=>"110000010",
  42547=>"010100000",
  42548=>"110011011",
  42549=>"011011011",
  42550=>"101101001",
  42551=>"101101000",
  42552=>"011110111",
  42553=>"101111100",
  42554=>"000111111",
  42555=>"010011111",
  42556=>"000101110",
  42557=>"011110011",
  42558=>"111110111",
  42559=>"011001111",
  42560=>"001110100",
  42561=>"100101010",
  42562=>"101010111",
  42563=>"110011100",
  42564=>"011100110",
  42565=>"001111011",
  42566=>"110001011",
  42567=>"001101011",
  42568=>"111111010",
  42569=>"000111000",
  42570=>"011010011",
  42571=>"001010111",
  42572=>"101000000",
  42573=>"000111111",
  42574=>"100111011",
  42575=>"011011111",
  42576=>"011101110",
  42577=>"100101010",
  42578=>"000001110",
  42579=>"000111100",
  42580=>"001100110",
  42581=>"100000001",
  42582=>"000101101",
  42583=>"111110100",
  42584=>"100000011",
  42585=>"111000111",
  42586=>"111011001",
  42587=>"000001010",
  42588=>"101011000",
  42589=>"111111110",
  42590=>"110000111",
  42591=>"101011100",
  42592=>"110100111",
  42593=>"010010101",
  42594=>"100101000",
  42595=>"001010100",
  42596=>"000100011",
  42597=>"110000100",
  42598=>"011111000",
  42599=>"111001110",
  42600=>"100111011",
  42601=>"011101010",
  42602=>"110010110",
  42603=>"100100000",
  42604=>"100010011",
  42605=>"100100001",
  42606=>"000011010",
  42607=>"111111001",
  42608=>"101001101",
  42609=>"000000010",
  42610=>"000011111",
  42611=>"111110001",
  42612=>"011001010",
  42613=>"001101101",
  42614=>"100000000",
  42615=>"100011001",
  42616=>"111111001",
  42617=>"001010101",
  42618=>"111110001",
  42619=>"000101011",
  42620=>"100010010",
  42621=>"001101000",
  42622=>"000001011",
  42623=>"011100001",
  42624=>"111110111",
  42625=>"001011001",
  42626=>"111111111",
  42627=>"111001011",
  42628=>"100001010",
  42629=>"101100011",
  42630=>"000101111",
  42631=>"001110001",
  42632=>"001001011",
  42633=>"011100000",
  42634=>"001011111",
  42635=>"010100000",
  42636=>"000100000",
  42637=>"111110010",
  42638=>"010000010",
  42639=>"111110001",
  42640=>"010100101",
  42641=>"111101101",
  42642=>"101000101",
  42643=>"000010111",
  42644=>"111100010",
  42645=>"001100100",
  42646=>"000100010",
  42647=>"011001111",
  42648=>"010101011",
  42649=>"110110111",
  42650=>"100100011",
  42651=>"101111101",
  42652=>"111011011",
  42653=>"100110110",
  42654=>"010000101",
  42655=>"101010110",
  42656=>"001110000",
  42657=>"111110001",
  42658=>"001010111",
  42659=>"011001101",
  42660=>"100101011",
  42661=>"101001000",
  42662=>"000010111",
  42663=>"011010010",
  42664=>"000110001",
  42665=>"110011100",
  42666=>"010101101",
  42667=>"010010110",
  42668=>"110010000",
  42669=>"110001011",
  42670=>"000111101",
  42671=>"000000101",
  42672=>"111111011",
  42673=>"111100101",
  42674=>"111000100",
  42675=>"101101000",
  42676=>"000110101",
  42677=>"001011001",
  42678=>"010101111",
  42679=>"101101001",
  42680=>"111001101",
  42681=>"011011110",
  42682=>"011100000",
  42683=>"001110110",
  42684=>"011000010",
  42685=>"100101101",
  42686=>"010010100",
  42687=>"011001100",
  42688=>"111101000",
  42689=>"110111100",
  42690=>"001001001",
  42691=>"100101101",
  42692=>"100110010",
  42693=>"100001100",
  42694=>"011001001",
  42695=>"111100001",
  42696=>"000000011",
  42697=>"010011100",
  42698=>"100100101",
  42699=>"100101111",
  42700=>"000000110",
  42701=>"110100001",
  42702=>"110001101",
  42703=>"000001100",
  42704=>"101010111",
  42705=>"101011100",
  42706=>"010010101",
  42707=>"011010011",
  42708=>"111011000",
  42709=>"101100010",
  42710=>"000010011",
  42711=>"011101010",
  42712=>"101001101",
  42713=>"001000000",
  42714=>"001001000",
  42715=>"110110100",
  42716=>"010110100",
  42717=>"111100111",
  42718=>"010110111",
  42719=>"001111011",
  42720=>"001100001",
  42721=>"010000001",
  42722=>"000000010",
  42723=>"011110111",
  42724=>"011001001",
  42725=>"000000100",
  42726=>"000010001",
  42727=>"000111010",
  42728=>"001001001",
  42729=>"011101100",
  42730=>"011010001",
  42731=>"010101000",
  42732=>"000110000",
  42733=>"101110110",
  42734=>"111101111",
  42735=>"101001100",
  42736=>"011101100",
  42737=>"011011100",
  42738=>"011100001",
  42739=>"000011110",
  42740=>"100000010",
  42741=>"110111111",
  42742=>"010111110",
  42743=>"111010111",
  42744=>"011010010",
  42745=>"100110101",
  42746=>"101111111",
  42747=>"000100101",
  42748=>"011010101",
  42749=>"100110001",
  42750=>"001101100",
  42751=>"011110001",
  42752=>"111100101",
  42753=>"010010100",
  42754=>"100100100",
  42755=>"110101101",
  42756=>"111100101",
  42757=>"110010011",
  42758=>"101000001",
  42759=>"001111001",
  42760=>"011001000",
  42761=>"011111111",
  42762=>"001111100",
  42763=>"111000001",
  42764=>"110000001",
  42765=>"101110111",
  42766=>"000110000",
  42767=>"101000110",
  42768=>"110110001",
  42769=>"001001101",
  42770=>"111100111",
  42771=>"100011100",
  42772=>"111100011",
  42773=>"101110110",
  42774=>"111001110",
  42775=>"001101111",
  42776=>"101001101",
  42777=>"011010001",
  42778=>"011101001",
  42779=>"001100001",
  42780=>"110110111",
  42781=>"010100010",
  42782=>"001000100",
  42783=>"111110010",
  42784=>"010010000",
  42785=>"011110110",
  42786=>"011011000",
  42787=>"000111100",
  42788=>"101010000",
  42789=>"001100100",
  42790=>"111110000",
  42791=>"110010111",
  42792=>"110101101",
  42793=>"001000001",
  42794=>"011001100",
  42795=>"000000010",
  42796=>"011001111",
  42797=>"001000001",
  42798=>"010111100",
  42799=>"011110111",
  42800=>"001101100",
  42801=>"010010100",
  42802=>"000101000",
  42803=>"110101011",
  42804=>"010000111",
  42805=>"011011010",
  42806=>"000101001",
  42807=>"111111000",
  42808=>"000001001",
  42809=>"011010100",
  42810=>"000010101",
  42811=>"010110110",
  42812=>"100001100",
  42813=>"100011000",
  42814=>"011001111",
  42815=>"011000000",
  42816=>"101001010",
  42817=>"011000001",
  42818=>"111000001",
  42819=>"100101000",
  42820=>"011111110",
  42821=>"011111000",
  42822=>"000110000",
  42823=>"111110000",
  42824=>"100100000",
  42825=>"110111100",
  42826=>"011100000",
  42827=>"011101100",
  42828=>"100110111",
  42829=>"110011110",
  42830=>"111010101",
  42831=>"101010110",
  42832=>"100100100",
  42833=>"111010110",
  42834=>"011001110",
  42835=>"001010110",
  42836=>"000011001",
  42837=>"110101101",
  42838=>"000001110",
  42839=>"010111100",
  42840=>"100010111",
  42841=>"101010110",
  42842=>"010001001",
  42843=>"001000110",
  42844=>"001100111",
  42845=>"101000000",
  42846=>"100101000",
  42847=>"101100100",
  42848=>"110100011",
  42849=>"010110111",
  42850=>"001100011",
  42851=>"110000001",
  42852=>"110110100",
  42853=>"000100110",
  42854=>"100111000",
  42855=>"010110001",
  42856=>"110011011",
  42857=>"001101111",
  42858=>"111100001",
  42859=>"011001000",
  42860=>"000110010",
  42861=>"100010110",
  42862=>"010100100",
  42863=>"011110111",
  42864=>"010010010",
  42865=>"111111110",
  42866=>"001011111",
  42867=>"001011010",
  42868=>"101011000",
  42869=>"000111000",
  42870=>"010110000",
  42871=>"100101100",
  42872=>"000010000",
  42873=>"111011100",
  42874=>"110011000",
  42875=>"000010011",
  42876=>"100010010",
  42877=>"111001111",
  42878=>"010111000",
  42879=>"010010000",
  42880=>"100011100",
  42881=>"011000110",
  42882=>"111100001",
  42883=>"110111011",
  42884=>"101110010",
  42885=>"100110000",
  42886=>"001010011",
  42887=>"010011100",
  42888=>"011110111",
  42889=>"110000110",
  42890=>"000101110",
  42891=>"111111100",
  42892=>"001100000",
  42893=>"100000000",
  42894=>"100011011",
  42895=>"101000100",
  42896=>"001100100",
  42897=>"011000011",
  42898=>"111111000",
  42899=>"110001101",
  42900=>"101101110",
  42901=>"001001101",
  42902=>"111001100",
  42903=>"000000010",
  42904=>"000110101",
  42905=>"001010001",
  42906=>"101011011",
  42907=>"011101100",
  42908=>"010100011",
  42909=>"100001000",
  42910=>"101101000",
  42911=>"111100011",
  42912=>"101001111",
  42913=>"011111111",
  42914=>"011101001",
  42915=>"100011000",
  42916=>"101110000",
  42917=>"011100111",
  42918=>"001110010",
  42919=>"111011101",
  42920=>"111101010",
  42921=>"010101101",
  42922=>"001101000",
  42923=>"111000110",
  42924=>"010101110",
  42925=>"000011001",
  42926=>"001101000",
  42927=>"001101010",
  42928=>"010010000",
  42929=>"100011001",
  42930=>"000011000",
  42931=>"010011000",
  42932=>"101100010",
  42933=>"100101101",
  42934=>"010111101",
  42935=>"000000001",
  42936=>"000000111",
  42937=>"001010000",
  42938=>"000101101",
  42939=>"110011111",
  42940=>"110001001",
  42941=>"010111111",
  42942=>"011000000",
  42943=>"110001111",
  42944=>"100011001",
  42945=>"000100100",
  42946=>"111100101",
  42947=>"111101111",
  42948=>"100100011",
  42949=>"010101101",
  42950=>"100111101",
  42951=>"100100111",
  42952=>"101000000",
  42953=>"010101110",
  42954=>"011011100",
  42955=>"000110110",
  42956=>"101000001",
  42957=>"110110010",
  42958=>"101111100",
  42959=>"100010111",
  42960=>"101010110",
  42961=>"111000111",
  42962=>"000100101",
  42963=>"001011101",
  42964=>"011010100",
  42965=>"100101100",
  42966=>"111101001",
  42967=>"111101000",
  42968=>"100000011",
  42969=>"001101010",
  42970=>"000110101",
  42971=>"010100111",
  42972=>"100001100",
  42973=>"101111010",
  42974=>"101010000",
  42975=>"101011010",
  42976=>"010111000",
  42977=>"111000111",
  42978=>"100011010",
  42979=>"011000101",
  42980=>"100001100",
  42981=>"101101001",
  42982=>"110010000",
  42983=>"111011011",
  42984=>"000000000",
  42985=>"001110011",
  42986=>"101111000",
  42987=>"111110110",
  42988=>"111011001",
  42989=>"111000010",
  42990=>"010011000",
  42991=>"000100101",
  42992=>"110001000",
  42993=>"101110110",
  42994=>"010111111",
  42995=>"000011101",
  42996=>"110101010",
  42997=>"001111011",
  42998=>"100111111",
  42999=>"100001101",
  43000=>"111000011",
  43001=>"110011100",
  43002=>"000111101",
  43003=>"000100000",
  43004=>"001011000",
  43005=>"010110011",
  43006=>"011010110",
  43007=>"110100100",
  43008=>"010101111",
  43009=>"001100101",
  43010=>"110000000",
  43011=>"100100010",
  43012=>"110110011",
  43013=>"010111010",
  43014=>"110101000",
  43015=>"011011110",
  43016=>"010101000",
  43017=>"110100011",
  43018=>"110100111",
  43019=>"011011111",
  43020=>"010010101",
  43021=>"000110111",
  43022=>"000100111",
  43023=>"111011011",
  43024=>"110010100",
  43025=>"011100010",
  43026=>"011011110",
  43027=>"100101110",
  43028=>"000000010",
  43029=>"010101100",
  43030=>"111110011",
  43031=>"000010111",
  43032=>"001100001",
  43033=>"111111000",
  43034=>"111010101",
  43035=>"111101000",
  43036=>"101000001",
  43037=>"010111000",
  43038=>"010010011",
  43039=>"011100010",
  43040=>"111000111",
  43041=>"101001111",
  43042=>"111100011",
  43043=>"100010100",
  43044=>"110011111",
  43045=>"100100110",
  43046=>"000100010",
  43047=>"000010110",
  43048=>"111110000",
  43049=>"100101000",
  43050=>"101010101",
  43051=>"001100111",
  43052=>"110000110",
  43053=>"001010011",
  43054=>"000011100",
  43055=>"111111111",
  43056=>"000110000",
  43057=>"001000100",
  43058=>"110011010",
  43059=>"011010001",
  43060=>"111101110",
  43061=>"000000001",
  43062=>"000111111",
  43063=>"101110011",
  43064=>"010101000",
  43065=>"010101010",
  43066=>"001000110",
  43067=>"101001011",
  43068=>"110011100",
  43069=>"011110010",
  43070=>"000010110",
  43071=>"011101100",
  43072=>"101100111",
  43073=>"100110100",
  43074=>"011010011",
  43075=>"000000111",
  43076=>"111001001",
  43077=>"111001110",
  43078=>"011110000",
  43079=>"110111000",
  43080=>"111110111",
  43081=>"110011111",
  43082=>"001011101",
  43083=>"001100011",
  43084=>"001100100",
  43085=>"100000011",
  43086=>"000110001",
  43087=>"111101000",
  43088=>"111111110",
  43089=>"111110100",
  43090=>"001110010",
  43091=>"000000110",
  43092=>"101101111",
  43093=>"001010110",
  43094=>"001100000",
  43095=>"011000100",
  43096=>"010111111",
  43097=>"001011101",
  43098=>"010110001",
  43099=>"011111110",
  43100=>"011010111",
  43101=>"110000100",
  43102=>"111001001",
  43103=>"001010101",
  43104=>"010000010",
  43105=>"101001110",
  43106=>"101101101",
  43107=>"110110010",
  43108=>"000100100",
  43109=>"100100010",
  43110=>"100110001",
  43111=>"111110110",
  43112=>"001010100",
  43113=>"111011001",
  43114=>"111000010",
  43115=>"011000010",
  43116=>"010000010",
  43117=>"000000000",
  43118=>"000000010",
  43119=>"010010101",
  43120=>"111001011",
  43121=>"010111101",
  43122=>"111010100",
  43123=>"111011100",
  43124=>"100101101",
  43125=>"111010100",
  43126=>"110010110",
  43127=>"110000011",
  43128=>"010001011",
  43129=>"000101100",
  43130=>"111110001",
  43131=>"010101100",
  43132=>"101011000",
  43133=>"010000001",
  43134=>"010101101",
  43135=>"111101111",
  43136=>"000110101",
  43137=>"111110111",
  43138=>"001001000",
  43139=>"111000101",
  43140=>"100001111",
  43141=>"011000000",
  43142=>"111100110",
  43143=>"011111111",
  43144=>"111000100",
  43145=>"101001100",
  43146=>"110010111",
  43147=>"111100111",
  43148=>"101100000",
  43149=>"000100100",
  43150=>"010110000",
  43151=>"000001000",
  43152=>"010001110",
  43153=>"100110001",
  43154=>"110001010",
  43155=>"010000000",
  43156=>"111111000",
  43157=>"011101111",
  43158=>"101101010",
  43159=>"101000100",
  43160=>"000111000",
  43161=>"001010010",
  43162=>"111100000",
  43163=>"110101000",
  43164=>"011111010",
  43165=>"011110111",
  43166=>"100110010",
  43167=>"100100111",
  43168=>"011111101",
  43169=>"011011001",
  43170=>"111101001",
  43171=>"111000011",
  43172=>"000101011",
  43173=>"111000001",
  43174=>"100010000",
  43175=>"001000000",
  43176=>"011111101",
  43177=>"000110010",
  43178=>"010000001",
  43179=>"010110100",
  43180=>"010010110",
  43181=>"011010100",
  43182=>"001000001",
  43183=>"111100110",
  43184=>"101100110",
  43185=>"000011111",
  43186=>"010000000",
  43187=>"010110011",
  43188=>"110010010",
  43189=>"111111010",
  43190=>"010100001",
  43191=>"110110111",
  43192=>"001100010",
  43193=>"110100101",
  43194=>"100010101",
  43195=>"011000110",
  43196=>"000010110",
  43197=>"100101100",
  43198=>"101100101",
  43199=>"110010001",
  43200=>"011110000",
  43201=>"100010110",
  43202=>"100101001",
  43203=>"001001101",
  43204=>"101111011",
  43205=>"101001100",
  43206=>"001111110",
  43207=>"000010110",
  43208=>"110101001",
  43209=>"001101110",
  43210=>"111111000",
  43211=>"110011010",
  43212=>"011101111",
  43213=>"011000110",
  43214=>"000100100",
  43215=>"111111110",
  43216=>"001110110",
  43217=>"010001001",
  43218=>"001100100",
  43219=>"011010011",
  43220=>"101101010",
  43221=>"011100110",
  43222=>"000011010",
  43223=>"110000101",
  43224=>"111111000",
  43225=>"011001110",
  43226=>"010001010",
  43227=>"000010101",
  43228=>"001001011",
  43229=>"100100101",
  43230=>"101010111",
  43231=>"110011001",
  43232=>"011100000",
  43233=>"110100000",
  43234=>"000011101",
  43235=>"100111110",
  43236=>"111110110",
  43237=>"001101010",
  43238=>"011101011",
  43239=>"011101011",
  43240=>"110100001",
  43241=>"100001101",
  43242=>"100011100",
  43243=>"011000011",
  43244=>"101001100",
  43245=>"000111011",
  43246=>"011000111",
  43247=>"000001000",
  43248=>"101101001",
  43249=>"001101100",
  43250=>"011100000",
  43251=>"010000111",
  43252=>"101111010",
  43253=>"101100110",
  43254=>"001100101",
  43255=>"000101110",
  43256=>"111110010",
  43257=>"100000101",
  43258=>"011110010",
  43259=>"100001011",
  43260=>"000111111",
  43261=>"100001001",
  43262=>"000111100",
  43263=>"111010001",
  43264=>"100101101",
  43265=>"100000110",
  43266=>"100111111",
  43267=>"111110100",
  43268=>"000011000",
  43269=>"000101111",
  43270=>"111011011",
  43271=>"001010110",
  43272=>"011101111",
  43273=>"111100111",
  43274=>"010001010",
  43275=>"111111001",
  43276=>"100110010",
  43277=>"100000011",
  43278=>"010010100",
  43279=>"001101100",
  43280=>"000000101",
  43281=>"110010011",
  43282=>"100010111",
  43283=>"111110010",
  43284=>"000000001",
  43285=>"110111111",
  43286=>"000110110",
  43287=>"010101101",
  43288=>"110110100",
  43289=>"100001100",
  43290=>"101010000",
  43291=>"101111101",
  43292=>"000110001",
  43293=>"001110101",
  43294=>"100000111",
  43295=>"010010110",
  43296=>"010010110",
  43297=>"100001111",
  43298=>"011001101",
  43299=>"111110001",
  43300=>"011111100",
  43301=>"110111000",
  43302=>"110101011",
  43303=>"001001101",
  43304=>"010010001",
  43305=>"101101011",
  43306=>"101001010",
  43307=>"110100101",
  43308=>"101000000",
  43309=>"100111011",
  43310=>"111111101",
  43311=>"010000110",
  43312=>"110011101",
  43313=>"000011110",
  43314=>"110100100",
  43315=>"010110001",
  43316=>"011110111",
  43317=>"111101011",
  43318=>"011101011",
  43319=>"001000000",
  43320=>"001000100",
  43321=>"101010011",
  43322=>"000111100",
  43323=>"000000110",
  43324=>"011101011",
  43325=>"101000100",
  43326=>"010001000",
  43327=>"000000101",
  43328=>"110000011",
  43329=>"001111001",
  43330=>"111010001",
  43331=>"110011100",
  43332=>"011100110",
  43333=>"000001110",
  43334=>"001110101",
  43335=>"001100100",
  43336=>"111001001",
  43337=>"100011000",
  43338=>"111101111",
  43339=>"110010110",
  43340=>"101001101",
  43341=>"011100010",
  43342=>"100101100",
  43343=>"101111111",
  43344=>"110101111",
  43345=>"111001011",
  43346=>"010100001",
  43347=>"100010110",
  43348=>"001001110",
  43349=>"100101111",
  43350=>"101000110",
  43351=>"100001110",
  43352=>"010110111",
  43353=>"000100111",
  43354=>"001101100",
  43355=>"000001100",
  43356=>"111100001",
  43357=>"111101000",
  43358=>"001100101",
  43359=>"100100110",
  43360=>"010000110",
  43361=>"101110001",
  43362=>"001011011",
  43363=>"010010100",
  43364=>"000111100",
  43365=>"110001000",
  43366=>"110001110",
  43367=>"010110000",
  43368=>"100000010",
  43369=>"001111111",
  43370=>"010101111",
  43371=>"110110111",
  43372=>"100110100",
  43373=>"010111111",
  43374=>"001001000",
  43375=>"111101101",
  43376=>"000010001",
  43377=>"011010100",
  43378=>"111010000",
  43379=>"111110100",
  43380=>"000000010",
  43381=>"010100011",
  43382=>"101010110",
  43383=>"011010100",
  43384=>"001001100",
  43385=>"010101110",
  43386=>"010101111",
  43387=>"000000010",
  43388=>"011010011",
  43389=>"100011011",
  43390=>"111011000",
  43391=>"100001111",
  43392=>"000001010",
  43393=>"000010011",
  43394=>"101100001",
  43395=>"101100001",
  43396=>"111101101",
  43397=>"101101100",
  43398=>"000100101",
  43399=>"000101011",
  43400=>"010110111",
  43401=>"100100101",
  43402=>"100001111",
  43403=>"101110101",
  43404=>"000110111",
  43405=>"000010000",
  43406=>"100100011",
  43407=>"100110101",
  43408=>"000001010",
  43409=>"011110111",
  43410=>"100011001",
  43411=>"111001101",
  43412=>"001011101",
  43413=>"010100101",
  43414=>"100011000",
  43415=>"110111101",
  43416=>"010111011",
  43417=>"111001111",
  43418=>"010011111",
  43419=>"101011001",
  43420=>"010111011",
  43421=>"011101010",
  43422=>"101110011",
  43423=>"010110100",
  43424=>"010011110",
  43425=>"011110001",
  43426=>"111101111",
  43427=>"010101101",
  43428=>"101110110",
  43429=>"000110100",
  43430=>"010001001",
  43431=>"010110000",
  43432=>"111111001",
  43433=>"001111111",
  43434=>"100001010",
  43435=>"000010111",
  43436=>"110100100",
  43437=>"001011000",
  43438=>"000100110",
  43439=>"001011110",
  43440=>"100011001",
  43441=>"000011011",
  43442=>"101101111",
  43443=>"010010010",
  43444=>"010011100",
  43445=>"101111011",
  43446=>"000101000",
  43447=>"100110100",
  43448=>"110111000",
  43449=>"000111110",
  43450=>"110000000",
  43451=>"100011000",
  43452=>"110111111",
  43453=>"000000011",
  43454=>"101100100",
  43455=>"111101000",
  43456=>"011110010",
  43457=>"001110110",
  43458=>"011001110",
  43459=>"001001000",
  43460=>"001110111",
  43461=>"101100111",
  43462=>"101001111",
  43463=>"010010011",
  43464=>"000010101",
  43465=>"011101110",
  43466=>"101000010",
  43467=>"111000111",
  43468=>"101000000",
  43469=>"010001110",
  43470=>"011000111",
  43471=>"110011000",
  43472=>"001101011",
  43473=>"111001111",
  43474=>"101000100",
  43475=>"110001110",
  43476=>"001101001",
  43477=>"101010000",
  43478=>"100110010",
  43479=>"100011011",
  43480=>"101110001",
  43481=>"010010001",
  43482=>"111110111",
  43483=>"011011000",
  43484=>"011100100",
  43485=>"011110011",
  43486=>"101111010",
  43487=>"011111011",
  43488=>"110111011",
  43489=>"001110111",
  43490=>"001101110",
  43491=>"101011010",
  43492=>"001011101",
  43493=>"011101010",
  43494=>"001111001",
  43495=>"111011101",
  43496=>"111111111",
  43497=>"110111111",
  43498=>"111110010",
  43499=>"111111011",
  43500=>"100010110",
  43501=>"101101111",
  43502=>"110111000",
  43503=>"001010100",
  43504=>"101110000",
  43505=>"011110100",
  43506=>"000110100",
  43507=>"001011101",
  43508=>"011011001",
  43509=>"101110011",
  43510=>"110110110",
  43511=>"010111110",
  43512=>"011001100",
  43513=>"011100000",
  43514=>"111111111",
  43515=>"100010101",
  43516=>"100001000",
  43517=>"111101111",
  43518=>"010101001",
  43519=>"010000000",
  43520=>"110101001",
  43521=>"011100101",
  43522=>"000011000",
  43523=>"011000101",
  43524=>"001001101",
  43525=>"011110001",
  43526=>"110111100",
  43527=>"111101010",
  43528=>"100110110",
  43529=>"100101100",
  43530=>"111000001",
  43531=>"111101100",
  43532=>"011010000",
  43533=>"100000001",
  43534=>"101110000",
  43535=>"000100001",
  43536=>"111111011",
  43537=>"000001100",
  43538=>"110111110",
  43539=>"001011110",
  43540=>"010000101",
  43541=>"001100000",
  43542=>"101001011",
  43543=>"100110101",
  43544=>"011001101",
  43545=>"111101000",
  43546=>"111000100",
  43547=>"001001001",
  43548=>"001100011",
  43549=>"110010100",
  43550=>"001101000",
  43551=>"111111100",
  43552=>"011011110",
  43553=>"011100010",
  43554=>"001001110",
  43555=>"101111100",
  43556=>"011110011",
  43557=>"110000000",
  43558=>"100011010",
  43559=>"000100110",
  43560=>"101011101",
  43561=>"100000110",
  43562=>"000101001",
  43563=>"001111011",
  43564=>"001000010",
  43565=>"001110110",
  43566=>"011000100",
  43567=>"111000100",
  43568=>"010111000",
  43569=>"101011111",
  43570=>"011001001",
  43571=>"001011000",
  43572=>"111000111",
  43573=>"011010001",
  43574=>"111110101",
  43575=>"100001111",
  43576=>"100101011",
  43577=>"001100110",
  43578=>"000001000",
  43579=>"000100110",
  43580=>"101110101",
  43581=>"000001111",
  43582=>"001001100",
  43583=>"001011010",
  43584=>"001100001",
  43585=>"111011010",
  43586=>"010011111",
  43587=>"100010010",
  43588=>"111010110",
  43589=>"101000101",
  43590=>"000000000",
  43591=>"110000100",
  43592=>"101100000",
  43593=>"100001101",
  43594=>"000000000",
  43595=>"001110011",
  43596=>"110101111",
  43597=>"001100000",
  43598=>"001111111",
  43599=>"101111110",
  43600=>"011111010",
  43601=>"010000100",
  43602=>"011111000",
  43603=>"001001110",
  43604=>"011111100",
  43605=>"000101000",
  43606=>"001110010",
  43607=>"011000001",
  43608=>"011000001",
  43609=>"011111100",
  43610=>"110010101",
  43611=>"000001001",
  43612=>"000011010",
  43613=>"001000000",
  43614=>"001010111",
  43615=>"111111010",
  43616=>"110010001",
  43617=>"001011101",
  43618=>"010000100",
  43619=>"011110111",
  43620=>"010101111",
  43621=>"101001101",
  43622=>"000111010",
  43623=>"110110100",
  43624=>"100011000",
  43625=>"011100000",
  43626=>"101010101",
  43627=>"100011111",
  43628=>"101010101",
  43629=>"110100110",
  43630=>"000010100",
  43631=>"011100001",
  43632=>"100100110",
  43633=>"000001011",
  43634=>"101000001",
  43635=>"000011111",
  43636=>"000000010",
  43637=>"001000100",
  43638=>"011111000",
  43639=>"111001101",
  43640=>"011101101",
  43641=>"111001111",
  43642=>"110101010",
  43643=>"100110101",
  43644=>"011001111",
  43645=>"101010101",
  43646=>"010110010",
  43647=>"000110101",
  43648=>"010001000",
  43649=>"111101000",
  43650=>"100011111",
  43651=>"001001000",
  43652=>"000110111",
  43653=>"001001000",
  43654=>"010101101",
  43655=>"000000000",
  43656=>"000110101",
  43657=>"101111111",
  43658=>"011110011",
  43659=>"101010010",
  43660=>"000001101",
  43661=>"000011000",
  43662=>"110011111",
  43663=>"010001001",
  43664=>"011100110",
  43665=>"101111110",
  43666=>"110011100",
  43667=>"010010111",
  43668=>"000010000",
  43669=>"110001001",
  43670=>"001000000",
  43671=>"101011101",
  43672=>"001001010",
  43673=>"011011000",
  43674=>"101100000",
  43675=>"101010110",
  43676=>"011111101",
  43677=>"110000100",
  43678=>"001000101",
  43679=>"100010010",
  43680=>"110000001",
  43681=>"000110110",
  43682=>"011111001",
  43683=>"011010100",
  43684=>"000110010",
  43685=>"010110000",
  43686=>"011111010",
  43687=>"110011110",
  43688=>"110001000",
  43689=>"000001100",
  43690=>"011100100",
  43691=>"111001010",
  43692=>"011111000",
  43693=>"010100001",
  43694=>"000101100",
  43695=>"111101111",
  43696=>"000001100",
  43697=>"011001110",
  43698=>"001101010",
  43699=>"110101110",
  43700=>"000111011",
  43701=>"101010010",
  43702=>"111111000",
  43703=>"111100001",
  43704=>"110111011",
  43705=>"011111111",
  43706=>"011101010",
  43707=>"010111000",
  43708=>"100001010",
  43709=>"101010000",
  43710=>"000010101",
  43711=>"011111110",
  43712=>"110010000",
  43713=>"000110111",
  43714=>"100110011",
  43715=>"000001000",
  43716=>"100011110",
  43717=>"000000100",
  43718=>"101010111",
  43719=>"010101011",
  43720=>"000001011",
  43721=>"110101110",
  43722=>"100001000",
  43723=>"001100010",
  43724=>"101000101",
  43725=>"010100101",
  43726=>"011010010",
  43727=>"110111101",
  43728=>"111111101",
  43729=>"000111111",
  43730=>"101110110",
  43731=>"100010000",
  43732=>"101101101",
  43733=>"010010000",
  43734=>"101011100",
  43735=>"111001010",
  43736=>"000011101",
  43737=>"111001010",
  43738=>"111110010",
  43739=>"000000100",
  43740=>"010011010",
  43741=>"110001001",
  43742=>"000101011",
  43743=>"110101111",
  43744=>"010010000",
  43745=>"000111011",
  43746=>"001110101",
  43747=>"111011111",
  43748=>"000001101",
  43749=>"010011010",
  43750=>"000000000",
  43751=>"011111001",
  43752=>"110011001",
  43753=>"000010000",
  43754=>"111111011",
  43755=>"100100010",
  43756=>"010110101",
  43757=>"010100100",
  43758=>"000101110",
  43759=>"110111100",
  43760=>"011010011",
  43761=>"110010011",
  43762=>"011000010",
  43763=>"011000100",
  43764=>"001000010",
  43765=>"110000000",
  43766=>"101111100",
  43767=>"100101110",
  43768=>"001001111",
  43769=>"010100001",
  43770=>"110011110",
  43771=>"111110000",
  43772=>"011111010",
  43773=>"010000110",
  43774=>"010001011",
  43775=>"001001000",
  43776=>"000011001",
  43777=>"000111001",
  43778=>"101111011",
  43779=>"101000011",
  43780=>"110111011",
  43781=>"100001100",
  43782=>"000100101",
  43783=>"111101110",
  43784=>"101010001",
  43785=>"011011011",
  43786=>"110011111",
  43787=>"101011001",
  43788=>"001110110",
  43789=>"001110101",
  43790=>"100111101",
  43791=>"001000101",
  43792=>"011100010",
  43793=>"110110001",
  43794=>"110110111",
  43795=>"111101110",
  43796=>"100111111",
  43797=>"011011010",
  43798=>"101011011",
  43799=>"100110000",
  43800=>"101001011",
  43801=>"101001010",
  43802=>"000000101",
  43803=>"100001010",
  43804=>"100100000",
  43805=>"000101111",
  43806=>"101110000",
  43807=>"101010011",
  43808=>"001100110",
  43809=>"111011111",
  43810=>"001101001",
  43811=>"111000000",
  43812=>"010000011",
  43813=>"110111001",
  43814=>"001011100",
  43815=>"100011100",
  43816=>"011000001",
  43817=>"001000000",
  43818=>"011001000",
  43819=>"101111111",
  43820=>"001100111",
  43821=>"000000000",
  43822=>"101011110",
  43823=>"000101100",
  43824=>"001001110",
  43825=>"111000001",
  43826=>"000001100",
  43827=>"001001000",
  43828=>"010110010",
  43829=>"111111010",
  43830=>"111001110",
  43831=>"101100111",
  43832=>"101011011",
  43833=>"010011110",
  43834=>"111111100",
  43835=>"101100011",
  43836=>"001100101",
  43837=>"100010110",
  43838=>"000001011",
  43839=>"011011101",
  43840=>"100100000",
  43841=>"000011001",
  43842=>"011010100",
  43843=>"101111100",
  43844=>"011010100",
  43845=>"110111000",
  43846=>"011111001",
  43847=>"100001111",
  43848=>"011010110",
  43849=>"000000000",
  43850=>"001111110",
  43851=>"101000100",
  43852=>"100111000",
  43853=>"100000001",
  43854=>"000000101",
  43855=>"000111011",
  43856=>"101101111",
  43857=>"100110110",
  43858=>"011100011",
  43859=>"100011001",
  43860=>"110101100",
  43861=>"000001000",
  43862=>"001001011",
  43863=>"100110111",
  43864=>"111010100",
  43865=>"001011000",
  43866=>"001100011",
  43867=>"111010011",
  43868=>"010100010",
  43869=>"111011010",
  43870=>"001111000",
  43871=>"101101110",
  43872=>"001100100",
  43873=>"110111111",
  43874=>"010111100",
  43875=>"100111000",
  43876=>"111001000",
  43877=>"111000010",
  43878=>"101011110",
  43879=>"000111011",
  43880=>"000001101",
  43881=>"001000100",
  43882=>"001001111",
  43883=>"001000010",
  43884=>"011000111",
  43885=>"000011001",
  43886=>"001101110",
  43887=>"101001100",
  43888=>"101100101",
  43889=>"000000101",
  43890=>"010110110",
  43891=>"001001101",
  43892=>"000101000",
  43893=>"000000100",
  43894=>"000111111",
  43895=>"010010111",
  43896=>"011001111",
  43897=>"010011000",
  43898=>"101111110",
  43899=>"100100010",
  43900=>"110101011",
  43901=>"101001011",
  43902=>"101011010",
  43903=>"101100010",
  43904=>"001000111",
  43905=>"010001101",
  43906=>"000100101",
  43907=>"111001001",
  43908=>"010101000",
  43909=>"101010100",
  43910=>"010111111",
  43911=>"100000000",
  43912=>"100000110",
  43913=>"111011111",
  43914=>"011010001",
  43915=>"111111111",
  43916=>"111001101",
  43917=>"011101100",
  43918=>"000111011",
  43919=>"001000100",
  43920=>"101011011",
  43921=>"100000100",
  43922=>"000010001",
  43923=>"000101100",
  43924=>"011000001",
  43925=>"100001000",
  43926=>"100111001",
  43927=>"110001100",
  43928=>"010100110",
  43929=>"111111110",
  43930=>"111010110",
  43931=>"001100101",
  43932=>"001110000",
  43933=>"100110001",
  43934=>"111101111",
  43935=>"111100011",
  43936=>"000010111",
  43937=>"011100000",
  43938=>"010100100",
  43939=>"100100110",
  43940=>"001011000",
  43941=>"110111000",
  43942=>"110010111",
  43943=>"110001000",
  43944=>"101101110",
  43945=>"100100000",
  43946=>"101100001",
  43947=>"000000010",
  43948=>"110010100",
  43949=>"011110010",
  43950=>"110000010",
  43951=>"000000001",
  43952=>"110001000",
  43953=>"010000110",
  43954=>"011110100",
  43955=>"010000111",
  43956=>"011100100",
  43957=>"000101111",
  43958=>"111111110",
  43959=>"001100001",
  43960=>"101100010",
  43961=>"101011111",
  43962=>"110111000",
  43963=>"000110111",
  43964=>"111101111",
  43965=>"000101111",
  43966=>"010101000",
  43967=>"000011111",
  43968=>"100011000",
  43969=>"101111011",
  43970=>"000000000",
  43971=>"001110111",
  43972=>"111000101",
  43973=>"001010010",
  43974=>"101101100",
  43975=>"100011000",
  43976=>"001011011",
  43977=>"001001100",
  43978=>"010100111",
  43979=>"100000111",
  43980=>"111011111",
  43981=>"011011110",
  43982=>"110100101",
  43983=>"000111011",
  43984=>"110100100",
  43985=>"011010000",
  43986=>"101000101",
  43987=>"001101101",
  43988=>"111110001",
  43989=>"111001000",
  43990=>"000100001",
  43991=>"111000100",
  43992=>"111100000",
  43993=>"111011111",
  43994=>"101000001",
  43995=>"011010101",
  43996=>"111100101",
  43997=>"110011111",
  43998=>"001010111",
  43999=>"110111110",
  44000=>"011100101",
  44001=>"001101000",
  44002=>"111110010",
  44003=>"111111100",
  44004=>"111111011",
  44005=>"001100100",
  44006=>"000111111",
  44007=>"001000111",
  44008=>"110000101",
  44009=>"011101111",
  44010=>"101101111",
  44011=>"100000100",
  44012=>"000011100",
  44013=>"111000111",
  44014=>"000001010",
  44015=>"001000110",
  44016=>"100110000",
  44017=>"110001000",
  44018=>"011001010",
  44019=>"000011111",
  44020=>"001101101",
  44021=>"110111100",
  44022=>"001000110",
  44023=>"000001001",
  44024=>"110111101",
  44025=>"011111100",
  44026=>"100011011",
  44027=>"111111100",
  44028=>"010000100",
  44029=>"110111110",
  44030=>"000001111",
  44031=>"011111010",
  44032=>"010000101",
  44033=>"111100100",
  44034=>"000000101",
  44035=>"111111001",
  44036=>"011001011",
  44037=>"000110101",
  44038=>"000010110",
  44039=>"011101101",
  44040=>"001001001",
  44041=>"101101101",
  44042=>"010000110",
  44043=>"110011100",
  44044=>"110100110",
  44045=>"001011100",
  44046=>"101110010",
  44047=>"100100000",
  44048=>"011100001",
  44049=>"000110011",
  44050=>"011110011",
  44051=>"010101110",
  44052=>"001000001",
  44053=>"111100000",
  44054=>"101101101",
  44055=>"101110100",
  44056=>"111110001",
  44057=>"101101110",
  44058=>"001100101",
  44059=>"110110011",
  44060=>"011110100",
  44061=>"011100100",
  44062=>"010011110",
  44063=>"110101001",
  44064=>"111001000",
  44065=>"110010111",
  44066=>"011101100",
  44067=>"111010001",
  44068=>"001001101",
  44069=>"111000011",
  44070=>"101101000",
  44071=>"101111111",
  44072=>"101111101",
  44073=>"101100100",
  44074=>"010101010",
  44075=>"101110010",
  44076=>"000111010",
  44077=>"000111011",
  44078=>"110100110",
  44079=>"111101011",
  44080=>"111001110",
  44081=>"111110100",
  44082=>"001111010",
  44083=>"011110011",
  44084=>"000000100",
  44085=>"100001100",
  44086=>"100101000",
  44087=>"111111001",
  44088=>"101101010",
  44089=>"100011011",
  44090=>"000111101",
  44091=>"000100101",
  44092=>"110110010",
  44093=>"000100101",
  44094=>"100111101",
  44095=>"101101110",
  44096=>"010101110",
  44097=>"101101000",
  44098=>"011010100",
  44099=>"001011101",
  44100=>"101101111",
  44101=>"100100110",
  44102=>"100101110",
  44103=>"000001001",
  44104=>"111001110",
  44105=>"111001010",
  44106=>"001100000",
  44107=>"111001111",
  44108=>"101100000",
  44109=>"011000011",
  44110=>"001111000",
  44111=>"101100111",
  44112=>"101000011",
  44113=>"000111111",
  44114=>"001110110",
  44115=>"100010111",
  44116=>"010110010",
  44117=>"111011000",
  44118=>"010010110",
  44119=>"101101111",
  44120=>"000011110",
  44121=>"101001110",
  44122=>"100100111",
  44123=>"010010010",
  44124=>"010010011",
  44125=>"110001001",
  44126=>"010001111",
  44127=>"011001000",
  44128=>"000001101",
  44129=>"001111010",
  44130=>"001101001",
  44131=>"000001011",
  44132=>"101101100",
  44133=>"001101000",
  44134=>"111100100",
  44135=>"011101000",
  44136=>"010001010",
  44137=>"001001011",
  44138=>"010011001",
  44139=>"000000111",
  44140=>"101100110",
  44141=>"010011100",
  44142=>"101000111",
  44143=>"001000100",
  44144=>"110001001",
  44145=>"010001000",
  44146=>"100011011",
  44147=>"001101110",
  44148=>"100001111",
  44149=>"001111100",
  44150=>"001110101",
  44151=>"000111000",
  44152=>"111101011",
  44153=>"101100111",
  44154=>"010000100",
  44155=>"101101101",
  44156=>"001001101",
  44157=>"101101101",
  44158=>"000100011",
  44159=>"000000101",
  44160=>"011011100",
  44161=>"101010000",
  44162=>"010111101",
  44163=>"001101100",
  44164=>"100110111",
  44165=>"100110011",
  44166=>"100001001",
  44167=>"110110101",
  44168=>"111100000",
  44169=>"000010011",
  44170=>"100110101",
  44171=>"010111101",
  44172=>"110100101",
  44173=>"011001001",
  44174=>"100000001",
  44175=>"111101101",
  44176=>"010111100",
  44177=>"101011101",
  44178=>"100101000",
  44179=>"001111001",
  44180=>"001100011",
  44181=>"100110010",
  44182=>"010011010",
  44183=>"101000010",
  44184=>"101001001",
  44185=>"100100010",
  44186=>"000000010",
  44187=>"001001111",
  44188=>"101101111",
  44189=>"111000010",
  44190=>"001001110",
  44191=>"001111001",
  44192=>"011010100",
  44193=>"001111011",
  44194=>"100000100",
  44195=>"000010100",
  44196=>"110000110",
  44197=>"001001100",
  44198=>"110101000",
  44199=>"011111110",
  44200=>"010001011",
  44201=>"101010010",
  44202=>"010110001",
  44203=>"001100011",
  44204=>"110010110",
  44205=>"001001100",
  44206=>"100110000",
  44207=>"010000011",
  44208=>"011011000",
  44209=>"101000110",
  44210=>"101010111",
  44211=>"101111011",
  44212=>"001100000",
  44213=>"010010001",
  44214=>"000000010",
  44215=>"100000000",
  44216=>"001111111",
  44217=>"011100111",
  44218=>"010011000",
  44219=>"100111101",
  44220=>"100001000",
  44221=>"011111001",
  44222=>"001011110",
  44223=>"001110110",
  44224=>"111001101",
  44225=>"101011100",
  44226=>"010111110",
  44227=>"111101101",
  44228=>"001110101",
  44229=>"111011111",
  44230=>"001110111",
  44231=>"000100111",
  44232=>"001000000",
  44233=>"111101111",
  44234=>"010111110",
  44235=>"111110110",
  44236=>"111111000",
  44237=>"000101110",
  44238=>"010001000",
  44239=>"010101000",
  44240=>"011011010",
  44241=>"100011000",
  44242=>"110010001",
  44243=>"100001101",
  44244=>"110001001",
  44245=>"010000111",
  44246=>"011011011",
  44247=>"011111010",
  44248=>"011110001",
  44249=>"100001101",
  44250=>"000111001",
  44251=>"100000100",
  44252=>"010000010",
  44253=>"011100111",
  44254=>"111110101",
  44255=>"010001110",
  44256=>"001110001",
  44257=>"000000010",
  44258=>"110010111",
  44259=>"000110110",
  44260=>"101100101",
  44261=>"011000010",
  44262=>"000101010",
  44263=>"000100011",
  44264=>"001100010",
  44265=>"001001100",
  44266=>"001110111",
  44267=>"010000000",
  44268=>"011010100",
  44269=>"010101100",
  44270=>"110010000",
  44271=>"111110101",
  44272=>"010100011",
  44273=>"001001000",
  44274=>"111001111",
  44275=>"011011100",
  44276=>"110011110",
  44277=>"001101101",
  44278=>"111110101",
  44279=>"010011010",
  44280=>"110001111",
  44281=>"111001000",
  44282=>"011010001",
  44283=>"010010010",
  44284=>"100000001",
  44285=>"111001001",
  44286=>"001100011",
  44287=>"111110000",
  44288=>"100100111",
  44289=>"010110100",
  44290=>"111110011",
  44291=>"001110111",
  44292=>"010000011",
  44293=>"001100001",
  44294=>"011011101",
  44295=>"000101110",
  44296=>"101010001",
  44297=>"100110011",
  44298=>"111110110",
  44299=>"100000000",
  44300=>"001110111",
  44301=>"101101100",
  44302=>"101011010",
  44303=>"110011111",
  44304=>"101001101",
  44305=>"010010101",
  44306=>"101111100",
  44307=>"110101010",
  44308=>"111110100",
  44309=>"100111111",
  44310=>"000110100",
  44311=>"110110011",
  44312=>"001001101",
  44313=>"011001001",
  44314=>"000110011",
  44315=>"011101111",
  44316=>"101111010",
  44317=>"110100000",
  44318=>"100001101",
  44319=>"001110101",
  44320=>"100100011",
  44321=>"100001000",
  44322=>"010001110",
  44323=>"111111011",
  44324=>"011011100",
  44325=>"100110010",
  44326=>"011010100",
  44327=>"111111010",
  44328=>"110100000",
  44329=>"100001101",
  44330=>"000011101",
  44331=>"001010011",
  44332=>"101101100",
  44333=>"100100000",
  44334=>"000100001",
  44335=>"110101001",
  44336=>"001001110",
  44337=>"000101011",
  44338=>"100000111",
  44339=>"001100010",
  44340=>"000010101",
  44341=>"110000100",
  44342=>"000100010",
  44343=>"101100011",
  44344=>"000011100",
  44345=>"111011010",
  44346=>"001111010",
  44347=>"110001000",
  44348=>"001010010",
  44349=>"000010001",
  44350=>"000111111",
  44351=>"100011100",
  44352=>"000100100",
  44353=>"100101110",
  44354=>"010001101",
  44355=>"011100000",
  44356=>"101101111",
  44357=>"111101011",
  44358=>"110101010",
  44359=>"100010001",
  44360=>"100010110",
  44361=>"110101110",
  44362=>"101001001",
  44363=>"011110001",
  44364=>"011111100",
  44365=>"100100101",
  44366=>"011011000",
  44367=>"010000011",
  44368=>"100101111",
  44369=>"001101100",
  44370=>"011110101",
  44371=>"000011111",
  44372=>"011101101",
  44373=>"000111000",
  44374=>"001100100",
  44375=>"011100001",
  44376=>"010000000",
  44377=>"110011101",
  44378=>"100010110",
  44379=>"111101101",
  44380=>"001000101",
  44381=>"011010010",
  44382=>"101001101",
  44383=>"011100110",
  44384=>"100110110",
  44385=>"101011011",
  44386=>"000011010",
  44387=>"111000111",
  44388=>"001011001",
  44389=>"000001011",
  44390=>"100101101",
  44391=>"001001101",
  44392=>"001111001",
  44393=>"001110010",
  44394=>"001001110",
  44395=>"001100010",
  44396=>"010010110",
  44397=>"000001010",
  44398=>"110111000",
  44399=>"010001101",
  44400=>"100000000",
  44401=>"100010010",
  44402=>"110000011",
  44403=>"001100001",
  44404=>"101100000",
  44405=>"110111010",
  44406=>"111000000",
  44407=>"100001011",
  44408=>"000011000",
  44409=>"011001000",
  44410=>"010001101",
  44411=>"011011010",
  44412=>"110011000",
  44413=>"011010100",
  44414=>"011100101",
  44415=>"000001011",
  44416=>"111111111",
  44417=>"100100000",
  44418=>"111101100",
  44419=>"111010000",
  44420=>"111100001",
  44421=>"010110000",
  44422=>"101111010",
  44423=>"100110110",
  44424=>"011101100",
  44425=>"111001010",
  44426=>"000010110",
  44427=>"000000001",
  44428=>"100001110",
  44429=>"101100101",
  44430=>"011000001",
  44431=>"110001110",
  44432=>"111110111",
  44433=>"101000001",
  44434=>"100000110",
  44435=>"110101110",
  44436=>"111001101",
  44437=>"000000110",
  44438=>"001000011",
  44439=>"011000000",
  44440=>"111100000",
  44441=>"010011000",
  44442=>"110101010",
  44443=>"111010011",
  44444=>"111001001",
  44445=>"011011000",
  44446=>"111011110",
  44447=>"011001001",
  44448=>"100001011",
  44449=>"000001100",
  44450=>"011111111",
  44451=>"110110000",
  44452=>"000100000",
  44453=>"100010010",
  44454=>"101000000",
  44455=>"110011000",
  44456=>"010011110",
  44457=>"011011000",
  44458=>"010111000",
  44459=>"100111110",
  44460=>"100011100",
  44461=>"101111100",
  44462=>"011101100",
  44463=>"010101110",
  44464=>"011011100",
  44465=>"110011100",
  44466=>"100111111",
  44467=>"000011000",
  44468=>"101110110",
  44469=>"111100001",
  44470=>"001011101",
  44471=>"100100111",
  44472=>"011000001",
  44473=>"101101101",
  44474=>"101000010",
  44475=>"110101010",
  44476=>"000110000",
  44477=>"000001010",
  44478=>"000101110",
  44479=>"010101111",
  44480=>"000110101",
  44481=>"000111101",
  44482=>"111100010",
  44483=>"110001000",
  44484=>"000011000",
  44485=>"011011100",
  44486=>"000001001",
  44487=>"010010101",
  44488=>"010100101",
  44489=>"010001111",
  44490=>"100010100",
  44491=>"110101100",
  44492=>"000000110",
  44493=>"101110100",
  44494=>"010011000",
  44495=>"000010110",
  44496=>"101011011",
  44497=>"011111100",
  44498=>"101010001",
  44499=>"010111000",
  44500=>"100111011",
  44501=>"101000001",
  44502=>"110001111",
  44503=>"011010101",
  44504=>"110011010",
  44505=>"001010011",
  44506=>"000000110",
  44507=>"100101001",
  44508=>"111101010",
  44509=>"110001101",
  44510=>"000001110",
  44511=>"101010110",
  44512=>"001111101",
  44513=>"010100000",
  44514=>"110100000",
  44515=>"111001111",
  44516=>"111011101",
  44517=>"001101101",
  44518=>"011011011",
  44519=>"011100010",
  44520=>"001101110",
  44521=>"011110101",
  44522=>"000010100",
  44523=>"011010100",
  44524=>"110101011",
  44525=>"110101000",
  44526=>"101111000",
  44527=>"101111011",
  44528=>"001110001",
  44529=>"111000101",
  44530=>"000100001",
  44531=>"000000000",
  44532=>"111011011",
  44533=>"001010110",
  44534=>"101000001",
  44535=>"000111100",
  44536=>"000000000",
  44537=>"110101010",
  44538=>"010000000",
  44539=>"110011010",
  44540=>"100001111",
  44541=>"011000001",
  44542=>"111111000",
  44543=>"111100110",
  44544=>"001001100",
  44545=>"011101101",
  44546=>"001100111",
  44547=>"110101001",
  44548=>"011010001",
  44549=>"101000011",
  44550=>"111000000",
  44551=>"111010101",
  44552=>"000110001",
  44553=>"101110010",
  44554=>"000111111",
  44555=>"101011101",
  44556=>"000100110",
  44557=>"110011111",
  44558=>"010010100",
  44559=>"101011001",
  44560=>"100100001",
  44561=>"110000110",
  44562=>"011011100",
  44563=>"101101001",
  44564=>"000000100",
  44565=>"000000100",
  44566=>"100111111",
  44567=>"001010100",
  44568=>"010001011",
  44569=>"111100011",
  44570=>"101000010",
  44571=>"000010111",
  44572=>"110011101",
  44573=>"100011000",
  44574=>"111111101",
  44575=>"000110111",
  44576=>"011111000",
  44577=>"101110110",
  44578=>"000110010",
  44579=>"000111000",
  44580=>"011100100",
  44581=>"011010110",
  44582=>"011001010",
  44583=>"101001001",
  44584=>"110111100",
  44585=>"110101101",
  44586=>"101111010",
  44587=>"010000010",
  44588=>"100000000",
  44589=>"111111010",
  44590=>"001101000",
  44591=>"101110011",
  44592=>"101111010",
  44593=>"001111001",
  44594=>"101010010",
  44595=>"001001001",
  44596=>"011111000",
  44597=>"111101100",
  44598=>"000010101",
  44599=>"100101000",
  44600=>"000001000",
  44601=>"000101100",
  44602=>"000101100",
  44603=>"100100001",
  44604=>"000000111",
  44605=>"110011011",
  44606=>"111100001",
  44607=>"110110100",
  44608=>"000111001",
  44609=>"100011010",
  44610=>"010100010",
  44611=>"110111110",
  44612=>"010100110",
  44613=>"110100000",
  44614=>"011010100",
  44615=>"111111111",
  44616=>"000100100",
  44617=>"101010100",
  44618=>"001000010",
  44619=>"101110001",
  44620=>"001101111",
  44621=>"101101010",
  44622=>"110111100",
  44623=>"001101101",
  44624=>"000101101",
  44625=>"110100101",
  44626=>"101100001",
  44627=>"011011111",
  44628=>"110001100",
  44629=>"000001000",
  44630=>"010101001",
  44631=>"000010111",
  44632=>"001111010",
  44633=>"101000101",
  44634=>"111010100",
  44635=>"011011010",
  44636=>"100000111",
  44637=>"011110100",
  44638=>"001000111",
  44639=>"111110101",
  44640=>"111100000",
  44641=>"101000001",
  44642=>"101011010",
  44643=>"110111011",
  44644=>"101000010",
  44645=>"111011110",
  44646=>"000011100",
  44647=>"111011001",
  44648=>"000010010",
  44649=>"000010000",
  44650=>"001000100",
  44651=>"001001101",
  44652=>"000101111",
  44653=>"001011100",
  44654=>"011100011",
  44655=>"011111000",
  44656=>"001100101",
  44657=>"001001000",
  44658=>"011111111",
  44659=>"011011011",
  44660=>"010100011",
  44661=>"110111111",
  44662=>"010101001",
  44663=>"000010010",
  44664=>"100101111",
  44665=>"011000010",
  44666=>"000101100",
  44667=>"010000100",
  44668=>"110001001",
  44669=>"101000100",
  44670=>"100101111",
  44671=>"011100110",
  44672=>"101100101",
  44673=>"100011001",
  44674=>"001100001",
  44675=>"000110011",
  44676=>"000110011",
  44677=>"000000011",
  44678=>"100010000",
  44679=>"101110111",
  44680=>"111100010",
  44681=>"000000101",
  44682=>"110011110",
  44683=>"100100101",
  44684=>"101011001",
  44685=>"110010111",
  44686=>"100010001",
  44687=>"101001111",
  44688=>"111100110",
  44689=>"101100101",
  44690=>"010111101",
  44691=>"010111100",
  44692=>"011011101",
  44693=>"010100011",
  44694=>"111111011",
  44695=>"001000011",
  44696=>"011011011",
  44697=>"111110110",
  44698=>"111110101",
  44699=>"101101111",
  44700=>"011001101",
  44701=>"010000001",
  44702=>"011010000",
  44703=>"001111110",
  44704=>"010011000",
  44705=>"000001010",
  44706=>"111110101",
  44707=>"001011101",
  44708=>"111101100",
  44709=>"010100100",
  44710=>"111101111",
  44711=>"001010101",
  44712=>"100010111",
  44713=>"000000010",
  44714=>"001110111",
  44715=>"010100001",
  44716=>"110010111",
  44717=>"011110100",
  44718=>"100110101",
  44719=>"011001011",
  44720=>"010111111",
  44721=>"000100111",
  44722=>"111111100",
  44723=>"011111101",
  44724=>"100000010",
  44725=>"010011001",
  44726=>"101100101",
  44727=>"100010001",
  44728=>"001100100",
  44729=>"111101000",
  44730=>"110011010",
  44731=>"111000000",
  44732=>"101111000",
  44733=>"100010010",
  44734=>"100000001",
  44735=>"111001111",
  44736=>"101100101",
  44737=>"100000001",
  44738=>"011110111",
  44739=>"100101111",
  44740=>"010011001",
  44741=>"000011011",
  44742=>"000101011",
  44743=>"000101010",
  44744=>"011000011",
  44745=>"010101111",
  44746=>"101111001",
  44747=>"101010101",
  44748=>"100010101",
  44749=>"000001101",
  44750=>"110100001",
  44751=>"100011100",
  44752=>"100000111",
  44753=>"000001110",
  44754=>"101110100",
  44755=>"011001011",
  44756=>"110101101",
  44757=>"110010000",
  44758=>"010000111",
  44759=>"011011000",
  44760=>"000001100",
  44761=>"000110010",
  44762=>"000011110",
  44763=>"001100100",
  44764=>"000001110",
  44765=>"000101001",
  44766=>"101000000",
  44767=>"111100101",
  44768=>"010111011",
  44769=>"110100001",
  44770=>"100111001",
  44771=>"000010111",
  44772=>"011010111",
  44773=>"001110101",
  44774=>"110101100",
  44775=>"010000111",
  44776=>"000100111",
  44777=>"011011101",
  44778=>"000100110",
  44779=>"101001111",
  44780=>"101101011",
  44781=>"000011010",
  44782=>"011110000",
  44783=>"011000001",
  44784=>"010101100",
  44785=>"010011000",
  44786=>"010100000",
  44787=>"111000111",
  44788=>"111000011",
  44789=>"000110100",
  44790=>"111101111",
  44791=>"000100011",
  44792=>"110001000",
  44793=>"111110110",
  44794=>"100001110",
  44795=>"001101010",
  44796=>"100011010",
  44797=>"011101000",
  44798=>"100010001",
  44799=>"010011000",
  44800=>"000101000",
  44801=>"000100101",
  44802=>"010110110",
  44803=>"100100001",
  44804=>"001010100",
  44805=>"101100000",
  44806=>"110110111",
  44807=>"111000000",
  44808=>"001100111",
  44809=>"001010000",
  44810=>"101001011",
  44811=>"110100101",
  44812=>"110010000",
  44813=>"101011000",
  44814=>"011101000",
  44815=>"110111011",
  44816=>"011110000",
  44817=>"000000100",
  44818=>"101111110",
  44819=>"111101011",
  44820=>"101100110",
  44821=>"111000111",
  44822=>"111010001",
  44823=>"110101001",
  44824=>"000101110",
  44825=>"111100101",
  44826=>"001000111",
  44827=>"001001100",
  44828=>"010101010",
  44829=>"010011000",
  44830=>"100010011",
  44831=>"110001010",
  44832=>"001011111",
  44833=>"111100111",
  44834=>"111010010",
  44835=>"111110000",
  44836=>"100011110",
  44837=>"000010010",
  44838=>"011011011",
  44839=>"111011001",
  44840=>"010010001",
  44841=>"111111001",
  44842=>"011111111",
  44843=>"101011100",
  44844=>"101000010",
  44845=>"000000010",
  44846=>"001011000",
  44847=>"110101101",
  44848=>"001011101",
  44849=>"011100010",
  44850=>"111110001",
  44851=>"001010100",
  44852=>"001000011",
  44853=>"110110011",
  44854=>"010000000",
  44855=>"100100011",
  44856=>"010000001",
  44857=>"000000010",
  44858=>"101110101",
  44859=>"010101100",
  44860=>"101100111",
  44861=>"110100010",
  44862=>"111011001",
  44863=>"001100011",
  44864=>"101010111",
  44865=>"001010110",
  44866=>"010001011",
  44867=>"000011111",
  44868=>"010111110",
  44869=>"110011000",
  44870=>"001101010",
  44871=>"010000111",
  44872=>"100100100",
  44873=>"111111111",
  44874=>"010110000",
  44875=>"001000100",
  44876=>"100000001",
  44877=>"110000100",
  44878=>"000111000",
  44879=>"111110010",
  44880=>"010000011",
  44881=>"111101011",
  44882=>"000110111",
  44883=>"101011100",
  44884=>"110110110",
  44885=>"011000101",
  44886=>"001100111",
  44887=>"000001011",
  44888=>"001000001",
  44889=>"011010011",
  44890=>"000101010",
  44891=>"101000100",
  44892=>"001010100",
  44893=>"001100111",
  44894=>"000010001",
  44895=>"001000100",
  44896=>"010010010",
  44897=>"100000111",
  44898=>"000000000",
  44899=>"000000110",
  44900=>"101010001",
  44901=>"011100000",
  44902=>"000010100",
  44903=>"110110111",
  44904=>"010101010",
  44905=>"100110101",
  44906=>"010110001",
  44907=>"011000110",
  44908=>"010001110",
  44909=>"111101111",
  44910=>"110100000",
  44911=>"011100110",
  44912=>"100111011",
  44913=>"111101101",
  44914=>"100100100",
  44915=>"001011001",
  44916=>"011010100",
  44917=>"011111010",
  44918=>"000000011",
  44919=>"000010011",
  44920=>"101001100",
  44921=>"001000010",
  44922=>"110001100",
  44923=>"101000011",
  44924=>"001110001",
  44925=>"000100011",
  44926=>"101100111",
  44927=>"101111111",
  44928=>"100110011",
  44929=>"110011001",
  44930=>"011011011",
  44931=>"001000101",
  44932=>"001101000",
  44933=>"101010010",
  44934=>"101100111",
  44935=>"001010001",
  44936=>"101001111",
  44937=>"001111110",
  44938=>"101000111",
  44939=>"100111011",
  44940=>"011110111",
  44941=>"001011100",
  44942=>"010010111",
  44943=>"111100110",
  44944=>"100101011",
  44945=>"111011001",
  44946=>"010001100",
  44947=>"111110001",
  44948=>"101100000",
  44949=>"010111100",
  44950=>"100110111",
  44951=>"011110001",
  44952=>"111010000",
  44953=>"000000100",
  44954=>"000101110",
  44955=>"000000000",
  44956=>"111111000",
  44957=>"110110000",
  44958=>"110010011",
  44959=>"000101111",
  44960=>"111100110",
  44961=>"100101011",
  44962=>"111001101",
  44963=>"011111000",
  44964=>"100110010",
  44965=>"010111010",
  44966=>"000000001",
  44967=>"110000000",
  44968=>"001001000",
  44969=>"010000011",
  44970=>"111010101",
  44971=>"100111110",
  44972=>"101000011",
  44973=>"011001011",
  44974=>"001011011",
  44975=>"110000101",
  44976=>"000010100",
  44977=>"001110010",
  44978=>"011110010",
  44979=>"100011010",
  44980=>"111011010",
  44981=>"001101000",
  44982=>"101110110",
  44983=>"011101111",
  44984=>"110010101",
  44985=>"001001010",
  44986=>"110111100",
  44987=>"011100101",
  44988=>"000001001",
  44989=>"111000101",
  44990=>"110100110",
  44991=>"110111101",
  44992=>"111000111",
  44993=>"101111110",
  44994=>"101000111",
  44995=>"111000000",
  44996=>"100000010",
  44997=>"010011111",
  44998=>"011000001",
  44999=>"000110101",
  45000=>"000110111",
  45001=>"011100000",
  45002=>"101010100",
  45003=>"111110111",
  45004=>"001110010",
  45005=>"101100011",
  45006=>"100100010",
  45007=>"011010101",
  45008=>"001111110",
  45009=>"100011011",
  45010=>"100101110",
  45011=>"100100001",
  45012=>"000011100",
  45013=>"101010110",
  45014=>"010100000",
  45015=>"010000110",
  45016=>"111101111",
  45017=>"101011000",
  45018=>"111100001",
  45019=>"000110010",
  45020=>"011110101",
  45021=>"010001101",
  45022=>"110010101",
  45023=>"110010010",
  45024=>"111010000",
  45025=>"101110100",
  45026=>"000011111",
  45027=>"001101000",
  45028=>"000101101",
  45029=>"110101110",
  45030=>"010010110",
  45031=>"111100001",
  45032=>"011011010",
  45033=>"000111111",
  45034=>"110001010",
  45035=>"110011111",
  45036=>"000100111",
  45037=>"101010011",
  45038=>"010001110",
  45039=>"001110110",
  45040=>"011001101",
  45041=>"110000101",
  45042=>"010000010",
  45043=>"011101001",
  45044=>"000111010",
  45045=>"100000010",
  45046=>"000000010",
  45047=>"110101111",
  45048=>"111111111",
  45049=>"111010100",
  45050=>"111011111",
  45051=>"111101001",
  45052=>"100110000",
  45053=>"011100001",
  45054=>"011110011",
  45055=>"001011011",
  45056=>"110101000",
  45057=>"101001001",
  45058=>"000010110",
  45059=>"101111100",
  45060=>"111101100",
  45061=>"110111100",
  45062=>"011010001",
  45063=>"000001000",
  45064=>"011010010",
  45065=>"000000011",
  45066=>"101001110",
  45067=>"110101001",
  45068=>"111111101",
  45069=>"010100011",
  45070=>"000011111",
  45071=>"101111001",
  45072=>"101001001",
  45073=>"110001100",
  45074=>"001111000",
  45075=>"000101111",
  45076=>"000011100",
  45077=>"000101011",
  45078=>"100111101",
  45079=>"011010011",
  45080=>"000111011",
  45081=>"111111110",
  45082=>"111100101",
  45083=>"110111001",
  45084=>"001001110",
  45085=>"011111011",
  45086=>"001001110",
  45087=>"011000000",
  45088=>"100010001",
  45089=>"100010101",
  45090=>"000110101",
  45091=>"001101100",
  45092=>"101100111",
  45093=>"001000010",
  45094=>"100000010",
  45095=>"011100001",
  45096=>"011011011",
  45097=>"000000101",
  45098=>"100101100",
  45099=>"100110001",
  45100=>"100010000",
  45101=>"111011101",
  45102=>"110111111",
  45103=>"100100001",
  45104=>"100011001",
  45105=>"111001100",
  45106=>"011010110",
  45107=>"100111101",
  45108=>"100011010",
  45109=>"101000010",
  45110=>"010000101",
  45111=>"101011101",
  45112=>"100101110",
  45113=>"110011011",
  45114=>"011011101",
  45115=>"111000100",
  45116=>"111110111",
  45117=>"111001111",
  45118=>"100101010",
  45119=>"010101010",
  45120=>"110011010",
  45121=>"010011001",
  45122=>"110111011",
  45123=>"100010000",
  45124=>"001010101",
  45125=>"110000101",
  45126=>"000000100",
  45127=>"011010101",
  45128=>"100110001",
  45129=>"111001101",
  45130=>"000001011",
  45131=>"000000100",
  45132=>"110000100",
  45133=>"110011101",
  45134=>"010010010",
  45135=>"000001101",
  45136=>"100111001",
  45137=>"111111111",
  45138=>"110011011",
  45139=>"100100110",
  45140=>"010000011",
  45141=>"001000001",
  45142=>"011110100",
  45143=>"000000001",
  45144=>"000011010",
  45145=>"001000011",
  45146=>"110010000",
  45147=>"001100001",
  45148=>"011010110",
  45149=>"100110010",
  45150=>"110101101",
  45151=>"000101110",
  45152=>"111000101",
  45153=>"100110011",
  45154=>"001101000",
  45155=>"001010001",
  45156=>"111100000",
  45157=>"001000000",
  45158=>"000101101",
  45159=>"011010101",
  45160=>"000001001",
  45161=>"001100101",
  45162=>"010101000",
  45163=>"001100010",
  45164=>"101010011",
  45165=>"100000011",
  45166=>"001101000",
  45167=>"100110000",
  45168=>"111001001",
  45169=>"101001010",
  45170=>"000010110",
  45171=>"000011111",
  45172=>"010000111",
  45173=>"111101111",
  45174=>"100100010",
  45175=>"100101111",
  45176=>"010100010",
  45177=>"000000111",
  45178=>"101111110",
  45179=>"111110100",
  45180=>"111110000",
  45181=>"100110010",
  45182=>"101110101",
  45183=>"110110101",
  45184=>"110010000",
  45185=>"000111110",
  45186=>"101100000",
  45187=>"001100000",
  45188=>"110101111",
  45189=>"000010011",
  45190=>"110101101",
  45191=>"101110000",
  45192=>"100110110",
  45193=>"101111001",
  45194=>"111100100",
  45195=>"000001111",
  45196=>"101001100",
  45197=>"101100101",
  45198=>"101100010",
  45199=>"001001101",
  45200=>"011110000",
  45201=>"111101101",
  45202=>"100011111",
  45203=>"011001011",
  45204=>"100100111",
  45205=>"101100001",
  45206=>"111000000",
  45207=>"110000111",
  45208=>"000101000",
  45209=>"111100111",
  45210=>"010111110",
  45211=>"000100000",
  45212=>"011000010",
  45213=>"111110000",
  45214=>"001011100",
  45215=>"010000100",
  45216=>"100001101",
  45217=>"000001000",
  45218=>"001100010",
  45219=>"100000010",
  45220=>"010010111",
  45221=>"100010000",
  45222=>"110000111",
  45223=>"101000101",
  45224=>"011111111",
  45225=>"000001011",
  45226=>"100000111",
  45227=>"111111111",
  45228=>"010011001",
  45229=>"010111111",
  45230=>"010101101",
  45231=>"010100001",
  45232=>"100100001",
  45233=>"001100001",
  45234=>"111101000",
  45235=>"111001000",
  45236=>"010010011",
  45237=>"110011010",
  45238=>"010111000",
  45239=>"001000001",
  45240=>"100110111",
  45241=>"100101100",
  45242=>"101100011",
  45243=>"011110111",
  45244=>"011001001",
  45245=>"100110001",
  45246=>"100000001",
  45247=>"000010101",
  45248=>"101001111",
  45249=>"101101110",
  45250=>"000111100",
  45251=>"011011000",
  45252=>"010110011",
  45253=>"110111011",
  45254=>"111011001",
  45255=>"101001110",
  45256=>"000010010",
  45257=>"010011000",
  45258=>"100110100",
  45259=>"110010100",
  45260=>"101011010",
  45261=>"110000110",
  45262=>"001111111",
  45263=>"011000001",
  45264=>"110010011",
  45265=>"111001101",
  45266=>"101000000",
  45267=>"111100111",
  45268=>"011110111",
  45269=>"111001111",
  45270=>"010011110",
  45271=>"001111011",
  45272=>"101010110",
  45273=>"011111010",
  45274=>"111000011",
  45275=>"100010111",
  45276=>"111010111",
  45277=>"100100010",
  45278=>"111111101",
  45279=>"011010101",
  45280=>"100000100",
  45281=>"111011100",
  45282=>"100100100",
  45283=>"111100101",
  45284=>"010100011",
  45285=>"011011100",
  45286=>"111111110",
  45287=>"111001110",
  45288=>"101010001",
  45289=>"111011101",
  45290=>"101110010",
  45291=>"000001100",
  45292=>"001101111",
  45293=>"111101111",
  45294=>"001100000",
  45295=>"101000000",
  45296=>"100011011",
  45297=>"101111011",
  45298=>"010111001",
  45299=>"000101000",
  45300=>"100100001",
  45301=>"111010101",
  45302=>"110111111",
  45303=>"001001001",
  45304=>"011001100",
  45305=>"111100101",
  45306=>"011111000",
  45307=>"000100000",
  45308=>"000001010",
  45309=>"011011010",
  45310=>"011000111",
  45311=>"100001001",
  45312=>"001100110",
  45313=>"001001001",
  45314=>"101000101",
  45315=>"101010110",
  45316=>"010101111",
  45317=>"010000110",
  45318=>"100010001",
  45319=>"101001101",
  45320=>"000100010",
  45321=>"001100000",
  45322=>"010010001",
  45323=>"110000000",
  45324=>"000100101",
  45325=>"011010000",
  45326=>"110000000",
  45327=>"101100100",
  45328=>"000001111",
  45329=>"010001101",
  45330=>"011101100",
  45331=>"011011000",
  45332=>"001010001",
  45333=>"100111000",
  45334=>"110010101",
  45335=>"110110110",
  45336=>"000001010",
  45337=>"001001001",
  45338=>"101010011",
  45339=>"100011111",
  45340=>"001100011",
  45341=>"001010111",
  45342=>"111110010",
  45343=>"000000001",
  45344=>"011000000",
  45345=>"010010011",
  45346=>"101111110",
  45347=>"101000101",
  45348=>"000101010",
  45349=>"000100011",
  45350=>"001101110",
  45351=>"111100001",
  45352=>"000101101",
  45353=>"001010100",
  45354=>"100000110",
  45355=>"100000110",
  45356=>"111111011",
  45357=>"000100001",
  45358=>"000100001",
  45359=>"101010101",
  45360=>"100011101",
  45361=>"100011111",
  45362=>"010100010",
  45363=>"100111100",
  45364=>"011110110",
  45365=>"001101100",
  45366=>"010010100",
  45367=>"010110011",
  45368=>"001000001",
  45369=>"000010001",
  45370=>"011100100",
  45371=>"000001010",
  45372=>"100011001",
  45373=>"101111000",
  45374=>"110101001",
  45375=>"111011100",
  45376=>"101010001",
  45377=>"101110000",
  45378=>"111100110",
  45379=>"000111111",
  45380=>"111111111",
  45381=>"011110111",
  45382=>"000001101",
  45383=>"000001100",
  45384=>"101001101",
  45385=>"110110101",
  45386=>"101011110",
  45387=>"111101101",
  45388=>"101010000",
  45389=>"101001011",
  45390=>"100111010",
  45391=>"000011001",
  45392=>"101000110",
  45393=>"011100000",
  45394=>"111010100",
  45395=>"000100100",
  45396=>"001001011",
  45397=>"000100100",
  45398=>"110001101",
  45399=>"101000111",
  45400=>"000010011",
  45401=>"100100010",
  45402=>"101001001",
  45403=>"111011001",
  45404=>"110111100",
  45405=>"011100011",
  45406=>"111010010",
  45407=>"110010111",
  45408=>"000111110",
  45409=>"001111110",
  45410=>"110011101",
  45411=>"100000110",
  45412=>"100110100",
  45413=>"111111101",
  45414=>"111111100",
  45415=>"100110111",
  45416=>"010110010",
  45417=>"010110001",
  45418=>"000010110",
  45419=>"101011100",
  45420=>"000100010",
  45421=>"001110000",
  45422=>"111101111",
  45423=>"010111011",
  45424=>"011100101",
  45425=>"000111010",
  45426=>"111101110",
  45427=>"000010110",
  45428=>"001010001",
  45429=>"010100110",
  45430=>"000111001",
  45431=>"001101011",
  45432=>"101111101",
  45433=>"101010110",
  45434=>"000010010",
  45435=>"000000011",
  45436=>"111110011",
  45437=>"111110100",
  45438=>"111101100",
  45439=>"100111100",
  45440=>"001111101",
  45441=>"001000110",
  45442=>"110100010",
  45443=>"100111110",
  45444=>"010111001",
  45445=>"000011110",
  45446=>"110111110",
  45447=>"100111001",
  45448=>"001011001",
  45449=>"111100011",
  45450=>"110011010",
  45451=>"101000001",
  45452=>"011101011",
  45453=>"111010110",
  45454=>"000000111",
  45455=>"111111011",
  45456=>"011000110",
  45457=>"111100000",
  45458=>"001111111",
  45459=>"010100001",
  45460=>"101110111",
  45461=>"101101111",
  45462=>"100100101",
  45463=>"111001111",
  45464=>"110000000",
  45465=>"000001010",
  45466=>"101010100",
  45467=>"111001110",
  45468=>"000101111",
  45469=>"111000011",
  45470=>"101000110",
  45471=>"010011100",
  45472=>"101100101",
  45473=>"010001000",
  45474=>"010001110",
  45475=>"000001000",
  45476=>"010010011",
  45477=>"111101000",
  45478=>"111111110",
  45479=>"101100110",
  45480=>"100010011",
  45481=>"010010001",
  45482=>"101011011",
  45483=>"100011000",
  45484=>"010110110",
  45485=>"101111000",
  45486=>"011001001",
  45487=>"011110011",
  45488=>"111111001",
  45489=>"101101110",
  45490=>"111111101",
  45491=>"001000001",
  45492=>"011100011",
  45493=>"101110100",
  45494=>"100110000",
  45495=>"111011011",
  45496=>"100011110",
  45497=>"001001110",
  45498=>"001011100",
  45499=>"010101110",
  45500=>"111110100",
  45501=>"010111011",
  45502=>"101000000",
  45503=>"100011010",
  45504=>"111010101",
  45505=>"010010010",
  45506=>"000101110",
  45507=>"110011110",
  45508=>"100001111",
  45509=>"110100011",
  45510=>"010000010",
  45511=>"000000100",
  45512=>"001001001",
  45513=>"101100000",
  45514=>"100101111",
  45515=>"111010011",
  45516=>"100111010",
  45517=>"010011111",
  45518=>"100000001",
  45519=>"001001111",
  45520=>"000000100",
  45521=>"111111101",
  45522=>"000010110",
  45523=>"100001101",
  45524=>"001011010",
  45525=>"110000111",
  45526=>"001010000",
  45527=>"111100101",
  45528=>"001100100",
  45529=>"011001100",
  45530=>"011111111",
  45531=>"111000110",
  45532=>"001010001",
  45533=>"111111110",
  45534=>"101100000",
  45535=>"100001001",
  45536=>"001011100",
  45537=>"110011001",
  45538=>"111000111",
  45539=>"101010001",
  45540=>"010011001",
  45541=>"101011101",
  45542=>"111100111",
  45543=>"000000000",
  45544=>"010101010",
  45545=>"110100101",
  45546=>"100100101",
  45547=>"001000111",
  45548=>"101011111",
  45549=>"001101111",
  45550=>"011010010",
  45551=>"000000010",
  45552=>"101000000",
  45553=>"001011111",
  45554=>"010111000",
  45555=>"001000001",
  45556=>"110100111",
  45557=>"000110001",
  45558=>"011101110",
  45559=>"100100100",
  45560=>"001111111",
  45561=>"111001111",
  45562=>"100101100",
  45563=>"101000101",
  45564=>"000100100",
  45565=>"000000111",
  45566=>"101011101",
  45567=>"010001101",
  45568=>"011100110",
  45569=>"000111111",
  45570=>"101111101",
  45571=>"001101101",
  45572=>"110000000",
  45573=>"010101000",
  45574=>"111010011",
  45575=>"111111011",
  45576=>"111011111",
  45577=>"011100010",
  45578=>"111010000",
  45579=>"000101001",
  45580=>"100100111",
  45581=>"010010011",
  45582=>"110001001",
  45583=>"011011001",
  45584=>"111010001",
  45585=>"010010110",
  45586=>"011010001",
  45587=>"011101101",
  45588=>"110011110",
  45589=>"011101110",
  45590=>"010100111",
  45591=>"011101110",
  45592=>"111010101",
  45593=>"101001101",
  45594=>"111001011",
  45595=>"111111110",
  45596=>"111001000",
  45597=>"000000010",
  45598=>"111100001",
  45599=>"110000110",
  45600=>"100000000",
  45601=>"110000011",
  45602=>"000010000",
  45603=>"000110111",
  45604=>"001100000",
  45605=>"110110100",
  45606=>"110010010",
  45607=>"001110110",
  45608=>"010111111",
  45609=>"101000100",
  45610=>"101100100",
  45611=>"001000110",
  45612=>"001101011",
  45613=>"101010111",
  45614=>"100100000",
  45615=>"100011100",
  45616=>"110110111",
  45617=>"100101100",
  45618=>"011110110",
  45619=>"111000010",
  45620=>"100111101",
  45621=>"110100110",
  45622=>"110011100",
  45623=>"010000110",
  45624=>"010011101",
  45625=>"110101111",
  45626=>"110110110",
  45627=>"001011110",
  45628=>"000100100",
  45629=>"100011111",
  45630=>"110101100",
  45631=>"101100100",
  45632=>"100000101",
  45633=>"100010110",
  45634=>"011001010",
  45635=>"010111001",
  45636=>"100010000",
  45637=>"111100011",
  45638=>"001000110",
  45639=>"111101011",
  45640=>"000000010",
  45641=>"001001110",
  45642=>"011101101",
  45643=>"101010000",
  45644=>"100110111",
  45645=>"100101100",
  45646=>"111111111",
  45647=>"000010010",
  45648=>"110011110",
  45649=>"010110100",
  45650=>"100111100",
  45651=>"010100111",
  45652=>"101110001",
  45653=>"010000100",
  45654=>"000101010",
  45655=>"010000111",
  45656=>"000010001",
  45657=>"000001100",
  45658=>"011111100",
  45659=>"000100001",
  45660=>"000001001",
  45661=>"000110000",
  45662=>"100000001",
  45663=>"000101111",
  45664=>"100101010",
  45665=>"001010001",
  45666=>"101000010",
  45667=>"010100001",
  45668=>"101001011",
  45669=>"000100100",
  45670=>"110101010",
  45671=>"101101110",
  45672=>"011001000",
  45673=>"110010000",
  45674=>"010001101",
  45675=>"100100001",
  45676=>"110010110",
  45677=>"000100110",
  45678=>"111100010",
  45679=>"010011111",
  45680=>"110001110",
  45681=>"110000010",
  45682=>"100010011",
  45683=>"011101011",
  45684=>"100001010",
  45685=>"010000111",
  45686=>"111100000",
  45687=>"010111011",
  45688=>"000010011",
  45689=>"101000110",
  45690=>"000111111",
  45691=>"100001110",
  45692=>"111000111",
  45693=>"011110101",
  45694=>"101110101",
  45695=>"110010001",
  45696=>"110010101",
  45697=>"001110111",
  45698=>"111101111",
  45699=>"100110100",
  45700=>"001101011",
  45701=>"111010000",
  45702=>"100000010",
  45703=>"110110000",
  45704=>"111101011",
  45705=>"111000011",
  45706=>"100000000",
  45707=>"011000011",
  45708=>"010101100",
  45709=>"010100010",
  45710=>"001100100",
  45711=>"000101000",
  45712=>"110010011",
  45713=>"110000111",
  45714=>"111101100",
  45715=>"100101000",
  45716=>"010100000",
  45717=>"110001000",
  45718=>"100000010",
  45719=>"101010010",
  45720=>"010101001",
  45721=>"010010011",
  45722=>"000111010",
  45723=>"001001111",
  45724=>"011010101",
  45725=>"100011111",
  45726=>"000111101",
  45727=>"011000111",
  45728=>"111101111",
  45729=>"100000111",
  45730=>"000011111",
  45731=>"000001110",
  45732=>"111001100",
  45733=>"010001000",
  45734=>"101100100",
  45735=>"101110010",
  45736=>"011011011",
  45737=>"011010011",
  45738=>"100110111",
  45739=>"101110010",
  45740=>"111011000",
  45741=>"110001010",
  45742=>"001001010",
  45743=>"001001011",
  45744=>"001010100",
  45745=>"000011000",
  45746=>"010101111",
  45747=>"100101110",
  45748=>"010111101",
  45749=>"110001011",
  45750=>"110011110",
  45751=>"010111011",
  45752=>"110100101",
  45753=>"111000010",
  45754=>"110111101",
  45755=>"110011100",
  45756=>"001000001",
  45757=>"011011101",
  45758=>"100001100",
  45759=>"111110000",
  45760=>"010100111",
  45761=>"000110101",
  45762=>"110001001",
  45763=>"001101101",
  45764=>"110100100",
  45765=>"000011001",
  45766=>"000110100",
  45767=>"110010001",
  45768=>"101000100",
  45769=>"000001000",
  45770=>"011101100",
  45771=>"010100001",
  45772=>"111100101",
  45773=>"100111001",
  45774=>"111010101",
  45775=>"011010000",
  45776=>"010011010",
  45777=>"110110000",
  45778=>"011101000",
  45779=>"001100001",
  45780=>"111100111",
  45781=>"010011011",
  45782=>"110010111",
  45783=>"110011001",
  45784=>"111111101",
  45785=>"000001011",
  45786=>"101010000",
  45787=>"110101101",
  45788=>"001000111",
  45789=>"110000101",
  45790=>"010011010",
  45791=>"101010011",
  45792=>"110000011",
  45793=>"100000100",
  45794=>"111101101",
  45795=>"111001000",
  45796=>"010011000",
  45797=>"110101010",
  45798=>"101010000",
  45799=>"000011110",
  45800=>"000110000",
  45801=>"100000010",
  45802=>"111000011",
  45803=>"011110011",
  45804=>"001001000",
  45805=>"101110001",
  45806=>"010011000",
  45807=>"001011011",
  45808=>"001010110",
  45809=>"000111010",
  45810=>"101111100",
  45811=>"100100100",
  45812=>"101100000",
  45813=>"000111111",
  45814=>"011000111",
  45815=>"011010010",
  45816=>"001101000",
  45817=>"010101010",
  45818=>"101000010",
  45819=>"011111110",
  45820=>"000101001",
  45821=>"011011101",
  45822=>"100010001",
  45823=>"101011110",
  45824=>"010010110",
  45825=>"000001011",
  45826=>"011110010",
  45827=>"101100010",
  45828=>"000010111",
  45829=>"101000000",
  45830=>"010110001",
  45831=>"110011100",
  45832=>"000111011",
  45833=>"100111000",
  45834=>"100101011",
  45835=>"100001010",
  45836=>"010100101",
  45837=>"000001011",
  45838=>"011011011",
  45839=>"111110111",
  45840=>"011010010",
  45841=>"101000110",
  45842=>"100100011",
  45843=>"011010111",
  45844=>"010001010",
  45845=>"110011001",
  45846=>"010100101",
  45847=>"001111010",
  45848=>"001001001",
  45849=>"110000101",
  45850=>"101111010",
  45851=>"000101101",
  45852=>"011110000",
  45853=>"100111111",
  45854=>"101101011",
  45855=>"001011001",
  45856=>"010000100",
  45857=>"111001010",
  45858=>"100010000",
  45859=>"100000100",
  45860=>"111100001",
  45861=>"111101111",
  45862=>"010010100",
  45863=>"010100011",
  45864=>"100010111",
  45865=>"001000000",
  45866=>"111100001",
  45867=>"000110001",
  45868=>"010101010",
  45869=>"011001101",
  45870=>"000111100",
  45871=>"110110110",
  45872=>"000100101",
  45873=>"000001011",
  45874=>"000101010",
  45875=>"010100100",
  45876=>"101011111",
  45877=>"001100101",
  45878=>"001110001",
  45879=>"011001000",
  45880=>"100101111",
  45881=>"001110000",
  45882=>"011111100",
  45883=>"111011010",
  45884=>"001100001",
  45885=>"000010011",
  45886=>"000000101",
  45887=>"111111110",
  45888=>"001110001",
  45889=>"101000010",
  45890=>"000000101",
  45891=>"100000100",
  45892=>"101110000",
  45893=>"111110111",
  45894=>"101100010",
  45895=>"000101001",
  45896=>"011100100",
  45897=>"001100111",
  45898=>"111110011",
  45899=>"001110101",
  45900=>"101010100",
  45901=>"110011011",
  45902=>"110011010",
  45903=>"111110011",
  45904=>"101101101",
  45905=>"100100010",
  45906=>"101010101",
  45907=>"000110111",
  45908=>"100010101",
  45909=>"000011010",
  45910=>"111000001",
  45911=>"100110101",
  45912=>"011100011",
  45913=>"101001100",
  45914=>"110101000",
  45915=>"101100111",
  45916=>"010011101",
  45917=>"110110011",
  45918=>"101011010",
  45919=>"100110110",
  45920=>"000000001",
  45921=>"111011001",
  45922=>"000010000",
  45923=>"001000001",
  45924=>"000000111",
  45925=>"110100101",
  45926=>"000010000",
  45927=>"010000011",
  45928=>"011001001",
  45929=>"011011110",
  45930=>"011000001",
  45931=>"100000110",
  45932=>"010000000",
  45933=>"000000001",
  45934=>"100110001",
  45935=>"000110010",
  45936=>"101010001",
  45937=>"110011000",
  45938=>"111111010",
  45939=>"000000011",
  45940=>"000001000",
  45941=>"101001110",
  45942=>"111100011",
  45943=>"011100000",
  45944=>"111010000",
  45945=>"100010100",
  45946=>"010010111",
  45947=>"011011011",
  45948=>"111101111",
  45949=>"110001101",
  45950=>"101100101",
  45951=>"100011101",
  45952=>"110011110",
  45953=>"100000100",
  45954=>"110001000",
  45955=>"101101011",
  45956=>"110001010",
  45957=>"011100011",
  45958=>"101000000",
  45959=>"001000001",
  45960=>"101010101",
  45961=>"001101011",
  45962=>"110100110",
  45963=>"010000110",
  45964=>"011011101",
  45965=>"010000100",
  45966=>"011011000",
  45967=>"010101100",
  45968=>"110110001",
  45969=>"111111111",
  45970=>"101101101",
  45971=>"100001101",
  45972=>"001011000",
  45973=>"010101100",
  45974=>"001001000",
  45975=>"100011011",
  45976=>"110110010",
  45977=>"001111111",
  45978=>"110011100",
  45979=>"100101101",
  45980=>"000001001",
  45981=>"000011000",
  45982=>"101111010",
  45983=>"100101010",
  45984=>"010010010",
  45985=>"010000101",
  45986=>"000100111",
  45987=>"000101100",
  45988=>"100110101",
  45989=>"010110111",
  45990=>"000110000",
  45991=>"100001000",
  45992=>"111101111",
  45993=>"000000100",
  45994=>"100101001",
  45995=>"000101111",
  45996=>"100010001",
  45997=>"110011111",
  45998=>"010100110",
  45999=>"110100111",
  46000=>"101001000",
  46001=>"111111011",
  46002=>"011011000",
  46003=>"001011011",
  46004=>"000111111",
  46005=>"011110111",
  46006=>"001011000",
  46007=>"111000010",
  46008=>"101100101",
  46009=>"010011110",
  46010=>"010011010",
  46011=>"011010000",
  46012=>"011000001",
  46013=>"110011101",
  46014=>"110110101",
  46015=>"001101001",
  46016=>"111011100",
  46017=>"101010010",
  46018=>"111110100",
  46019=>"000001001",
  46020=>"000010110",
  46021=>"011111001",
  46022=>"110101101",
  46023=>"100010001",
  46024=>"010000011",
  46025=>"000101001",
  46026=>"100011001",
  46027=>"100010101",
  46028=>"111101100",
  46029=>"100111100",
  46030=>"000100000",
  46031=>"110010111",
  46032=>"101110011",
  46033=>"110110010",
  46034=>"101111001",
  46035=>"101010000",
  46036=>"111111111",
  46037=>"101011011",
  46038=>"111101011",
  46039=>"001110100",
  46040=>"110110000",
  46041=>"001101110",
  46042=>"101011000",
  46043=>"100110101",
  46044=>"001000100",
  46045=>"010000001",
  46046=>"100010110",
  46047=>"101110000",
  46048=>"101010011",
  46049=>"001011100",
  46050=>"001110111",
  46051=>"100010111",
  46052=>"101001111",
  46053=>"101101001",
  46054=>"100000110",
  46055=>"111101010",
  46056=>"000001010",
  46057=>"011001010",
  46058=>"101001111",
  46059=>"101000110",
  46060=>"000011010",
  46061=>"011001001",
  46062=>"011011111",
  46063=>"100011010",
  46064=>"001001111",
  46065=>"111101000",
  46066=>"111010111",
  46067=>"010101000",
  46068=>"101110100",
  46069=>"000000111",
  46070=>"101110111",
  46071=>"001010010",
  46072=>"001000100",
  46073=>"001100011",
  46074=>"000101100",
  46075=>"010011111",
  46076=>"101111111",
  46077=>"010000011",
  46078=>"010000001",
  46079=>"000001000",
  46080=>"111010111",
  46081=>"100100010",
  46082=>"001011011",
  46083=>"000011011",
  46084=>"101000001",
  46085=>"100101000",
  46086=>"010010000",
  46087=>"000000101",
  46088=>"011100000",
  46089=>"111000100",
  46090=>"101100101",
  46091=>"110011100",
  46092=>"000000000",
  46093=>"000100100",
  46094=>"001100111",
  46095=>"101101001",
  46096=>"000110001",
  46097=>"101101110",
  46098=>"110011110",
  46099=>"110001100",
  46100=>"000101101",
  46101=>"101011001",
  46102=>"100011100",
  46103=>"011101001",
  46104=>"110100110",
  46105=>"110000010",
  46106=>"001111001",
  46107=>"101101100",
  46108=>"011000111",
  46109=>"001100111",
  46110=>"011111100",
  46111=>"000100011",
  46112=>"001011100",
  46113=>"101001100",
  46114=>"101111101",
  46115=>"011100001",
  46116=>"000000011",
  46117=>"011101000",
  46118=>"111111011",
  46119=>"001001011",
  46120=>"011010100",
  46121=>"100000010",
  46122=>"010000001",
  46123=>"110110010",
  46124=>"011010100",
  46125=>"111111101",
  46126=>"000110000",
  46127=>"010110111",
  46128=>"111111101",
  46129=>"101111101",
  46130=>"100000110",
  46131=>"101100111",
  46132=>"110101000",
  46133=>"001000000",
  46134=>"111110110",
  46135=>"100100010",
  46136=>"110001101",
  46137=>"101101100",
  46138=>"100000111",
  46139=>"110010111",
  46140=>"111000101",
  46141=>"111011100",
  46142=>"011001100",
  46143=>"010101000",
  46144=>"101110000",
  46145=>"000011010",
  46146=>"100111100",
  46147=>"110100010",
  46148=>"000111111",
  46149=>"100111011",
  46150=>"000001111",
  46151=>"111001011",
  46152=>"010101000",
  46153=>"000001000",
  46154=>"010010110",
  46155=>"100010101",
  46156=>"101101101",
  46157=>"111101100",
  46158=>"000010100",
  46159=>"110001001",
  46160=>"010001001",
  46161=>"110000101",
  46162=>"000101110",
  46163=>"000010001",
  46164=>"001100010",
  46165=>"111000111",
  46166=>"000011110",
  46167=>"101001110",
  46168=>"010011001",
  46169=>"100011100",
  46170=>"010010111",
  46171=>"000111110",
  46172=>"100001011",
  46173=>"001000010",
  46174=>"100011101",
  46175=>"110011001",
  46176=>"001101000",
  46177=>"001110111",
  46178=>"100111010",
  46179=>"101011001",
  46180=>"010010010",
  46181=>"101011001",
  46182=>"111100101",
  46183=>"000011010",
  46184=>"101110101",
  46185=>"010101110",
  46186=>"000011010",
  46187=>"100010000",
  46188=>"011100101",
  46189=>"000001111",
  46190=>"110111011",
  46191=>"111101101",
  46192=>"001100011",
  46193=>"010100001",
  46194=>"101011001",
  46195=>"101110111",
  46196=>"110111000",
  46197=>"010000111",
  46198=>"110111101",
  46199=>"010111001",
  46200=>"010011000",
  46201=>"011001010",
  46202=>"101010001",
  46203=>"010001101",
  46204=>"011010000",
  46205=>"100000010",
  46206=>"111101111",
  46207=>"110001111",
  46208=>"010011110",
  46209=>"100101111",
  46210=>"001011000",
  46211=>"101001001",
  46212=>"111111111",
  46213=>"010001000",
  46214=>"010100101",
  46215=>"101100100",
  46216=>"100101111",
  46217=>"000111010",
  46218=>"110000000",
  46219=>"101011001",
  46220=>"101111101",
  46221=>"001010100",
  46222=>"110011011",
  46223=>"110111000",
  46224=>"101000111",
  46225=>"000010111",
  46226=>"111111011",
  46227=>"100110100",
  46228=>"101001111",
  46229=>"100110110",
  46230=>"010000010",
  46231=>"001011001",
  46232=>"010101000",
  46233=>"010001000",
  46234=>"111111100",
  46235=>"110011010",
  46236=>"101010010",
  46237=>"110011101",
  46238=>"000011111",
  46239=>"100000011",
  46240=>"010110010",
  46241=>"111111000",
  46242=>"011110111",
  46243=>"010000100",
  46244=>"000111010",
  46245=>"000100111",
  46246=>"110000011",
  46247=>"011100110",
  46248=>"111110100",
  46249=>"100001111",
  46250=>"110100100",
  46251=>"101111110",
  46252=>"100010001",
  46253=>"010010101",
  46254=>"111110001",
  46255=>"000001100",
  46256=>"010010111",
  46257=>"000000101",
  46258=>"010111101",
  46259=>"010100100",
  46260=>"010101110",
  46261=>"110110010",
  46262=>"101101000",
  46263=>"100100011",
  46264=>"010011010",
  46265=>"011101110",
  46266=>"000001101",
  46267=>"111111100",
  46268=>"100011000",
  46269=>"111000101",
  46270=>"000111111",
  46271=>"111000011",
  46272=>"010011011",
  46273=>"010100010",
  46274=>"011111111",
  46275=>"101000101",
  46276=>"101100111",
  46277=>"011010010",
  46278=>"100100010",
  46279=>"001000111",
  46280=>"110111111",
  46281=>"110111010",
  46282=>"001111100",
  46283=>"111001101",
  46284=>"010000001",
  46285=>"011011000",
  46286=>"110110111",
  46287=>"100011110",
  46288=>"101000111",
  46289=>"000100001",
  46290=>"001011011",
  46291=>"001111000",
  46292=>"101011011",
  46293=>"010000110",
  46294=>"100001001",
  46295=>"011100001",
  46296=>"100010101",
  46297=>"010010011",
  46298=>"000001011",
  46299=>"010011111",
  46300=>"011110001",
  46301=>"101100100",
  46302=>"111011101",
  46303=>"111100000",
  46304=>"000101111",
  46305=>"000101101",
  46306=>"111011100",
  46307=>"001011000",
  46308=>"010001111",
  46309=>"010001010",
  46310=>"000000100",
  46311=>"010101000",
  46312=>"111000111",
  46313=>"110101100",
  46314=>"001010000",
  46315=>"111101110",
  46316=>"100011010",
  46317=>"101111010",
  46318=>"111111101",
  46319=>"001110110",
  46320=>"101111011",
  46321=>"001010000",
  46322=>"010100100",
  46323=>"010010011",
  46324=>"111101000",
  46325=>"101101000",
  46326=>"010110111",
  46327=>"110100111",
  46328=>"111010010",
  46329=>"011100111",
  46330=>"101101110",
  46331=>"100101110",
  46332=>"110100010",
  46333=>"001110000",
  46334=>"110000100",
  46335=>"011111111",
  46336=>"110100100",
  46337=>"010001100",
  46338=>"100100111",
  46339=>"110100001",
  46340=>"001110111",
  46341=>"100100101",
  46342=>"010010111",
  46343=>"001111000",
  46344=>"101010110",
  46345=>"101010010",
  46346=>"110110111",
  46347=>"011010001",
  46348=>"111011110",
  46349=>"000001111",
  46350=>"100110101",
  46351=>"111000011",
  46352=>"111110010",
  46353=>"011101011",
  46354=>"011101001",
  46355=>"110111100",
  46356=>"100111110",
  46357=>"000111101",
  46358=>"000100100",
  46359=>"111111000",
  46360=>"011011010",
  46361=>"111100010",
  46362=>"011110010",
  46363=>"010010101",
  46364=>"101000110",
  46365=>"110110001",
  46366=>"000110011",
  46367=>"011010101",
  46368=>"101101010",
  46369=>"011100001",
  46370=>"001011011",
  46371=>"011000000",
  46372=>"101001001",
  46373=>"101100001",
  46374=>"001110100",
  46375=>"010011011",
  46376=>"101110100",
  46377=>"101001000",
  46378=>"111100010",
  46379=>"010010001",
  46380=>"010010100",
  46381=>"100000000",
  46382=>"100000110",
  46383=>"110110101",
  46384=>"000111011",
  46385=>"010101000",
  46386=>"010111011",
  46387=>"011001111",
  46388=>"010010111",
  46389=>"101010111",
  46390=>"011100110",
  46391=>"101111011",
  46392=>"000101000",
  46393=>"110000101",
  46394=>"001111011",
  46395=>"111111010",
  46396=>"111001011",
  46397=>"110100000",
  46398=>"011110000",
  46399=>"010101010",
  46400=>"110110000",
  46401=>"001010010",
  46402=>"001000100",
  46403=>"000100000",
  46404=>"011011001",
  46405=>"110010001",
  46406=>"111100011",
  46407=>"111101110",
  46408=>"000001100",
  46409=>"011000000",
  46410=>"011101110",
  46411=>"111000110",
  46412=>"111110000",
  46413=>"001000000",
  46414=>"000000011",
  46415=>"000010010",
  46416=>"010000011",
  46417=>"101001110",
  46418=>"101011111",
  46419=>"101011011",
  46420=>"110000000",
  46421=>"010000111",
  46422=>"101001100",
  46423=>"000000001",
  46424=>"110000111",
  46425=>"110110011",
  46426=>"010101101",
  46427=>"110001010",
  46428=>"001100111",
  46429=>"000100110",
  46430=>"111100101",
  46431=>"000010000",
  46432=>"000110001",
  46433=>"011101111",
  46434=>"110100010",
  46435=>"101010011",
  46436=>"100011100",
  46437=>"000001010",
  46438=>"100000111",
  46439=>"000111001",
  46440=>"000110100",
  46441=>"100100101",
  46442=>"001011111",
  46443=>"000001110",
  46444=>"110001100",
  46445=>"101000000",
  46446=>"101011001",
  46447=>"111000111",
  46448=>"001110001",
  46449=>"000100110",
  46450=>"010000110",
  46451=>"000110101",
  46452=>"110000001",
  46453=>"100010111",
  46454=>"110011100",
  46455=>"101110111",
  46456=>"000110111",
  46457=>"011110000",
  46458=>"010010010",
  46459=>"111010010",
  46460=>"000000100",
  46461=>"000010100",
  46462=>"001101100",
  46463=>"110101001",
  46464=>"000011110",
  46465=>"010000000",
  46466=>"110011101",
  46467=>"010010111",
  46468=>"111011100",
  46469=>"100101111",
  46470=>"101111111",
  46471=>"000111100",
  46472=>"010001110",
  46473=>"110111100",
  46474=>"011111011",
  46475=>"011000000",
  46476=>"011010111",
  46477=>"000011111",
  46478=>"011111111",
  46479=>"011101101",
  46480=>"100111000",
  46481=>"011101100",
  46482=>"001000111",
  46483=>"100010110",
  46484=>"010010010",
  46485=>"101010110",
  46486=>"110000101",
  46487=>"110111001",
  46488=>"001100101",
  46489=>"011000000",
  46490=>"010101000",
  46491=>"010101111",
  46492=>"101111101",
  46493=>"011101110",
  46494=>"001101001",
  46495=>"100001011",
  46496=>"001101101",
  46497=>"011100000",
  46498=>"001000110",
  46499=>"100001101",
  46500=>"101110000",
  46501=>"010010101",
  46502=>"010100111",
  46503=>"000001110",
  46504=>"100011011",
  46505=>"111001110",
  46506=>"001001010",
  46507=>"001110011",
  46508=>"011001001",
  46509=>"110101100",
  46510=>"001000100",
  46511=>"001011101",
  46512=>"111100100",
  46513=>"100101010",
  46514=>"100101100",
  46515=>"000000110",
  46516=>"011101010",
  46517=>"001001100",
  46518=>"011000110",
  46519=>"111101111",
  46520=>"001110010",
  46521=>"010110101",
  46522=>"000000100",
  46523=>"100100011",
  46524=>"101111111",
  46525=>"111001101",
  46526=>"110011011",
  46527=>"101111111",
  46528=>"101010110",
  46529=>"111110000",
  46530=>"101001001",
  46531=>"111111100",
  46532=>"101110111",
  46533=>"001110001",
  46534=>"010101000",
  46535=>"000000100",
  46536=>"101111000",
  46537=>"111110011",
  46538=>"101000011",
  46539=>"010111000",
  46540=>"000000110",
  46541=>"001100111",
  46542=>"000101000",
  46543=>"101101101",
  46544=>"101101101",
  46545=>"110010011",
  46546=>"110010011",
  46547=>"111110110",
  46548=>"001111011",
  46549=>"100100101",
  46550=>"000101101",
  46551=>"101000001",
  46552=>"111011000",
  46553=>"101001000",
  46554=>"000101100",
  46555=>"111100000",
  46556=>"111100010",
  46557=>"111001001",
  46558=>"010011011",
  46559=>"000111101",
  46560=>"100000111",
  46561=>"101111111",
  46562=>"101100100",
  46563=>"001000101",
  46564=>"001111001",
  46565=>"011100111",
  46566=>"111001101",
  46567=>"101001011",
  46568=>"111000011",
  46569=>"001001001",
  46570=>"100001011",
  46571=>"010110100",
  46572=>"010101110",
  46573=>"011010100",
  46574=>"101010000",
  46575=>"001000100",
  46576=>"110000011",
  46577=>"001000111",
  46578=>"010100010",
  46579=>"111101011",
  46580=>"111111011",
  46581=>"110110010",
  46582=>"011100001",
  46583=>"110000111",
  46584=>"000101001",
  46585=>"000010010",
  46586=>"001010001",
  46587=>"000000100",
  46588=>"000001100",
  46589=>"011011111",
  46590=>"001111000",
  46591=>"010000001",
  46592=>"011011000",
  46593=>"011111111",
  46594=>"111000111",
  46595=>"100101010",
  46596=>"011000100",
  46597=>"101001101",
  46598=>"000100101",
  46599=>"010100001",
  46600=>"001001101",
  46601=>"010001011",
  46602=>"110111101",
  46603=>"000110000",
  46604=>"010000001",
  46605=>"000000111",
  46606=>"111001111",
  46607=>"011001001",
  46608=>"001111011",
  46609=>"001100011",
  46610=>"011110000",
  46611=>"010001111",
  46612=>"010001011",
  46613=>"010000111",
  46614=>"100111111",
  46615=>"011111011",
  46616=>"100110100",
  46617=>"011000001",
  46618=>"110011001",
  46619=>"111000010",
  46620=>"110111110",
  46621=>"001010100",
  46622=>"111010001",
  46623=>"000100001",
  46624=>"111010111",
  46625=>"010001100",
  46626=>"101011010",
  46627=>"010110010",
  46628=>"011010111",
  46629=>"011000111",
  46630=>"101010011",
  46631=>"011000011",
  46632=>"101100111",
  46633=>"001000101",
  46634=>"010110001",
  46635=>"000111101",
  46636=>"001010101",
  46637=>"100100000",
  46638=>"000000001",
  46639=>"000001000",
  46640=>"101100110",
  46641=>"101101010",
  46642=>"001010110",
  46643=>"011100111",
  46644=>"110010001",
  46645=>"011100000",
  46646=>"101010000",
  46647=>"100100111",
  46648=>"010001111",
  46649=>"110001100",
  46650=>"011100000",
  46651=>"100101110",
  46652=>"100001000",
  46653=>"111100101",
  46654=>"111101110",
  46655=>"111011001",
  46656=>"011011100",
  46657=>"001110001",
  46658=>"101100110",
  46659=>"010010000",
  46660=>"011010111",
  46661=>"011101001",
  46662=>"111101001",
  46663=>"001101110",
  46664=>"110011100",
  46665=>"111110000",
  46666=>"001110101",
  46667=>"000110001",
  46668=>"111101011",
  46669=>"000101100",
  46670=>"101101000",
  46671=>"100100010",
  46672=>"001101100",
  46673=>"010111011",
  46674=>"110001010",
  46675=>"010100001",
  46676=>"100011101",
  46677=>"010010010",
  46678=>"000100010",
  46679=>"110010101",
  46680=>"111001101",
  46681=>"101001110",
  46682=>"101011001",
  46683=>"101011011",
  46684=>"101100011",
  46685=>"101101100",
  46686=>"111111100",
  46687=>"001011111",
  46688=>"000100001",
  46689=>"010010110",
  46690=>"100011111",
  46691=>"011010010",
  46692=>"100100011",
  46693=>"001010101",
  46694=>"010000000",
  46695=>"011010000",
  46696=>"101110001",
  46697=>"011111011",
  46698=>"011000111",
  46699=>"011100011",
  46700=>"111111110",
  46701=>"000100110",
  46702=>"101101101",
  46703=>"101110100",
  46704=>"000100010",
  46705=>"010100001",
  46706=>"001000010",
  46707=>"111001000",
  46708=>"010100010",
  46709=>"110010111",
  46710=>"101001001",
  46711=>"010011011",
  46712=>"110100011",
  46713=>"101000000",
  46714=>"011110111",
  46715=>"010010010",
  46716=>"110010001",
  46717=>"010111010",
  46718=>"010001101",
  46719=>"110000001",
  46720=>"100011001",
  46721=>"111000000",
  46722=>"111110111",
  46723=>"011000011",
  46724=>"000010100",
  46725=>"100000001",
  46726=>"010001010",
  46727=>"010010100",
  46728=>"110111000",
  46729=>"000000011",
  46730=>"101110101",
  46731=>"101111110",
  46732=>"000010011",
  46733=>"001011001",
  46734=>"101010000",
  46735=>"010000110",
  46736=>"110101000",
  46737=>"011101010",
  46738=>"000111011",
  46739=>"101100011",
  46740=>"101101001",
  46741=>"011110100",
  46742=>"111110110",
  46743=>"111000101",
  46744=>"011010111",
  46745=>"010100110",
  46746=>"101111010",
  46747=>"110001111",
  46748=>"100000001",
  46749=>"010011000",
  46750=>"010011010",
  46751=>"100010011",
  46752=>"100110011",
  46753=>"101101100",
  46754=>"111000100",
  46755=>"111100101",
  46756=>"100110110",
  46757=>"000100110",
  46758=>"010010100",
  46759=>"000001110",
  46760=>"010100100",
  46761=>"000000101",
  46762=>"100001110",
  46763=>"110011001",
  46764=>"100100110",
  46765=>"100101011",
  46766=>"110100111",
  46767=>"100001011",
  46768=>"100100010",
  46769=>"011000101",
  46770=>"110101011",
  46771=>"110101001",
  46772=>"001011000",
  46773=>"101000101",
  46774=>"000110000",
  46775=>"010011101",
  46776=>"100110100",
  46777=>"011111011",
  46778=>"001100001",
  46779=>"100010110",
  46780=>"110001100",
  46781=>"010000000",
  46782=>"011000010",
  46783=>"111111110",
  46784=>"100000111",
  46785=>"100011010",
  46786=>"100101110",
  46787=>"011110010",
  46788=>"011001110",
  46789=>"000101111",
  46790=>"111110100",
  46791=>"100011110",
  46792=>"111001101",
  46793=>"001010110",
  46794=>"101000001",
  46795=>"111100001",
  46796=>"111111010",
  46797=>"010000000",
  46798=>"011000001",
  46799=>"100101011",
  46800=>"111000010",
  46801=>"101011110",
  46802=>"000010000",
  46803=>"101001001",
  46804=>"011101101",
  46805=>"000010110",
  46806=>"010010000",
  46807=>"011001101",
  46808=>"110000111",
  46809=>"111110010",
  46810=>"101000100",
  46811=>"101010000",
  46812=>"111011011",
  46813=>"010100111",
  46814=>"101010110",
  46815=>"001111100",
  46816=>"100011000",
  46817=>"001110101",
  46818=>"101001100",
  46819=>"100010000",
  46820=>"011111001",
  46821=>"001000111",
  46822=>"101101001",
  46823=>"101110001",
  46824=>"111001000",
  46825=>"101111011",
  46826=>"010111000",
  46827=>"001000111",
  46828=>"011100101",
  46829=>"111101010",
  46830=>"100001111",
  46831=>"100010010",
  46832=>"110110000",
  46833=>"110000001",
  46834=>"000010100",
  46835=>"101010111",
  46836=>"110011001",
  46837=>"011101100",
  46838=>"110011111",
  46839=>"000001000",
  46840=>"011111111",
  46841=>"100100001",
  46842=>"001100111",
  46843=>"101101000",
  46844=>"101110100",
  46845=>"111011001",
  46846=>"001011001",
  46847=>"010110001",
  46848=>"010101010",
  46849=>"111100011",
  46850=>"100101110",
  46851=>"000100001",
  46852=>"011111111",
  46853=>"100100111",
  46854=>"110001010",
  46855=>"101001111",
  46856=>"000101111",
  46857=>"000100000",
  46858=>"110000101",
  46859=>"101010010",
  46860=>"110010111",
  46861=>"000011110",
  46862=>"011010110",
  46863=>"011001111",
  46864=>"010110000",
  46865=>"101101000",
  46866=>"100101110",
  46867=>"100001101",
  46868=>"100110111",
  46869=>"000110000",
  46870=>"111111110",
  46871=>"100001110",
  46872=>"100111101",
  46873=>"110101100",
  46874=>"100101011",
  46875=>"101000011",
  46876=>"100110011",
  46877=>"010111001",
  46878=>"100100101",
  46879=>"100100010",
  46880=>"110011010",
  46881=>"000101101",
  46882=>"000110010",
  46883=>"110100000",
  46884=>"001000101",
  46885=>"000000000",
  46886=>"001001000",
  46887=>"100001110",
  46888=>"111011110",
  46889=>"110111011",
  46890=>"011010110",
  46891=>"110110110",
  46892=>"001001110",
  46893=>"011111111",
  46894=>"111010010",
  46895=>"100100111",
  46896=>"101101000",
  46897=>"000010000",
  46898=>"100100100",
  46899=>"001101000",
  46900=>"011000000",
  46901=>"111000011",
  46902=>"010010111",
  46903=>"101101111",
  46904=>"001001010",
  46905=>"100001101",
  46906=>"100010011",
  46907=>"000011010",
  46908=>"001011100",
  46909=>"110000110",
  46910=>"111001110",
  46911=>"000000010",
  46912=>"100000001",
  46913=>"101111101",
  46914=>"111011110",
  46915=>"100000101",
  46916=>"010111110",
  46917=>"100111011",
  46918=>"000001000",
  46919=>"001001010",
  46920=>"100000000",
  46921=>"010010001",
  46922=>"011011111",
  46923=>"001100101",
  46924=>"011000100",
  46925=>"011110011",
  46926=>"010101101",
  46927=>"000111101",
  46928=>"000001111",
  46929=>"100100001",
  46930=>"100001110",
  46931=>"011001011",
  46932=>"011111110",
  46933=>"000000011",
  46934=>"100001110",
  46935=>"101111011",
  46936=>"101000100",
  46937=>"111011110",
  46938=>"011010001",
  46939=>"110001100",
  46940=>"100001011",
  46941=>"000100000",
  46942=>"110010111",
  46943=>"110110001",
  46944=>"100000111",
  46945=>"010000110",
  46946=>"100001101",
  46947=>"101011110",
  46948=>"101011110",
  46949=>"001000111",
  46950=>"111101101",
  46951=>"010100010",
  46952=>"111111100",
  46953=>"011100100",
  46954=>"010000101",
  46955=>"011010110",
  46956=>"100001101",
  46957=>"101111001",
  46958=>"011001001",
  46959=>"000000000",
  46960=>"011011111",
  46961=>"001011001",
  46962=>"100010010",
  46963=>"100010010",
  46964=>"011111111",
  46965=>"010010000",
  46966=>"110010010",
  46967=>"011000111",
  46968=>"110111111",
  46969=>"000010011",
  46970=>"111111011",
  46971=>"111111100",
  46972=>"111111101",
  46973=>"000110101",
  46974=>"010011110",
  46975=>"111111100",
  46976=>"101001101",
  46977=>"100001110",
  46978=>"100010000",
  46979=>"110100111",
  46980=>"010110101",
  46981=>"101011001",
  46982=>"010000101",
  46983=>"110000011",
  46984=>"111010101",
  46985=>"111111100",
  46986=>"111101010",
  46987=>"111001011",
  46988=>"010011101",
  46989=>"100111011",
  46990=>"011001000",
  46991=>"001101000",
  46992=>"000110110",
  46993=>"001001001",
  46994=>"001000110",
  46995=>"000000100",
  46996=>"000000011",
  46997=>"001100100",
  46998=>"110100110",
  46999=>"011111100",
  47000=>"111010110",
  47001=>"000000100",
  47002=>"000010001",
  47003=>"110111110",
  47004=>"111011101",
  47005=>"111010100",
  47006=>"101100111",
  47007=>"001100101",
  47008=>"110001111",
  47009=>"011001010",
  47010=>"000011101",
  47011=>"011000000",
  47012=>"101101001",
  47013=>"001011010",
  47014=>"100010010",
  47015=>"011011101",
  47016=>"000001110",
  47017=>"100101011",
  47018=>"011100111",
  47019=>"000010010",
  47020=>"011000000",
  47021=>"101100011",
  47022=>"111111000",
  47023=>"111111000",
  47024=>"110111011",
  47025=>"101110000",
  47026=>"100100111",
  47027=>"010000100",
  47028=>"111010001",
  47029=>"011100110",
  47030=>"010001010",
  47031=>"110101110",
  47032=>"110001010",
  47033=>"010101000",
  47034=>"111011001",
  47035=>"110011000",
  47036=>"010001001",
  47037=>"000011011",
  47038=>"000100101",
  47039=>"111110110",
  47040=>"101101111",
  47041=>"110000101",
  47042=>"111101001",
  47043=>"011001101",
  47044=>"011111001",
  47045=>"110110101",
  47046=>"111111001",
  47047=>"100110110",
  47048=>"000100011",
  47049=>"110011011",
  47050=>"101101110",
  47051=>"111111000",
  47052=>"001100110",
  47053=>"111010100",
  47054=>"000101101",
  47055=>"101101011",
  47056=>"110100101",
  47057=>"101110010",
  47058=>"000110101",
  47059=>"010001100",
  47060=>"111111001",
  47061=>"111110000",
  47062=>"000010000",
  47063=>"000100111",
  47064=>"011000001",
  47065=>"111100000",
  47066=>"010111110",
  47067=>"010100010",
  47068=>"111100001",
  47069=>"001000010",
  47070=>"111011110",
  47071=>"111000101",
  47072=>"001000111",
  47073=>"010010001",
  47074=>"111111110",
  47075=>"010010111",
  47076=>"010010000",
  47077=>"100000001",
  47078=>"011100101",
  47079=>"000100110",
  47080=>"000000000",
  47081=>"100100001",
  47082=>"101001111",
  47083=>"011001101",
  47084=>"011010010",
  47085=>"101011100",
  47086=>"010100010",
  47087=>"000000110",
  47088=>"011010010",
  47089=>"110000000",
  47090=>"011010101",
  47091=>"010010101",
  47092=>"101100001",
  47093=>"011110000",
  47094=>"000000100",
  47095=>"000111111",
  47096=>"111101111",
  47097=>"100011111",
  47098=>"111011111",
  47099=>"010010000",
  47100=>"010001011",
  47101=>"100111000",
  47102=>"111001100",
  47103=>"110000011",
  47104=>"110010010",
  47105=>"000001110",
  47106=>"001010111",
  47107=>"001100110",
  47108=>"000000100",
  47109=>"001100111",
  47110=>"011110101",
  47111=>"100000000",
  47112=>"101111100",
  47113=>"100111101",
  47114=>"111101110",
  47115=>"011100101",
  47116=>"000101110",
  47117=>"100001010",
  47118=>"010010011",
  47119=>"000110010",
  47120=>"110101011",
  47121=>"111110000",
  47122=>"100101100",
  47123=>"101001000",
  47124=>"001100110",
  47125=>"100000010",
  47126=>"101110100",
  47127=>"000101011",
  47128=>"001010110",
  47129=>"101010011",
  47130=>"110001010",
  47131=>"011100101",
  47132=>"011011001",
  47133=>"000000110",
  47134=>"100010111",
  47135=>"100100010",
  47136=>"000001110",
  47137=>"101000001",
  47138=>"010011110",
  47139=>"000011101",
  47140=>"101101011",
  47141=>"011001001",
  47142=>"000101011",
  47143=>"001000100",
  47144=>"011011110",
  47145=>"111011111",
  47146=>"000111101",
  47147=>"000011011",
  47148=>"011110101",
  47149=>"010101101",
  47150=>"011000011",
  47151=>"101001000",
  47152=>"110010110",
  47153=>"110100110",
  47154=>"101000001",
  47155=>"101010100",
  47156=>"111110100",
  47157=>"111011100",
  47158=>"000101110",
  47159=>"001011101",
  47160=>"000110001",
  47161=>"110000011",
  47162=>"000011010",
  47163=>"011010101",
  47164=>"111101100",
  47165=>"010111000",
  47166=>"100000010",
  47167=>"000001010",
  47168=>"000000000",
  47169=>"001000010",
  47170=>"011000000",
  47171=>"000100011",
  47172=>"010101110",
  47173=>"110000000",
  47174=>"110101101",
  47175=>"010000000",
  47176=>"110010100",
  47177=>"100110010",
  47178=>"111100001",
  47179=>"101000010",
  47180=>"000011111",
  47181=>"001110011",
  47182=>"111110011",
  47183=>"111000111",
  47184=>"111011101",
  47185=>"010111100",
  47186=>"011101110",
  47187=>"100101001",
  47188=>"000101100",
  47189=>"110011010",
  47190=>"000011101",
  47191=>"110000010",
  47192=>"010011111",
  47193=>"001101111",
  47194=>"100010100",
  47195=>"011010010",
  47196=>"011011100",
  47197=>"000010101",
  47198=>"000101011",
  47199=>"010001001",
  47200=>"110001101",
  47201=>"100100111",
  47202=>"100000100",
  47203=>"000000100",
  47204=>"000001011",
  47205=>"111011110",
  47206=>"110100010",
  47207=>"010101101",
  47208=>"011001010",
  47209=>"100111110",
  47210=>"100000110",
  47211=>"011001000",
  47212=>"011111101",
  47213=>"100011000",
  47214=>"010101011",
  47215=>"001000111",
  47216=>"110010000",
  47217=>"110010010",
  47218=>"100100001",
  47219=>"000010001",
  47220=>"101100100",
  47221=>"001100110",
  47222=>"001011110",
  47223=>"100111101",
  47224=>"101000000",
  47225=>"000100000",
  47226=>"110010100",
  47227=>"000001100",
  47228=>"000011001",
  47229=>"110100111",
  47230=>"000000110",
  47231=>"101000110",
  47232=>"001010111",
  47233=>"011111001",
  47234=>"001111000",
  47235=>"111110101",
  47236=>"110111011",
  47237=>"111101001",
  47238=>"011010011",
  47239=>"001001010",
  47240=>"000010011",
  47241=>"000100101",
  47242=>"000111101",
  47243=>"111101001",
  47244=>"000000000",
  47245=>"111101000",
  47246=>"011100010",
  47247=>"000101010",
  47248=>"000011110",
  47249=>"110111101",
  47250=>"111111011",
  47251=>"110100001",
  47252=>"000010011",
  47253=>"000011011",
  47254=>"110011011",
  47255=>"110110011",
  47256=>"000100110",
  47257=>"111010100",
  47258=>"001001110",
  47259=>"110110011",
  47260=>"000110001",
  47261=>"011001011",
  47262=>"110010100",
  47263=>"010001100",
  47264=>"001010101",
  47265=>"101001101",
  47266=>"100101000",
  47267=>"100101000",
  47268=>"101011111",
  47269=>"100010110",
  47270=>"011011001",
  47271=>"100010101",
  47272=>"111011110",
  47273=>"111111110",
  47274=>"000011001",
  47275=>"101001110",
  47276=>"000111110",
  47277=>"101011111",
  47278=>"010000011",
  47279=>"100010001",
  47280=>"010111010",
  47281=>"010011101",
  47282=>"100000100",
  47283=>"100100011",
  47284=>"011110000",
  47285=>"010101011",
  47286=>"110111011",
  47287=>"000001001",
  47288=>"100000101",
  47289=>"000010011",
  47290=>"100111111",
  47291=>"101100000",
  47292=>"010101101",
  47293=>"110010100",
  47294=>"000001010",
  47295=>"001000100",
  47296=>"011000111",
  47297=>"010010000",
  47298=>"100000100",
  47299=>"101010111",
  47300=>"000111011",
  47301=>"011010100",
  47302=>"011110011",
  47303=>"100011010",
  47304=>"011111101",
  47305=>"000000010",
  47306=>"101111000",
  47307=>"111110110",
  47308=>"011111000",
  47309=>"111100011",
  47310=>"010010100",
  47311=>"000111111",
  47312=>"111100011",
  47313=>"101011110",
  47314=>"000100111",
  47315=>"000011111",
  47316=>"100111000",
  47317=>"110001111",
  47318=>"110011101",
  47319=>"100011100",
  47320=>"001001001",
  47321=>"001110000",
  47322=>"000110001",
  47323=>"101000110",
  47324=>"101011001",
  47325=>"110110111",
  47326=>"010011110",
  47327=>"010000010",
  47328=>"110010010",
  47329=>"111011101",
  47330=>"010101110",
  47331=>"010100000",
  47332=>"110101111",
  47333=>"101011001",
  47334=>"000101010",
  47335=>"000010111",
  47336=>"111001000",
  47337=>"110110001",
  47338=>"101000001",
  47339=>"010000110",
  47340=>"011111000",
  47341=>"100100100",
  47342=>"110110011",
  47343=>"011101110",
  47344=>"011011000",
  47345=>"111001100",
  47346=>"000001111",
  47347=>"011100011",
  47348=>"000010001",
  47349=>"101100101",
  47350=>"001010100",
  47351=>"101100011",
  47352=>"011001000",
  47353=>"111000101",
  47354=>"000010011",
  47355=>"010000000",
  47356=>"011010001",
  47357=>"010000110",
  47358=>"111001101",
  47359=>"100001110",
  47360=>"011001111",
  47361=>"110110101",
  47362=>"001010101",
  47363=>"000000111",
  47364=>"100110111",
  47365=>"001110110",
  47366=>"111111110",
  47367=>"011101101",
  47368=>"100101110",
  47369=>"101100010",
  47370=>"110111111",
  47371=>"110110111",
  47372=>"001000010",
  47373=>"100111011",
  47374=>"010111001",
  47375=>"101000100",
  47376=>"110000000",
  47377=>"100011000",
  47378=>"001101111",
  47379=>"010001100",
  47380=>"010011110",
  47381=>"000110011",
  47382=>"101001110",
  47383=>"100110001",
  47384=>"111010001",
  47385=>"000000110",
  47386=>"110100001",
  47387=>"010011011",
  47388=>"000110101",
  47389=>"011101001",
  47390=>"000010001",
  47391=>"001100101",
  47392=>"101001100",
  47393=>"000111010",
  47394=>"010001010",
  47395=>"011001001",
  47396=>"001010011",
  47397=>"110000110",
  47398=>"110101000",
  47399=>"110011110",
  47400=>"101010001",
  47401=>"110100010",
  47402=>"001011100",
  47403=>"111000111",
  47404=>"011001101",
  47405=>"001000111",
  47406=>"000000000",
  47407=>"100110110",
  47408=>"001010011",
  47409=>"010001110",
  47410=>"100110001",
  47411=>"011111011",
  47412=>"001101001",
  47413=>"010001111",
  47414=>"111101010",
  47415=>"000110111",
  47416=>"010010100",
  47417=>"001001001",
  47418=>"111011111",
  47419=>"010100100",
  47420=>"110011010",
  47421=>"010100100",
  47422=>"010011011",
  47423=>"111111010",
  47424=>"100101000",
  47425=>"011001001",
  47426=>"010101100",
  47427=>"100001011",
  47428=>"011000011",
  47429=>"111110101",
  47430=>"100000011",
  47431=>"001101111",
  47432=>"110011110",
  47433=>"010000011",
  47434=>"101001101",
  47435=>"010011000",
  47436=>"110001100",
  47437=>"110100011",
  47438=>"010101001",
  47439=>"001001101",
  47440=>"100001010",
  47441=>"101111000",
  47442=>"000110000",
  47443=>"011001000",
  47444=>"010010100",
  47445=>"110111000",
  47446=>"101100100",
  47447=>"011011110",
  47448=>"011101100",
  47449=>"110100001",
  47450=>"010100111",
  47451=>"001101000",
  47452=>"100111001",
  47453=>"111111011",
  47454=>"000011100",
  47455=>"000000101",
  47456=>"000101101",
  47457=>"111011111",
  47458=>"001110111",
  47459=>"000100010",
  47460=>"110001100",
  47461=>"100001010",
  47462=>"010110011",
  47463=>"001110101",
  47464=>"100011101",
  47465=>"010110010",
  47466=>"111101001",
  47467=>"100010100",
  47468=>"011100000",
  47469=>"010000011",
  47470=>"001001001",
  47471=>"101111101",
  47472=>"010101010",
  47473=>"000001111",
  47474=>"110010001",
  47475=>"100001101",
  47476=>"001001100",
  47477=>"001011100",
  47478=>"101110100",
  47479=>"011000010",
  47480=>"110111100",
  47481=>"100101110",
  47482=>"100010000",
  47483=>"001111011",
  47484=>"101000000",
  47485=>"011011110",
  47486=>"111001011",
  47487=>"110000100",
  47488=>"100100111",
  47489=>"001100000",
  47490=>"110001110",
  47491=>"101001000",
  47492=>"110101001",
  47493=>"110001000",
  47494=>"011010010",
  47495=>"011011100",
  47496=>"100000100",
  47497=>"001111010",
  47498=>"010111100",
  47499=>"000000101",
  47500=>"001110011",
  47501=>"100111111",
  47502=>"010011101",
  47503=>"100000011",
  47504=>"011101001",
  47505=>"010001111",
  47506=>"011001000",
  47507=>"101001011",
  47508=>"001111100",
  47509=>"111000000",
  47510=>"001010100",
  47511=>"101001001",
  47512=>"111110111",
  47513=>"010010100",
  47514=>"010101001",
  47515=>"001101000",
  47516=>"000100110",
  47517=>"010010100",
  47518=>"011110111",
  47519=>"100011101",
  47520=>"011000001",
  47521=>"010111111",
  47522=>"010001111",
  47523=>"111111111",
  47524=>"000011001",
  47525=>"000100100",
  47526=>"011010001",
  47527=>"111010111",
  47528=>"000000001",
  47529=>"000010110",
  47530=>"101101110",
  47531=>"100111011",
  47532=>"110010111",
  47533=>"101001101",
  47534=>"011001100",
  47535=>"001011000",
  47536=>"011010110",
  47537=>"110000011",
  47538=>"000010010",
  47539=>"011001100",
  47540=>"100011111",
  47541=>"011110101",
  47542=>"010100010",
  47543=>"101111001",
  47544=>"110110010",
  47545=>"010000110",
  47546=>"111010101",
  47547=>"010100100",
  47548=>"011001000",
  47549=>"111001000",
  47550=>"111011000",
  47551=>"000001101",
  47552=>"000001000",
  47553=>"000010010",
  47554=>"101010000",
  47555=>"101000110",
  47556=>"100101110",
  47557=>"010111110",
  47558=>"111011000",
  47559=>"010000000",
  47560=>"000111011",
  47561=>"100110111",
  47562=>"100101100",
  47563=>"111001111",
  47564=>"010100000",
  47565=>"000110110",
  47566=>"101001011",
  47567=>"011001110",
  47568=>"111100110",
  47569=>"011011010",
  47570=>"101101101",
  47571=>"011111111",
  47572=>"001010111",
  47573=>"100111010",
  47574=>"100011111",
  47575=>"111011111",
  47576=>"101101011",
  47577=>"011011101",
  47578=>"100111111",
  47579=>"000001111",
  47580=>"101110010",
  47581=>"000110011",
  47582=>"010100001",
  47583=>"101111000",
  47584=>"110111011",
  47585=>"101010110",
  47586=>"011001000",
  47587=>"010100001",
  47588=>"111101010",
  47589=>"001110000",
  47590=>"011101011",
  47591=>"010011101",
  47592=>"101010010",
  47593=>"100101001",
  47594=>"101000000",
  47595=>"101100000",
  47596=>"100110010",
  47597=>"111001010",
  47598=>"110011010",
  47599=>"100011011",
  47600=>"010111000",
  47601=>"111001111",
  47602=>"110110110",
  47603=>"110000010",
  47604=>"001000001",
  47605=>"010100011",
  47606=>"110000010",
  47607=>"111011101",
  47608=>"101000001",
  47609=>"101001100",
  47610=>"011111001",
  47611=>"111110011",
  47612=>"110110111",
  47613=>"111111101",
  47614=>"001101111",
  47615=>"100010101",
  47616=>"000110101",
  47617=>"100101000",
  47618=>"110101111",
  47619=>"001101000",
  47620=>"110100010",
  47621=>"101001110",
  47622=>"011110111",
  47623=>"000000011",
  47624=>"011111000",
  47625=>"001011011",
  47626=>"101111010",
  47627=>"110001011",
  47628=>"000000011",
  47629=>"110000111",
  47630=>"000000000",
  47631=>"011011100",
  47632=>"101011001",
  47633=>"111010100",
  47634=>"111011100",
  47635=>"110101101",
  47636=>"001100100",
  47637=>"110110100",
  47638=>"000011011",
  47639=>"100101001",
  47640=>"100110010",
  47641=>"000001000",
  47642=>"000010001",
  47643=>"010100100",
  47644=>"010011100",
  47645=>"010000100",
  47646=>"011111000",
  47647=>"100111011",
  47648=>"101001011",
  47649=>"000011010",
  47650=>"011000000",
  47651=>"101010101",
  47652=>"010011001",
  47653=>"100000000",
  47654=>"100111111",
  47655=>"101110111",
  47656=>"111010001",
  47657=>"000100001",
  47658=>"110111001",
  47659=>"011001010",
  47660=>"101010100",
  47661=>"111111000",
  47662=>"000101001",
  47663=>"011101000",
  47664=>"011100001",
  47665=>"101110010",
  47666=>"101000001",
  47667=>"100010101",
  47668=>"111000101",
  47669=>"000010101",
  47670=>"011110111",
  47671=>"100100010",
  47672=>"111011110",
  47673=>"011010101",
  47674=>"001000000",
  47675=>"011100011",
  47676=>"101010011",
  47677=>"110110010",
  47678=>"101111100",
  47679=>"010001110",
  47680=>"000111111",
  47681=>"011000001",
  47682=>"110010010",
  47683=>"110010000",
  47684=>"000000111",
  47685=>"010111001",
  47686=>"000100011",
  47687=>"010101000",
  47688=>"101101101",
  47689=>"101010111",
  47690=>"010101000",
  47691=>"100001000",
  47692=>"110111000",
  47693=>"100001000",
  47694=>"000001000",
  47695=>"110110001",
  47696=>"011110110",
  47697=>"100001000",
  47698=>"001010111",
  47699=>"101100111",
  47700=>"110011110",
  47701=>"000110000",
  47702=>"101001111",
  47703=>"001101000",
  47704=>"110100010",
  47705=>"001011000",
  47706=>"111100011",
  47707=>"000001101",
  47708=>"001111010",
  47709=>"010010010",
  47710=>"100001010",
  47711=>"011011100",
  47712=>"000011100",
  47713=>"111000010",
  47714=>"001110001",
  47715=>"010111101",
  47716=>"011100111",
  47717=>"100101000",
  47718=>"001011100",
  47719=>"001100001",
  47720=>"101001010",
  47721=>"100110100",
  47722=>"011111111",
  47723=>"100100101",
  47724=>"001010011",
  47725=>"101001011",
  47726=>"000101110",
  47727=>"000111110",
  47728=>"100100101",
  47729=>"000000100",
  47730=>"110111010",
  47731=>"110011001",
  47732=>"010111000",
  47733=>"100101011",
  47734=>"001110010",
  47735=>"110100110",
  47736=>"000101101",
  47737=>"111111101",
  47738=>"111111011",
  47739=>"001001101",
  47740=>"001010111",
  47741=>"101000111",
  47742=>"100000011",
  47743=>"001011111",
  47744=>"010000001",
  47745=>"111111100",
  47746=>"101001001",
  47747=>"010011001",
  47748=>"100101110",
  47749=>"001010000",
  47750=>"011011011",
  47751=>"001010000",
  47752=>"110000000",
  47753=>"000010000",
  47754=>"110010010",
  47755=>"011110101",
  47756=>"001000100",
  47757=>"010001010",
  47758=>"110100011",
  47759=>"100110010",
  47760=>"010110100",
  47761=>"111010000",
  47762=>"010010001",
  47763=>"101001011",
  47764=>"011101110",
  47765=>"011101011",
  47766=>"010010111",
  47767=>"000111110",
  47768=>"101011000",
  47769=>"111101001",
  47770=>"111001000",
  47771=>"101010011",
  47772=>"110011100",
  47773=>"010010110",
  47774=>"000101110",
  47775=>"110111111",
  47776=>"110111100",
  47777=>"111000101",
  47778=>"010000011",
  47779=>"010100001",
  47780=>"111011010",
  47781=>"110111110",
  47782=>"010001000",
  47783=>"101000000",
  47784=>"110100000",
  47785=>"111011111",
  47786=>"101110000",
  47787=>"101000000",
  47788=>"001000111",
  47789=>"100110010",
  47790=>"100101111",
  47791=>"111110000",
  47792=>"101011111",
  47793=>"010000101",
  47794=>"010001101",
  47795=>"111001011",
  47796=>"111001110",
  47797=>"001010011",
  47798=>"111111010",
  47799=>"000111001",
  47800=>"000011111",
  47801=>"010110101",
  47802=>"101101101",
  47803=>"100001011",
  47804=>"111101000",
  47805=>"011010001",
  47806=>"000001000",
  47807=>"010000100",
  47808=>"010010001",
  47809=>"010000000",
  47810=>"111000000",
  47811=>"011000011",
  47812=>"000010000",
  47813=>"000000100",
  47814=>"101011111",
  47815=>"100111011",
  47816=>"011100010",
  47817=>"111001011",
  47818=>"111111001",
  47819=>"010000111",
  47820=>"001110011",
  47821=>"001101010",
  47822=>"001100001",
  47823=>"011011111",
  47824=>"011001111",
  47825=>"001000100",
  47826=>"010111100",
  47827=>"111001101",
  47828=>"011001000",
  47829=>"001101101",
  47830=>"001111111",
  47831=>"010110110",
  47832=>"100101000",
  47833=>"001101000",
  47834=>"110110111",
  47835=>"101111010",
  47836=>"100001110",
  47837=>"001110111",
  47838=>"010011101",
  47839=>"100001101",
  47840=>"111001111",
  47841=>"110010111",
  47842=>"011010011",
  47843=>"111111011",
  47844=>"011000010",
  47845=>"011010011",
  47846=>"100011111",
  47847=>"110101101",
  47848=>"100011000",
  47849=>"100000000",
  47850=>"000100100",
  47851=>"001000011",
  47852=>"001011010",
  47853=>"000100001",
  47854=>"100011111",
  47855=>"100110010",
  47856=>"110010001",
  47857=>"110100111",
  47858=>"011001101",
  47859=>"010110111",
  47860=>"110101110",
  47861=>"011010001",
  47862=>"101001110",
  47863=>"001010001",
  47864=>"101110110",
  47865=>"111110101",
  47866=>"001100101",
  47867=>"001100001",
  47868=>"011110000",
  47869=>"111001101",
  47870=>"010110101",
  47871=>"010100101",
  47872=>"000110011",
  47873=>"110010011",
  47874=>"000001000",
  47875=>"010000001",
  47876=>"011111001",
  47877=>"110011001",
  47878=>"100100110",
  47879=>"000011001",
  47880=>"111000011",
  47881=>"001010011",
  47882=>"111111000",
  47883=>"101110101",
  47884=>"010111001",
  47885=>"110101101",
  47886=>"001110010",
  47887=>"010001010",
  47888=>"000100011",
  47889=>"010011000",
  47890=>"000011111",
  47891=>"001110110",
  47892=>"110111110",
  47893=>"001001011",
  47894=>"001000001",
  47895=>"000001011",
  47896=>"000001010",
  47897=>"010100001",
  47898=>"000010110",
  47899=>"011111010",
  47900=>"000111110",
  47901=>"100111100",
  47902=>"111100010",
  47903=>"101101010",
  47904=>"011000111",
  47905=>"001000011",
  47906=>"010101101",
  47907=>"101000001",
  47908=>"000101010",
  47909=>"010101001",
  47910=>"100110011",
  47911=>"110010010",
  47912=>"010000001",
  47913=>"100111100",
  47914=>"011111001",
  47915=>"000111010",
  47916=>"000011111",
  47917=>"011011010",
  47918=>"011100011",
  47919=>"000000111",
  47920=>"011110110",
  47921=>"010111110",
  47922=>"010010100",
  47923=>"111111011",
  47924=>"001011000",
  47925=>"100101111",
  47926=>"111001011",
  47927=>"000100111",
  47928=>"010111100",
  47929=>"111110111",
  47930=>"001001000",
  47931=>"111100010",
  47932=>"111110001",
  47933=>"101001011",
  47934=>"111111111",
  47935=>"001001111",
  47936=>"000010101",
  47937=>"010000001",
  47938=>"110100101",
  47939=>"100001001",
  47940=>"000001010",
  47941=>"010010010",
  47942=>"111011001",
  47943=>"010110000",
  47944=>"110110011",
  47945=>"000111011",
  47946=>"101000100",
  47947=>"110001001",
  47948=>"101001100",
  47949=>"101000011",
  47950=>"001001100",
  47951=>"001011100",
  47952=>"101101100",
  47953=>"001010010",
  47954=>"011100000",
  47955=>"011001101",
  47956=>"100100100",
  47957=>"110001010",
  47958=>"001000000",
  47959=>"001000111",
  47960=>"111111011",
  47961=>"001011111",
  47962=>"000110101",
  47963=>"100001011",
  47964=>"101110011",
  47965=>"111111111",
  47966=>"011111010",
  47967=>"000010011",
  47968=>"010010101",
  47969=>"101101100",
  47970=>"001000111",
  47971=>"000100010",
  47972=>"010001000",
  47973=>"110111100",
  47974=>"111111011",
  47975=>"100100011",
  47976=>"101100011",
  47977=>"111011111",
  47978=>"110010101",
  47979=>"101101001",
  47980=>"001001011",
  47981=>"100001010",
  47982=>"000001111",
  47983=>"110110101",
  47984=>"110000011",
  47985=>"010101011",
  47986=>"110101111",
  47987=>"011000000",
  47988=>"000100000",
  47989=>"000101001",
  47990=>"001100110",
  47991=>"101001001",
  47992=>"111111011",
  47993=>"111111110",
  47994=>"000100001",
  47995=>"011000101",
  47996=>"000000100",
  47997=>"111000010",
  47998=>"011000011",
  47999=>"111101000",
  48000=>"000010110",
  48001=>"000110010",
  48002=>"111000000",
  48003=>"001100110",
  48004=>"000010001",
  48005=>"000100011",
  48006=>"101100111",
  48007=>"001100110",
  48008=>"100011100",
  48009=>"101111100",
  48010=>"011100100",
  48011=>"000010101",
  48012=>"000011000",
  48013=>"011000101",
  48014=>"110000011",
  48015=>"100110100",
  48016=>"111110011",
  48017=>"101111101",
  48018=>"111111010",
  48019=>"011101010",
  48020=>"111011101",
  48021=>"111010100",
  48022=>"001110001",
  48023=>"100010111",
  48024=>"110001010",
  48025=>"010001010",
  48026=>"000001101",
  48027=>"000110001",
  48028=>"111010101",
  48029=>"110101111",
  48030=>"011111111",
  48031=>"010111000",
  48032=>"111001101",
  48033=>"001101101",
  48034=>"111001010",
  48035=>"001100101",
  48036=>"000011010",
  48037=>"110110100",
  48038=>"010000101",
  48039=>"010001011",
  48040=>"000000101",
  48041=>"001010111",
  48042=>"011101000",
  48043=>"111010100",
  48044=>"001100101",
  48045=>"001000010",
  48046=>"111110000",
  48047=>"000000101",
  48048=>"100100000",
  48049=>"010110111",
  48050=>"100100001",
  48051=>"000101110",
  48052=>"001011000",
  48053=>"111101000",
  48054=>"110010111",
  48055=>"011111000",
  48056=>"011011000",
  48057=>"001010000",
  48058=>"110101110",
  48059=>"010010101",
  48060=>"101000111",
  48061=>"001101100",
  48062=>"111101101",
  48063=>"101010011",
  48064=>"001010111",
  48065=>"111100110",
  48066=>"000100110",
  48067=>"100101111",
  48068=>"111100000",
  48069=>"010011111",
  48070=>"101001000",
  48071=>"011110111",
  48072=>"111000000",
  48073=>"010011101",
  48074=>"100011001",
  48075=>"000000010",
  48076=>"101001100",
  48077=>"001011000",
  48078=>"101010111",
  48079=>"010110000",
  48080=>"101011100",
  48081=>"100000010",
  48082=>"011111000",
  48083=>"011100011",
  48084=>"001100000",
  48085=>"100010110",
  48086=>"110001010",
  48087=>"011110011",
  48088=>"011110010",
  48089=>"010101110",
  48090=>"110111100",
  48091=>"001101101",
  48092=>"100010001",
  48093=>"000011010",
  48094=>"011110000",
  48095=>"001101001",
  48096=>"010010010",
  48097=>"000101011",
  48098=>"101001000",
  48099=>"100101110",
  48100=>"010010001",
  48101=>"001000110",
  48102=>"110111000",
  48103=>"001000100",
  48104=>"100001100",
  48105=>"101001110",
  48106=>"000001110",
  48107=>"011011110",
  48108=>"111000010",
  48109=>"001010110",
  48110=>"111110000",
  48111=>"001010011",
  48112=>"001010011",
  48113=>"001000010",
  48114=>"101111000",
  48115=>"101101010",
  48116=>"010001101",
  48117=>"011000010",
  48118=>"100000111",
  48119=>"000110110",
  48120=>"011010101",
  48121=>"001010101",
  48122=>"100111100",
  48123=>"000111110",
  48124=>"100110010",
  48125=>"100000011",
  48126=>"010010001",
  48127=>"010001101",
  48128=>"011011111",
  48129=>"110110101",
  48130=>"110111110",
  48131=>"010101010",
  48132=>"001111000",
  48133=>"101000011",
  48134=>"011010011",
  48135=>"001000100",
  48136=>"000101101",
  48137=>"100011011",
  48138=>"110010000",
  48139=>"011000000",
  48140=>"111100011",
  48141=>"000110110",
  48142=>"010110001",
  48143=>"001110101",
  48144=>"010000010",
  48145=>"110111001",
  48146=>"110011111",
  48147=>"010100000",
  48148=>"100101001",
  48149=>"100101111",
  48150=>"000010001",
  48151=>"001101101",
  48152=>"101000111",
  48153=>"010010111",
  48154=>"010111110",
  48155=>"100001010",
  48156=>"010001011",
  48157=>"101100111",
  48158=>"100101011",
  48159=>"000001111",
  48160=>"110101001",
  48161=>"000001001",
  48162=>"011111000",
  48163=>"001011110",
  48164=>"101001100",
  48165=>"000011001",
  48166=>"100000011",
  48167=>"101011110",
  48168=>"111111001",
  48169=>"011001001",
  48170=>"011110111",
  48171=>"100101100",
  48172=>"111110111",
  48173=>"010101000",
  48174=>"010001001",
  48175=>"010111100",
  48176=>"100000010",
  48177=>"001101100",
  48178=>"010011011",
  48179=>"001101100",
  48180=>"010010001",
  48181=>"101110010",
  48182=>"111111011",
  48183=>"110011001",
  48184=>"000101100",
  48185=>"010011100",
  48186=>"000101001",
  48187=>"110111011",
  48188=>"011000011",
  48189=>"010010011",
  48190=>"110111011",
  48191=>"111011110",
  48192=>"101000010",
  48193=>"100000101",
  48194=>"000000101",
  48195=>"001011010",
  48196=>"100000110",
  48197=>"001010100",
  48198=>"110101111",
  48199=>"010111101",
  48200=>"111010000",
  48201=>"011010111",
  48202=>"100010001",
  48203=>"001000000",
  48204=>"100011011",
  48205=>"110000001",
  48206=>"110010010",
  48207=>"111011110",
  48208=>"001110101",
  48209=>"111111101",
  48210=>"000001001",
  48211=>"110101100",
  48212=>"010001000",
  48213=>"101001011",
  48214=>"100111000",
  48215=>"110010010",
  48216=>"010111011",
  48217=>"000010011",
  48218=>"001001001",
  48219=>"000100101",
  48220=>"000110100",
  48221=>"100100100",
  48222=>"111011010",
  48223=>"010011001",
  48224=>"111010010",
  48225=>"001110101",
  48226=>"111110001",
  48227=>"001001111",
  48228=>"111000110",
  48229=>"110101000",
  48230=>"000001000",
  48231=>"101101001",
  48232=>"001000110",
  48233=>"010100000",
  48234=>"000001011",
  48235=>"100010100",
  48236=>"110111010",
  48237=>"110100010",
  48238=>"001011010",
  48239=>"111101100",
  48240=>"100010110",
  48241=>"111011111",
  48242=>"101110110",
  48243=>"011001011",
  48244=>"100100111",
  48245=>"111000111",
  48246=>"000000110",
  48247=>"111001111",
  48248=>"110100111",
  48249=>"000010111",
  48250=>"111000010",
  48251=>"100011001",
  48252=>"111001010",
  48253=>"100001010",
  48254=>"011101111",
  48255=>"100111100",
  48256=>"101010000",
  48257=>"101101111",
  48258=>"010001010",
  48259=>"010001010",
  48260=>"111111011",
  48261=>"111101100",
  48262=>"001000111",
  48263=>"011111001",
  48264=>"011000100",
  48265=>"100001111",
  48266=>"010011111",
  48267=>"101010100",
  48268=>"000010101",
  48269=>"010101000",
  48270=>"101010001",
  48271=>"101101101",
  48272=>"010110111",
  48273=>"011110100",
  48274=>"111001111",
  48275=>"110011101",
  48276=>"000100100",
  48277=>"010000111",
  48278=>"010010000",
  48279=>"011010000",
  48280=>"001111010",
  48281=>"001100000",
  48282=>"010110101",
  48283=>"010111100",
  48284=>"001010100",
  48285=>"011001000",
  48286=>"100111011",
  48287=>"001000000",
  48288=>"001100110",
  48289=>"100010101",
  48290=>"110010011",
  48291=>"100100001",
  48292=>"111011001",
  48293=>"110001010",
  48294=>"100010011",
  48295=>"110011111",
  48296=>"010010011",
  48297=>"000110000",
  48298=>"111101010",
  48299=>"001101000",
  48300=>"110011111",
  48301=>"001000111",
  48302=>"000101101",
  48303=>"010101011",
  48304=>"101001001",
  48305=>"001001000",
  48306=>"111110101",
  48307=>"100000101",
  48308=>"110100010",
  48309=>"111101101",
  48310=>"111000110",
  48311=>"010001111",
  48312=>"010010000",
  48313=>"001101001",
  48314=>"101011011",
  48315=>"111100000",
  48316=>"011110010",
  48317=>"111111011",
  48318=>"101011100",
  48319=>"011111111",
  48320=>"110011111",
  48321=>"101000011",
  48322=>"101111111",
  48323=>"000100101",
  48324=>"010000110",
  48325=>"010001000",
  48326=>"010011011",
  48327=>"111001100",
  48328=>"000101101",
  48329=>"111001101",
  48330=>"010110110",
  48331=>"011101100",
  48332=>"010000010",
  48333=>"010100111",
  48334=>"011110001",
  48335=>"101111000",
  48336=>"111111101",
  48337=>"101001111",
  48338=>"001101101",
  48339=>"111100011",
  48340=>"001101010",
  48341=>"011110010",
  48342=>"001001011",
  48343=>"000101001",
  48344=>"100101010",
  48345=>"010111100",
  48346=>"000101001",
  48347=>"111000110",
  48348=>"110110010",
  48349=>"101011111",
  48350=>"011111101",
  48351=>"101010010",
  48352=>"111111011",
  48353=>"110111111",
  48354=>"001000001",
  48355=>"110100010",
  48356=>"011111001",
  48357=>"010100100",
  48358=>"111001101",
  48359=>"111001001",
  48360=>"000100010",
  48361=>"010110001",
  48362=>"111111101",
  48363=>"001001000",
  48364=>"011010110",
  48365=>"111110100",
  48366=>"000101110",
  48367=>"110111101",
  48368=>"000000110",
  48369=>"000001000",
  48370=>"101001010",
  48371=>"001000110",
  48372=>"011000110",
  48373=>"100110100",
  48374=>"000110101",
  48375=>"111101101",
  48376=>"101011111",
  48377=>"101010000",
  48378=>"010101011",
  48379=>"011100110",
  48380=>"001000001",
  48381=>"000111011",
  48382=>"111000111",
  48383=>"011011100",
  48384=>"000111001",
  48385=>"110100010",
  48386=>"100111011",
  48387=>"011010111",
  48388=>"010000000",
  48389=>"110001010",
  48390=>"011100101",
  48391=>"111110110",
  48392=>"000011010",
  48393=>"101101111",
  48394=>"110011100",
  48395=>"111011011",
  48396=>"011001001",
  48397=>"000111100",
  48398=>"101011010",
  48399=>"011110010",
  48400=>"001101011",
  48401=>"010110101",
  48402=>"111111111",
  48403=>"000101011",
  48404=>"101101110",
  48405=>"001110111",
  48406=>"010001111",
  48407=>"011111111",
  48408=>"101100011",
  48409=>"001011111",
  48410=>"111010000",
  48411=>"111110001",
  48412=>"000011101",
  48413=>"011000011",
  48414=>"111100101",
  48415=>"010000100",
  48416=>"110101000",
  48417=>"011010101",
  48418=>"001001001",
  48419=>"011101101",
  48420=>"100111110",
  48421=>"010110101",
  48422=>"001101111",
  48423=>"010011001",
  48424=>"000001111",
  48425=>"111111111",
  48426=>"001110011",
  48427=>"110010100",
  48428=>"110011001",
  48429=>"100010001",
  48430=>"000000001",
  48431=>"000110100",
  48432=>"000001010",
  48433=>"111001101",
  48434=>"111101011",
  48435=>"000101001",
  48436=>"100001100",
  48437=>"100000000",
  48438=>"111000110",
  48439=>"110101111",
  48440=>"110001011",
  48441=>"000011001",
  48442=>"111100010",
  48443=>"010011110",
  48444=>"100110110",
  48445=>"000111110",
  48446=>"001011110",
  48447=>"011001000",
  48448=>"100001100",
  48449=>"110010100",
  48450=>"111101101",
  48451=>"110100011",
  48452=>"111111111",
  48453=>"110101111",
  48454=>"110000010",
  48455=>"000110101",
  48456=>"010000110",
  48457=>"000011101",
  48458=>"011111011",
  48459=>"010001000",
  48460=>"100011111",
  48461=>"000011001",
  48462=>"000001011",
  48463=>"000100110",
  48464=>"010011000",
  48465=>"100100111",
  48466=>"110010000",
  48467=>"100100000",
  48468=>"110111000",
  48469=>"111111111",
  48470=>"011011110",
  48471=>"001110010",
  48472=>"100010000",
  48473=>"101001011",
  48474=>"010010100",
  48475=>"000000010",
  48476=>"110111100",
  48477=>"100001110",
  48478=>"011010101",
  48479=>"111100100",
  48480=>"110100110",
  48481=>"100001011",
  48482=>"011000011",
  48483=>"110010000",
  48484=>"100011000",
  48485=>"000111110",
  48486=>"100111011",
  48487=>"111010100",
  48488=>"000001000",
  48489=>"010011101",
  48490=>"000110110",
  48491=>"100111111",
  48492=>"001100011",
  48493=>"010100101",
  48494=>"000000011",
  48495=>"111101000",
  48496=>"111111111",
  48497=>"101110011",
  48498=>"101001000",
  48499=>"011010100",
  48500=>"101100110",
  48501=>"100100010",
  48502=>"011010100",
  48503=>"011000111",
  48504=>"001000110",
  48505=>"101001011",
  48506=>"011111000",
  48507=>"111100000",
  48508=>"011110111",
  48509=>"111000010",
  48510=>"111100100",
  48511=>"110110101",
  48512=>"111110000",
  48513=>"101111010",
  48514=>"010001100",
  48515=>"000100110",
  48516=>"110000000",
  48517=>"100101010",
  48518=>"110011111",
  48519=>"000000001",
  48520=>"110010010",
  48521=>"010001101",
  48522=>"101100010",
  48523=>"101101101",
  48524=>"000001111",
  48525=>"100100011",
  48526=>"001100101",
  48527=>"000010000",
  48528=>"010100101",
  48529=>"000111000",
  48530=>"000010111",
  48531=>"011001001",
  48532=>"100001101",
  48533=>"100000110",
  48534=>"101111110",
  48535=>"010000010",
  48536=>"001000100",
  48537=>"011011101",
  48538=>"100110111",
  48539=>"111111000",
  48540=>"011011111",
  48541=>"111011101",
  48542=>"101101111",
  48543=>"101010110",
  48544=>"110100111",
  48545=>"111001010",
  48546=>"111010111",
  48547=>"110000001",
  48548=>"001110101",
  48549=>"010000000",
  48550=>"101001100",
  48551=>"001001100",
  48552=>"111001111",
  48553=>"100010100",
  48554=>"000100010",
  48555=>"010110010",
  48556=>"110000100",
  48557=>"111000001",
  48558=>"110110011",
  48559=>"011011000",
  48560=>"101001101",
  48561=>"100101001",
  48562=>"110000010",
  48563=>"110100001",
  48564=>"011010001",
  48565=>"001010001",
  48566=>"110101001",
  48567=>"111101101",
  48568=>"001110110",
  48569=>"100011111",
  48570=>"010010000",
  48571=>"101001001",
  48572=>"000000000",
  48573=>"001010100",
  48574=>"000101010",
  48575=>"000100100",
  48576=>"110010010",
  48577=>"101110111",
  48578=>"110110011",
  48579=>"110011010",
  48580=>"111001101",
  48581=>"011100110",
  48582=>"011110010",
  48583=>"101010101",
  48584=>"000000111",
  48585=>"100000100",
  48586=>"111010110",
  48587=>"010000000",
  48588=>"101000100",
  48589=>"011010000",
  48590=>"111110101",
  48591=>"000000010",
  48592=>"010110110",
  48593=>"010001001",
  48594=>"101101111",
  48595=>"111101001",
  48596=>"010110101",
  48597=>"110100010",
  48598=>"100001100",
  48599=>"000010100",
  48600=>"000111111",
  48601=>"101000000",
  48602=>"101111101",
  48603=>"110110001",
  48604=>"101001010",
  48605=>"000110001",
  48606=>"111111100",
  48607=>"001000011",
  48608=>"110000111",
  48609=>"111111110",
  48610=>"011010000",
  48611=>"000000111",
  48612=>"000010000",
  48613=>"111010111",
  48614=>"111011111",
  48615=>"000011010",
  48616=>"111111111",
  48617=>"011010111",
  48618=>"000011110",
  48619=>"010101011",
  48620=>"110000001",
  48621=>"101110010",
  48622=>"000000001",
  48623=>"111111001",
  48624=>"000000000",
  48625=>"000100010",
  48626=>"000101000",
  48627=>"111001011",
  48628=>"111011111",
  48629=>"101101100",
  48630=>"110000100",
  48631=>"001100010",
  48632=>"100101111",
  48633=>"000001100",
  48634=>"000000111",
  48635=>"100101101",
  48636=>"000011100",
  48637=>"100101101",
  48638=>"011111010",
  48639=>"010111010",
  48640=>"000010111",
  48641=>"001011100",
  48642=>"110111110",
  48643=>"111101001",
  48644=>"010101000",
  48645=>"101010010",
  48646=>"011001001",
  48647=>"011111100",
  48648=>"000110010",
  48649=>"100101010",
  48650=>"111110010",
  48651=>"000001100",
  48652=>"100000111",
  48653=>"000101001",
  48654=>"111101011",
  48655=>"100101001",
  48656=>"111100010",
  48657=>"001111000",
  48658=>"011101101",
  48659=>"100110011",
  48660=>"010111101",
  48661=>"110101111",
  48662=>"100010110",
  48663=>"101111110",
  48664=>"101001111",
  48665=>"010110100",
  48666=>"011010001",
  48667=>"100001001",
  48668=>"111010110",
  48669=>"000010110",
  48670=>"010011011",
  48671=>"000010001",
  48672=>"001000110",
  48673=>"100110011",
  48674=>"001001000",
  48675=>"110000111",
  48676=>"011001100",
  48677=>"110111110",
  48678=>"100110110",
  48679=>"011000001",
  48680=>"100111111",
  48681=>"110111100",
  48682=>"000000010",
  48683=>"101101101",
  48684=>"011100001",
  48685=>"110000010",
  48686=>"111100000",
  48687=>"111010111",
  48688=>"011011011",
  48689=>"010100101",
  48690=>"001000010",
  48691=>"011010001",
  48692=>"000100010",
  48693=>"000101110",
  48694=>"111110010",
  48695=>"101100001",
  48696=>"001100000",
  48697=>"001001110",
  48698=>"001101010",
  48699=>"110000011",
  48700=>"111100000",
  48701=>"101111100",
  48702=>"111101110",
  48703=>"000110110",
  48704=>"101000101",
  48705=>"101101010",
  48706=>"011100110",
  48707=>"110110111",
  48708=>"100001011",
  48709=>"001000010",
  48710=>"000011111",
  48711=>"010010000",
  48712=>"010110101",
  48713=>"101100110",
  48714=>"000111111",
  48715=>"011101001",
  48716=>"111111111",
  48717=>"001111111",
  48718=>"100000000",
  48719=>"100001011",
  48720=>"100111001",
  48721=>"000111110",
  48722=>"100001000",
  48723=>"011110001",
  48724=>"110101110",
  48725=>"010010111",
  48726=>"000000001",
  48727=>"000001111",
  48728=>"011111001",
  48729=>"110000001",
  48730=>"110000111",
  48731=>"000001001",
  48732=>"000110100",
  48733=>"111001011",
  48734=>"101001110",
  48735=>"100100110",
  48736=>"011100000",
  48737=>"001110011",
  48738=>"001001010",
  48739=>"010111000",
  48740=>"001000010",
  48741=>"000001101",
  48742=>"101010010",
  48743=>"000001000",
  48744=>"001111110",
  48745=>"100101000",
  48746=>"000110100",
  48747=>"101110101",
  48748=>"000110101",
  48749=>"100111111",
  48750=>"010001111",
  48751=>"110000010",
  48752=>"010011010",
  48753=>"010110000",
  48754=>"010011001",
  48755=>"101110111",
  48756=>"001100011",
  48757=>"000101111",
  48758=>"000010110",
  48759=>"111110111",
  48760=>"100010101",
  48761=>"111000000",
  48762=>"011000001",
  48763=>"010101000",
  48764=>"010100100",
  48765=>"010000011",
  48766=>"100111110",
  48767=>"110010110",
  48768=>"001000000",
  48769=>"000011011",
  48770=>"111001011",
  48771=>"000011011",
  48772=>"000100010",
  48773=>"101010000",
  48774=>"101011100",
  48775=>"111011010",
  48776=>"101101001",
  48777=>"110100110",
  48778=>"101111011",
  48779=>"101010000",
  48780=>"110101110",
  48781=>"010110000",
  48782=>"111110111",
  48783=>"111111011",
  48784=>"010110100",
  48785=>"000000000",
  48786=>"101001001",
  48787=>"100011101",
  48788=>"000000101",
  48789=>"000011001",
  48790=>"000111000",
  48791=>"011100011",
  48792=>"001010001",
  48793=>"100110000",
  48794=>"001110111",
  48795=>"010101000",
  48796=>"101011000",
  48797=>"100011100",
  48798=>"101011011",
  48799=>"110110110",
  48800=>"001010110",
  48801=>"100001111",
  48802=>"000001001",
  48803=>"110110010",
  48804=>"010011111",
  48805=>"011001000",
  48806=>"000111000",
  48807=>"000111111",
  48808=>"001010111",
  48809=>"101000000",
  48810=>"011100001",
  48811=>"001011010",
  48812=>"010111111",
  48813=>"000001001",
  48814=>"000001010",
  48815=>"011001100",
  48816=>"111110001",
  48817=>"011010110",
  48818=>"000100110",
  48819=>"010001001",
  48820=>"000011011",
  48821=>"001011100",
  48822=>"110001011",
  48823=>"010001000",
  48824=>"100001110",
  48825=>"011111111",
  48826=>"010011001",
  48827=>"110000001",
  48828=>"101111101",
  48829=>"010001001",
  48830=>"011001001",
  48831=>"001001000",
  48832=>"101110101",
  48833=>"100101000",
  48834=>"010101100",
  48835=>"111111000",
  48836=>"101000101",
  48837=>"010100010",
  48838=>"101100010",
  48839=>"000100000",
  48840=>"111101100",
  48841=>"011001111",
  48842=>"000001000",
  48843=>"010101110",
  48844=>"111110100",
  48845=>"001101010",
  48846=>"010000101",
  48847=>"011110111",
  48848=>"110110111",
  48849=>"100101010",
  48850=>"000110001",
  48851=>"010001010",
  48852=>"000111000",
  48853=>"101011001",
  48854=>"011010101",
  48855=>"110010110",
  48856=>"000100010",
  48857=>"101010100",
  48858=>"100111000",
  48859=>"000010011",
  48860=>"101110001",
  48861=>"110000100",
  48862=>"000111000",
  48863=>"010000010",
  48864=>"010010010",
  48865=>"000111101",
  48866=>"000011011",
  48867=>"010010010",
  48868=>"010100001",
  48869=>"000100001",
  48870=>"111100000",
  48871=>"010100100",
  48872=>"011010010",
  48873=>"111010010",
  48874=>"011111000",
  48875=>"011101000",
  48876=>"110110111",
  48877=>"011010100",
  48878=>"000000101",
  48879=>"010111100",
  48880=>"101101111",
  48881=>"110100001",
  48882=>"101011101",
  48883=>"110100101",
  48884=>"111100000",
  48885=>"000000111",
  48886=>"000001111",
  48887=>"111111011",
  48888=>"011100001",
  48889=>"001000111",
  48890=>"000010011",
  48891=>"111011001",
  48892=>"101000011",
  48893=>"100000010",
  48894=>"101010110",
  48895=>"110000011",
  48896=>"010110111",
  48897=>"001111111",
  48898=>"111100101",
  48899=>"000000011",
  48900=>"111101010",
  48901=>"111001101",
  48902=>"010000110",
  48903=>"101101001",
  48904=>"010000001",
  48905=>"101001101",
  48906=>"100111111",
  48907=>"100011111",
  48908=>"000110111",
  48909=>"100110110",
  48910=>"111000111",
  48911=>"001011001",
  48912=>"100011000",
  48913=>"000011000",
  48914=>"011000010",
  48915=>"011101001",
  48916=>"111100010",
  48917=>"010000011",
  48918=>"110010111",
  48919=>"110011001",
  48920=>"001011011",
  48921=>"000110011",
  48922=>"011001000",
  48923=>"011000001",
  48924=>"000000110",
  48925=>"011001011",
  48926=>"100100100",
  48927=>"000100001",
  48928=>"110101110",
  48929=>"011011000",
  48930=>"100111010",
  48931=>"110000000",
  48932=>"100010111",
  48933=>"111110011",
  48934=>"110100001",
  48935=>"111011010",
  48936=>"011011100",
  48937=>"001001101",
  48938=>"110001001",
  48939=>"110101000",
  48940=>"000001100",
  48941=>"000001000",
  48942=>"011100010",
  48943=>"000000001",
  48944=>"000001111",
  48945=>"110001001",
  48946=>"001110001",
  48947=>"000011100",
  48948=>"101111000",
  48949=>"110101111",
  48950=>"111100110",
  48951=>"000110111",
  48952=>"011011100",
  48953=>"111011000",
  48954=>"000011100",
  48955=>"000101011",
  48956=>"001001011",
  48957=>"000010001",
  48958=>"000010001",
  48959=>"010111000",
  48960=>"001110100",
  48961=>"111111011",
  48962=>"111111111",
  48963=>"111111011",
  48964=>"001110010",
  48965=>"010111101",
  48966=>"101110000",
  48967=>"101111001",
  48968=>"000110110",
  48969=>"101100001",
  48970=>"010110001",
  48971=>"100111100",
  48972=>"011010000",
  48973=>"011111000",
  48974=>"001001110",
  48975=>"010110000",
  48976=>"101001000",
  48977=>"110010100",
  48978=>"010000110",
  48979=>"101000101",
  48980=>"000001000",
  48981=>"010010000",
  48982=>"100001001",
  48983=>"110100000",
  48984=>"101000100",
  48985=>"000101010",
  48986=>"100100110",
  48987=>"010111010",
  48988=>"110110011",
  48989=>"010001001",
  48990=>"100010001",
  48991=>"101100110",
  48992=>"001101010",
  48993=>"001011111",
  48994=>"011000001",
  48995=>"000101011",
  48996=>"100000100",
  48997=>"000100011",
  48998=>"110110101",
  48999=>"011010010",
  49000=>"110011011",
  49001=>"101100110",
  49002=>"101011100",
  49003=>"010001001",
  49004=>"000000000",
  49005=>"110010100",
  49006=>"001111101",
  49007=>"110111011",
  49008=>"011101111",
  49009=>"001110111",
  49010=>"000011011",
  49011=>"010101100",
  49012=>"001010000",
  49013=>"001001001",
  49014=>"011000100",
  49015=>"101011000",
  49016=>"101110010",
  49017=>"100000111",
  49018=>"110011111",
  49019=>"011110101",
  49020=>"000000001",
  49021=>"010101000",
  49022=>"110010101",
  49023=>"111111111",
  49024=>"010101111",
  49025=>"101011000",
  49026=>"001100001",
  49027=>"001011000",
  49028=>"100001011",
  49029=>"010001001",
  49030=>"111101101",
  49031=>"001100011",
  49032=>"111001110",
  49033=>"010110010",
  49034=>"010011000",
  49035=>"111011001",
  49036=>"100100000",
  49037=>"011001110",
  49038=>"101100001",
  49039=>"001001100",
  49040=>"100111111",
  49041=>"100001010",
  49042=>"001111111",
  49043=>"101100001",
  49044=>"110111011",
  49045=>"011010001",
  49046=>"011001010",
  49047=>"010111110",
  49048=>"010111111",
  49049=>"111111000",
  49050=>"010101011",
  49051=>"010000110",
  49052=>"000000010",
  49053=>"000100110",
  49054=>"100111011",
  49055=>"011110100",
  49056=>"010110011",
  49057=>"000110000",
  49058=>"110101111",
  49059=>"011010110",
  49060=>"001000010",
  49061=>"110001001",
  49062=>"101100110",
  49063=>"011011010",
  49064=>"101000001",
  49065=>"000000110",
  49066=>"000001011",
  49067=>"111011010",
  49068=>"100100011",
  49069=>"110111111",
  49070=>"110010101",
  49071=>"111110001",
  49072=>"100111111",
  49073=>"110000101",
  49074=>"100111110",
  49075=>"000110001",
  49076=>"011111101",
  49077=>"111101001",
  49078=>"101100011",
  49079=>"000001010",
  49080=>"100000100",
  49081=>"110110100",
  49082=>"100100100",
  49083=>"100010001",
  49084=>"101101010",
  49085=>"111110100",
  49086=>"111000100",
  49087=>"110100000",
  49088=>"000110001",
  49089=>"010101011",
  49090=>"110111000",
  49091=>"000100000",
  49092=>"001111000",
  49093=>"101101110",
  49094=>"100011010",
  49095=>"111101000",
  49096=>"100110010",
  49097=>"100100010",
  49098=>"111011001",
  49099=>"001100110",
  49100=>"101011011",
  49101=>"111111111",
  49102=>"000010000",
  49103=>"010000000",
  49104=>"111101001",
  49105=>"111000111",
  49106=>"111001110",
  49107=>"001110111",
  49108=>"001111101",
  49109=>"111110000",
  49110=>"011001111",
  49111=>"000101111",
  49112=>"001000001",
  49113=>"101101100",
  49114=>"000000000",
  49115=>"011110010",
  49116=>"101011110",
  49117=>"010101100",
  49118=>"000000000",
  49119=>"010100110",
  49120=>"111111010",
  49121=>"010111100",
  49122=>"011001011",
  49123=>"011100110",
  49124=>"101000101",
  49125=>"000001101",
  49126=>"111100010",
  49127=>"100110000",
  49128=>"101100000",
  49129=>"000111111",
  49130=>"101010000",
  49131=>"011100000",
  49132=>"011000001",
  49133=>"011001100",
  49134=>"010111011",
  49135=>"011100011",
  49136=>"011111011",
  49137=>"011111111",
  49138=>"010100001",
  49139=>"100010100",
  49140=>"000011101",
  49141=>"110010100",
  49142=>"011101010",
  49143=>"110101100",
  49144=>"100110001",
  49145=>"010000011",
  49146=>"001001001",
  49147=>"100110010",
  49148=>"010011101",
  49149=>"011000101",
  49150=>"100110111",
  49151=>"011000001",
  49152=>"010001001",
  49153=>"000010000",
  49154=>"011001101",
  49155=>"110111001",
  49156=>"110111011",
  49157=>"011101111",
  49158=>"000001011",
  49159=>"101110010",
  49160=>"110000110",
  49161=>"101010010",
  49162=>"100010010",
  49163=>"010010010",
  49164=>"010101110",
  49165=>"111111011",
  49166=>"001001010",
  49167=>"011111100",
  49168=>"111111100",
  49169=>"010000011",
  49170=>"101111100",
  49171=>"101101110",
  49172=>"001010100",
  49173=>"100000000",
  49174=>"010110100",
  49175=>"011110111",
  49176=>"000001011",
  49177=>"101101000",
  49178=>"011001111",
  49179=>"110111110",
  49180=>"101111010",
  49181=>"011111110",
  49182=>"010011001",
  49183=>"001011101",
  49184=>"110011011",
  49185=>"101111110",
  49186=>"101001101",
  49187=>"100011111",
  49188=>"010011111",
  49189=>"010000111",
  49190=>"111001111",
  49191=>"011001000",
  49192=>"011101101",
  49193=>"001110101",
  49194=>"111001000",
  49195=>"110100110",
  49196=>"000000000",
  49197=>"010000110",
  49198=>"111100100",
  49199=>"110001011",
  49200=>"100001110",
  49201=>"100010011",
  49202=>"000101000",
  49203=>"111111110",
  49204=>"101000010",
  49205=>"111011010",
  49206=>"111010001",
  49207=>"001011110",
  49208=>"101110000",
  49209=>"111101010",
  49210=>"001001111",
  49211=>"100011111",
  49212=>"001010010",
  49213=>"010000011",
  49214=>"110001011",
  49215=>"100001101",
  49216=>"010110000",
  49217=>"000001100",
  49218=>"001111000",
  49219=>"101000100",
  49220=>"001110001",
  49221=>"111000001",
  49222=>"100000110",
  49223=>"011111001",
  49224=>"010110111",
  49225=>"110111010",
  49226=>"010101001",
  49227=>"010011010",
  49228=>"011110010",
  49229=>"011011011",
  49230=>"010111101",
  49231=>"101110000",
  49232=>"111110110",
  49233=>"101101101",
  49234=>"101111000",
  49235=>"111110011",
  49236=>"101100110",
  49237=>"001101010",
  49238=>"011000010",
  49239=>"001010011",
  49240=>"101111110",
  49241=>"011001011",
  49242=>"111111110",
  49243=>"001100000",
  49244=>"011010000",
  49245=>"000000101",
  49246=>"010110110",
  49247=>"010000110",
  49248=>"010011000",
  49249=>"110001101",
  49250=>"000001111",
  49251=>"100010000",
  49252=>"100011010",
  49253=>"010111011",
  49254=>"111100110",
  49255=>"000001000",
  49256=>"000101001",
  49257=>"111110001",
  49258=>"001001111",
  49259=>"001111000",
  49260=>"000110011",
  49261=>"110000111",
  49262=>"000110101",
  49263=>"000100110",
  49264=>"101001101",
  49265=>"100001100",
  49266=>"110100111",
  49267=>"000001111",
  49268=>"100110000",
  49269=>"111110011",
  49270=>"110011100",
  49271=>"111010000",
  49272=>"101101100",
  49273=>"000111010",
  49274=>"011010001",
  49275=>"010001101",
  49276=>"011110111",
  49277=>"110011001",
  49278=>"000001001",
  49279=>"001110100",
  49280=>"101011101",
  49281=>"101110111",
  49282=>"000000000",
  49283=>"010101111",
  49284=>"111111110",
  49285=>"110000000",
  49286=>"110100001",
  49287=>"101011011",
  49288=>"000000000",
  49289=>"101000110",
  49290=>"111111101",
  49291=>"000101111",
  49292=>"010101100",
  49293=>"100100001",
  49294=>"010110011",
  49295=>"001100101",
  49296=>"010110001",
  49297=>"011010000",
  49298=>"001000001",
  49299=>"101011010",
  49300=>"110001000",
  49301=>"001100010",
  49302=>"011110111",
  49303=>"000110000",
  49304=>"000011000",
  49305=>"001111110",
  49306=>"110110110",
  49307=>"011011100",
  49308=>"100111101",
  49309=>"010101111",
  49310=>"110001011",
  49311=>"010101001",
  49312=>"011101111",
  49313=>"101011110",
  49314=>"111010100",
  49315=>"110010000",
  49316=>"101110101",
  49317=>"111100010",
  49318=>"001100000",
  49319=>"010101101",
  49320=>"111101111",
  49321=>"000000010",
  49322=>"001110001",
  49323=>"101010001",
  49324=>"001101110",
  49325=>"110100101",
  49326=>"100101110",
  49327=>"011011110",
  49328=>"101001010",
  49329=>"000101111",
  49330=>"000010010",
  49331=>"000000001",
  49332=>"010101001",
  49333=>"101100011",
  49334=>"100101001",
  49335=>"010011000",
  49336=>"010010111",
  49337=>"010010001",
  49338=>"010001101",
  49339=>"010010111",
  49340=>"010100000",
  49341=>"111100100",
  49342=>"111100011",
  49343=>"101011111",
  49344=>"010011110",
  49345=>"100000100",
  49346=>"011000101",
  49347=>"100001101",
  49348=>"000011100",
  49349=>"000001100",
  49350=>"110111101",
  49351=>"010000010",
  49352=>"010010011",
  49353=>"011111000",
  49354=>"100011011",
  49355=>"001100010",
  49356=>"100010101",
  49357=>"001110100",
  49358=>"010001010",
  49359=>"011001100",
  49360=>"101010001",
  49361=>"110011011",
  49362=>"111001100",
  49363=>"011010101",
  49364=>"110100101",
  49365=>"011011111",
  49366=>"000011001",
  49367=>"011010001",
  49368=>"101010100",
  49369=>"101100110",
  49370=>"010101101",
  49371=>"110000011",
  49372=>"110101011",
  49373=>"001110111",
  49374=>"101000011",
  49375=>"111000100",
  49376=>"010011000",
  49377=>"011001110",
  49378=>"001001010",
  49379=>"001111000",
  49380=>"100110101",
  49381=>"011110010",
  49382=>"111000000",
  49383=>"111100100",
  49384=>"110100010",
  49385=>"110110100",
  49386=>"001110110",
  49387=>"100100100",
  49388=>"100110110",
  49389=>"100001111",
  49390=>"100101010",
  49391=>"111011001",
  49392=>"010011111",
  49393=>"011000100",
  49394=>"010101010",
  49395=>"011010000",
  49396=>"111100101",
  49397=>"110001010",
  49398=>"101000000",
  49399=>"110110100",
  49400=>"101001001",
  49401=>"001111001",
  49402=>"110011011",
  49403=>"000010100",
  49404=>"000000101",
  49405=>"001000100",
  49406=>"110000001",
  49407=>"100010110",
  49408=>"000111001",
  49409=>"111101001",
  49410=>"110010010",
  49411=>"111111011",
  49412=>"111110111",
  49413=>"000000011",
  49414=>"101100000",
  49415=>"001101110",
  49416=>"101011110",
  49417=>"110111100",
  49418=>"110111011",
  49419=>"101000010",
  49420=>"011111000",
  49421=>"111110010",
  49422=>"101100001",
  49423=>"101100111",
  49424=>"010111001",
  49425=>"110111101",
  49426=>"011110110",
  49427=>"100110111",
  49428=>"101000101",
  49429=>"100010001",
  49430=>"000011000",
  49431=>"001001100",
  49432=>"000011010",
  49433=>"110001010",
  49434=>"011100100",
  49435=>"101100011",
  49436=>"101111011",
  49437=>"000100110",
  49438=>"110111111",
  49439=>"110011010",
  49440=>"100000111",
  49441=>"001011110",
  49442=>"010001111",
  49443=>"011101010",
  49444=>"111010011",
  49445=>"011010101",
  49446=>"010000101",
  49447=>"100110101",
  49448=>"111111100",
  49449=>"010100111",
  49450=>"001101101",
  49451=>"011110111",
  49452=>"011010111",
  49453=>"110111101",
  49454=>"101101010",
  49455=>"100111111",
  49456=>"000101010",
  49457=>"111001101",
  49458=>"011100001",
  49459=>"010101010",
  49460=>"001111011",
  49461=>"001100011",
  49462=>"100000100",
  49463=>"100100001",
  49464=>"010110100",
  49465=>"110000111",
  49466=>"101110101",
  49467=>"100101011",
  49468=>"010000111",
  49469=>"010100010",
  49470=>"110011001",
  49471=>"100000111",
  49472=>"111010010",
  49473=>"101100011",
  49474=>"111010100",
  49475=>"010100110",
  49476=>"111111100",
  49477=>"100110110",
  49478=>"010110011",
  49479=>"000000011",
  49480=>"101001001",
  49481=>"001000110",
  49482=>"011000000",
  49483=>"100001110",
  49484=>"001011100",
  49485=>"001011011",
  49486=>"000101010",
  49487=>"011001001",
  49488=>"011010001",
  49489=>"100111101",
  49490=>"010110000",
  49491=>"001101101",
  49492=>"100011100",
  49493=>"101010001",
  49494=>"111110110",
  49495=>"000001000",
  49496=>"110011100",
  49497=>"001000000",
  49498=>"011010100",
  49499=>"101100010",
  49500=>"110011100",
  49501=>"000000011",
  49502=>"010000111",
  49503=>"000000100",
  49504=>"000010111",
  49505=>"101000110",
  49506=>"010001111",
  49507=>"100101111",
  49508=>"011011001",
  49509=>"011110000",
  49510=>"011001100",
  49511=>"000000010",
  49512=>"101111011",
  49513=>"101000000",
  49514=>"010101100",
  49515=>"110110000",
  49516=>"111010110",
  49517=>"000100111",
  49518=>"001000110",
  49519=>"101101100",
  49520=>"101001010",
  49521=>"111000011",
  49522=>"101101001",
  49523=>"110110111",
  49524=>"100000110",
  49525=>"011100010",
  49526=>"000110011",
  49527=>"111010110",
  49528=>"111000010",
  49529=>"000010011",
  49530=>"111101011",
  49531=>"011100010",
  49532=>"111001000",
  49533=>"011011001",
  49534=>"101110001",
  49535=>"110010110",
  49536=>"010000100",
  49537=>"100100010",
  49538=>"110010111",
  49539=>"000100001",
  49540=>"101011001",
  49541=>"010000111",
  49542=>"011110110",
  49543=>"010111010",
  49544=>"001111100",
  49545=>"101000000",
  49546=>"000000111",
  49547=>"011110111",
  49548=>"000100111",
  49549=>"010110100",
  49550=>"111101100",
  49551=>"111100110",
  49552=>"101101000",
  49553=>"010010011",
  49554=>"011000001",
  49555=>"010111001",
  49556=>"101011101",
  49557=>"000100111",
  49558=>"011100011",
  49559=>"010111110",
  49560=>"101001000",
  49561=>"001100001",
  49562=>"100100101",
  49563=>"001100111",
  49564=>"110110010",
  49565=>"000011000",
  49566=>"001000101",
  49567=>"100000010",
  49568=>"010100001",
  49569=>"010000000",
  49570=>"011010110",
  49571=>"101011001",
  49572=>"011011001",
  49573=>"100001000",
  49574=>"010111100",
  49575=>"001010110",
  49576=>"000101111",
  49577=>"100010010",
  49578=>"100000101",
  49579=>"001011001",
  49580=>"010101001",
  49581=>"010010010",
  49582=>"110010011",
  49583=>"101100001",
  49584=>"100111101",
  49585=>"010110101",
  49586=>"101100010",
  49587=>"001100011",
  49588=>"100010101",
  49589=>"011010100",
  49590=>"010110010",
  49591=>"011010100",
  49592=>"100000000",
  49593=>"000000100",
  49594=>"000010011",
  49595=>"100011000",
  49596=>"111100111",
  49597=>"111110101",
  49598=>"100101001",
  49599=>"110001110",
  49600=>"010001011",
  49601=>"011000101",
  49602=>"000001010",
  49603=>"000010010",
  49604=>"010101000",
  49605=>"110001100",
  49606=>"111110111",
  49607=>"000100111",
  49608=>"100011100",
  49609=>"110101110",
  49610=>"110000110",
  49611=>"110001000",
  49612=>"001010010",
  49613=>"000000010",
  49614=>"101010101",
  49615=>"000000100",
  49616=>"111010000",
  49617=>"011110110",
  49618=>"010011011",
  49619=>"110001001",
  49620=>"011100001",
  49621=>"101001000",
  49622=>"110101110",
  49623=>"101000101",
  49624=>"001001000",
  49625=>"111111101",
  49626=>"101111010",
  49627=>"111010111",
  49628=>"111001000",
  49629=>"111011001",
  49630=>"010111011",
  49631=>"110011100",
  49632=>"000110001",
  49633=>"100011100",
  49634=>"110000000",
  49635=>"001111100",
  49636=>"100111100",
  49637=>"100011100",
  49638=>"110001000",
  49639=>"100011001",
  49640=>"011010111",
  49641=>"100101001",
  49642=>"100000100",
  49643=>"010100101",
  49644=>"101110100",
  49645=>"011010111",
  49646=>"000010100",
  49647=>"111001010",
  49648=>"001010000",
  49649=>"010011111",
  49650=>"111000101",
  49651=>"100001011",
  49652=>"111101100",
  49653=>"000101000",
  49654=>"100101001",
  49655=>"001111111",
  49656=>"011000101",
  49657=>"111100000",
  49658=>"100101111",
  49659=>"010110100",
  49660=>"111010001",
  49661=>"111111110",
  49662=>"100011101",
  49663=>"111011110",
  49664=>"101101011",
  49665=>"010001010",
  49666=>"100000001",
  49667=>"101001010",
  49668=>"011111100",
  49669=>"101110100",
  49670=>"000100100",
  49671=>"010011001",
  49672=>"001011011",
  49673=>"010010001",
  49674=>"100111101",
  49675=>"110010010",
  49676=>"011000011",
  49677=>"110000100",
  49678=>"100001011",
  49679=>"100010011",
  49680=>"100001110",
  49681=>"000011101",
  49682=>"000011110",
  49683=>"100110100",
  49684=>"110100001",
  49685=>"000111010",
  49686=>"100000010",
  49687=>"000101111",
  49688=>"000011000",
  49689=>"111110010",
  49690=>"001000110",
  49691=>"010011100",
  49692=>"000010010",
  49693=>"110111001",
  49694=>"011101111",
  49695=>"001011101",
  49696=>"110001111",
  49697=>"010000010",
  49698=>"100010000",
  49699=>"011110101",
  49700=>"110101110",
  49701=>"010011101",
  49702=>"011101110",
  49703=>"110011001",
  49704=>"000000011",
  49705=>"000110000",
  49706=>"111010000",
  49707=>"000011100",
  49708=>"111110101",
  49709=>"111100010",
  49710=>"000000100",
  49711=>"000011000",
  49712=>"001010111",
  49713=>"010001001",
  49714=>"100001001",
  49715=>"000110000",
  49716=>"011101001",
  49717=>"101100000",
  49718=>"001000100",
  49719=>"101110110",
  49720=>"001100111",
  49721=>"100111100",
  49722=>"111000101",
  49723=>"011000010",
  49724=>"010011111",
  49725=>"000000110",
  49726=>"101101111",
  49727=>"111000001",
  49728=>"111000100",
  49729=>"100001000",
  49730=>"110110010",
  49731=>"001101111",
  49732=>"100011100",
  49733=>"000011111",
  49734=>"100000001",
  49735=>"011110001",
  49736=>"011001111",
  49737=>"101001110",
  49738=>"001100100",
  49739=>"100110100",
  49740=>"111000100",
  49741=>"100000110",
  49742=>"010001100",
  49743=>"010000011",
  49744=>"001001000",
  49745=>"100101110",
  49746=>"000101111",
  49747=>"010011000",
  49748=>"010000011",
  49749=>"010011001",
  49750=>"001000110",
  49751=>"001001111",
  49752=>"001111010",
  49753=>"100110011",
  49754=>"101101110",
  49755=>"010011010",
  49756=>"010001000",
  49757=>"101010010",
  49758=>"000010111",
  49759=>"011110001",
  49760=>"100000010",
  49761=>"010010000",
  49762=>"011001101",
  49763=>"010011010",
  49764=>"101100000",
  49765=>"101100111",
  49766=>"110001111",
  49767=>"100101000",
  49768=>"001001110",
  49769=>"010001111",
  49770=>"100000111",
  49771=>"011000011",
  49772=>"100010000",
  49773=>"111100000",
  49774=>"010101100",
  49775=>"011100010",
  49776=>"000100000",
  49777=>"000010110",
  49778=>"011010111",
  49779=>"101101001",
  49780=>"000111011",
  49781=>"000101000",
  49782=>"000110111",
  49783=>"011000110",
  49784=>"101001011",
  49785=>"000011111",
  49786=>"110000000",
  49787=>"000010011",
  49788=>"101101010",
  49789=>"001101011",
  49790=>"000110000",
  49791=>"101011110",
  49792=>"011110110",
  49793=>"111010011",
  49794=>"010000000",
  49795=>"010000011",
  49796=>"001010111",
  49797=>"111100100",
  49798=>"010110101",
  49799=>"100100000",
  49800=>"011011101",
  49801=>"100000011",
  49802=>"111001000",
  49803=>"100111111",
  49804=>"111111010",
  49805=>"000011110",
  49806=>"100111000",
  49807=>"001111110",
  49808=>"001101111",
  49809=>"110110000",
  49810=>"111011101",
  49811=>"110101110",
  49812=>"011110011",
  49813=>"110111010",
  49814=>"011001011",
  49815=>"011011010",
  49816=>"111100100",
  49817=>"111111111",
  49818=>"001100110",
  49819=>"000011100",
  49820=>"001010011",
  49821=>"001001000",
  49822=>"011111101",
  49823=>"111000111",
  49824=>"100101001",
  49825=>"010001111",
  49826=>"010000111",
  49827=>"011101000",
  49828=>"011011011",
  49829=>"101000101",
  49830=>"000101010",
  49831=>"000001000",
  49832=>"110101011",
  49833=>"101111001",
  49834=>"001000111",
  49835=>"100001111",
  49836=>"000011000",
  49837=>"100100110",
  49838=>"110110101",
  49839=>"110100000",
  49840=>"101000001",
  49841=>"010110011",
  49842=>"011100111",
  49843=>"010011101",
  49844=>"100111011",
  49845=>"010001101",
  49846=>"001000000",
  49847=>"100001010",
  49848=>"110000100",
  49849=>"000011111",
  49850=>"010001011",
  49851=>"001111101",
  49852=>"110010101",
  49853=>"000101011",
  49854=>"100101001",
  49855=>"010010010",
  49856=>"010011010",
  49857=>"111000111",
  49858=>"101001101",
  49859=>"010000101",
  49860=>"001111111",
  49861=>"101100110",
  49862=>"111110011",
  49863=>"011101011",
  49864=>"100000001",
  49865=>"010101000",
  49866=>"110000110",
  49867=>"110111101",
  49868=>"000000010",
  49869=>"011101111",
  49870=>"010000011",
  49871=>"001011000",
  49872=>"000111011",
  49873=>"101000111",
  49874=>"101110010",
  49875=>"000001100",
  49876=>"111000011",
  49877=>"100001010",
  49878=>"010100111",
  49879=>"001010001",
  49880=>"000001111",
  49881=>"110100010",
  49882=>"001010010",
  49883=>"111101001",
  49884=>"001000100",
  49885=>"111010000",
  49886=>"000110100",
  49887=>"001111010",
  49888=>"001000000",
  49889=>"000111100",
  49890=>"010011010",
  49891=>"010100110",
  49892=>"101011101",
  49893=>"001001111",
  49894=>"100000000",
  49895=>"010100011",
  49896=>"000011000",
  49897=>"101010111",
  49898=>"101010011",
  49899=>"101000101",
  49900=>"110100111",
  49901=>"101000101",
  49902=>"111101110",
  49903=>"001101110",
  49904=>"111100000",
  49905=>"101100010",
  49906=>"101010000",
  49907=>"110110101",
  49908=>"110000110",
  49909=>"110100110",
  49910=>"010100101",
  49911=>"011011011",
  49912=>"000000111",
  49913=>"100111010",
  49914=>"100110111",
  49915=>"010101011",
  49916=>"000111010",
  49917=>"101001111",
  49918=>"100000011",
  49919=>"000100110",
  49920=>"100111001",
  49921=>"010011111",
  49922=>"001101110",
  49923=>"010000100",
  49924=>"010000001",
  49925=>"010111100",
  49926=>"000100111",
  49927=>"111011111",
  49928=>"100000100",
  49929=>"111101100",
  49930=>"100101000",
  49931=>"110101110",
  49932=>"110100001",
  49933=>"010111111",
  49934=>"011111001",
  49935=>"101011011",
  49936=>"101101001",
  49937=>"010111111",
  49938=>"011011111",
  49939=>"001101110",
  49940=>"110000000",
  49941=>"011101100",
  49942=>"110111111",
  49943=>"100110111",
  49944=>"101001100",
  49945=>"000011100",
  49946=>"010111101",
  49947=>"000101100",
  49948=>"011001110",
  49949=>"100000101",
  49950=>"010100010",
  49951=>"101000111",
  49952=>"000101000",
  49953=>"100100010",
  49954=>"011110000",
  49955=>"110101011",
  49956=>"111011110",
  49957=>"101001011",
  49958=>"001101000",
  49959=>"000000001",
  49960=>"110110110",
  49961=>"100001000",
  49962=>"100110110",
  49963=>"111111010",
  49964=>"000110001",
  49965=>"001000001",
  49966=>"011101000",
  49967=>"100010010",
  49968=>"110011000",
  49969=>"000011110",
  49970=>"000110110",
  49971=>"000101001",
  49972=>"010011010",
  49973=>"010100111",
  49974=>"011100100",
  49975=>"001000110",
  49976=>"110011001",
  49977=>"000000011",
  49978=>"001110100",
  49979=>"001011001",
  49980=>"110100000",
  49981=>"110000110",
  49982=>"011001011",
  49983=>"100101111",
  49984=>"110001001",
  49985=>"101000110",
  49986=>"111010100",
  49987=>"001000101",
  49988=>"001000101",
  49989=>"010010000",
  49990=>"011001100",
  49991=>"000101101",
  49992=>"101001100",
  49993=>"100100110",
  49994=>"111111110",
  49995=>"001001101",
  49996=>"000111011",
  49997=>"011100100",
  49998=>"111100000",
  49999=>"001011101",
  50000=>"011000101",
  50001=>"110011111",
  50002=>"000001010",
  50003=>"001100001",
  50004=>"101001100",
  50005=>"001000100",
  50006=>"010111110",
  50007=>"001100100",
  50008=>"001110100",
  50009=>"101011111",
  50010=>"000011001",
  50011=>"001110110",
  50012=>"100101110",
  50013=>"101000001",
  50014=>"000111110",
  50015=>"001110010",
  50016=>"111100101",
  50017=>"001100001",
  50018=>"000111111",
  50019=>"010100101",
  50020=>"100000001",
  50021=>"001110011",
  50022=>"100001110",
  50023=>"101011100",
  50024=>"100001000",
  50025=>"010001011",
  50026=>"111100010",
  50027=>"000101010",
  50028=>"100000110",
  50029=>"000011011",
  50030=>"011000000",
  50031=>"001001010",
  50032=>"001111010",
  50033=>"101101001",
  50034=>"011100000",
  50035=>"110101100",
  50036=>"000110111",
  50037=>"011001011",
  50038=>"000101101",
  50039=>"010100100",
  50040=>"001110110",
  50041=>"000001100",
  50042=>"010010001",
  50043=>"001000011",
  50044=>"000110001",
  50045=>"111111000",
  50046=>"000110101",
  50047=>"101111101",
  50048=>"010001101",
  50049=>"110110011",
  50050=>"010110001",
  50051=>"000001010",
  50052=>"010000001",
  50053=>"101110110",
  50054=>"100100111",
  50055=>"011100001",
  50056=>"011010101",
  50057=>"111111101",
  50058=>"001000101",
  50059=>"010110100",
  50060=>"001001110",
  50061=>"011001101",
  50062=>"011100010",
  50063=>"100010111",
  50064=>"101001011",
  50065=>"101011011",
  50066=>"110000001",
  50067=>"101100100",
  50068=>"000100110",
  50069=>"101011111",
  50070=>"100011101",
  50071=>"111100101",
  50072=>"111111110",
  50073=>"010011100",
  50074=>"011100001",
  50075=>"111001100",
  50076=>"010010101",
  50077=>"110111001",
  50078=>"111011000",
  50079=>"010101011",
  50080=>"011001010",
  50081=>"101111000",
  50082=>"010000010",
  50083=>"010101100",
  50084=>"100000110",
  50085=>"001100010",
  50086=>"000000100",
  50087=>"001111110",
  50088=>"100110011",
  50089=>"110110101",
  50090=>"101011110",
  50091=>"001100100",
  50092=>"000101011",
  50093=>"010110011",
  50094=>"011000010",
  50095=>"111011011",
  50096=>"111100110",
  50097=>"110111101",
  50098=>"001111110",
  50099=>"100011001",
  50100=>"101110000",
  50101=>"100100110",
  50102=>"010100110",
  50103=>"011011011",
  50104=>"110110101",
  50105=>"101000010",
  50106=>"100101000",
  50107=>"010001010",
  50108=>"101101000",
  50109=>"011111100",
  50110=>"111000000",
  50111=>"100000011",
  50112=>"000010100",
  50113=>"100100001",
  50114=>"100000111",
  50115=>"000000100",
  50116=>"000001111",
  50117=>"001111010",
  50118=>"001111010",
  50119=>"001000000",
  50120=>"111010011",
  50121=>"111100101",
  50122=>"110100111",
  50123=>"111110100",
  50124=>"001001101",
  50125=>"010100010",
  50126=>"100100001",
  50127=>"101000000",
  50128=>"101000100",
  50129=>"101000010",
  50130=>"000010110",
  50131=>"100010101",
  50132=>"011000111",
  50133=>"111001001",
  50134=>"111111000",
  50135=>"100100111",
  50136=>"100100100",
  50137=>"010100000",
  50138=>"111111000",
  50139=>"111010001",
  50140=>"010101010",
  50141=>"111110111",
  50142=>"010001000",
  50143=>"011000010",
  50144=>"000010011",
  50145=>"100110101",
  50146=>"000110010",
  50147=>"010100000",
  50148=>"011000011",
  50149=>"010001010",
  50150=>"001101011",
  50151=>"110100100",
  50152=>"000100000",
  50153=>"011101110",
  50154=>"100110010",
  50155=>"001110000",
  50156=>"011101011",
  50157=>"011001111",
  50158=>"110101100",
  50159=>"000001111",
  50160=>"001001111",
  50161=>"001011010",
  50162=>"000010011",
  50163=>"011000000",
  50164=>"100111101",
  50165=>"000011011",
  50166=>"101110001",
  50167=>"001100011",
  50168=>"000111100",
  50169=>"111000111",
  50170=>"000100001",
  50171=>"111100111",
  50172=>"010101110",
  50173=>"100100111",
  50174=>"001101111",
  50175=>"000010100",
  50176=>"011111100",
  50177=>"001000110",
  50178=>"001100110",
  50179=>"000010110",
  50180=>"100100100",
  50181=>"110100110",
  50182=>"001001100",
  50183=>"101000010",
  50184=>"100000110",
  50185=>"000001100",
  50186=>"001101101",
  50187=>"101000010",
  50188=>"011011010",
  50189=>"101111110",
  50190=>"110011110",
  50191=>"111001010",
  50192=>"111010000",
  50193=>"001011011",
  50194=>"010000010",
  50195=>"011111011",
  50196=>"001101100",
  50197=>"110000000",
  50198=>"000011000",
  50199=>"110000100",
  50200=>"100011011",
  50201=>"101101011",
  50202=>"100000011",
  50203=>"110101111",
  50204=>"010000101",
  50205=>"110000001",
  50206=>"111011000",
  50207=>"010100000",
  50208=>"111110001",
  50209=>"000010111",
  50210=>"101100001",
  50211=>"110010110",
  50212=>"011010010",
  50213=>"010110101",
  50214=>"000011001",
  50215=>"110000101",
  50216=>"111010011",
  50217=>"011001000",
  50218=>"111001111",
  50219=>"010111111",
  50220=>"111100001",
  50221=>"100101010",
  50222=>"010010001",
  50223=>"011011011",
  50224=>"110111000",
  50225=>"000101011",
  50226=>"000010101",
  50227=>"001000100",
  50228=>"001100110",
  50229=>"111001000",
  50230=>"101110000",
  50231=>"110001001",
  50232=>"100110100",
  50233=>"000000110",
  50234=>"100011000",
  50235=>"100010110",
  50236=>"000111010",
  50237=>"111100101",
  50238=>"111110000",
  50239=>"011110011",
  50240=>"110100110",
  50241=>"101101110",
  50242=>"101011110",
  50243=>"111110000",
  50244=>"100001011",
  50245=>"111111011",
  50246=>"100101111",
  50247=>"111110110",
  50248=>"010010100",
  50249=>"100011100",
  50250=>"101011001",
  50251=>"010000001",
  50252=>"111111001",
  50253=>"010010011",
  50254=>"011100011",
  50255=>"011111010",
  50256=>"000110000",
  50257=>"100000000",
  50258=>"111011111",
  50259=>"110101000",
  50260=>"111001010",
  50261=>"111110111",
  50262=>"010100101",
  50263=>"111111010",
  50264=>"001011000",
  50265=>"000101001",
  50266=>"010111110",
  50267=>"010001000",
  50268=>"101011110",
  50269=>"000010010",
  50270=>"100111111",
  50271=>"110111111",
  50272=>"010101001",
  50273=>"111111001",
  50274=>"000001001",
  50275=>"101111101",
  50276=>"100111000",
  50277=>"111100001",
  50278=>"100000001",
  50279=>"000011000",
  50280=>"011010100",
  50281=>"110111010",
  50282=>"111010101",
  50283=>"010111100",
  50284=>"100001111",
  50285=>"000100000",
  50286=>"011000100",
  50287=>"000111011",
  50288=>"110101011",
  50289=>"110000111",
  50290=>"101110011",
  50291=>"011110110",
  50292=>"011111000",
  50293=>"110011111",
  50294=>"101101001",
  50295=>"000010011",
  50296=>"011101100",
  50297=>"110011000",
  50298=>"110010000",
  50299=>"011001010",
  50300=>"110000111",
  50301=>"100111011",
  50302=>"000110100",
  50303=>"100100111",
  50304=>"011001010",
  50305=>"010000110",
  50306=>"100011100",
  50307=>"100000111",
  50308=>"101010011",
  50309=>"010111011",
  50310=>"100111100",
  50311=>"110011110",
  50312=>"010001000",
  50313=>"000111111",
  50314=>"000110101",
  50315=>"110101100",
  50316=>"110110010",
  50317=>"100010010",
  50318=>"111000110",
  50319=>"111100100",
  50320=>"000110110",
  50321=>"010111111",
  50322=>"001110000",
  50323=>"100110100",
  50324=>"000111000",
  50325=>"101100011",
  50326=>"001011111",
  50327=>"000010111",
  50328=>"010010010",
  50329=>"100100010",
  50330=>"011110100",
  50331=>"010100111",
  50332=>"111111000",
  50333=>"110101010",
  50334=>"011110110",
  50335=>"100101111",
  50336=>"010001001",
  50337=>"000010001",
  50338=>"000101011",
  50339=>"001001100",
  50340=>"010010000",
  50341=>"000011110",
  50342=>"011001111",
  50343=>"100110000",
  50344=>"100011011",
  50345=>"000010110",
  50346=>"111010110",
  50347=>"011001110",
  50348=>"010100000",
  50349=>"111111111",
  50350=>"101010111",
  50351=>"000110010",
  50352=>"010001011",
  50353=>"001111110",
  50354=>"110111110",
  50355=>"011000111",
  50356=>"111011001",
  50357=>"110001001",
  50358=>"101101100",
  50359=>"000000110",
  50360=>"011110000",
  50361=>"001111010",
  50362=>"101101010",
  50363=>"100100001",
  50364=>"011110001",
  50365=>"000011010",
  50366=>"011000001",
  50367=>"001011000",
  50368=>"110100000",
  50369=>"101001110",
  50370=>"100011000",
  50371=>"101010100",
  50372=>"111011001",
  50373=>"000001011",
  50374=>"100101000",
  50375=>"011110101",
  50376=>"100101001",
  50377=>"001001101",
  50378=>"110000010",
  50379=>"110100111",
  50380=>"101010010",
  50381=>"001000011",
  50382=>"000001000",
  50383=>"000111000",
  50384=>"111100010",
  50385=>"101110100",
  50386=>"101000010",
  50387=>"100010101",
  50388=>"001000011",
  50389=>"010100000",
  50390=>"011000011",
  50391=>"001011110",
  50392=>"111101011",
  50393=>"000101100",
  50394=>"100111010",
  50395=>"111110001",
  50396=>"100000101",
  50397=>"111000001",
  50398=>"000100011",
  50399=>"010100101",
  50400=>"010111110",
  50401=>"110000100",
  50402=>"001011010",
  50403=>"111111111",
  50404=>"001101011",
  50405=>"100101110",
  50406=>"010001111",
  50407=>"000111111",
  50408=>"000001001",
  50409=>"110000000",
  50410=>"000111001",
  50411=>"110101101",
  50412=>"101110001",
  50413=>"000010011",
  50414=>"010001101",
  50415=>"111110111",
  50416=>"110111110",
  50417=>"000101101",
  50418=>"110101100",
  50419=>"100101011",
  50420=>"101010000",
  50421=>"001110110",
  50422=>"001000100",
  50423=>"100001000",
  50424=>"101101101",
  50425=>"111001010",
  50426=>"110101011",
  50427=>"101010111",
  50428=>"101010101",
  50429=>"101010001",
  50430=>"111101111",
  50431=>"000110101",
  50432=>"100000000",
  50433=>"101010111",
  50434=>"110011010",
  50435=>"011001011",
  50436=>"101111101",
  50437=>"100110010",
  50438=>"111000101",
  50439=>"001001100",
  50440=>"111110011",
  50441=>"011000000",
  50442=>"111100001",
  50443=>"101100001",
  50444=>"010011101",
  50445=>"010100010",
  50446=>"111011101",
  50447=>"110101101",
  50448=>"100111101",
  50449=>"100000100",
  50450=>"101011001",
  50451=>"100101111",
  50452=>"100101000",
  50453=>"111101000",
  50454=>"101100000",
  50455=>"011000100",
  50456=>"000110110",
  50457=>"011111111",
  50458=>"110010001",
  50459=>"101101010",
  50460=>"111110001",
  50461=>"100111101",
  50462=>"100010010",
  50463=>"000100000",
  50464=>"001011011",
  50465=>"000101110",
  50466=>"010111011",
  50467=>"011001101",
  50468=>"110011111",
  50469=>"111110000",
  50470=>"010010100",
  50471=>"111111110",
  50472=>"111111100",
  50473=>"101110110",
  50474=>"110010101",
  50475=>"000100101",
  50476=>"000100000",
  50477=>"110111111",
  50478=>"011001110",
  50479=>"011111000",
  50480=>"000010100",
  50481=>"010001110",
  50482=>"111010110",
  50483=>"010000110",
  50484=>"101001000",
  50485=>"100111101",
  50486=>"000010101",
  50487=>"010100110",
  50488=>"110110110",
  50489=>"111011100",
  50490=>"110001101",
  50491=>"100010111",
  50492=>"100000010",
  50493=>"101110001",
  50494=>"000110011",
  50495=>"110101011",
  50496=>"010011000",
  50497=>"111111111",
  50498=>"110100111",
  50499=>"010000010",
  50500=>"110011110",
  50501=>"111001111",
  50502=>"101011101",
  50503=>"111001010",
  50504=>"010001100",
  50505=>"111001100",
  50506=>"110111011",
  50507=>"001010011",
  50508=>"010011100",
  50509=>"010001000",
  50510=>"101111110",
  50511=>"010101001",
  50512=>"001011000",
  50513=>"101101111",
  50514=>"011011011",
  50515=>"100110001",
  50516=>"001110010",
  50517=>"110011011",
  50518=>"011011001",
  50519=>"111001010",
  50520=>"010000011",
  50521=>"000100100",
  50522=>"001111011",
  50523=>"010100101",
  50524=>"101101000",
  50525=>"110101111",
  50526=>"010010110",
  50527=>"101101100",
  50528=>"110101111",
  50529=>"111110010",
  50530=>"001101001",
  50531=>"100110001",
  50532=>"100110101",
  50533=>"111010100",
  50534=>"001001000",
  50535=>"101001100",
  50536=>"111110011",
  50537=>"111000111",
  50538=>"100001100",
  50539=>"101100010",
  50540=>"100011010",
  50541=>"111000111",
  50542=>"011100000",
  50543=>"110100110",
  50544=>"011101010",
  50545=>"101010101",
  50546=>"101011111",
  50547=>"111101101",
  50548=>"001000100",
  50549=>"000010101",
  50550=>"010000001",
  50551=>"111110000",
  50552=>"001110010",
  50553=>"001000101",
  50554=>"101101101",
  50555=>"111000011",
  50556=>"100001011",
  50557=>"000001011",
  50558=>"000100110",
  50559=>"111101111",
  50560=>"111001111",
  50561=>"001110010",
  50562=>"000001100",
  50563=>"011000101",
  50564=>"011000011",
  50565=>"000101110",
  50566=>"110101111",
  50567=>"000111000",
  50568=>"001000000",
  50569=>"000011010",
  50570=>"000101100",
  50571=>"000000110",
  50572=>"111001000",
  50573=>"001010100",
  50574=>"011000000",
  50575=>"010000100",
  50576=>"010101110",
  50577=>"000000110",
  50578=>"001110111",
  50579=>"111001000",
  50580=>"101100110",
  50581=>"010111110",
  50582=>"011111110",
  50583=>"010001001",
  50584=>"000101110",
  50585=>"011001000",
  50586=>"001011100",
  50587=>"101000101",
  50588=>"011100110",
  50589=>"111011110",
  50590=>"100111011",
  50591=>"111011100",
  50592=>"000011110",
  50593=>"111101000",
  50594=>"000010101",
  50595=>"000000000",
  50596=>"000111110",
  50597=>"111111001",
  50598=>"011010001",
  50599=>"010010000",
  50600=>"000100001",
  50601=>"101010101",
  50602=>"010111011",
  50603=>"100000000",
  50604=>"101110101",
  50605=>"011001001",
  50606=>"100010110",
  50607=>"110111000",
  50608=>"011110110",
  50609=>"001111001",
  50610=>"010101100",
  50611=>"011110010",
  50612=>"000100010",
  50613=>"010100010",
  50614=>"011010110",
  50615=>"010011111",
  50616=>"100100010",
  50617=>"111110110",
  50618=>"100000011",
  50619=>"101100011",
  50620=>"010110110",
  50621=>"000000101",
  50622=>"110111110",
  50623=>"101010010",
  50624=>"000000111",
  50625=>"011110010",
  50626=>"001100000",
  50627=>"110010001",
  50628=>"011101110",
  50629=>"000111110",
  50630=>"001100101",
  50631=>"000000010",
  50632=>"110100000",
  50633=>"111001110",
  50634=>"110111101",
  50635=>"101001011",
  50636=>"010111101",
  50637=>"111110000",
  50638=>"100101001",
  50639=>"100110110",
  50640=>"110101000",
  50641=>"000011011",
  50642=>"010111010",
  50643=>"000101100",
  50644=>"110010100",
  50645=>"101101111",
  50646=>"000111110",
  50647=>"111101111",
  50648=>"010110000",
  50649=>"100001111",
  50650=>"111111001",
  50651=>"001000001",
  50652=>"111101010",
  50653=>"100010011",
  50654=>"111101000",
  50655=>"011001110",
  50656=>"101111001",
  50657=>"000110000",
  50658=>"001110011",
  50659=>"011001100",
  50660=>"111111100",
  50661=>"010100000",
  50662=>"101000101",
  50663=>"011111000",
  50664=>"100110000",
  50665=>"010111001",
  50666=>"111011010",
  50667=>"111111111",
  50668=>"011001101",
  50669=>"001000000",
  50670=>"101011010",
  50671=>"001000001",
  50672=>"001110010",
  50673=>"001011000",
  50674=>"101100010",
  50675=>"101000001",
  50676=>"111111011",
  50677=>"101010010",
  50678=>"001011100",
  50679=>"000011100",
  50680=>"110001010",
  50681=>"011010001",
  50682=>"000011000",
  50683=>"011100011",
  50684=>"111110100",
  50685=>"111111111",
  50686=>"001111000",
  50687=>"100101001",
  50688=>"000110001",
  50689=>"001101100",
  50690=>"111111011",
  50691=>"010110111",
  50692=>"010000111",
  50693=>"001111010",
  50694=>"001100100",
  50695=>"011101011",
  50696=>"000010111",
  50697=>"101111010",
  50698=>"110110011",
  50699=>"111110000",
  50700=>"111010000",
  50701=>"011000010",
  50702=>"111010000",
  50703=>"100100111",
  50704=>"110101110",
  50705=>"101111101",
  50706=>"000010111",
  50707=>"010100010",
  50708=>"000010110",
  50709=>"110010000",
  50710=>"001101011",
  50711=>"100000000",
  50712=>"100111101",
  50713=>"011001011",
  50714=>"101011000",
  50715=>"010000010",
  50716=>"010110100",
  50717=>"111110110",
  50718=>"100100110",
  50719=>"010011011",
  50720=>"010001000",
  50721=>"000000111",
  50722=>"001010010",
  50723=>"000011000",
  50724=>"111110000",
  50725=>"010001111",
  50726=>"001011111",
  50727=>"101010100",
  50728=>"100010001",
  50729=>"000101001",
  50730=>"010101011",
  50731=>"100001001",
  50732=>"001111000",
  50733=>"011110110",
  50734=>"101010000",
  50735=>"111110010",
  50736=>"001000111",
  50737=>"011001010",
  50738=>"111011000",
  50739=>"000000110",
  50740=>"011001101",
  50741=>"111000001",
  50742=>"111000011",
  50743=>"000110110",
  50744=>"011001100",
  50745=>"101110010",
  50746=>"110001101",
  50747=>"111011000",
  50748=>"110000110",
  50749=>"001001000",
  50750=>"000101001",
  50751=>"000001000",
  50752=>"110011111",
  50753=>"100000000",
  50754=>"011010000",
  50755=>"011000000",
  50756=>"011100110",
  50757=>"111100001",
  50758=>"011010000",
  50759=>"001010001",
  50760=>"000000000",
  50761=>"101000000",
  50762=>"000010011",
  50763=>"111000101",
  50764=>"011000011",
  50765=>"101000100",
  50766=>"101011001",
  50767=>"001101111",
  50768=>"010111101",
  50769=>"010011001",
  50770=>"100110110",
  50771=>"000110000",
  50772=>"000010001",
  50773=>"000001101",
  50774=>"010111100",
  50775=>"111111010",
  50776=>"000011000",
  50777=>"000101111",
  50778=>"111111110",
  50779=>"000011101",
  50780=>"110110111",
  50781=>"000101100",
  50782=>"000101101",
  50783=>"110011010",
  50784=>"011101010",
  50785=>"001110100",
  50786=>"000010111",
  50787=>"000011111",
  50788=>"111110100",
  50789=>"101101000",
  50790=>"010111000",
  50791=>"000010100",
  50792=>"111001101",
  50793=>"101111010",
  50794=>"111010111",
  50795=>"111000111",
  50796=>"111000001",
  50797=>"000000110",
  50798=>"111100001",
  50799=>"100000010",
  50800=>"110101000",
  50801=>"000001000",
  50802=>"101110010",
  50803=>"001010100",
  50804=>"101111001",
  50805=>"111100101",
  50806=>"101001111",
  50807=>"000010110",
  50808=>"111111010",
  50809=>"010011111",
  50810=>"111001011",
  50811=>"110000010",
  50812=>"011000101",
  50813=>"010111110",
  50814=>"011111001",
  50815=>"100000110",
  50816=>"000100101",
  50817=>"110100010",
  50818=>"010100001",
  50819=>"001101110",
  50820=>"011101001",
  50821=>"000111100",
  50822=>"011001101",
  50823=>"101000000",
  50824=>"100111000",
  50825=>"010001100",
  50826=>"100010101",
  50827=>"001001110",
  50828=>"000000010",
  50829=>"000011101",
  50830=>"111011100",
  50831=>"101111010",
  50832=>"111110000",
  50833=>"110010011",
  50834=>"111001110",
  50835=>"100110110",
  50836=>"111100001",
  50837=>"000101101",
  50838=>"101011011",
  50839=>"100000111",
  50840=>"100101001",
  50841=>"000010110",
  50842=>"101101101",
  50843=>"101101110",
  50844=>"010001000",
  50845=>"010011001",
  50846=>"000010110",
  50847=>"101011101",
  50848=>"001111101",
  50849=>"010010010",
  50850=>"111110100",
  50851=>"110100100",
  50852=>"100000010",
  50853=>"100110111",
  50854=>"010011000",
  50855=>"010000011",
  50856=>"101111111",
  50857=>"101110101",
  50858=>"100000000",
  50859=>"110000000",
  50860=>"000101100",
  50861=>"001111010",
  50862=>"000110111",
  50863=>"010010011",
  50864=>"010110111",
  50865=>"001010100",
  50866=>"000000010",
  50867=>"101100101",
  50868=>"110101111",
  50869=>"111100100",
  50870=>"100101010",
  50871=>"110110111",
  50872=>"100000000",
  50873=>"011111010",
  50874=>"001001111",
  50875=>"010111000",
  50876=>"100010000",
  50877=>"111100100",
  50878=>"110010111",
  50879=>"001011100",
  50880=>"111101101",
  50881=>"000011100",
  50882=>"101101111",
  50883=>"010101101",
  50884=>"110010110",
  50885=>"000001011",
  50886=>"100010101",
  50887=>"011010000",
  50888=>"000001111",
  50889=>"110010001",
  50890=>"111101101",
  50891=>"101000001",
  50892=>"101100001",
  50893=>"010100100",
  50894=>"111011001",
  50895=>"111000110",
  50896=>"001100000",
  50897=>"011011100",
  50898=>"000011110",
  50899=>"010010010",
  50900=>"110000001",
  50901=>"101010111",
  50902=>"011011101",
  50903=>"010100010",
  50904=>"011010011",
  50905=>"101001010",
  50906=>"001110011",
  50907=>"111000101",
  50908=>"011101100",
  50909=>"010010110",
  50910=>"111000100",
  50911=>"101101100",
  50912=>"101111111",
  50913=>"001011001",
  50914=>"010110111",
  50915=>"001011010",
  50916=>"111010000",
  50917=>"100110110",
  50918=>"001100111",
  50919=>"000100001",
  50920=>"101100000",
  50921=>"001011000",
  50922=>"010000110",
  50923=>"001111110",
  50924=>"110101111",
  50925=>"110110110",
  50926=>"110010110",
  50927=>"100000110",
  50928=>"011100010",
  50929=>"001001110",
  50930=>"001100111",
  50931=>"101000100",
  50932=>"000001011",
  50933=>"100010001",
  50934=>"101001011",
  50935=>"000001000",
  50936=>"010101101",
  50937=>"010001100",
  50938=>"001011010",
  50939=>"001000000",
  50940=>"110011101",
  50941=>"111010100",
  50942=>"110110000",
  50943=>"110000010",
  50944=>"100011001",
  50945=>"011000101",
  50946=>"011011000",
  50947=>"001011001",
  50948=>"001111010",
  50949=>"000001001",
  50950=>"101010100",
  50951=>"110111111",
  50952=>"010000111",
  50953=>"111110110",
  50954=>"111110000",
  50955=>"111001110",
  50956=>"101101110",
  50957=>"100011110",
  50958=>"011110010",
  50959=>"001000110",
  50960=>"101100010",
  50961=>"100001010",
  50962=>"001101110",
  50963=>"010001001",
  50964=>"101100110",
  50965=>"110000101",
  50966=>"110110101",
  50967=>"000001110",
  50968=>"011110111",
  50969=>"111001101",
  50970=>"101000101",
  50971=>"100101010",
  50972=>"100100011",
  50973=>"011101111",
  50974=>"110110001",
  50975=>"110010100",
  50976=>"010100111",
  50977=>"111101101",
  50978=>"100001000",
  50979=>"111100100",
  50980=>"000010000",
  50981=>"111110000",
  50982=>"111111100",
  50983=>"010010101",
  50984=>"110000101",
  50985=>"100011000",
  50986=>"101000110",
  50987=>"000010111",
  50988=>"111111000",
  50989=>"010110001",
  50990=>"000000110",
  50991=>"000101001",
  50992=>"010101010",
  50993=>"101000011",
  50994=>"110111110",
  50995=>"110000010",
  50996=>"000110011",
  50997=>"101101011",
  50998=>"111110111",
  50999=>"100110111",
  51000=>"011010100",
  51001=>"100001010",
  51002=>"010111010",
  51003=>"011001000",
  51004=>"011101110",
  51005=>"011110100",
  51006=>"111001111",
  51007=>"111001110",
  51008=>"101011000",
  51009=>"001010010",
  51010=>"010001010",
  51011=>"111011011",
  51012=>"011101111",
  51013=>"000100101",
  51014=>"100101110",
  51015=>"001100100",
  51016=>"111000010",
  51017=>"111111011",
  51018=>"101011110",
  51019=>"000010011",
  51020=>"100110111",
  51021=>"011011110",
  51022=>"111111101",
  51023=>"011101001",
  51024=>"000000001",
  51025=>"010100001",
  51026=>"001100110",
  51027=>"100010100",
  51028=>"000000011",
  51029=>"000100100",
  51030=>"111101110",
  51031=>"011111100",
  51032=>"111001100",
  51033=>"000000110",
  51034=>"011000110",
  51035=>"101101010",
  51036=>"111010101",
  51037=>"111001111",
  51038=>"000001111",
  51039=>"011110110",
  51040=>"100000000",
  51041=>"010101000",
  51042=>"001011111",
  51043=>"001000010",
  51044=>"010100100",
  51045=>"111110111",
  51046=>"000001011",
  51047=>"100010111",
  51048=>"001000010",
  51049=>"010001001",
  51050=>"101101001",
  51051=>"110001011",
  51052=>"111000111",
  51053=>"011010110",
  51054=>"100001111",
  51055=>"110110010",
  51056=>"100111000",
  51057=>"111011110",
  51058=>"101011010",
  51059=>"011100001",
  51060=>"111001001",
  51061=>"000000111",
  51062=>"111001000",
  51063=>"000001111",
  51064=>"111010110",
  51065=>"011100111",
  51066=>"011100100",
  51067=>"101001111",
  51068=>"110110000",
  51069=>"000000100",
  51070=>"000100011",
  51071=>"000011110",
  51072=>"011101100",
  51073=>"110100011",
  51074=>"000101001",
  51075=>"000000010",
  51076=>"011000101",
  51077=>"010011011",
  51078=>"101001110",
  51079=>"100001000",
  51080=>"101000110",
  51081=>"001110011",
  51082=>"000110101",
  51083=>"001100011",
  51084=>"001000001",
  51085=>"011110000",
  51086=>"000011011",
  51087=>"010100110",
  51088=>"110000010",
  51089=>"001111111",
  51090=>"000001001",
  51091=>"000110000",
  51092=>"110100011",
  51093=>"011101100",
  51094=>"111101010",
  51095=>"000101111",
  51096=>"101100000",
  51097=>"000100010",
  51098=>"110100010",
  51099=>"011010011",
  51100=>"101010110",
  51101=>"110010001",
  51102=>"010001001",
  51103=>"110000011",
  51104=>"111100110",
  51105=>"110000110",
  51106=>"110011011",
  51107=>"101010011",
  51108=>"001010100",
  51109=>"110000011",
  51110=>"001111000",
  51111=>"100100110",
  51112=>"011011010",
  51113=>"100100001",
  51114=>"011100001",
  51115=>"111000001",
  51116=>"101101111",
  51117=>"101110111",
  51118=>"111010100",
  51119=>"001010110",
  51120=>"110001000",
  51121=>"110110010",
  51122=>"110010100",
  51123=>"111000101",
  51124=>"010111111",
  51125=>"011010110",
  51126=>"100101110",
  51127=>"001110001",
  51128=>"000100000",
  51129=>"110001101",
  51130=>"110111110",
  51131=>"100000011",
  51132=>"010101110",
  51133=>"000000100",
  51134=>"000000100",
  51135=>"011011000",
  51136=>"101111101",
  51137=>"111100101",
  51138=>"100000000",
  51139=>"111110101",
  51140=>"001011111",
  51141=>"000001001",
  51142=>"000011111",
  51143=>"010000000",
  51144=>"001010010",
  51145=>"110100110",
  51146=>"100110110",
  51147=>"111110101",
  51148=>"000100111",
  51149=>"010101001",
  51150=>"000100100",
  51151=>"100001011",
  51152=>"110111111",
  51153=>"110011110",
  51154=>"100101011",
  51155=>"111100001",
  51156=>"111101000",
  51157=>"111010010",
  51158=>"111111001",
  51159=>"000011101",
  51160=>"000000001",
  51161=>"000110100",
  51162=>"001010111",
  51163=>"001000010",
  51164=>"001010111",
  51165=>"000010000",
  51166=>"111011010",
  51167=>"000110101",
  51168=>"111101000",
  51169=>"111100101",
  51170=>"001001001",
  51171=>"011011101",
  51172=>"010000000",
  51173=>"000111110",
  51174=>"000010011",
  51175=>"000001000",
  51176=>"101101000",
  51177=>"010001011",
  51178=>"000001011",
  51179=>"001011111",
  51180=>"101001111",
  51181=>"111001100",
  51182=>"000001100",
  51183=>"001111111",
  51184=>"101100111",
  51185=>"010010100",
  51186=>"001001111",
  51187=>"001001001",
  51188=>"011100110",
  51189=>"010100001",
  51190=>"000111100",
  51191=>"000000000",
  51192=>"101000111",
  51193=>"101101000",
  51194=>"110000110",
  51195=>"010111101",
  51196=>"011011100",
  51197=>"101100001",
  51198=>"100111001",
  51199=>"101100111",
  51200=>"000110010",
  51201=>"111000001",
  51202=>"000110110",
  51203=>"101110110",
  51204=>"011111010",
  51205=>"000101101",
  51206=>"010110000",
  51207=>"101101011",
  51208=>"011001110",
  51209=>"011010101",
  51210=>"010001001",
  51211=>"010010000",
  51212=>"000011111",
  51213=>"101100111",
  51214=>"001110100",
  51215=>"000011011",
  51216=>"011110001",
  51217=>"011101110",
  51218=>"010011000",
  51219=>"010111000",
  51220=>"100011110",
  51221=>"000100110",
  51222=>"100000001",
  51223=>"010000000",
  51224=>"110111100",
  51225=>"001010010",
  51226=>"000000010",
  51227=>"100000010",
  51228=>"010010101",
  51229=>"111011100",
  51230=>"100000011",
  51231=>"000100100",
  51232=>"000001110",
  51233=>"100110100",
  51234=>"000101011",
  51235=>"010010001",
  51236=>"010010100",
  51237=>"101001100",
  51238=>"001111001",
  51239=>"111011010",
  51240=>"111011100",
  51241=>"000110000",
  51242=>"010101110",
  51243=>"000111101",
  51244=>"011010110",
  51245=>"001011001",
  51246=>"111001010",
  51247=>"011101110",
  51248=>"101110011",
  51249=>"100100000",
  51250=>"111010111",
  51251=>"110111101",
  51252=>"010010011",
  51253=>"111000011",
  51254=>"110111000",
  51255=>"000000111",
  51256=>"010100111",
  51257=>"110100001",
  51258=>"100100011",
  51259=>"110010100",
  51260=>"001001110",
  51261=>"011010111",
  51262=>"111100010",
  51263=>"000110100",
  51264=>"000110011",
  51265=>"000101010",
  51266=>"100110100",
  51267=>"011001100",
  51268=>"100101101",
  51269=>"101011000",
  51270=>"001101010",
  51271=>"000100001",
  51272=>"100110010",
  51273=>"001110100",
  51274=>"000100101",
  51275=>"001001011",
  51276=>"100011100",
  51277=>"101111100",
  51278=>"111111000",
  51279=>"010111000",
  51280=>"100000111",
  51281=>"100000000",
  51282=>"111111101",
  51283=>"011100100",
  51284=>"011000000",
  51285=>"001111010",
  51286=>"101010011",
  51287=>"000011010",
  51288=>"001101101",
  51289=>"010000100",
  51290=>"001110101",
  51291=>"110101001",
  51292=>"011111101",
  51293=>"001000000",
  51294=>"010011000",
  51295=>"010001011",
  51296=>"111011000",
  51297=>"100110111",
  51298=>"100101000",
  51299=>"000101001",
  51300=>"110111100",
  51301=>"111111110",
  51302=>"111110100",
  51303=>"010000111",
  51304=>"010101011",
  51305=>"001100010",
  51306=>"001101110",
  51307=>"011001011",
  51308=>"010101011",
  51309=>"101110100",
  51310=>"011000000",
  51311=>"001011111",
  51312=>"011001001",
  51313=>"010110000",
  51314=>"000001001",
  51315=>"100100010",
  51316=>"011100010",
  51317=>"000000010",
  51318=>"110110101",
  51319=>"110110010",
  51320=>"110110100",
  51321=>"110010111",
  51322=>"110001100",
  51323=>"100000010",
  51324=>"010111100",
  51325=>"010110111",
  51326=>"000001001",
  51327=>"001010101",
  51328=>"101001000",
  51329=>"000111010",
  51330=>"011001111",
  51331=>"011001111",
  51332=>"000110101",
  51333=>"000000111",
  51334=>"100010011",
  51335=>"011100101",
  51336=>"011101011",
  51337=>"011110001",
  51338=>"001001000",
  51339=>"000000101",
  51340=>"100100100",
  51341=>"001100110",
  51342=>"011011100",
  51343=>"011101011",
  51344=>"010111011",
  51345=>"000111001",
  51346=>"111101110",
  51347=>"011011010",
  51348=>"100011010",
  51349=>"100010100",
  51350=>"000011011",
  51351=>"101011101",
  51352=>"110000101",
  51353=>"110010011",
  51354=>"001011101",
  51355=>"111011010",
  51356=>"100101100",
  51357=>"110110110",
  51358=>"010100111",
  51359=>"101011111",
  51360=>"000101000",
  51361=>"110110111",
  51362=>"110100100",
  51363=>"111001010",
  51364=>"100011111",
  51365=>"100011101",
  51366=>"101111111",
  51367=>"101101011",
  51368=>"100100110",
  51369=>"100111110",
  51370=>"111101111",
  51371=>"111010000",
  51372=>"101011111",
  51373=>"111000110",
  51374=>"000110110",
  51375=>"101001101",
  51376=>"110111110",
  51377=>"001100011",
  51378=>"111100100",
  51379=>"000000001",
  51380=>"011011011",
  51381=>"101110011",
  51382=>"000110011",
  51383=>"111111000",
  51384=>"100100000",
  51385=>"011000000",
  51386=>"101100010",
  51387=>"111001011",
  51388=>"101110101",
  51389=>"111111101",
  51390=>"000000000",
  51391=>"010001100",
  51392=>"110111010",
  51393=>"001111010",
  51394=>"010100001",
  51395=>"111000100",
  51396=>"111110011",
  51397=>"010100101",
  51398=>"001101100",
  51399=>"001011111",
  51400=>"011100011",
  51401=>"001111110",
  51402=>"000100100",
  51403=>"101011111",
  51404=>"111100001",
  51405=>"011011101",
  51406=>"000011100",
  51407=>"111011101",
  51408=>"101101000",
  51409=>"101101001",
  51410=>"101011111",
  51411=>"011001100",
  51412=>"101101001",
  51413=>"100100101",
  51414=>"001110011",
  51415=>"011100000",
  51416=>"100001111",
  51417=>"100111100",
  51418=>"010101110",
  51419=>"111101000",
  51420=>"011000000",
  51421=>"010010111",
  51422=>"000000101",
  51423=>"101110111",
  51424=>"100001111",
  51425=>"101011111",
  51426=>"010100111",
  51427=>"000100101",
  51428=>"110110010",
  51429=>"000011011",
  51430=>"000001100",
  51431=>"000110011",
  51432=>"010001100",
  51433=>"001000110",
  51434=>"000011111",
  51435=>"110101010",
  51436=>"110011011",
  51437=>"000111001",
  51438=>"110000000",
  51439=>"000001101",
  51440=>"011010011",
  51441=>"111100111",
  51442=>"100000111",
  51443=>"000111101",
  51444=>"100000011",
  51445=>"110110111",
  51446=>"001010010",
  51447=>"000110000",
  51448=>"101000011",
  51449=>"101111011",
  51450=>"100101000",
  51451=>"100101001",
  51452=>"110000010",
  51453=>"000110011",
  51454=>"101010111",
  51455=>"100011101",
  51456=>"001010000",
  51457=>"101000000",
  51458=>"101101111",
  51459=>"010011000",
  51460=>"001110001",
  51461=>"001001010",
  51462=>"000010000",
  51463=>"000110000",
  51464=>"000011000",
  51465=>"001000100",
  51466=>"110111001",
  51467=>"001100000",
  51468=>"010010101",
  51469=>"011111010",
  51470=>"011100101",
  51471=>"010010011",
  51472=>"011001111",
  51473=>"011101100",
  51474=>"110010101",
  51475=>"100110110",
  51476=>"010000100",
  51477=>"010101111",
  51478=>"111010001",
  51479=>"011101101",
  51480=>"100111000",
  51481=>"000100111",
  51482=>"110100111",
  51483=>"000000110",
  51484=>"000000010",
  51485=>"010001100",
  51486=>"001100010",
  51487=>"110100100",
  51488=>"010001001",
  51489=>"001010000",
  51490=>"001101101",
  51491=>"000101111",
  51492=>"101011000",
  51493=>"001010000",
  51494=>"001000000",
  51495=>"110100010",
  51496=>"010000010",
  51497=>"100001100",
  51498=>"110000001",
  51499=>"110010010",
  51500=>"111111010",
  51501=>"000000111",
  51502=>"000100000",
  51503=>"001001010",
  51504=>"001000111",
  51505=>"010111001",
  51506=>"001000100",
  51507=>"010011000",
  51508=>"011001000",
  51509=>"100001000",
  51510=>"101010000",
  51511=>"010011100",
  51512=>"000000110",
  51513=>"100100001",
  51514=>"011000000",
  51515=>"100111100",
  51516=>"011010011",
  51517=>"010100010",
  51518=>"101011000",
  51519=>"010010000",
  51520=>"100101100",
  51521=>"110000110",
  51522=>"100000110",
  51523=>"001111101",
  51524=>"111111100",
  51525=>"001010111",
  51526=>"010100010",
  51527=>"100100100",
  51528=>"001101110",
  51529=>"100010110",
  51530=>"011010111",
  51531=>"001111001",
  51532=>"111010110",
  51533=>"111111101",
  51534=>"100010010",
  51535=>"110110011",
  51536=>"111101111",
  51537=>"000111010",
  51538=>"011010101",
  51539=>"000101101",
  51540=>"011101100",
  51541=>"000010111",
  51542=>"010010011",
  51543=>"101011011",
  51544=>"011000101",
  51545=>"100110011",
  51546=>"001110101",
  51547=>"001101111",
  51548=>"111100111",
  51549=>"011000110",
  51550=>"111110111",
  51551=>"000001111",
  51552=>"111111011",
  51553=>"001000001",
  51554=>"010111000",
  51555=>"001001000",
  51556=>"001000100",
  51557=>"000011100",
  51558=>"011100110",
  51559=>"000101011",
  51560=>"111110010",
  51561=>"100100010",
  51562=>"000010101",
  51563=>"100011011",
  51564=>"011000100",
  51565=>"101010110",
  51566=>"100101001",
  51567=>"000111111",
  51568=>"110110100",
  51569=>"011010100",
  51570=>"111110111",
  51571=>"101010010",
  51572=>"110001111",
  51573=>"001001000",
  51574=>"000110100",
  51575=>"010010110",
  51576=>"011111100",
  51577=>"011110111",
  51578=>"010011111",
  51579=>"100100100",
  51580=>"000100100",
  51581=>"100101010",
  51582=>"001110011",
  51583=>"000010111",
  51584=>"010010010",
  51585=>"011010011",
  51586=>"111000010",
  51587=>"010011001",
  51588=>"010110101",
  51589=>"110100000",
  51590=>"110101100",
  51591=>"111011010",
  51592=>"000000110",
  51593=>"001110101",
  51594=>"011101001",
  51595=>"100111101",
  51596=>"111001100",
  51597=>"101111101",
  51598=>"000100000",
  51599=>"110110010",
  51600=>"010110011",
  51601=>"010001100",
  51602=>"000001010",
  51603=>"111110110",
  51604=>"010000001",
  51605=>"111110000",
  51606=>"111101000",
  51607=>"110000100",
  51608=>"100000100",
  51609=>"011000000",
  51610=>"110010011",
  51611=>"101111010",
  51612=>"010111001",
  51613=>"000001110",
  51614=>"001111011",
  51615=>"010000011",
  51616=>"010100100",
  51617=>"000011101",
  51618=>"110010100",
  51619=>"110110110",
  51620=>"111101010",
  51621=>"000100110",
  51622=>"010010111",
  51623=>"110010010",
  51624=>"111100011",
  51625=>"011010100",
  51626=>"011010011",
  51627=>"000000100",
  51628=>"000111000",
  51629=>"111100111",
  51630=>"101111011",
  51631=>"010101101",
  51632=>"101000100",
  51633=>"011010111",
  51634=>"111001100",
  51635=>"000011111",
  51636=>"110010011",
  51637=>"011010001",
  51638=>"001010111",
  51639=>"001011010",
  51640=>"000000111",
  51641=>"000010010",
  51642=>"001010101",
  51643=>"111101010",
  51644=>"011110000",
  51645=>"000000001",
  51646=>"100011100",
  51647=>"111010010",
  51648=>"010100011",
  51649=>"000010101",
  51650=>"001100010",
  51651=>"001101000",
  51652=>"000011011",
  51653=>"001011100",
  51654=>"110100110",
  51655=>"110101000",
  51656=>"101000001",
  51657=>"000001001",
  51658=>"110010010",
  51659=>"011010000",
  51660=>"101111101",
  51661=>"010000001",
  51662=>"110110100",
  51663=>"111001110",
  51664=>"111001000",
  51665=>"010001000",
  51666=>"101010001",
  51667=>"010100010",
  51668=>"000010010",
  51669=>"001100001",
  51670=>"110011110",
  51671=>"011001100",
  51672=>"110000011",
  51673=>"100111101",
  51674=>"001110011",
  51675=>"011111101",
  51676=>"001011000",
  51677=>"110111001",
  51678=>"111010011",
  51679=>"001110110",
  51680=>"001101110",
  51681=>"000011111",
  51682=>"000001001",
  51683=>"110001111",
  51684=>"111101000",
  51685=>"110111111",
  51686=>"000011110",
  51687=>"110001100",
  51688=>"010111100",
  51689=>"010010101",
  51690=>"001010000",
  51691=>"001110101",
  51692=>"000011101",
  51693=>"111110100",
  51694=>"010010100",
  51695=>"101100111",
  51696=>"110001000",
  51697=>"111110010",
  51698=>"111011101",
  51699=>"111100111",
  51700=>"111111000",
  51701=>"100101101",
  51702=>"100110110",
  51703=>"111101110",
  51704=>"000011101",
  51705=>"010000001",
  51706=>"011011111",
  51707=>"001101001",
  51708=>"110100111",
  51709=>"110100111",
  51710=>"001111100",
  51711=>"001001011",
  51712=>"101000011",
  51713=>"001001101",
  51714=>"111101001",
  51715=>"110101001",
  51716=>"111001110",
  51717=>"110101011",
  51718=>"100001101",
  51719=>"010000110",
  51720=>"111100010",
  51721=>"100101101",
  51722=>"011000111",
  51723=>"000101000",
  51724=>"100001001",
  51725=>"110100110",
  51726=>"111111000",
  51727=>"010101110",
  51728=>"110011110",
  51729=>"001111110",
  51730=>"101100011",
  51731=>"110000010",
  51732=>"000011011",
  51733=>"010000001",
  51734=>"100000001",
  51735=>"011111101",
  51736=>"101010101",
  51737=>"101110011",
  51738=>"111011110",
  51739=>"100001100",
  51740=>"001101101",
  51741=>"100011010",
  51742=>"000101001",
  51743=>"000000000",
  51744=>"111101111",
  51745=>"010101101",
  51746=>"000010001",
  51747=>"101000011",
  51748=>"101011001",
  51749=>"010001101",
  51750=>"011110110",
  51751=>"111001100",
  51752=>"010000100",
  51753=>"011001100",
  51754=>"010001010",
  51755=>"101011101",
  51756=>"111011111",
  51757=>"111110001",
  51758=>"100001111",
  51759=>"011111110",
  51760=>"011101100",
  51761=>"111011111",
  51762=>"000110101",
  51763=>"010100111",
  51764=>"010101010",
  51765=>"101000001",
  51766=>"000010110",
  51767=>"000111100",
  51768=>"110100000",
  51769=>"111101100",
  51770=>"011000010",
  51771=>"010000100",
  51772=>"011001111",
  51773=>"010010010",
  51774=>"101101000",
  51775=>"100101100",
  51776=>"001001010",
  51777=>"000100100",
  51778=>"011001100",
  51779=>"101001010",
  51780=>"100011001",
  51781=>"000100110",
  51782=>"000011000",
  51783=>"101000001",
  51784=>"100110001",
  51785=>"010101010",
  51786=>"111111111",
  51787=>"101101011",
  51788=>"001000111",
  51789=>"010010110",
  51790=>"000100110",
  51791=>"100000111",
  51792=>"011011000",
  51793=>"110101000",
  51794=>"010100100",
  51795=>"000101011",
  51796=>"110110110",
  51797=>"010101110",
  51798=>"111011010",
  51799=>"001011011",
  51800=>"000110101",
  51801=>"110101011",
  51802=>"010010010",
  51803=>"000100000",
  51804=>"011111101",
  51805=>"110010111",
  51806=>"111111101",
  51807=>"011111011",
  51808=>"110101011",
  51809=>"000011011",
  51810=>"010000010",
  51811=>"111001111",
  51812=>"111101100",
  51813=>"100001101",
  51814=>"000110101",
  51815=>"000010101",
  51816=>"110000001",
  51817=>"001110001",
  51818=>"100000001",
  51819=>"011111110",
  51820=>"100100100",
  51821=>"111001111",
  51822=>"101111110",
  51823=>"100000111",
  51824=>"101111000",
  51825=>"011111101",
  51826=>"000001001",
  51827=>"111001001",
  51828=>"101011101",
  51829=>"100101110",
  51830=>"101110001",
  51831=>"111100011",
  51832=>"110100111",
  51833=>"010101010",
  51834=>"101000001",
  51835=>"010011000",
  51836=>"100000001",
  51837=>"001101111",
  51838=>"010100000",
  51839=>"011101100",
  51840=>"111110011",
  51841=>"000101000",
  51842=>"000111000",
  51843=>"100111010",
  51844=>"111011010",
  51845=>"110101011",
  51846=>"001001001",
  51847=>"000100000",
  51848=>"001001101",
  51849=>"101010100",
  51850=>"100111111",
  51851=>"001000110",
  51852=>"000011011",
  51853=>"011000011",
  51854=>"011111110",
  51855=>"111100001",
  51856=>"011010111",
  51857=>"111110101",
  51858=>"111111111",
  51859=>"110001101",
  51860=>"101011110",
  51861=>"101101111",
  51862=>"000110001",
  51863=>"100000110",
  51864=>"101001111",
  51865=>"001000000",
  51866=>"100010000",
  51867=>"101110010",
  51868=>"011010110",
  51869=>"000001000",
  51870=>"010000000",
  51871=>"110111101",
  51872=>"101001001",
  51873=>"100000110",
  51874=>"001010010",
  51875=>"000101001",
  51876=>"010110011",
  51877=>"001100011",
  51878=>"001100110",
  51879=>"001100000",
  51880=>"001110001",
  51881=>"000011001",
  51882=>"011001110",
  51883=>"010001000",
  51884=>"111000110",
  51885=>"010000000",
  51886=>"010010100",
  51887=>"111001010",
  51888=>"110100010",
  51889=>"101010001",
  51890=>"110111100",
  51891=>"001111011",
  51892=>"010110011",
  51893=>"001011011",
  51894=>"011101011",
  51895=>"100100011",
  51896=>"000010010",
  51897=>"101010100",
  51898=>"100000101",
  51899=>"101111110",
  51900=>"000010000",
  51901=>"000000101",
  51902=>"000000111",
  51903=>"011001001",
  51904=>"110110100",
  51905=>"001110010",
  51906=>"000010010",
  51907=>"101000110",
  51908=>"110011011",
  51909=>"101011010",
  51910=>"100111011",
  51911=>"001000010",
  51912=>"000110011",
  51913=>"001010001",
  51914=>"111101010",
  51915=>"010111010",
  51916=>"000000001",
  51917=>"010011100",
  51918=>"111101001",
  51919=>"000001011",
  51920=>"110101100",
  51921=>"111110100",
  51922=>"001001110",
  51923=>"011001011",
  51924=>"110001000",
  51925=>"000111001",
  51926=>"000001011",
  51927=>"011110011",
  51928=>"001000101",
  51929=>"111010101",
  51930=>"010111000",
  51931=>"110010001",
  51932=>"000010000",
  51933=>"011111111",
  51934=>"110101110",
  51935=>"110110010",
  51936=>"100100010",
  51937=>"010100111",
  51938=>"010111110",
  51939=>"111101001",
  51940=>"001001101",
  51941=>"001101010",
  51942=>"101001101",
  51943=>"001010001",
  51944=>"110110001",
  51945=>"011001011",
  51946=>"111100111",
  51947=>"111111100",
  51948=>"010100000",
  51949=>"111100101",
  51950=>"110110101",
  51951=>"000100100",
  51952=>"101100011",
  51953=>"111101000",
  51954=>"011000100",
  51955=>"101110000",
  51956=>"000001110",
  51957=>"111100101",
  51958=>"111101000",
  51959=>"110001101",
  51960=>"001110110",
  51961=>"001000101",
  51962=>"101000101",
  51963=>"010000110",
  51964=>"000110100",
  51965=>"011111110",
  51966=>"000110110",
  51967=>"001111110",
  51968=>"100000001",
  51969=>"011010111",
  51970=>"100010001",
  51971=>"111101010",
  51972=>"101100000",
  51973=>"110011010",
  51974=>"001010101",
  51975=>"111111001",
  51976=>"110111101",
  51977=>"001101100",
  51978=>"111101101",
  51979=>"001001010",
  51980=>"010000101",
  51981=>"011110111",
  51982=>"100011001",
  51983=>"011101101",
  51984=>"001011111",
  51985=>"011010000",
  51986=>"111110001",
  51987=>"100110110",
  51988=>"010010101",
  51989=>"101100000",
  51990=>"110001010",
  51991=>"100111011",
  51992=>"011000101",
  51993=>"000011100",
  51994=>"000110110",
  51995=>"101111001",
  51996=>"110111111",
  51997=>"111011011",
  51998=>"100111000",
  51999=>"011000011",
  52000=>"111111010",
  52001=>"011000100",
  52002=>"111110110",
  52003=>"010110111",
  52004=>"010100101",
  52005=>"111010101",
  52006=>"001001101",
  52007=>"000001101",
  52008=>"010110011",
  52009=>"101101101",
  52010=>"100000111",
  52011=>"101000101",
  52012=>"100101111",
  52013=>"111011101",
  52014=>"010100010",
  52015=>"100000100",
  52016=>"100011101",
  52017=>"001001100",
  52018=>"010001010",
  52019=>"110000110",
  52020=>"111001011",
  52021=>"000001010",
  52022=>"001010101",
  52023=>"000010010",
  52024=>"001001100",
  52025=>"011011011",
  52026=>"110010001",
  52027=>"001100110",
  52028=>"001111000",
  52029=>"000011000",
  52030=>"101100100",
  52031=>"110000111",
  52032=>"000110111",
  52033=>"000110111",
  52034=>"100011010",
  52035=>"111100001",
  52036=>"100101100",
  52037=>"010000010",
  52038=>"110101100",
  52039=>"011111010",
  52040=>"100010010",
  52041=>"011111110",
  52042=>"110111001",
  52043=>"110100010",
  52044=>"001111100",
  52045=>"011010100",
  52046=>"100000000",
  52047=>"111111110",
  52048=>"000101010",
  52049=>"100111000",
  52050=>"101010001",
  52051=>"000100011",
  52052=>"100011010",
  52053=>"101110010",
  52054=>"001011101",
  52055=>"000101101",
  52056=>"010011000",
  52057=>"010010101",
  52058=>"111110010",
  52059=>"101010111",
  52060=>"111101111",
  52061=>"011000001",
  52062=>"111101001",
  52063=>"100110000",
  52064=>"100010001",
  52065=>"010001101",
  52066=>"100011100",
  52067=>"111010010",
  52068=>"110000000",
  52069=>"100111000",
  52070=>"110010001",
  52071=>"001101011",
  52072=>"010010110",
  52073=>"010000110",
  52074=>"110001111",
  52075=>"110010000",
  52076=>"111111110",
  52077=>"101100111",
  52078=>"111010100",
  52079=>"010001010",
  52080=>"100111011",
  52081=>"010101111",
  52082=>"000001111",
  52083=>"011101101",
  52084=>"111010000",
  52085=>"100101100",
  52086=>"001001100",
  52087=>"100111010",
  52088=>"110010101",
  52089=>"000100101",
  52090=>"001101110",
  52091=>"100110101",
  52092=>"000000000",
  52093=>"000011101",
  52094=>"111011111",
  52095=>"100010110",
  52096=>"111000101",
  52097=>"001111010",
  52098=>"100000100",
  52099=>"000010000",
  52100=>"010110110",
  52101=>"010110001",
  52102=>"001000110",
  52103=>"110111011",
  52104=>"100111111",
  52105=>"010100111",
  52106=>"100111011",
  52107=>"011101111",
  52108=>"110110111",
  52109=>"000101110",
  52110=>"001001111",
  52111=>"110010111",
  52112=>"100000010",
  52113=>"011001001",
  52114=>"000010000",
  52115=>"111011100",
  52116=>"000101001",
  52117=>"101111001",
  52118=>"111111000",
  52119=>"101111111",
  52120=>"110010101",
  52121=>"111001010",
  52122=>"111001111",
  52123=>"010000001",
  52124=>"000101110",
  52125=>"011111010",
  52126=>"111010011",
  52127=>"001010100",
  52128=>"001001001",
  52129=>"111101101",
  52130=>"011110101",
  52131=>"010100100",
  52132=>"110010100",
  52133=>"001000010",
  52134=>"000110010",
  52135=>"011101010",
  52136=>"101111000",
  52137=>"100110010",
  52138=>"010101010",
  52139=>"101110010",
  52140=>"000010011",
  52141=>"111001111",
  52142=>"000101000",
  52143=>"011011111",
  52144=>"100100001",
  52145=>"111101011",
  52146=>"110001111",
  52147=>"111111011",
  52148=>"110010100",
  52149=>"110010110",
  52150=>"000001111",
  52151=>"001011011",
  52152=>"010101100",
  52153=>"010000111",
  52154=>"001111100",
  52155=>"110001100",
  52156=>"101001000",
  52157=>"101110010",
  52158=>"110010010",
  52159=>"001001001",
  52160=>"110001010",
  52161=>"111110010",
  52162=>"000101010",
  52163=>"110111100",
  52164=>"001101111",
  52165=>"110101011",
  52166=>"011011001",
  52167=>"000111001",
  52168=>"010110000",
  52169=>"101101010",
  52170=>"111101110",
  52171=>"000000110",
  52172=>"110000011",
  52173=>"000110011",
  52174=>"100011111",
  52175=>"001011111",
  52176=>"101100011",
  52177=>"111011111",
  52178=>"001000101",
  52179=>"010001000",
  52180=>"010110001",
  52181=>"111011111",
  52182=>"010110011",
  52183=>"000010010",
  52184=>"000011101",
  52185=>"001000011",
  52186=>"101001001",
  52187=>"010001101",
  52188=>"111000100",
  52189=>"110110010",
  52190=>"111011101",
  52191=>"000001000",
  52192=>"000000111",
  52193=>"010111001",
  52194=>"110100111",
  52195=>"111111001",
  52196=>"010000100",
  52197=>"110000101",
  52198=>"110100001",
  52199=>"100110001",
  52200=>"000100010",
  52201=>"010010001",
  52202=>"001101111",
  52203=>"011110001",
  52204=>"111100001",
  52205=>"000011101",
  52206=>"101001010",
  52207=>"000010110",
  52208=>"011101001",
  52209=>"111100010",
  52210=>"100000011",
  52211=>"111110110",
  52212=>"111010001",
  52213=>"011011010",
  52214=>"100011100",
  52215=>"001010100",
  52216=>"000010000",
  52217=>"011110011",
  52218=>"010111000",
  52219=>"101000111",
  52220=>"001001100",
  52221=>"100111011",
  52222=>"000000001",
  52223=>"000101101",
  52224=>"100111010",
  52225=>"010110110",
  52226=>"010100010",
  52227=>"110000100",
  52228=>"000110101",
  52229=>"001100100",
  52230=>"100010101",
  52231=>"110100110",
  52232=>"111001010",
  52233=>"010000000",
  52234=>"101100111",
  52235=>"000011101",
  52236=>"001010010",
  52237=>"111001111",
  52238=>"010110010",
  52239=>"000010111",
  52240=>"001100000",
  52241=>"000000001",
  52242=>"111111011",
  52243=>"111100000",
  52244=>"111111010",
  52245=>"100001101",
  52246=>"100010110",
  52247=>"101010101",
  52248=>"110111101",
  52249=>"111110111",
  52250=>"011101010",
  52251=>"011000100",
  52252=>"000010111",
  52253=>"100111000",
  52254=>"010001100",
  52255=>"010010011",
  52256=>"010111000",
  52257=>"111010000",
  52258=>"100100111",
  52259=>"011000000",
  52260=>"111100000",
  52261=>"001101010",
  52262=>"011100101",
  52263=>"011010100",
  52264=>"000111001",
  52265=>"111011111",
  52266=>"001101111",
  52267=>"011011100",
  52268=>"001100001",
  52269=>"000100100",
  52270=>"111010100",
  52271=>"110011010",
  52272=>"011111110",
  52273=>"100001001",
  52274=>"011000100",
  52275=>"111111111",
  52276=>"011010010",
  52277=>"000110111",
  52278=>"000111011",
  52279=>"010111100",
  52280=>"110110011",
  52281=>"110010000",
  52282=>"011111001",
  52283=>"001010110",
  52284=>"010100100",
  52285=>"011101001",
  52286=>"110010000",
  52287=>"111100111",
  52288=>"010100110",
  52289=>"111010001",
  52290=>"100111010",
  52291=>"001111011",
  52292=>"111100101",
  52293=>"101100011",
  52294=>"001000000",
  52295=>"101110010",
  52296=>"011011010",
  52297=>"011010110",
  52298=>"101100111",
  52299=>"100001110",
  52300=>"010001001",
  52301=>"011101001",
  52302=>"111011000",
  52303=>"011101110",
  52304=>"100010011",
  52305=>"100100011",
  52306=>"001011010",
  52307=>"010000000",
  52308=>"101111111",
  52309=>"100111111",
  52310=>"011101110",
  52311=>"000011010",
  52312=>"001010100",
  52313=>"011001110",
  52314=>"100100000",
  52315=>"011111001",
  52316=>"000100110",
  52317=>"001111010",
  52318=>"111000110",
  52319=>"100000001",
  52320=>"111100100",
  52321=>"111101001",
  52322=>"100101001",
  52323=>"001111110",
  52324=>"000011000",
  52325=>"111110010",
  52326=>"111101100",
  52327=>"011100101",
  52328=>"111010110",
  52329=>"111000110",
  52330=>"111111111",
  52331=>"010000111",
  52332=>"011010011",
  52333=>"111001100",
  52334=>"000100001",
  52335=>"101000111",
  52336=>"011111000",
  52337=>"101001000",
  52338=>"011101100",
  52339=>"101101001",
  52340=>"101001001",
  52341=>"100001100",
  52342=>"010111010",
  52343=>"110110000",
  52344=>"110111011",
  52345=>"000010001",
  52346=>"000000000",
  52347=>"100001000",
  52348=>"100100000",
  52349=>"010101100",
  52350=>"010000000",
  52351=>"100001011",
  52352=>"110101011",
  52353=>"110110001",
  52354=>"110100000",
  52355=>"110000100",
  52356=>"001011011",
  52357=>"111011011",
  52358=>"110011010",
  52359=>"000010000",
  52360=>"101011001",
  52361=>"110111110",
  52362=>"110101000",
  52363=>"011000010",
  52364=>"011100111",
  52365=>"110100100",
  52366=>"000100010",
  52367=>"000110001",
  52368=>"011000000",
  52369=>"011101011",
  52370=>"001000011",
  52371=>"011001101",
  52372=>"101010101",
  52373=>"001001000",
  52374=>"011000011",
  52375=>"010010011",
  52376=>"010001110",
  52377=>"111100111",
  52378=>"000011000",
  52379=>"000010000",
  52380=>"001011111",
  52381=>"100001101",
  52382=>"001110001",
  52383=>"000000010",
  52384=>"010011000",
  52385=>"010001101",
  52386=>"101110001",
  52387=>"001100110",
  52388=>"100111110",
  52389=>"100001000",
  52390=>"000110100",
  52391=>"100010001",
  52392=>"000101000",
  52393=>"110010111",
  52394=>"110010110",
  52395=>"000001001",
  52396=>"000001000",
  52397=>"101101100",
  52398=>"000001100",
  52399=>"110101001",
  52400=>"111000000",
  52401=>"101100001",
  52402=>"001101111",
  52403=>"101010100",
  52404=>"001000010",
  52405=>"000101111",
  52406=>"111101001",
  52407=>"101000011",
  52408=>"010110111",
  52409=>"001111000",
  52410=>"100000100",
  52411=>"010101111",
  52412=>"011101011",
  52413=>"000011101",
  52414=>"110110100",
  52415=>"100110010",
  52416=>"010000010",
  52417=>"100000110",
  52418=>"111100011",
  52419=>"000010010",
  52420=>"111110010",
  52421=>"111000000",
  52422=>"000000001",
  52423=>"111000001",
  52424=>"000001110",
  52425=>"000000001",
  52426=>"010001111",
  52427=>"110010111",
  52428=>"111011001",
  52429=>"010110001",
  52430=>"011010010",
  52431=>"111111111",
  52432=>"101100110",
  52433=>"011100101",
  52434=>"000000011",
  52435=>"111011101",
  52436=>"001101011",
  52437=>"101000110",
  52438=>"011101100",
  52439=>"010100011",
  52440=>"100011010",
  52441=>"111100100",
  52442=>"101101000",
  52443=>"110000000",
  52444=>"000101010",
  52445=>"111001000",
  52446=>"000010001",
  52447=>"110110100",
  52448=>"111110010",
  52449=>"101101011",
  52450=>"011010010",
  52451=>"111000111",
  52452=>"000110000",
  52453=>"110101101",
  52454=>"110101111",
  52455=>"111010000",
  52456=>"011110100",
  52457=>"100000000",
  52458=>"010001000",
  52459=>"000001100",
  52460=>"000010000",
  52461=>"111000100",
  52462=>"111011001",
  52463=>"101001011",
  52464=>"101010001",
  52465=>"011111111",
  52466=>"001100101",
  52467=>"100001000",
  52468=>"101011000",
  52469=>"101000110",
  52470=>"000011101",
  52471=>"000101101",
  52472=>"010100000",
  52473=>"001010111",
  52474=>"100010101",
  52475=>"001111101",
  52476=>"100011000",
  52477=>"000111010",
  52478=>"011111101",
  52479=>"001101001",
  52480=>"110010011",
  52481=>"101000111",
  52482=>"100011101",
  52483=>"111100100",
  52484=>"111110010",
  52485=>"000001100",
  52486=>"110011001",
  52487=>"111110101",
  52488=>"110011111",
  52489=>"010100101",
  52490=>"001001110",
  52491=>"100001101",
  52492=>"110000111",
  52493=>"110001011",
  52494=>"101000010",
  52495=>"110100010",
  52496=>"000101100",
  52497=>"011010011",
  52498=>"001000110",
  52499=>"101001001",
  52500=>"111001110",
  52501=>"011111001",
  52502=>"101100101",
  52503=>"001101101",
  52504=>"001100010",
  52505=>"100100001",
  52506=>"101011010",
  52507=>"110000010",
  52508=>"001111000",
  52509=>"101011101",
  52510=>"100011010",
  52511=>"011000010",
  52512=>"111111011",
  52513=>"110011111",
  52514=>"101111001",
  52515=>"111101010",
  52516=>"110110001",
  52517=>"001101101",
  52518=>"000010001",
  52519=>"100000000",
  52520=>"000111110",
  52521=>"001101000",
  52522=>"001100001",
  52523=>"110110110",
  52524=>"110111011",
  52525=>"000101101",
  52526=>"010011011",
  52527=>"110001010",
  52528=>"101000000",
  52529=>"000000100",
  52530=>"110001100",
  52531=>"110010110",
  52532=>"101001101",
  52533=>"110000000",
  52534=>"001110111",
  52535=>"111011001",
  52536=>"111110000",
  52537=>"011100110",
  52538=>"111011101",
  52539=>"001001111",
  52540=>"101001111",
  52541=>"001111010",
  52542=>"100111101",
  52543=>"111011000",
  52544=>"100111000",
  52545=>"110101011",
  52546=>"111001010",
  52547=>"001110101",
  52548=>"110000100",
  52549=>"000001010",
  52550=>"100010001",
  52551=>"000001101",
  52552=>"111100000",
  52553=>"111000011",
  52554=>"000001011",
  52555=>"000110110",
  52556=>"111010011",
  52557=>"000011111",
  52558=>"110010110",
  52559=>"111011011",
  52560=>"111001100",
  52561=>"011001101",
  52562=>"101010000",
  52563=>"101011111",
  52564=>"100111111",
  52565=>"011111111",
  52566=>"111010101",
  52567=>"101110110",
  52568=>"000000100",
  52569=>"011010010",
  52570=>"010010001",
  52571=>"000010001",
  52572=>"110111001",
  52573=>"111101010",
  52574=>"010011011",
  52575=>"100001111",
  52576=>"011000100",
  52577=>"001110110",
  52578=>"101110100",
  52579=>"010001010",
  52580=>"111000010",
  52581=>"101101111",
  52582=>"110001100",
  52583=>"001000000",
  52584=>"010001001",
  52585=>"001010001",
  52586=>"010101011",
  52587=>"111000111",
  52588=>"100010000",
  52589=>"100000011",
  52590=>"001101110",
  52591=>"111100110",
  52592=>"011010111",
  52593=>"100001000",
  52594=>"110111100",
  52595=>"101011110",
  52596=>"101100000",
  52597=>"101000000",
  52598=>"101101000",
  52599=>"001000011",
  52600=>"110110111",
  52601=>"001010100",
  52602=>"111110110",
  52603=>"011100100",
  52604=>"010000000",
  52605=>"001110111",
  52606=>"011101111",
  52607=>"010001110",
  52608=>"111111111",
  52609=>"010100010",
  52610=>"000010000",
  52611=>"001010000",
  52612=>"000111000",
  52613=>"100101001",
  52614=>"001100101",
  52615=>"101100101",
  52616=>"110000001",
  52617=>"011110110",
  52618=>"100110001",
  52619=>"101101100",
  52620=>"000111100",
  52621=>"111000011",
  52622=>"100011000",
  52623=>"101110001",
  52624=>"110011010",
  52625=>"000111010",
  52626=>"111110100",
  52627=>"101000110",
  52628=>"111110011",
  52629=>"011100110",
  52630=>"101000111",
  52631=>"001010010",
  52632=>"111001101",
  52633=>"001011000",
  52634=>"001111101",
  52635=>"011110101",
  52636=>"010100111",
  52637=>"010000001",
  52638=>"011100110",
  52639=>"100100011",
  52640=>"111110100",
  52641=>"000110100",
  52642=>"011001001",
  52643=>"011100000",
  52644=>"010111110",
  52645=>"111011110",
  52646=>"010010010",
  52647=>"001000111",
  52648=>"110111111",
  52649=>"000011111",
  52650=>"011000001",
  52651=>"100010111",
  52652=>"111111101",
  52653=>"100000110",
  52654=>"101000000",
  52655=>"011011110",
  52656=>"010101010",
  52657=>"010100111",
  52658=>"111100100",
  52659=>"011011101",
  52660=>"000110100",
  52661=>"010101001",
  52662=>"010011101",
  52663=>"100110010",
  52664=>"111111111",
  52665=>"101111110",
  52666=>"111101111",
  52667=>"110101111",
  52668=>"111110101",
  52669=>"001111001",
  52670=>"001111011",
  52671=>"100100111",
  52672=>"000011111",
  52673=>"110111011",
  52674=>"000010110",
  52675=>"100111011",
  52676=>"110101011",
  52677=>"111001011",
  52678=>"001100101",
  52679=>"101000010",
  52680=>"000110101",
  52681=>"100110101",
  52682=>"001101010",
  52683=>"111010011",
  52684=>"111000001",
  52685=>"100010100",
  52686=>"011101100",
  52687=>"110101101",
  52688=>"110011100",
  52689=>"011110011",
  52690=>"100001111",
  52691=>"010000011",
  52692=>"111011101",
  52693=>"010101111",
  52694=>"000000110",
  52695=>"110011010",
  52696=>"011110111",
  52697=>"110000111",
  52698=>"111100001",
  52699=>"001010000",
  52700=>"000111100",
  52701=>"000001100",
  52702=>"000100011",
  52703=>"000001101",
  52704=>"011110110",
  52705=>"011110010",
  52706=>"100000111",
  52707=>"101000100",
  52708=>"010000011",
  52709=>"000111000",
  52710=>"011000101",
  52711=>"011010101",
  52712=>"111100011",
  52713=>"101101111",
  52714=>"101011001",
  52715=>"101100011",
  52716=>"010010011",
  52717=>"110011000",
  52718=>"011001111",
  52719=>"100010111",
  52720=>"111111011",
  52721=>"101100010",
  52722=>"101101101",
  52723=>"110011010",
  52724=>"010101100",
  52725=>"111110100",
  52726=>"111110000",
  52727=>"111001111",
  52728=>"010011000",
  52729=>"100110010",
  52730=>"111000010",
  52731=>"000011000",
  52732=>"001110111",
  52733=>"001110000",
  52734=>"000111110",
  52735=>"010011010",
  52736=>"000010101",
  52737=>"000010000",
  52738=>"110010110",
  52739=>"001100110",
  52740=>"101111101",
  52741=>"100111011",
  52742=>"100110101",
  52743=>"000011110",
  52744=>"110000010",
  52745=>"001111010",
  52746=>"111011111",
  52747=>"010000000",
  52748=>"010000110",
  52749=>"100011000",
  52750=>"000101111",
  52751=>"110100000",
  52752=>"110110110",
  52753=>"111001100",
  52754=>"000000101",
  52755=>"101110010",
  52756=>"001101110",
  52757=>"000000011",
  52758=>"100001111",
  52759=>"010001000",
  52760=>"001010000",
  52761=>"100001001",
  52762=>"111001001",
  52763=>"010110110",
  52764=>"011000000",
  52765=>"111010011",
  52766=>"000011100",
  52767=>"000110011",
  52768=>"000101011",
  52769=>"011100001",
  52770=>"110000010",
  52771=>"101110101",
  52772=>"110100010",
  52773=>"010011001",
  52774=>"110101100",
  52775=>"010110100",
  52776=>"100000010",
  52777=>"000111000",
  52778=>"100100011",
  52779=>"110010110",
  52780=>"001001000",
  52781=>"010000000",
  52782=>"110111011",
  52783=>"100101110",
  52784=>"101000001",
  52785=>"010101100",
  52786=>"100010011",
  52787=>"001011011",
  52788=>"110110100",
  52789=>"010001001",
  52790=>"100000100",
  52791=>"001001110",
  52792=>"100110011",
  52793=>"100000110",
  52794=>"110101101",
  52795=>"001111010",
  52796=>"011100111",
  52797=>"101000000",
  52798=>"111111010",
  52799=>"110111100",
  52800=>"100100001",
  52801=>"001101000",
  52802=>"011101100",
  52803=>"001001011",
  52804=>"110001010",
  52805=>"111010100",
  52806=>"011001110",
  52807=>"000000110",
  52808=>"000100001",
  52809=>"100000110",
  52810=>"110100011",
  52811=>"110011011",
  52812=>"000011111",
  52813=>"011101100",
  52814=>"111000000",
  52815=>"111111001",
  52816=>"111100010",
  52817=>"010001100",
  52818=>"100100101",
  52819=>"100011101",
  52820=>"110010101",
  52821=>"111110111",
  52822=>"100000010",
  52823=>"111011111",
  52824=>"011101101",
  52825=>"010010100",
  52826=>"001010001",
  52827=>"101000000",
  52828=>"001011001",
  52829=>"111110101",
  52830=>"011011110",
  52831=>"010101111",
  52832=>"111001100",
  52833=>"010110000",
  52834=>"100100101",
  52835=>"010100001",
  52836=>"001101001",
  52837=>"001101010",
  52838=>"000010111",
  52839=>"000111101",
  52840=>"001000100",
  52841=>"110011100",
  52842=>"010101010",
  52843=>"110101100",
  52844=>"011001111",
  52845=>"101001010",
  52846=>"001000101",
  52847=>"010101110",
  52848=>"101011111",
  52849=>"001001110",
  52850=>"010100010",
  52851=>"110101011",
  52852=>"111100001",
  52853=>"111110010",
  52854=>"110111000",
  52855=>"101100011",
  52856=>"111011111",
  52857=>"110101100",
  52858=>"111110100",
  52859=>"010101101",
  52860=>"010000000",
  52861=>"000111010",
  52862=>"101111111",
  52863=>"100010110",
  52864=>"100011000",
  52865=>"010001011",
  52866=>"010110011",
  52867=>"001000011",
  52868=>"100000111",
  52869=>"100010101",
  52870=>"111101110",
  52871=>"110010111",
  52872=>"111000011",
  52873=>"000101111",
  52874=>"010011000",
  52875=>"110111110",
  52876=>"101010111",
  52877=>"000001110",
  52878=>"111110111",
  52879=>"001100111",
  52880=>"100010011",
  52881=>"100010100",
  52882=>"001000110",
  52883=>"111100101",
  52884=>"011111110",
  52885=>"011000100",
  52886=>"110010111",
  52887=>"001101000",
  52888=>"110110100",
  52889=>"100000010",
  52890=>"111010001",
  52891=>"111001111",
  52892=>"011111011",
  52893=>"110001111",
  52894=>"011110100",
  52895=>"000000111",
  52896=>"000010111",
  52897=>"010011111",
  52898=>"001110010",
  52899=>"010100000",
  52900=>"010100101",
  52901=>"111111011",
  52902=>"011101011",
  52903=>"011111000",
  52904=>"001010101",
  52905=>"000110110",
  52906=>"011001101",
  52907=>"110010110",
  52908=>"000000000",
  52909=>"001101111",
  52910=>"000000001",
  52911=>"101110111",
  52912=>"000110111",
  52913=>"100101111",
  52914=>"001010101",
  52915=>"101111101",
  52916=>"110010001",
  52917=>"001001110",
  52918=>"101000001",
  52919=>"100111100",
  52920=>"011111010",
  52921=>"100011001",
  52922=>"001101111",
  52923=>"000010111",
  52924=>"011011001",
  52925=>"100100001",
  52926=>"101011010",
  52927=>"010010100",
  52928=>"100100110",
  52929=>"001001001",
  52930=>"111010000",
  52931=>"100110101",
  52932=>"001101010",
  52933=>"011000110",
  52934=>"101101011",
  52935=>"101000001",
  52936=>"011010011",
  52937=>"101100110",
  52938=>"001110101",
  52939=>"011110011",
  52940=>"011000000",
  52941=>"010100101",
  52942=>"110111010",
  52943=>"111101011",
  52944=>"000000100",
  52945=>"110100110",
  52946=>"001001010",
  52947=>"000010010",
  52948=>"011000111",
  52949=>"000011000",
  52950=>"011011010",
  52951=>"101101010",
  52952=>"111010100",
  52953=>"001100011",
  52954=>"011101100",
  52955=>"110011011",
  52956=>"001111111",
  52957=>"101111000",
  52958=>"010001000",
  52959=>"000101110",
  52960=>"001000010",
  52961=>"101101100",
  52962=>"011110110",
  52963=>"100110010",
  52964=>"110100011",
  52965=>"000111000",
  52966=>"000110111",
  52967=>"101111110",
  52968=>"101110100",
  52969=>"001111101",
  52970=>"010110000",
  52971=>"010010101",
  52972=>"010011100",
  52973=>"000101001",
  52974=>"011111101",
  52975=>"010010010",
  52976=>"111011110",
  52977=>"101001100",
  52978=>"111101111",
  52979=>"100001101",
  52980=>"101011110",
  52981=>"110010110",
  52982=>"111110100",
  52983=>"101101010",
  52984=>"001000101",
  52985=>"110011111",
  52986=>"010001011",
  52987=>"000001001",
  52988=>"001111101",
  52989=>"100101101",
  52990=>"001011000",
  52991=>"001001101",
  52992=>"111001000",
  52993=>"111100101",
  52994=>"111101000",
  52995=>"011111110",
  52996=>"100101110",
  52997=>"000010010",
  52998=>"000000101",
  52999=>"011011001",
  53000=>"011001111",
  53001=>"001000111",
  53002=>"001111100",
  53003=>"000011100",
  53004=>"001001000",
  53005=>"001100001",
  53006=>"011000101",
  53007=>"010010010",
  53008=>"001010101",
  53009=>"101001010",
  53010=>"000010011",
  53011=>"101101100",
  53012=>"101000011",
  53013=>"101110011",
  53014=>"000010011",
  53015=>"100001101",
  53016=>"011011000",
  53017=>"100010100",
  53018=>"001000010",
  53019=>"111110010",
  53020=>"100001001",
  53021=>"100111011",
  53022=>"010001001",
  53023=>"011100010",
  53024=>"011101110",
  53025=>"011110001",
  53026=>"000011101",
  53027=>"011010010",
  53028=>"001010100",
  53029=>"000001011",
  53030=>"110111000",
  53031=>"001100011",
  53032=>"111111100",
  53033=>"000000001",
  53034=>"001110000",
  53035=>"110101111",
  53036=>"101000101",
  53037=>"111000000",
  53038=>"001000010",
  53039=>"010101111",
  53040=>"000101110",
  53041=>"001010100",
  53042=>"001111100",
  53043=>"011100111",
  53044=>"101101011",
  53045=>"111110101",
  53046=>"011011111",
  53047=>"101111011",
  53048=>"001110111",
  53049=>"001111101",
  53050=>"001100111",
  53051=>"011001100",
  53052=>"111000111",
  53053=>"001101111",
  53054=>"000010010",
  53055=>"110010000",
  53056=>"011000110",
  53057=>"010100010",
  53058=>"111101010",
  53059=>"011011001",
  53060=>"110001101",
  53061=>"001010001",
  53062=>"100010100",
  53063=>"100000001",
  53064=>"010010111",
  53065=>"010011110",
  53066=>"101000000",
  53067=>"010000100",
  53068=>"101111101",
  53069=>"110011010",
  53070=>"001000100",
  53071=>"101010011",
  53072=>"001101111",
  53073=>"010101001",
  53074=>"000100100",
  53075=>"001100011",
  53076=>"001010000",
  53077=>"101110100",
  53078=>"010011001",
  53079=>"111010001",
  53080=>"000100100",
  53081=>"100000011",
  53082=>"110101010",
  53083=>"011001001",
  53084=>"001011010",
  53085=>"001000111",
  53086=>"011101100",
  53087=>"000001111",
  53088=>"110100001",
  53089=>"000110110",
  53090=>"101110110",
  53091=>"011111111",
  53092=>"000101000",
  53093=>"001100001",
  53094=>"001101110",
  53095=>"111110010",
  53096=>"100010010",
  53097=>"010001001",
  53098=>"101111100",
  53099=>"101010100",
  53100=>"001000100",
  53101=>"010000001",
  53102=>"101110101",
  53103=>"010010101",
  53104=>"010000101",
  53105=>"000010010",
  53106=>"000011011",
  53107=>"011101111",
  53108=>"001010010",
  53109=>"011100101",
  53110=>"101010010",
  53111=>"101010000",
  53112=>"111111101",
  53113=>"001100111",
  53114=>"111100111",
  53115=>"010000011",
  53116=>"111111000",
  53117=>"010001000",
  53118=>"000001001",
  53119=>"000000001",
  53120=>"011100111",
  53121=>"110110110",
  53122=>"001001100",
  53123=>"010010111",
  53124=>"101110110",
  53125=>"110000001",
  53126=>"101100000",
  53127=>"001010010",
  53128=>"110111010",
  53129=>"010101001",
  53130=>"100110101",
  53131=>"000101110",
  53132=>"000110000",
  53133=>"001000100",
  53134=>"000101011",
  53135=>"101000111",
  53136=>"100001000",
  53137=>"110100111",
  53138=>"001011001",
  53139=>"011011101",
  53140=>"010001110",
  53141=>"011001010",
  53142=>"100100010",
  53143=>"000111101",
  53144=>"111100000",
  53145=>"010111000",
  53146=>"111110010",
  53147=>"010100101",
  53148=>"110001111",
  53149=>"000010011",
  53150=>"101101101",
  53151=>"011001101",
  53152=>"101000010",
  53153=>"101100111",
  53154=>"111100111",
  53155=>"000001011",
  53156=>"000001010",
  53157=>"111101011",
  53158=>"111001110",
  53159=>"111100110",
  53160=>"000011010",
  53161=>"011010000",
  53162=>"000011000",
  53163=>"001011100",
  53164=>"000000011",
  53165=>"100000000",
  53166=>"001000111",
  53167=>"101010010",
  53168=>"001010101",
  53169=>"101000011",
  53170=>"111000001",
  53171=>"111101101",
  53172=>"111110101",
  53173=>"111000011",
  53174=>"011110001",
  53175=>"000101111",
  53176=>"001010101",
  53177=>"010111001",
  53178=>"111110110",
  53179=>"001010011",
  53180=>"111111000",
  53181=>"100001011",
  53182=>"000011001",
  53183=>"000001010",
  53184=>"011000101",
  53185=>"100101111",
  53186=>"110011100",
  53187=>"000110101",
  53188=>"101110001",
  53189=>"100100000",
  53190=>"110001001",
  53191=>"111011001",
  53192=>"000000100",
  53193=>"101001001",
  53194=>"000011001",
  53195=>"100111100",
  53196=>"010111010",
  53197=>"100001111",
  53198=>"111010010",
  53199=>"100111011",
  53200=>"000011001",
  53201=>"011110011",
  53202=>"111111010",
  53203=>"100000000",
  53204=>"111111000",
  53205=>"001111011",
  53206=>"000000110",
  53207=>"001001000",
  53208=>"010010001",
  53209=>"100011010",
  53210=>"100000011",
  53211=>"101000001",
  53212=>"110001100",
  53213=>"001000011",
  53214=>"111011001",
  53215=>"000011001",
  53216=>"010001010",
  53217=>"010000111",
  53218=>"011000010",
  53219=>"000000011",
  53220=>"000111100",
  53221=>"010001011",
  53222=>"000100000",
  53223=>"010011001",
  53224=>"001001111",
  53225=>"111001110",
  53226=>"110000001",
  53227=>"000100101",
  53228=>"010000100",
  53229=>"001011011",
  53230=>"001101100",
  53231=>"000010110",
  53232=>"001011001",
  53233=>"101101000",
  53234=>"000101010",
  53235=>"110111110",
  53236=>"101000111",
  53237=>"110100001",
  53238=>"100010111",
  53239=>"011100010",
  53240=>"001001010",
  53241=>"100101000",
  53242=>"010011001",
  53243=>"011000110",
  53244=>"100110100",
  53245=>"011111100",
  53246=>"001110111",
  53247=>"011001111",
  53248=>"111011011",
  53249=>"011110100",
  53250=>"000101111",
  53251=>"001010100",
  53252=>"011110101",
  53253=>"110010111",
  53254=>"100100010",
  53255=>"111101101",
  53256=>"001111100",
  53257=>"101000100",
  53258=>"001011010",
  53259=>"010110100",
  53260=>"000001000",
  53261=>"000101100",
  53262=>"110111110",
  53263=>"001000110",
  53264=>"101011110",
  53265=>"000010100",
  53266=>"101010001",
  53267=>"000101000",
  53268=>"011010101",
  53269=>"100111110",
  53270=>"111001111",
  53271=>"000101011",
  53272=>"111011000",
  53273=>"001110001",
  53274=>"010000011",
  53275=>"001100111",
  53276=>"000111000",
  53277=>"111010000",
  53278=>"100000001",
  53279=>"111100101",
  53280=>"110001101",
  53281=>"010110101",
  53282=>"111101111",
  53283=>"111100100",
  53284=>"101101110",
  53285=>"001100101",
  53286=>"010100011",
  53287=>"000100011",
  53288=>"110011101",
  53289=>"001101011",
  53290=>"111110100",
  53291=>"011110010",
  53292=>"111111010",
  53293=>"011101000",
  53294=>"101101100",
  53295=>"000001111",
  53296=>"111110101",
  53297=>"110100111",
  53298=>"010001110",
  53299=>"111001101",
  53300=>"100101110",
  53301=>"101000010",
  53302=>"001101101",
  53303=>"010010011",
  53304=>"000001110",
  53305=>"101110101",
  53306=>"001001011",
  53307=>"110000001",
  53308=>"011011000",
  53309=>"101011110",
  53310=>"101101100",
  53311=>"000000101",
  53312=>"000011010",
  53313=>"111000000",
  53314=>"101010110",
  53315=>"100101001",
  53316=>"101011001",
  53317=>"001001001",
  53318=>"011110011",
  53319=>"011111111",
  53320=>"001100010",
  53321=>"101011111",
  53322=>"011011011",
  53323=>"100111111",
  53324=>"001111011",
  53325=>"110101101",
  53326=>"101000000",
  53327=>"111111100",
  53328=>"000100011",
  53329=>"111111110",
  53330=>"100100101",
  53331=>"010111011",
  53332=>"111011110",
  53333=>"100110010",
  53334=>"000011111",
  53335=>"111001001",
  53336=>"101111111",
  53337=>"110001110",
  53338=>"011001011",
  53339=>"100100010",
  53340=>"100101001",
  53341=>"110100000",
  53342=>"101100100",
  53343=>"000001110",
  53344=>"011011101",
  53345=>"101100101",
  53346=>"011100000",
  53347=>"110011101",
  53348=>"110101001",
  53349=>"001111101",
  53350=>"100101111",
  53351=>"100111110",
  53352=>"000011010",
  53353=>"110111011",
  53354=>"101101101",
  53355=>"001110010",
  53356=>"110111110",
  53357=>"111110000",
  53358=>"001001000",
  53359=>"100110101",
  53360=>"111100011",
  53361=>"110110111",
  53362=>"001100101",
  53363=>"001010110",
  53364=>"001000100",
  53365=>"000101111",
  53366=>"000110011",
  53367=>"000101010",
  53368=>"011011110",
  53369=>"000111101",
  53370=>"111100010",
  53371=>"100001000",
  53372=>"101000001",
  53373=>"101010100",
  53374=>"010000010",
  53375=>"110110100",
  53376=>"001101010",
  53377=>"010111100",
  53378=>"000110100",
  53379=>"100000100",
  53380=>"010101001",
  53381=>"100010101",
  53382=>"000101100",
  53383=>"001111110",
  53384=>"011011000",
  53385=>"001011001",
  53386=>"010100010",
  53387=>"000011101",
  53388=>"100011110",
  53389=>"000010000",
  53390=>"111001011",
  53391=>"111100111",
  53392=>"001010111",
  53393=>"000100000",
  53394=>"000101100",
  53395=>"011100111",
  53396=>"001111000",
  53397=>"100001000",
  53398=>"110001100",
  53399=>"111110011",
  53400=>"001011010",
  53401=>"010110110",
  53402=>"110110010",
  53403=>"111010001",
  53404=>"010000111",
  53405=>"101011000",
  53406=>"110101011",
  53407=>"110011110",
  53408=>"101000001",
  53409=>"111100111",
  53410=>"001010000",
  53411=>"010101011",
  53412=>"111110001",
  53413=>"010001100",
  53414=>"011100111",
  53415=>"110001001",
  53416=>"101000011",
  53417=>"010101011",
  53418=>"110010001",
  53419=>"001100101",
  53420=>"011100111",
  53421=>"111000100",
  53422=>"100110000",
  53423=>"111011111",
  53424=>"100010101",
  53425=>"010001100",
  53426=>"111000000",
  53427=>"111110010",
  53428=>"010011000",
  53429=>"011110010",
  53430=>"000100110",
  53431=>"010001011",
  53432=>"000001110",
  53433=>"110000100",
  53434=>"000100101",
  53435=>"010110100",
  53436=>"101110111",
  53437=>"110010001",
  53438=>"000111101",
  53439=>"000100100",
  53440=>"010111011",
  53441=>"100000000",
  53442=>"000000011",
  53443=>"110111111",
  53444=>"111111011",
  53445=>"000010111",
  53446=>"000011001",
  53447=>"010101000",
  53448=>"101110111",
  53449=>"111001100",
  53450=>"111010001",
  53451=>"101110101",
  53452=>"101111101",
  53453=>"010101010",
  53454=>"010001010",
  53455=>"111111001",
  53456=>"011110101",
  53457=>"011000000",
  53458=>"011100000",
  53459=>"111011011",
  53460=>"110101011",
  53461=>"100001011",
  53462=>"110011001",
  53463=>"111110110",
  53464=>"010000001",
  53465=>"101111101",
  53466=>"001001010",
  53467=>"111001000",
  53468=>"111010101",
  53469=>"111010101",
  53470=>"100110100",
  53471=>"001110100",
  53472=>"100010010",
  53473=>"100111111",
  53474=>"100001100",
  53475=>"011001100",
  53476=>"000011101",
  53477=>"010010101",
  53478=>"111000111",
  53479=>"010100111",
  53480=>"000000010",
  53481=>"110000011",
  53482=>"000100110",
  53483=>"110100101",
  53484=>"000010001",
  53485=>"000110001",
  53486=>"000000010",
  53487=>"110010010",
  53488=>"000010001",
  53489=>"110010000",
  53490=>"100000110",
  53491=>"110000001",
  53492=>"110101100",
  53493=>"000110001",
  53494=>"011111111",
  53495=>"100011100",
  53496=>"001111000",
  53497=>"111101000",
  53498=>"000010010",
  53499=>"001010011",
  53500=>"100000111",
  53501=>"001000100",
  53502=>"110010100",
  53503=>"010011111",
  53504=>"000101111",
  53505=>"100001011",
  53506=>"110011110",
  53507=>"000101000",
  53508=>"100111100",
  53509=>"101100111",
  53510=>"001001000",
  53511=>"001101101",
  53512=>"000011000",
  53513=>"001000100",
  53514=>"001110101",
  53515=>"000110110",
  53516=>"010100110",
  53517=>"000001000",
  53518=>"111010010",
  53519=>"000101100",
  53520=>"000010100",
  53521=>"101100111",
  53522=>"000111100",
  53523=>"000110001",
  53524=>"111101100",
  53525=>"011010111",
  53526=>"111110101",
  53527=>"000100000",
  53528=>"001001001",
  53529=>"001111110",
  53530=>"100111101",
  53531=>"010110000",
  53532=>"001001000",
  53533=>"111110010",
  53534=>"010010000",
  53535=>"000100011",
  53536=>"001001000",
  53537=>"000011110",
  53538=>"000100101",
  53539=>"010011010",
  53540=>"110001010",
  53541=>"101110001",
  53542=>"101010100",
  53543=>"100111100",
  53544=>"001010011",
  53545=>"000111111",
  53546=>"011000100",
  53547=>"000010010",
  53548=>"001010110",
  53549=>"000111100",
  53550=>"100110101",
  53551=>"000001000",
  53552=>"110100100",
  53553=>"110111110",
  53554=>"100000111",
  53555=>"011101100",
  53556=>"010010100",
  53557=>"010000100",
  53558=>"000110010",
  53559=>"111110101",
  53560=>"001001110",
  53561=>"100001000",
  53562=>"000110010",
  53563=>"111111110",
  53564=>"011100011",
  53565=>"101100100",
  53566=>"011010001",
  53567=>"111100011",
  53568=>"110000100",
  53569=>"000100011",
  53570=>"100000010",
  53571=>"000111110",
  53572=>"011101101",
  53573=>"110100111",
  53574=>"111001001",
  53575=>"001001001",
  53576=>"110110000",
  53577=>"110010001",
  53578=>"011111000",
  53579=>"000100101",
  53580=>"101011000",
  53581=>"001000101",
  53582=>"100111000",
  53583=>"001001101",
  53584=>"111000100",
  53585=>"100111110",
  53586=>"101001111",
  53587=>"101011110",
  53588=>"110001110",
  53589=>"010100011",
  53590=>"100000000",
  53591=>"000001111",
  53592=>"000110011",
  53593=>"010010100",
  53594=>"010011110",
  53595=>"001010111",
  53596=>"001010100",
  53597=>"110111001",
  53598=>"010000001",
  53599=>"101001111",
  53600=>"001101110",
  53601=>"101000110",
  53602=>"001101101",
  53603=>"111000010",
  53604=>"110010000",
  53605=>"001000101",
  53606=>"101001010",
  53607=>"100100111",
  53608=>"100011000",
  53609=>"110011011",
  53610=>"011101101",
  53611=>"100110001",
  53612=>"111000110",
  53613=>"001011100",
  53614=>"000100100",
  53615=>"010111010",
  53616=>"101100110",
  53617=>"101001100",
  53618=>"001011111",
  53619=>"100110111",
  53620=>"000010111",
  53621=>"100010100",
  53622=>"001111011",
  53623=>"000001000",
  53624=>"000110010",
  53625=>"111110011",
  53626=>"100010010",
  53627=>"001101101",
  53628=>"001110100",
  53629=>"110110001",
  53630=>"010101001",
  53631=>"000100000",
  53632=>"101100101",
  53633=>"100101010",
  53634=>"000000011",
  53635=>"000110111",
  53636=>"101101110",
  53637=>"101100100",
  53638=>"100111111",
  53639=>"000110100",
  53640=>"010000000",
  53641=>"010110000",
  53642=>"101010001",
  53643=>"110000001",
  53644=>"001010110",
  53645=>"011110100",
  53646=>"110001000",
  53647=>"110011101",
  53648=>"000110001",
  53649=>"101010001",
  53650=>"000011001",
  53651=>"000110101",
  53652=>"110000000",
  53653=>"001100011",
  53654=>"010100111",
  53655=>"011101010",
  53656=>"000100101",
  53657=>"110100100",
  53658=>"001001101",
  53659=>"000111010",
  53660=>"001100110",
  53661=>"111010101",
  53662=>"001110001",
  53663=>"000001011",
  53664=>"010100000",
  53665=>"100001000",
  53666=>"111011110",
  53667=>"111000001",
  53668=>"110100011",
  53669=>"010100000",
  53670=>"000110111",
  53671=>"101110011",
  53672=>"100101010",
  53673=>"001001010",
  53674=>"001001001",
  53675=>"101111101",
  53676=>"000101010",
  53677=>"011010000",
  53678=>"011111110",
  53679=>"000010111",
  53680=>"100100100",
  53681=>"011010111",
  53682=>"000101000",
  53683=>"001011111",
  53684=>"100000111",
  53685=>"110100001",
  53686=>"111000101",
  53687=>"101000101",
  53688=>"101110111",
  53689=>"010111101",
  53690=>"100010001",
  53691=>"100000110",
  53692=>"011101110",
  53693=>"100000000",
  53694=>"111001111",
  53695=>"101001101",
  53696=>"000010111",
  53697=>"001101001",
  53698=>"101100101",
  53699=>"011101001",
  53700=>"010000011",
  53701=>"110110100",
  53702=>"111011111",
  53703=>"111111100",
  53704=>"011011001",
  53705=>"101011011",
  53706=>"111111000",
  53707=>"000011000",
  53708=>"100000011",
  53709=>"111101111",
  53710=>"111000000",
  53711=>"010101110",
  53712=>"101101000",
  53713=>"011011111",
  53714=>"100010001",
  53715=>"001001011",
  53716=>"100100100",
  53717=>"001000010",
  53718=>"101101011",
  53719=>"111010100",
  53720=>"100100111",
  53721=>"110000010",
  53722=>"111101110",
  53723=>"111011101",
  53724=>"110011010",
  53725=>"011011010",
  53726=>"000001000",
  53727=>"011011010",
  53728=>"010000010",
  53729=>"101000010",
  53730=>"010110001",
  53731=>"011010101",
  53732=>"001000111",
  53733=>"000010101",
  53734=>"010011101",
  53735=>"000101100",
  53736=>"001001010",
  53737=>"011101101",
  53738=>"111110011",
  53739=>"101100101",
  53740=>"111001011",
  53741=>"111000000",
  53742=>"000101100",
  53743=>"110000110",
  53744=>"010100111",
  53745=>"010101111",
  53746=>"111100011",
  53747=>"011100000",
  53748=>"011011001",
  53749=>"101100010",
  53750=>"100100000",
  53751=>"100100101",
  53752=>"011110000",
  53753=>"110000001",
  53754=>"101010111",
  53755=>"100001010",
  53756=>"101110010",
  53757=>"100111100",
  53758=>"101001110",
  53759=>"110000111",
  53760=>"101011111",
  53761=>"001110100",
  53762=>"111110110",
  53763=>"000100110",
  53764=>"001111001",
  53765=>"110100111",
  53766=>"110011000",
  53767=>"101001000",
  53768=>"010100000",
  53769=>"011111110",
  53770=>"001101010",
  53771=>"010000000",
  53772=>"100100110",
  53773=>"011100010",
  53774=>"100100111",
  53775=>"000111011",
  53776=>"111111101",
  53777=>"111000100",
  53778=>"101010101",
  53779=>"011000100",
  53780=>"011010001",
  53781=>"010110100",
  53782=>"100110011",
  53783=>"001011101",
  53784=>"001000000",
  53785=>"110110011",
  53786=>"010101101",
  53787=>"000111100",
  53788=>"111110100",
  53789=>"001010111",
  53790=>"100111101",
  53791=>"100111010",
  53792=>"111111101",
  53793=>"010110011",
  53794=>"000000001",
  53795=>"110001101",
  53796=>"110001000",
  53797=>"000011110",
  53798=>"011011000",
  53799=>"111001111",
  53800=>"111110000",
  53801=>"011001100",
  53802=>"101010101",
  53803=>"010100100",
  53804=>"000011101",
  53805=>"111110010",
  53806=>"111111011",
  53807=>"000011110",
  53808=>"011000000",
  53809=>"111110110",
  53810=>"011100101",
  53811=>"110100101",
  53812=>"100101111",
  53813=>"010010110",
  53814=>"100100001",
  53815=>"010100001",
  53816=>"011110011",
  53817=>"111110000",
  53818=>"100110110",
  53819=>"011110100",
  53820=>"000111010",
  53821=>"001011110",
  53822=>"101010111",
  53823=>"000001011",
  53824=>"011101011",
  53825=>"110000110",
  53826=>"000001011",
  53827=>"011100010",
  53828=>"110011010",
  53829=>"110101000",
  53830=>"011111111",
  53831=>"010110111",
  53832=>"101010000",
  53833=>"111110011",
  53834=>"000100110",
  53835=>"110010011",
  53836=>"010100010",
  53837=>"001001100",
  53838=>"011001010",
  53839=>"010001001",
  53840=>"111101110",
  53841=>"010010000",
  53842=>"010110110",
  53843=>"101100000",
  53844=>"010001011",
  53845=>"100000101",
  53846=>"101010000",
  53847=>"011011000",
  53848=>"111100111",
  53849=>"001011101",
  53850=>"100011011",
  53851=>"101100001",
  53852=>"111111011",
  53853=>"011111000",
  53854=>"100100010",
  53855=>"110111101",
  53856=>"011001000",
  53857=>"000001111",
  53858=>"001110111",
  53859=>"110100101",
  53860=>"011101110",
  53861=>"101111111",
  53862=>"010010100",
  53863=>"111101111",
  53864=>"000000001",
  53865=>"010011010",
  53866=>"001101110",
  53867=>"101010100",
  53868=>"111110011",
  53869=>"001010101",
  53870=>"010101111",
  53871=>"101000100",
  53872=>"010110101",
  53873=>"110000111",
  53874=>"000010101",
  53875=>"010010010",
  53876=>"110110010",
  53877=>"010000100",
  53878=>"110010000",
  53879=>"110011000",
  53880=>"101110111",
  53881=>"011000101",
  53882=>"111110011",
  53883=>"100100100",
  53884=>"000101101",
  53885=>"010111110",
  53886=>"111001100",
  53887=>"001010110",
  53888=>"101000000",
  53889=>"011011001",
  53890=>"111101111",
  53891=>"100100111",
  53892=>"000001100",
  53893=>"010000100",
  53894=>"111100101",
  53895=>"000001001",
  53896=>"000000011",
  53897=>"111100010",
  53898=>"000000101",
  53899=>"011011110",
  53900=>"001110101",
  53901=>"111001111",
  53902=>"000110111",
  53903=>"011110011",
  53904=>"100000001",
  53905=>"011101011",
  53906=>"001010000",
  53907=>"110000101",
  53908=>"101111001",
  53909=>"010111001",
  53910=>"111011001",
  53911=>"100001000",
  53912=>"001110000",
  53913=>"011001001",
  53914=>"110110110",
  53915=>"001100111",
  53916=>"111110001",
  53917=>"000010010",
  53918=>"000110011",
  53919=>"011010111",
  53920=>"000000000",
  53921=>"011110010",
  53922=>"110101001",
  53923=>"100010011",
  53924=>"100111100",
  53925=>"111010001",
  53926=>"101010101",
  53927=>"010101100",
  53928=>"011110010",
  53929=>"110001010",
  53930=>"011110001",
  53931=>"101011100",
  53932=>"001001010",
  53933=>"011000000",
  53934=>"100001000",
  53935=>"100001000",
  53936=>"101101101",
  53937=>"001000011",
  53938=>"111111011",
  53939=>"100011110",
  53940=>"110001011",
  53941=>"010001100",
  53942=>"110101111",
  53943=>"001011001",
  53944=>"111100001",
  53945=>"110011001",
  53946=>"110111110",
  53947=>"110110000",
  53948=>"000000011",
  53949=>"111100001",
  53950=>"101101000",
  53951=>"010011100",
  53952=>"100100110",
  53953=>"111110000",
  53954=>"111110001",
  53955=>"011010100",
  53956=>"010000111",
  53957=>"000011101",
  53958=>"111111110",
  53959=>"111001111",
  53960=>"111110111",
  53961=>"100001100",
  53962=>"110010000",
  53963=>"111101100",
  53964=>"111100110",
  53965=>"100000111",
  53966=>"010101100",
  53967=>"110000111",
  53968=>"010101011",
  53969=>"000010000",
  53970=>"010011010",
  53971=>"111000001",
  53972=>"100101010",
  53973=>"001000110",
  53974=>"111010011",
  53975=>"001000111",
  53976=>"000001010",
  53977=>"111111010",
  53978=>"110100110",
  53979=>"111111111",
  53980=>"101101100",
  53981=>"000111010",
  53982=>"000101010",
  53983=>"110000001",
  53984=>"100000010",
  53985=>"010010001",
  53986=>"000000011",
  53987=>"110010111",
  53988=>"000001111",
  53989=>"001010110",
  53990=>"001011000",
  53991=>"010110001",
  53992=>"001101111",
  53993=>"110101110",
  53994=>"000100000",
  53995=>"101111100",
  53996=>"011101000",
  53997=>"100110001",
  53998=>"110111000",
  53999=>"011100110",
  54000=>"000111010",
  54001=>"000111001",
  54002=>"110001101",
  54003=>"111101001",
  54004=>"000100100",
  54005=>"111000011",
  54006=>"111100111",
  54007=>"101100111",
  54008=>"101110111",
  54009=>"001100100",
  54010=>"011010000",
  54011=>"000101111",
  54012=>"000011111",
  54013=>"101111110",
  54014=>"110000011",
  54015=>"000010011",
  54016=>"110101010",
  54017=>"000001110",
  54018=>"101100010",
  54019=>"100000010",
  54020=>"111111111",
  54021=>"000000000",
  54022=>"110000001",
  54023=>"100011111",
  54024=>"110000010",
  54025=>"001111111",
  54026=>"001110011",
  54027=>"111111001",
  54028=>"100100000",
  54029=>"100000000",
  54030=>"110101010",
  54031=>"111101011",
  54032=>"101001110",
  54033=>"101111010",
  54034=>"111110001",
  54035=>"001110010",
  54036=>"011100001",
  54037=>"001000101",
  54038=>"000010100",
  54039=>"111100111",
  54040=>"111100010",
  54041=>"110111101",
  54042=>"000001001",
  54043=>"000010011",
  54044=>"101110010",
  54045=>"010110111",
  54046=>"011101001",
  54047=>"000011111",
  54048=>"010001110",
  54049=>"110011111",
  54050=>"111001101",
  54051=>"101001011",
  54052=>"001000001",
  54053=>"000000111",
  54054=>"000000001",
  54055=>"000100101",
  54056=>"110110000",
  54057=>"111110100",
  54058=>"010110011",
  54059=>"001100010",
  54060=>"100101100",
  54061=>"000100001",
  54062=>"000101000",
  54063=>"000101111",
  54064=>"101011110",
  54065=>"110100011",
  54066=>"000011010",
  54067=>"010001111",
  54068=>"110100000",
  54069=>"101010110",
  54070=>"111100101",
  54071=>"010101001",
  54072=>"010010001",
  54073=>"010001110",
  54074=>"000101000",
  54075=>"100111110",
  54076=>"011110000",
  54077=>"110000100",
  54078=>"101101110",
  54079=>"011111010",
  54080=>"010110011",
  54081=>"011100010",
  54082=>"111000010",
  54083=>"111001100",
  54084=>"000101110",
  54085=>"110011001",
  54086=>"001101001",
  54087=>"000000101",
  54088=>"111111101",
  54089=>"101110001",
  54090=>"001101110",
  54091=>"010001101",
  54092=>"101110011",
  54093=>"111000011",
  54094=>"010010101",
  54095=>"001110101",
  54096=>"110000110",
  54097=>"111010101",
  54098=>"111111010",
  54099=>"011000111",
  54100=>"110110100",
  54101=>"010110100",
  54102=>"010111100",
  54103=>"011000000",
  54104=>"110100100",
  54105=>"111000010",
  54106=>"011110111",
  54107=>"010101000",
  54108=>"100111010",
  54109=>"100011100",
  54110=>"000100001",
  54111=>"001000001",
  54112=>"111101100",
  54113=>"011111110",
  54114=>"100000001",
  54115=>"000111101",
  54116=>"111101101",
  54117=>"011111011",
  54118=>"100100101",
  54119=>"010101110",
  54120=>"110011000",
  54121=>"110100001",
  54122=>"111000010",
  54123=>"110101011",
  54124=>"000010111",
  54125=>"110100010",
  54126=>"101011010",
  54127=>"011111001",
  54128=>"011011001",
  54129=>"000001001",
  54130=>"011011011",
  54131=>"001010100",
  54132=>"010101011",
  54133=>"000101010",
  54134=>"011101001",
  54135=>"111001101",
  54136=>"000010011",
  54137=>"100001001",
  54138=>"110100000",
  54139=>"110001100",
  54140=>"000000100",
  54141=>"110011100",
  54142=>"111100100",
  54143=>"001100010",
  54144=>"011001100",
  54145=>"110000101",
  54146=>"001011110",
  54147=>"010010001",
  54148=>"000110001",
  54149=>"010100100",
  54150=>"100000010",
  54151=>"000101011",
  54152=>"111100000",
  54153=>"010010011",
  54154=>"000101001",
  54155=>"111101011",
  54156=>"111011010",
  54157=>"100000111",
  54158=>"010011010",
  54159=>"101000111",
  54160=>"101110000",
  54161=>"011001000",
  54162=>"001010111",
  54163=>"101111001",
  54164=>"111111101",
  54165=>"001100000",
  54166=>"110000011",
  54167=>"000111101",
  54168=>"010011000",
  54169=>"001010100",
  54170=>"000100001",
  54171=>"101011010",
  54172=>"000001000",
  54173=>"011011110",
  54174=>"111001111",
  54175=>"100101000",
  54176=>"100000110",
  54177=>"101111000",
  54178=>"001010001",
  54179=>"101101000",
  54180=>"011000000",
  54181=>"010110100",
  54182=>"110001000",
  54183=>"000000000",
  54184=>"001110010",
  54185=>"101000001",
  54186=>"101010011",
  54187=>"010101100",
  54188=>"101111001",
  54189=>"101010001",
  54190=>"000010010",
  54191=>"100010110",
  54192=>"100010100",
  54193=>"100010111",
  54194=>"100011101",
  54195=>"010000010",
  54196=>"011011010",
  54197=>"101101001",
  54198=>"011011110",
  54199=>"010000001",
  54200=>"101100110",
  54201=>"111010010",
  54202=>"101001011",
  54203=>"110111011",
  54204=>"111001110",
  54205=>"011010000",
  54206=>"010101001",
  54207=>"100100100",
  54208=>"000100001",
  54209=>"001000101",
  54210=>"000000101",
  54211=>"110100000",
  54212=>"011100111",
  54213=>"001111101",
  54214=>"110001101",
  54215=>"100000100",
  54216=>"101000000",
  54217=>"110101111",
  54218=>"100100001",
  54219=>"011110110",
  54220=>"101100011",
  54221=>"111100100",
  54222=>"000010001",
  54223=>"011110100",
  54224=>"101100111",
  54225=>"110100110",
  54226=>"110101110",
  54227=>"111101000",
  54228=>"110110111",
  54229=>"010011001",
  54230=>"011001110",
  54231=>"100010011",
  54232=>"010110111",
  54233=>"101011111",
  54234=>"110010110",
  54235=>"101000101",
  54236=>"111000011",
  54237=>"011111010",
  54238=>"100100110",
  54239=>"100000011",
  54240=>"100001100",
  54241=>"010100110",
  54242=>"000110001",
  54243=>"110010100",
  54244=>"111001001",
  54245=>"111100111",
  54246=>"010101110",
  54247=>"101110111",
  54248=>"100010010",
  54249=>"000010111",
  54250=>"000010010",
  54251=>"100110111",
  54252=>"100011010",
  54253=>"000100010",
  54254=>"011100111",
  54255=>"111101110",
  54256=>"010000100",
  54257=>"010010010",
  54258=>"001001010",
  54259=>"011011010",
  54260=>"111010010",
  54261=>"111000000",
  54262=>"000100110",
  54263=>"110101110",
  54264=>"001011010",
  54265=>"011111000",
  54266=>"100011001",
  54267=>"101001011",
  54268=>"111110110",
  54269=>"011111100",
  54270=>"001000100",
  54271=>"111111101",
  54272=>"110100010",
  54273=>"000011010",
  54274=>"010111100",
  54275=>"011100000",
  54276=>"000000110",
  54277=>"000000111",
  54278=>"101110011",
  54279=>"101000010",
  54280=>"100000001",
  54281=>"011010111",
  54282=>"001101100",
  54283=>"111110010",
  54284=>"000110101",
  54285=>"101101001",
  54286=>"011100000",
  54287=>"111111010",
  54288=>"001001110",
  54289=>"000100101",
  54290=>"010001001",
  54291=>"101110010",
  54292=>"001100001",
  54293=>"111000011",
  54294=>"111101000",
  54295=>"010000011",
  54296=>"001110010",
  54297=>"001110111",
  54298=>"001010011",
  54299=>"101101110",
  54300=>"100010110",
  54301=>"001010000",
  54302=>"110110010",
  54303=>"000000100",
  54304=>"000100010",
  54305=>"100101111",
  54306=>"001010100",
  54307=>"001101010",
  54308=>"001110010",
  54309=>"000011100",
  54310=>"000111011",
  54311=>"011001001",
  54312=>"011110000",
  54313=>"011101110",
  54314=>"011111111",
  54315=>"101000000",
  54316=>"100100000",
  54317=>"101101100",
  54318=>"010010101",
  54319=>"001010011",
  54320=>"110110111",
  54321=>"001110011",
  54322=>"110110100",
  54323=>"110100111",
  54324=>"000011001",
  54325=>"011010101",
  54326=>"011010110",
  54327=>"110001111",
  54328=>"100010101",
  54329=>"111011001",
  54330=>"110101011",
  54331=>"100000101",
  54332=>"100010000",
  54333=>"011100001",
  54334=>"101000010",
  54335=>"001100101",
  54336=>"100111111",
  54337=>"101100001",
  54338=>"100001011",
  54339=>"000101001",
  54340=>"100101101",
  54341=>"101000000",
  54342=>"011100010",
  54343=>"010111000",
  54344=>"010111100",
  54345=>"010101000",
  54346=>"001100110",
  54347=>"101001000",
  54348=>"001000110",
  54349=>"101111101",
  54350=>"101100101",
  54351=>"010101010",
  54352=>"101010110",
  54353=>"100101110",
  54354=>"110110010",
  54355=>"110111100",
  54356=>"001010001",
  54357=>"010111101",
  54358=>"101111010",
  54359=>"000100110",
  54360=>"011001010",
  54361=>"000101011",
  54362=>"110101000",
  54363=>"010000101",
  54364=>"111101000",
  54365=>"001101000",
  54366=>"011001111",
  54367=>"010000111",
  54368=>"100101100",
  54369=>"011110011",
  54370=>"111110110",
  54371=>"000000011",
  54372=>"101110001",
  54373=>"111011111",
  54374=>"101110111",
  54375=>"010111000",
  54376=>"101111110",
  54377=>"101110011",
  54378=>"011011110",
  54379=>"111010001",
  54380=>"111011001",
  54381=>"010000100",
  54382=>"000100000",
  54383=>"110001111",
  54384=>"011001101",
  54385=>"011011111",
  54386=>"000010011",
  54387=>"010100100",
  54388=>"001000101",
  54389=>"010010110",
  54390=>"101000101",
  54391=>"101001110",
  54392=>"100111011",
  54393=>"101111100",
  54394=>"000100000",
  54395=>"001000011",
  54396=>"010000010",
  54397=>"101101011",
  54398=>"000010100",
  54399=>"110001010",
  54400=>"000000001",
  54401=>"111110000",
  54402=>"011100111",
  54403=>"110001001",
  54404=>"001000011",
  54405=>"001100111",
  54406=>"010100100",
  54407=>"000001111",
  54408=>"011101111",
  54409=>"011110100",
  54410=>"100010010",
  54411=>"011101111",
  54412=>"001001010",
  54413=>"111100011",
  54414=>"001111000",
  54415=>"111010100",
  54416=>"000111010",
  54417=>"001000011",
  54418=>"101011010",
  54419=>"011001000",
  54420=>"010000001",
  54421=>"101001100",
  54422=>"010100000",
  54423=>"101011101",
  54424=>"101110010",
  54425=>"111011111",
  54426=>"110100110",
  54427=>"000000010",
  54428=>"000100100",
  54429=>"111000001",
  54430=>"001010010",
  54431=>"101010100",
  54432=>"100010101",
  54433=>"110000001",
  54434=>"011111011",
  54435=>"111110011",
  54436=>"101101111",
  54437=>"001110101",
  54438=>"111000011",
  54439=>"100001011",
  54440=>"011110101",
  54441=>"001010100",
  54442=>"011101001",
  54443=>"111110000",
  54444=>"101010110",
  54445=>"011000110",
  54446=>"101110001",
  54447=>"000100110",
  54448=>"110101001",
  54449=>"111101111",
  54450=>"100100101",
  54451=>"010010010",
  54452=>"101111001",
  54453=>"001101110",
  54454=>"010100010",
  54455=>"001110010",
  54456=>"000000100",
  54457=>"000100110",
  54458=>"111001010",
  54459=>"011001100",
  54460=>"100100110",
  54461=>"110011110",
  54462=>"111000111",
  54463=>"100100111",
  54464=>"111000000",
  54465=>"011001110",
  54466=>"011000010",
  54467=>"000100110",
  54468=>"001000000",
  54469=>"000011010",
  54470=>"001100101",
  54471=>"010101001",
  54472=>"011111011",
  54473=>"101001110",
  54474=>"011110001",
  54475=>"111110111",
  54476=>"110011011",
  54477=>"111110000",
  54478=>"001100000",
  54479=>"100011101",
  54480=>"000000101",
  54481=>"001110110",
  54482=>"001110100",
  54483=>"010001101",
  54484=>"100010000",
  54485=>"110101111",
  54486=>"101110011",
  54487=>"101110001",
  54488=>"101111011",
  54489=>"111111010",
  54490=>"110111010",
  54491=>"011101101",
  54492=>"001000011",
  54493=>"100000100",
  54494=>"001010100",
  54495=>"101110010",
  54496=>"010011111",
  54497=>"011011100",
  54498=>"001111001",
  54499=>"000110111",
  54500=>"100101010",
  54501=>"011010010",
  54502=>"001010010",
  54503=>"101101010",
  54504=>"000101111",
  54505=>"000101000",
  54506=>"110110011",
  54507=>"001110101",
  54508=>"010100011",
  54509=>"101010100",
  54510=>"010000110",
  54511=>"101001101",
  54512=>"111001100",
  54513=>"001111110",
  54514=>"000100011",
  54515=>"010010111",
  54516=>"010101010",
  54517=>"111000010",
  54518=>"100111101",
  54519=>"001011011",
  54520=>"100111001",
  54521=>"111011010",
  54522=>"011100101",
  54523=>"010110000",
  54524=>"001110100",
  54525=>"011110101",
  54526=>"101001100",
  54527=>"111001100",
  54528=>"010001011",
  54529=>"110000000",
  54530=>"101101100",
  54531=>"000110011",
  54532=>"000101100",
  54533=>"011110011",
  54534=>"001111111",
  54535=>"011000101",
  54536=>"110010001",
  54537=>"010110101",
  54538=>"001010011",
  54539=>"010100010",
  54540=>"001111011",
  54541=>"001010111",
  54542=>"110010110",
  54543=>"010100100",
  54544=>"001001000",
  54545=>"000101011",
  54546=>"111101111",
  54547=>"011000100",
  54548=>"111001010",
  54549=>"001000110",
  54550=>"110011110",
  54551=>"111101001",
  54552=>"110011101",
  54553=>"011000100",
  54554=>"100101110",
  54555=>"000110101",
  54556=>"111011000",
  54557=>"010000101",
  54558=>"011011101",
  54559=>"001011101",
  54560=>"011101000",
  54561=>"100110101",
  54562=>"011010000",
  54563=>"001110100",
  54564=>"001010011",
  54565=>"101011011",
  54566=>"001101011",
  54567=>"101100110",
  54568=>"001011010",
  54569=>"110000010",
  54570=>"001110110",
  54571=>"111011110",
  54572=>"111011001",
  54573=>"000000010",
  54574=>"000000010",
  54575=>"101101101",
  54576=>"001000110",
  54577=>"001000101",
  54578=>"101110111",
  54579=>"011000000",
  54580=>"111111101",
  54581=>"001000111",
  54582=>"101100000",
  54583=>"001101001",
  54584=>"110101111",
  54585=>"101100010",
  54586=>"010111111",
  54587=>"010111010",
  54588=>"111110111",
  54589=>"110001001",
  54590=>"010010000",
  54591=>"111101011",
  54592=>"000011001",
  54593=>"000011010",
  54594=>"101000110",
  54595=>"110101111",
  54596=>"001000111",
  54597=>"011111110",
  54598=>"110010100",
  54599=>"011001110",
  54600=>"101101101",
  54601=>"111100011",
  54602=>"000110011",
  54603=>"000101111",
  54604=>"000011110",
  54605=>"011011111",
  54606=>"110001111",
  54607=>"001100101",
  54608=>"101100010",
  54609=>"001011001",
  54610=>"010000110",
  54611=>"111100111",
  54612=>"101010010",
  54613=>"110010110",
  54614=>"110011101",
  54615=>"011110101",
  54616=>"011001110",
  54617=>"100001010",
  54618=>"101101001",
  54619=>"101100000",
  54620=>"110010011",
  54621=>"110010111",
  54622=>"101010100",
  54623=>"001101111",
  54624=>"010110110",
  54625=>"001100100",
  54626=>"100000000",
  54627=>"100000000",
  54628=>"001101101",
  54629=>"110110101",
  54630=>"111001000",
  54631=>"100110000",
  54632=>"001001000",
  54633=>"010101100",
  54634=>"101101111",
  54635=>"010111000",
  54636=>"010111010",
  54637=>"010001110",
  54638=>"110001001",
  54639=>"011010000",
  54640=>"001100111",
  54641=>"101111101",
  54642=>"010111111",
  54643=>"101010101",
  54644=>"000011011",
  54645=>"100101111",
  54646=>"101001101",
  54647=>"000110111",
  54648=>"010110001",
  54649=>"000110011",
  54650=>"011010011",
  54651=>"011101000",
  54652=>"011011011",
  54653=>"101111110",
  54654=>"110111010",
  54655=>"000011001",
  54656=>"010110111",
  54657=>"100011000",
  54658=>"011010100",
  54659=>"100000001",
  54660=>"100001101",
  54661=>"001000110",
  54662=>"111101100",
  54663=>"010001011",
  54664=>"000001110",
  54665=>"000001101",
  54666=>"101111001",
  54667=>"111001110",
  54668=>"101110110",
  54669=>"111011000",
  54670=>"001001001",
  54671=>"011011000",
  54672=>"100011111",
  54673=>"110000111",
  54674=>"111111000",
  54675=>"010001000",
  54676=>"000010011",
  54677=>"110000000",
  54678=>"010010101",
  54679=>"011111111",
  54680=>"011000101",
  54681=>"010011101",
  54682=>"110000111",
  54683=>"110110011",
  54684=>"100001101",
  54685=>"101111011",
  54686=>"011110011",
  54687=>"000101101",
  54688=>"100010101",
  54689=>"011010111",
  54690=>"111101001",
  54691=>"111111111",
  54692=>"110101001",
  54693=>"111001101",
  54694=>"111101110",
  54695=>"000101010",
  54696=>"000100111",
  54697=>"000101110",
  54698=>"101011000",
  54699=>"001010100",
  54700=>"110000001",
  54701=>"011011100",
  54702=>"101100111",
  54703=>"001101101",
  54704=>"110010011",
  54705=>"101010111",
  54706=>"000100101",
  54707=>"001011010",
  54708=>"001010011",
  54709=>"011110011",
  54710=>"001111100",
  54711=>"001110101",
  54712=>"101010010",
  54713=>"011001101",
  54714=>"011000010",
  54715=>"110101011",
  54716=>"101110010",
  54717=>"111001011",
  54718=>"111010001",
  54719=>"010101001",
  54720=>"011100110",
  54721=>"011000111",
  54722=>"000101100",
  54723=>"111000111",
  54724=>"010010000",
  54725=>"011001110",
  54726=>"111010100",
  54727=>"000101011",
  54728=>"010001010",
  54729=>"110001111",
  54730=>"100000000",
  54731=>"010111100",
  54732=>"100000111",
  54733=>"000000001",
  54734=>"101000000",
  54735=>"001000101",
  54736=>"101010000",
  54737=>"110101110",
  54738=>"100000100",
  54739=>"000000101",
  54740=>"101011001",
  54741=>"010011110",
  54742=>"011111101",
  54743=>"000010000",
  54744=>"101000110",
  54745=>"011111011",
  54746=>"011101001",
  54747=>"101010101",
  54748=>"011100101",
  54749=>"010101100",
  54750=>"110100010",
  54751=>"101111101",
  54752=>"111011111",
  54753=>"000011100",
  54754=>"011000111",
  54755=>"101000000",
  54756=>"111101010",
  54757=>"011010000",
  54758=>"001001011",
  54759=>"100110111",
  54760=>"011110001",
  54761=>"110100001",
  54762=>"000001111",
  54763=>"100110010",
  54764=>"111111111",
  54765=>"010011101",
  54766=>"010001100",
  54767=>"010000010",
  54768=>"101011111",
  54769=>"011100000",
  54770=>"001101111",
  54771=>"000011011",
  54772=>"100001110",
  54773=>"001101011",
  54774=>"100101011",
  54775=>"110000110",
  54776=>"100010000",
  54777=>"110011100",
  54778=>"011001011",
  54779=>"010101101",
  54780=>"000110100",
  54781=>"101000011",
  54782=>"111110001",
  54783=>"001001010",
  54784=>"111010100",
  54785=>"101000000",
  54786=>"111011110",
  54787=>"110010111",
  54788=>"101110111",
  54789=>"011111011",
  54790=>"011000101",
  54791=>"100110110",
  54792=>"001001010",
  54793=>"111100010",
  54794=>"101011011",
  54795=>"000010001",
  54796=>"110010101",
  54797=>"100011101",
  54798=>"001010001",
  54799=>"010111011",
  54800=>"101000100",
  54801=>"000111101",
  54802=>"111110110",
  54803=>"101010000",
  54804=>"001100011",
  54805=>"110000011",
  54806=>"111101111",
  54807=>"110100100",
  54808=>"100001010",
  54809=>"100111010",
  54810=>"001011000",
  54811=>"100111000",
  54812=>"001011111",
  54813=>"100100111",
  54814=>"000111000",
  54815=>"011111101",
  54816=>"010000001",
  54817=>"010001100",
  54818=>"000000110",
  54819=>"110000101",
  54820=>"010100011",
  54821=>"101110011",
  54822=>"111110001",
  54823=>"110111011",
  54824=>"010111110",
  54825=>"100000001",
  54826=>"010001001",
  54827=>"000010100",
  54828=>"000100011",
  54829=>"111001110",
  54830=>"000011111",
  54831=>"111011000",
  54832=>"111111001",
  54833=>"110000101",
  54834=>"011010010",
  54835=>"001010000",
  54836=>"110000000",
  54837=>"100100011",
  54838=>"001001111",
  54839=>"011000111",
  54840=>"101011111",
  54841=>"101101110",
  54842=>"100000011",
  54843=>"110100010",
  54844=>"101001110",
  54845=>"100000000",
  54846=>"110001100",
  54847=>"001000010",
  54848=>"010001110",
  54849=>"101010101",
  54850=>"101100111",
  54851=>"110011000",
  54852=>"011011011",
  54853=>"111001010",
  54854=>"011101011",
  54855=>"111001110",
  54856=>"110011111",
  54857=>"111101111",
  54858=>"100000101",
  54859=>"000111111",
  54860=>"011011111",
  54861=>"101011110",
  54862=>"011111000",
  54863=>"110100111",
  54864=>"000011110",
  54865=>"100111000",
  54866=>"110110001",
  54867=>"011101001",
  54868=>"100001100",
  54869=>"000110001",
  54870=>"110010111",
  54871=>"001000010",
  54872=>"100001011",
  54873=>"110000100",
  54874=>"001110100",
  54875=>"101001001",
  54876=>"011110100",
  54877=>"000000100",
  54878=>"100011010",
  54879=>"110000101",
  54880=>"000100101",
  54881=>"100000001",
  54882=>"011000101",
  54883=>"100100110",
  54884=>"000000001",
  54885=>"001001001",
  54886=>"100100111",
  54887=>"110011100",
  54888=>"001111100",
  54889=>"001001111",
  54890=>"011100100",
  54891=>"010001111",
  54892=>"111100111",
  54893=>"001010000",
  54894=>"101011100",
  54895=>"100011110",
  54896=>"001000110",
  54897=>"101000011",
  54898=>"001010011",
  54899=>"111100101",
  54900=>"110011111",
  54901=>"100100001",
  54902=>"110110010",
  54903=>"010111000",
  54904=>"100110101",
  54905=>"110100000",
  54906=>"011110111",
  54907=>"100001111",
  54908=>"010000001",
  54909=>"101100100",
  54910=>"010010110",
  54911=>"001110111",
  54912=>"101110011",
  54913=>"111101100",
  54914=>"010001010",
  54915=>"111011001",
  54916=>"010100111",
  54917=>"111011000",
  54918=>"000011100",
  54919=>"000100000",
  54920=>"000000101",
  54921=>"000000110",
  54922=>"111011110",
  54923=>"110111011",
  54924=>"000000010",
  54925=>"111110010",
  54926=>"101111010",
  54927=>"011110101",
  54928=>"100110101",
  54929=>"011001011",
  54930=>"110010010",
  54931=>"110000100",
  54932=>"101110111",
  54933=>"111011000",
  54934=>"000010100",
  54935=>"011001000",
  54936=>"101011000",
  54937=>"101011001",
  54938=>"101001101",
  54939=>"111111001",
  54940=>"001100010",
  54941=>"001011010",
  54942=>"111110110",
  54943=>"010101111",
  54944=>"110000101",
  54945=>"111010101",
  54946=>"011010100",
  54947=>"001001000",
  54948=>"101010001",
  54949=>"011010001",
  54950=>"100000000",
  54951=>"001011001",
  54952=>"001011111",
  54953=>"000010101",
  54954=>"000000010",
  54955=>"000101101",
  54956=>"100011011",
  54957=>"000001100",
  54958=>"000010011",
  54959=>"011111001",
  54960=>"000011000",
  54961=>"010001110",
  54962=>"101000100",
  54963=>"010101000",
  54964=>"111100101",
  54965=>"010000101",
  54966=>"001010111",
  54967=>"010001101",
  54968=>"000000000",
  54969=>"101001010",
  54970=>"101111110",
  54971=>"011001001",
  54972=>"100001110",
  54973=>"111010010",
  54974=>"000010000",
  54975=>"110111010",
  54976=>"111101010",
  54977=>"110000001",
  54978=>"001101010",
  54979=>"000011110",
  54980=>"001011111",
  54981=>"000110101",
  54982=>"001101101",
  54983=>"100111000",
  54984=>"010101010",
  54985=>"000000101",
  54986=>"100110110",
  54987=>"000000100",
  54988=>"100110001",
  54989=>"111001111",
  54990=>"000000100",
  54991=>"101010011",
  54992=>"110011000",
  54993=>"110111110",
  54994=>"010100011",
  54995=>"000000110",
  54996=>"010011000",
  54997=>"000000100",
  54998=>"010001100",
  54999=>"110101001",
  55000=>"100001110",
  55001=>"001111000",
  55002=>"100100000",
  55003=>"101100000",
  55004=>"110010001",
  55005=>"101110010",
  55006=>"111111111",
  55007=>"110111001",
  55008=>"001000101",
  55009=>"001111001",
  55010=>"010110000",
  55011=>"010101001",
  55012=>"001010011",
  55013=>"100100101",
  55014=>"100001011",
  55015=>"110100100",
  55016=>"101100111",
  55017=>"111011111",
  55018=>"011111101",
  55019=>"010011111",
  55020=>"001100010",
  55021=>"000001111",
  55022=>"101011111",
  55023=>"000111011",
  55024=>"100001011",
  55025=>"011101100",
  55026=>"100000000",
  55027=>"110100001",
  55028=>"111101000",
  55029=>"101001010",
  55030=>"111000001",
  55031=>"100000110",
  55032=>"101111101",
  55033=>"111100101",
  55034=>"111000000",
  55035=>"001001111",
  55036=>"111010101",
  55037=>"001101111",
  55038=>"000010110",
  55039=>"000001000",
  55040=>"111001001",
  55041=>"110111010",
  55042=>"100011010",
  55043=>"001100111",
  55044=>"100111000",
  55045=>"100101001",
  55046=>"110001101",
  55047=>"010001000",
  55048=>"011000101",
  55049=>"100100100",
  55050=>"100000111",
  55051=>"011100100",
  55052=>"000101101",
  55053=>"100000011",
  55054=>"111010011",
  55055=>"000100001",
  55056=>"010010000",
  55057=>"111100001",
  55058=>"111011010",
  55059=>"100010110",
  55060=>"001000110",
  55061=>"101110100",
  55062=>"010110000",
  55063=>"111110010",
  55064=>"101011011",
  55065=>"000110111",
  55066=>"000001000",
  55067=>"110001110",
  55068=>"011001001",
  55069=>"110101100",
  55070=>"111000011",
  55071=>"001010011",
  55072=>"111111101",
  55073=>"101111111",
  55074=>"110110000",
  55075=>"111001111",
  55076=>"010000000",
  55077=>"111001101",
  55078=>"000010101",
  55079=>"001100010",
  55080=>"011100111",
  55081=>"001010000",
  55082=>"011011110",
  55083=>"010000011",
  55084=>"001010001",
  55085=>"010100000",
  55086=>"010010100",
  55087=>"100011100",
  55088=>"101111011",
  55089=>"100001001",
  55090=>"101111001",
  55091=>"111000010",
  55092=>"001000000",
  55093=>"011000001",
  55094=>"001101110",
  55095=>"000000110",
  55096=>"011010001",
  55097=>"000001000",
  55098=>"101000000",
  55099=>"001001111",
  55100=>"011000001",
  55101=>"010111001",
  55102=>"000111100",
  55103=>"000111110",
  55104=>"100001110",
  55105=>"000001000",
  55106=>"010100101",
  55107=>"111111010",
  55108=>"111001000",
  55109=>"010000110",
  55110=>"010001100",
  55111=>"101100000",
  55112=>"011010101",
  55113=>"101110011",
  55114=>"011100100",
  55115=>"010010101",
  55116=>"000110011",
  55117=>"110000011",
  55118=>"011111011",
  55119=>"110000011",
  55120=>"101000111",
  55121=>"010101110",
  55122=>"000010010",
  55123=>"001010101",
  55124=>"000100011",
  55125=>"111011011",
  55126=>"001000001",
  55127=>"100000101",
  55128=>"000101111",
  55129=>"111101111",
  55130=>"110110001",
  55131=>"001100000",
  55132=>"011110000",
  55133=>"100100111",
  55134=>"111001000",
  55135=>"110111111",
  55136=>"010110000",
  55137=>"110111111",
  55138=>"011000101",
  55139=>"110011011",
  55140=>"100010000",
  55141=>"011001111",
  55142=>"010110101",
  55143=>"100101000",
  55144=>"111010100",
  55145=>"000001011",
  55146=>"011000110",
  55147=>"000011011",
  55148=>"000101001",
  55149=>"011100000",
  55150=>"000101010",
  55151=>"010101001",
  55152=>"010111001",
  55153=>"010101011",
  55154=>"111110111",
  55155=>"111010111",
  55156=>"100110110",
  55157=>"011011001",
  55158=>"100010000",
  55159=>"000000100",
  55160=>"101111011",
  55161=>"001111001",
  55162=>"000100111",
  55163=>"000010101",
  55164=>"011001011",
  55165=>"001110001",
  55166=>"000000010",
  55167=>"111100100",
  55168=>"010011010",
  55169=>"011101100",
  55170=>"011111011",
  55171=>"000101011",
  55172=>"100110000",
  55173=>"000110101",
  55174=>"111011101",
  55175=>"000001001",
  55176=>"111100011",
  55177=>"111111001",
  55178=>"101110011",
  55179=>"101101101",
  55180=>"000000011",
  55181=>"000111100",
  55182=>"000001110",
  55183=>"100001001",
  55184=>"111101101",
  55185=>"011100000",
  55186=>"000011001",
  55187=>"010000111",
  55188=>"111011010",
  55189=>"010111111",
  55190=>"001000001",
  55191=>"101010000",
  55192=>"000001111",
  55193=>"001010110",
  55194=>"000001011",
  55195=>"101001010",
  55196=>"001010101",
  55197=>"101011100",
  55198=>"101010001",
  55199=>"000001001",
  55200=>"011011110",
  55201=>"111111101",
  55202=>"101010111",
  55203=>"010001100",
  55204=>"100001010",
  55205=>"011101110",
  55206=>"100110010",
  55207=>"010110110",
  55208=>"100001100",
  55209=>"010011000",
  55210=>"110111010",
  55211=>"101111001",
  55212=>"101110110",
  55213=>"000011111",
  55214=>"010100000",
  55215=>"000001100",
  55216=>"011101101",
  55217=>"101010001",
  55218=>"110001101",
  55219=>"101010100",
  55220=>"100111001",
  55221=>"110111111",
  55222=>"110100011",
  55223=>"010010100",
  55224=>"011100111",
  55225=>"101000011",
  55226=>"110010101",
  55227=>"001100000",
  55228=>"001011101",
  55229=>"111000110",
  55230=>"100011000",
  55231=>"001001011",
  55232=>"000001010",
  55233=>"101100110",
  55234=>"010000110",
  55235=>"111100100",
  55236=>"111100101",
  55237=>"100101011",
  55238=>"101110000",
  55239=>"101110100",
  55240=>"000001100",
  55241=>"001110010",
  55242=>"101011111",
  55243=>"100000010",
  55244=>"010000010",
  55245=>"000110111",
  55246=>"111011010",
  55247=>"100101010",
  55248=>"110010000",
  55249=>"010100011",
  55250=>"111000011",
  55251=>"010000000",
  55252=>"010100111",
  55253=>"111001111",
  55254=>"001001100",
  55255=>"001010101",
  55256=>"010100001",
  55257=>"011111011",
  55258=>"111100111",
  55259=>"011011100",
  55260=>"100100011",
  55261=>"001001000",
  55262=>"111001101",
  55263=>"110110001",
  55264=>"111111011",
  55265=>"101100111",
  55266=>"011001011",
  55267=>"110011100",
  55268=>"000100000",
  55269=>"011101110",
  55270=>"011101010",
  55271=>"100000011",
  55272=>"101101100",
  55273=>"101111100",
  55274=>"001101110",
  55275=>"000101000",
  55276=>"011001000",
  55277=>"010001011",
  55278=>"001001011",
  55279=>"101011100",
  55280=>"010110000",
  55281=>"100101001",
  55282=>"111101101",
  55283=>"011010100",
  55284=>"110101001",
  55285=>"110111001",
  55286=>"111001000",
  55287=>"000110101",
  55288=>"010010110",
  55289=>"111100011",
  55290=>"110000111",
  55291=>"011110101",
  55292=>"100100010",
  55293=>"100100101",
  55294=>"000100000",
  55295=>"110011110",
  55296=>"110010100",
  55297=>"000100001",
  55298=>"111111100",
  55299=>"001001110",
  55300=>"101111111",
  55301=>"101001000",
  55302=>"111100110",
  55303=>"001000011",
  55304=>"100100110",
  55305=>"000001000",
  55306=>"001001010",
  55307=>"011010110",
  55308=>"011011000",
  55309=>"011111000",
  55310=>"001011001",
  55311=>"010100011",
  55312=>"110001100",
  55313=>"110011000",
  55314=>"101101001",
  55315=>"000000000",
  55316=>"001111101",
  55317=>"101111010",
  55318=>"110011101",
  55319=>"001100110",
  55320=>"010110000",
  55321=>"001010100",
  55322=>"011110111",
  55323=>"000000011",
  55324=>"000101010",
  55325=>"101000000",
  55326=>"000101101",
  55327=>"011000011",
  55328=>"110011000",
  55329=>"000101010",
  55330=>"010010100",
  55331=>"001101010",
  55332=>"101010111",
  55333=>"110111011",
  55334=>"111110001",
  55335=>"011111111",
  55336=>"100011011",
  55337=>"010100100",
  55338=>"011110111",
  55339=>"101011011",
  55340=>"000000000",
  55341=>"101001100",
  55342=>"111101111",
  55343=>"001101011",
  55344=>"100000010",
  55345=>"000000011",
  55346=>"100001000",
  55347=>"010001010",
  55348=>"000111001",
  55349=>"111110001",
  55350=>"000000110",
  55351=>"001010100",
  55352=>"101100111",
  55353=>"101100100",
  55354=>"111001010",
  55355=>"011100000",
  55356=>"010010001",
  55357=>"111111010",
  55358=>"011101000",
  55359=>"000110101",
  55360=>"000011000",
  55361=>"000011110",
  55362=>"000111111",
  55363=>"101111110",
  55364=>"111010011",
  55365=>"011100111",
  55366=>"110011101",
  55367=>"101010110",
  55368=>"000000010",
  55369=>"000001000",
  55370=>"000110001",
  55371=>"111011000",
  55372=>"001110100",
  55373=>"101111101",
  55374=>"111111111",
  55375=>"001110101",
  55376=>"100010001",
  55377=>"000111111",
  55378=>"100011000",
  55379=>"111011110",
  55380=>"010010010",
  55381=>"011101111",
  55382=>"111100001",
  55383=>"011100101",
  55384=>"011010100",
  55385=>"011001111",
  55386=>"001001100",
  55387=>"000000010",
  55388=>"100000101",
  55389=>"000011100",
  55390=>"100011100",
  55391=>"001100101",
  55392=>"000001101",
  55393=>"101101100",
  55394=>"010101101",
  55395=>"010011011",
  55396=>"100110000",
  55397=>"101011111",
  55398=>"101001111",
  55399=>"000111110",
  55400=>"010101001",
  55401=>"100111100",
  55402=>"101101111",
  55403=>"010111001",
  55404=>"110110001",
  55405=>"010000010",
  55406=>"110011001",
  55407=>"000101101",
  55408=>"001000001",
  55409=>"110100111",
  55410=>"100001001",
  55411=>"100101101",
  55412=>"010100010",
  55413=>"010010101",
  55414=>"010010001",
  55415=>"100111011",
  55416=>"111001110",
  55417=>"011010000",
  55418=>"011011010",
  55419=>"101111100",
  55420=>"011100001",
  55421=>"101111010",
  55422=>"010100000",
  55423=>"010010000",
  55424=>"111001001",
  55425=>"010100001",
  55426=>"010110011",
  55427=>"011100011",
  55428=>"001011000",
  55429=>"110101011",
  55430=>"110001010",
  55431=>"100011010",
  55432=>"101110010",
  55433=>"111101001",
  55434=>"101010101",
  55435=>"110110000",
  55436=>"001101101",
  55437=>"000000110",
  55438=>"101010111",
  55439=>"101000001",
  55440=>"110000101",
  55441=>"000111001",
  55442=>"110011010",
  55443=>"111011101",
  55444=>"100111000",
  55445=>"010100010",
  55446=>"010000011",
  55447=>"101101100",
  55448=>"000101100",
  55449=>"111111101",
  55450=>"100101010",
  55451=>"110110011",
  55452=>"000010000",
  55453=>"100111101",
  55454=>"100101101",
  55455=>"000001111",
  55456=>"100110111",
  55457=>"011110010",
  55458=>"100110001",
  55459=>"111101000",
  55460=>"110100100",
  55461=>"101000110",
  55462=>"000101110",
  55463=>"000100111",
  55464=>"011011110",
  55465=>"100000000",
  55466=>"111110011",
  55467=>"000111110",
  55468=>"101100101",
  55469=>"011001101",
  55470=>"001100001",
  55471=>"100011101",
  55472=>"011000010",
  55473=>"000110100",
  55474=>"000101010",
  55475=>"101100011",
  55476=>"000011101",
  55477=>"000111100",
  55478=>"101100101",
  55479=>"101011110",
  55480=>"100010101",
  55481=>"100011111",
  55482=>"001000000",
  55483=>"010111010",
  55484=>"111110110",
  55485=>"111000111",
  55486=>"001001001",
  55487=>"110001001",
  55488=>"000110011",
  55489=>"100111011",
  55490=>"100000110",
  55491=>"011000110",
  55492=>"111010110",
  55493=>"000011100",
  55494=>"100011010",
  55495=>"001001000",
  55496=>"100010110",
  55497=>"001010001",
  55498=>"000111001",
  55499=>"000101010",
  55500=>"110100100",
  55501=>"110111101",
  55502=>"011000101",
  55503=>"110010010",
  55504=>"011010110",
  55505=>"001011000",
  55506=>"010011011",
  55507=>"111100010",
  55508=>"000101110",
  55509=>"010000100",
  55510=>"011101001",
  55511=>"010001110",
  55512=>"001110001",
  55513=>"110111010",
  55514=>"000000111",
  55515=>"110001010",
  55516=>"000010000",
  55517=>"110001100",
  55518=>"001000000",
  55519=>"100011110",
  55520=>"111010000",
  55521=>"000110000",
  55522=>"100001110",
  55523=>"000000000",
  55524=>"100001110",
  55525=>"000001111",
  55526=>"100010001",
  55527=>"001001101",
  55528=>"000001101",
  55529=>"011100101",
  55530=>"001110100",
  55531=>"011101011",
  55532=>"100101101",
  55533=>"000100100",
  55534=>"110000011",
  55535=>"110101001",
  55536=>"110000000",
  55537=>"011011101",
  55538=>"001001000",
  55539=>"111111100",
  55540=>"010110000",
  55541=>"000001010",
  55542=>"011011101",
  55543=>"101000100",
  55544=>"110010110",
  55545=>"101101010",
  55546=>"010001111",
  55547=>"101100100",
  55548=>"001011110",
  55549=>"011010100",
  55550=>"000000011",
  55551=>"010100001",
  55552=>"100111101",
  55553=>"101111011",
  55554=>"111000111",
  55555=>"011110110",
  55556=>"110100111",
  55557=>"011000111",
  55558=>"010110101",
  55559=>"011000010",
  55560=>"111010111",
  55561=>"011010110",
  55562=>"110111110",
  55563=>"100111101",
  55564=>"000101111",
  55565=>"001110110",
  55566=>"001011110",
  55567=>"000111110",
  55568=>"101101011",
  55569=>"101101110",
  55570=>"010111001",
  55571=>"000001011",
  55572=>"100110011",
  55573=>"101010000",
  55574=>"001101111",
  55575=>"010111011",
  55576=>"010001010",
  55577=>"101101011",
  55578=>"111100110",
  55579=>"111100011",
  55580=>"111101101",
  55581=>"001001001",
  55582=>"001010011",
  55583=>"101110110",
  55584=>"001100100",
  55585=>"111000110",
  55586=>"001011111",
  55587=>"000100000",
  55588=>"001111011",
  55589=>"011011011",
  55590=>"011001100",
  55591=>"000111000",
  55592=>"100111100",
  55593=>"000101000",
  55594=>"111100011",
  55595=>"110011010",
  55596=>"101000111",
  55597=>"000110111",
  55598=>"110000101",
  55599=>"000101111",
  55600=>"101011111",
  55601=>"111001000",
  55602=>"100011111",
  55603=>"000001011",
  55604=>"010100101",
  55605=>"111000101",
  55606=>"001011010",
  55607=>"110111010",
  55608=>"100101110",
  55609=>"111111000",
  55610=>"100000100",
  55611=>"111110100",
  55612=>"101111100",
  55613=>"000101111",
  55614=>"110101111",
  55615=>"111010011",
  55616=>"101110101",
  55617=>"110100001",
  55618=>"101001100",
  55619=>"011101100",
  55620=>"110010111",
  55621=>"001000100",
  55622=>"000000100",
  55623=>"111000010",
  55624=>"101100111",
  55625=>"101100010",
  55626=>"110001000",
  55627=>"101011010",
  55628=>"011111110",
  55629=>"011000000",
  55630=>"001110100",
  55631=>"001100100",
  55632=>"111111100",
  55633=>"011001011",
  55634=>"000110111",
  55635=>"101111011",
  55636=>"101000111",
  55637=>"100101101",
  55638=>"011101101",
  55639=>"011010011",
  55640=>"101001110",
  55641=>"100011100",
  55642=>"110110011",
  55643=>"000100000",
  55644=>"000011000",
  55645=>"100011000",
  55646=>"010010011",
  55647=>"100000010",
  55648=>"001111011",
  55649=>"100011011",
  55650=>"000110101",
  55651=>"010101011",
  55652=>"000101101",
  55653=>"000101101",
  55654=>"001101011",
  55655=>"100001011",
  55656=>"010100101",
  55657=>"000100111",
  55658=>"010000101",
  55659=>"011001101",
  55660=>"110100100",
  55661=>"011101001",
  55662=>"000000100",
  55663=>"010010000",
  55664=>"000001010",
  55665=>"011101010",
  55666=>"010111101",
  55667=>"111110110",
  55668=>"100000110",
  55669=>"000001111",
  55670=>"101000010",
  55671=>"011110110",
  55672=>"110000111",
  55673=>"100010010",
  55674=>"110100111",
  55675=>"101101000",
  55676=>"011111101",
  55677=>"000110110",
  55678=>"100101101",
  55679=>"001100000",
  55680=>"010000111",
  55681=>"100001111",
  55682=>"001001110",
  55683=>"100010011",
  55684=>"000000111",
  55685=>"000000010",
  55686=>"000000100",
  55687=>"100100111",
  55688=>"011101100",
  55689=>"011111110",
  55690=>"110110100",
  55691=>"011000111",
  55692=>"110101110",
  55693=>"001111110",
  55694=>"111001011",
  55695=>"011101001",
  55696=>"110110100",
  55697=>"000010101",
  55698=>"010011111",
  55699=>"010010001",
  55700=>"100000010",
  55701=>"000100100",
  55702=>"100110111",
  55703=>"000100001",
  55704=>"000001110",
  55705=>"010010001",
  55706=>"001100001",
  55707=>"000000000",
  55708=>"000000001",
  55709=>"011010110",
  55710=>"001011010",
  55711=>"001011000",
  55712=>"101100010",
  55713=>"111111001",
  55714=>"000001000",
  55715=>"011011001",
  55716=>"100110111",
  55717=>"101001110",
  55718=>"010000100",
  55719=>"101001001",
  55720=>"010111110",
  55721=>"101100111",
  55722=>"000001101",
  55723=>"101101100",
  55724=>"011000001",
  55725=>"111110111",
  55726=>"000000011",
  55727=>"111101110",
  55728=>"001111000",
  55729=>"011100011",
  55730=>"011100101",
  55731=>"111111110",
  55732=>"110110110",
  55733=>"011100100",
  55734=>"011101001",
  55735=>"110111010",
  55736=>"000100100",
  55737=>"000100011",
  55738=>"000010110",
  55739=>"100011100",
  55740=>"101101000",
  55741=>"011011001",
  55742=>"000111110",
  55743=>"101000101",
  55744=>"100101111",
  55745=>"101110011",
  55746=>"011100101",
  55747=>"101100101",
  55748=>"000110111",
  55749=>"011101111",
  55750=>"000001010",
  55751=>"111011110",
  55752=>"111111110",
  55753=>"001000110",
  55754=>"000011100",
  55755=>"000101101",
  55756=>"010101010",
  55757=>"000100110",
  55758=>"000000100",
  55759=>"111000010",
  55760=>"111101100",
  55761=>"011000111",
  55762=>"110011100",
  55763=>"101011111",
  55764=>"010111110",
  55765=>"110111000",
  55766=>"111001000",
  55767=>"100110101",
  55768=>"110100010",
  55769=>"110000111",
  55770=>"100011110",
  55771=>"101100000",
  55772=>"101001100",
  55773=>"000110001",
  55774=>"101110110",
  55775=>"111001010",
  55776=>"110011011",
  55777=>"010000100",
  55778=>"101110101",
  55779=>"100100000",
  55780=>"001001110",
  55781=>"101101111",
  55782=>"001110010",
  55783=>"010101100",
  55784=>"001111010",
  55785=>"010110100",
  55786=>"111001001",
  55787=>"010101100",
  55788=>"110111110",
  55789=>"001000001",
  55790=>"100001010",
  55791=>"110001110",
  55792=>"001000010",
  55793=>"110111101",
  55794=>"101010001",
  55795=>"000100011",
  55796=>"000010011",
  55797=>"001100100",
  55798=>"110010101",
  55799=>"101011001",
  55800=>"110010010",
  55801=>"001101110",
  55802=>"011010000",
  55803=>"110101010",
  55804=>"011100010",
  55805=>"101011100",
  55806=>"001000011",
  55807=>"001111000",
  55808=>"100011010",
  55809=>"111001001",
  55810=>"111011000",
  55811=>"111100110",
  55812=>"010110110",
  55813=>"000100101",
  55814=>"000110111",
  55815=>"000011010",
  55816=>"000000001",
  55817=>"110101011",
  55818=>"100001010",
  55819=>"010000011",
  55820=>"000010000",
  55821=>"010110101",
  55822=>"111000111",
  55823=>"001011011",
  55824=>"000110101",
  55825=>"001111010",
  55826=>"110100001",
  55827=>"001101001",
  55828=>"011110110",
  55829=>"001101111",
  55830=>"011010111",
  55831=>"111010110",
  55832=>"010000010",
  55833=>"110101101",
  55834=>"110100100",
  55835=>"101001001",
  55836=>"101100010",
  55837=>"100000110",
  55838=>"101101100",
  55839=>"011001100",
  55840=>"101100110",
  55841=>"101001111",
  55842=>"000001010",
  55843=>"010001101",
  55844=>"111011111",
  55845=>"101110001",
  55846=>"011011110",
  55847=>"010010111",
  55848=>"111111001",
  55849=>"000011010",
  55850=>"000101011",
  55851=>"100100011",
  55852=>"100111100",
  55853=>"000001010",
  55854=>"000111000",
  55855=>"000000001",
  55856=>"110111010",
  55857=>"111000111",
  55858=>"100111100",
  55859=>"100110110",
  55860=>"110010110",
  55861=>"100110100",
  55862=>"000011010",
  55863=>"110011010",
  55864=>"010001001",
  55865=>"010001011",
  55866=>"000111111",
  55867=>"110001111",
  55868=>"001011011",
  55869=>"010000010",
  55870=>"011111000",
  55871=>"011110010",
  55872=>"101111110",
  55873=>"000000001",
  55874=>"001001110",
  55875=>"100011001",
  55876=>"011011000",
  55877=>"011011010",
  55878=>"101000011",
  55879=>"000101010",
  55880=>"111111111",
  55881=>"101100101",
  55882=>"111101100",
  55883=>"010101111",
  55884=>"010001000",
  55885=>"010000101",
  55886=>"110101000",
  55887=>"101101010",
  55888=>"010101001",
  55889=>"111110111",
  55890=>"110100101",
  55891=>"010001111",
  55892=>"110000111",
  55893=>"100101101",
  55894=>"100111101",
  55895=>"110100100",
  55896=>"110010101",
  55897=>"001011000",
  55898=>"001111001",
  55899=>"001010100",
  55900=>"011001001",
  55901=>"110010101",
  55902=>"010001010",
  55903=>"111111101",
  55904=>"010001010",
  55905=>"111010101",
  55906=>"001100000",
  55907=>"011001010",
  55908=>"101011001",
  55909=>"011000110",
  55910=>"010110100",
  55911=>"101001111",
  55912=>"110100001",
  55913=>"010010110",
  55914=>"010111101",
  55915=>"000000110",
  55916=>"000100010",
  55917=>"011010001",
  55918=>"101000101",
  55919=>"101001111",
  55920=>"100101000",
  55921=>"110100110",
  55922=>"111111010",
  55923=>"011001110",
  55924=>"111000011",
  55925=>"001000011",
  55926=>"101100101",
  55927=>"110101110",
  55928=>"111010100",
  55929=>"110110111",
  55930=>"000100000",
  55931=>"011000000",
  55932=>"001000100",
  55933=>"010101010",
  55934=>"000100100",
  55935=>"001110100",
  55936=>"010000110",
  55937=>"100000111",
  55938=>"110001010",
  55939=>"010010100",
  55940=>"100000000",
  55941=>"110000000",
  55942=>"100111001",
  55943=>"011010010",
  55944=>"000111000",
  55945=>"001001111",
  55946=>"011101101",
  55947=>"110100100",
  55948=>"110111001",
  55949=>"001100101",
  55950=>"110001100",
  55951=>"000010110",
  55952=>"011101011",
  55953=>"010111010",
  55954=>"111011101",
  55955=>"111010110",
  55956=>"001000000",
  55957=>"001101001",
  55958=>"001000100",
  55959=>"010100001",
  55960=>"110111101",
  55961=>"010110001",
  55962=>"011101111",
  55963=>"000011001",
  55964=>"110001011",
  55965=>"101010011",
  55966=>"111111010",
  55967=>"101111110",
  55968=>"111000010",
  55969=>"111110011",
  55970=>"010110010",
  55971=>"111101111",
  55972=>"111101110",
  55973=>"000100011",
  55974=>"000111100",
  55975=>"010000100",
  55976=>"010101000",
  55977=>"111010110",
  55978=>"000100111",
  55979=>"101001101",
  55980=>"000110111",
  55981=>"000001110",
  55982=>"100111101",
  55983=>"001110011",
  55984=>"010011111",
  55985=>"001001011",
  55986=>"101101001",
  55987=>"111010100",
  55988=>"000010011",
  55989=>"010110100",
  55990=>"111101101",
  55991=>"010000010",
  55992=>"011001110",
  55993=>"010010000",
  55994=>"011011001",
  55995=>"101111101",
  55996=>"011010011",
  55997=>"001100110",
  55998=>"100111010",
  55999=>"101100111",
  56000=>"110001010",
  56001=>"100001000",
  56002=>"000100001",
  56003=>"111011011",
  56004=>"011101010",
  56005=>"111000011",
  56006=>"001110000",
  56007=>"101100011",
  56008=>"010001110",
  56009=>"101001000",
  56010=>"010111001",
  56011=>"111011100",
  56012=>"000111010",
  56013=>"010100001",
  56014=>"110100110",
  56015=>"000100110",
  56016=>"001000111",
  56017=>"011000001",
  56018=>"011000110",
  56019=>"000110110",
  56020=>"100100011",
  56021=>"000000110",
  56022=>"001100111",
  56023=>"101000111",
  56024=>"101100010",
  56025=>"011111000",
  56026=>"110111000",
  56027=>"011001000",
  56028=>"110110101",
  56029=>"010110001",
  56030=>"011000110",
  56031=>"100010111",
  56032=>"110100101",
  56033=>"100000000",
  56034=>"100101111",
  56035=>"100101111",
  56036=>"000000011",
  56037=>"100011011",
  56038=>"101011110",
  56039=>"100100110",
  56040=>"000010110",
  56041=>"101100100",
  56042=>"111110001",
  56043=>"101110110",
  56044=>"111010110",
  56045=>"001010111",
  56046=>"110000111",
  56047=>"000010010",
  56048=>"001010010",
  56049=>"001111101",
  56050=>"010100001",
  56051=>"000111101",
  56052=>"001100000",
  56053=>"100100000",
  56054=>"111010110",
  56055=>"110110101",
  56056=>"110110000",
  56057=>"111100001",
  56058=>"100110100",
  56059=>"000010000",
  56060=>"111100010",
  56061=>"100010101",
  56062=>"000010101",
  56063=>"100110010",
  56064=>"100000000",
  56065=>"101001011",
  56066=>"011000110",
  56067=>"101000000",
  56068=>"001001000",
  56069=>"011100111",
  56070=>"101010100",
  56071=>"001011100",
  56072=>"000101100",
  56073=>"110111011",
  56074=>"000111111",
  56075=>"111100100",
  56076=>"111110100",
  56077=>"011100000",
  56078=>"010101100",
  56079=>"100000001",
  56080=>"010011000",
  56081=>"111010011",
  56082=>"110001011",
  56083=>"111001010",
  56084=>"001001111",
  56085=>"000011010",
  56086=>"001111000",
  56087=>"000000111",
  56088=>"100111000",
  56089=>"111110110",
  56090=>"000000001",
  56091=>"100011001",
  56092=>"010001101",
  56093=>"110010000",
  56094=>"111011101",
  56095=>"111110101",
  56096=>"101010100",
  56097=>"111111000",
  56098=>"111110101",
  56099=>"011100111",
  56100=>"010110011",
  56101=>"101011001",
  56102=>"100001001",
  56103=>"001000011",
  56104=>"001000101",
  56105=>"010011000",
  56106=>"001111010",
  56107=>"110101001",
  56108=>"000010001",
  56109=>"011001100",
  56110=>"111111001",
  56111=>"101111111",
  56112=>"101000001",
  56113=>"000010010",
  56114=>"110111000",
  56115=>"010010010",
  56116=>"101001111",
  56117=>"100110000",
  56118=>"110000011",
  56119=>"011101010",
  56120=>"001100001",
  56121=>"110100111",
  56122=>"100010001",
  56123=>"110001100",
  56124=>"111110101",
  56125=>"111001010",
  56126=>"111101000",
  56127=>"010111101",
  56128=>"111011111",
  56129=>"101110001",
  56130=>"001010101",
  56131=>"110101111",
  56132=>"000010101",
  56133=>"111110010",
  56134=>"111101101",
  56135=>"111101011",
  56136=>"111010000",
  56137=>"110001101",
  56138=>"001001101",
  56139=>"100010011",
  56140=>"000110111",
  56141=>"111101010",
  56142=>"111101111",
  56143=>"111101001",
  56144=>"100010000",
  56145=>"111111011",
  56146=>"100101000",
  56147=>"110100110",
  56148=>"101110011",
  56149=>"100011001",
  56150=>"000011011",
  56151=>"100100011",
  56152=>"011010001",
  56153=>"101111110",
  56154=>"100010111",
  56155=>"111011001",
  56156=>"011010001",
  56157=>"001111101",
  56158=>"010000110",
  56159=>"011000010",
  56160=>"001010010",
  56161=>"010101000",
  56162=>"001111111",
  56163=>"010000000",
  56164=>"000110000",
  56165=>"011001000",
  56166=>"110110100",
  56167=>"001010010",
  56168=>"111001001",
  56169=>"110111001",
  56170=>"001010010",
  56171=>"101011100",
  56172=>"111000000",
  56173=>"001100101",
  56174=>"000001001",
  56175=>"001010111",
  56176=>"100010010",
  56177=>"011111110",
  56178=>"000100110",
  56179=>"010001010",
  56180=>"101100101",
  56181=>"001011111",
  56182=>"000011011",
  56183=>"110010100",
  56184=>"011010110",
  56185=>"111010100",
  56186=>"111011010",
  56187=>"101010110",
  56188=>"010001111",
  56189=>"011000011",
  56190=>"110001110",
  56191=>"001010111",
  56192=>"000001110",
  56193=>"111110011",
  56194=>"011000111",
  56195=>"010111010",
  56196=>"011011000",
  56197=>"010010000",
  56198=>"000101110",
  56199=>"111011001",
  56200=>"101111001",
  56201=>"001110101",
  56202=>"001110000",
  56203=>"000011010",
  56204=>"111101010",
  56205=>"111101000",
  56206=>"101011101",
  56207=>"111001111",
  56208=>"101110001",
  56209=>"000101010",
  56210=>"101000101",
  56211=>"111101000",
  56212=>"101011110",
  56213=>"101011111",
  56214=>"011101000",
  56215=>"110001000",
  56216=>"101000100",
  56217=>"111100101",
  56218=>"001000111",
  56219=>"010010111",
  56220=>"110101100",
  56221=>"110001010",
  56222=>"101001011",
  56223=>"001111001",
  56224=>"110011000",
  56225=>"011000010",
  56226=>"000101101",
  56227=>"001001000",
  56228=>"011010100",
  56229=>"100010111",
  56230=>"100110111",
  56231=>"011010110",
  56232=>"110001111",
  56233=>"100110111",
  56234=>"000110110",
  56235=>"110001111",
  56236=>"010110100",
  56237=>"001011101",
  56238=>"111010010",
  56239=>"000011101",
  56240=>"000011110",
  56241=>"010010101",
  56242=>"011110111",
  56243=>"100000100",
  56244=>"000111110",
  56245=>"010010010",
  56246=>"000001110",
  56247=>"111110000",
  56248=>"101011011",
  56249=>"010101110",
  56250=>"101000000",
  56251=>"100101100",
  56252=>"010101010",
  56253=>"011011001",
  56254=>"101010111",
  56255=>"111111110",
  56256=>"100101111",
  56257=>"011101001",
  56258=>"101010111",
  56259=>"111000001",
  56260=>"001110001",
  56261=>"011010111",
  56262=>"100101000",
  56263=>"101111001",
  56264=>"000000001",
  56265=>"000001010",
  56266=>"001100110",
  56267=>"100000000",
  56268=>"111011111",
  56269=>"000111110",
  56270=>"000000100",
  56271=>"011000110",
  56272=>"001010111",
  56273=>"100111111",
  56274=>"011111110",
  56275=>"111110100",
  56276=>"000000001",
  56277=>"001111100",
  56278=>"010001001",
  56279=>"000111100",
  56280=>"011010100",
  56281=>"011111000",
  56282=>"010011010",
  56283=>"000000001",
  56284=>"001110110",
  56285=>"001000010",
  56286=>"011111000",
  56287=>"000011011",
  56288=>"101010101",
  56289=>"000011011",
  56290=>"100011111",
  56291=>"100011010",
  56292=>"110110100",
  56293=>"000000000",
  56294=>"100010011",
  56295=>"111101000",
  56296=>"001110111",
  56297=>"011011001",
  56298=>"010000000",
  56299=>"100010011",
  56300=>"111011010",
  56301=>"100001110",
  56302=>"100011001",
  56303=>"100011000",
  56304=>"100001110",
  56305=>"010110110",
  56306=>"000000000",
  56307=>"010101101",
  56308=>"001110101",
  56309=>"111101001",
  56310=>"000101110",
  56311=>"101001111",
  56312=>"011011100",
  56313=>"011001111",
  56314=>"111100101",
  56315=>"100011100",
  56316=>"011100011",
  56317=>"100101001",
  56318=>"110011000",
  56319=>"011101111",
  56320=>"111100110",
  56321=>"000000101",
  56322=>"101111010",
  56323=>"101101001",
  56324=>"011000010",
  56325=>"110111001",
  56326=>"101000111",
  56327=>"101101111",
  56328=>"111011101",
  56329=>"000001001",
  56330=>"111101110",
  56331=>"110100010",
  56332=>"101000010",
  56333=>"001000110",
  56334=>"100101110",
  56335=>"011001010",
  56336=>"010111011",
  56337=>"110001001",
  56338=>"011100000",
  56339=>"010111100",
  56340=>"111111110",
  56341=>"000010100",
  56342=>"111010100",
  56343=>"000010111",
  56344=>"000001000",
  56345=>"111110010",
  56346=>"101111000",
  56347=>"011000110",
  56348=>"110000011",
  56349=>"101100101",
  56350=>"010100111",
  56351=>"111100010",
  56352=>"100011011",
  56353=>"010011101",
  56354=>"100011000",
  56355=>"010101010",
  56356=>"110101111",
  56357=>"000000100",
  56358=>"010001010",
  56359=>"111110101",
  56360=>"110010010",
  56361=>"001001001",
  56362=>"011001100",
  56363=>"000110111",
  56364=>"001110110",
  56365=>"001100101",
  56366=>"111011111",
  56367=>"101111001",
  56368=>"111111010",
  56369=>"000100110",
  56370=>"011010101",
  56371=>"101010000",
  56372=>"111110011",
  56373=>"001010011",
  56374=>"010101110",
  56375=>"010111010",
  56376=>"100000001",
  56377=>"011010011",
  56378=>"100010110",
  56379=>"110010001",
  56380=>"000001010",
  56381=>"010011111",
  56382=>"011100100",
  56383=>"100010101",
  56384=>"100010001",
  56385=>"011000111",
  56386=>"001000011",
  56387=>"001000000",
  56388=>"000010100",
  56389=>"101100101",
  56390=>"111100000",
  56391=>"000111011",
  56392=>"011100100",
  56393=>"111111011",
  56394=>"001000111",
  56395=>"001001000",
  56396=>"010100101",
  56397=>"111011101",
  56398=>"001110101",
  56399=>"101111001",
  56400=>"011000010",
  56401=>"000011111",
  56402=>"110101101",
  56403=>"000001100",
  56404=>"001000110",
  56405=>"101100100",
  56406=>"110001101",
  56407=>"000101110",
  56408=>"111110011",
  56409=>"101111001",
  56410=>"100110101",
  56411=>"101110100",
  56412=>"111101001",
  56413=>"101101111",
  56414=>"111011101",
  56415=>"100111000",
  56416=>"110000100",
  56417=>"010100001",
  56418=>"000100100",
  56419=>"110100100",
  56420=>"001100110",
  56421=>"001100100",
  56422=>"100101010",
  56423=>"111000111",
  56424=>"010111010",
  56425=>"100101001",
  56426=>"011000001",
  56427=>"001111000",
  56428=>"100101000",
  56429=>"001100110",
  56430=>"101000010",
  56431=>"011100100",
  56432=>"100111100",
  56433=>"011000010",
  56434=>"010100000",
  56435=>"001111010",
  56436=>"100110100",
  56437=>"010110000",
  56438=>"110000010",
  56439=>"011000000",
  56440=>"100001100",
  56441=>"101110001",
  56442=>"111011010",
  56443=>"001001110",
  56444=>"000101000",
  56445=>"011100101",
  56446=>"111111000",
  56447=>"001110001",
  56448=>"101000111",
  56449=>"111011110",
  56450=>"101001010",
  56451=>"111011010",
  56452=>"001100110",
  56453=>"001101010",
  56454=>"110000011",
  56455=>"110101101",
  56456=>"110101110",
  56457=>"101011100",
  56458=>"100000110",
  56459=>"110010111",
  56460=>"000100100",
  56461=>"110001011",
  56462=>"001110111",
  56463=>"011000110",
  56464=>"011101100",
  56465=>"001010101",
  56466=>"101000010",
  56467=>"110011011",
  56468=>"110101100",
  56469=>"101001010",
  56470=>"001110111",
  56471=>"111010010",
  56472=>"000111110",
  56473=>"110100000",
  56474=>"100010101",
  56475=>"110111011",
  56476=>"010001000",
  56477=>"101111100",
  56478=>"011110010",
  56479=>"011110001",
  56480=>"011011111",
  56481=>"101110101",
  56482=>"100110010",
  56483=>"110110000",
  56484=>"111110111",
  56485=>"001010110",
  56486=>"011001100",
  56487=>"110000011",
  56488=>"110000010",
  56489=>"101010001",
  56490=>"111110000",
  56491=>"010000010",
  56492=>"101110101",
  56493=>"000101111",
  56494=>"000101110",
  56495=>"110010010",
  56496=>"010001011",
  56497=>"010001000",
  56498=>"001101100",
  56499=>"111101011",
  56500=>"001110000",
  56501=>"000110000",
  56502=>"111010101",
  56503=>"010011111",
  56504=>"001110110",
  56505=>"000000001",
  56506=>"111000100",
  56507=>"001011000",
  56508=>"010111011",
  56509=>"000010101",
  56510=>"110100101",
  56511=>"001011101",
  56512=>"010110011",
  56513=>"101000110",
  56514=>"101100110",
  56515=>"001010101",
  56516=>"111100010",
  56517=>"000010000",
  56518=>"000111010",
  56519=>"001100011",
  56520=>"001111110",
  56521=>"100010000",
  56522=>"011100111",
  56523=>"110110101",
  56524=>"011011111",
  56525=>"101001111",
  56526=>"000110000",
  56527=>"001001000",
  56528=>"011100110",
  56529=>"010000010",
  56530=>"101001010",
  56531=>"101100100",
  56532=>"111001001",
  56533=>"111101111",
  56534=>"101101001",
  56535=>"000111110",
  56536=>"010011110",
  56537=>"000010000",
  56538=>"111100101",
  56539=>"100000111",
  56540=>"010000010",
  56541=>"011111110",
  56542=>"111101110",
  56543=>"001011100",
  56544=>"101001100",
  56545=>"111111010",
  56546=>"101111100",
  56547=>"101111010",
  56548=>"010101000",
  56549=>"100100110",
  56550=>"110011100",
  56551=>"010111100",
  56552=>"110100000",
  56553=>"000010011",
  56554=>"000010011",
  56555=>"000011011",
  56556=>"101011001",
  56557=>"110111001",
  56558=>"010011011",
  56559=>"010101111",
  56560=>"101000011",
  56561=>"101000101",
  56562=>"111011100",
  56563=>"011100100",
  56564=>"000000000",
  56565=>"011000100",
  56566=>"011110011",
  56567=>"001110111",
  56568=>"011101100",
  56569=>"100100001",
  56570=>"111000111",
  56571=>"011100110",
  56572=>"011011100",
  56573=>"111100110",
  56574=>"101110111",
  56575=>"101001011",
  56576=>"010111000",
  56577=>"011010111",
  56578=>"101000011",
  56579=>"010111100",
  56580=>"100100111",
  56581=>"000000001",
  56582=>"111110000",
  56583=>"110100000",
  56584=>"011110101",
  56585=>"011101100",
  56586=>"000011011",
  56587=>"010000001",
  56588=>"100011000",
  56589=>"110110011",
  56590=>"100000011",
  56591=>"110100001",
  56592=>"010000000",
  56593=>"110010101",
  56594=>"111101101",
  56595=>"010101010",
  56596=>"110101110",
  56597=>"011110000",
  56598=>"111111011",
  56599=>"000010101",
  56600=>"000100110",
  56601=>"011111001",
  56602=>"011111011",
  56603=>"101010110",
  56604=>"110101011",
  56605=>"000000101",
  56606=>"111000001",
  56607=>"000001010",
  56608=>"100011011",
  56609=>"100011110",
  56610=>"111110101",
  56611=>"010101000",
  56612=>"111101001",
  56613=>"001000000",
  56614=>"111000011",
  56615=>"001001001",
  56616=>"100101011",
  56617=>"111100100",
  56618=>"001101111",
  56619=>"011000100",
  56620=>"001011011",
  56621=>"000000101",
  56622=>"011000101",
  56623=>"110010010",
  56624=>"011100101",
  56625=>"110000001",
  56626=>"100100101",
  56627=>"011010000",
  56628=>"101101110",
  56629=>"010011101",
  56630=>"001000110",
  56631=>"011111001",
  56632=>"001001100",
  56633=>"011001100",
  56634=>"111111000",
  56635=>"011000101",
  56636=>"111101101",
  56637=>"101101101",
  56638=>"110011001",
  56639=>"110010001",
  56640=>"110101001",
  56641=>"011100110",
  56642=>"110100000",
  56643=>"010101110",
  56644=>"010100111",
  56645=>"011110001",
  56646=>"000000101",
  56647=>"000100000",
  56648=>"010011000",
  56649=>"111010000",
  56650=>"111001100",
  56651=>"100111011",
  56652=>"000011011",
  56653=>"011111100",
  56654=>"001001000",
  56655=>"010010000",
  56656=>"001111100",
  56657=>"111001110",
  56658=>"001100011",
  56659=>"011000011",
  56660=>"010100001",
  56661=>"010000001",
  56662=>"001000110",
  56663=>"010011001",
  56664=>"011111001",
  56665=>"001010111",
  56666=>"010010110",
  56667=>"001000110",
  56668=>"111111100",
  56669=>"110011000",
  56670=>"001101000",
  56671=>"111000010",
  56672=>"000110110",
  56673=>"001011000",
  56674=>"010100000",
  56675=>"001000011",
  56676=>"011001100",
  56677=>"011101010",
  56678=>"001111000",
  56679=>"010110001",
  56680=>"001111100",
  56681=>"001110011",
  56682=>"111111101",
  56683=>"001001110",
  56684=>"101110101",
  56685=>"111110101",
  56686=>"100000010",
  56687=>"000101110",
  56688=>"000101011",
  56689=>"110111110",
  56690=>"111000010",
  56691=>"110010101",
  56692=>"101100111",
  56693=>"111111011",
  56694=>"011100100",
  56695=>"111011001",
  56696=>"111000010",
  56697=>"111001010",
  56698=>"100111101",
  56699=>"000011101",
  56700=>"001010100",
  56701=>"100110000",
  56702=>"110110101",
  56703=>"110110111",
  56704=>"111101101",
  56705=>"001000011",
  56706=>"101111100",
  56707=>"100000000",
  56708=>"011100000",
  56709=>"011010001",
  56710=>"001110111",
  56711=>"110000110",
  56712=>"100010101",
  56713=>"000100100",
  56714=>"111011000",
  56715=>"000010100",
  56716=>"010111110",
  56717=>"000100111",
  56718=>"001101111",
  56719=>"011011101",
  56720=>"101110101",
  56721=>"000011010",
  56722=>"110101000",
  56723=>"001000001",
  56724=>"100010011",
  56725=>"001100100",
  56726=>"111101000",
  56727=>"011001000",
  56728=>"011010100",
  56729=>"001011001",
  56730=>"101011010",
  56731=>"111000011",
  56732=>"000010110",
  56733=>"011010001",
  56734=>"111011111",
  56735=>"110101010",
  56736=>"110100010",
  56737=>"000000100",
  56738=>"000010110",
  56739=>"010000000",
  56740=>"111110001",
  56741=>"001000000",
  56742=>"111111000",
  56743=>"010101101",
  56744=>"011111110",
  56745=>"101111111",
  56746=>"000000110",
  56747=>"100011011",
  56748=>"011110111",
  56749=>"101011110",
  56750=>"000010000",
  56751=>"001010101",
  56752=>"110100010",
  56753=>"000001000",
  56754=>"011100101",
  56755=>"111111100",
  56756=>"001011010",
  56757=>"110010000",
  56758=>"011111110",
  56759=>"001000001",
  56760=>"100101010",
  56761=>"111000110",
  56762=>"001011101",
  56763=>"001011101",
  56764=>"010000000",
  56765=>"011101000",
  56766=>"000110010",
  56767=>"101110001",
  56768=>"001011111",
  56769=>"110111000",
  56770=>"100000100",
  56771=>"000000100",
  56772=>"001100110",
  56773=>"000100101",
  56774=>"001000100",
  56775=>"111010010",
  56776=>"111101101",
  56777=>"000100010",
  56778=>"011100110",
  56779=>"110001110",
  56780=>"100100111",
  56781=>"001011010",
  56782=>"000111001",
  56783=>"000001110",
  56784=>"010010001",
  56785=>"010111111",
  56786=>"011001111",
  56787=>"101111110",
  56788=>"011101011",
  56789=>"101011111",
  56790=>"100110111",
  56791=>"011111001",
  56792=>"010010111",
  56793=>"010101101",
  56794=>"010101011",
  56795=>"100111100",
  56796=>"100101100",
  56797=>"100100001",
  56798=>"000101011",
  56799=>"000100111",
  56800=>"011111000",
  56801=>"100101011",
  56802=>"100111001",
  56803=>"001010010",
  56804=>"110111010",
  56805=>"011010100",
  56806=>"000001000",
  56807=>"101100000",
  56808=>"001111110",
  56809=>"001110110",
  56810=>"010111100",
  56811=>"000001110",
  56812=>"010110010",
  56813=>"010111010",
  56814=>"101100010",
  56815=>"111100110",
  56816=>"000111001",
  56817=>"000100111",
  56818=>"110111100",
  56819=>"101100111",
  56820=>"000000100",
  56821=>"000000101",
  56822=>"100100101",
  56823=>"100111011",
  56824=>"100101111",
  56825=>"111111110",
  56826=>"100000110",
  56827=>"000001010",
  56828=>"001000000",
  56829=>"101110000",
  56830=>"011100000",
  56831=>"000010000",
  56832=>"011100001",
  56833=>"000001010",
  56834=>"000101110",
  56835=>"110000001",
  56836=>"011010000",
  56837=>"000000001",
  56838=>"110010011",
  56839=>"000101111",
  56840=>"000001110",
  56841=>"010111110",
  56842=>"101001101",
  56843=>"010111000",
  56844=>"001001101",
  56845=>"010001111",
  56846=>"000001011",
  56847=>"100100110",
  56848=>"111001001",
  56849=>"011001000",
  56850=>"001101000",
  56851=>"000000111",
  56852=>"001001100",
  56853=>"100001000",
  56854=>"100010010",
  56855=>"111001001",
  56856=>"100010001",
  56857=>"001000100",
  56858=>"000001000",
  56859=>"110110110",
  56860=>"001101110",
  56861=>"011010111",
  56862=>"110101100",
  56863=>"010110111",
  56864=>"000100000",
  56865=>"101010000",
  56866=>"100000000",
  56867=>"111100001",
  56868=>"001001100",
  56869=>"111011110",
  56870=>"010100110",
  56871=>"010101001",
  56872=>"000101011",
  56873=>"010011110",
  56874=>"111011100",
  56875=>"111101110",
  56876=>"101000010",
  56877=>"101101100",
  56878=>"010111011",
  56879=>"111001001",
  56880=>"110101111",
  56881=>"100110001",
  56882=>"101000000",
  56883=>"101101001",
  56884=>"001111001",
  56885=>"011110010",
  56886=>"101101101",
  56887=>"000100011",
  56888=>"010110101",
  56889=>"110001111",
  56890=>"001000001",
  56891=>"110101111",
  56892=>"010100000",
  56893=>"001010011",
  56894=>"001000000",
  56895=>"000010110",
  56896=>"101111111",
  56897=>"011110100",
  56898=>"011110011",
  56899=>"000001000",
  56900=>"011010100",
  56901=>"100101001",
  56902=>"101110000",
  56903=>"110000101",
  56904=>"010101000",
  56905=>"100010010",
  56906=>"010010110",
  56907=>"110100011",
  56908=>"010010000",
  56909=>"100100011",
  56910=>"011011111",
  56911=>"000000001",
  56912=>"110101101",
  56913=>"101101010",
  56914=>"100100010",
  56915=>"001000101",
  56916=>"111101100",
  56917=>"001011011",
  56918=>"010111000",
  56919=>"110011011",
  56920=>"111001111",
  56921=>"111111100",
  56922=>"111101010",
  56923=>"100101100",
  56924=>"010100010",
  56925=>"000000100",
  56926=>"000011010",
  56927=>"111111111",
  56928=>"010100001",
  56929=>"010001000",
  56930=>"111011000",
  56931=>"110111101",
  56932=>"111111111",
  56933=>"000011000",
  56934=>"001100111",
  56935=>"010001000",
  56936=>"000110100",
  56937=>"010101010",
  56938=>"100110101",
  56939=>"100100101",
  56940=>"010100110",
  56941=>"100001100",
  56942=>"110001000",
  56943=>"100101110",
  56944=>"110010001",
  56945=>"101011100",
  56946=>"010000110",
  56947=>"111111100",
  56948=>"011001110",
  56949=>"001000111",
  56950=>"101011100",
  56951=>"001110111",
  56952=>"101010000",
  56953=>"101110111",
  56954=>"001101011",
  56955=>"010011101",
  56956=>"101001000",
  56957=>"010011111",
  56958=>"110110110",
  56959=>"111111111",
  56960=>"000100110",
  56961=>"111010100",
  56962=>"110111100",
  56963=>"101111000",
  56964=>"100001011",
  56965=>"000100011",
  56966=>"011110011",
  56967=>"110011010",
  56968=>"101010111",
  56969=>"111111000",
  56970=>"111011111",
  56971=>"110110111",
  56972=>"010001110",
  56973=>"000000111",
  56974=>"000000001",
  56975=>"111100101",
  56976=>"101110011",
  56977=>"111110010",
  56978=>"001001111",
  56979=>"011110101",
  56980=>"011001100",
  56981=>"010111111",
  56982=>"011111110",
  56983=>"101111110",
  56984=>"011100100",
  56985=>"011011100",
  56986=>"101111100",
  56987=>"110100110",
  56988=>"110100101",
  56989=>"000110010",
  56990=>"000000101",
  56991=>"111000101",
  56992=>"111001010",
  56993=>"010011101",
  56994=>"101001111",
  56995=>"000110100",
  56996=>"010101001",
  56997=>"100100011",
  56998=>"110110100",
  56999=>"100000000",
  57000=>"011011101",
  57001=>"110110000",
  57002=>"101101011",
  57003=>"001001100",
  57004=>"111010100",
  57005=>"101110000",
  57006=>"010100110",
  57007=>"011100000",
  57008=>"100111001",
  57009=>"111000011",
  57010=>"011100000",
  57011=>"111111001",
  57012=>"010111010",
  57013=>"010001110",
  57014=>"000101111",
  57015=>"000000001",
  57016=>"001010001",
  57017=>"001001011",
  57018=>"101111011",
  57019=>"001001111",
  57020=>"111011101",
  57021=>"001001110",
  57022=>"000100111",
  57023=>"110011001",
  57024=>"101110010",
  57025=>"010110111",
  57026=>"110100101",
  57027=>"110101000",
  57028=>"111111011",
  57029=>"000011011",
  57030=>"000001101",
  57031=>"001100000",
  57032=>"001110101",
  57033=>"101010011",
  57034=>"000110010",
  57035=>"111000111",
  57036=>"010000111",
  57037=>"110001101",
  57038=>"000100000",
  57039=>"000000001",
  57040=>"100000110",
  57041=>"100010101",
  57042=>"111001111",
  57043=>"100010110",
  57044=>"101001101",
  57045=>"100011000",
  57046=>"111000100",
  57047=>"010011000",
  57048=>"101011000",
  57049=>"011000011",
  57050=>"111111001",
  57051=>"001001111",
  57052=>"000101001",
  57053=>"110001010",
  57054=>"010011011",
  57055=>"011111111",
  57056=>"000010000",
  57057=>"000100010",
  57058=>"110111011",
  57059=>"010101001",
  57060=>"100110101",
  57061=>"011100111",
  57062=>"101101011",
  57063=>"101010101",
  57064=>"001010100",
  57065=>"110100011",
  57066=>"111011101",
  57067=>"111110011",
  57068=>"011001010",
  57069=>"000100110",
  57070=>"001101110",
  57071=>"000001001",
  57072=>"110011110",
  57073=>"001011110",
  57074=>"110011010",
  57075=>"110010101",
  57076=>"101100011",
  57077=>"111100111",
  57078=>"011101011",
  57079=>"001001110",
  57080=>"111100011",
  57081=>"000011101",
  57082=>"000001111",
  57083=>"111100000",
  57084=>"000000000",
  57085=>"000111010",
  57086=>"101111110",
  57087=>"110000011",
  57088=>"110100000",
  57089=>"001000010",
  57090=>"101101100",
  57091=>"111011000",
  57092=>"110010000",
  57093=>"101001010",
  57094=>"111100111",
  57095=>"010011111",
  57096=>"001100000",
  57097=>"000100001",
  57098=>"110100111",
  57099=>"000000001",
  57100=>"111110011",
  57101=>"111011101",
  57102=>"110010001",
  57103=>"101110010",
  57104=>"111111010",
  57105=>"010101011",
  57106=>"001001111",
  57107=>"111011110",
  57108=>"010101110",
  57109=>"001011010",
  57110=>"011111111",
  57111=>"001111001",
  57112=>"001110101",
  57113=>"011000111",
  57114=>"111100001",
  57115=>"000000010",
  57116=>"100000000",
  57117=>"101011101",
  57118=>"111111111",
  57119=>"011001100",
  57120=>"101110111",
  57121=>"010110111",
  57122=>"000001110",
  57123=>"101010101",
  57124=>"111101100",
  57125=>"111000101",
  57126=>"100110011",
  57127=>"010010000",
  57128=>"100000000",
  57129=>"000101010",
  57130=>"000011001",
  57131=>"001110110",
  57132=>"111101001",
  57133=>"000000011",
  57134=>"001010001",
  57135=>"101111110",
  57136=>"000001100",
  57137=>"100100110",
  57138=>"000001011",
  57139=>"001010010",
  57140=>"011001000",
  57141=>"110001011",
  57142=>"001100111",
  57143=>"011100001",
  57144=>"011110110",
  57145=>"110010010",
  57146=>"010100010",
  57147=>"100000101",
  57148=>"111111100",
  57149=>"000000000",
  57150=>"010000011",
  57151=>"010010100",
  57152=>"000110011",
  57153=>"110110111",
  57154=>"011000000",
  57155=>"101100100",
  57156=>"001011010",
  57157=>"110010000",
  57158=>"101001010",
  57159=>"110101001",
  57160=>"010000111",
  57161=>"110111111",
  57162=>"011000110",
  57163=>"000100010",
  57164=>"000000111",
  57165=>"001001110",
  57166=>"101000101",
  57167=>"101010000",
  57168=>"111101011",
  57169=>"110111111",
  57170=>"110100000",
  57171=>"000000001",
  57172=>"101101011",
  57173=>"111110100",
  57174=>"001100001",
  57175=>"011011100",
  57176=>"110001101",
  57177=>"101010001",
  57178=>"001111101",
  57179=>"011010101",
  57180=>"010111110",
  57181=>"001100100",
  57182=>"110000111",
  57183=>"001011110",
  57184=>"010110001",
  57185=>"000011010",
  57186=>"010001111",
  57187=>"110111000",
  57188=>"001011001",
  57189=>"000110111",
  57190=>"110101011",
  57191=>"110001000",
  57192=>"111001010",
  57193=>"111111010",
  57194=>"011010001",
  57195=>"000100011",
  57196=>"000010110",
  57197=>"100100011",
  57198=>"100110100",
  57199=>"111010110",
  57200=>"011011110",
  57201=>"111111100",
  57202=>"001000100",
  57203=>"010011001",
  57204=>"000000000",
  57205=>"000101000",
  57206=>"100000100",
  57207=>"100010000",
  57208=>"001000011",
  57209=>"100011100",
  57210=>"110001010",
  57211=>"111111101",
  57212=>"101011110",
  57213=>"010000101",
  57214=>"011011010",
  57215=>"110100010",
  57216=>"101101111",
  57217=>"110100111",
  57218=>"011001000",
  57219=>"111101100",
  57220=>"011011000",
  57221=>"111100110",
  57222=>"001010010",
  57223=>"111110111",
  57224=>"000011110",
  57225=>"001001011",
  57226=>"010111000",
  57227=>"100000010",
  57228=>"010010100",
  57229=>"101011110",
  57230=>"001011111",
  57231=>"001010111",
  57232=>"010000011",
  57233=>"110010010",
  57234=>"101110101",
  57235=>"111101100",
  57236=>"011010011",
  57237=>"111111101",
  57238=>"001001111",
  57239=>"011100101",
  57240=>"001101000",
  57241=>"010000000",
  57242=>"100111010",
  57243=>"110111011",
  57244=>"001111110",
  57245=>"010110110",
  57246=>"110101001",
  57247=>"100100100",
  57248=>"000001111",
  57249=>"000100111",
  57250=>"111010000",
  57251=>"101110110",
  57252=>"101100110",
  57253=>"010111111",
  57254=>"000110000",
  57255=>"100101110",
  57256=>"001001001",
  57257=>"000011010",
  57258=>"001110110",
  57259=>"111110101",
  57260=>"111000010",
  57261=>"000101011",
  57262=>"110100010",
  57263=>"110101001",
  57264=>"111100111",
  57265=>"000111010",
  57266=>"100101011",
  57267=>"100000000",
  57268=>"000000101",
  57269=>"101011011",
  57270=>"110100110",
  57271=>"000011110",
  57272=>"110111001",
  57273=>"110111101",
  57274=>"000100010",
  57275=>"001010000",
  57276=>"110111111",
  57277=>"111010111",
  57278=>"110111011",
  57279=>"100011000",
  57280=>"110001111",
  57281=>"010101000",
  57282=>"110101101",
  57283=>"101000011",
  57284=>"010110101",
  57285=>"111000000",
  57286=>"100001010",
  57287=>"110111011",
  57288=>"010101000",
  57289=>"011101111",
  57290=>"110110100",
  57291=>"101101101",
  57292=>"101100011",
  57293=>"011000000",
  57294=>"100111000",
  57295=>"101110010",
  57296=>"110100000",
  57297=>"110110000",
  57298=>"111011001",
  57299=>"010010100",
  57300=>"101001100",
  57301=>"001001010",
  57302=>"011100111",
  57303=>"010110011",
  57304=>"100001010",
  57305=>"001110111",
  57306=>"110111010",
  57307=>"001110000",
  57308=>"001011110",
  57309=>"001100001",
  57310=>"001011001",
  57311=>"010111010",
  57312=>"000111111",
  57313=>"001000010",
  57314=>"111110011",
  57315=>"101111001",
  57316=>"100000001",
  57317=>"111110111",
  57318=>"000101000",
  57319=>"001110001",
  57320=>"100001000",
  57321=>"000001111",
  57322=>"000100100",
  57323=>"010100100",
  57324=>"110110101",
  57325=>"011001000",
  57326=>"100100111",
  57327=>"011010110",
  57328=>"100010110",
  57329=>"101111001",
  57330=>"001110011",
  57331=>"101000111",
  57332=>"101001110",
  57333=>"011010000",
  57334=>"100111001",
  57335=>"100101111",
  57336=>"001000110",
  57337=>"101011111",
  57338=>"001010111",
  57339=>"100111100",
  57340=>"101000101",
  57341=>"111000000",
  57342=>"100100011",
  57343=>"000001001",
  57344=>"001001011",
  57345=>"000011001",
  57346=>"111111110",
  57347=>"000001011",
  57348=>"000100010",
  57349=>"000111010",
  57350=>"000010101",
  57351=>"101101001",
  57352=>"010011010",
  57353=>"101000010",
  57354=>"110111100",
  57355=>"101000100",
  57356=>"011111100",
  57357=>"100111001",
  57358=>"101110000",
  57359=>"101101110",
  57360=>"000000110",
  57361=>"001111111",
  57362=>"000110110",
  57363=>"110111101",
  57364=>"010000100",
  57365=>"100100100",
  57366=>"011100100",
  57367=>"001101001",
  57368=>"100000011",
  57369=>"011111001",
  57370=>"100000101",
  57371=>"001010111",
  57372=>"100110100",
  57373=>"011010011",
  57374=>"111010001",
  57375=>"010010000",
  57376=>"100100001",
  57377=>"011110010",
  57378=>"010100011",
  57379=>"000010101",
  57380=>"110001001",
  57381=>"100110100",
  57382=>"110010100",
  57383=>"010111000",
  57384=>"010000100",
  57385=>"100011000",
  57386=>"001011100",
  57387=>"011011100",
  57388=>"111100010",
  57389=>"011000111",
  57390=>"100101110",
  57391=>"010101110",
  57392=>"111001101",
  57393=>"100010011",
  57394=>"101110111",
  57395=>"110111011",
  57396=>"101100000",
  57397=>"011010010",
  57398=>"001010111",
  57399=>"110011011",
  57400=>"111111110",
  57401=>"001110100",
  57402=>"111101011",
  57403=>"100111001",
  57404=>"110000010",
  57405=>"010100101",
  57406=>"101011100",
  57407=>"001000000",
  57408=>"110101010",
  57409=>"111001001",
  57410=>"011100000",
  57411=>"001000101",
  57412=>"000101001",
  57413=>"110111001",
  57414=>"100011101",
  57415=>"011100110",
  57416=>"111111011",
  57417=>"001010000",
  57418=>"010000000",
  57419=>"110100101",
  57420=>"110001111",
  57421=>"001010110",
  57422=>"110000000",
  57423=>"000011110",
  57424=>"010110001",
  57425=>"110011011",
  57426=>"111011101",
  57427=>"000111111",
  57428=>"110110001",
  57429=>"101100110",
  57430=>"010101011",
  57431=>"000000001",
  57432=>"001000101",
  57433=>"110101001",
  57434=>"101000001",
  57435=>"011000000",
  57436=>"110011011",
  57437=>"001000111",
  57438=>"001001001",
  57439=>"100000011",
  57440=>"100101000",
  57441=>"001001111",
  57442=>"101110101",
  57443=>"110000001",
  57444=>"101110010",
  57445=>"110111010",
  57446=>"110001110",
  57447=>"110001011",
  57448=>"001101100",
  57449=>"110101110",
  57450=>"101010100",
  57451=>"001110001",
  57452=>"101011001",
  57453=>"100100100",
  57454=>"111011011",
  57455=>"001100001",
  57456=>"100101001",
  57457=>"010111011",
  57458=>"011011111",
  57459=>"010111001",
  57460=>"100011011",
  57461=>"000110010",
  57462=>"011111000",
  57463=>"111100111",
  57464=>"001001001",
  57465=>"110111111",
  57466=>"010101000",
  57467=>"011000000",
  57468=>"001110011",
  57469=>"000000111",
  57470=>"101101010",
  57471=>"101001111",
  57472=>"110111001",
  57473=>"101011110",
  57474=>"010000001",
  57475=>"110010100",
  57476=>"000000000",
  57477=>"010101011",
  57478=>"010010111",
  57479=>"000110101",
  57480=>"011110100",
  57481=>"000011000",
  57482=>"010010100",
  57483=>"101001000",
  57484=>"100001011",
  57485=>"011011110",
  57486=>"111010000",
  57487=>"000001001",
  57488=>"110110011",
  57489=>"000100110",
  57490=>"101011111",
  57491=>"000011100",
  57492=>"001010111",
  57493=>"100100000",
  57494=>"000110010",
  57495=>"100110110",
  57496=>"111100101",
  57497=>"000000001",
  57498=>"011001111",
  57499=>"001001110",
  57500=>"110001010",
  57501=>"101000010",
  57502=>"000111011",
  57503=>"101100100",
  57504=>"111100010",
  57505=>"110010111",
  57506=>"110101011",
  57507=>"010010000",
  57508=>"010111111",
  57509=>"100100011",
  57510=>"000110001",
  57511=>"010110001",
  57512=>"111011001",
  57513=>"011110010",
  57514=>"000001000",
  57515=>"010000100",
  57516=>"011110000",
  57517=>"000010111",
  57518=>"101111111",
  57519=>"101100001",
  57520=>"110000010",
  57521=>"011100000",
  57522=>"110000001",
  57523=>"110101100",
  57524=>"011011011",
  57525=>"000011000",
  57526=>"110000110",
  57527=>"111111100",
  57528=>"000110010",
  57529=>"101110111",
  57530=>"000110000",
  57531=>"010011010",
  57532=>"110110010",
  57533=>"001111000",
  57534=>"011000110",
  57535=>"000110101",
  57536=>"000000001",
  57537=>"001111101",
  57538=>"010100110",
  57539=>"110101110",
  57540=>"000001100",
  57541=>"111000110",
  57542=>"000000010",
  57543=>"110010111",
  57544=>"010100010",
  57545=>"111010110",
  57546=>"100001110",
  57547=>"110111100",
  57548=>"100101100",
  57549=>"011110101",
  57550=>"110011000",
  57551=>"001110110",
  57552=>"010111110",
  57553=>"111010111",
  57554=>"010000110",
  57555=>"111000010",
  57556=>"010101010",
  57557=>"101111110",
  57558=>"011011111",
  57559=>"101100101",
  57560=>"101100101",
  57561=>"000001011",
  57562=>"000110110",
  57563=>"101100011",
  57564=>"011111001",
  57565=>"010111011",
  57566=>"010111100",
  57567=>"101111011",
  57568=>"101111011",
  57569=>"011010011",
  57570=>"001000110",
  57571=>"111000000",
  57572=>"001100111",
  57573=>"101111110",
  57574=>"101100111",
  57575=>"011001110",
  57576=>"101101010",
  57577=>"100111011",
  57578=>"010010100",
  57579=>"010111110",
  57580=>"101111001",
  57581=>"111100000",
  57582=>"010001101",
  57583=>"111101000",
  57584=>"001011001",
  57585=>"000101110",
  57586=>"110111110",
  57587=>"101010001",
  57588=>"010101111",
  57589=>"000111101",
  57590=>"100111101",
  57591=>"111110110",
  57592=>"010000100",
  57593=>"010010011",
  57594=>"101101010",
  57595=>"100010101",
  57596=>"000010111",
  57597=>"001101100",
  57598=>"001110100",
  57599=>"001001000",
  57600=>"000000100",
  57601=>"111111111",
  57602=>"000100000",
  57603=>"111001100",
  57604=>"000110110",
  57605=>"001001011",
  57606=>"110111001",
  57607=>"110110000",
  57608=>"011001100",
  57609=>"011101001",
  57610=>"100101000",
  57611=>"001000101",
  57612=>"100101000",
  57613=>"011101100",
  57614=>"101110101",
  57615=>"100110101",
  57616=>"111010001",
  57617=>"100101001",
  57618=>"011111100",
  57619=>"011010110",
  57620=>"111110000",
  57621=>"101110001",
  57622=>"000111011",
  57623=>"100100110",
  57624=>"010111100",
  57625=>"010110001",
  57626=>"000100011",
  57627=>"010000001",
  57628=>"010011010",
  57629=>"110111111",
  57630=>"011111001",
  57631=>"011011001",
  57632=>"000000110",
  57633=>"001010100",
  57634=>"001010110",
  57635=>"111100011",
  57636=>"110101101",
  57637=>"010001000",
  57638=>"100000110",
  57639=>"010000100",
  57640=>"101001011",
  57641=>"011111011",
  57642=>"011110111",
  57643=>"110000100",
  57644=>"001100001",
  57645=>"000000100",
  57646=>"000000001",
  57647=>"110110111",
  57648=>"011000101",
  57649=>"101011010",
  57650=>"000010010",
  57651=>"111101101",
  57652=>"100001000",
  57653=>"010000100",
  57654=>"111011111",
  57655=>"001001010",
  57656=>"011000001",
  57657=>"100001110",
  57658=>"000111101",
  57659=>"111110001",
  57660=>"110011010",
  57661=>"011100101",
  57662=>"010011000",
  57663=>"011101011",
  57664=>"001001001",
  57665=>"111101001",
  57666=>"010011011",
  57667=>"011110101",
  57668=>"000100110",
  57669=>"011000010",
  57670=>"101101101",
  57671=>"100000100",
  57672=>"001001000",
  57673=>"110001101",
  57674=>"110100111",
  57675=>"010010100",
  57676=>"001100101",
  57677=>"001011110",
  57678=>"001100000",
  57679=>"000001101",
  57680=>"111110010",
  57681=>"101101101",
  57682=>"110100001",
  57683=>"110111110",
  57684=>"111000001",
  57685=>"111111011",
  57686=>"101011001",
  57687=>"000110001",
  57688=>"010001011",
  57689=>"101011001",
  57690=>"000110000",
  57691=>"001110100",
  57692=>"100111001",
  57693=>"000001000",
  57694=>"100100000",
  57695=>"000111110",
  57696=>"000100111",
  57697=>"111011000",
  57698=>"111111100",
  57699=>"001000111",
  57700=>"110010101",
  57701=>"110011110",
  57702=>"001111111",
  57703=>"100011111",
  57704=>"010110011",
  57705=>"110001110",
  57706=>"111010100",
  57707=>"010011011",
  57708=>"011010110",
  57709=>"010011000",
  57710=>"111101101",
  57711=>"110010011",
  57712=>"101011111",
  57713=>"001111101",
  57714=>"001010111",
  57715=>"000111010",
  57716=>"010110010",
  57717=>"001111010",
  57718=>"010110110",
  57719=>"111110011",
  57720=>"000100010",
  57721=>"000010111",
  57722=>"110100100",
  57723=>"010110010",
  57724=>"011111000",
  57725=>"010011110",
  57726=>"000110111",
  57727=>"000100111",
  57728=>"100010110",
  57729=>"001010000",
  57730=>"001111110",
  57731=>"100100101",
  57732=>"000011101",
  57733=>"000000101",
  57734=>"111001011",
  57735=>"110011110",
  57736=>"111001000",
  57737=>"001000101",
  57738=>"100111100",
  57739=>"110000111",
  57740=>"110100101",
  57741=>"111110100",
  57742=>"110010010",
  57743=>"101001001",
  57744=>"111111100",
  57745=>"100110001",
  57746=>"000101101",
  57747=>"101001010",
  57748=>"100010010",
  57749=>"100011100",
  57750=>"101111100",
  57751=>"001110110",
  57752=>"101010001",
  57753=>"000011010",
  57754=>"001010001",
  57755=>"011011010",
  57756=>"001011111",
  57757=>"000101111",
  57758=>"111001101",
  57759=>"111000111",
  57760=>"101111000",
  57761=>"011111111",
  57762=>"010001000",
  57763=>"111011100",
  57764=>"100101101",
  57765=>"010000011",
  57766=>"000001100",
  57767=>"110101011",
  57768=>"010101000",
  57769=>"001100000",
  57770=>"000011111",
  57771=>"001000110",
  57772=>"011000001",
  57773=>"000100111",
  57774=>"001011111",
  57775=>"010010000",
  57776=>"000100001",
  57777=>"000011111",
  57778=>"000010100",
  57779=>"000011110",
  57780=>"000010010",
  57781=>"111000111",
  57782=>"000111010",
  57783=>"111010110",
  57784=>"001010001",
  57785=>"110000001",
  57786=>"001001000",
  57787=>"110010100",
  57788=>"110010001",
  57789=>"111111001",
  57790=>"011100100",
  57791=>"001001111",
  57792=>"110010000",
  57793=>"100011001",
  57794=>"100010111",
  57795=>"101101111",
  57796=>"000011000",
  57797=>"011101100",
  57798=>"000101010",
  57799=>"111001001",
  57800=>"110111000",
  57801=>"001000001",
  57802=>"010011011",
  57803=>"011110010",
  57804=>"000001000",
  57805=>"110000001",
  57806=>"000000100",
  57807=>"011011101",
  57808=>"100000110",
  57809=>"010101000",
  57810=>"101011100",
  57811=>"100011111",
  57812=>"100011110",
  57813=>"100101100",
  57814=>"011001110",
  57815=>"010110011",
  57816=>"011001101",
  57817=>"010101000",
  57818=>"110001001",
  57819=>"101010110",
  57820=>"111000010",
  57821=>"011111111",
  57822=>"101010011",
  57823=>"011101011",
  57824=>"101000101",
  57825=>"111011001",
  57826=>"101111001",
  57827=>"000101101",
  57828=>"001011101",
  57829=>"110100000",
  57830=>"100000100",
  57831=>"111001001",
  57832=>"010011000",
  57833=>"100111100",
  57834=>"000010000",
  57835=>"110010011",
  57836=>"000001011",
  57837=>"110000000",
  57838=>"110100100",
  57839=>"101011010",
  57840=>"000011001",
  57841=>"100110101",
  57842=>"001000001",
  57843=>"011000000",
  57844=>"101111011",
  57845=>"101001111",
  57846=>"000000100",
  57847=>"110101001",
  57848=>"010110011",
  57849=>"011001100",
  57850=>"110001111",
  57851=>"101000010",
  57852=>"101001001",
  57853=>"110011010",
  57854=>"111100100",
  57855=>"010001011",
  57856=>"111101110",
  57857=>"100100100",
  57858=>"111011001",
  57859=>"101000010",
  57860=>"010101001",
  57861=>"011010011",
  57862=>"101100110",
  57863=>"110000011",
  57864=>"011101111",
  57865=>"001001110",
  57866=>"001100100",
  57867=>"010110110",
  57868=>"000001101",
  57869=>"101010111",
  57870=>"111010010",
  57871=>"000001101",
  57872=>"101100101",
  57873=>"110010110",
  57874=>"011100110",
  57875=>"111011000",
  57876=>"010010010",
  57877=>"110101100",
  57878=>"011000011",
  57879=>"111001000",
  57880=>"010011011",
  57881=>"001001010",
  57882=>"010011000",
  57883=>"101010100",
  57884=>"000011110",
  57885=>"010000010",
  57886=>"110111101",
  57887=>"001000101",
  57888=>"101011100",
  57889=>"101001101",
  57890=>"011011000",
  57891=>"110111010",
  57892=>"001000011",
  57893=>"101001011",
  57894=>"101001111",
  57895=>"111110011",
  57896=>"000010000",
  57897=>"100101011",
  57898=>"010101000",
  57899=>"010100010",
  57900=>"010100111",
  57901=>"100101011",
  57902=>"010010111",
  57903=>"011010110",
  57904=>"000110110",
  57905=>"001001001",
  57906=>"111000010",
  57907=>"001100111",
  57908=>"111001000",
  57909=>"110000000",
  57910=>"011111110",
  57911=>"101101001",
  57912=>"111111100",
  57913=>"101010110",
  57914=>"101110001",
  57915=>"000100100",
  57916=>"010110010",
  57917=>"001110001",
  57918=>"100001000",
  57919=>"110100111",
  57920=>"010001011",
  57921=>"101110111",
  57922=>"111101111",
  57923=>"111101110",
  57924=>"101000111",
  57925=>"001100011",
  57926=>"011100101",
  57927=>"011001000",
  57928=>"010011011",
  57929=>"110010011",
  57930=>"111111100",
  57931=>"110101011",
  57932=>"100000100",
  57933=>"100001100",
  57934=>"000101100",
  57935=>"001000010",
  57936=>"001000010",
  57937=>"011100111",
  57938=>"000001000",
  57939=>"110001110",
  57940=>"101000111",
  57941=>"010000000",
  57942=>"010001100",
  57943=>"101101101",
  57944=>"011100111",
  57945=>"011100100",
  57946=>"101111011",
  57947=>"011101111",
  57948=>"110100010",
  57949=>"001000000",
  57950=>"111010011",
  57951=>"001000110",
  57952=>"000111111",
  57953=>"101101100",
  57954=>"010010111",
  57955=>"001101101",
  57956=>"100000001",
  57957=>"100111111",
  57958=>"000101010",
  57959=>"010110101",
  57960=>"001100100",
  57961=>"101101010",
  57962=>"110000101",
  57963=>"101000000",
  57964=>"001011101",
  57965=>"101101100",
  57966=>"001101001",
  57967=>"010110001",
  57968=>"100001000",
  57969=>"001000000",
  57970=>"110101111",
  57971=>"100110001",
  57972=>"110111110",
  57973=>"110000000",
  57974=>"010000010",
  57975=>"111010111",
  57976=>"110111010",
  57977=>"000101010",
  57978=>"110000111",
  57979=>"011100001",
  57980=>"100010011",
  57981=>"000110111",
  57982=>"111100000",
  57983=>"100001001",
  57984=>"111111101",
  57985=>"101100011",
  57986=>"001111001",
  57987=>"100100011",
  57988=>"100000000",
  57989=>"100000001",
  57990=>"001101011",
  57991=>"011111100",
  57992=>"111101111",
  57993=>"111110010",
  57994=>"111101010",
  57995=>"011100100",
  57996=>"001101111",
  57997=>"100000110",
  57998=>"000100010",
  57999=>"001011011",
  58000=>"101101111",
  58001=>"101011100",
  58002=>"101110111",
  58003=>"011011000",
  58004=>"101101000",
  58005=>"110011101",
  58006=>"011011111",
  58007=>"011011001",
  58008=>"100100011",
  58009=>"100101110",
  58010=>"001101100",
  58011=>"101010110",
  58012=>"100111110",
  58013=>"001110011",
  58014=>"001011111",
  58015=>"100101110",
  58016=>"100111110",
  58017=>"101100011",
  58018=>"110011101",
  58019=>"111000100",
  58020=>"111011100",
  58021=>"101100001",
  58022=>"110110000",
  58023=>"001000000",
  58024=>"001001000",
  58025=>"100100110",
  58026=>"110001110",
  58027=>"011100000",
  58028=>"000000100",
  58029=>"011011010",
  58030=>"111001111",
  58031=>"000110001",
  58032=>"011010010",
  58033=>"101100001",
  58034=>"000001100",
  58035=>"100010100",
  58036=>"010000010",
  58037=>"101010101",
  58038=>"000001101",
  58039=>"001010000",
  58040=>"000100100",
  58041=>"001101010",
  58042=>"010111010",
  58043=>"101011000",
  58044=>"110001100",
  58045=>"100111000",
  58046=>"011101000",
  58047=>"010000100",
  58048=>"111101100",
  58049=>"011011110",
  58050=>"001010101",
  58051=>"110011001",
  58052=>"110101111",
  58053=>"101111011",
  58054=>"111001010",
  58055=>"110101100",
  58056=>"000010000",
  58057=>"000101000",
  58058=>"011010001",
  58059=>"001001010",
  58060=>"101010011",
  58061=>"100111111",
  58062=>"110000011",
  58063=>"101001001",
  58064=>"000011000",
  58065=>"001011001",
  58066=>"000001101",
  58067=>"000011110",
  58068=>"000100101",
  58069=>"011000100",
  58070=>"011011011",
  58071=>"111001000",
  58072=>"111111100",
  58073=>"001001110",
  58074=>"010000000",
  58075=>"100010000",
  58076=>"100101111",
  58077=>"111011011",
  58078=>"001000111",
  58079=>"010101100",
  58080=>"000010101",
  58081=>"100000010",
  58082=>"010011111",
  58083=>"001111100",
  58084=>"011100010",
  58085=>"011100111",
  58086=>"100100000",
  58087=>"010010111",
  58088=>"000100000",
  58089=>"101001110",
  58090=>"000100010",
  58091=>"010010011",
  58092=>"000011001",
  58093=>"101010101",
  58094=>"101000010",
  58095=>"111000101",
  58096=>"010110111",
  58097=>"100100001",
  58098=>"000111100",
  58099=>"100111111",
  58100=>"000000011",
  58101=>"100011101",
  58102=>"111100001",
  58103=>"010101100",
  58104=>"100010001",
  58105=>"000111010",
  58106=>"111110001",
  58107=>"111010000",
  58108=>"011111011",
  58109=>"100010000",
  58110=>"001001001",
  58111=>"000111001",
  58112=>"011111010",
  58113=>"111011011",
  58114=>"000111100",
  58115=>"111010111",
  58116=>"101011000",
  58117=>"000000000",
  58118=>"111010100",
  58119=>"010010100",
  58120=>"110000101",
  58121=>"011010111",
  58122=>"011111100",
  58123=>"001011101",
  58124=>"111010010",
  58125=>"011010110",
  58126=>"100000010",
  58127=>"111000001",
  58128=>"101110100",
  58129=>"000111010",
  58130=>"111011110",
  58131=>"010001101",
  58132=>"011011000",
  58133=>"010100101",
  58134=>"110000010",
  58135=>"000110110",
  58136=>"001011011",
  58137=>"000000101",
  58138=>"010111111",
  58139=>"100101101",
  58140=>"000011100",
  58141=>"110100100",
  58142=>"111000000",
  58143=>"000001101",
  58144=>"110011100",
  58145=>"100011010",
  58146=>"000001110",
  58147=>"010010011",
  58148=>"010010000",
  58149=>"001000000",
  58150=>"011111100",
  58151=>"110111010",
  58152=>"101110110",
  58153=>"110001011",
  58154=>"101000000",
  58155=>"100101110",
  58156=>"111101001",
  58157=>"100010011",
  58158=>"100011010",
  58159=>"110101110",
  58160=>"100010100",
  58161=>"110011010",
  58162=>"010000101",
  58163=>"111111000",
  58164=>"010100011",
  58165=>"110011011",
  58166=>"001001100",
  58167=>"001110111",
  58168=>"100010010",
  58169=>"101110101",
  58170=>"111100001",
  58171=>"111001001",
  58172=>"111111001",
  58173=>"011001000",
  58174=>"010001110",
  58175=>"010001110",
  58176=>"101010001",
  58177=>"101000111",
  58178=>"000001110",
  58179=>"000101110",
  58180=>"100001000",
  58181=>"111101100",
  58182=>"111111011",
  58183=>"001110001",
  58184=>"010111001",
  58185=>"101010111",
  58186=>"001101101",
  58187=>"011101011",
  58188=>"100101000",
  58189=>"000101101",
  58190=>"100001000",
  58191=>"000000100",
  58192=>"000111100",
  58193=>"001000001",
  58194=>"110100001",
  58195=>"011100011",
  58196=>"110101110",
  58197=>"001111111",
  58198=>"011001001",
  58199=>"010110010",
  58200=>"111110011",
  58201=>"011111001",
  58202=>"101100000",
  58203=>"011101000",
  58204=>"000011100",
  58205=>"011011100",
  58206=>"100101111",
  58207=>"010100101",
  58208=>"000001101",
  58209=>"001010111",
  58210=>"010000000",
  58211=>"000010010",
  58212=>"011100111",
  58213=>"111010001",
  58214=>"110100101",
  58215=>"001111111",
  58216=>"100101110",
  58217=>"101111111",
  58218=>"100111100",
  58219=>"000011111",
  58220=>"011111001",
  58221=>"000001000",
  58222=>"111011001",
  58223=>"111101011",
  58224=>"100001111",
  58225=>"010001111",
  58226=>"011111011",
  58227=>"111011011",
  58228=>"100101110",
  58229=>"111001011",
  58230=>"000010010",
  58231=>"001000101",
  58232=>"101010000",
  58233=>"010011100",
  58234=>"000011101",
  58235=>"110110110",
  58236=>"010001000",
  58237=>"111010110",
  58238=>"001010000",
  58239=>"100100010",
  58240=>"000000010",
  58241=>"010001111",
  58242=>"001010111",
  58243=>"101101000",
  58244=>"011010000",
  58245=>"110000110",
  58246=>"000110010",
  58247=>"011001010",
  58248=>"110000111",
  58249=>"000101100",
  58250=>"111011001",
  58251=>"001111000",
  58252=>"001000001",
  58253=>"010011101",
  58254=>"101111110",
  58255=>"011001110",
  58256=>"000110011",
  58257=>"110000011",
  58258=>"000001000",
  58259=>"000100100",
  58260=>"100101111",
  58261=>"101101111",
  58262=>"101110000",
  58263=>"001100010",
  58264=>"000000110",
  58265=>"010111101",
  58266=>"000101101",
  58267=>"110011010",
  58268=>"100011011",
  58269=>"001010101",
  58270=>"011100010",
  58271=>"111010011",
  58272=>"110101010",
  58273=>"101010001",
  58274=>"111101101",
  58275=>"101111001",
  58276=>"011001000",
  58277=>"111101011",
  58278=>"000000010",
  58279=>"100100111",
  58280=>"010011101",
  58281=>"111111111",
  58282=>"111110110",
  58283=>"101011011",
  58284=>"001100110",
  58285=>"101001000",
  58286=>"010000000",
  58287=>"111001011",
  58288=>"010100101",
  58289=>"101000011",
  58290=>"100111100",
  58291=>"001111110",
  58292=>"111100000",
  58293=>"110001101",
  58294=>"101101110",
  58295=>"000011111",
  58296=>"111001110",
  58297=>"000110100",
  58298=>"000010010",
  58299=>"111000010",
  58300=>"101100010",
  58301=>"001111011",
  58302=>"011000111",
  58303=>"010001000",
  58304=>"010001000",
  58305=>"000100101",
  58306=>"101001010",
  58307=>"100110111",
  58308=>"001100001",
  58309=>"110110010",
  58310=>"100100011",
  58311=>"011001001",
  58312=>"100101101",
  58313=>"100001001",
  58314=>"001101011",
  58315=>"101111101",
  58316=>"101010110",
  58317=>"000001110",
  58318=>"000110000",
  58319=>"110101110",
  58320=>"100010011",
  58321=>"100010110",
  58322=>"111010100",
  58323=>"000100101",
  58324=>"000101010",
  58325=>"100000000",
  58326=>"110000001",
  58327=>"101100100",
  58328=>"111111100",
  58329=>"000011111",
  58330=>"000111111",
  58331=>"001001001",
  58332=>"001001110",
  58333=>"011111111",
  58334=>"000110000",
  58335=>"010011000",
  58336=>"100111100",
  58337=>"001010000",
  58338=>"101110010",
  58339=>"010010101",
  58340=>"000111000",
  58341=>"111011110",
  58342=>"010001010",
  58343=>"100110101",
  58344=>"000100010",
  58345=>"011101111",
  58346=>"101011100",
  58347=>"101110100",
  58348=>"111100101",
  58349=>"111111000",
  58350=>"011111000",
  58351=>"101110001",
  58352=>"111101010",
  58353=>"000000011",
  58354=>"100010101",
  58355=>"010111000",
  58356=>"111011100",
  58357=>"000100001",
  58358=>"101001010",
  58359=>"000100101",
  58360=>"100100101",
  58361=>"101011010",
  58362=>"100010000",
  58363=>"101111101",
  58364=>"000010001",
  58365=>"010011010",
  58366=>"101111000",
  58367=>"101101101",
  58368=>"010011000",
  58369=>"000110010",
  58370=>"011010000",
  58371=>"100101001",
  58372=>"011110100",
  58373=>"000000111",
  58374=>"100010010",
  58375=>"011111110",
  58376=>"001000101",
  58377=>"011011001",
  58378=>"000110000",
  58379=>"011011101",
  58380=>"100111011",
  58381=>"011100001",
  58382=>"011010100",
  58383=>"010011000",
  58384=>"000111110",
  58385=>"100101010",
  58386=>"110100100",
  58387=>"011100110",
  58388=>"101101110",
  58389=>"000111011",
  58390=>"001101101",
  58391=>"111100010",
  58392=>"010101110",
  58393=>"101111101",
  58394=>"010001110",
  58395=>"110011110",
  58396=>"011110111",
  58397=>"011101100",
  58398=>"101110100",
  58399=>"101100100",
  58400=>"101000101",
  58401=>"011001011",
  58402=>"010110101",
  58403=>"011000011",
  58404=>"101011111",
  58405=>"111100000",
  58406=>"111110110",
  58407=>"110100100",
  58408=>"001101100",
  58409=>"010001001",
  58410=>"001110101",
  58411=>"010011010",
  58412=>"111111111",
  58413=>"011011101",
  58414=>"000110001",
  58415=>"101110001",
  58416=>"110011101",
  58417=>"111010011",
  58418=>"111011000",
  58419=>"011101001",
  58420=>"001000100",
  58421=>"011101111",
  58422=>"110101010",
  58423=>"101100000",
  58424=>"001001001",
  58425=>"011001101",
  58426=>"001000010",
  58427=>"000100100",
  58428=>"010010001",
  58429=>"111100000",
  58430=>"001011110",
  58431=>"001111011",
  58432=>"111101100",
  58433=>"000100000",
  58434=>"100101101",
  58435=>"001100011",
  58436=>"110000000",
  58437=>"111001000",
  58438=>"100001001",
  58439=>"100000100",
  58440=>"011011011",
  58441=>"010110111",
  58442=>"001010101",
  58443=>"111100111",
  58444=>"010001000",
  58445=>"110010001",
  58446=>"110000111",
  58447=>"111001001",
  58448=>"001100100",
  58449=>"110100100",
  58450=>"000001101",
  58451=>"000111001",
  58452=>"110111101",
  58453=>"001001111",
  58454=>"001000001",
  58455=>"010101001",
  58456=>"101100111",
  58457=>"011100000",
  58458=>"111011010",
  58459=>"011111100",
  58460=>"101001001",
  58461=>"000111000",
  58462=>"111111010",
  58463=>"000101110",
  58464=>"111000011",
  58465=>"111111100",
  58466=>"000111101",
  58467=>"010100101",
  58468=>"101110111",
  58469=>"011111100",
  58470=>"110000010",
  58471=>"010011101",
  58472=>"010001111",
  58473=>"111100010",
  58474=>"111101010",
  58475=>"100010110",
  58476=>"101001011",
  58477=>"000110100",
  58478=>"001100011",
  58479=>"000101000",
  58480=>"011101111",
  58481=>"111110110",
  58482=>"111100011",
  58483=>"101010000",
  58484=>"010101101",
  58485=>"010110000",
  58486=>"101010111",
  58487=>"111011111",
  58488=>"101011000",
  58489=>"011010010",
  58490=>"000101101",
  58491=>"010010000",
  58492=>"001111011",
  58493=>"000101100",
  58494=>"000010000",
  58495=>"010010111",
  58496=>"001010000",
  58497=>"000011010",
  58498=>"111110011",
  58499=>"110101111",
  58500=>"110010011",
  58501=>"001100001",
  58502=>"011101010",
  58503=>"001101100",
  58504=>"000001110",
  58505=>"010001011",
  58506=>"101010010",
  58507=>"100010111",
  58508=>"100110010",
  58509=>"010010110",
  58510=>"111110001",
  58511=>"100011110",
  58512=>"101111010",
  58513=>"100101101",
  58514=>"001100011",
  58515=>"001101111",
  58516=>"100100001",
  58517=>"110101111",
  58518=>"101110011",
  58519=>"011110110",
  58520=>"111010000",
  58521=>"110101100",
  58522=>"111010000",
  58523=>"000110011",
  58524=>"110000001",
  58525=>"011000101",
  58526=>"010011010",
  58527=>"111001100",
  58528=>"110011100",
  58529=>"001010100",
  58530=>"001000011",
  58531=>"010011101",
  58532=>"101110111",
  58533=>"001101111",
  58534=>"010011001",
  58535=>"110001010",
  58536=>"101011010",
  58537=>"010111010",
  58538=>"110110000",
  58539=>"010110010",
  58540=>"011000010",
  58541=>"110010001",
  58542=>"111000111",
  58543=>"101100110",
  58544=>"010001001",
  58545=>"110101010",
  58546=>"011000100",
  58547=>"111001000",
  58548=>"000110100",
  58549=>"111111101",
  58550=>"111001011",
  58551=>"110100111",
  58552=>"011010010",
  58553=>"010111110",
  58554=>"001100000",
  58555=>"010010100",
  58556=>"111101000",
  58557=>"000010010",
  58558=>"101001111",
  58559=>"111101101",
  58560=>"011101111",
  58561=>"000111101",
  58562=>"001100000",
  58563=>"001110101",
  58564=>"010101011",
  58565=>"101100111",
  58566=>"101000001",
  58567=>"111011111",
  58568=>"000001110",
  58569=>"011100111",
  58570=>"011111110",
  58571=>"000110100",
  58572=>"000101100",
  58573=>"001011110",
  58574=>"000101111",
  58575=>"111011001",
  58576=>"110100101",
  58577=>"010001111",
  58578=>"011000001",
  58579=>"110110100",
  58580=>"001001001",
  58581=>"011110011",
  58582=>"111101100",
  58583=>"100001110",
  58584=>"110101001",
  58585=>"110011100",
  58586=>"010010001",
  58587=>"101110011",
  58588=>"100101101",
  58589=>"001001111",
  58590=>"100011000",
  58591=>"001110100",
  58592=>"100010000",
  58593=>"111000011",
  58594=>"110101001",
  58595=>"101010101",
  58596=>"000001111",
  58597=>"010010111",
  58598=>"000110110",
  58599=>"001111001",
  58600=>"100001010",
  58601=>"000110011",
  58602=>"111010111",
  58603=>"111110111",
  58604=>"111011000",
  58605=>"000011110",
  58606=>"000010000",
  58607=>"000000001",
  58608=>"001100111",
  58609=>"111110110",
  58610=>"011001100",
  58611=>"110010011",
  58612=>"101110101",
  58613=>"010101101",
  58614=>"010011001",
  58615=>"110100010",
  58616=>"100010100",
  58617=>"010100011",
  58618=>"100101101",
  58619=>"100111000",
  58620=>"001011101",
  58621=>"100100111",
  58622=>"111000100",
  58623=>"101011110",
  58624=>"000001110",
  58625=>"010110101",
  58626=>"100011110",
  58627=>"001000101",
  58628=>"110011111",
  58629=>"101101001",
  58630=>"101100010",
  58631=>"110010111",
  58632=>"100001000",
  58633=>"000011100",
  58634=>"110110000",
  58635=>"001010100",
  58636=>"100010110",
  58637=>"111100000",
  58638=>"011001011",
  58639=>"101101001",
  58640=>"010111000",
  58641=>"011000111",
  58642=>"000011001",
  58643=>"100010101",
  58644=>"001100001",
  58645=>"010110101",
  58646=>"110000010",
  58647=>"000011011",
  58648=>"101011001",
  58649=>"100101110",
  58650=>"001111011",
  58651=>"110101100",
  58652=>"100000111",
  58653=>"011101010",
  58654=>"011110011",
  58655=>"100010010",
  58656=>"100101011",
  58657=>"000000001",
  58658=>"100001100",
  58659=>"010110010",
  58660=>"001101010",
  58661=>"011011111",
  58662=>"100011111",
  58663=>"100000101",
  58664=>"100011110",
  58665=>"100101110",
  58666=>"101000101",
  58667=>"101101110",
  58668=>"111011010",
  58669=>"011011000",
  58670=>"000101000",
  58671=>"111001111",
  58672=>"110110000",
  58673=>"011110101",
  58674=>"111111110",
  58675=>"000110110",
  58676=>"001100011",
  58677=>"010001000",
  58678=>"011010100",
  58679=>"110010101",
  58680=>"011100100",
  58681=>"011001000",
  58682=>"110110010",
  58683=>"011010100",
  58684=>"000100100",
  58685=>"011101100",
  58686=>"110011100",
  58687=>"011111110",
  58688=>"100101011",
  58689=>"101101101",
  58690=>"111111111",
  58691=>"100110011",
  58692=>"110100110",
  58693=>"011100101",
  58694=>"110000100",
  58695=>"001101011",
  58696=>"010100100",
  58697=>"010010000",
  58698=>"110110011",
  58699=>"100010110",
  58700=>"011010101",
  58701=>"101100010",
  58702=>"011001111",
  58703=>"110010100",
  58704=>"110001001",
  58705=>"100010111",
  58706=>"101101110",
  58707=>"000001010",
  58708=>"100101001",
  58709=>"110111100",
  58710=>"111111001",
  58711=>"010000100",
  58712=>"101111100",
  58713=>"100110010",
  58714=>"100101111",
  58715=>"001100011",
  58716=>"111100010",
  58717=>"011011000",
  58718=>"100111100",
  58719=>"110010011",
  58720=>"011011000",
  58721=>"001001111",
  58722=>"110000011",
  58723=>"101011001",
  58724=>"111011110",
  58725=>"101101111",
  58726=>"001000011",
  58727=>"111010110",
  58728=>"111011001",
  58729=>"110001000",
  58730=>"011011011",
  58731=>"110110110",
  58732=>"100111100",
  58733=>"111101100",
  58734=>"000010111",
  58735=>"111111100",
  58736=>"101100000",
  58737=>"010011011",
  58738=>"010001011",
  58739=>"001111000",
  58740=>"011101000",
  58741=>"010101010",
  58742=>"101001010",
  58743=>"001111011",
  58744=>"000000101",
  58745=>"001001011",
  58746=>"101000111",
  58747=>"111111001",
  58748=>"011100111",
  58749=>"101111111",
  58750=>"010011111",
  58751=>"000010010",
  58752=>"000100010",
  58753=>"000110001",
  58754=>"110111010",
  58755=>"000101101",
  58756=>"011101101",
  58757=>"101000000",
  58758=>"001100100",
  58759=>"000010110",
  58760=>"000101001",
  58761=>"101100101",
  58762=>"111001000",
  58763=>"100011110",
  58764=>"001011000",
  58765=>"000101101",
  58766=>"011110011",
  58767=>"101011011",
  58768=>"110100010",
  58769=>"100010011",
  58770=>"000000011",
  58771=>"111011111",
  58772=>"111111001",
  58773=>"010100011",
  58774=>"111000000",
  58775=>"011011101",
  58776=>"101100101",
  58777=>"011001100",
  58778=>"000111110",
  58779=>"111101110",
  58780=>"010110101",
  58781=>"111100001",
  58782=>"111010111",
  58783=>"000111111",
  58784=>"001001000",
  58785=>"100001001",
  58786=>"001110000",
  58787=>"010101101",
  58788=>"000010100",
  58789=>"001001100",
  58790=>"010010000",
  58791=>"001100011",
  58792=>"100111111",
  58793=>"110111000",
  58794=>"000110111",
  58795=>"010001100",
  58796=>"010011101",
  58797=>"001010010",
  58798=>"111101011",
  58799=>"110011000",
  58800=>"001000101",
  58801=>"010011011",
  58802=>"110101000",
  58803=>"111100101",
  58804=>"100011101",
  58805=>"100000111",
  58806=>"110100100",
  58807=>"111000111",
  58808=>"011000110",
  58809=>"100010010",
  58810=>"111010111",
  58811=>"010001001",
  58812=>"010111101",
  58813=>"111010000",
  58814=>"110000001",
  58815=>"101111100",
  58816=>"111001000",
  58817=>"101010100",
  58818=>"101000011",
  58819=>"011100001",
  58820=>"111010001",
  58821=>"010110000",
  58822=>"111111101",
  58823=>"100000000",
  58824=>"000010011",
  58825=>"101100011",
  58826=>"101000000",
  58827=>"000111111",
  58828=>"101001010",
  58829=>"100110011",
  58830=>"000111000",
  58831=>"000100011",
  58832=>"001101011",
  58833=>"100010100",
  58834=>"000111110",
  58835=>"110111001",
  58836=>"010001110",
  58837=>"101110101",
  58838=>"010110100",
  58839=>"010001001",
  58840=>"110001100",
  58841=>"001010111",
  58842=>"100110100",
  58843=>"111010000",
  58844=>"101001111",
  58845=>"101110000",
  58846=>"000101011",
  58847=>"011110011",
  58848=>"100010001",
  58849=>"000011001",
  58850=>"011111100",
  58851=>"100010000",
  58852=>"101010110",
  58853=>"110011010",
  58854=>"110110010",
  58855=>"001011000",
  58856=>"100111101",
  58857=>"001110101",
  58858=>"111011101",
  58859=>"100110001",
  58860=>"000110000",
  58861=>"001101000",
  58862=>"100111010",
  58863=>"110001000",
  58864=>"010110011",
  58865=>"100001011",
  58866=>"100110000",
  58867=>"100000001",
  58868=>"101110111",
  58869=>"111111000",
  58870=>"001101011",
  58871=>"001001000",
  58872=>"011001000",
  58873=>"101010111",
  58874=>"010001000",
  58875=>"110000000",
  58876=>"111010111",
  58877=>"000110001",
  58878=>"100001000",
  58879=>"000001111",
  58880=>"111110001",
  58881=>"100010100",
  58882=>"001011011",
  58883=>"000000110",
  58884=>"100110100",
  58885=>"010101111",
  58886=>"000011110",
  58887=>"000000000",
  58888=>"110010010",
  58889=>"001110110",
  58890=>"110011000",
  58891=>"111110010",
  58892=>"001110001",
  58893=>"001100000",
  58894=>"111000001",
  58895=>"111110100",
  58896=>"101011110",
  58897=>"010010101",
  58898=>"011000010",
  58899=>"001100000",
  58900=>"001001110",
  58901=>"111000010",
  58902=>"110001100",
  58903=>"011011000",
  58904=>"110010000",
  58905=>"000101001",
  58906=>"101100110",
  58907=>"010100110",
  58908=>"010001010",
  58909=>"111011110",
  58910=>"001011100",
  58911=>"000000010",
  58912=>"000010111",
  58913=>"001101111",
  58914=>"000001000",
  58915=>"010101100",
  58916=>"110101110",
  58917=>"011000001",
  58918=>"100010010",
  58919=>"111010011",
  58920=>"100110110",
  58921=>"001010100",
  58922=>"001100000",
  58923=>"111001101",
  58924=>"100101111",
  58925=>"101111101",
  58926=>"001000001",
  58927=>"101010010",
  58928=>"001110011",
  58929=>"001100110",
  58930=>"001101101",
  58931=>"110011010",
  58932=>"001100010",
  58933=>"110011101",
  58934=>"101010101",
  58935=>"001001001",
  58936=>"111010011",
  58937=>"000100000",
  58938=>"010001101",
  58939=>"111100010",
  58940=>"011010100",
  58941=>"011101010",
  58942=>"110101010",
  58943=>"001010100",
  58944=>"111000010",
  58945=>"001100100",
  58946=>"000010110",
  58947=>"010111010",
  58948=>"110010111",
  58949=>"101000000",
  58950=>"011001000",
  58951=>"010101110",
  58952=>"011100110",
  58953=>"100110111",
  58954=>"100110100",
  58955=>"110101110",
  58956=>"100001100",
  58957=>"101110111",
  58958=>"000010110",
  58959=>"001100011",
  58960=>"100011100",
  58961=>"011100000",
  58962=>"011000010",
  58963=>"100010111",
  58964=>"011110010",
  58965=>"101100110",
  58966=>"110000010",
  58967=>"100010010",
  58968=>"001110110",
  58969=>"101001110",
  58970=>"101110110",
  58971=>"000001001",
  58972=>"001010001",
  58973=>"011000010",
  58974=>"011110001",
  58975=>"100000000",
  58976=>"110011101",
  58977=>"011001011",
  58978=>"011111101",
  58979=>"111110000",
  58980=>"111110010",
  58981=>"010110111",
  58982=>"100101111",
  58983=>"001111000",
  58984=>"010111111",
  58985=>"111101011",
  58986=>"111111101",
  58987=>"001010000",
  58988=>"000000001",
  58989=>"000100100",
  58990=>"011101100",
  58991=>"000101111",
  58992=>"000001000",
  58993=>"010000000",
  58994=>"101101111",
  58995=>"010000111",
  58996=>"011011100",
  58997=>"100000001",
  58998=>"011100101",
  58999=>"110001111",
  59000=>"000101000",
  59001=>"110011100",
  59002=>"010100001",
  59003=>"100110111",
  59004=>"100100101",
  59005=>"100101101",
  59006=>"100011010",
  59007=>"111100010",
  59008=>"011111100",
  59009=>"000100110",
  59010=>"001100000",
  59011=>"011111010",
  59012=>"010001001",
  59013=>"100101101",
  59014=>"000100011",
  59015=>"111111111",
  59016=>"011001000",
  59017=>"011010000",
  59018=>"010111100",
  59019=>"010100101",
  59020=>"110010001",
  59021=>"000100000",
  59022=>"110110010",
  59023=>"101100000",
  59024=>"011011100",
  59025=>"011001101",
  59026=>"010011110",
  59027=>"010111001",
  59028=>"110011101",
  59029=>"100011110",
  59030=>"110111011",
  59031=>"011111110",
  59032=>"011001010",
  59033=>"000111111",
  59034=>"100001000",
  59035=>"101010001",
  59036=>"111111001",
  59037=>"100111100",
  59038=>"101011011",
  59039=>"110111011",
  59040=>"000101010",
  59041=>"000010100",
  59042=>"110001001",
  59043=>"001101000",
  59044=>"111010100",
  59045=>"010001110",
  59046=>"000001100",
  59047=>"001000000",
  59048=>"111110001",
  59049=>"111000000",
  59050=>"010001101",
  59051=>"010101011",
  59052=>"001110111",
  59053=>"101001011",
  59054=>"111000110",
  59055=>"000100000",
  59056=>"100000001",
  59057=>"110001111",
  59058=>"001101000",
  59059=>"001100110",
  59060=>"011110100",
  59061=>"111101000",
  59062=>"000111100",
  59063=>"011111011",
  59064=>"001001011",
  59065=>"101000001",
  59066=>"011001011",
  59067=>"010000111",
  59068=>"010000011",
  59069=>"100001100",
  59070=>"111011011",
  59071=>"111000010",
  59072=>"111101100",
  59073=>"101110110",
  59074=>"011001111",
  59075=>"101010110",
  59076=>"100001100",
  59077=>"111111110",
  59078=>"001000100",
  59079=>"101000101",
  59080=>"011010000",
  59081=>"101000011",
  59082=>"110001011",
  59083=>"000000100",
  59084=>"000000010",
  59085=>"110101111",
  59086=>"010001001",
  59087=>"000001010",
  59088=>"000110111",
  59089=>"001000101",
  59090=>"011101100",
  59091=>"100000100",
  59092=>"101001010",
  59093=>"001000011",
  59094=>"011011000",
  59095=>"110000001",
  59096=>"000000000",
  59097=>"101000111",
  59098=>"101001110",
  59099=>"111110000",
  59100=>"101111000",
  59101=>"100100101",
  59102=>"000011111",
  59103=>"010101011",
  59104=>"000010111",
  59105=>"111000000",
  59106=>"000111010",
  59107=>"010100000",
  59108=>"110100110",
  59109=>"001101111",
  59110=>"000000000",
  59111=>"001010111",
  59112=>"000110100",
  59113=>"100011110",
  59114=>"010111111",
  59115=>"111101100",
  59116=>"001110001",
  59117=>"000000101",
  59118=>"000000001",
  59119=>"110100110",
  59120=>"100001001",
  59121=>"010101000",
  59122=>"110100000",
  59123=>"010000111",
  59124=>"011001001",
  59125=>"110010010",
  59126=>"110110001",
  59127=>"111001101",
  59128=>"101001100",
  59129=>"111010100",
  59130=>"100000100",
  59131=>"000111100",
  59132=>"111110110",
  59133=>"000110000",
  59134=>"000101000",
  59135=>"001111010",
  59136=>"110111111",
  59137=>"000011001",
  59138=>"000100011",
  59139=>"011110101",
  59140=>"100001000",
  59141=>"001000001",
  59142=>"110010001",
  59143=>"010010011",
  59144=>"001110111",
  59145=>"110000111",
  59146=>"010000001",
  59147=>"001010011",
  59148=>"000010001",
  59149=>"001001111",
  59150=>"110101111",
  59151=>"111101101",
  59152=>"111100100",
  59153=>"010011011",
  59154=>"101001001",
  59155=>"001100110",
  59156=>"101011010",
  59157=>"000110101",
  59158=>"001110010",
  59159=>"100001111",
  59160=>"001101101",
  59161=>"010110000",
  59162=>"000110011",
  59163=>"000100100",
  59164=>"111010100",
  59165=>"011000101",
  59166=>"111011011",
  59167=>"100111000",
  59168=>"110110011",
  59169=>"101101001",
  59170=>"000001110",
  59171=>"011110000",
  59172=>"001100110",
  59173=>"011000111",
  59174=>"000110011",
  59175=>"101110110",
  59176=>"000110010",
  59177=>"111110110",
  59178=>"011110110",
  59179=>"101011000",
  59180=>"010111100",
  59181=>"000001111",
  59182=>"100111100",
  59183=>"000110100",
  59184=>"001101111",
  59185=>"111001001",
  59186=>"111000111",
  59187=>"110010111",
  59188=>"101111110",
  59189=>"110110101",
  59190=>"101110000",
  59191=>"111101111",
  59192=>"011010110",
  59193=>"001001011",
  59194=>"001001100",
  59195=>"110000010",
  59196=>"111100110",
  59197=>"111011001",
  59198=>"101001011",
  59199=>"011110001",
  59200=>"010001000",
  59201=>"100100100",
  59202=>"011000100",
  59203=>"011101110",
  59204=>"010010000",
  59205=>"011110111",
  59206=>"111011101",
  59207=>"110101000",
  59208=>"001010010",
  59209=>"000101100",
  59210=>"101111101",
  59211=>"100101111",
  59212=>"110100001",
  59213=>"101011100",
  59214=>"010000001",
  59215=>"110010111",
  59216=>"101101000",
  59217=>"100000000",
  59218=>"110101100",
  59219=>"111001100",
  59220=>"100000001",
  59221=>"110001010",
  59222=>"010110011",
  59223=>"011011111",
  59224=>"100111110",
  59225=>"101111000",
  59226=>"010110011",
  59227=>"111101111",
  59228=>"110100011",
  59229=>"001100110",
  59230=>"010110011",
  59231=>"000100111",
  59232=>"101101111",
  59233=>"111011011",
  59234=>"100000000",
  59235=>"100110111",
  59236=>"011010110",
  59237=>"100010001",
  59238=>"100011110",
  59239=>"101110011",
  59240=>"111001001",
  59241=>"000011000",
  59242=>"111010101",
  59243=>"011001100",
  59244=>"101110110",
  59245=>"100101101",
  59246=>"101100110",
  59247=>"100101100",
  59248=>"100110000",
  59249=>"000101100",
  59250=>"110110011",
  59251=>"001000101",
  59252=>"110000111",
  59253=>"001111010",
  59254=>"001000011",
  59255=>"001000000",
  59256=>"001111101",
  59257=>"010100100",
  59258=>"010100100",
  59259=>"011111010",
  59260=>"001010000",
  59261=>"001000011",
  59262=>"101000100",
  59263=>"100010110",
  59264=>"000010010",
  59265=>"100011010",
  59266=>"000101101",
  59267=>"001001111",
  59268=>"010111000",
  59269=>"101011111",
  59270=>"010100001",
  59271=>"000110010",
  59272=>"100101111",
  59273=>"000001001",
  59274=>"100110010",
  59275=>"010000100",
  59276=>"110000000",
  59277=>"001000100",
  59278=>"110100011",
  59279=>"011101101",
  59280=>"100110011",
  59281=>"000010010",
  59282=>"111100111",
  59283=>"011000110",
  59284=>"000011110",
  59285=>"111100100",
  59286=>"111010101",
  59287=>"001001110",
  59288=>"000110100",
  59289=>"000001001",
  59290=>"001010000",
  59291=>"010110111",
  59292=>"100000001",
  59293=>"110001111",
  59294=>"011110101",
  59295=>"111111111",
  59296=>"011100101",
  59297=>"111100011",
  59298=>"110011110",
  59299=>"001001000",
  59300=>"011001001",
  59301=>"111100111",
  59302=>"000111100",
  59303=>"000010001",
  59304=>"001110110",
  59305=>"101110000",
  59306=>"010011101",
  59307=>"101010111",
  59308=>"010111000",
  59309=>"111111100",
  59310=>"010101010",
  59311=>"111111010",
  59312=>"101011010",
  59313=>"100111000",
  59314=>"110011101",
  59315=>"010100010",
  59316=>"001100101",
  59317=>"100010001",
  59318=>"110010101",
  59319=>"010001010",
  59320=>"011001001",
  59321=>"001000010",
  59322=>"101000111",
  59323=>"110001001",
  59324=>"001010100",
  59325=>"001110101",
  59326=>"010001110",
  59327=>"000001001",
  59328=>"001110000",
  59329=>"111111111",
  59330=>"101110001",
  59331=>"100110001",
  59332=>"010010001",
  59333=>"000101110",
  59334=>"110011010",
  59335=>"100110110",
  59336=>"101100010",
  59337=>"101001101",
  59338=>"011101010",
  59339=>"100000001",
  59340=>"001000000",
  59341=>"011100101",
  59342=>"010011111",
  59343=>"110011001",
  59344=>"001101000",
  59345=>"010110000",
  59346=>"010110001",
  59347=>"100010001",
  59348=>"111111110",
  59349=>"010101110",
  59350=>"010100010",
  59351=>"101110110",
  59352=>"011011011",
  59353=>"110110101",
  59354=>"011100011",
  59355=>"110110100",
  59356=>"001000000",
  59357=>"001000101",
  59358=>"111101001",
  59359=>"011000110",
  59360=>"011001100",
  59361=>"010011100",
  59362=>"000110110",
  59363=>"110100000",
  59364=>"001011010",
  59365=>"111100111",
  59366=>"001000100",
  59367=>"010111010",
  59368=>"010100110",
  59369=>"110011101",
  59370=>"000101110",
  59371=>"000100000",
  59372=>"010010011",
  59373=>"110000100",
  59374=>"110000111",
  59375=>"110101000",
  59376=>"010000000",
  59377=>"111010000",
  59378=>"100111110",
  59379=>"011110111",
  59380=>"001111010",
  59381=>"011000111",
  59382=>"001111100",
  59383=>"001100111",
  59384=>"110001011",
  59385=>"001100001",
  59386=>"110110010",
  59387=>"110110011",
  59388=>"110000010",
  59389=>"110101111",
  59390=>"111000111",
  59391=>"010100001",
  59392=>"010000010",
  59393=>"010101010",
  59394=>"111111010",
  59395=>"001000001",
  59396=>"110111010",
  59397=>"000011001",
  59398=>"111010111",
  59399=>"101010011",
  59400=>"000000100",
  59401=>"101000000",
  59402=>"110011111",
  59403=>"010010100",
  59404=>"011000010",
  59405=>"111101000",
  59406=>"101111011",
  59407=>"001011001",
  59408=>"001100011",
  59409=>"011001000",
  59410=>"010111100",
  59411=>"100111011",
  59412=>"010100000",
  59413=>"110011011",
  59414=>"110001011",
  59415=>"010111001",
  59416=>"010010010",
  59417=>"101011011",
  59418=>"101011000",
  59419=>"011010111",
  59420=>"111101101",
  59421=>"001001110",
  59422=>"011101000",
  59423=>"101111011",
  59424=>"010101001",
  59425=>"010100111",
  59426=>"110111100",
  59427=>"110111110",
  59428=>"000000000",
  59429=>"111011100",
  59430=>"011000100",
  59431=>"111101111",
  59432=>"110101110",
  59433=>"001110011",
  59434=>"001101011",
  59435=>"100100101",
  59436=>"110000111",
  59437=>"101110000",
  59438=>"101100011",
  59439=>"111001101",
  59440=>"001011101",
  59441=>"111100100",
  59442=>"010000011",
  59443=>"000000110",
  59444=>"100000000",
  59445=>"111110100",
  59446=>"010001100",
  59447=>"111110000",
  59448=>"001100000",
  59449=>"101011111",
  59450=>"001001000",
  59451=>"000111011",
  59452=>"100001100",
  59453=>"101000010",
  59454=>"100001101",
  59455=>"110000100",
  59456=>"001010000",
  59457=>"011100011",
  59458=>"110001011",
  59459=>"101000000",
  59460=>"111010010",
  59461=>"010001010",
  59462=>"000100111",
  59463=>"000010011",
  59464=>"101010011",
  59465=>"001111101",
  59466=>"001101010",
  59467=>"000010101",
  59468=>"000111000",
  59469=>"000000101",
  59470=>"101111101",
  59471=>"001100000",
  59472=>"111111000",
  59473=>"010000100",
  59474=>"100100101",
  59475=>"001011011",
  59476=>"011001010",
  59477=>"001101101",
  59478=>"011010010",
  59479=>"111011010",
  59480=>"101000110",
  59481=>"000010010",
  59482=>"011010011",
  59483=>"110101011",
  59484=>"100010111",
  59485=>"101100011",
  59486=>"011011110",
  59487=>"100010010",
  59488=>"000100000",
  59489=>"100101111",
  59490=>"110011010",
  59491=>"000111111",
  59492=>"000000001",
  59493=>"100010010",
  59494=>"101110011",
  59495=>"111010100",
  59496=>"011001101",
  59497=>"111101000",
  59498=>"110101010",
  59499=>"111101110",
  59500=>"101001101",
  59501=>"000111110",
  59502=>"010000000",
  59503=>"111010110",
  59504=>"111111111",
  59505=>"111000001",
  59506=>"101001110",
  59507=>"000111000",
  59508=>"100110001",
  59509=>"011100100",
  59510=>"101010000",
  59511=>"001111111",
  59512=>"001010111",
  59513=>"011110010",
  59514=>"101011101",
  59515=>"100011111",
  59516=>"011111100",
  59517=>"010111110",
  59518=>"000011000",
  59519=>"000011101",
  59520=>"110111111",
  59521=>"010111011",
  59522=>"101000000",
  59523=>"100001111",
  59524=>"001001111",
  59525=>"011001011",
  59526=>"010110001",
  59527=>"111100010",
  59528=>"000111000",
  59529=>"101101000",
  59530=>"101001110",
  59531=>"010110110",
  59532=>"110111101",
  59533=>"110100110",
  59534=>"111111010",
  59535=>"111101010",
  59536=>"110101100",
  59537=>"101110110",
  59538=>"011100110",
  59539=>"100010001",
  59540=>"111001101",
  59541=>"100011110",
  59542=>"100010011",
  59543=>"111110101",
  59544=>"110010011",
  59545=>"010011010",
  59546=>"000100100",
  59547=>"010101111",
  59548=>"011010000",
  59549=>"101011111",
  59550=>"000000110",
  59551=>"011011001",
  59552=>"001001011",
  59553=>"101010100",
  59554=>"110010000",
  59555=>"100111001",
  59556=>"011111110",
  59557=>"111001010",
  59558=>"010010000",
  59559=>"011000101",
  59560=>"111010101",
  59561=>"111111011",
  59562=>"110111110",
  59563=>"110100110",
  59564=>"100111011",
  59565=>"111001001",
  59566=>"111010001",
  59567=>"110111100",
  59568=>"000101101",
  59569=>"000001101",
  59570=>"001100000",
  59571=>"101000000",
  59572=>"111101101",
  59573=>"110001001",
  59574=>"100001001",
  59575=>"001100000",
  59576=>"001001011",
  59577=>"011010000",
  59578=>"000111110",
  59579=>"000101101",
  59580=>"010110111",
  59581=>"101100001",
  59582=>"000101001",
  59583=>"010110001",
  59584=>"111010011",
  59585=>"111101000",
  59586=>"110110111",
  59587=>"010000111",
  59588=>"001111111",
  59589=>"001100011",
  59590=>"010010010",
  59591=>"010010100",
  59592=>"110101100",
  59593=>"100111111",
  59594=>"111001100",
  59595=>"111101001",
  59596=>"000000011",
  59597=>"011110100",
  59598=>"000001010",
  59599=>"100101101",
  59600=>"011111010",
  59601=>"110111101",
  59602=>"101001111",
  59603=>"000011001",
  59604=>"111100111",
  59605=>"010010100",
  59606=>"110001010",
  59607=>"011101000",
  59608=>"000011001",
  59609=>"111010010",
  59610=>"100000001",
  59611=>"111100111",
  59612=>"100110001",
  59613=>"100100001",
  59614=>"000101100",
  59615=>"101100111",
  59616=>"100000110",
  59617=>"001000011",
  59618=>"010110100",
  59619=>"001100110",
  59620=>"110011011",
  59621=>"001010001",
  59622=>"010101100",
  59623=>"001111000",
  59624=>"100100000",
  59625=>"111101001",
  59626=>"011001010",
  59627=>"100100011",
  59628=>"100011110",
  59629=>"010011100",
  59630=>"000000100",
  59631=>"000001101",
  59632=>"110110100",
  59633=>"110100111",
  59634=>"010101001",
  59635=>"110111001",
  59636=>"011001101",
  59637=>"111000110",
  59638=>"111100101",
  59639=>"000000110",
  59640=>"101110000",
  59641=>"100011110",
  59642=>"100101010",
  59643=>"001101001",
  59644=>"100000110",
  59645=>"111111100",
  59646=>"111100110",
  59647=>"100000111",
  59648=>"100011111",
  59649=>"010101011",
  59650=>"001111000",
  59651=>"011100010",
  59652=>"000100110",
  59653=>"111001110",
  59654=>"110100100",
  59655=>"101110000",
  59656=>"101110110",
  59657=>"000000100",
  59658=>"111010011",
  59659=>"000110000",
  59660=>"100101001",
  59661=>"001101000",
  59662=>"011100101",
  59663=>"100000010",
  59664=>"011001101",
  59665=>"110110100",
  59666=>"100111001",
  59667=>"011111011",
  59668=>"010000101",
  59669=>"110010010",
  59670=>"000010010",
  59671=>"110100010",
  59672=>"000010000",
  59673=>"101110000",
  59674=>"001111010",
  59675=>"011101001",
  59676=>"011100010",
  59677=>"100110100",
  59678=>"101111000",
  59679=>"001010100",
  59680=>"010000111",
  59681=>"110001010",
  59682=>"001001000",
  59683=>"001100010",
  59684=>"010001110",
  59685=>"111110100",
  59686=>"111111110",
  59687=>"110101010",
  59688=>"101100110",
  59689=>"111010111",
  59690=>"101111111",
  59691=>"010111011",
  59692=>"001100000",
  59693=>"011000101",
  59694=>"001100011",
  59695=>"000101101",
  59696=>"011111100",
  59697=>"000010111",
  59698=>"011001100",
  59699=>"000100111",
  59700=>"110100000",
  59701=>"001010011",
  59702=>"001011101",
  59703=>"011111010",
  59704=>"110100011",
  59705=>"001000111",
  59706=>"000011001",
  59707=>"111110001",
  59708=>"011101100",
  59709=>"111101010",
  59710=>"011001110",
  59711=>"010010110",
  59712=>"101101111",
  59713=>"000000000",
  59714=>"101110010",
  59715=>"001101011",
  59716=>"101100111",
  59717=>"110011001",
  59718=>"010111011",
  59719=>"111100110",
  59720=>"010110011",
  59721=>"111100010",
  59722=>"011111110",
  59723=>"110011011",
  59724=>"100010010",
  59725=>"100100101",
  59726=>"111110110",
  59727=>"101010001",
  59728=>"101011000",
  59729=>"001010110",
  59730=>"011100111",
  59731=>"001010011",
  59732=>"000000110",
  59733=>"011110001",
  59734=>"110100110",
  59735=>"110000101",
  59736=>"000011101",
  59737=>"010101100",
  59738=>"011001111",
  59739=>"100101111",
  59740=>"110010111",
  59741=>"001100011",
  59742=>"000000011",
  59743=>"100100111",
  59744=>"100111000",
  59745=>"110011101",
  59746=>"100101010",
  59747=>"010011100",
  59748=>"000100100",
  59749=>"010011111",
  59750=>"111100101",
  59751=>"010001101",
  59752=>"110000100",
  59753=>"001111001",
  59754=>"100100110",
  59755=>"000000111",
  59756=>"101000100",
  59757=>"000000011",
  59758=>"011100001",
  59759=>"110011011",
  59760=>"001111101",
  59761=>"001110101",
  59762=>"111001101",
  59763=>"000101111",
  59764=>"001010111",
  59765=>"010101100",
  59766=>"110000011",
  59767=>"010100000",
  59768=>"101100000",
  59769=>"101110010",
  59770=>"101000010",
  59771=>"101100110",
  59772=>"111010111",
  59773=>"101110110",
  59774=>"100011011",
  59775=>"100100100",
  59776=>"100110111",
  59777=>"100011001",
  59778=>"100011110",
  59779=>"011110010",
  59780=>"000000100",
  59781=>"000011001",
  59782=>"010001110",
  59783=>"010000010",
  59784=>"101101001",
  59785=>"001101011",
  59786=>"011111110",
  59787=>"101000010",
  59788=>"101101010",
  59789=>"000100110",
  59790=>"000001011",
  59791=>"010111111",
  59792=>"111011010",
  59793=>"011010001",
  59794=>"100011100",
  59795=>"000011101",
  59796=>"001100010",
  59797=>"100011000",
  59798=>"100100100",
  59799=>"100111010",
  59800=>"011010000",
  59801=>"000000111",
  59802=>"100110100",
  59803=>"100100101",
  59804=>"111100001",
  59805=>"111111101",
  59806=>"001011101",
  59807=>"100010010",
  59808=>"111011000",
  59809=>"000111011",
  59810=>"100110010",
  59811=>"111011001",
  59812=>"111110101",
  59813=>"010010000",
  59814=>"011111101",
  59815=>"000110111",
  59816=>"100111111",
  59817=>"000110101",
  59818=>"110000000",
  59819=>"011000001",
  59820=>"001101001",
  59821=>"010000000",
  59822=>"110100111",
  59823=>"100110001",
  59824=>"010011000",
  59825=>"011000111",
  59826=>"100101110",
  59827=>"001010010",
  59828=>"011000100",
  59829=>"000100010",
  59830=>"010001100",
  59831=>"001111011",
  59832=>"000111111",
  59833=>"001001101",
  59834=>"100011100",
  59835=>"110001101",
  59836=>"010110100",
  59837=>"011010011",
  59838=>"100100001",
  59839=>"110100100",
  59840=>"010101100",
  59841=>"000011110",
  59842=>"110010100",
  59843=>"001010000",
  59844=>"000000100",
  59845=>"101111000",
  59846=>"101001100",
  59847=>"010111000",
  59848=>"101101100",
  59849=>"101001100",
  59850=>"100000111",
  59851=>"111111110",
  59852=>"010001101",
  59853=>"100100001",
  59854=>"010000100",
  59855=>"111100000",
  59856=>"101100110",
  59857=>"000100011",
  59858=>"101101001",
  59859=>"000000111",
  59860=>"100011000",
  59861=>"001000110",
  59862=>"101110111",
  59863=>"010111111",
  59864=>"001010010",
  59865=>"000101000",
  59866=>"100001100",
  59867=>"100100100",
  59868=>"011010111",
  59869=>"001110100",
  59870=>"110000000",
  59871=>"111110100",
  59872=>"011101111",
  59873=>"101001101",
  59874=>"101101101",
  59875=>"101101101",
  59876=>"001100110",
  59877=>"100011011",
  59878=>"100000001",
  59879=>"001001100",
  59880=>"001011100",
  59881=>"000001111",
  59882=>"101000001",
  59883=>"100101111",
  59884=>"000001010",
  59885=>"001110000",
  59886=>"001001100",
  59887=>"111001100",
  59888=>"110110100",
  59889=>"101011110",
  59890=>"100011110",
  59891=>"101010011",
  59892=>"111000100",
  59893=>"111101100",
  59894=>"101110110",
  59895=>"101110011",
  59896=>"001110000",
  59897=>"001111111",
  59898=>"110000110",
  59899=>"001100111",
  59900=>"000110011",
  59901=>"111111111",
  59902=>"011110000",
  59903=>"000101110",
  59904=>"100101111",
  59905=>"011101111",
  59906=>"000001110",
  59907=>"010100100",
  59908=>"100101101",
  59909=>"110110100",
  59910=>"000101100",
  59911=>"011101011",
  59912=>"111011001",
  59913=>"100110100",
  59914=>"000100101",
  59915=>"101011110",
  59916=>"111001010",
  59917=>"111100001",
  59918=>"111111001",
  59919=>"100111100",
  59920=>"010101100",
  59921=>"100001111",
  59922=>"111001100",
  59923=>"101100101",
  59924=>"101010000",
  59925=>"001111000",
  59926=>"001111110",
  59927=>"011101001",
  59928=>"010110001",
  59929=>"000110010",
  59930=>"101000011",
  59931=>"000010000",
  59932=>"001001011",
  59933=>"101100100",
  59934=>"011011110",
  59935=>"101000111",
  59936=>"111011011",
  59937=>"100101001",
  59938=>"011001010",
  59939=>"001001110",
  59940=>"010000111",
  59941=>"111011000",
  59942=>"110011110",
  59943=>"101001000",
  59944=>"001110100",
  59945=>"101000001",
  59946=>"101010100",
  59947=>"100111111",
  59948=>"001011010",
  59949=>"000001001",
  59950=>"111111011",
  59951=>"000100000",
  59952=>"010011111",
  59953=>"101011010",
  59954=>"111011000",
  59955=>"110001111",
  59956=>"000100000",
  59957=>"011111101",
  59958=>"010001110",
  59959=>"101000000",
  59960=>"111110000",
  59961=>"010100011",
  59962=>"000001100",
  59963=>"100111111",
  59964=>"010000011",
  59965=>"100000001",
  59966=>"111110000",
  59967=>"011110000",
  59968=>"000000111",
  59969=>"001101110",
  59970=>"001000001",
  59971=>"101010111",
  59972=>"001111111",
  59973=>"011011010",
  59974=>"000000010",
  59975=>"110001110",
  59976=>"111011000",
  59977=>"010001010",
  59978=>"101111111",
  59979=>"111100110",
  59980=>"010100100",
  59981=>"011001001",
  59982=>"001100001",
  59983=>"110100011",
  59984=>"000011000",
  59985=>"010110001",
  59986=>"110111010",
  59987=>"111000100",
  59988=>"000101100",
  59989=>"111011000",
  59990=>"011000000",
  59991=>"110100110",
  59992=>"111001110",
  59993=>"010100011",
  59994=>"111001001",
  59995=>"001000001",
  59996=>"100010110",
  59997=>"111111110",
  59998=>"010010001",
  59999=>"101101101",
  60000=>"110010111",
  60001=>"000011101",
  60002=>"001101111",
  60003=>"101001011",
  60004=>"110011011",
  60005=>"001010110",
  60006=>"111000001",
  60007=>"111100010",
  60008=>"011100100",
  60009=>"000011011",
  60010=>"110110011",
  60011=>"010010010",
  60012=>"010010100",
  60013=>"010011101",
  60014=>"110101011",
  60015=>"111110110",
  60016=>"011000000",
  60017=>"001100011",
  60018=>"111111101",
  60019=>"101011111",
  60020=>"000010011",
  60021=>"111110101",
  60022=>"010110111",
  60023=>"101100000",
  60024=>"111011110",
  60025=>"010100001",
  60026=>"011010000",
  60027=>"111100110",
  60028=>"111101001",
  60029=>"001011011",
  60030=>"100111110",
  60031=>"101011100",
  60032=>"010111100",
  60033=>"000011010",
  60034=>"001100011",
  60035=>"000001101",
  60036=>"001010110",
  60037=>"111000110",
  60038=>"001100011",
  60039=>"101101110",
  60040=>"000100000",
  60041=>"000100101",
  60042=>"100000111",
  60043=>"011101110",
  60044=>"101011100",
  60045=>"101010100",
  60046=>"011001101",
  60047=>"100101100",
  60048=>"010111001",
  60049=>"001101001",
  60050=>"100100000",
  60051=>"010000011",
  60052=>"100010001",
  60053=>"111110100",
  60054=>"001010100",
  60055=>"100110100",
  60056=>"100000011",
  60057=>"001101010",
  60058=>"100101111",
  60059=>"001000101",
  60060=>"111010111",
  60061=>"111101001",
  60062=>"101011100",
  60063=>"011110101",
  60064=>"010110001",
  60065=>"101011101",
  60066=>"101100010",
  60067=>"010010111",
  60068=>"111010000",
  60069=>"011100001",
  60070=>"101010010",
  60071=>"101001110",
  60072=>"010110001",
  60073=>"101010100",
  60074=>"000011001",
  60075=>"110000000",
  60076=>"101010011",
  60077=>"110111101",
  60078=>"111101101",
  60079=>"110110000",
  60080=>"000011111",
  60081=>"000010001",
  60082=>"011011000",
  60083=>"000010010",
  60084=>"011100011",
  60085=>"101001010",
  60086=>"110011100",
  60087=>"010111111",
  60088=>"111100100",
  60089=>"010101010",
  60090=>"101000010",
  60091=>"011001101",
  60092=>"111001100",
  60093=>"001001000",
  60094=>"101110011",
  60095=>"011110001",
  60096=>"101001101",
  60097=>"110101101",
  60098=>"011110001",
  60099=>"111110111",
  60100=>"010001001",
  60101=>"100101010",
  60102=>"101000001",
  60103=>"111101111",
  60104=>"011010001",
  60105=>"010001101",
  60106=>"010110000",
  60107=>"001111100",
  60108=>"000001111",
  60109=>"010010010",
  60110=>"101101000",
  60111=>"110001000",
  60112=>"010000101",
  60113=>"011011100",
  60114=>"010111010",
  60115=>"001111011",
  60116=>"011110101",
  60117=>"010000111",
  60118=>"110001111",
  60119=>"010110011",
  60120=>"001011101",
  60121=>"100100000",
  60122=>"011111000",
  60123=>"010010000",
  60124=>"111110000",
  60125=>"010110110",
  60126=>"110101101",
  60127=>"001001001",
  60128=>"000111101",
  60129=>"010000110",
  60130=>"111010001",
  60131=>"001001000",
  60132=>"100110111",
  60133=>"010101010",
  60134=>"010111101",
  60135=>"011100011",
  60136=>"011010000",
  60137=>"001100000",
  60138=>"101111000",
  60139=>"001000111",
  60140=>"100000110",
  60141=>"000111110",
  60142=>"010001111",
  60143=>"001101000",
  60144=>"000111000",
  60145=>"111011011",
  60146=>"111111010",
  60147=>"110101000",
  60148=>"101001101",
  60149=>"111110110",
  60150=>"111101000",
  60151=>"110011111",
  60152=>"101011100",
  60153=>"001011100",
  60154=>"110101010",
  60155=>"101010001",
  60156=>"010010010",
  60157=>"011010111",
  60158=>"010110110",
  60159=>"100110100",
  60160=>"000000001",
  60161=>"100001001",
  60162=>"110011110",
  60163=>"011011000",
  60164=>"001011010",
  60165=>"000110000",
  60166=>"101001000",
  60167=>"001010111",
  60168=>"001011001",
  60169=>"110010110",
  60170=>"101001000",
  60171=>"000010110",
  60172=>"101101100",
  60173=>"000100101",
  60174=>"000101011",
  60175=>"111110101",
  60176=>"001100110",
  60177=>"001011010",
  60178=>"011100100",
  60179=>"001111110",
  60180=>"111000100",
  60181=>"111111010",
  60182=>"011110001",
  60183=>"011010000",
  60184=>"111100000",
  60185=>"011000001",
  60186=>"000101111",
  60187=>"101011100",
  60188=>"111100101",
  60189=>"000000001",
  60190=>"011111010",
  60191=>"000000110",
  60192=>"011010101",
  60193=>"100111011",
  60194=>"110001111",
  60195=>"010010010",
  60196=>"000101110",
  60197=>"101001001",
  60198=>"010000000",
  60199=>"011000111",
  60200=>"011111001",
  60201=>"001101011",
  60202=>"111110100",
  60203=>"010110001",
  60204=>"110110110",
  60205=>"110100111",
  60206=>"100001001",
  60207=>"010111101",
  60208=>"110001111",
  60209=>"001000101",
  60210=>"110100111",
  60211=>"101001001",
  60212=>"010001101",
  60213=>"010110000",
  60214=>"011110110",
  60215=>"001101000",
  60216=>"100100101",
  60217=>"001101111",
  60218=>"100000101",
  60219=>"110100010",
  60220=>"010111100",
  60221=>"111111010",
  60222=>"101010111",
  60223=>"110110111",
  60224=>"000110111",
  60225=>"100111101",
  60226=>"101010110",
  60227=>"111010110",
  60228=>"100100000",
  60229=>"110100010",
  60230=>"110101110",
  60231=>"110001001",
  60232=>"101100100",
  60233=>"001011111",
  60234=>"000001110",
  60235=>"011111100",
  60236=>"010011001",
  60237=>"110001100",
  60238=>"111011110",
  60239=>"101111010",
  60240=>"101011000",
  60241=>"001000000",
  60242=>"011100001",
  60243=>"101011100",
  60244=>"111110000",
  60245=>"101000110",
  60246=>"110010010",
  60247=>"111000001",
  60248=>"010111010",
  60249=>"011111100",
  60250=>"000101010",
  60251=>"010110101",
  60252=>"001010010",
  60253=>"000111100",
  60254=>"101111010",
  60255=>"100000000",
  60256=>"010011101",
  60257=>"100110010",
  60258=>"001000010",
  60259=>"110101110",
  60260=>"000001101",
  60261=>"011011111",
  60262=>"010100010",
  60263=>"010101011",
  60264=>"101100001",
  60265=>"001100001",
  60266=>"111001011",
  60267=>"111111110",
  60268=>"111110111",
  60269=>"001110100",
  60270=>"000101111",
  60271=>"000101101",
  60272=>"111011101",
  60273=>"011111011",
  60274=>"101111011",
  60275=>"101110000",
  60276=>"100010010",
  60277=>"100100100",
  60278=>"001001101",
  60279=>"000010100",
  60280=>"001100101",
  60281=>"111110001",
  60282=>"001011111",
  60283=>"110001001",
  60284=>"110000001",
  60285=>"111001111",
  60286=>"100110110",
  60287=>"001001010",
  60288=>"111101011",
  60289=>"001111111",
  60290=>"001000000",
  60291=>"011011000",
  60292=>"111111111",
  60293=>"010110001",
  60294=>"000100011",
  60295=>"000101001",
  60296=>"011111000",
  60297=>"111010100",
  60298=>"110111101",
  60299=>"111100000",
  60300=>"100010100",
  60301=>"010101001",
  60302=>"110111110",
  60303=>"100001010",
  60304=>"111010001",
  60305=>"111111101",
  60306=>"111101100",
  60307=>"110011010",
  60308=>"100111010",
  60309=>"100011010",
  60310=>"111000000",
  60311=>"010010100",
  60312=>"001111101",
  60313=>"000100000",
  60314=>"101000010",
  60315=>"010001011",
  60316=>"011101011",
  60317=>"011110011",
  60318=>"110100010",
  60319=>"110010100",
  60320=>"111101010",
  60321=>"100111000",
  60322=>"001100010",
  60323=>"000000011",
  60324=>"101111110",
  60325=>"111100101",
  60326=>"101000111",
  60327=>"110100000",
  60328=>"001000011",
  60329=>"111000000",
  60330=>"000111100",
  60331=>"100111101",
  60332=>"001000011",
  60333=>"000101111",
  60334=>"011110110",
  60335=>"001000101",
  60336=>"011111101",
  60337=>"010100000",
  60338=>"101011110",
  60339=>"111101100",
  60340=>"101000100",
  60341=>"111100101",
  60342=>"011011001",
  60343=>"011110011",
  60344=>"101101101",
  60345=>"111100110",
  60346=>"010000111",
  60347=>"010001000",
  60348=>"110010100",
  60349=>"010000000",
  60350=>"101011110",
  60351=>"110100101",
  60352=>"010001110",
  60353=>"110100011",
  60354=>"000010100",
  60355=>"010010000",
  60356=>"011001010",
  60357=>"001000000",
  60358=>"101110111",
  60359=>"011111001",
  60360=>"010010011",
  60361=>"000110001",
  60362=>"110111101",
  60363=>"011111010",
  60364=>"101001001",
  60365=>"110101101",
  60366=>"110001001",
  60367=>"100101000",
  60368=>"110110001",
  60369=>"101001110",
  60370=>"000111000",
  60371=>"011011000",
  60372=>"100100100",
  60373=>"101001101",
  60374=>"010111100",
  60375=>"000001101",
  60376=>"010000010",
  60377=>"101111000",
  60378=>"011110111",
  60379=>"110110100",
  60380=>"000101111",
  60381=>"110010101",
  60382=>"100001111",
  60383=>"110010000",
  60384=>"110100100",
  60385=>"100111101",
  60386=>"110100101",
  60387=>"101010000",
  60388=>"111101011",
  60389=>"101100011",
  60390=>"011011111",
  60391=>"101000111",
  60392=>"111011010",
  60393=>"000001110",
  60394=>"000100000",
  60395=>"100000011",
  60396=>"001111110",
  60397=>"001010000",
  60398=>"111000000",
  60399=>"110101011",
  60400=>"001001010",
  60401=>"101000011",
  60402=>"000111100",
  60403=>"011000111",
  60404=>"011110111",
  60405=>"110110100",
  60406=>"000110100",
  60407=>"011001100",
  60408=>"001000110",
  60409=>"001000111",
  60410=>"011110110",
  60411=>"111111011",
  60412=>"101100000",
  60413=>"000011101",
  60414=>"011001011",
  60415=>"100110000",
  60416=>"011000000",
  60417=>"101111001",
  60418=>"011000101",
  60419=>"101011001",
  60420=>"010100010",
  60421=>"001000110",
  60422=>"111110011",
  60423=>"010011000",
  60424=>"110011111",
  60425=>"101000001",
  60426=>"010100001",
  60427=>"110010111",
  60428=>"001111100",
  60429=>"001100000",
  60430=>"001000101",
  60431=>"110110010",
  60432=>"111111010",
  60433=>"001010110",
  60434=>"111011000",
  60435=>"110001011",
  60436=>"001001000",
  60437=>"001010000",
  60438=>"111010010",
  60439=>"000000111",
  60440=>"010110100",
  60441=>"101011110",
  60442=>"001111000",
  60443=>"100011001",
  60444=>"111110001",
  60445=>"101100101",
  60446=>"100110001",
  60447=>"110110110",
  60448=>"110010101",
  60449=>"001010010",
  60450=>"000000000",
  60451=>"010001111",
  60452=>"101000001",
  60453=>"110101000",
  60454=>"101000010",
  60455=>"101010001",
  60456=>"010101010",
  60457=>"100010100",
  60458=>"010101011",
  60459=>"001100101",
  60460=>"111111010",
  60461=>"110110010",
  60462=>"011100011",
  60463=>"111110001",
  60464=>"110001110",
  60465=>"000110100",
  60466=>"101001010",
  60467=>"110011010",
  60468=>"110111010",
  60469=>"000011000",
  60470=>"100010101",
  60471=>"101111111",
  60472=>"001110111",
  60473=>"111110010",
  60474=>"000111101",
  60475=>"001000011",
  60476=>"100001001",
  60477=>"001100001",
  60478=>"111011101",
  60479=>"111000010",
  60480=>"010000100",
  60481=>"100111001",
  60482=>"100101000",
  60483=>"011101000",
  60484=>"010010000",
  60485=>"011101110",
  60486=>"100010100",
  60487=>"011111100",
  60488=>"001000100",
  60489=>"001110011",
  60490=>"010101101",
  60491=>"100100111",
  60492=>"101010101",
  60493=>"100110111",
  60494=>"110100100",
  60495=>"111110010",
  60496=>"111110101",
  60497=>"011010000",
  60498=>"011110110",
  60499=>"101011100",
  60500=>"101111010",
  60501=>"110000100",
  60502=>"011011001",
  60503=>"110011110",
  60504=>"101111110",
  60505=>"100000111",
  60506=>"101001001",
  60507=>"010000011",
  60508=>"101001001",
  60509=>"100011111",
  60510=>"001011010",
  60511=>"100001101",
  60512=>"100010011",
  60513=>"110000000",
  60514=>"100010000",
  60515=>"100101100",
  60516=>"100111101",
  60517=>"111110110",
  60518=>"100001001",
  60519=>"110010000",
  60520=>"001110100",
  60521=>"110110011",
  60522=>"101001000",
  60523=>"111101011",
  60524=>"001001101",
  60525=>"001101111",
  60526=>"000010010",
  60527=>"000101111",
  60528=>"110010010",
  60529=>"000000000",
  60530=>"111110101",
  60531=>"110000001",
  60532=>"100111111",
  60533=>"110101110",
  60534=>"000110000",
  60535=>"001101010",
  60536=>"101110110",
  60537=>"011010110",
  60538=>"110001110",
  60539=>"101111101",
  60540=>"111101100",
  60541=>"111111001",
  60542=>"100101000",
  60543=>"111101100",
  60544=>"110110011",
  60545=>"011111111",
  60546=>"010001110",
  60547=>"100100000",
  60548=>"110000110",
  60549=>"001011100",
  60550=>"000110010",
  60551=>"100010000",
  60552=>"001000010",
  60553=>"100110100",
  60554=>"000101100",
  60555=>"111101100",
  60556=>"000110011",
  60557=>"110101111",
  60558=>"110001001",
  60559=>"000010000",
  60560=>"110110100",
  60561=>"010001000",
  60562=>"000001010",
  60563=>"001100111",
  60564=>"011101001",
  60565=>"111011110",
  60566=>"010101011",
  60567=>"011001101",
  60568=>"111100101",
  60569=>"111011000",
  60570=>"001110111",
  60571=>"011011100",
  60572=>"100011001",
  60573=>"110101000",
  60574=>"111000000",
  60575=>"001011001",
  60576=>"000100101",
  60577=>"110110111",
  60578=>"011101100",
  60579=>"000000001",
  60580=>"101111011",
  60581=>"011110011",
  60582=>"001010001",
  60583=>"111001000",
  60584=>"111010100",
  60585=>"111001100",
  60586=>"001110001",
  60587=>"000011000",
  60588=>"101010011",
  60589=>"011110000",
  60590=>"110101101",
  60591=>"111101110",
  60592=>"011001010",
  60593=>"101110001",
  60594=>"101010110",
  60595=>"010110100",
  60596=>"011100001",
  60597=>"101001001",
  60598=>"101010001",
  60599=>"010000011",
  60600=>"101010100",
  60601=>"111001000",
  60602=>"000010000",
  60603=>"110010000",
  60604=>"001010000",
  60605=>"100110011",
  60606=>"101000100",
  60607=>"111011101",
  60608=>"000101000",
  60609=>"010011011",
  60610=>"010101000",
  60611=>"111111111",
  60612=>"011001111",
  60613=>"111111110",
  60614=>"001010110",
  60615=>"101101110",
  60616=>"000101011",
  60617=>"000000001",
  60618=>"111100101",
  60619=>"110110011",
  60620=>"100010100",
  60621=>"000000101",
  60622=>"011101010",
  60623=>"010010100",
  60624=>"100111110",
  60625=>"010110110",
  60626=>"010100110",
  60627=>"011001101",
  60628=>"110110011",
  60629=>"001100011",
  60630=>"110110000",
  60631=>"001100010",
  60632=>"001100010",
  60633=>"010001111",
  60634=>"100000100",
  60635=>"000000001",
  60636=>"110100000",
  60637=>"010110001",
  60638=>"011110011",
  60639=>"101110010",
  60640=>"101101000",
  60641=>"111010001",
  60642=>"111111011",
  60643=>"000100101",
  60644=>"001110011",
  60645=>"001000001",
  60646=>"111101000",
  60647=>"010001110",
  60648=>"010100010",
  60649=>"111110001",
  60650=>"010010010",
  60651=>"000011100",
  60652=>"010011100",
  60653=>"011010011",
  60654=>"001100110",
  60655=>"101000000",
  60656=>"101000111",
  60657=>"111110101",
  60658=>"111011001",
  60659=>"111100010",
  60660=>"110111000",
  60661=>"010010101",
  60662=>"001010011",
  60663=>"000001110",
  60664=>"101111101",
  60665=>"111111101",
  60666=>"101001000",
  60667=>"010000001",
  60668=>"011000100",
  60669=>"110110101",
  60670=>"100000001",
  60671=>"111110110",
  60672=>"010000010",
  60673=>"010111010",
  60674=>"110011011",
  60675=>"111110110",
  60676=>"000101000",
  60677=>"110100011",
  60678=>"101110010",
  60679=>"000100101",
  60680=>"101001000",
  60681=>"100000110",
  60682=>"111010011",
  60683=>"101000010",
  60684=>"100100011",
  60685=>"000100000",
  60686=>"001010110",
  60687=>"011011110",
  60688=>"001110000",
  60689=>"000010010",
  60690=>"010010010",
  60691=>"011000001",
  60692=>"000011000",
  60693=>"101101010",
  60694=>"010011100",
  60695=>"001101010",
  60696=>"101101110",
  60697=>"000010100",
  60698=>"000001110",
  60699=>"110011100",
  60700=>"111100111",
  60701=>"110100000",
  60702=>"001011100",
  60703=>"001111011",
  60704=>"011011011",
  60705=>"010010000",
  60706=>"010110000",
  60707=>"111011000",
  60708=>"011101001",
  60709=>"010101101",
  60710=>"000001101",
  60711=>"010111111",
  60712=>"110000111",
  60713=>"110111100",
  60714=>"101111110",
  60715=>"011101010",
  60716=>"011101001",
  60717=>"101110000",
  60718=>"001111111",
  60719=>"111100100",
  60720=>"011101111",
  60721=>"011000000",
  60722=>"001011000",
  60723=>"010000100",
  60724=>"100001010",
  60725=>"010111110",
  60726=>"011101101",
  60727=>"100010001",
  60728=>"000011000",
  60729=>"110000010",
  60730=>"101100100",
  60731=>"000111110",
  60732=>"100000110",
  60733=>"110000001",
  60734=>"011010000",
  60735=>"001010101",
  60736=>"100101110",
  60737=>"011110110",
  60738=>"001111011",
  60739=>"011100101",
  60740=>"100001101",
  60741=>"110001110",
  60742=>"110011000",
  60743=>"000000001",
  60744=>"011011111",
  60745=>"111000110",
  60746=>"111100111",
  60747=>"111011001",
  60748=>"000000110",
  60749=>"001011010",
  60750=>"001100000",
  60751=>"010001101",
  60752=>"101001100",
  60753=>"111111001",
  60754=>"100100011",
  60755=>"111101000",
  60756=>"100010110",
  60757=>"001001101",
  60758=>"011111101",
  60759=>"010000000",
  60760=>"010111001",
  60761=>"100101000",
  60762=>"100100010",
  60763=>"010100000",
  60764=>"111111100",
  60765=>"101100100",
  60766=>"100001001",
  60767=>"111000001",
  60768=>"110000101",
  60769=>"001110101",
  60770=>"010001111",
  60771=>"001101100",
  60772=>"001000111",
  60773=>"000111110",
  60774=>"011011010",
  60775=>"010110111",
  60776=>"110111110",
  60777=>"000110100",
  60778=>"111111000",
  60779=>"110100000",
  60780=>"101010011",
  60781=>"011010011",
  60782=>"000100000",
  60783=>"011100001",
  60784=>"010001001",
  60785=>"101101111",
  60786=>"101110101",
  60787=>"110011101",
  60788=>"110101011",
  60789=>"111111101",
  60790=>"011111001",
  60791=>"011010010",
  60792=>"010101010",
  60793=>"011111110",
  60794=>"000100101",
  60795=>"110010111",
  60796=>"011000000",
  60797=>"110000011",
  60798=>"000001101",
  60799=>"110111000",
  60800=>"100101111",
  60801=>"011100110",
  60802=>"101001011",
  60803=>"001010111",
  60804=>"000011010",
  60805=>"011001110",
  60806=>"100100010",
  60807=>"000010001",
  60808=>"001010101",
  60809=>"100100110",
  60810=>"001010010",
  60811=>"000001100",
  60812=>"101101001",
  60813=>"111101110",
  60814=>"000000010",
  60815=>"010111001",
  60816=>"001101101",
  60817=>"011100110",
  60818=>"110001110",
  60819=>"000000100",
  60820=>"011000101",
  60821=>"001111100",
  60822=>"011000000",
  60823=>"000101010",
  60824=>"010011101",
  60825=>"110100111",
  60826=>"110100011",
  60827=>"011000100",
  60828=>"100000010",
  60829=>"011001001",
  60830=>"100100010",
  60831=>"001100000",
  60832=>"010111110",
  60833=>"011111010",
  60834=>"011100001",
  60835=>"000100100",
  60836=>"100111001",
  60837=>"010011000",
  60838=>"110001010",
  60839=>"100001100",
  60840=>"011101010",
  60841=>"011111111",
  60842=>"001100001",
  60843=>"000110010",
  60844=>"111111000",
  60845=>"000100001",
  60846=>"100101010",
  60847=>"001111000",
  60848=>"001000000",
  60849=>"110111010",
  60850=>"100010001",
  60851=>"110000001",
  60852=>"011110101",
  60853=>"101100100",
  60854=>"110111011",
  60855=>"010001110",
  60856=>"101001010",
  60857=>"101000111",
  60858=>"011100110",
  60859=>"100001111",
  60860=>"101100100",
  60861=>"000000101",
  60862=>"101111110",
  60863=>"111000000",
  60864=>"111111000",
  60865=>"010011101",
  60866=>"110100010",
  60867=>"010100010",
  60868=>"000001110",
  60869=>"010110011",
  60870=>"010100110",
  60871=>"100000001",
  60872=>"110001101",
  60873=>"100010001",
  60874=>"001101101",
  60875=>"011101011",
  60876=>"000010000",
  60877=>"111000001",
  60878=>"111100001",
  60879=>"100100110",
  60880=>"100110111",
  60881=>"000100111",
  60882=>"001111010",
  60883=>"001010110",
  60884=>"100011100",
  60885=>"100001100",
  60886=>"110000010",
  60887=>"001001111",
  60888=>"101000000",
  60889=>"010101101",
  60890=>"010011100",
  60891=>"111010010",
  60892=>"001000001",
  60893=>"110100101",
  60894=>"101111110",
  60895=>"101111100",
  60896=>"010010100",
  60897=>"101011010",
  60898=>"100101001",
  60899=>"010000111",
  60900=>"111101000",
  60901=>"100000000",
  60902=>"010100011",
  60903=>"001000011",
  60904=>"001111101",
  60905=>"010110010",
  60906=>"000011011",
  60907=>"111001000",
  60908=>"010100111",
  60909=>"010000100",
  60910=>"001010111",
  60911=>"011101011",
  60912=>"111110100",
  60913=>"001010001",
  60914=>"011001100",
  60915=>"110101011",
  60916=>"000110000",
  60917=>"011000101",
  60918=>"101100010",
  60919=>"000100100",
  60920=>"000010110",
  60921=>"011010100",
  60922=>"010110000",
  60923=>"101001111",
  60924=>"111010001",
  60925=>"000001100",
  60926=>"111110111",
  60927=>"101000100",
  60928=>"010100111",
  60929=>"110001010",
  60930=>"011011001",
  60931=>"111111011",
  60932=>"010001110",
  60933=>"000010011",
  60934=>"101001001",
  60935=>"000011110",
  60936=>"100010000",
  60937=>"010111111",
  60938=>"001000010",
  60939=>"010010110",
  60940=>"110000011",
  60941=>"111000001",
  60942=>"101110110",
  60943=>"111111011",
  60944=>"011010000",
  60945=>"011110011",
  60946=>"110100111",
  60947=>"110000111",
  60948=>"010010011",
  60949=>"001110010",
  60950=>"111101110",
  60951=>"001110000",
  60952=>"000100010",
  60953=>"001111001",
  60954=>"010001110",
  60955=>"000000111",
  60956=>"101111100",
  60957=>"001111011",
  60958=>"111001111",
  60959=>"001111001",
  60960=>"001101001",
  60961=>"100100010",
  60962=>"101101000",
  60963=>"100000110",
  60964=>"000110001",
  60965=>"010011011",
  60966=>"100000011",
  60967=>"001101111",
  60968=>"111000100",
  60969=>"001001010",
  60970=>"101110111",
  60971=>"100010100",
  60972=>"011000100",
  60973=>"010110111",
  60974=>"000001001",
  60975=>"111111101",
  60976=>"110100010",
  60977=>"001010100",
  60978=>"000100101",
  60979=>"001001111",
  60980=>"101100000",
  60981=>"100111111",
  60982=>"101111011",
  60983=>"011001101",
  60984=>"010010001",
  60985=>"010000010",
  60986=>"101000101",
  60987=>"000000111",
  60988=>"100101001",
  60989=>"100100101",
  60990=>"000101010",
  60991=>"001101110",
  60992=>"101011000",
  60993=>"110111010",
  60994=>"110011111",
  60995=>"001101011",
  60996=>"001011111",
  60997=>"011011011",
  60998=>"100100010",
  60999=>"011100100",
  61000=>"101010001",
  61001=>"100011111",
  61002=>"111011111",
  61003=>"100011100",
  61004=>"000001000",
  61005=>"101001011",
  61006=>"100010110",
  61007=>"010010101",
  61008=>"010100011",
  61009=>"111001011",
  61010=>"101111011",
  61011=>"000000000",
  61012=>"111010001",
  61013=>"010010100",
  61014=>"010001001",
  61015=>"110010111",
  61016=>"010111011",
  61017=>"110101000",
  61018=>"110110111",
  61019=>"010010010",
  61020=>"000100111",
  61021=>"111101001",
  61022=>"101100000",
  61023=>"111010011",
  61024=>"110001000",
  61025=>"101101101",
  61026=>"100110110",
  61027=>"001110111",
  61028=>"111010101",
  61029=>"101000100",
  61030=>"010110000",
  61031=>"101101001",
  61032=>"100100011",
  61033=>"000111100",
  61034=>"101100110",
  61035=>"101011001",
  61036=>"111101110",
  61037=>"000101000",
  61038=>"010110110",
  61039=>"101011100",
  61040=>"001000101",
  61041=>"000001010",
  61042=>"001100101",
  61043=>"100100111",
  61044=>"111010110",
  61045=>"111100100",
  61046=>"111001000",
  61047=>"111010101",
  61048=>"101010100",
  61049=>"001101011",
  61050=>"000110001",
  61051=>"010011100",
  61052=>"101000110",
  61053=>"011001011",
  61054=>"011001101",
  61055=>"011111011",
  61056=>"101100000",
  61057=>"010001110",
  61058=>"001010001",
  61059=>"110111001",
  61060=>"110110010",
  61061=>"010011111",
  61062=>"011001100",
  61063=>"100011010",
  61064=>"010111100",
  61065=>"011000001",
  61066=>"110010010",
  61067=>"101001101",
  61068=>"100010110",
  61069=>"000000001",
  61070=>"101101110",
  61071=>"001001100",
  61072=>"100110010",
  61073=>"001011010",
  61074=>"001110001",
  61075=>"100110111",
  61076=>"011010111",
  61077=>"100101111",
  61078=>"000110011",
  61079=>"000010001",
  61080=>"000011001",
  61081=>"001101001",
  61082=>"000011111",
  61083=>"001110011",
  61084=>"110101001",
  61085=>"100011110",
  61086=>"110000101",
  61087=>"100100010",
  61088=>"100111101",
  61089=>"001111100",
  61090=>"000111111",
  61091=>"110011100",
  61092=>"000011101",
  61093=>"101101001",
  61094=>"001101000",
  61095=>"010101001",
  61096=>"011011000",
  61097=>"110100010",
  61098=>"011001100",
  61099=>"111111110",
  61100=>"011111111",
  61101=>"001100011",
  61102=>"111010100",
  61103=>"001101110",
  61104=>"001010101",
  61105=>"000111111",
  61106=>"111001110",
  61107=>"101100111",
  61108=>"101000001",
  61109=>"111000000",
  61110=>"010010011",
  61111=>"111111100",
  61112=>"010001010",
  61113=>"001100010",
  61114=>"110011101",
  61115=>"101010101",
  61116=>"001111111",
  61117=>"111011000",
  61118=>"000111110",
  61119=>"100111000",
  61120=>"001010100",
  61121=>"011011010",
  61122=>"100001000",
  61123=>"010001000",
  61124=>"101010111",
  61125=>"000001000",
  61126=>"011000111",
  61127=>"101011010",
  61128=>"110101100",
  61129=>"110111011",
  61130=>"110110111",
  61131=>"111010101",
  61132=>"111100011",
  61133=>"011110111",
  61134=>"101111000",
  61135=>"101010010",
  61136=>"010010011",
  61137=>"000110100",
  61138=>"011011100",
  61139=>"100000001",
  61140=>"000101110",
  61141=>"011010101",
  61142=>"011011010",
  61143=>"101001101",
  61144=>"001000011",
  61145=>"010001101",
  61146=>"101011001",
  61147=>"110100001",
  61148=>"100011010",
  61149=>"000011110",
  61150=>"011011000",
  61151=>"110000011",
  61152=>"000000000",
  61153=>"000110100",
  61154=>"111100011",
  61155=>"000010100",
  61156=>"111010111",
  61157=>"001110110",
  61158=>"011100101",
  61159=>"010011111",
  61160=>"110101100",
  61161=>"001101011",
  61162=>"111011010",
  61163=>"010110000",
  61164=>"000001011",
  61165=>"001110101",
  61166=>"011110111",
  61167=>"110101001",
  61168=>"110111111",
  61169=>"100111000",
  61170=>"110110100",
  61171=>"110010111",
  61172=>"101010101",
  61173=>"111101011",
  61174=>"010100011",
  61175=>"000000111",
  61176=>"110110110",
  61177=>"000010000",
  61178=>"110011001",
  61179=>"000000010",
  61180=>"101010011",
  61181=>"000111111",
  61182=>"011101100",
  61183=>"011000001",
  61184=>"111010111",
  61185=>"110100100",
  61186=>"000011000",
  61187=>"010010000",
  61188=>"011111001",
  61189=>"011010100",
  61190=>"111111000",
  61191=>"000100101",
  61192=>"000110111",
  61193=>"111000110",
  61194=>"000010111",
  61195=>"111100111",
  61196=>"011110111",
  61197=>"100111010",
  61198=>"001000011",
  61199=>"111110111",
  61200=>"100001100",
  61201=>"110011101",
  61202=>"100011000",
  61203=>"110011000",
  61204=>"100011001",
  61205=>"011100010",
  61206=>"100010100",
  61207=>"011001101",
  61208=>"011101010",
  61209=>"001010001",
  61210=>"111011001",
  61211=>"111100010",
  61212=>"000100110",
  61213=>"100111111",
  61214=>"000000000",
  61215=>"110001111",
  61216=>"111111100",
  61217=>"110101101",
  61218=>"000010100",
  61219=>"000101011",
  61220=>"111001001",
  61221=>"100000000",
  61222=>"100001001",
  61223=>"010110000",
  61224=>"000000011",
  61225=>"110100001",
  61226=>"100111001",
  61227=>"010001000",
  61228=>"000011011",
  61229=>"000000000",
  61230=>"001111011",
  61231=>"010000000",
  61232=>"011100111",
  61233=>"111100011",
  61234=>"000011100",
  61235=>"111110100",
  61236=>"100111000",
  61237=>"111000101",
  61238=>"100100011",
  61239=>"000100111",
  61240=>"101111111",
  61241=>"111000110",
  61242=>"000100111",
  61243=>"011101111",
  61244=>"001110101",
  61245=>"001101000",
  61246=>"100000111",
  61247=>"000000010",
  61248=>"101111010",
  61249=>"110110100",
  61250=>"000101011",
  61251=>"101010111",
  61252=>"101011000",
  61253=>"100011100",
  61254=>"000000110",
  61255=>"011111111",
  61256=>"001010110",
  61257=>"001000100",
  61258=>"101000100",
  61259=>"100000011",
  61260=>"011100110",
  61261=>"001000001",
  61262=>"100010001",
  61263=>"001110110",
  61264=>"100010000",
  61265=>"001001000",
  61266=>"000101011",
  61267=>"101011010",
  61268=>"101101111",
  61269=>"001100000",
  61270=>"001000100",
  61271=>"010100000",
  61272=>"110100101",
  61273=>"111010110",
  61274=>"011010000",
  61275=>"010100100",
  61276=>"010101001",
  61277=>"101100111",
  61278=>"011110111",
  61279=>"001010011",
  61280=>"001111110",
  61281=>"111011101",
  61282=>"110111011",
  61283=>"101001001",
  61284=>"011000010",
  61285=>"110001101",
  61286=>"100001010",
  61287=>"001101000",
  61288=>"110101110",
  61289=>"100111001",
  61290=>"001001001",
  61291=>"010011110",
  61292=>"001000110",
  61293=>"001001010",
  61294=>"011000001",
  61295=>"010011100",
  61296=>"110010110",
  61297=>"111100101",
  61298=>"010011011",
  61299=>"001011000",
  61300=>"111101101",
  61301=>"010111111",
  61302=>"100010000",
  61303=>"100001011",
  61304=>"000001001",
  61305=>"111100111",
  61306=>"111110010",
  61307=>"110110111",
  61308=>"101101011",
  61309=>"100000011",
  61310=>"001111110",
  61311=>"010111101",
  61312=>"010011111",
  61313=>"101111001",
  61314=>"110101000",
  61315=>"111100101",
  61316=>"101011100",
  61317=>"110010000",
  61318=>"001000110",
  61319=>"010001010",
  61320=>"100011001",
  61321=>"111000111",
  61322=>"110111000",
  61323=>"101100100",
  61324=>"010101110",
  61325=>"001110110",
  61326=>"110011101",
  61327=>"101111000",
  61328=>"101101100",
  61329=>"001011110",
  61330=>"000000111",
  61331=>"010011010",
  61332=>"000100110",
  61333=>"010111001",
  61334=>"011001010",
  61335=>"011000111",
  61336=>"000011110",
  61337=>"011101101",
  61338=>"011101101",
  61339=>"000001010",
  61340=>"001110001",
  61341=>"000001100",
  61342=>"010101001",
  61343=>"110100011",
  61344=>"000000011",
  61345=>"000001101",
  61346=>"001101011",
  61347=>"101110100",
  61348=>"001000010",
  61349=>"011110010",
  61350=>"110100100",
  61351=>"100000000",
  61352=>"001100010",
  61353=>"010110110",
  61354=>"010010011",
  61355=>"101010111",
  61356=>"000000010",
  61357=>"110101100",
  61358=>"010010010",
  61359=>"011100010",
  61360=>"010100100",
  61361=>"111110100",
  61362=>"001010011",
  61363=>"000100101",
  61364=>"000001100",
  61365=>"001010001",
  61366=>"111011010",
  61367=>"111011110",
  61368=>"111001111",
  61369=>"011101100",
  61370=>"110101100",
  61371=>"010110010",
  61372=>"010110110",
  61373=>"001101101",
  61374=>"110000011",
  61375=>"101001101",
  61376=>"011100000",
  61377=>"001110110",
  61378=>"100100111",
  61379=>"111001100",
  61380=>"100000010",
  61381=>"110010001",
  61382=>"110000010",
  61383=>"101101000",
  61384=>"111101111",
  61385=>"100110101",
  61386=>"010100000",
  61387=>"111101111",
  61388=>"000000110",
  61389=>"010000110",
  61390=>"001110011",
  61391=>"110111010",
  61392=>"111001111",
  61393=>"000001110",
  61394=>"000011110",
  61395=>"110111011",
  61396=>"001100001",
  61397=>"000101110",
  61398=>"001111000",
  61399=>"110111001",
  61400=>"110100010",
  61401=>"111100110",
  61402=>"110010010",
  61403=>"001101011",
  61404=>"011100101",
  61405=>"100110010",
  61406=>"101001101",
  61407=>"001011000",
  61408=>"011111111",
  61409=>"011001000",
  61410=>"101110101",
  61411=>"001110000",
  61412=>"001110010",
  61413=>"011010000",
  61414=>"000111111",
  61415=>"110010000",
  61416=>"011011100",
  61417=>"111110001",
  61418=>"010110011",
  61419=>"001110010",
  61420=>"110011010",
  61421=>"000011111",
  61422=>"000000110",
  61423=>"100100001",
  61424=>"101010011",
  61425=>"000111111",
  61426=>"010110100",
  61427=>"111101100",
  61428=>"110010011",
  61429=>"111011101",
  61430=>"100111001",
  61431=>"000111111",
  61432=>"010011011",
  61433=>"110100100",
  61434=>"110111100",
  61435=>"100110101",
  61436=>"111000100",
  61437=>"101010110",
  61438=>"000000110",
  61439=>"101100011",
  61440=>"001001001",
  61441=>"100101111",
  61442=>"111011100",
  61443=>"101110011",
  61444=>"000010011",
  61445=>"000110001",
  61446=>"011011001",
  61447=>"011101101",
  61448=>"011101111",
  61449=>"000100110",
  61450=>"010000110",
  61451=>"111101011",
  61452=>"101001100",
  61453=>"010000100",
  61454=>"000010000",
  61455=>"101010101",
  61456=>"100011011",
  61457=>"010010000",
  61458=>"010101000",
  61459=>"001111110",
  61460=>"010000000",
  61461=>"011100010",
  61462=>"111001100",
  61463=>"110011100",
  61464=>"100110111",
  61465=>"010110111",
  61466=>"010010110",
  61467=>"100101011",
  61468=>"111000010",
  61469=>"100001011",
  61470=>"110101001",
  61471=>"001110000",
  61472=>"100000001",
  61473=>"011110001",
  61474=>"001110110",
  61475=>"000001000",
  61476=>"101011010",
  61477=>"110010010",
  61478=>"111110111",
  61479=>"111001110",
  61480=>"010000110",
  61481=>"101111011",
  61482=>"100001001",
  61483=>"110101000",
  61484=>"100111100",
  61485=>"000001111",
  61486=>"000111111",
  61487=>"100010111",
  61488=>"000001110",
  61489=>"111111111",
  61490=>"111011010",
  61491=>"001000100",
  61492=>"000010010",
  61493=>"101000100",
  61494=>"010000011",
  61495=>"000110011",
  61496=>"001000011",
  61497=>"000001010",
  61498=>"111001011",
  61499=>"010101111",
  61500=>"111010001",
  61501=>"100000110",
  61502=>"100011001",
  61503=>"000100100",
  61504=>"100000101",
  61505=>"110000011",
  61506=>"001001111",
  61507=>"010001101",
  61508=>"110110001",
  61509=>"001111110",
  61510=>"011010011",
  61511=>"110111101",
  61512=>"011110010",
  61513=>"000011000",
  61514=>"110010111",
  61515=>"100101101",
  61516=>"110100011",
  61517=>"100000111",
  61518=>"100011100",
  61519=>"111110111",
  61520=>"000001001",
  61521=>"010011100",
  61522=>"001111110",
  61523=>"000111110",
  61524=>"101011110",
  61525=>"110010110",
  61526=>"101001000",
  61527=>"111000100",
  61528=>"011000000",
  61529=>"001111100",
  61530=>"100110100",
  61531=>"100000001",
  61532=>"111101011",
  61533=>"000101111",
  61534=>"010010001",
  61535=>"111001111",
  61536=>"100110100",
  61537=>"101000110",
  61538=>"000111101",
  61539=>"001101011",
  61540=>"110000101",
  61541=>"000001101",
  61542=>"111001101",
  61543=>"101111101",
  61544=>"100111110",
  61545=>"100011111",
  61546=>"110010000",
  61547=>"110111010",
  61548=>"011000001",
  61549=>"111101011",
  61550=>"001000100",
  61551=>"000100000",
  61552=>"010011110",
  61553=>"110111111",
  61554=>"001010100",
  61555=>"100110110",
  61556=>"111010100",
  61557=>"000000100",
  61558=>"001110111",
  61559=>"001111010",
  61560=>"000111101",
  61561=>"100000111",
  61562=>"110100111",
  61563=>"000011101",
  61564=>"101010110",
  61565=>"110101000",
  61566=>"011101010",
  61567=>"111001000",
  61568=>"001111100",
  61569=>"110100000",
  61570=>"110111100",
  61571=>"101010101",
  61572=>"010010000",
  61573=>"110001101",
  61574=>"010101000",
  61575=>"100100001",
  61576=>"001001111",
  61577=>"001111011",
  61578=>"000000011",
  61579=>"000001011",
  61580=>"000111001",
  61581=>"010101010",
  61582=>"111000110",
  61583=>"101000110",
  61584=>"101011100",
  61585=>"000111100",
  61586=>"100000011",
  61587=>"100001111",
  61588=>"000111011",
  61589=>"000011001",
  61590=>"100001111",
  61591=>"110101001",
  61592=>"000000110",
  61593=>"001101011",
  61594=>"101110111",
  61595=>"101010010",
  61596=>"100000000",
  61597=>"111101001",
  61598=>"110100001",
  61599=>"100001001",
  61600=>"000100000",
  61601=>"011010000",
  61602=>"111100000",
  61603=>"100111000",
  61604=>"110001001",
  61605=>"000011100",
  61606=>"110101010",
  61607=>"111100000",
  61608=>"011000110",
  61609=>"111000100",
  61610=>"011001100",
  61611=>"001110101",
  61612=>"000000101",
  61613=>"111011001",
  61614=>"011111001",
  61615=>"111010100",
  61616=>"110010011",
  61617=>"001011110",
  61618=>"000110110",
  61619=>"110010101",
  61620=>"110011000",
  61621=>"000110001",
  61622=>"001101011",
  61623=>"001111101",
  61624=>"011100110",
  61625=>"111001011",
  61626=>"000100100",
  61627=>"010010110",
  61628=>"001011100",
  61629=>"010010000",
  61630=>"101110010",
  61631=>"011110011",
  61632=>"010001001",
  61633=>"011001101",
  61634=>"010011100",
  61635=>"000100010",
  61636=>"111010011",
  61637=>"111111101",
  61638=>"011110111",
  61639=>"011111101",
  61640=>"001110100",
  61641=>"010101111",
  61642=>"011011011",
  61643=>"111010011",
  61644=>"000001001",
  61645=>"011000001",
  61646=>"001111000",
  61647=>"100111110",
  61648=>"100010010",
  61649=>"101101011",
  61650=>"011100010",
  61651=>"110001110",
  61652=>"000110001",
  61653=>"010111110",
  61654=>"110011101",
  61655=>"101111000",
  61656=>"110010110",
  61657=>"110101110",
  61658=>"000000101",
  61659=>"100101001",
  61660=>"101010001",
  61661=>"101101011",
  61662=>"000110111",
  61663=>"111011000",
  61664=>"011011010",
  61665=>"011000100",
  61666=>"101011001",
  61667=>"000000011",
  61668=>"001110101",
  61669=>"001111111",
  61670=>"011110010",
  61671=>"000010000",
  61672=>"100011110",
  61673=>"101010000",
  61674=>"010110111",
  61675=>"100000011",
  61676=>"001000000",
  61677=>"101010010",
  61678=>"001100110",
  61679=>"001000100",
  61680=>"110111010",
  61681=>"110101000",
  61682=>"001101010",
  61683=>"001101010",
  61684=>"111001011",
  61685=>"011010101",
  61686=>"101010100",
  61687=>"111001001",
  61688=>"000110111",
  61689=>"111010010",
  61690=>"010000110",
  61691=>"010110001",
  61692=>"111101111",
  61693=>"110100010",
  61694=>"011111010",
  61695=>"001110101",
  61696=>"011100000",
  61697=>"000111110",
  61698=>"010100000",
  61699=>"111100001",
  61700=>"001101110",
  61701=>"000100111",
  61702=>"101001111",
  61703=>"101011000",
  61704=>"001001100",
  61705=>"010111011",
  61706=>"111101010",
  61707=>"011111001",
  61708=>"000100111",
  61709=>"101000110",
  61710=>"000101000",
  61711=>"001011000",
  61712=>"111110000",
  61713=>"100110101",
  61714=>"000011001",
  61715=>"100111100",
  61716=>"011011101",
  61717=>"001100100",
  61718=>"100101000",
  61719=>"010100110",
  61720=>"111010100",
  61721=>"111001100",
  61722=>"000010110",
  61723=>"001110010",
  61724=>"000111110",
  61725=>"100100110",
  61726=>"010000010",
  61727=>"000111010",
  61728=>"010010000",
  61729=>"110011000",
  61730=>"001101010",
  61731=>"110000101",
  61732=>"111001001",
  61733=>"011000010",
  61734=>"000000110",
  61735=>"110001100",
  61736=>"010101111",
  61737=>"001001001",
  61738=>"100111110",
  61739=>"111101011",
  61740=>"111011001",
  61741=>"010000010",
  61742=>"000001111",
  61743=>"011011101",
  61744=>"011011011",
  61745=>"111111100",
  61746=>"001011110",
  61747=>"110101100",
  61748=>"000101011",
  61749=>"010000001",
  61750=>"101111010",
  61751=>"011010000",
  61752=>"110101110",
  61753=>"111011010",
  61754=>"001101110",
  61755=>"000110101",
  61756=>"100111001",
  61757=>"101011011",
  61758=>"000110000",
  61759=>"000100000",
  61760=>"100001100",
  61761=>"000111111",
  61762=>"010000110",
  61763=>"100011101",
  61764=>"010001011",
  61765=>"111101101",
  61766=>"101000101",
  61767=>"000110000",
  61768=>"101000111",
  61769=>"110110010",
  61770=>"101001101",
  61771=>"001000000",
  61772=>"001110101",
  61773=>"011011100",
  61774=>"011000110",
  61775=>"101011101",
  61776=>"000000001",
  61777=>"101000011",
  61778=>"000010111",
  61779=>"011000011",
  61780=>"011111110",
  61781=>"100111111",
  61782=>"011100101",
  61783=>"000011011",
  61784=>"101001010",
  61785=>"010001011",
  61786=>"110011101",
  61787=>"100100111",
  61788=>"001100000",
  61789=>"110110010",
  61790=>"101101100",
  61791=>"110000100",
  61792=>"000101010",
  61793=>"111110000",
  61794=>"001111111",
  61795=>"011100110",
  61796=>"101101110",
  61797=>"000000000",
  61798=>"110001010",
  61799=>"110100000",
  61800=>"111011100",
  61801=>"010100110",
  61802=>"100101110",
  61803=>"000110001",
  61804=>"000001010",
  61805=>"001101010",
  61806=>"110000010",
  61807=>"010010111",
  61808=>"101110110",
  61809=>"110110110",
  61810=>"001011110",
  61811=>"000001111",
  61812=>"011101110",
  61813=>"110010000",
  61814=>"111000000",
  61815=>"010001111",
  61816=>"000000100",
  61817=>"001000000",
  61818=>"011001001",
  61819=>"000101011",
  61820=>"110011101",
  61821=>"001011011",
  61822=>"100000100",
  61823=>"010100010",
  61824=>"101110100",
  61825=>"001000010",
  61826=>"000100001",
  61827=>"001100100",
  61828=>"010001000",
  61829=>"011101000",
  61830=>"100011000",
  61831=>"000000010",
  61832=>"111100011",
  61833=>"000001010",
  61834=>"011000001",
  61835=>"001000111",
  61836=>"001011110",
  61837=>"001111100",
  61838=>"111110000",
  61839=>"101001110",
  61840=>"001110011",
  61841=>"010000100",
  61842=>"000000111",
  61843=>"100111111",
  61844=>"111100101",
  61845=>"001000011",
  61846=>"010111011",
  61847=>"000000000",
  61848=>"001101110",
  61849=>"001101001",
  61850=>"010110001",
  61851=>"000110011",
  61852=>"000010000",
  61853=>"001000101",
  61854=>"010101111",
  61855=>"100101100",
  61856=>"000101110",
  61857=>"011010000",
  61858=>"000110000",
  61859=>"111101100",
  61860=>"111111010",
  61861=>"101001001",
  61862=>"101010011",
  61863=>"101010011",
  61864=>"001101000",
  61865=>"110011111",
  61866=>"000010011",
  61867=>"100111011",
  61868=>"011101110",
  61869=>"011000101",
  61870=>"101100011",
  61871=>"101001000",
  61872=>"101010110",
  61873=>"111110111",
  61874=>"001111111",
  61875=>"101101101",
  61876=>"111010111",
  61877=>"011011100",
  61878=>"000011100",
  61879=>"111000110",
  61880=>"010111110",
  61881=>"000101000",
  61882=>"001101010",
  61883=>"011010010",
  61884=>"000010110",
  61885=>"001111110",
  61886=>"010111001",
  61887=>"011110010",
  61888=>"000011011",
  61889=>"101110001",
  61890=>"011001111",
  61891=>"000001110",
  61892=>"011011100",
  61893=>"111111101",
  61894=>"000101010",
  61895=>"101011111",
  61896=>"111011101",
  61897=>"101011100",
  61898=>"000001001",
  61899=>"000100101",
  61900=>"000111110",
  61901=>"100111001",
  61902=>"000101010",
  61903=>"001001000",
  61904=>"001010101",
  61905=>"000001111",
  61906=>"001100011",
  61907=>"000100111",
  61908=>"100110111",
  61909=>"001011000",
  61910=>"011011100",
  61911=>"111101000",
  61912=>"110000001",
  61913=>"100011100",
  61914=>"001100111",
  61915=>"010110000",
  61916=>"001101111",
  61917=>"101010101",
  61918=>"111111111",
  61919=>"110111111",
  61920=>"000000101",
  61921=>"000011001",
  61922=>"010001001",
  61923=>"110101101",
  61924=>"000111011",
  61925=>"011100111",
  61926=>"000111101",
  61927=>"101101101",
  61928=>"110110100",
  61929=>"111111101",
  61930=>"000010101",
  61931=>"000010010",
  61932=>"111000111",
  61933=>"000011000",
  61934=>"100000000",
  61935=>"000010111",
  61936=>"100011111",
  61937=>"000100111",
  61938=>"000000000",
  61939=>"111010110",
  61940=>"111010100",
  61941=>"101000010",
  61942=>"001001000",
  61943=>"101111001",
  61944=>"110110111",
  61945=>"001100000",
  61946=>"001111001",
  61947=>"011101110",
  61948=>"001011110",
  61949=>"000001100",
  61950=>"111110000",
  61951=>"101000001",
  61952=>"101101010",
  61953=>"111000111",
  61954=>"101001000",
  61955=>"000001110",
  61956=>"001110011",
  61957=>"111011010",
  61958=>"011101011",
  61959=>"101100101",
  61960=>"001111100",
  61961=>"000110001",
  61962=>"001101010",
  61963=>"000111011",
  61964=>"100011010",
  61965=>"011111001",
  61966=>"001010011",
  61967=>"010011010",
  61968=>"111010100",
  61969=>"110101111",
  61970=>"000000101",
  61971=>"011111101",
  61972=>"011011101",
  61973=>"111111100",
  61974=>"001001111",
  61975=>"000110000",
  61976=>"001010100",
  61977=>"101010010",
  61978=>"100000110",
  61979=>"000110010",
  61980=>"110011011",
  61981=>"000010100",
  61982=>"100100000",
  61983=>"001011110",
  61984=>"100000010",
  61985=>"011011010",
  61986=>"010110100",
  61987=>"010100000",
  61988=>"111111011",
  61989=>"100010010",
  61990=>"100110110",
  61991=>"100001011",
  61992=>"001101000",
  61993=>"101111000",
  61994=>"011010001",
  61995=>"100000000",
  61996=>"100001110",
  61997=>"010110100",
  61998=>"110111101",
  61999=>"100001111",
  62000=>"000010110",
  62001=>"011000111",
  62002=>"000001001",
  62003=>"110011110",
  62004=>"010111001",
  62005=>"111101110",
  62006=>"000100011",
  62007=>"101011110",
  62008=>"010000000",
  62009=>"010111010",
  62010=>"101110001",
  62011=>"000100011",
  62012=>"001111010",
  62013=>"000000010",
  62014=>"010010111",
  62015=>"110101110",
  62016=>"101001011",
  62017=>"110000111",
  62018=>"101000110",
  62019=>"111001100",
  62020=>"011111010",
  62021=>"111101001",
  62022=>"111011110",
  62023=>"101110011",
  62024=>"011111011",
  62025=>"011101100",
  62026=>"110110001",
  62027=>"110110110",
  62028=>"100110111",
  62029=>"000011011",
  62030=>"101101011",
  62031=>"100101010",
  62032=>"100011111",
  62033=>"000111111",
  62034=>"111110001",
  62035=>"011001000",
  62036=>"010100010",
  62037=>"000110111",
  62038=>"111010110",
  62039=>"101001001",
  62040=>"111010010",
  62041=>"000100110",
  62042=>"001100111",
  62043=>"011000110",
  62044=>"011000110",
  62045=>"011010111",
  62046=>"001101100",
  62047=>"001000010",
  62048=>"111110110",
  62049=>"111011110",
  62050=>"001000010",
  62051=>"101010101",
  62052=>"000100011",
  62053=>"000110001",
  62054=>"000100010",
  62055=>"001011100",
  62056=>"101110101",
  62057=>"101001000",
  62058=>"101110101",
  62059=>"011100000",
  62060=>"000001111",
  62061=>"110110110",
  62062=>"100010001",
  62063=>"101000111",
  62064=>"010000000",
  62065=>"111000110",
  62066=>"101011100",
  62067=>"010011110",
  62068=>"001011001",
  62069=>"101001111",
  62070=>"101011001",
  62071=>"010010100",
  62072=>"011010010",
  62073=>"111100100",
  62074=>"010011111",
  62075=>"110100001",
  62076=>"100101110",
  62077=>"100100011",
  62078=>"111100000",
  62079=>"011000101",
  62080=>"010110011",
  62081=>"111111011",
  62082=>"110000010",
  62083=>"111001100",
  62084=>"100110001",
  62085=>"011111001",
  62086=>"000100011",
  62087=>"111110000",
  62088=>"001010001",
  62089=>"011101111",
  62090=>"011110111",
  62091=>"111110011",
  62092=>"100110100",
  62093=>"001101110",
  62094=>"101010011",
  62095=>"101011110",
  62096=>"000001101",
  62097=>"111111011",
  62098=>"000010110",
  62099=>"111111010",
  62100=>"101001110",
  62101=>"110000100",
  62102=>"100111110",
  62103=>"010101111",
  62104=>"011011111",
  62105=>"100001100",
  62106=>"101011001",
  62107=>"011001110",
  62108=>"001000101",
  62109=>"010110011",
  62110=>"100100100",
  62111=>"001011011",
  62112=>"100111110",
  62113=>"000101101",
  62114=>"110010101",
  62115=>"000011000",
  62116=>"000001101",
  62117=>"001001101",
  62118=>"011000110",
  62119=>"100111010",
  62120=>"110110000",
  62121=>"001100101",
  62122=>"100110011",
  62123=>"010011001",
  62124=>"000100001",
  62125=>"011011001",
  62126=>"111000110",
  62127=>"101111110",
  62128=>"101011000",
  62129=>"011010101",
  62130=>"110001000",
  62131=>"000011011",
  62132=>"000110111",
  62133=>"000000110",
  62134=>"110010100",
  62135=>"111000100",
  62136=>"110001111",
  62137=>"011001101",
  62138=>"110110001",
  62139=>"110101010",
  62140=>"111100111",
  62141=>"010111111",
  62142=>"111001010",
  62143=>"010101000",
  62144=>"101010000",
  62145=>"101110110",
  62146=>"001010101",
  62147=>"110111111",
  62148=>"101101010",
  62149=>"010100000",
  62150=>"101011100",
  62151=>"110010111",
  62152=>"110010000",
  62153=>"110010010",
  62154=>"100010011",
  62155=>"100000111",
  62156=>"110010111",
  62157=>"111111010",
  62158=>"010011100",
  62159=>"010110011",
  62160=>"100010001",
  62161=>"111010000",
  62162=>"110111001",
  62163=>"111111101",
  62164=>"100000100",
  62165=>"001001010",
  62166=>"000000100",
  62167=>"000011001",
  62168=>"001110010",
  62169=>"100111111",
  62170=>"000010100",
  62171=>"110011011",
  62172=>"000011100",
  62173=>"000110000",
  62174=>"000010000",
  62175=>"101010001",
  62176=>"110000101",
  62177=>"100000111",
  62178=>"011010011",
  62179=>"000110100",
  62180=>"000000011",
  62181=>"011011000",
  62182=>"000000000",
  62183=>"000111111",
  62184=>"100011001",
  62185=>"101010011",
  62186=>"100111010",
  62187=>"011110100",
  62188=>"000000011",
  62189=>"010000000",
  62190=>"110111110",
  62191=>"001011011",
  62192=>"001011110",
  62193=>"001010010",
  62194=>"001000001",
  62195=>"111111101",
  62196=>"010110000",
  62197=>"000011010",
  62198=>"001000000",
  62199=>"000111100",
  62200=>"001000101",
  62201=>"110110111",
  62202=>"100011100",
  62203=>"001001000",
  62204=>"100011001",
  62205=>"010001011",
  62206=>"110000000",
  62207=>"011000100",
  62208=>"111011110",
  62209=>"110000001",
  62210=>"110101111",
  62211=>"101010001",
  62212=>"100100100",
  62213=>"100010110",
  62214=>"111000110",
  62215=>"010011101",
  62216=>"100000000",
  62217=>"100110111",
  62218=>"100110001",
  62219=>"110010010",
  62220=>"101000001",
  62221=>"111100100",
  62222=>"100000000",
  62223=>"110011001",
  62224=>"001010001",
  62225=>"010111000",
  62226=>"011101110",
  62227=>"011100011",
  62228=>"110100101",
  62229=>"000111101",
  62230=>"011000001",
  62231=>"011011000",
  62232=>"100010001",
  62233=>"111101010",
  62234=>"001000110",
  62235=>"001011100",
  62236=>"101100101",
  62237=>"001101100",
  62238=>"000000111",
  62239=>"000101011",
  62240=>"100110011",
  62241=>"100000011",
  62242=>"011001011",
  62243=>"111111011",
  62244=>"100100100",
  62245=>"111000110",
  62246=>"111111011",
  62247=>"000011111",
  62248=>"110110000",
  62249=>"101100101",
  62250=>"111110101",
  62251=>"010000100",
  62252=>"110000101",
  62253=>"100000010",
  62254=>"010000111",
  62255=>"111111110",
  62256=>"001010001",
  62257=>"000001111",
  62258=>"101110000",
  62259=>"110010010",
  62260=>"000000011",
  62261=>"010010110",
  62262=>"111010100",
  62263=>"100100001",
  62264=>"011100000",
  62265=>"000011011",
  62266=>"101000100",
  62267=>"111011011",
  62268=>"110000000",
  62269=>"011010100",
  62270=>"111001011",
  62271=>"110110010",
  62272=>"001100100",
  62273=>"100000000",
  62274=>"100000101",
  62275=>"000100001",
  62276=>"110000100",
  62277=>"101010011",
  62278=>"010110011",
  62279=>"110101101",
  62280=>"110010111",
  62281=>"111000110",
  62282=>"001001000",
  62283=>"100110000",
  62284=>"011011001",
  62285=>"111100100",
  62286=>"111101101",
  62287=>"001011001",
  62288=>"001010000",
  62289=>"001011011",
  62290=>"011110101",
  62291=>"110100110",
  62292=>"111011000",
  62293=>"111011111",
  62294=>"001000011",
  62295=>"111100111",
  62296=>"011010010",
  62297=>"111100000",
  62298=>"000011111",
  62299=>"000001111",
  62300=>"000010100",
  62301=>"010001101",
  62302=>"000001000",
  62303=>"011011000",
  62304=>"110001111",
  62305=>"100011010",
  62306=>"000110110",
  62307=>"110000010",
  62308=>"001000011",
  62309=>"011011111",
  62310=>"000011111",
  62311=>"000101000",
  62312=>"010011001",
  62313=>"101101010",
  62314=>"110000111",
  62315=>"110100101",
  62316=>"100010101",
  62317=>"110000010",
  62318=>"000110000",
  62319=>"011011100",
  62320=>"101010110",
  62321=>"101111110",
  62322=>"111001000",
  62323=>"010111000",
  62324=>"011110101",
  62325=>"010111001",
  62326=>"100100011",
  62327=>"100111111",
  62328=>"111111010",
  62329=>"010011110",
  62330=>"000010010",
  62331=>"011110110",
  62332=>"001001000",
  62333=>"010000000",
  62334=>"111010111",
  62335=>"001100110",
  62336=>"101000000",
  62337=>"110100111",
  62338=>"000111111",
  62339=>"001011011",
  62340=>"000011010",
  62341=>"001010001",
  62342=>"000001110",
  62343=>"111001101",
  62344=>"111100101",
  62345=>"001001001",
  62346=>"001011001",
  62347=>"000110010",
  62348=>"111011101",
  62349=>"010010100",
  62350=>"001001101",
  62351=>"111000110",
  62352=>"010011111",
  62353=>"111101000",
  62354=>"111001111",
  62355=>"101010011",
  62356=>"001100001",
  62357=>"001100000",
  62358=>"110111010",
  62359=>"100000001",
  62360=>"001000010",
  62361=>"010010010",
  62362=>"100110011",
  62363=>"100011011",
  62364=>"011010100",
  62365=>"001000101",
  62366=>"101111110",
  62367=>"111101000",
  62368=>"101000000",
  62369=>"010110101",
  62370=>"111111101",
  62371=>"010000011",
  62372=>"010001110",
  62373=>"101100111",
  62374=>"000001010",
  62375=>"011000011",
  62376=>"001100010",
  62377=>"000100100",
  62378=>"110010010",
  62379=>"110101111",
  62380=>"100010011",
  62381=>"000100111",
  62382=>"110010101",
  62383=>"001101001",
  62384=>"000111001",
  62385=>"100011100",
  62386=>"001101000",
  62387=>"000101100",
  62388=>"110001001",
  62389=>"011110010",
  62390=>"101101111",
  62391=>"110111101",
  62392=>"011100111",
  62393=>"111001010",
  62394=>"111101101",
  62395=>"111011100",
  62396=>"110110110",
  62397=>"000000010",
  62398=>"011011011",
  62399=>"110110011",
  62400=>"111011001",
  62401=>"001110111",
  62402=>"111101000",
  62403=>"110001111",
  62404=>"010100001",
  62405=>"110110101",
  62406=>"010101100",
  62407=>"010000010",
  62408=>"000100010",
  62409=>"001110100",
  62410=>"011101111",
  62411=>"011010110",
  62412=>"110001110",
  62413=>"010000011",
  62414=>"110011001",
  62415=>"010100100",
  62416=>"100111000",
  62417=>"110001011",
  62418=>"001100001",
  62419=>"100011000",
  62420=>"000111111",
  62421=>"000011010",
  62422=>"110100100",
  62423=>"011101011",
  62424=>"000010111",
  62425=>"010101110",
  62426=>"111001011",
  62427=>"010010000",
  62428=>"000010000",
  62429=>"000100110",
  62430=>"100001111",
  62431=>"011000001",
  62432=>"000110011",
  62433=>"001010000",
  62434=>"000010101",
  62435=>"010111111",
  62436=>"010010000",
  62437=>"111110111",
  62438=>"110111111",
  62439=>"010111001",
  62440=>"111000000",
  62441=>"000000010",
  62442=>"001111011",
  62443=>"011110111",
  62444=>"111001101",
  62445=>"111111110",
  62446=>"011100010",
  62447=>"111001111",
  62448=>"100100110",
  62449=>"111101011",
  62450=>"100101110",
  62451=>"101100110",
  62452=>"011001111",
  62453=>"101010111",
  62454=>"001000010",
  62455=>"001111111",
  62456=>"101111111",
  62457=>"100000110",
  62458=>"111000010",
  62459=>"001000110",
  62460=>"100101000",
  62461=>"100100000",
  62462=>"000111101",
  62463=>"000110110",
  62464=>"010100110",
  62465=>"111011011",
  62466=>"101101011",
  62467=>"000010110",
  62468=>"101000100",
  62469=>"110010100",
  62470=>"001100011",
  62471=>"001000111",
  62472=>"000100101",
  62473=>"111100000",
  62474=>"100110010",
  62475=>"001000010",
  62476=>"101001011",
  62477=>"111101011",
  62478=>"101011010",
  62479=>"011110010",
  62480=>"010001011",
  62481=>"000011000",
  62482=>"101111110",
  62483=>"100000000",
  62484=>"111111011",
  62485=>"110110100",
  62486=>"011111111",
  62487=>"100111000",
  62488=>"100101010",
  62489=>"100110000",
  62490=>"011000001",
  62491=>"110101111",
  62492=>"001110011",
  62493=>"101101100",
  62494=>"111110101",
  62495=>"000001001",
  62496=>"000010110",
  62497=>"111111001",
  62498=>"000110001",
  62499=>"101010010",
  62500=>"110001110",
  62501=>"010001110",
  62502=>"011010011",
  62503=>"010101001",
  62504=>"001111001",
  62505=>"111000000",
  62506=>"001001010",
  62507=>"101111100",
  62508=>"000000010",
  62509=>"110001101",
  62510=>"011100000",
  62511=>"100000010",
  62512=>"010110000",
  62513=>"111100011",
  62514=>"110110101",
  62515=>"111111000",
  62516=>"000000100",
  62517=>"001101100",
  62518=>"000110001",
  62519=>"100000110",
  62520=>"111110100",
  62521=>"111111011",
  62522=>"011111001",
  62523=>"110010110",
  62524=>"000000001",
  62525=>"000110100",
  62526=>"100100010",
  62527=>"001001011",
  62528=>"011010101",
  62529=>"101010100",
  62530=>"100010001",
  62531=>"100001010",
  62532=>"001001100",
  62533=>"110001010",
  62534=>"111011000",
  62535=>"001111010",
  62536=>"110011010",
  62537=>"000100011",
  62538=>"001000110",
  62539=>"111110010",
  62540=>"000100001",
  62541=>"110010101",
  62542=>"110111111",
  62543=>"010011010",
  62544=>"110100110",
  62545=>"110110111",
  62546=>"101000110",
  62547=>"000101010",
  62548=>"111111000",
  62549=>"110101000",
  62550=>"111100100",
  62551=>"100111110",
  62552=>"111000111",
  62553=>"101111011",
  62554=>"000110010",
  62555=>"110010011",
  62556=>"001110100",
  62557=>"011000000",
  62558=>"101101010",
  62559=>"100101101",
  62560=>"110001011",
  62561=>"010110000",
  62562=>"010111111",
  62563=>"101101111",
  62564=>"010000010",
  62565=>"101001010",
  62566=>"111100110",
  62567=>"001010110",
  62568=>"000010110",
  62569=>"011111001",
  62570=>"011001111",
  62571=>"001001100",
  62572=>"101100111",
  62573=>"010000100",
  62574=>"001001100",
  62575=>"000011011",
  62576=>"011101101",
  62577=>"110100010",
  62578=>"010000111",
  62579=>"111110000",
  62580=>"110110100",
  62581=>"000111111",
  62582=>"111101000",
  62583=>"010110100",
  62584=>"101000110",
  62585=>"010001100",
  62586=>"000000101",
  62587=>"010110001",
  62588=>"111110101",
  62589=>"000010111",
  62590=>"111001000",
  62591=>"000011101",
  62592=>"010000010",
  62593=>"100100000",
  62594=>"010100100",
  62595=>"111100101",
  62596=>"011001100",
  62597=>"010000110",
  62598=>"000000100",
  62599=>"001001010",
  62600=>"011101101",
  62601=>"110111000",
  62602=>"001100000",
  62603=>"010000110",
  62604=>"111101011",
  62605=>"101001100",
  62606=>"101000000",
  62607=>"100111100",
  62608=>"010011011",
  62609=>"001010101",
  62610=>"001110111",
  62611=>"111111010",
  62612=>"110111111",
  62613=>"111010100",
  62614=>"001111110",
  62615=>"101100111",
  62616=>"000100000",
  62617=>"111110001",
  62618=>"001011001",
  62619=>"101100011",
  62620=>"100111000",
  62621=>"000011011",
  62622=>"000010111",
  62623=>"011011001",
  62624=>"111010100",
  62625=>"100000100",
  62626=>"101011111",
  62627=>"011011000",
  62628=>"110010011",
  62629=>"110001000",
  62630=>"011101011",
  62631=>"101011000",
  62632=>"100000010",
  62633=>"011001110",
  62634=>"110011010",
  62635=>"101110111",
  62636=>"110010100",
  62637=>"101110000",
  62638=>"100000110",
  62639=>"100100100",
  62640=>"100100000",
  62641=>"100110101",
  62642=>"000000000",
  62643=>"100011010",
  62644=>"100100000",
  62645=>"110000101",
  62646=>"110010110",
  62647=>"101111110",
  62648=>"010010100",
  62649=>"001011010",
  62650=>"010000010",
  62651=>"111011100",
  62652=>"101010000",
  62653=>"111011101",
  62654=>"011000010",
  62655=>"101000001",
  62656=>"010101011",
  62657=>"011010111",
  62658=>"000000001",
  62659=>"000011001",
  62660=>"011010010",
  62661=>"110010000",
  62662=>"000110111",
  62663=>"000001011",
  62664=>"110111101",
  62665=>"111011100",
  62666=>"000000100",
  62667=>"101011010",
  62668=>"001100111",
  62669=>"000000111",
  62670=>"000100100",
  62671=>"110111110",
  62672=>"101101110",
  62673=>"001010001",
  62674=>"000111111",
  62675=>"000001100",
  62676=>"110011100",
  62677=>"000001000",
  62678=>"001101000",
  62679=>"100000000",
  62680=>"100010001",
  62681=>"001001100",
  62682=>"101000001",
  62683=>"011010011",
  62684=>"001000011",
  62685=>"011001010",
  62686=>"000100011",
  62687=>"000011001",
  62688=>"001000011",
  62689=>"011011110",
  62690=>"101010110",
  62691=>"100010101",
  62692=>"001000100",
  62693=>"011101001",
  62694=>"100111111",
  62695=>"111001101",
  62696=>"000001010",
  62697=>"101001010",
  62698=>"110000010",
  62699=>"101101011",
  62700=>"011110000",
  62701=>"000001110",
  62702=>"111010110",
  62703=>"011010000",
  62704=>"010110101",
  62705=>"110111100",
  62706=>"110001101",
  62707=>"000111100",
  62708=>"000010110",
  62709=>"100110010",
  62710=>"110101110",
  62711=>"000111000",
  62712=>"110101000",
  62713=>"100101010",
  62714=>"011001000",
  62715=>"110111100",
  62716=>"010101101",
  62717=>"111010101",
  62718=>"100000100",
  62719=>"111111000",
  62720=>"101010110",
  62721=>"010000110",
  62722=>"101100111",
  62723=>"010000110",
  62724=>"010001010",
  62725=>"110111111",
  62726=>"101000111",
  62727=>"100111000",
  62728=>"001000001",
  62729=>"011110000",
  62730=>"110101101",
  62731=>"011100010",
  62732=>"110100011",
  62733=>"001110000",
  62734=>"111100011",
  62735=>"000100010",
  62736=>"010001101",
  62737=>"001101000",
  62738=>"101100001",
  62739=>"100010101",
  62740=>"001000001",
  62741=>"111100100",
  62742=>"000101111",
  62743=>"101010011",
  62744=>"111011100",
  62745=>"000000010",
  62746=>"011000110",
  62747=>"011001111",
  62748=>"000000101",
  62749=>"101010001",
  62750=>"011001000",
  62751=>"000101110",
  62752=>"000101100",
  62753=>"111110101",
  62754=>"111110001",
  62755=>"100001100",
  62756=>"111110110",
  62757=>"100011100",
  62758=>"100101000",
  62759=>"000000001",
  62760=>"000001010",
  62761=>"011001100",
  62762=>"001000100",
  62763=>"100111000",
  62764=>"011110001",
  62765=>"010000010",
  62766=>"011010000",
  62767=>"111110100",
  62768=>"010010011",
  62769=>"011110001",
  62770=>"110101010",
  62771=>"101101100",
  62772=>"011111010",
  62773=>"111010000",
  62774=>"010000001",
  62775=>"100000000",
  62776=>"110001000",
  62777=>"111101100",
  62778=>"011011011",
  62779=>"100111010",
  62780=>"110110110",
  62781=>"011101100",
  62782=>"011001011",
  62783=>"111001001",
  62784=>"001111001",
  62785=>"001011011",
  62786=>"011011111",
  62787=>"100101001",
  62788=>"110110101",
  62789=>"011011110",
  62790=>"001101000",
  62791=>"010111111",
  62792=>"001010110",
  62793=>"011010010",
  62794=>"001001111",
  62795=>"110111110",
  62796=>"110011000",
  62797=>"000110100",
  62798=>"000010111",
  62799=>"011011010",
  62800=>"011100110",
  62801=>"101011010",
  62802=>"001000010",
  62803=>"101000110",
  62804=>"010001111",
  62805=>"010110001",
  62806=>"011011111",
  62807=>"011110110",
  62808=>"001100000",
  62809=>"110010111",
  62810=>"111110010",
  62811=>"011000011",
  62812=>"100101011",
  62813=>"011100111",
  62814=>"001000010",
  62815=>"010000001",
  62816=>"001101000",
  62817=>"010000100",
  62818=>"000010110",
  62819=>"000100101",
  62820=>"100110110",
  62821=>"110011110",
  62822=>"110010110",
  62823=>"000001010",
  62824=>"100101010",
  62825=>"100001001",
  62826=>"110101001",
  62827=>"100010011",
  62828=>"010111101",
  62829=>"110001111",
  62830=>"111110010",
  62831=>"001101010",
  62832=>"100000001",
  62833=>"000000001",
  62834=>"111101111",
  62835=>"011110010",
  62836=>"001010111",
  62837=>"101110100",
  62838=>"000110011",
  62839=>"000101111",
  62840=>"101001010",
  62841=>"011101100",
  62842=>"000111111",
  62843=>"011010101",
  62844=>"010010111",
  62845=>"001111010",
  62846=>"000010110",
  62847=>"100000100",
  62848=>"101010010",
  62849=>"011110111",
  62850=>"101101010",
  62851=>"101001111",
  62852=>"111100111",
  62853=>"001011110",
  62854=>"101111001",
  62855=>"110100010",
  62856=>"000010100",
  62857=>"111000110",
  62858=>"110010100",
  62859=>"011101101",
  62860=>"111101100",
  62861=>"100110111",
  62862=>"010101111",
  62863=>"111101101",
  62864=>"011010011",
  62865=>"000000000",
  62866=>"100111001",
  62867=>"001111111",
  62868=>"100011101",
  62869=>"001111000",
  62870=>"111110101",
  62871=>"010101011",
  62872=>"001111000",
  62873=>"001100011",
  62874=>"000111011",
  62875=>"010111110",
  62876=>"001110100",
  62877=>"100110011",
  62878=>"101100100",
  62879=>"001110011",
  62880=>"011100100",
  62881=>"001000010",
  62882=>"110001011",
  62883=>"010101100",
  62884=>"001011011",
  62885=>"001100000",
  62886=>"000110111",
  62887=>"111110001",
  62888=>"011000111",
  62889=>"011100110",
  62890=>"111010000",
  62891=>"001000000",
  62892=>"000111101",
  62893=>"010010001",
  62894=>"111001101",
  62895=>"010001110",
  62896=>"000110000",
  62897=>"000010100",
  62898=>"011001101",
  62899=>"101000110",
  62900=>"000000100",
  62901=>"110000011",
  62902=>"100100000",
  62903=>"010110101",
  62904=>"011011100",
  62905=>"100000110",
  62906=>"100011101",
  62907=>"001101011",
  62908=>"011010000",
  62909=>"010010100",
  62910=>"111000011",
  62911=>"110110001",
  62912=>"001011010",
  62913=>"100110100",
  62914=>"000011001",
  62915=>"111010001",
  62916=>"110101010",
  62917=>"000110110",
  62918=>"111101100",
  62919=>"000101001",
  62920=>"001110100",
  62921=>"001100110",
  62922=>"001010011",
  62923=>"110000010",
  62924=>"111101011",
  62925=>"101111011",
  62926=>"101111101",
  62927=>"011000110",
  62928=>"000011110",
  62929=>"100001101",
  62930=>"010101111",
  62931=>"101010011",
  62932=>"011001010",
  62933=>"100000000",
  62934=>"001010000",
  62935=>"001100011",
  62936=>"000101110",
  62937=>"011111011",
  62938=>"101100000",
  62939=>"000110011",
  62940=>"110101010",
  62941=>"000110010",
  62942=>"110101101",
  62943=>"000101100",
  62944=>"000000011",
  62945=>"100110010",
  62946=>"111111100",
  62947=>"110100101",
  62948=>"001010110",
  62949=>"101000111",
  62950=>"111001001",
  62951=>"100101000",
  62952=>"100110000",
  62953=>"100101000",
  62954=>"001101010",
  62955=>"001100100",
  62956=>"010010101",
  62957=>"011010000",
  62958=>"010001010",
  62959=>"010000111",
  62960=>"111010010",
  62961=>"110001010",
  62962=>"001011101",
  62963=>"101111011",
  62964=>"101110111",
  62965=>"100100110",
  62966=>"101011111",
  62967=>"110100000",
  62968=>"100010000",
  62969=>"000110000",
  62970=>"101001110",
  62971=>"000110110",
  62972=>"111111110",
  62973=>"000111001",
  62974=>"001010011",
  62975=>"100110001",
  62976=>"101011011",
  62977=>"000000011",
  62978=>"010011101",
  62979=>"100001001",
  62980=>"011100111",
  62981=>"001111010",
  62982=>"010111001",
  62983=>"101101000",
  62984=>"100100001",
  62985=>"111110111",
  62986=>"011100100",
  62987=>"010011101",
  62988=>"110111011",
  62989=>"000010011",
  62990=>"001111000",
  62991=>"110101111",
  62992=>"011110011",
  62993=>"010001110",
  62994=>"010000101",
  62995=>"010100101",
  62996=>"101111111",
  62997=>"000000001",
  62998=>"001111001",
  62999=>"010010001",
  63000=>"111110100",
  63001=>"111101011",
  63002=>"001001001",
  63003=>"000010100",
  63004=>"000000000",
  63005=>"011101000",
  63006=>"000100110",
  63007=>"011011101",
  63008=>"000100000",
  63009=>"001011110",
  63010=>"000111001",
  63011=>"001100001",
  63012=>"111011100",
  63013=>"011010001",
  63014=>"111011010",
  63015=>"011000000",
  63016=>"100001111",
  63017=>"010110101",
  63018=>"100010101",
  63019=>"011111110",
  63020=>"000010111",
  63021=>"011100001",
  63022=>"100101010",
  63023=>"000001100",
  63024=>"110111100",
  63025=>"110111000",
  63026=>"111111101",
  63027=>"111110001",
  63028=>"110010001",
  63029=>"001000101",
  63030=>"001011010",
  63031=>"111111110",
  63032=>"001100101",
  63033=>"101101101",
  63034=>"010101011",
  63035=>"010010011",
  63036=>"100000111",
  63037=>"111111101",
  63038=>"011110000",
  63039=>"010000010",
  63040=>"110110010",
  63041=>"001110010",
  63042=>"111000011",
  63043=>"011100011",
  63044=>"001100011",
  63045=>"111011011",
  63046=>"000110010",
  63047=>"110100111",
  63048=>"100110001",
  63049=>"001000110",
  63050=>"001001101",
  63051=>"111111111",
  63052=>"011011011",
  63053=>"001010000",
  63054=>"101100010",
  63055=>"010110011",
  63056=>"101001010",
  63057=>"001111011",
  63058=>"111100000",
  63059=>"110000011",
  63060=>"110000000",
  63061=>"111111011",
  63062=>"110101111",
  63063=>"110010110",
  63064=>"010010001",
  63065=>"000011000",
  63066=>"100011101",
  63067=>"100000010",
  63068=>"111000100",
  63069=>"100110100",
  63070=>"111011100",
  63071=>"011100011",
  63072=>"101101001",
  63073=>"001111001",
  63074=>"001011111",
  63075=>"101000100",
  63076=>"110011001",
  63077=>"101100110",
  63078=>"010001101",
  63079=>"111000111",
  63080=>"010110100",
  63081=>"011010010",
  63082=>"011111110",
  63083=>"001001000",
  63084=>"111110000",
  63085=>"110110000",
  63086=>"101100101",
  63087=>"010100011",
  63088=>"000110011",
  63089=>"001111110",
  63090=>"101110101",
  63091=>"110101010",
  63092=>"010010100",
  63093=>"111110001",
  63094=>"101011111",
  63095=>"010011011",
  63096=>"000010010",
  63097=>"101111110",
  63098=>"000001110",
  63099=>"100111111",
  63100=>"010000110",
  63101=>"010110101",
  63102=>"111010000",
  63103=>"011001001",
  63104=>"111011000",
  63105=>"101111010",
  63106=>"100110000",
  63107=>"001001101",
  63108=>"000110001",
  63109=>"111100101",
  63110=>"010011111",
  63111=>"011011010",
  63112=>"011010101",
  63113=>"100100001",
  63114=>"100011011",
  63115=>"111101000",
  63116=>"011001100",
  63117=>"010111010",
  63118=>"010010100",
  63119=>"110100001",
  63120=>"001100110",
  63121=>"000100110",
  63122=>"000110000",
  63123=>"010000111",
  63124=>"110010111",
  63125=>"100111011",
  63126=>"010001100",
  63127=>"001111110",
  63128=>"001010011",
  63129=>"001100111",
  63130=>"110110100",
  63131=>"001110100",
  63132=>"111111010",
  63133=>"110001101",
  63134=>"000011001",
  63135=>"011010000",
  63136=>"011110101",
  63137=>"000000001",
  63138=>"110011101",
  63139=>"001010000",
  63140=>"100110100",
  63141=>"011010011",
  63142=>"111101010",
  63143=>"001110010",
  63144=>"111100101",
  63145=>"100000111",
  63146=>"010011010",
  63147=>"010101001",
  63148=>"011101000",
  63149=>"111011100",
  63150=>"001101101",
  63151=>"000011001",
  63152=>"111011100",
  63153=>"011000011",
  63154=>"001110111",
  63155=>"110011110",
  63156=>"001111001",
  63157=>"111011011",
  63158=>"010100110",
  63159=>"111000010",
  63160=>"100111001",
  63161=>"000101000",
  63162=>"100111111",
  63163=>"011001110",
  63164=>"010000011",
  63165=>"001111001",
  63166=>"000011111",
  63167=>"011111111",
  63168=>"001001001",
  63169=>"111101000",
  63170=>"111100001",
  63171=>"111101001",
  63172=>"010100000",
  63173=>"100101111",
  63174=>"101010000",
  63175=>"110111111",
  63176=>"111100000",
  63177=>"100110000",
  63178=>"101101010",
  63179=>"100101101",
  63180=>"000100011",
  63181=>"100010010",
  63182=>"110011010",
  63183=>"000111001",
  63184=>"111000001",
  63185=>"111011110",
  63186=>"100101000",
  63187=>"001000110",
  63188=>"001001110",
  63189=>"001101110",
  63190=>"100111010",
  63191=>"000110011",
  63192=>"000010010",
  63193=>"001000110",
  63194=>"010111110",
  63195=>"001100000",
  63196=>"111110101",
  63197=>"101001111",
  63198=>"010010111",
  63199=>"000010011",
  63200=>"100000111",
  63201=>"101000100",
  63202=>"001100001",
  63203=>"001011011",
  63204=>"111101001",
  63205=>"010000111",
  63206=>"101100000",
  63207=>"010011111",
  63208=>"000000000",
  63209=>"100000001",
  63210=>"100111110",
  63211=>"110010010",
  63212=>"101110100",
  63213=>"101000011",
  63214=>"011001011",
  63215=>"101011011",
  63216=>"111110110",
  63217=>"011001100",
  63218=>"111100111",
  63219=>"010110011",
  63220=>"010100001",
  63221=>"001000010",
  63222=>"011110110",
  63223=>"110101001",
  63224=>"011100000",
  63225=>"101100000",
  63226=>"100101100",
  63227=>"000100100",
  63228=>"111001100",
  63229=>"011001011",
  63230=>"011000111",
  63231=>"000000010",
  63232=>"010001101",
  63233=>"111111111",
  63234=>"101010101",
  63235=>"101100010",
  63236=>"110101110",
  63237=>"001110001",
  63238=>"010000101",
  63239=>"110101000",
  63240=>"111000011",
  63241=>"101111100",
  63242=>"110100100",
  63243=>"000100010",
  63244=>"010001000",
  63245=>"011010101",
  63246=>"101010100",
  63247=>"011111100",
  63248=>"110011001",
  63249=>"010011101",
  63250=>"100000011",
  63251=>"111000000",
  63252=>"010010111",
  63253=>"110000111",
  63254=>"111110011",
  63255=>"100110001",
  63256=>"010110001",
  63257=>"010010110",
  63258=>"010011010",
  63259=>"111011110",
  63260=>"001110000",
  63261=>"111100100",
  63262=>"101010101",
  63263=>"111111011",
  63264=>"011001011",
  63265=>"100101001",
  63266=>"001011010",
  63267=>"001110101",
  63268=>"000011111",
  63269=>"111001100",
  63270=>"110010011",
  63271=>"001100011",
  63272=>"110111111",
  63273=>"010100001",
  63274=>"011011111",
  63275=>"110001100",
  63276=>"011001001",
  63277=>"000110111",
  63278=>"110000010",
  63279=>"100010011",
  63280=>"101001111",
  63281=>"010000111",
  63282=>"110011111",
  63283=>"110001100",
  63284=>"100111110",
  63285=>"100000101",
  63286=>"111101110",
  63287=>"100111101",
  63288=>"101000010",
  63289=>"110100011",
  63290=>"110111000",
  63291=>"101111101",
  63292=>"001000100",
  63293=>"110110111",
  63294=>"111001101",
  63295=>"110011111",
  63296=>"000001110",
  63297=>"101001100",
  63298=>"110101111",
  63299=>"010111000",
  63300=>"111000101",
  63301=>"001101110",
  63302=>"101011010",
  63303=>"111110111",
  63304=>"010101111",
  63305=>"000111100",
  63306=>"011011110",
  63307=>"001110011",
  63308=>"100111001",
  63309=>"000001010",
  63310=>"111110111",
  63311=>"001111010",
  63312=>"111010101",
  63313=>"000010010",
  63314=>"001101110",
  63315=>"010010101",
  63316=>"100110001",
  63317=>"110010111",
  63318=>"000100100",
  63319=>"101100010",
  63320=>"000101101",
  63321=>"100010101",
  63322=>"101001011",
  63323=>"011001111",
  63324=>"110101100",
  63325=>"001000110",
  63326=>"100110100",
  63327=>"111011101",
  63328=>"001111110",
  63329=>"110110111",
  63330=>"101011111",
  63331=>"011010110",
  63332=>"011101101",
  63333=>"010111000",
  63334=>"010101000",
  63335=>"101110111",
  63336=>"001000100",
  63337=>"010110001",
  63338=>"000100000",
  63339=>"110011110",
  63340=>"100010110",
  63341=>"001100100",
  63342=>"110110100",
  63343=>"100111011",
  63344=>"001001001",
  63345=>"000010111",
  63346=>"110000111",
  63347=>"110011100",
  63348=>"111111100",
  63349=>"101100100",
  63350=>"101111011",
  63351=>"011110000",
  63352=>"110011101",
  63353=>"000111000",
  63354=>"000111111",
  63355=>"111111011",
  63356=>"110110001",
  63357=>"111111101",
  63358=>"111010010",
  63359=>"011111100",
  63360=>"001110110",
  63361=>"011111010",
  63362=>"100000011",
  63363=>"001010111",
  63364=>"010110011",
  63365=>"101111100",
  63366=>"000100100",
  63367=>"101110010",
  63368=>"011101001",
  63369=>"011011010",
  63370=>"110011001",
  63371=>"101100100",
  63372=>"001010110",
  63373=>"110101010",
  63374=>"010100100",
  63375=>"111001011",
  63376=>"100111011",
  63377=>"010000100",
  63378=>"010110000",
  63379=>"111111010",
  63380=>"100111000",
  63381=>"001110010",
  63382=>"001110010",
  63383=>"111000000",
  63384=>"111101001",
  63385=>"000100010",
  63386=>"111111100",
  63387=>"110101000",
  63388=>"010100101",
  63389=>"010000001",
  63390=>"110101010",
  63391=>"001100101",
  63392=>"001100111",
  63393=>"100010111",
  63394=>"001000110",
  63395=>"100010111",
  63396=>"000011001",
  63397=>"110001000",
  63398=>"111111111",
  63399=>"100110000",
  63400=>"000000100",
  63401=>"111100001",
  63402=>"011010000",
  63403=>"110101000",
  63404=>"000111000",
  63405=>"000101110",
  63406=>"101111101",
  63407=>"000001110",
  63408=>"001011101",
  63409=>"111111100",
  63410=>"001010100",
  63411=>"110101011",
  63412=>"100110011",
  63413=>"100011110",
  63414=>"000010001",
  63415=>"100100110",
  63416=>"001000000",
  63417=>"101100011",
  63418=>"101010010",
  63419=>"011010010",
  63420=>"101011110",
  63421=>"101011001",
  63422=>"010010001",
  63423=>"111110011",
  63424=>"011010000",
  63425=>"000110000",
  63426=>"000011011",
  63427=>"000010101",
  63428=>"011000001",
  63429=>"111110000",
  63430=>"000110010",
  63431=>"000001010",
  63432=>"000001001",
  63433=>"000110101",
  63434=>"001010111",
  63435=>"010001101",
  63436=>"101110101",
  63437=>"101110010",
  63438=>"101011100",
  63439=>"111000011",
  63440=>"000001000",
  63441=>"111101111",
  63442=>"001001010",
  63443=>"011000010",
  63444=>"101110111",
  63445=>"111100111",
  63446=>"010001000",
  63447=>"000110001",
  63448=>"001101110",
  63449=>"100000010",
  63450=>"010100101",
  63451=>"100000000",
  63452=>"010110001",
  63453=>"000110001",
  63454=>"011011001",
  63455=>"011001010",
  63456=>"010001111",
  63457=>"101001101",
  63458=>"111000001",
  63459=>"101011111",
  63460=>"101010000",
  63461=>"101010001",
  63462=>"101100111",
  63463=>"010100100",
  63464=>"000100011",
  63465=>"110111011",
  63466=>"000101001",
  63467=>"111110110",
  63468=>"111111101",
  63469=>"011110011",
  63470=>"011101110",
  63471=>"111001011",
  63472=>"011010110",
  63473=>"000101000",
  63474=>"110110001",
  63475=>"000110110",
  63476=>"001000111",
  63477=>"000100100",
  63478=>"010111010",
  63479=>"000010000",
  63480=>"111101101",
  63481=>"110010110",
  63482=>"011000000",
  63483=>"111101001",
  63484=>"001100001",
  63485=>"000000010",
  63486=>"111110100",
  63487=>"000000001",
  63488=>"110100111",
  63489=>"011000000",
  63490=>"110101101",
  63491=>"100011111",
  63492=>"100111010",
  63493=>"101110110",
  63494=>"001011111",
  63495=>"000001010",
  63496=>"110100000",
  63497=>"001111011",
  63498=>"010001111",
  63499=>"001011110",
  63500=>"110110100",
  63501=>"010111011",
  63502=>"100101001",
  63503=>"110110011",
  63504=>"100111110",
  63505=>"101111110",
  63506=>"101010110",
  63507=>"000101101",
  63508=>"000110100",
  63509=>"100110000",
  63510=>"110100011",
  63511=>"111001111",
  63512=>"001100111",
  63513=>"101011011",
  63514=>"111111001",
  63515=>"001100100",
  63516=>"110110111",
  63517=>"100010001",
  63518=>"111011000",
  63519=>"000010001",
  63520=>"101010100",
  63521=>"101000001",
  63522=>"010110100",
  63523=>"110101100",
  63524=>"110011010",
  63525=>"000000010",
  63526=>"000001010",
  63527=>"111111010",
  63528=>"100010001",
  63529=>"100000111",
  63530=>"111110011",
  63531=>"111111111",
  63532=>"011110011",
  63533=>"100010101",
  63534=>"100110111",
  63535=>"110000101",
  63536=>"000110010",
  63537=>"010001001",
  63538=>"110000000",
  63539=>"000011010",
  63540=>"111110001",
  63541=>"101001100",
  63542=>"101010111",
  63543=>"101100010",
  63544=>"010111111",
  63545=>"100111001",
  63546=>"011111011",
  63547=>"111101110",
  63548=>"111000010",
  63549=>"010111111",
  63550=>"100010101",
  63551=>"011100010",
  63552=>"001001111",
  63553=>"011101011",
  63554=>"100011101",
  63555=>"011001111",
  63556=>"111010111",
  63557=>"100111111",
  63558=>"101101000",
  63559=>"010011110",
  63560=>"010010001",
  63561=>"111001011",
  63562=>"001011010",
  63563=>"100010110",
  63564=>"101110000",
  63565=>"010111110",
  63566=>"111010100",
  63567=>"010010000",
  63568=>"010010001",
  63569=>"001010010",
  63570=>"111110000",
  63571=>"000001100",
  63572=>"111110001",
  63573=>"101100110",
  63574=>"110100001",
  63575=>"000101101",
  63576=>"100010010",
  63577=>"101101001",
  63578=>"100010001",
  63579=>"011000010",
  63580=>"111010101",
  63581=>"101100001",
  63582=>"110101101",
  63583=>"100000101",
  63584=>"011110100",
  63585=>"111110100",
  63586=>"111111010",
  63587=>"010100101",
  63588=>"010111010",
  63589=>"001111111",
  63590=>"110110111",
  63591=>"111111100",
  63592=>"100010100",
  63593=>"011100010",
  63594=>"010111110",
  63595=>"000000100",
  63596=>"011101111",
  63597=>"001001000",
  63598=>"100001010",
  63599=>"110000000",
  63600=>"010100101",
  63601=>"011010010",
  63602=>"010011010",
  63603=>"001101100",
  63604=>"110011101",
  63605=>"000100111",
  63606=>"000110000",
  63607=>"000000001",
  63608=>"010100011",
  63609=>"100000011",
  63610=>"111000111",
  63611=>"001000001",
  63612=>"110000101",
  63613=>"101000110",
  63614=>"001010101",
  63615=>"001100100",
  63616=>"010010101",
  63617=>"101100111",
  63618=>"110010000",
  63619=>"001111000",
  63620=>"001110111",
  63621=>"101100101",
  63622=>"010011101",
  63623=>"100010000",
  63624=>"011011011",
  63625=>"000011001",
  63626=>"010011111",
  63627=>"101001100",
  63628=>"010000110",
  63629=>"101111100",
  63630=>"110110000",
  63631=>"101001010",
  63632=>"111101001",
  63633=>"111110101",
  63634=>"100000011",
  63635=>"101110001",
  63636=>"111001011",
  63637=>"011110010",
  63638=>"011111111",
  63639=>"000111100",
  63640=>"101101100",
  63641=>"101111111",
  63642=>"100101001",
  63643=>"011001001",
  63644=>"010111000",
  63645=>"000001010",
  63646=>"100000101",
  63647=>"001011100",
  63648=>"101011100",
  63649=>"000000110",
  63650=>"001010000",
  63651=>"101110011",
  63652=>"011011001",
  63653=>"001100010",
  63654=>"110110000",
  63655=>"011010010",
  63656=>"101101010",
  63657=>"001111100",
  63658=>"011000010",
  63659=>"110010100",
  63660=>"100111001",
  63661=>"001101011",
  63662=>"001000001",
  63663=>"000010101",
  63664=>"011000111",
  63665=>"000001010",
  63666=>"010001000",
  63667=>"101110110",
  63668=>"110011101",
  63669=>"101110001",
  63670=>"111010100",
  63671=>"000110001",
  63672=>"111100011",
  63673=>"010110011",
  63674=>"100010010",
  63675=>"110011000",
  63676=>"000010011",
  63677=>"000001001",
  63678=>"111001000",
  63679=>"111111111",
  63680=>"100100001",
  63681=>"011110001",
  63682=>"010001100",
  63683=>"100100010",
  63684=>"111011110",
  63685=>"101001001",
  63686=>"100110110",
  63687=>"101101101",
  63688=>"000100010",
  63689=>"001001001",
  63690=>"010111111",
  63691=>"100100011",
  63692=>"000101100",
  63693=>"000010000",
  63694=>"011001010",
  63695=>"101000000",
  63696=>"001000011",
  63697=>"100011100",
  63698=>"101111110",
  63699=>"101001000",
  63700=>"010011011",
  63701=>"011001011",
  63702=>"000101111",
  63703=>"110101000",
  63704=>"100010100",
  63705=>"100011100",
  63706=>"010001001",
  63707=>"000101110",
  63708=>"100001101",
  63709=>"100011010",
  63710=>"000000010",
  63711=>"101000100",
  63712=>"100000000",
  63713=>"000110010",
  63714=>"011111010",
  63715=>"100000000",
  63716=>"110001010",
  63717=>"010000011",
  63718=>"001010100",
  63719=>"111001011",
  63720=>"011110001",
  63721=>"000100110",
  63722=>"000011110",
  63723=>"101011100",
  63724=>"001101000",
  63725=>"010011110",
  63726=>"001000011",
  63727=>"001010110",
  63728=>"110000001",
  63729=>"101110111",
  63730=>"110011011",
  63731=>"010000010",
  63732=>"011101001",
  63733=>"001101110",
  63734=>"000111010",
  63735=>"010111010",
  63736=>"011101110",
  63737=>"111001101",
  63738=>"001111000",
  63739=>"111011111",
  63740=>"011111001",
  63741=>"011001001",
  63742=>"100011011",
  63743=>"100110000",
  63744=>"000100010",
  63745=>"001000001",
  63746=>"001101010",
  63747=>"101100001",
  63748=>"001010010",
  63749=>"001101101",
  63750=>"100111010",
  63751=>"110111111",
  63752=>"110001001",
  63753=>"010111001",
  63754=>"000000110",
  63755=>"000101000",
  63756=>"010111000",
  63757=>"110010010",
  63758=>"011110110",
  63759=>"100100001",
  63760=>"100110001",
  63761=>"001010000",
  63762=>"001100000",
  63763=>"101001110",
  63764=>"110111110",
  63765=>"111011010",
  63766=>"010100100",
  63767=>"101110100",
  63768=>"111110110",
  63769=>"100101110",
  63770=>"011110000",
  63771=>"101100100",
  63772=>"010100111",
  63773=>"111111010",
  63774=>"001000001",
  63775=>"111010111",
  63776=>"010010100",
  63777=>"011111000",
  63778=>"100001001",
  63779=>"011100001",
  63780=>"011001010",
  63781=>"001000011",
  63782=>"010000100",
  63783=>"100010000",
  63784=>"100101111",
  63785=>"011101001",
  63786=>"010111100",
  63787=>"100111010",
  63788=>"101110010",
  63789=>"010000000",
  63790=>"100111111",
  63791=>"110111000",
  63792=>"110011011",
  63793=>"101011111",
  63794=>"001001000",
  63795=>"010000001",
  63796=>"011011111",
  63797=>"111111001",
  63798=>"101010001",
  63799=>"000011010",
  63800=>"010101011",
  63801=>"010111110",
  63802=>"000111101",
  63803=>"111011011",
  63804=>"010010010",
  63805=>"001010101",
  63806=>"100011111",
  63807=>"100000001",
  63808=>"001000011",
  63809=>"001010010",
  63810=>"001100001",
  63811=>"000000110",
  63812=>"000111110",
  63813=>"110101100",
  63814=>"010110111",
  63815=>"011111000",
  63816=>"101011011",
  63817=>"010010100",
  63818=>"100101011",
  63819=>"100010110",
  63820=>"001001010",
  63821=>"100001010",
  63822=>"110011011",
  63823=>"111111001",
  63824=>"100001101",
  63825=>"001000010",
  63826=>"001011101",
  63827=>"001000111",
  63828=>"100111000",
  63829=>"111100101",
  63830=>"010001010",
  63831=>"010011001",
  63832=>"001011101",
  63833=>"010111000",
  63834=>"010001100",
  63835=>"111010001",
  63836=>"110100101",
  63837=>"101000011",
  63838=>"011101001",
  63839=>"001001001",
  63840=>"111010100",
  63841=>"100001010",
  63842=>"000101100",
  63843=>"010000011",
  63844=>"001100011",
  63845=>"101001100",
  63846=>"111111111",
  63847=>"000010001",
  63848=>"111111010",
  63849=>"101011101",
  63850=>"110101011",
  63851=>"000111100",
  63852=>"011100001",
  63853=>"001000110",
  63854=>"110010010",
  63855=>"001010100",
  63856=>"000101100",
  63857=>"101010010",
  63858=>"100001100",
  63859=>"101011101",
  63860=>"111111000",
  63861=>"110111111",
  63862=>"010110010",
  63863=>"010000111",
  63864=>"000101100",
  63865=>"000110101",
  63866=>"011000100",
  63867=>"100100111",
  63868=>"100011100",
  63869=>"111100110",
  63870=>"011111100",
  63871=>"001100101",
  63872=>"011010111",
  63873=>"010101010",
  63874=>"101001101",
  63875=>"100100011",
  63876=>"111111001",
  63877=>"100001110",
  63878=>"100100011",
  63879=>"010111000",
  63880=>"100001100",
  63881=>"011100010",
  63882=>"011001010",
  63883=>"001101010",
  63884=>"000011001",
  63885=>"111011001",
  63886=>"001110100",
  63887=>"001100011",
  63888=>"100101110",
  63889=>"000001001",
  63890=>"011110101",
  63891=>"011101001",
  63892=>"111000100",
  63893=>"111001001",
  63894=>"000000000",
  63895=>"010011101",
  63896=>"100011100",
  63897=>"000001101",
  63898=>"110110100",
  63899=>"110010000",
  63900=>"011010000",
  63901=>"000100011",
  63902=>"111101001",
  63903=>"101011101",
  63904=>"110110011",
  63905=>"010010010",
  63906=>"010101101",
  63907=>"101011111",
  63908=>"111001110",
  63909=>"011011011",
  63910=>"110001010",
  63911=>"110110100",
  63912=>"111001110",
  63913=>"000011101",
  63914=>"000100110",
  63915=>"010111011",
  63916=>"001111110",
  63917=>"110011111",
  63918=>"001001110",
  63919=>"000001100",
  63920=>"010110000",
  63921=>"001100111",
  63922=>"011110001",
  63923=>"000011010",
  63924=>"010010011",
  63925=>"000011111",
  63926=>"111010010",
  63927=>"110101011",
  63928=>"111010110",
  63929=>"001001110",
  63930=>"001000001",
  63931=>"101101011",
  63932=>"100111111",
  63933=>"110011010",
  63934=>"100101011",
  63935=>"110101010",
  63936=>"100101101",
  63937=>"101011100",
  63938=>"001101011",
  63939=>"011110101",
  63940=>"110111111",
  63941=>"001000000",
  63942=>"111111110",
  63943=>"010110100",
  63944=>"011000010",
  63945=>"011110010",
  63946=>"110111010",
  63947=>"011010000",
  63948=>"101011100",
  63949=>"010111111",
  63950=>"010101000",
  63951=>"010100100",
  63952=>"000110001",
  63953=>"100011001",
  63954=>"001110001",
  63955=>"010001100",
  63956=>"101001111",
  63957=>"101000111",
  63958=>"011001010",
  63959=>"010011001",
  63960=>"010101111",
  63961=>"100011011",
  63962=>"001000110",
  63963=>"110101000",
  63964=>"111000010",
  63965=>"010000110",
  63966=>"000000110",
  63967=>"111101001",
  63968=>"110111111",
  63969=>"011100111",
  63970=>"000111001",
  63971=>"100001101",
  63972=>"110000010",
  63973=>"111011010",
  63974=>"111111110",
  63975=>"100000100",
  63976=>"010000010",
  63977=>"011000101",
  63978=>"100101001",
  63979=>"000110101",
  63980=>"100001110",
  63981=>"001001101",
  63982=>"100101010",
  63983=>"111011010",
  63984=>"001010100",
  63985=>"101111110",
  63986=>"101011110",
  63987=>"011110100",
  63988=>"100010110",
  63989=>"101100101",
  63990=>"010001000",
  63991=>"101101101",
  63992=>"000010001",
  63993=>"011100100",
  63994=>"110101101",
  63995=>"011110101",
  63996=>"001011101",
  63997=>"001010001",
  63998=>"010101111",
  63999=>"110101000",
  64000=>"000010100",
  64001=>"010110001",
  64002=>"010110001",
  64003=>"001010111",
  64004=>"001100101",
  64005=>"111110111",
  64006=>"101010001",
  64007=>"000010101",
  64008=>"000011000",
  64009=>"010001111",
  64010=>"111100101",
  64011=>"001000001",
  64012=>"111100001",
  64013=>"101011011",
  64014=>"000010011",
  64015=>"001111111",
  64016=>"001001011",
  64017=>"110101110",
  64018=>"010100100",
  64019=>"001000110",
  64020=>"101011101",
  64021=>"101101101",
  64022=>"000010111",
  64023=>"111001111",
  64024=>"011000101",
  64025=>"100100111",
  64026=>"101100010",
  64027=>"000111100",
  64028=>"101110101",
  64029=>"110110011",
  64030=>"100001000",
  64031=>"011111000",
  64032=>"110110110",
  64033=>"001011110",
  64034=>"000100011",
  64035=>"100010111",
  64036=>"111001101",
  64037=>"111101000",
  64038=>"100000101",
  64039=>"111110010",
  64040=>"010100101",
  64041=>"101110000",
  64042=>"011101110",
  64043=>"010001110",
  64044=>"010101100",
  64045=>"101110100",
  64046=>"000000010",
  64047=>"000011100",
  64048=>"100001110",
  64049=>"011111110",
  64050=>"101100101",
  64051=>"110111011",
  64052=>"011010001",
  64053=>"011011000",
  64054=>"001111010",
  64055=>"001101110",
  64056=>"000110111",
  64057=>"110010110",
  64058=>"001110010",
  64059=>"100011110",
  64060=>"101111111",
  64061=>"111110101",
  64062=>"110011110",
  64063=>"011011001",
  64064=>"110101001",
  64065=>"000001101",
  64066=>"101010111",
  64067=>"111101110",
  64068=>"101111100",
  64069=>"111010111",
  64070=>"001111100",
  64071=>"001010111",
  64072=>"100101100",
  64073=>"110001010",
  64074=>"110110100",
  64075=>"010111011",
  64076=>"001101111",
  64077=>"010111011",
  64078=>"111111111",
  64079=>"011110111",
  64080=>"000111001",
  64081=>"000110011",
  64082=>"100010011",
  64083=>"000100100",
  64084=>"000001000",
  64085=>"110011011",
  64086=>"100001101",
  64087=>"010000110",
  64088=>"110000011",
  64089=>"011111000",
  64090=>"110100100",
  64091=>"000011111",
  64092=>"100100001",
  64093=>"101101000",
  64094=>"001111001",
  64095=>"100110111",
  64096=>"110111100",
  64097=>"000111000",
  64098=>"011111001",
  64099=>"000111010",
  64100=>"101100010",
  64101=>"111010110",
  64102=>"010100100",
  64103=>"111110110",
  64104=>"100011101",
  64105=>"010000010",
  64106=>"111000011",
  64107=>"000101100",
  64108=>"000100100",
  64109=>"010010110",
  64110=>"000101011",
  64111=>"110100111",
  64112=>"111011101",
  64113=>"000011000",
  64114=>"111101101",
  64115=>"011100110",
  64116=>"011010111",
  64117=>"101110111",
  64118=>"011110000",
  64119=>"111000011",
  64120=>"001111101",
  64121=>"010011011",
  64122=>"000100011",
  64123=>"000001000",
  64124=>"111011101",
  64125=>"001011000",
  64126=>"110001010",
  64127=>"111000010",
  64128=>"000111010",
  64129=>"001010110",
  64130=>"100011101",
  64131=>"000001000",
  64132=>"110101100",
  64133=>"000100100",
  64134=>"000001101",
  64135=>"000110000",
  64136=>"100011111",
  64137=>"100110011",
  64138=>"110110100",
  64139=>"111100111",
  64140=>"001010011",
  64141=>"111001001",
  64142=>"111110011",
  64143=>"000000100",
  64144=>"111111110",
  64145=>"000110111",
  64146=>"010001001",
  64147=>"100100101",
  64148=>"000110110",
  64149=>"110000100",
  64150=>"000000011",
  64151=>"101010100",
  64152=>"010000010",
  64153=>"111000100",
  64154=>"110010010",
  64155=>"010110100",
  64156=>"110000110",
  64157=>"100000010",
  64158=>"110001011",
  64159=>"011100011",
  64160=>"001000100",
  64161=>"100111110",
  64162=>"001111001",
  64163=>"101001010",
  64164=>"110010100",
  64165=>"011110111",
  64166=>"111100011",
  64167=>"000000001",
  64168=>"010001010",
  64169=>"001001110",
  64170=>"011110000",
  64171=>"011001000",
  64172=>"101011011",
  64173=>"111111111",
  64174=>"010101101",
  64175=>"111110010",
  64176=>"001010111",
  64177=>"100010011",
  64178=>"001010110",
  64179=>"000000100",
  64180=>"001010100",
  64181=>"111101001",
  64182=>"110010001",
  64183=>"111111111",
  64184=>"110000110",
  64185=>"100000000",
  64186=>"100000010",
  64187=>"000001001",
  64188=>"001010111",
  64189=>"001000010",
  64190=>"000010010",
  64191=>"101100111",
  64192=>"111010010",
  64193=>"101011110",
  64194=>"110000000",
  64195=>"000000011",
  64196=>"111011010",
  64197=>"100011000",
  64198=>"111001111",
  64199=>"101000101",
  64200=>"000000110",
  64201=>"001011111",
  64202=>"101111000",
  64203=>"010000101",
  64204=>"011001111",
  64205=>"111100011",
  64206=>"010000100",
  64207=>"101110111",
  64208=>"010101001",
  64209=>"111111100",
  64210=>"111011010",
  64211=>"000101000",
  64212=>"111101111",
  64213=>"001001101",
  64214=>"100000011",
  64215=>"001111111",
  64216=>"000011101",
  64217=>"100011101",
  64218=>"011001111",
  64219=>"010011010",
  64220=>"011011010",
  64221=>"010000000",
  64222=>"000011111",
  64223=>"111111010",
  64224=>"100010110",
  64225=>"100000001",
  64226=>"111101011",
  64227=>"000001101",
  64228=>"101101000",
  64229=>"010000110",
  64230=>"100011111",
  64231=>"001000110",
  64232=>"111001000",
  64233=>"100101011",
  64234=>"001100110",
  64235=>"010110111",
  64236=>"000010110",
  64237=>"010000011",
  64238=>"011110001",
  64239=>"111011000",
  64240=>"101000000",
  64241=>"111100011",
  64242=>"100111011",
  64243=>"100010101",
  64244=>"001001101",
  64245=>"100101001",
  64246=>"011101001",
  64247=>"001000111",
  64248=>"011110001",
  64249=>"101000101",
  64250=>"100010000",
  64251=>"000001111",
  64252=>"000111101",
  64253=>"000011011",
  64254=>"111001000",
  64255=>"100100010",
  64256=>"110110110",
  64257=>"101001000",
  64258=>"000000000",
  64259=>"100111001",
  64260=>"101111100",
  64261=>"000111000",
  64262=>"010100010",
  64263=>"100000010",
  64264=>"111000001",
  64265=>"001010101",
  64266=>"000001111",
  64267=>"011110011",
  64268=>"000000001",
  64269=>"110001001",
  64270=>"010110011",
  64271=>"111111110",
  64272=>"000110010",
  64273=>"100100000",
  64274=>"111101100",
  64275=>"110010010",
  64276=>"001111010",
  64277=>"000111000",
  64278=>"000110110",
  64279=>"000010110",
  64280=>"111000111",
  64281=>"001100000",
  64282=>"100111110",
  64283=>"111110110",
  64284=>"100000011",
  64285=>"100111101",
  64286=>"000010010",
  64287=>"011100110",
  64288=>"010000010",
  64289=>"110101010",
  64290=>"111001100",
  64291=>"000001101",
  64292=>"011011111",
  64293=>"000100001",
  64294=>"001001110",
  64295=>"110010001",
  64296=>"110101011",
  64297=>"111000011",
  64298=>"100110000",
  64299=>"000010100",
  64300=>"101111101",
  64301=>"000101010",
  64302=>"000101000",
  64303=>"010010000",
  64304=>"000111000",
  64305=>"010111000",
  64306=>"000110101",
  64307=>"110111010",
  64308=>"101000111",
  64309=>"000101110",
  64310=>"001110001",
  64311=>"011001111",
  64312=>"011011000",
  64313=>"000101000",
  64314=>"111111001",
  64315=>"111000100",
  64316=>"111011010",
  64317=>"000000001",
  64318=>"100110000",
  64319=>"001011100",
  64320=>"110110001",
  64321=>"011000010",
  64322=>"010100010",
  64323=>"100000010",
  64324=>"110101100",
  64325=>"011001000",
  64326=>"011110110",
  64327=>"111011001",
  64328=>"000000000",
  64329=>"011000101",
  64330=>"000001000",
  64331=>"111100001",
  64332=>"010011101",
  64333=>"000101110",
  64334=>"110000000",
  64335=>"001101000",
  64336=>"000011101",
  64337=>"000011000",
  64338=>"000101001",
  64339=>"000111011",
  64340=>"100110100",
  64341=>"110110001",
  64342=>"100110010",
  64343=>"101100011",
  64344=>"010101101",
  64345=>"001000011",
  64346=>"101110110",
  64347=>"101001111",
  64348=>"111001000",
  64349=>"000010011",
  64350=>"001010000",
  64351=>"110111111",
  64352=>"010000000",
  64353=>"100000011",
  64354=>"101111101",
  64355=>"000110110",
  64356=>"001111100",
  64357=>"100000001",
  64358=>"100111110",
  64359=>"001111000",
  64360=>"011111110",
  64361=>"001111001",
  64362=>"000001101",
  64363=>"110000101",
  64364=>"001100001",
  64365=>"001000110",
  64366=>"111011110",
  64367=>"010000110",
  64368=>"111111100",
  64369=>"100000011",
  64370=>"101100000",
  64371=>"000101001",
  64372=>"010100010",
  64373=>"001010010",
  64374=>"100110000",
  64375=>"001001000",
  64376=>"101001011",
  64377=>"111000001",
  64378=>"100010111",
  64379=>"001010001",
  64380=>"010000011",
  64381=>"000101001",
  64382=>"000011101",
  64383=>"111011101",
  64384=>"100011111",
  64385=>"011010101",
  64386=>"001001101",
  64387=>"001010001",
  64388=>"110000001",
  64389=>"011000000",
  64390=>"101011111",
  64391=>"101010100",
  64392=>"111001001",
  64393=>"010101000",
  64394=>"100000010",
  64395=>"101001011",
  64396=>"110101000",
  64397=>"110101101",
  64398=>"000001001",
  64399=>"000010110",
  64400=>"011000111",
  64401=>"010010000",
  64402=>"101101001",
  64403=>"001000010",
  64404=>"110101101",
  64405=>"110011100",
  64406=>"101110011",
  64407=>"001110100",
  64408=>"111100111",
  64409=>"011100111",
  64410=>"011001111",
  64411=>"101000011",
  64412=>"000011000",
  64413=>"001001001",
  64414=>"001000110",
  64415=>"000110011",
  64416=>"100000001",
  64417=>"101110111",
  64418=>"001101001",
  64419=>"001101000",
  64420=>"001000001",
  64421=>"101010101",
  64422=>"110010101",
  64423=>"111100111",
  64424=>"111100001",
  64425=>"000011000",
  64426=>"101010010",
  64427=>"010001100",
  64428=>"100101000",
  64429=>"011101001",
  64430=>"101010011",
  64431=>"001000101",
  64432=>"000101111",
  64433=>"101111000",
  64434=>"101010010",
  64435=>"011111110",
  64436=>"100010000",
  64437=>"011000101",
  64438=>"111011111",
  64439=>"110100010",
  64440=>"111011110",
  64441=>"010001111",
  64442=>"001101010",
  64443=>"101011011",
  64444=>"110110010",
  64445=>"110101101",
  64446=>"001011000",
  64447=>"100110111",
  64448=>"001011101",
  64449=>"100000000",
  64450=>"100001100",
  64451=>"100100010",
  64452=>"111111000",
  64453=>"111111010",
  64454=>"111111111",
  64455=>"101101100",
  64456=>"100111110",
  64457=>"100101000",
  64458=>"111110001",
  64459=>"001011110",
  64460=>"100100010",
  64461=>"100100111",
  64462=>"100000100",
  64463=>"101110110",
  64464=>"010011100",
  64465=>"010010000",
  64466=>"100110010",
  64467=>"011111101",
  64468=>"000000100",
  64469=>"110101000",
  64470=>"000010000",
  64471=>"101101011",
  64472=>"000001100",
  64473=>"110011101",
  64474=>"001000010",
  64475=>"110101011",
  64476=>"101110010",
  64477=>"010011001",
  64478=>"001101101",
  64479=>"000001000",
  64480=>"100101010",
  64481=>"111011100",
  64482=>"100011111",
  64483=>"011011010",
  64484=>"111001110",
  64485=>"111100111",
  64486=>"000000100",
  64487=>"010010110",
  64488=>"001111011",
  64489=>"010110100",
  64490=>"101110000",
  64491=>"111100110",
  64492=>"011000000",
  64493=>"110101101",
  64494=>"010000100",
  64495=>"000011110",
  64496=>"000011010",
  64497=>"110110111",
  64498=>"010111100",
  64499=>"110100010",
  64500=>"100011110",
  64501=>"010110110",
  64502=>"010000000",
  64503=>"101000010",
  64504=>"001000110",
  64505=>"111111011",
  64506=>"001100111",
  64507=>"000001001",
  64508=>"111110110",
  64509=>"011100101",
  64510=>"010110001",
  64511=>"111001001",
  64512=>"000100100",
  64513=>"101100000",
  64514=>"000100110",
  64515=>"011001001",
  64516=>"110010101",
  64517=>"100010110",
  64518=>"001101111",
  64519=>"000001000",
  64520=>"100111010",
  64521=>"111100111",
  64522=>"100010010",
  64523=>"101011111",
  64524=>"011110010",
  64525=>"010000110",
  64526=>"010000000",
  64527=>"001011101",
  64528=>"010110111",
  64529=>"001100001",
  64530=>"110110011",
  64531=>"111000100",
  64532=>"001110111",
  64533=>"111110100",
  64534=>"110110100",
  64535=>"101001001",
  64536=>"110010001",
  64537=>"110011101",
  64538=>"111110000",
  64539=>"010000011",
  64540=>"101111100",
  64541=>"111100011",
  64542=>"001110110",
  64543=>"100110000",
  64544=>"001010110",
  64545=>"010100110",
  64546=>"110010001",
  64547=>"110010010",
  64548=>"111100110",
  64549=>"110111111",
  64550=>"101100001",
  64551=>"011101001",
  64552=>"001000101",
  64553=>"000011110",
  64554=>"111100011",
  64555=>"010110011",
  64556=>"110000101",
  64557=>"101110010",
  64558=>"100001011",
  64559=>"100000000",
  64560=>"101001011",
  64561=>"000010000",
  64562=>"110110001",
  64563=>"000010001",
  64564=>"101001000",
  64565=>"100000101",
  64566=>"111010100",
  64567=>"011100010",
  64568=>"100100111",
  64569=>"101010001",
  64570=>"010011010",
  64571=>"011010101",
  64572=>"000110000",
  64573=>"110100010",
  64574=>"011010000",
  64575=>"111011101",
  64576=>"101111011",
  64577=>"010000001",
  64578=>"100101000",
  64579=>"101000001",
  64580=>"001111011",
  64581=>"011000000",
  64582=>"001100100",
  64583=>"101100100",
  64584=>"011101010",
  64585=>"111010110",
  64586=>"011111110",
  64587=>"100001100",
  64588=>"011100100",
  64589=>"101001100",
  64590=>"111101001",
  64591=>"100011110",
  64592=>"001000001",
  64593=>"100010100",
  64594=>"000100110",
  64595=>"001011110",
  64596=>"110010110",
  64597=>"001101011",
  64598=>"101110011",
  64599=>"000001110",
  64600=>"011010110",
  64601=>"010101111",
  64602=>"001110011",
  64603=>"011010010",
  64604=>"110011010",
  64605=>"110100101",
  64606=>"101100000",
  64607=>"111010010",
  64608=>"110111011",
  64609=>"000000110",
  64610=>"001001100",
  64611=>"001001000",
  64612=>"000000000",
  64613=>"000101101",
  64614=>"001100110",
  64615=>"100000111",
  64616=>"111101001",
  64617=>"100000001",
  64618=>"010000111",
  64619=>"100110011",
  64620=>"010010001",
  64621=>"111001110",
  64622=>"111011111",
  64623=>"001111111",
  64624=>"101110000",
  64625=>"101110101",
  64626=>"101010111",
  64627=>"000100000",
  64628=>"111110110",
  64629=>"100010001",
  64630=>"100111011",
  64631=>"100011011",
  64632=>"000010111",
  64633=>"110000111",
  64634=>"000111110",
  64635=>"111001011",
  64636=>"101110110",
  64637=>"101111011",
  64638=>"011111111",
  64639=>"101111100",
  64640=>"100101010",
  64641=>"100001000",
  64642=>"110000110",
  64643=>"000101110",
  64644=>"110010001",
  64645=>"001110101",
  64646=>"000111001",
  64647=>"000010001",
  64648=>"101110111",
  64649=>"000100011",
  64650=>"001000011",
  64651=>"100100110",
  64652=>"110110111",
  64653=>"101101100",
  64654=>"100000011",
  64655=>"011101111",
  64656=>"110101011",
  64657=>"000100110",
  64658=>"000001110",
  64659=>"111011111",
  64660=>"110101011",
  64661=>"010100101",
  64662=>"011100000",
  64663=>"110110100",
  64664=>"101111011",
  64665=>"101100111",
  64666=>"001000011",
  64667=>"110101010",
  64668=>"010111101",
  64669=>"011011100",
  64670=>"011000011",
  64671=>"111011110",
  64672=>"011111111",
  64673=>"011000001",
  64674=>"000111011",
  64675=>"100111111",
  64676=>"011111011",
  64677=>"010101000",
  64678=>"011100001",
  64679=>"011111000",
  64680=>"000110110",
  64681=>"111100001",
  64682=>"000111101",
  64683=>"110010000",
  64684=>"000010100",
  64685=>"000111110",
  64686=>"111101100",
  64687=>"010101000",
  64688=>"000100011",
  64689=>"000101101",
  64690=>"110001000",
  64691=>"100010100",
  64692=>"110100001",
  64693=>"111111001",
  64694=>"010010010",
  64695=>"111111101",
  64696=>"100011010",
  64697=>"011010011",
  64698=>"000000110",
  64699=>"011001011",
  64700=>"110100011",
  64701=>"111011011",
  64702=>"011010011",
  64703=>"110010101",
  64704=>"110101111",
  64705=>"010110000",
  64706=>"110000110",
  64707=>"000110111",
  64708=>"000000001",
  64709=>"101000111",
  64710=>"100100001",
  64711=>"110000111",
  64712=>"101100001",
  64713=>"000111110",
  64714=>"000101000",
  64715=>"111010100",
  64716=>"001101111",
  64717=>"011001001",
  64718=>"000110001",
  64719=>"101101110",
  64720=>"010001010",
  64721=>"001011001",
  64722=>"010000000",
  64723=>"110100110",
  64724=>"110101000",
  64725=>"011000011",
  64726=>"110111100",
  64727=>"101001001",
  64728=>"000000000",
  64729=>"100011000",
  64730=>"000000010",
  64731=>"001110000",
  64732=>"101011011",
  64733=>"100001110",
  64734=>"101000101",
  64735=>"111110111",
  64736=>"110001000",
  64737=>"000010010",
  64738=>"011111111",
  64739=>"010100010",
  64740=>"011011000",
  64741=>"100010011",
  64742=>"111110101",
  64743=>"001010100",
  64744=>"010111010",
  64745=>"001101110",
  64746=>"001100110",
  64747=>"110000011",
  64748=>"011000100",
  64749=>"111011110",
  64750=>"100000100",
  64751=>"001101100",
  64752=>"010011111",
  64753=>"100001110",
  64754=>"101100100",
  64755=>"100100001",
  64756=>"101110000",
  64757=>"001110010",
  64758=>"010100101",
  64759=>"001100010",
  64760=>"100100100",
  64761=>"110001110",
  64762=>"110111011",
  64763=>"101100000",
  64764=>"010110110",
  64765=>"001000110",
  64766=>"110101111",
  64767=>"011001000",
  64768=>"110001010",
  64769=>"110101111",
  64770=>"001011110",
  64771=>"111011000",
  64772=>"011001011",
  64773=>"110101001",
  64774=>"100111000",
  64775=>"101000100",
  64776=>"001001111",
  64777=>"101000011",
  64778=>"001101001",
  64779=>"001110010",
  64780=>"111101101",
  64781=>"011010100",
  64782=>"011101100",
  64783=>"100001101",
  64784=>"111100100",
  64785=>"111101010",
  64786=>"100001000",
  64787=>"100111011",
  64788=>"101100110",
  64789=>"011010110",
  64790=>"101110001",
  64791=>"001011011",
  64792=>"100101011",
  64793=>"110000100",
  64794=>"000001101",
  64795=>"101010101",
  64796=>"010010010",
  64797=>"110001001",
  64798=>"001110100",
  64799=>"000000100",
  64800=>"000111000",
  64801=>"110010000",
  64802=>"100110101",
  64803=>"010010000",
  64804=>"010001110",
  64805=>"001000111",
  64806=>"101001111",
  64807=>"000010101",
  64808=>"001101110",
  64809=>"111010001",
  64810=>"101010000",
  64811=>"111001010",
  64812=>"110110111",
  64813=>"111100101",
  64814=>"100110010",
  64815=>"000111001",
  64816=>"011111100",
  64817=>"101111110",
  64818=>"101010001",
  64819=>"100000111",
  64820=>"000010110",
  64821=>"011101100",
  64822=>"111101111",
  64823=>"001111001",
  64824=>"000001100",
  64825=>"110000111",
  64826=>"111011011",
  64827=>"010100101",
  64828=>"000001001",
  64829=>"001100000",
  64830=>"111110000",
  64831=>"001010100",
  64832=>"011010100",
  64833=>"111010100",
  64834=>"011101110",
  64835=>"010011000",
  64836=>"010010000",
  64837=>"111100101",
  64838=>"001000010",
  64839=>"110110001",
  64840=>"101101010",
  64841=>"101011110",
  64842=>"011000100",
  64843=>"111000000",
  64844=>"010101010",
  64845=>"011011000",
  64846=>"011101010",
  64847=>"101000000",
  64848=>"101100110",
  64849=>"110011000",
  64850=>"111010111",
  64851=>"111010011",
  64852=>"100000111",
  64853=>"111011010",
  64854=>"110001111",
  64855=>"110011101",
  64856=>"000110001",
  64857=>"110000001",
  64858=>"000100011",
  64859=>"110110001",
  64860=>"010111010",
  64861=>"011001100",
  64862=>"101100110",
  64863=>"010011000",
  64864=>"001001110",
  64865=>"100000110",
  64866=>"010010111",
  64867=>"010011100",
  64868=>"011000110",
  64869=>"010101111",
  64870=>"000010100",
  64871=>"010100111",
  64872=>"001110111",
  64873=>"010001001",
  64874=>"101110110",
  64875=>"010110100",
  64876=>"111100100",
  64877=>"111001111",
  64878=>"011110011",
  64879=>"101101011",
  64880=>"110100001",
  64881=>"101110010",
  64882=>"001000100",
  64883=>"000001100",
  64884=>"011100001",
  64885=>"110011101",
  64886=>"011000110",
  64887=>"000101100",
  64888=>"111001111",
  64889=>"011110100",
  64890=>"111010110",
  64891=>"101101110",
  64892=>"001101011",
  64893=>"111111100",
  64894=>"100000010",
  64895=>"100100110",
  64896=>"000010000",
  64897=>"110111001",
  64898=>"111110011",
  64899=>"101111100",
  64900=>"000010110",
  64901=>"101010011",
  64902=>"011101010",
  64903=>"011101001",
  64904=>"000101010",
  64905=>"110101011",
  64906=>"011001101",
  64907=>"100110011",
  64908=>"101011011",
  64909=>"000000101",
  64910=>"001000011",
  64911=>"101111001",
  64912=>"100101011",
  64913=>"100011000",
  64914=>"110100011",
  64915=>"100101110",
  64916=>"001010010",
  64917=>"000011000",
  64918=>"010000110",
  64919=>"010101001",
  64920=>"010010100",
  64921=>"000000000",
  64922=>"111011001",
  64923=>"000101111",
  64924=>"100111101",
  64925=>"010010011",
  64926=>"101001000",
  64927=>"010110011",
  64928=>"100111001",
  64929=>"001010101",
  64930=>"111010010",
  64931=>"011001001",
  64932=>"110001101",
  64933=>"100010000",
  64934=>"100011100",
  64935=>"111110000",
  64936=>"111011001",
  64937=>"011110111",
  64938=>"001101101",
  64939=>"001000010",
  64940=>"000111100",
  64941=>"101010011",
  64942=>"101100111",
  64943=>"000101001",
  64944=>"110011100",
  64945=>"010100111",
  64946=>"110100000",
  64947=>"000000111",
  64948=>"111111110",
  64949=>"010101000",
  64950=>"000001111",
  64951=>"100010011",
  64952=>"111110111",
  64953=>"100101000",
  64954=>"001110110",
  64955=>"010100001",
  64956=>"111101100",
  64957=>"101101011",
  64958=>"000000000",
  64959=>"000111010",
  64960=>"110000010",
  64961=>"100011101",
  64962=>"000001101",
  64963=>"110111111",
  64964=>"011101010",
  64965=>"010110000",
  64966=>"110111101",
  64967=>"101000001",
  64968=>"000010010",
  64969=>"011011000",
  64970=>"110101011",
  64971=>"011110101",
  64972=>"000110111",
  64973=>"010010100",
  64974=>"000000111",
  64975=>"111100101",
  64976=>"111101111",
  64977=>"100011011",
  64978=>"110110100",
  64979=>"111111001",
  64980=>"100010100",
  64981=>"001100001",
  64982=>"010111001",
  64983=>"110000000",
  64984=>"110110111",
  64985=>"010001000",
  64986=>"001100111",
  64987=>"000011011",
  64988=>"100110011",
  64989=>"101000000",
  64990=>"001000111",
  64991=>"011110011",
  64992=>"000000000",
  64993=>"000111100",
  64994=>"100010010",
  64995=>"011111010",
  64996=>"110011010",
  64997=>"001001111",
  64998=>"110100010",
  64999=>"100000000",
  65000=>"111100111",
  65001=>"001111011",
  65002=>"011011111",
  65003=>"010111000",
  65004=>"001011001",
  65005=>"110010100",
  65006=>"110000011",
  65007=>"001010000",
  65008=>"001101110",
  65009=>"100100010",
  65010=>"000111100",
  65011=>"000000000",
  65012=>"111010000",
  65013=>"111010011",
  65014=>"001010101",
  65015=>"000000001",
  65016=>"010111111",
  65017=>"100001010",
  65018=>"000111001",
  65019=>"111001110",
  65020=>"001011010",
  65021=>"001100100",
  65022=>"101010100",
  65023=>"011001001",
  65024=>"011111111",
  65025=>"101110011",
  65026=>"110111100",
  65027=>"111010110",
  65028=>"010001000",
  65029=>"000010101",
  65030=>"001110001",
  65031=>"010100111",
  65032=>"010100011",
  65033=>"010111110",
  65034=>"010000110",
  65035=>"101011010",
  65036=>"000011101",
  65037=>"110100110",
  65038=>"111000000",
  65039=>"001011111",
  65040=>"110110001",
  65041=>"011110111",
  65042=>"001001110",
  65043=>"010011010",
  65044=>"000100001",
  65045=>"011110000",
  65046=>"100011000",
  65047=>"010010000",
  65048=>"111110111",
  65049=>"110010001",
  65050=>"100100110",
  65051=>"101010101",
  65052=>"000010001",
  65053=>"100000011",
  65054=>"111111001",
  65055=>"100100000",
  65056=>"111001001",
  65057=>"110000001",
  65058=>"011100010",
  65059=>"001110010",
  65060=>"100001101",
  65061=>"111111111",
  65062=>"111001010",
  65063=>"101111001",
  65064=>"010010000",
  65065=>"111010110",
  65066=>"111001101",
  65067=>"111110011",
  65068=>"110100111",
  65069=>"001100101",
  65070=>"101010000",
  65071=>"010001100",
  65072=>"111110001",
  65073=>"110000010",
  65074=>"100011000",
  65075=>"011011000",
  65076=>"100010100",
  65077=>"010110111",
  65078=>"111001000",
  65079=>"011110100",
  65080=>"011100111",
  65081=>"011111101",
  65082=>"001111110",
  65083=>"100110101",
  65084=>"101101000",
  65085=>"010001001",
  65086=>"011110010",
  65087=>"101101000",
  65088=>"110000001",
  65089=>"011001110",
  65090=>"010011000",
  65091=>"110111101",
  65092=>"110000010",
  65093=>"111011111",
  65094=>"101100001",
  65095=>"001000111",
  65096=>"110001111",
  65097=>"101000000",
  65098=>"111111000",
  65099=>"010010111",
  65100=>"110011110",
  65101=>"001010110",
  65102=>"110010110",
  65103=>"011111010",
  65104=>"010010000",
  65105=>"101101100",
  65106=>"010000010",
  65107=>"010110001",
  65108=>"000000010",
  65109=>"010110101",
  65110=>"000011011",
  65111=>"010001011",
  65112=>"111101011",
  65113=>"101111011",
  65114=>"101110101",
  65115=>"000000010",
  65116=>"001111000",
  65117=>"010011101",
  65118=>"011110101",
  65119=>"011011100",
  65120=>"110001101",
  65121=>"010010110",
  65122=>"000111000",
  65123=>"011010011",
  65124=>"011001001",
  65125=>"100101100",
  65126=>"111010100",
  65127=>"110001111",
  65128=>"111000011",
  65129=>"011111111",
  65130=>"011000000",
  65131=>"000110100",
  65132=>"110011000",
  65133=>"000010100",
  65134=>"001100000",
  65135=>"000100010",
  65136=>"110011101",
  65137=>"001000000",
  65138=>"111001101",
  65139=>"100100010",
  65140=>"011111001",
  65141=>"010100101",
  65142=>"011000001",
  65143=>"001110101",
  65144=>"000001000",
  65145=>"110000011",
  65146=>"010001100",
  65147=>"110111111",
  65148=>"001010101",
  65149=>"001011011",
  65150=>"011000101",
  65151=>"011101110",
  65152=>"111101001",
  65153=>"111110101",
  65154=>"100100000",
  65155=>"110001111",
  65156=>"100011101",
  65157=>"100100110",
  65158=>"101100001",
  65159=>"001111010",
  65160=>"010101011",
  65161=>"000110011",
  65162=>"000000010",
  65163=>"001100111",
  65164=>"001101011",
  65165=>"101011001",
  65166=>"111110100",
  65167=>"010110001",
  65168=>"111011001",
  65169=>"111011010",
  65170=>"001100101",
  65171=>"100011101",
  65172=>"001011011",
  65173=>"101001111",
  65174=>"110101110",
  65175=>"111000111",
  65176=>"111100000",
  65177=>"111111111",
  65178=>"010101000",
  65179=>"101110101",
  65180=>"111101001",
  65181=>"000001101",
  65182=>"110100110",
  65183=>"001110111",
  65184=>"001101110",
  65185=>"100111110",
  65186=>"001000100",
  65187=>"010110100",
  65188=>"101110111",
  65189=>"010110101",
  65190=>"010100011",
  65191=>"000110000",
  65192=>"101011101",
  65193=>"010000010",
  65194=>"110100110",
  65195=>"111111000",
  65196=>"011001000",
  65197=>"100101111",
  65198=>"011111101",
  65199=>"100010010",
  65200=>"110101101",
  65201=>"011010100",
  65202=>"100001001",
  65203=>"110111010",
  65204=>"100110100",
  65205=>"110101011",
  65206=>"100111101",
  65207=>"111101000",
  65208=>"010000100",
  65209=>"000000010",
  65210=>"101111000",
  65211=>"111011010",
  65212=>"111110000",
  65213=>"100110001",
  65214=>"110011010",
  65215=>"000011011",
  65216=>"001001101",
  65217=>"101101001",
  65218=>"100011101",
  65219=>"000000111",
  65220=>"100000100",
  65221=>"010101010",
  65222=>"110001100",
  65223=>"000000011",
  65224=>"000111001",
  65225=>"100001001",
  65226=>"010010010",
  65227=>"110100100",
  65228=>"000011000",
  65229=>"010111001",
  65230=>"011111001",
  65231=>"101111011",
  65232=>"101101010",
  65233=>"100111100",
  65234=>"011001000",
  65235=>"110100100",
  65236=>"000010101",
  65237=>"010101000",
  65238=>"000001101",
  65239=>"100001110",
  65240=>"110110111",
  65241=>"111110101",
  65242=>"111111100",
  65243=>"010001100",
  65244=>"100011101",
  65245=>"001101100",
  65246=>"000110111",
  65247=>"001101101",
  65248=>"100110000",
  65249=>"011000001",
  65250=>"001110000",
  65251=>"001001110",
  65252=>"101001110",
  65253=>"001001110",
  65254=>"100000100",
  65255=>"100011110",
  65256=>"010010110",
  65257=>"010010110",
  65258=>"001101001",
  65259=>"001010100",
  65260=>"110000000",
  65261=>"000101010",
  65262=>"001101001",
  65263=>"111000111",
  65264=>"110000110",
  65265=>"100100000",
  65266=>"010111010",
  65267=>"111101111",
  65268=>"000000001",
  65269=>"010101001",
  65270=>"100011001",
  65271=>"110100000",
  65272=>"011100111",
  65273=>"101000100",
  65274=>"100001000",
  65275=>"001000100",
  65276=>"000110101",
  65277=>"011011001",
  65278=>"011000101",
  65279=>"000101100",
  65280=>"010111011",
  65281=>"001100101",
  65282=>"001011010",
  65283=>"111110001",
  65284=>"111111110",
  65285=>"101010011",
  65286=>"101111001",
  65287=>"010100011",
  65288=>"000000111",
  65289=>"101100011",
  65290=>"010011010",
  65291=>"000001100",
  65292=>"000101101",
  65293=>"100110110",
  65294=>"101000010",
  65295=>"010111111",
  65296=>"111110101",
  65297=>"001001000",
  65298=>"000101011",
  65299=>"001000011",
  65300=>"001010000",
  65301=>"110001110",
  65302=>"010000010",
  65303=>"111000010",
  65304=>"101100100",
  65305=>"010100100",
  65306=>"000100111",
  65307=>"010000100",
  65308=>"101101111",
  65309=>"110001111",
  65310=>"110011110",
  65311=>"111011001",
  65312=>"001001011",
  65313=>"001110111",
  65314=>"100100001",
  65315=>"010000001",
  65316=>"100100100",
  65317=>"110110000",
  65318=>"111111100",
  65319=>"010101001",
  65320=>"000110110",
  65321=>"011110000",
  65322=>"101111110",
  65323=>"011100010",
  65324=>"101001111",
  65325=>"001110111",
  65326=>"000000100",
  65327=>"011110110",
  65328=>"010110101",
  65329=>"011011001",
  65330=>"010001000",
  65331=>"000101000",
  65332=>"000010110",
  65333=>"000000000",
  65334=>"001110111",
  65335=>"000111000",
  65336=>"010110101",
  65337=>"011010010",
  65338=>"101001001",
  65339=>"011100110",
  65340=>"100111111",
  65341=>"100000100",
  65342=>"010111001",
  65343=>"010010101",
  65344=>"000000001",
  65345=>"100110010",
  65346=>"000010111",
  65347=>"001100001",
  65348=>"110110010",
  65349=>"100111110",
  65350=>"111110010",
  65351=>"101010110",
  65352=>"101011001",
  65353=>"110110000",
  65354=>"111001011",
  65355=>"111101111",
  65356=>"110010011",
  65357=>"100101110",
  65358=>"110101000",
  65359=>"011111111",
  65360=>"000011011",
  65361=>"000100001",
  65362=>"110110001",
  65363=>"001101111",
  65364=>"101001000",
  65365=>"100111111",
  65366=>"101000101",
  65367=>"100010001",
  65368=>"011101011",
  65369=>"110000011",
  65370=>"011101001",
  65371=>"011110011",
  65372=>"000100000",
  65373=>"110000000",
  65374=>"001100100",
  65375=>"010110010",
  65376=>"000111010",
  65377=>"111100101",
  65378=>"111001111",
  65379=>"000111110",
  65380=>"101011111",
  65381=>"111011011",
  65382=>"111011100",
  65383=>"010100001",
  65384=>"011101000",
  65385=>"010011111",
  65386=>"000101100",
  65387=>"100111101",
  65388=>"010100101",
  65389=>"101111101",
  65390=>"111100011",
  65391=>"001011100",
  65392=>"101111000",
  65393=>"001110011",
  65394=>"010101000",
  65395=>"110110010",
  65396=>"010000000",
  65397=>"000111000",
  65398=>"110100000",
  65399=>"111111000",
  65400=>"110010011",
  65401=>"010010111",
  65402=>"010001001",
  65403=>"011100000",
  65404=>"011001010",
  65405=>"001010001",
  65406=>"010111101",
  65407=>"011111001",
  65408=>"000111000",
  65409=>"111000001",
  65410=>"000000010",
  65411=>"100100010",
  65412=>"101011101",
  65413=>"101101100",
  65414=>"101110001",
  65415=>"001101000",
  65416=>"001101110",
  65417=>"110111110",
  65418=>"111101010",
  65419=>"110011001",
  65420=>"001010110",
  65421=>"101001111",
  65422=>"101000111",
  65423=>"010111110",
  65424=>"001000010",
  65425=>"111111111",
  65426=>"101100011",
  65427=>"101101110",
  65428=>"111110000",
  65429=>"011010111",
  65430=>"110100111",
  65431=>"000000101",
  65432=>"010010000",
  65433=>"011010000",
  65434=>"000001011",
  65435=>"001010100",
  65436=>"110010111",
  65437=>"101011110",
  65438=>"101000110",
  65439=>"000001111",
  65440=>"001001100",
  65441=>"100110101",
  65442=>"010101101",
  65443=>"111100010",
  65444=>"011101101",
  65445=>"001101011",
  65446=>"000100111",
  65447=>"000101000",
  65448=>"010010010",
  65449=>"010010101",
  65450=>"111111101",
  65451=>"101111111",
  65452=>"010010100",
  65453=>"000100011",
  65454=>"010001011",
  65455=>"001000110",
  65456=>"111111001",
  65457=>"001101010",
  65458=>"000000111",
  65459=>"101111110",
  65460=>"111000010",
  65461=>"001010001",
  65462=>"111101111",
  65463=>"000000100",
  65464=>"000100110",
  65465=>"011110000",
  65466=>"101000000",
  65467=>"101111110",
  65468=>"111111111",
  65469=>"011100010",
  65470=>"010001010",
  65471=>"111000110",
  65472=>"101001000",
  65473=>"000001011",
  65474=>"111010111",
  65475=>"010000010",
  65476=>"000111000",
  65477=>"100110110",
  65478=>"001111110",
  65479=>"011010010",
  65480=>"010010110",
  65481=>"101010111",
  65482=>"100100000",
  65483=>"101101100",
  65484=>"010111010",
  65485=>"010111000",
  65486=>"110111000",
  65487=>"000110100",
  65488=>"101101000",
  65489=>"011011010",
  65490=>"011110111",
  65491=>"011010010",
  65492=>"101000110",
  65493=>"001111101",
  65494=>"100001001",
  65495=>"111100001",
  65496=>"000111101",
  65497=>"000000000",
  65498=>"101110000",
  65499=>"011100000",
  65500=>"001011000",
  65501=>"110110101",
  65502=>"010111110",
  65503=>"110001111",
  65504=>"000011000",
  65505=>"010010001",
  65506=>"001001000",
  65507=>"011101010",
  65508=>"011010100",
  65509=>"101101111",
  65510=>"100110010",
  65511=>"011111100",
  65512=>"100101010",
  65513=>"011000101",
  65514=>"110010010",
  65515=>"100010010",
  65516=>"000000001",
  65517=>"101010110",
  65518=>"110110000",
  65519=>"100011011",
  65520=>"000000110",
  65521=>"000000111",
  65522=>"100000011",
  65523=>"111011100",
  65524=>"100000011",
  65525=>"000001001",
  65526=>"100101111",
  65527=>"001101100",
  65528=>"111100000",
  65529=>"111010000",
  65530=>"101011000",
  65531=>"000010110",
  65532=>"011101011",
  65533=>"011010000",
  65534=>"010011001",
  65535=>"000101010");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;