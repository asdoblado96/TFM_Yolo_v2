LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L6_2_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(7 DOWNTO 0));
END L6_2_BNROM;

ARCHITECTURE RTL OF L6_2_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 255) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"1111010011010110"&"0001011010110000",
  1=>"1110110001010010"&"0001100011110010",
  2=>"1110111110100011"&"0001111000001101",
  3=>"1111010010001110"&"0001101011101010",
  4=>"1110111110001001"&"0010011001000100",
  5=>"1111111101000111"&"0001101101100100",
  6=>"1110111110011110"&"0010011101000000",
  7=>"1110100111011010"&"0010010001000001",
  8=>"1111011100111110"&"0001110111001100",
  9=>"1111001010101011"&"0001100001101011",
  10=>"1111101000110000"&"0001101010111000",
  11=>"1111011111000000"&"0001111001000111",
  12=>"1111100101101110"&"0001011001010001",
  13=>"1111100010100100"&"0001100110110001",
  14=>"1111000100010000"&"0010001010010010",
  15=>"1111000110101010"&"0001110100111100",
  16=>"1110111111101101"&"0001110100000000",
  17=>"1111010101100000"&"0001011011010011",
  18=>"1111110001000101"&"0001001111111100",
  19=>"1111011111011001"&"0001100011010110",
  20=>"1111011011110101"&"0001011110111110",
  21=>"1111011101100010"&"0001100101000011",
  22=>"1111110110101100"&"0001100100110010",
  23=>"1111011001000100"&"0001100111000000",
  24=>"0000010011111111"&"0001001110111101",
  25=>"1111010111011000"&"0010001001111000",
  26=>"1111101100110010"&"0001010110010101",
  27=>"1111100111100101"&"0001011011101110",
  28=>"1111110001101100"&"0001101010100011",
  29=>"1111110000101010"&"0001010111110110",
  30=>"1111100010101100"&"0001001000101001",
  31=>"0000001100110101"&"0001100000000101",
  32=>"1111000101001001"&"0001111110101110",
  33=>"1111011001100011"&"0001111100110000",
  34=>"1111010001001001"&"0001111000001101",
  35=>"1111000110001101"&"0001111110000111",
  36=>"1110110001000110"&"0010010101011010",
  37=>"1111010100101111"&"0001110101011011",
  38=>"1111011011100101"&"0001100100110111",
  39=>"1111001110110110"&"0001110101111101",
  40=>"1111011101010111"&"0001101101000110",
  41=>"0000001010100100"&"0001001000001101",
  42=>"1111001001101010"&"0001110000101011",
  43=>"0000000010110010"&"0001001011100110",
  44=>"1111100011101110"&"0001100010011010",
  45=>"1111011010011100"&"0001100110111111",
  46=>"1111000001001110"&"0001010000110100",
  47=>"1111000101110001"&"0001001011011100",
  48=>"1111110111100100"&"0001100011011101",
  49=>"1111101011111000"&"0001010100000010",
  50=>"1111101101110100"&"0001101100100011",
  51=>"1111011000011101"&"0001111000000111",
  52=>"1111011110101101"&"0001101011010111",
  53=>"1111011000100101"&"0001101000100010",
  54=>"1110111010011010"&"0001101110110100",
  55=>"1111010110010111"&"0001110000001000",
  56=>"1111011010000101"&"0001010001110111",
  57=>"1111010010001010"&"0001111001110100",
  58=>"1111100011100001"&"0001011000111011",
  59=>"1111011000000100"&"0001100010100001",
  60=>"1111100000101010"&"0001001111110100",
  61=>"1111010010001101"&"0001100110011010",
  62=>"1111110111100001"&"0001011110001011",
  63=>"1111010010111100"&"0001101010011011",
  64=>"1111100111111110"&"0001010011001101",
  65=>"1111101110001000"&"0001111100110101",
  66=>"1111110001100100"&"0001100100001110",
  67=>"1111111010010000"&"0001101010110001",
  68=>"1111010110100101"&"0001110101001001",
  69=>"1111100001101000"&"0001101001001101",
  70=>"1111010111100001"&"0001010011111000",
  71=>"1111101001000010"&"0001010000001111",
  72=>"1111011110111111"&"0001000000110000",
  73=>"1111111100111100"&"0001010111111101",
  74=>"1111100100110000"&"0010000000100110",
  75=>"1111011001110101"&"0001111100100011",
  76=>"1111101011011101"&"0001011110101101",
  77=>"1111101110010011"&"0001011010010000",
  78=>"1111001101100111"&"0001110110111000",
  79=>"1111011011100011"&"0001100000111010",
  80=>"1111001110110100"&"0001101100000101",
  81=>"1110011101110110"&"0010001101011000",
  82=>"1111101101100001"&"0001100010000001",
  83=>"1111100100111000"&"0001100101010001",
  84=>"1111110011010000"&"0001011010100110",
  85=>"1111111001100010"&"0000111110111011",
  86=>"1111100110000111"&"0001100010100101",
  87=>"1111111011100010"&"0001001111100010",
  88=>"1111111011001110"&"0001101110101000",
  89=>"1111100111011100"&"0001001011100001",
  90=>"1111101001100001"&"0001011110001011",
  91=>"1111000010010111"&"0010010111000001",
  92=>"1111100101011000"&"0001001100011000",
  93=>"1111110111010111"&"0001000010001010",
  94=>"1111100111101001"&"0001110000101010",
  95=>"1111011010111101"&"0010001100101011",
  96=>"1111001110111010"&"0001101010011011",
  97=>"1111111011000000"&"0001000100110111",
  98=>"1111011100100100"&"0001110001000000",
  99=>"1111110100010110"&"0001001101011001",
  100=>"1111111011100000"&"0001011000001101",
  101=>"1111100010101001"&"0000111010011111",
  102=>"1111100110100111"&"0001001010010110",
  103=>"1111000110101001"&"0001101111000101",
  104=>"1111100010110010"&"0010000011000010",
  105=>"1111000000100001"&"0010000111000011",
  106=>"1111110111111001"&"0001010000110101",
  107=>"1111011000100101"&"0001100010111101",
  108=>"1111101100001111"&"0001100001100000",
  109=>"1111001100011110"&"0001111101110101",
  110=>"1111010111001100"&"0001011100110011",
  111=>"1111011101110010"&"0001001001000100",
  112=>"1111001100001000"&"0001010110101001",
  113=>"1111010110000110"&"0001010000001111",
  114=>"1111100000001111"&"0001101111000001",
  115=>"1111111101111101"&"0001011111011100",
  116=>"1111010011100011"&"0001100010001101",
  117=>"1110100101011101"&"0010010001110110",
  118=>"1111011101001010"&"0001110001100010",
  119=>"1111001111101010"&"0001100101011100",
  120=>"1111101111001001"&"0001001000000000",
  121=>"1111101111011101"&"0001001111000101",
  122=>"1111111111011100"&"0001001101010001",
  123=>"1111011111100000"&"0001110111100100",
  124=>"1111010010111110"&"0001101100001111",
  125=>"1111101000111100"&"0010000100100111",
  126=>"1111001010010110"&"0001100100010011",
  127=>"1111111001011110"&"0001000101001101",
  128=>"1111001000100111"&"0001110110110111",
  129=>"1111011010101110"&"0001110101011000",
  130=>"1111101111011001"&"0001001101110000",
  131=>"1111111010000101"&"0001011000001000",
  132=>"1111110010000100"&"0001101001011011",
  133=>"1111011011101111"&"0001011010101011",
  134=>"1111011110110010"&"0001111000101111",
  135=>"1111000111101101"&"0001110100011011",
  136=>"0000001010101101"&"0001001001110111",
  137=>"1111001100110100"&"0010000110110100",
  138=>"1111100110001110"&"0001101010000001",
  139=>"1111110000000010"&"0001100110010111",
  140=>"0000011001101001"&"0001010010111100",
  141=>"1111011011110110"&"0001101010110110",
  142=>"1111011001011000"&"0001111000001100",
  143=>"1111011110000010"&"0001010111011011",
  144=>"1111101001001011"&"0000110101110001",
  145=>"1111101110101011"&"0001101001110111",
  146=>"1111110011011001"&"0001100010110001",
  147=>"1111101000011111"&"0001001011101010",
  148=>"1111111010100000"&"0001100001001110",
  149=>"1111100110111001"&"0001000110101001",
  150=>"1110101111001000"&"0010001001010011",
  151=>"1111010101101001"&"0001101010000111",
  152=>"1111111100001010"&"0001011000100100",
  153=>"1111101010000011"&"0001110100011000",
  154=>"1111001001010000"&"0010001100011111",
  155=>"1111101011001111"&"0010000011101001",
  156=>"1111011101011011"&"0001100111111110",
  157=>"1111101101011000"&"0001100110111110",
  158=>"1111100101110111"&"0001011010011111",
  159=>"1111100000010111"&"0001011101001111",
  160=>"1111100000010000"&"0001100000100011",
  161=>"1111011101110111"&"0001101011011101",
  162=>"1110011111011101"&"0010010101010110",
  163=>"1111100101001011"&"0001001110010101",
  164=>"1110001001110010"&"0010110011001000",
  165=>"1111111001101111"&"0001011011000100",
  166=>"1111110001101001"&"0001010011100101",
  167=>"1111110100101101"&"0001011001011010",
  168=>"1111010101010101"&"0001010110111111",
  169=>"1111000111111100"&"0010000001000111",
  170=>"1111101010010111"&"0001100110111101",
  171=>"1111110100111100"&"0001011111010110",
  172=>"1111011011100000"&"0001000011110100",
  173=>"1110100000100100"&"0010001000011100",
  174=>"1111001000011101"&"0001110110010110",
  175=>"1111101001010101"&"0001011101011001",
  176=>"1111011100010100"&"0001100111101000",
  177=>"0000000010100111"&"0001001110100010",
  178=>"1111010011101101"&"0001011010111011",
  179=>"1111110110010000"&"0001001010110101",
  180=>"1111100001001110"&"0001100010111100",
  181=>"1110101000101110"&"0010010110110011",
  182=>"1110100101111101"&"0011001000101110",
  183=>"1111100001011111"&"0001010101010100",
  184=>"1111010000101000"&"0001011000100101",
  185=>"1111100010000011"&"0001011010101001",
  186=>"1110110000001110"&"0001110111100010",
  187=>"1110110001001110"&"0010011101001111",
  188=>"1111111100101011"&"0001010101000001",
  189=>"1110101000101101"&"0010101101111110",
  190=>"1111011100111000"&"0001011001011100",
  191=>"1110111011111001"&"0001100000010010",
  192=>"1111100000110000"&"0001100010001010",
  193=>"0000001110100110"&"0001000101100000",
  194=>"1111111001010001"&"0000011011100001",
  195=>"1111100010111000"&"0001010001011001",
  196=>"1110011101001010"&"0010100011010101",
  197=>"1111000000111001"&"0010001110001100",
  198=>"1111001010011110"&"0001011000111011",
  199=>"1111010001111111"&"0001100100111101",
  200=>"1110111111010011"&"0001110010110001",
  201=>"1111011100011110"&"0001111000111011",
  202=>"1110110100011111"&"0001010100011010",
  203=>"1111011011000111"&"0001011001100100",
  204=>"1111010011010011"&"0001100001010111",
  205=>"1111111000111001"&"0001011011110111",
  206=>"1111010000011111"&"0001101111100000",
  207=>"1111101110001111"&"0001110111000110",
  208=>"1111011001010000"&"0001011000010001",
  209=>"1111110110111111"&"0001111011111100",
  210=>"1111011111111000"&"0001110000110110",
  211=>"1111110000110110"&"0001010011100000",
  212=>"1111100101011011"&"0001110100010111",
  213=>"1110101100100000"&"0010001101111101",
  214=>"1111001111011001"&"0001100111110101",
  215=>"1111101001101010"&"0001011010111100",
  216=>"1111000010001001"&"0001011100101111",
  217=>"1111100010010111"&"0001011010010001",
  218=>"1111100111100011"&"0001010111111001",
  219=>"1110110101000101"&"0010010001100101",
  220=>"1111011100110000"&"0001101101001100",
  221=>"1111011000100001"&"0001111000100011",
  222=>"1111100011111011"&"0001011110111100",
  223=>"1111011000000110"&"0001100011101000",
  224=>"1111100101011000"&"0001010101110101",
  225=>"1111010010000101"&"0001100111100111",
  226=>"1111100101001110"&"0001100011110001",
  227=>"1111001010111101"&"0001111110111000",
  228=>"1111111001111111"&"0001010100100111",
  229=>"1111011111110010"&"0001110000110010",
  230=>"1111000011010011"&"0001111001001101",
  231=>"1111100101001011"&"0001001010111011",
  232=>"1111010011111110"&"0001110100010011",
  233=>"1111100001001001"&"0001101110101000",
  234=>"1110110110101001"&"0010010011110010",
  235=>"1111101001000010"&"0001100100111000",
  236=>"1111010010001010"&"0001111011101101",
  237=>"1111011011011001"&"0001100000111010",
  238=>"0000001111100111"&"0001000000100110",
  239=>"1111100011100000"&"0010000000111011",
  240=>"1111010010100111"&"0001001010010001",
  241=>"1111110110011111"&"0001011100000110",
  242=>"1111010110100111"&"0001110000110111",
  243=>"1111100011100011"&"0001010000011000",
  244=>"1111110011110011"&"0001100001111000",
  245=>"1111010001100111"&"0001011111010101",
  246=>"1111100010011011"&"0001110001001011",
  247=>"1111000011100110"&"0010000010110000",
  248=>"1111000110010100"&"0001101100101111",
  249=>"1110111010110100"&"0001011010001101",
  250=>"1111110110110010"&"0001100101111111",
  251=>"0000001000111111"&"0001000110001000",
  252=>"1111100101000111"&"0001101111001100",
  253=>"1111101010100010"&"0001101100110010",
  254=>"1111011011001011"&"0001011010010111",
  255=>"1111100001000111"&"0001110001111001");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;