LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_5_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_5_BNROM;

ARCHITECTURE RTL OF L8_5_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0000111100010101"&"0001111101000101",
  1=>"0001100101011010"&"0010010101111101",
  2=>"0001110111010111"&"0010001111011001",
  3=>"0001100011100100"&"0010010001101000",
  4=>"0011010000111111"&"0001110010110010",
  5=>"0001011000001100"&"0010010001000100",
  6=>"0000110010001010"&"0010010000111100",
  7=>"0000100010000000"&"0010011000001011",
  8=>"0001000010000000"&"0010000111001011",
  9=>"0001110100010000"&"0010010100101011",
  10=>"0010011000000111"&"0010001101000110",
  11=>"0001111000001001"&"0010000110101110",
  12=>"0010111011010110"&"0010001010010000",
  13=>"0000001111110111"&"0010011000000110",
  14=>"0001000001000101"&"0001111010101101",
  15=>"0000101001111001"&"0010001100011111",
  16=>"0000011110011110"&"0010010101101011",
  17=>"0000110001111110"&"0010010111010111",
  18=>"0001111000101010"&"0010001000110010",
  19=>"0001000110101001"&"0010010010111000",
  20=>"0000111111011101"&"0010001101100111",
  21=>"0000101101100010"&"0001101011000111",
  22=>"0001111110101010"&"0010000111000111",
  23=>"0001101001010010"&"0010010000111111",
  24=>"0010001000110010"&"0010010010111100",
  25=>"1111000000110010"&"0001101001100010",
  26=>"0000001010011010"&"0001100111100000",
  27=>"0010000110010010"&"0001111010011000",
  28=>"0000100000011000"&"0010000110000110",
  29=>"1111110001111010"&"0001111100011000",
  30=>"0001011001110111"&"0010001110010010",
  31=>"0001101010011101"&"0010001111010000",
  32=>"0000110101110010"&"0001111000001001",
  33=>"0011000011100111"&"0010011000011111",
  34=>"0010010111110101"&"0001110010111010",
  35=>"1111110000011110"&"0001110110000101",
  36=>"0000111101011110"&"0010010101000001",
  37=>"0010111111000101"&"0010001110010111",
  38=>"0001001011011011"&"0001111111011100",
  39=>"0001001101010000"&"0001110110101111",
  40=>"0001100001000000"&"0010001000001001",
  41=>"0001011101110000"&"0010000010101101",
  42=>"0000100111110111"&"0010001100000100",
  43=>"0001110010100001"&"0010010101010000",
  44=>"0000111111011011"&"0010010110001001",
  45=>"0010001011111010"&"0001101011001101",
  46=>"1110111100001011"&"0001111110111010",
  47=>"1111101010011001"&"0010001101100110",
  48=>"0011000001101000"&"0010000111110001",
  49=>"0001110100100111"&"0001111001011000",
  50=>"1111110010011101"&"0010000011011010",
  51=>"0001010110100101"&"0010010101101011",
  52=>"0001011111010111"&"0010010011000111",
  53=>"1111010010111010"&"0001110100001000",
  54=>"0000111101111100"&"0010010011001001",
  55=>"0001111011111111"&"0010000111111011",
  56=>"0001001101001110"&"0010010110011110",
  57=>"1111111010110100"&"0010011011111010",
  58=>"0000000100001110"&"0001010100100100",
  59=>"0001101110011101"&"0010000011001100",
  60=>"0000100000110001"&"0001111111000010",
  61=>"0000101001010100"&"0010011011011001",
  62=>"0000001011010011"&"0010011110111111",
  63=>"0001111110001110"&"0001111100111101");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;