LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L9_1_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(9)-1 DOWNTO 0));
END L9_1_WROM;

ARCHITECTURE RTL OF L9_1_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 64511) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"00000000",
  1=>"00000010",
  2=>"00000011",
  3=>"11111111",
  4=>"00000010",
  5=>"11111111",
  6=>"11111110",
  7=>"00000000",
  8=>"11111111",
  9=>"11111111",
  10=>"00000010",
  11=>"11111111",
  12=>"11111111",
  13=>"00000000",
  14=>"11111111",
  15=>"11111111",
  16=>"00000010",
  17=>"00000001",
  18=>"00000000",
  19=>"11111111",
  20=>"00000000",
  21=>"00000000",
  22=>"11111111",
  23=>"11111111",
  24=>"00000000",
  25=>"11111110",
  26=>"00000001",
  27=>"11111111",
  28=>"00000000",
  29=>"00000000",
  30=>"00000001",
  31=>"00000001",
  32=>"00000001",
  33=>"00000000",
  34=>"00000001",
  35=>"11111110",
  36=>"00000010",
  37=>"00000010",
  38=>"00000000",
  39=>"00000010",
  40=>"11111111",
  41=>"00000000",
  42=>"00000001",
  43=>"11111111",
  44=>"11111110",
  45=>"11111110",
  46=>"00000000",
  47=>"11111110",
  48=>"11111110",
  49=>"00000010",
  50=>"00000000",
  51=>"00000000",
  52=>"00000000",
  53=>"00000000",
  54=>"00000001",
  55=>"11111111",
  56=>"00000000",
  57=>"00000001",
  58=>"11111111",
  59=>"00000010",
  60=>"11111110",
  61=>"00000011",
  62=>"00000010",
  63=>"00000000",
  64=>"00000000",
  65=>"00000001",
  66=>"00000010",
  67=>"00000000",
  68=>"00000001",
  69=>"11111111",
  70=>"00000000",
  71=>"00000000",
  72=>"00000010",
  73=>"00000000",
  74=>"00000010",
  75=>"00000010",
  76=>"00000000",
  77=>"00000000",
  78=>"00000010",
  79=>"00000001",
  80=>"11111111",
  81=>"11111110",
  82=>"11111110",
  83=>"00000001",
  84=>"00000010",
  85=>"11111110",
  86=>"00000001",
  87=>"11111111",
  88=>"00000000",
  89=>"11111111",
  90=>"00000000",
  91=>"00000001",
  92=>"11111110",
  93=>"11111110",
  94=>"11111111",
  95=>"00000000",
  96=>"00000001",
  97=>"11111111",
  98=>"11111111",
  99=>"11111111",
  100=>"00000001",
  101=>"00000000",
  102=>"11111111",
  103=>"00000001",
  104=>"00000000",
  105=>"00000001",
  106=>"00000001",
  107=>"11111111",
  108=>"11111111",
  109=>"00000001",
  110=>"00000010",
  111=>"00000001",
  112=>"00000010",
  113=>"00000010",
  114=>"00000000",
  115=>"00000001",
  116=>"00000010",
  117=>"11111111",
  118=>"11111111",
  119=>"00000001",
  120=>"00000001",
  121=>"00000001",
  122=>"11111111",
  123=>"00000001",
  124=>"00000010",
  125=>"00000010",
  126=>"11111111",
  127=>"00000001",
  128=>"00000000",
  129=>"11111111",
  130=>"11111111",
  131=>"11111110",
  132=>"00000010",
  133=>"11111111",
  134=>"00000001",
  135=>"11111111",
  136=>"11111110",
  137=>"11111111",
  138=>"00000000",
  139=>"00000000",
  140=>"11111111",
  141=>"11111111",
  142=>"11111110",
  143=>"00000001",
  144=>"11111110",
  145=>"00000000",
  146=>"00000000",
  147=>"11111111",
  148=>"00000001",
  149=>"00000001",
  150=>"00000001",
  151=>"00000000",
  152=>"00000000",
  153=>"11111110",
  154=>"11111111",
  155=>"11111111",
  156=>"11111110",
  157=>"11111111",
  158=>"11111110",
  159=>"00000000",
  160=>"00000001",
  161=>"11111111",
  162=>"00000000",
  163=>"00000000",
  164=>"11111111",
  165=>"11111111",
  166=>"00000010",
  167=>"11111111",
  168=>"00000000",
  169=>"11111111",
  170=>"00000010",
  171=>"00000001",
  172=>"00000000",
  173=>"00000011",
  174=>"00000000",
  175=>"00000011",
  176=>"00000000",
  177=>"11111110",
  178=>"11111110",
  179=>"00000000",
  180=>"00000010",
  181=>"00000001",
  182=>"11111101",
  183=>"00000000",
  184=>"00000010",
  185=>"00000000",
  186=>"00000010",
  187=>"00000010",
  188=>"00000001",
  189=>"00000001",
  190=>"11111111",
  191=>"00000001",
  192=>"00000010",
  193=>"00000001",
  194=>"11111111",
  195=>"11111111",
  196=>"11111111",
  197=>"11111110",
  198=>"00000001",
  199=>"00000000",
  200=>"11111111",
  201=>"00000000",
  202=>"00000000",
  203=>"11111110",
  204=>"11111111",
  205=>"00000010",
  206=>"11111110",
  207=>"00000010",
  208=>"11111111",
  209=>"11111111",
  210=>"00000000",
  211=>"11111111",
  212=>"11111110",
  213=>"11111111",
  214=>"00000001",
  215=>"11111110",
  216=>"00000001",
  217=>"00000000",
  218=>"11111110",
  219=>"00000000",
  220=>"11111110",
  221=>"11111111",
  222=>"11111110",
  223=>"11111110",
  224=>"11111111",
  225=>"11111110",
  226=>"11111111",
  227=>"11111111",
  228=>"11111111",
  229=>"00000010",
  230=>"00000010",
  231=>"00000000",
  232=>"00000001",
  233=>"00000000",
  234=>"00000010",
  235=>"11111101",
  236=>"11111111",
  237=>"11111110",
  238=>"00000010",
  239=>"00000000",
  240=>"00000001",
  241=>"11111111",
  242=>"00000001",
  243=>"00000001",
  244=>"00000001",
  245=>"11111111",
  246=>"00000010",
  247=>"11111111",
  248=>"00000001",
  249=>"00000010",
  250=>"00000010",
  251=>"00000010",
  252=>"11111111",
  253=>"00000010",
  254=>"00000010",
  255=>"00000000",
  256=>"00000010",
  257=>"11111111",
  258=>"00000001",
  259=>"11111110",
  260=>"11111110",
  261=>"00000001",
  262=>"00000001",
  263=>"00000001",
  264=>"11111110",
  265=>"00000000",
  266=>"00000000",
  267=>"00000000",
  268=>"00000001",
  269=>"00000001",
  270=>"11111110",
  271=>"11111111",
  272=>"11111111",
  273=>"00000001",
  274=>"00000001",
  275=>"00000001",
  276=>"11111110",
  277=>"11111111",
  278=>"11111111",
  279=>"00000010",
  280=>"11111111",
  281=>"00000010",
  282=>"00000001",
  283=>"11111111",
  284=>"00000000",
  285=>"00000000",
  286=>"00000010",
  287=>"00000000",
  288=>"00000001",
  289=>"00000001",
  290=>"00000001",
  291=>"00000010",
  292=>"00000000",
  293=>"11111111",
  294=>"00000001",
  295=>"00000001",
  296=>"00000011",
  297=>"11111111",
  298=>"00000010",
  299=>"00000000",
  300=>"11111111",
  301=>"00000010",
  302=>"00000001",
  303=>"11111110",
  304=>"00000000",
  305=>"11111111",
  306=>"00000001",
  307=>"00000001",
  308=>"00000001",
  309=>"00000010",
  310=>"11111110",
  311=>"00000010",
  312=>"00000001",
  313=>"11111111",
  314=>"00000000",
  315=>"00000000",
  316=>"00000001",
  317=>"00000000",
  318=>"11111110",
  319=>"00000000",
  320=>"11111110",
  321=>"00000001",
  322=>"00000000",
  323=>"00000001",
  324=>"11111110",
  325=>"11111111",
  326=>"00000010",
  327=>"11111110",
  328=>"00000001",
  329=>"00000010",
  330=>"00000000",
  331=>"00000001",
  332=>"00000010",
  333=>"00000000",
  334=>"00000010",
  335=>"11111111",
  336=>"00000010",
  337=>"00000010",
  338=>"11111111",
  339=>"00000001",
  340=>"00000001",
  341=>"00000001",
  342=>"00000000",
  343=>"00000001",
  344=>"11111110",
  345=>"11111110",
  346=>"11111110",
  347=>"00000000",
  348=>"00000000",
  349=>"11111110",
  350=>"11111111",
  351=>"00000000",
  352=>"00000001",
  353=>"00000001",
  354=>"00000010",
  355=>"11111101",
  356=>"00000001",
  357=>"00000010",
  358=>"11111111",
  359=>"00000000",
  360=>"00000001",
  361=>"00000001",
  362=>"11111110",
  363=>"00000001",
  364=>"00000000",
  365=>"11111110",
  366=>"11111110",
  367=>"11111111",
  368=>"00000001",
  369=>"11111111",
  370=>"00000010",
  371=>"00000000",
  372=>"11111111",
  373=>"00000001",
  374=>"00000011",
  375=>"11111110",
  376=>"00000000",
  377=>"11111111",
  378=>"00000010",
  379=>"11111110",
  380=>"11111110",
  381=>"11111111",
  382=>"00000000",
  383=>"11111111",
  384=>"00000001",
  385=>"00000001",
  386=>"11111110",
  387=>"00000001",
  388=>"11111110",
  389=>"00000000",
  390=>"11111111",
  391=>"00000001",
  392=>"11111111",
  393=>"00000000",
  394=>"11111111",
  395=>"11111111",
  396=>"00000001",
  397=>"00000000",
  398=>"00000001",
  399=>"00000000",
  400=>"00000001",
  401=>"00000001",
  402=>"00000010",
  403=>"00000001",
  404=>"11111111",
  405=>"00000001",
  406=>"00000010",
  407=>"00000011",
  408=>"00000001",
  409=>"00000001",
  410=>"00000010",
  411=>"11111110",
  412=>"00000010",
  413=>"00000000",
  414=>"11111101",
  415=>"00000001",
  416=>"00000001",
  417=>"11111111",
  418=>"00000001",
  419=>"11111110",
  420=>"00000000",
  421=>"11111110",
  422=>"11111110",
  423=>"00000001",
  424=>"00000000",
  425=>"00000000",
  426=>"11111110",
  427=>"11111111",
  428=>"11111101",
  429=>"00000001",
  430=>"00000000",
  431=>"00000010",
  432=>"00000000",
  433=>"11111111",
  434=>"00000000",
  435=>"00000010",
  436=>"11111110",
  437=>"00000001",
  438=>"00000001",
  439=>"00000010",
  440=>"11111111",
  441=>"00000010",
  442=>"11111111",
  443=>"11111110",
  444=>"11111111",
  445=>"11111110",
  446=>"11111110",
  447=>"11111111",
  448=>"00000001",
  449=>"00000001",
  450=>"00000000",
  451=>"11111110",
  452=>"00000001",
  453=>"00000001",
  454=>"00000001",
  455=>"00000000",
  456=>"11111111",
  457=>"00000010",
  458=>"00000001",
  459=>"11111111",
  460=>"00000001",
  461=>"11111110",
  462=>"11111110",
  463=>"00000001",
  464=>"00000000",
  465=>"00000001",
  466=>"00000000",
  467=>"00000000",
  468=>"11111111",
  469=>"00000000",
  470=>"00000000",
  471=>"00000000",
  472=>"00000000",
  473=>"00000000",
  474=>"00000001",
  475=>"00000000",
  476=>"00000010",
  477=>"00000001",
  478=>"11111110",
  479=>"11111111",
  480=>"00000000",
  481=>"00000000",
  482=>"00000000",
  483=>"00000000",
  484=>"11111111",
  485=>"11111111",
  486=>"00000010",
  487=>"11111111",
  488=>"11111111",
  489=>"11111111",
  490=>"00000001",
  491=>"11111111",
  492=>"11111111",
  493=>"11111111",
  494=>"00000010",
  495=>"00000001",
  496=>"11111110",
  497=>"00000000",
  498=>"11111110",
  499=>"00000000",
  500=>"11111110",
  501=>"00000001",
  502=>"00000010",
  503=>"00000000",
  504=>"00000000",
  505=>"00000001",
  506=>"11111110",
  507=>"11111111",
  508=>"00000001",
  509=>"11111110",
  510=>"00000000",
  511=>"00000000",
  512=>"00000001",
  513=>"00000001",
  514=>"00000010",
  515=>"00000001",
  516=>"11111111",
  517=>"00000001",
  518=>"11111111",
  519=>"00000000",
  520=>"11111110",
  521=>"00000010",
  522=>"00000010",
  523=>"00000000",
  524=>"11111111",
  525=>"00000001",
  526=>"11111111",
  527=>"00000000",
  528=>"11111111",
  529=>"11111111",
  530=>"00000001",
  531=>"00000000",
  532=>"11111111",
  533=>"00000001",
  534=>"00000001",
  535=>"11111111",
  536=>"00000000",
  537=>"00000001",
  538=>"11111111",
  539=>"11111111",
  540=>"00000010",
  541=>"00000000",
  542=>"00000001",
  543=>"00000000",
  544=>"00000001",
  545=>"00000001",
  546=>"11111111",
  547=>"00000010",
  548=>"00000001",
  549=>"00000001",
  550=>"00000001",
  551=>"00000000",
  552=>"11111111",
  553=>"00000000",
  554=>"11111110",
  555=>"00000001",
  556=>"11111111",
  557=>"11111111",
  558=>"11111111",
  559=>"00000000",
  560=>"00000001",
  561=>"11111110",
  562=>"00000001",
  563=>"00000010",
  564=>"00000001",
  565=>"11111111",
  566=>"00000010",
  567=>"00000000",
  568=>"11111111",
  569=>"00000000",
  570=>"00000001",
  571=>"11111111",
  572=>"00000010",
  573=>"00000000",
  574=>"00000010",
  575=>"00000001",
  576=>"00000000",
  577=>"00000000",
  578=>"00000000",
  579=>"00000010",
  580=>"11111110",
  581=>"11111111",
  582=>"00000000",
  583=>"00000000",
  584=>"00000001",
  585=>"00000001",
  586=>"11111111",
  587=>"00000010",
  588=>"11111111",
  589=>"00000000",
  590=>"11111111",
  591=>"00000010",
  592=>"00000000",
  593=>"11111111",
  594=>"00000001",
  595=>"11111111",
  596=>"00000001",
  597=>"00000001",
  598=>"00000000",
  599=>"00000001",
  600=>"00000001",
  601=>"00000000",
  602=>"11111111",
  603=>"00000010",
  604=>"00000010",
  605=>"11111111",
  606=>"00000000",
  607=>"11111110",
  608=>"00000001",
  609=>"11111110",
  610=>"00000011",
  611=>"00000001",
  612=>"11111111",
  613=>"00000000",
  614=>"11111111",
  615=>"11111110",
  616=>"11111111",
  617=>"00000001",
  618=>"11111111",
  619=>"11111111",
  620=>"11111110",
  621=>"00000000",
  622=>"11111111",
  623=>"00000000",
  624=>"00000010",
  625=>"00000001",
  626=>"00000001",
  627=>"11111111",
  628=>"00000000",
  629=>"11111111",
  630=>"11111111",
  631=>"00000000",
  632=>"00000001",
  633=>"00000001",
  634=>"11111111",
  635=>"00000000",
  636=>"00000000",
  637=>"00000001",
  638=>"00000000",
  639=>"11111111",
  640=>"00000010",
  641=>"00000000",
  642=>"00000011",
  643=>"00000000",
  644=>"00000001",
  645=>"11111111",
  646=>"00000000",
  647=>"11111110",
  648=>"00000001",
  649=>"00000000",
  650=>"00000001",
  651=>"00000010",
  652=>"00000001",
  653=>"00000001",
  654=>"11111111",
  655=>"00000000",
  656=>"00000001",
  657=>"11111110",
  658=>"00000001",
  659=>"11111110",
  660=>"00000000",
  661=>"00000010",
  662=>"00000000",
  663=>"00000011",
  664=>"11111111",
  665=>"00000001",
  666=>"00000000",
  667=>"11111111",
  668=>"11111111",
  669=>"00000011",
  670=>"00000000",
  671=>"00000000",
  672=>"00000000",
  673=>"11111111",
  674=>"00000001",
  675=>"00000000",
  676=>"00000001",
  677=>"00000010",
  678=>"00000000",
  679=>"00000000",
  680=>"11111111",
  681=>"11111110",
  682=>"11111111",
  683=>"11111110",
  684=>"00000001",
  685=>"00000001",
  686=>"00000000",
  687=>"00000001",
  688=>"00000001",
  689=>"11111111",
  690=>"00000001",
  691=>"11111110",
  692=>"11111110",
  693=>"11111111",
  694=>"11111110",
  695=>"00000000",
  696=>"11111110",
  697=>"00000000",
  698=>"00000010",
  699=>"00000001",
  700=>"00000000",
  701=>"11111111",
  702=>"00000001",
  703=>"11111110",
  704=>"00000000",
  705=>"00000000",
  706=>"00000000",
  707=>"11111110",
  708=>"00000000",
  709=>"11111111",
  710=>"00000010",
  711=>"00000010",
  712=>"11111111",
  713=>"11111111",
  714=>"00000001",
  715=>"00000000",
  716=>"11111111",
  717=>"00000000",
  718=>"00000010",
  719=>"00000010",
  720=>"00000000",
  721=>"00000010",
  722=>"11111101",
  723=>"00000000",
  724=>"11111110",
  725=>"11111110",
  726=>"11111111",
  727=>"11111111",
  728=>"00000001",
  729=>"11111110",
  730=>"00000001",
  731=>"11111111",
  732=>"00000000",
  733=>"00000000",
  734=>"11111111",
  735=>"11111110",
  736=>"11111111",
  737=>"00000001",
  738=>"00000000",
  739=>"00000001",
  740=>"11111110",
  741=>"11111111",
  742=>"11111111",
  743=>"11111111",
  744=>"00000001",
  745=>"11111110",
  746=>"00000001",
  747=>"00000001",
  748=>"00000000",
  749=>"00000001",
  750=>"00000000",
  751=>"00000001",
  752=>"00000000",
  753=>"00000001",
  754=>"00000000",
  755=>"00000000",
  756=>"00000001",
  757=>"00000010",
  758=>"00000001",
  759=>"00000000",
  760=>"11111110",
  761=>"11111111",
  762=>"00000010",
  763=>"00000000",
  764=>"00000001",
  765=>"11111111",
  766=>"00000000",
  767=>"00000010",
  768=>"11111110",
  769=>"00000001",
  770=>"11111111",
  771=>"11111110",
  772=>"11111111",
  773=>"00000010",
  774=>"00000001",
  775=>"00000001",
  776=>"11111110",
  777=>"11111111",
  778=>"11111111",
  779=>"00000000",
  780=>"00000010",
  781=>"00000010",
  782=>"00000000",
  783=>"11111111",
  784=>"00000000",
  785=>"11111110",
  786=>"00000010",
  787=>"11111111",
  788=>"11111110",
  789=>"11111111",
  790=>"00000010",
  791=>"11111110",
  792=>"00000010",
  793=>"00000001",
  794=>"00000000",
  795=>"00000000",
  796=>"11111111",
  797=>"11111111",
  798=>"00000000",
  799=>"11111111",
  800=>"00000010",
  801=>"11111111",
  802=>"00000000",
  803=>"00000010",
  804=>"00000010",
  805=>"00000010",
  806=>"00000000",
  807=>"11111111",
  808=>"11111111",
  809=>"00000001",
  810=>"00000000",
  811=>"11111110",
  812=>"00000010",
  813=>"11111110",
  814=>"11111111",
  815=>"00000000",
  816=>"11111111",
  817=>"11111110",
  818=>"00000001",
  819=>"11111111",
  820=>"00000000",
  821=>"00000001",
  822=>"00000000",
  823=>"11111111",
  824=>"00000000",
  825=>"11111110",
  826=>"00000001",
  827=>"00000001",
  828=>"11111110",
  829=>"00000000",
  830=>"00000001",
  831=>"00000001",
  832=>"00000000",
  833=>"11111111",
  834=>"00000001",
  835=>"00000000",
  836=>"11111111",
  837=>"00000000",
  838=>"00000000",
  839=>"00000000",
  840=>"11111111",
  841=>"11111110",
  842=>"11111111",
  843=>"00000000",
  844=>"11111111",
  845=>"00000010",
  846=>"00000001",
  847=>"00000000",
  848=>"11111110",
  849=>"00000001",
  850=>"00000000",
  851=>"00000000",
  852=>"00000000",
  853=>"11111110",
  854=>"00000010",
  855=>"11111111",
  856=>"11111111",
  857=>"00000001",
  858=>"00000000",
  859=>"11111110",
  860=>"11111111",
  861=>"00000000",
  862=>"11111111",
  863=>"00000001",
  864=>"00000001",
  865=>"00000011",
  866=>"11111111",
  867=>"00000001",
  868=>"11111111",
  869=>"00000001",
  870=>"00000000",
  871=>"00000010",
  872=>"00000010",
  873=>"00000001",
  874=>"11111110",
  875=>"11111110",
  876=>"00000000",
  877=>"00000001",
  878=>"00000000",
  879=>"00000001",
  880=>"00000000",
  881=>"11111110",
  882=>"11111111",
  883=>"11111111",
  884=>"11111110",
  885=>"11111111",
  886=>"11111111",
  887=>"11111111",
  888=>"11111110",
  889=>"00000001",
  890=>"00000000",
  891=>"00000000",
  892=>"11111110",
  893=>"00000001",
  894=>"00000000",
  895=>"00000001",
  896=>"00000000",
  897=>"00000001",
  898=>"00000000",
  899=>"00000001",
  900=>"00000000",
  901=>"00000010",
  902=>"00000000",
  903=>"00000000",
  904=>"00000000",
  905=>"00000000",
  906=>"00000001",
  907=>"11111111",
  908=>"00000001",
  909=>"11111110",
  910=>"11111111",
  911=>"00000000",
  912=>"11111111",
  913=>"00000000",
  914=>"00000000",
  915=>"11111111",
  916=>"00000010",
  917=>"00000001",
  918=>"00000001",
  919=>"11111111",
  920=>"11111111",
  921=>"11111110",
  922=>"00000001",
  923=>"00000000",
  924=>"00000000",
  925=>"11111110",
  926=>"11111111",
  927=>"11111110",
  928=>"00000001",
  929=>"00000001",
  930=>"11111110",
  931=>"00000000",
  932=>"00000001",
  933=>"00000001",
  934=>"11111101",
  935=>"11111110",
  936=>"00000000",
  937=>"00000001",
  938=>"11111111",
  939=>"11111111",
  940=>"00000001",
  941=>"00000000",
  942=>"00000001",
  943=>"00000001",
  944=>"11111110",
  945=>"11111111",
  946=>"11111110",
  947=>"00000001",
  948=>"00000001",
  949=>"00000000",
  950=>"11111110",
  951=>"00000011",
  952=>"00000000",
  953=>"00000001",
  954=>"11111111",
  955=>"00000001",
  956=>"00000001",
  957=>"00000000",
  958=>"00000000",
  959=>"00000000",
  960=>"11111110",
  961=>"00000001",
  962=>"11111110",
  963=>"00000001",
  964=>"11111111",
  965=>"11111110",
  966=>"00000001",
  967=>"00000001",
  968=>"00000001",
  969=>"11111110",
  970=>"11111110",
  971=>"00000001",
  972=>"00000000",
  973=>"00000001",
  974=>"00000000",
  975=>"00000000",
  976=>"00000010",
  977=>"00000000",
  978=>"00000001",
  979=>"00000010",
  980=>"00000011",
  981=>"00000001",
  982=>"00000000",
  983=>"00000000",
  984=>"00000000",
  985=>"00000010",
  986=>"00000001",
  987=>"11111111",
  988=>"00000000",
  989=>"11111111",
  990=>"00000010",
  991=>"00000000",
  992=>"00000001",
  993=>"11111110",
  994=>"11111111",
  995=>"00000010",
  996=>"11111110",
  997=>"00000010",
  998=>"00000000",
  999=>"00000010",
  1000=>"11111111",
  1001=>"00000001",
  1002=>"11111111",
  1003=>"00000010",
  1004=>"00000000",
  1005=>"00000001",
  1006=>"00000000",
  1007=>"00000000",
  1008=>"11111110",
  1009=>"11111110",
  1010=>"11111110",
  1011=>"11111110",
  1012=>"00000000",
  1013=>"00000001",
  1014=>"00000001",
  1015=>"11111111",
  1016=>"00000001",
  1017=>"00000000",
  1018=>"00000000",
  1019=>"00000011",
  1020=>"00000001",
  1021=>"00000000",
  1022=>"00000001",
  1023=>"00000000",
  1024=>"00000001",
  1025=>"00000001",
  1026=>"11111111",
  1027=>"00000000",
  1028=>"00000001",
  1029=>"00000010",
  1030=>"00000000",
  1031=>"00000001",
  1032=>"00000001",
  1033=>"00000011",
  1034=>"00000001",
  1035=>"11111110",
  1036=>"00000001",
  1037=>"11111110",
  1038=>"00000000",
  1039=>"00000001",
  1040=>"11111110",
  1041=>"00000001",
  1042=>"00000000",
  1043=>"00000001",
  1044=>"11111111",
  1045=>"11111111",
  1046=>"11111110",
  1047=>"00000001",
  1048=>"00000001",
  1049=>"00000000",
  1050=>"00000001",
  1051=>"00000001",
  1052=>"11111110",
  1053=>"11111111",
  1054=>"00000001",
  1055=>"00000001",
  1056=>"11111101",
  1057=>"11111111",
  1058=>"11111110",
  1059=>"00000010",
  1060=>"00000011",
  1061=>"00000011",
  1062=>"00000000",
  1063=>"00000000",
  1064=>"00000010",
  1065=>"11111111",
  1066=>"00000001",
  1067=>"00000000",
  1068=>"11111111",
  1069=>"11111110",
  1070=>"11111110",
  1071=>"11111110",
  1072=>"00000010",
  1073=>"00000010",
  1074=>"11111111",
  1075=>"11111110",
  1076=>"11111101",
  1077=>"11111110",
  1078=>"00000001",
  1079=>"00000011",
  1080=>"00000000",
  1081=>"00000000",
  1082=>"00000000",
  1083=>"00000010",
  1084=>"00000001",
  1085=>"11111111",
  1086=>"00000000",
  1087=>"00000001",
  1088=>"00000000",
  1089=>"00000001",
  1090=>"00000000",
  1091=>"00000000",
  1092=>"00000000",
  1093=>"11111101",
  1094=>"00000010",
  1095=>"00000000",
  1096=>"11111101",
  1097=>"00000001",
  1098=>"00000010",
  1099=>"11111110",
  1100=>"00000010",
  1101=>"11111110",
  1102=>"00000000",
  1103=>"00000010",
  1104=>"00000011",
  1105=>"00000000",
  1106=>"00000001",
  1107=>"11111111",
  1108=>"00000001",
  1109=>"00000001",
  1110=>"11111110",
  1111=>"00000000",
  1112=>"11111110",
  1113=>"00000000",
  1114=>"11111110",
  1115=>"00000001",
  1116=>"00000001",
  1117=>"00000000",
  1118=>"00000000",
  1119=>"11111111",
  1120=>"11111111",
  1121=>"11111110",
  1122=>"00000001",
  1123=>"00000001",
  1124=>"11111110",
  1125=>"00000001",
  1126=>"00000000",
  1127=>"11111111",
  1128=>"00000000",
  1129=>"11111111",
  1130=>"00000000",
  1131=>"11111111",
  1132=>"00000000",
  1133=>"11111111",
  1134=>"11111111",
  1135=>"00000000",
  1136=>"00000000",
  1137=>"11111111",
  1138=>"00000000",
  1139=>"11111110",
  1140=>"11111111",
  1141=>"00000001",
  1142=>"00000000",
  1143=>"00000001",
  1144=>"11111111",
  1145=>"00000001",
  1146=>"00000001",
  1147=>"11111110",
  1148=>"11111110",
  1149=>"11111111",
  1150=>"00000001",
  1151=>"11111110",
  1152=>"11111111",
  1153=>"11111111",
  1154=>"11111110",
  1155=>"11111110",
  1156=>"11111110",
  1157=>"11111111",
  1158=>"00000000",
  1159=>"00000001",
  1160=>"00000000",
  1161=>"00000010",
  1162=>"11111110",
  1163=>"11111110",
  1164=>"11111110",
  1165=>"11111110",
  1166=>"00000001",
  1167=>"00000000",
  1168=>"11111111",
  1169=>"11111110",
  1170=>"00000010",
  1171=>"11111111",
  1172=>"00000010",
  1173=>"11111111",
  1174=>"00000001",
  1175=>"00000010",
  1176=>"11111111",
  1177=>"00000000",
  1178=>"11111111",
  1179=>"11111110",
  1180=>"11111111",
  1181=>"00000000",
  1182=>"11111110",
  1183=>"00000001",
  1184=>"00000010",
  1185=>"00000000",
  1186=>"00000010",
  1187=>"11111110",
  1188=>"00000001",
  1189=>"11111111",
  1190=>"00000001",
  1191=>"11111111",
  1192=>"11111111",
  1193=>"00000001",
  1194=>"00000000",
  1195=>"11111111",
  1196=>"00000010",
  1197=>"00000010",
  1198=>"00000010",
  1199=>"00000000",
  1200=>"00000010",
  1201=>"00000010",
  1202=>"00000000",
  1203=>"00000001",
  1204=>"11111110",
  1205=>"11111111",
  1206=>"00000000",
  1207=>"00000000",
  1208=>"00000000",
  1209=>"00000000",
  1210=>"00000000",
  1211=>"11111111",
  1212=>"11111110",
  1213=>"00000001",
  1214=>"00000000",
  1215=>"11111111",
  1216=>"11111111",
  1217=>"00000001",
  1218=>"11111111",
  1219=>"00000010",
  1220=>"00000011",
  1221=>"00000010",
  1222=>"11111111",
  1223=>"11111110",
  1224=>"00000000",
  1225=>"00000001",
  1226=>"00000001",
  1227=>"00000001",
  1228=>"00000000",
  1229=>"11111111",
  1230=>"00000001",
  1231=>"00000000",
  1232=>"11111111",
  1233=>"11111111",
  1234=>"11111110",
  1235=>"00000001",
  1236=>"11111111",
  1237=>"00000001",
  1238=>"00000010",
  1239=>"11111110",
  1240=>"11111111",
  1241=>"00000000",
  1242=>"11111110",
  1243=>"00000000",
  1244=>"11111111",
  1245=>"00000010",
  1246=>"00000001",
  1247=>"00000001",
  1248=>"00000000",
  1249=>"11111111",
  1250=>"11111111",
  1251=>"00000000",
  1252=>"11111111",
  1253=>"11111111",
  1254=>"00000000",
  1255=>"00000010",
  1256=>"11111110",
  1257=>"11111111",
  1258=>"11111111",
  1259=>"00000001",
  1260=>"11111111",
  1261=>"11111111",
  1262=>"00000011",
  1263=>"00000000",
  1264=>"11111111",
  1265=>"11111110",
  1266=>"00000000",
  1267=>"00000010",
  1268=>"00000001",
  1269=>"11111111",
  1270=>"00000010",
  1271=>"11111110",
  1272=>"00000001",
  1273=>"11111110",
  1274=>"00000001",
  1275=>"11111110",
  1276=>"00000010",
  1277=>"00000001",
  1278=>"00000000",
  1279=>"11111111",
  1280=>"00000010",
  1281=>"00000001",
  1282=>"00000001",
  1283=>"11111110",
  1284=>"11111111",
  1285=>"11111111",
  1286=>"00000000",
  1287=>"11111111",
  1288=>"11111110",
  1289=>"11111111",
  1290=>"00000010",
  1291=>"00000000",
  1292=>"11111110",
  1293=>"00000010",
  1294=>"00000000",
  1295=>"00000001",
  1296=>"00000001",
  1297=>"00000001",
  1298=>"00000001",
  1299=>"00000001",
  1300=>"11111101",
  1301=>"00000001",
  1302=>"00000010",
  1303=>"00000001",
  1304=>"00000010",
  1305=>"00000000",
  1306=>"00000001",
  1307=>"00000000",
  1308=>"11111111",
  1309=>"11111111",
  1310=>"00000010",
  1311=>"00000010",
  1312=>"11111111",
  1313=>"11111111",
  1314=>"00000100",
  1315=>"00000001",
  1316=>"00000001",
  1317=>"00000001",
  1318=>"00000001",
  1319=>"00000001",
  1320=>"00000010",
  1321=>"00000011",
  1322=>"00000000",
  1323=>"11111110",
  1324=>"00000001",
  1325=>"00000011",
  1326=>"00000001",
  1327=>"00000001",
  1328=>"00000001",
  1329=>"00000001",
  1330=>"11111111",
  1331=>"00000001",
  1332=>"11111111",
  1333=>"11111110",
  1334=>"00000001",
  1335=>"00000011",
  1336=>"00000000",
  1337=>"11111111",
  1338=>"00000000",
  1339=>"00000001",
  1340=>"00000001",
  1341=>"00000000",
  1342=>"00000000",
  1343=>"00000011",
  1344=>"00000001",
  1345=>"00000001",
  1346=>"00000000",
  1347=>"11111111",
  1348=>"00000000",
  1349=>"00000000",
  1350=>"00000000",
  1351=>"11111111",
  1352=>"11111111",
  1353=>"00000001",
  1354=>"00000000",
  1355=>"11111110",
  1356=>"00000010",
  1357=>"00000000",
  1358=>"00000001",
  1359=>"00000000",
  1360=>"00000001",
  1361=>"11111110",
  1362=>"00000000",
  1363=>"11111111",
  1364=>"11111101",
  1365=>"00000010",
  1366=>"11111111",
  1367=>"00000001",
  1368=>"11111111",
  1369=>"00000000",
  1370=>"00000000",
  1371=>"11111111",
  1372=>"11111111",
  1373=>"00000011",
  1374=>"11111110",
  1375=>"00000010",
  1376=>"00000000",
  1377=>"00000001",
  1378=>"00000000",
  1379=>"00000011",
  1380=>"00000011",
  1381=>"00000001",
  1382=>"11111111",
  1383=>"11111111",
  1384=>"11111111",
  1385=>"00000001",
  1386=>"11111111",
  1387=>"00000000",
  1388=>"11111101",
  1389=>"11111110",
  1390=>"00000010",
  1391=>"11111101",
  1392=>"11111110",
  1393=>"11111110",
  1394=>"11111111",
  1395=>"11111110",
  1396=>"11111110",
  1397=>"00000000",
  1398=>"00000001",
  1399=>"00000000",
  1400=>"11111111",
  1401=>"11111111",
  1402=>"00000000",
  1403=>"11111110",
  1404=>"11111111",
  1405=>"00000000",
  1406=>"11111110",
  1407=>"00000001",
  1408=>"11111111",
  1409=>"11111111",
  1410=>"00000001",
  1411=>"11111110",
  1412=>"11111111",
  1413=>"11111110",
  1414=>"00000000",
  1415=>"00000001",
  1416=>"00000000",
  1417=>"00000001",
  1418=>"00000010",
  1419=>"00000010",
  1420=>"00000001",
  1421=>"00000010",
  1422=>"00000010",
  1423=>"00000001",
  1424=>"00000010",
  1425=>"11111110",
  1426=>"00000001",
  1427=>"11111110",
  1428=>"00000000",
  1429=>"00000001",
  1430=>"00000000",
  1431=>"11111111",
  1432=>"00000001",
  1433=>"00000010",
  1434=>"00000000",
  1435=>"11111111",
  1436=>"11111111",
  1437=>"00000001",
  1438=>"00000010",
  1439=>"00000000",
  1440=>"11111111",
  1441=>"00000000",
  1442=>"00000000",
  1443=>"11111111",
  1444=>"00000001",
  1445=>"00000010",
  1446=>"11111110",
  1447=>"11111111",
  1448=>"00000000",
  1449=>"11111111",
  1450=>"11111111",
  1451=>"11111111",
  1452=>"00000010",
  1453=>"11111110",
  1454=>"00000010",
  1455=>"00000001",
  1456=>"11111110",
  1457=>"00000001",
  1458=>"00000001",
  1459=>"00000000",
  1460=>"11111111",
  1461=>"11111111",
  1462=>"11111110",
  1463=>"11111111",
  1464=>"11111111",
  1465=>"00000001",
  1466=>"00000000",
  1467=>"00000001",
  1468=>"11111111",
  1469=>"11111111",
  1470=>"00000010",
  1471=>"00000000",
  1472=>"00000001",
  1473=>"11111111",
  1474=>"00000010",
  1475=>"00000000",
  1476=>"11111111",
  1477=>"11111110",
  1478=>"00000001",
  1479=>"00000010",
  1480=>"11111110",
  1481=>"00000001",
  1482=>"00000001",
  1483=>"00000010",
  1484=>"00000010",
  1485=>"00000001",
  1486=>"00000001",
  1487=>"00000010",
  1488=>"00000001",
  1489=>"00000000",
  1490=>"00000000",
  1491=>"00000001",
  1492=>"00000010",
  1493=>"00000000",
  1494=>"11111110",
  1495=>"00000001",
  1496=>"11111111",
  1497=>"00000000",
  1498=>"11111111",
  1499=>"00000000",
  1500=>"00000001",
  1501=>"11111111",
  1502=>"11111111",
  1503=>"00000001",
  1504=>"00000001",
  1505=>"11111111",
  1506=>"00000011",
  1507=>"00000001",
  1508=>"11111110",
  1509=>"00000001",
  1510=>"00000001",
  1511=>"11111111",
  1512=>"00000000",
  1513=>"11111111",
  1514=>"11111111",
  1515=>"00000000",
  1516=>"00000010",
  1517=>"11111110",
  1518=>"11111111",
  1519=>"11111111",
  1520=>"00000001",
  1521=>"00000010",
  1522=>"11111110",
  1523=>"00000001",
  1524=>"00000000",
  1525=>"11111110",
  1526=>"11111111",
  1527=>"00000000",
  1528=>"00000001",
  1529=>"00000001",
  1530=>"11111111",
  1531=>"11111111",
  1532=>"11111110",
  1533=>"00000000",
  1534=>"00000011",
  1535=>"00000000",
  1536=>"00000001",
  1537=>"00000010",
  1538=>"00000000",
  1539=>"11111101",
  1540=>"00000000",
  1541=>"11111110",
  1542=>"00000001",
  1543=>"11111110",
  1544=>"11111111",
  1545=>"00000001",
  1546=>"00000001",
  1547=>"11111111",
  1548=>"00000010",
  1549=>"11111110",
  1550=>"00000000",
  1551=>"00000000",
  1552=>"00000010",
  1553=>"00000000",
  1554=>"11111101",
  1555=>"00000000",
  1556=>"00000000",
  1557=>"00000000",
  1558=>"00000010",
  1559=>"11111111",
  1560=>"11111111",
  1561=>"11111111",
  1562=>"00000000",
  1563=>"11111111",
  1564=>"00000010",
  1565=>"00000000",
  1566=>"11111110",
  1567=>"00000000",
  1568=>"00000000",
  1569=>"00000010",
  1570=>"00000001",
  1571=>"11111111",
  1572=>"00000001",
  1573=>"11111101",
  1574=>"00000000",
  1575=>"00000011",
  1576=>"00000010",
  1577=>"11111111",
  1578=>"11111110",
  1579=>"00000010",
  1580=>"11111111",
  1581=>"00000000",
  1582=>"11111111",
  1583=>"11111110",
  1584=>"00000010",
  1585=>"00000000",
  1586=>"00000000",
  1587=>"00000000",
  1588=>"00000010",
  1589=>"11111111",
  1590=>"00000000",
  1591=>"00000010",
  1592=>"00000001",
  1593=>"00000000",
  1594=>"11111111",
  1595=>"11111111",
  1596=>"00000001",
  1597=>"11111111",
  1598=>"00000001",
  1599=>"11111111",
  1600=>"00000010",
  1601=>"11111111",
  1602=>"00000000",
  1603=>"00000000",
  1604=>"00000000",
  1605=>"11111111",
  1606=>"00000000",
  1607=>"11111111",
  1608=>"11111110",
  1609=>"00000000",
  1610=>"11111110",
  1611=>"11111111",
  1612=>"11111111",
  1613=>"11111110",
  1614=>"11111111",
  1615=>"11111110",
  1616=>"00000000",
  1617=>"00000010",
  1618=>"11111111",
  1619=>"11111111",
  1620=>"11111110",
  1621=>"11111110",
  1622=>"00000000",
  1623=>"00000000",
  1624=>"11111111",
  1625=>"00000001",
  1626=>"11111110",
  1627=>"11111110",
  1628=>"11111110",
  1629=>"00000011",
  1630=>"00000000",
  1631=>"11111101",
  1632=>"00000000",
  1633=>"11111110",
  1634=>"00000001",
  1635=>"00000001",
  1636=>"11111111",
  1637=>"11111111",
  1638=>"11111111",
  1639=>"11111111",
  1640=>"00000001",
  1641=>"11111110",
  1642=>"00000000",
  1643=>"00000001",
  1644=>"00000000",
  1645=>"00000010",
  1646=>"11111110",
  1647=>"11111111",
  1648=>"00000001",
  1649=>"00000001",
  1650=>"00000000",
  1651=>"00000001",
  1652=>"00000001",
  1653=>"11111110",
  1654=>"00000000",
  1655=>"11111111",
  1656=>"00000010",
  1657=>"11111111",
  1658=>"11111111",
  1659=>"00000011",
  1660=>"00000000",
  1661=>"00000001",
  1662=>"00000001",
  1663=>"00000001",
  1664=>"00000011",
  1665=>"00000001",
  1666=>"11111111",
  1667=>"11111110",
  1668=>"00000001",
  1669=>"00000001",
  1670=>"11111111",
  1671=>"11111111",
  1672=>"00000010",
  1673=>"00000011",
  1674=>"11111111",
  1675=>"00000000",
  1676=>"00000010",
  1677=>"00000000",
  1678=>"00000010",
  1679=>"00000000",
  1680=>"11111110",
  1681=>"00000000",
  1682=>"00000000",
  1683=>"00000001",
  1684=>"00000000",
  1685=>"00000001",
  1686=>"00000010",
  1687=>"00000000",
  1688=>"11111110",
  1689=>"11111111",
  1690=>"11111111",
  1691=>"00000000",
  1692=>"00000001",
  1693=>"11111110",
  1694=>"00000000",
  1695=>"00000001",
  1696=>"00000000",
  1697=>"00000001",
  1698=>"00000011",
  1699=>"00000000",
  1700=>"00000000",
  1701=>"11111110",
  1702=>"00000001",
  1703=>"11111111",
  1704=>"11111110",
  1705=>"00000000",
  1706=>"00000001",
  1707=>"11111110",
  1708=>"00000010",
  1709=>"00000000",
  1710=>"00000001",
  1711=>"11111110",
  1712=>"00000010",
  1713=>"11111110",
  1714=>"00000001",
  1715=>"11111111",
  1716=>"00000010",
  1717=>"00000001",
  1718=>"00000011",
  1719=>"11111111",
  1720=>"00000001",
  1721=>"11111111",
  1722=>"00000000",
  1723=>"11111111",
  1724=>"00000000",
  1725=>"00000001",
  1726=>"11111111",
  1727=>"00000010",
  1728=>"00000000",
  1729=>"11111110",
  1730=>"11111110",
  1731=>"00000010",
  1732=>"11111110",
  1733=>"11111111",
  1734=>"00000000",
  1735=>"11111111",
  1736=>"00000001",
  1737=>"11111110",
  1738=>"11111110",
  1739=>"00000000",
  1740=>"00000001",
  1741=>"11111111",
  1742=>"00000000",
  1743=>"00000001",
  1744=>"11111111",
  1745=>"11111110",
  1746=>"11111110",
  1747=>"00000010",
  1748=>"00000010",
  1749=>"11111101",
  1750=>"11111110",
  1751=>"00000000",
  1752=>"11111111",
  1753=>"00000000",
  1754=>"00000010",
  1755=>"00000000",
  1756=>"11111111",
  1757=>"11111111",
  1758=>"11111111",
  1759=>"00000010",
  1760=>"11111111",
  1761=>"00000000",
  1762=>"00000011",
  1763=>"11111111",
  1764=>"00000001",
  1765=>"11111101",
  1766=>"00000001",
  1767=>"00000000",
  1768=>"11111111",
  1769=>"11111111",
  1770=>"00000001",
  1771=>"00000010",
  1772=>"11111111",
  1773=>"00000000",
  1774=>"00000001",
  1775=>"00000000",
  1776=>"00000000",
  1777=>"00000010",
  1778=>"00000000",
  1779=>"00000000",
  1780=>"00000001",
  1781=>"00000000",
  1782=>"11111110",
  1783=>"11111101",
  1784=>"11111110",
  1785=>"00000010",
  1786=>"11111111",
  1787=>"11111111",
  1788=>"11111110",
  1789=>"00000001",
  1790=>"11111111",
  1791=>"11111111",
  1792=>"11111111",
  1793=>"00000000",
  1794=>"00000000",
  1795=>"11111110",
  1796=>"00000000",
  1797=>"00000000",
  1798=>"11111111",
  1799=>"00000001",
  1800=>"00000000",
  1801=>"11111111",
  1802=>"00000001",
  1803=>"00000001",
  1804=>"00000001",
  1805=>"00000000",
  1806=>"00000000",
  1807=>"11111110",
  1808=>"11111110",
  1809=>"00000000",
  1810=>"00000001",
  1811=>"00000010",
  1812=>"11111110",
  1813=>"00000001",
  1814=>"00000001",
  1815=>"11111110",
  1816=>"00000000",
  1817=>"00000001",
  1818=>"00000000",
  1819=>"00000010",
  1820=>"11111111",
  1821=>"11111110",
  1822=>"11111110",
  1823=>"00000001",
  1824=>"11111110",
  1825=>"00000010",
  1826=>"00000001",
  1827=>"00000001",
  1828=>"11111101",
  1829=>"11111110",
  1830=>"00000001",
  1831=>"00000000",
  1832=>"11111111",
  1833=>"00000000",
  1834=>"11111111",
  1835=>"00000001",
  1836=>"00000001",
  1837=>"00000001",
  1838=>"00000001",
  1839=>"00000010",
  1840=>"00000000",
  1841=>"00000000",
  1842=>"00000001",
  1843=>"11111111",
  1844=>"11111111",
  1845=>"00000001",
  1846=>"00000000",
  1847=>"00000010",
  1848=>"11111110",
  1849=>"11111101",
  1850=>"00000001",
  1851=>"11111111",
  1852=>"11111111",
  1853=>"00000001",
  1854=>"00000001",
  1855=>"00000000",
  1856=>"11111111",
  1857=>"00000000",
  1858=>"11111111",
  1859=>"11111111",
  1860=>"11111111",
  1861=>"11111110",
  1862=>"00000010",
  1863=>"00000001",
  1864=>"00000000",
  1865=>"11111111",
  1866=>"00000000",
  1867=>"11111110",
  1868=>"00000010",
  1869=>"11111110",
  1870=>"00000001",
  1871=>"11111111",
  1872=>"00000001",
  1873=>"00000000",
  1874=>"00000000",
  1875=>"00000010",
  1876=>"11111111",
  1877=>"11111111",
  1878=>"00000001",
  1879=>"11111110",
  1880=>"00000001",
  1881=>"11111111",
  1882=>"00000000",
  1883=>"00000001",
  1884=>"00000010",
  1885=>"11111111",
  1886=>"11111111",
  1887=>"11111111",
  1888=>"00000001",
  1889=>"00000000",
  1890=>"00000000",
  1891=>"11111111",
  1892=>"00000000",
  1893=>"11111110",
  1894=>"00000001",
  1895=>"00000001",
  1896=>"00000000",
  1897=>"11111110",
  1898=>"00000011",
  1899=>"00000000",
  1900=>"00000000",
  1901=>"00000001",
  1902=>"00000001",
  1903=>"00000010",
  1904=>"00000000",
  1905=>"11111111",
  1906=>"00000010",
  1907=>"00000000",
  1908=>"00000000",
  1909=>"00000010",
  1910=>"00000010",
  1911=>"00000011",
  1912=>"11111110",
  1913=>"00000000",
  1914=>"00000000",
  1915=>"00000011",
  1916=>"00000000",
  1917=>"00000001",
  1918=>"11111110",
  1919=>"11111110",
  1920=>"11111111",
  1921=>"00000000",
  1922=>"00000000",
  1923=>"00000001",
  1924=>"00000001",
  1925=>"11111111",
  1926=>"00000001",
  1927=>"00000000",
  1928=>"11111110",
  1929=>"00000010",
  1930=>"00000001",
  1931=>"00000000",
  1932=>"00000000",
  1933=>"00000000",
  1934=>"00000000",
  1935=>"00000001",
  1936=>"00000001",
  1937=>"11111110",
  1938=>"11111111",
  1939=>"11111111",
  1940=>"11111110",
  1941=>"00000000",
  1942=>"11111110",
  1943=>"11111101",
  1944=>"00000010",
  1945=>"00000001",
  1946=>"11111110",
  1947=>"00000000",
  1948=>"11111111",
  1949=>"11111111",
  1950=>"00000000",
  1951=>"00000001",
  1952=>"00000010",
  1953=>"11111110",
  1954=>"00000000",
  1955=>"00000001",
  1956=>"00000000",
  1957=>"11111111",
  1958=>"11111110",
  1959=>"00000001",
  1960=>"00000010",
  1961=>"00000001",
  1962=>"11111111",
  1963=>"00000000",
  1964=>"00000000",
  1965=>"00000000",
  1966=>"11111111",
  1967=>"00000001",
  1968=>"00000010",
  1969=>"00000001",
  1970=>"11111110",
  1971=>"00000011",
  1972=>"00000000",
  1973=>"11111111",
  1974=>"11111110",
  1975=>"11111111",
  1976=>"11111110",
  1977=>"11111111",
  1978=>"00000000",
  1979=>"00000000",
  1980=>"00000000",
  1981=>"11111111",
  1982=>"11111110",
  1983=>"11111111",
  1984=>"00000000",
  1985=>"00000001",
  1986=>"00000010",
  1987=>"11111110",
  1988=>"11111111",
  1989=>"00000001",
  1990=>"00000000",
  1991=>"00000011",
  1992=>"00000001",
  1993=>"00000010",
  1994=>"00000000",
  1995=>"00000010",
  1996=>"11111110",
  1997=>"00000001",
  1998=>"00000010",
  1999=>"00000001",
  2000=>"00000001",
  2001=>"00000011",
  2002=>"00000010",
  2003=>"11111110",
  2004=>"11111111",
  2005=>"00000001",
  2006=>"00000000",
  2007=>"11111111",
  2008=>"11111101",
  2009=>"11111111",
  2010=>"00000010",
  2011=>"11111111",
  2012=>"00000000",
  2013=>"11111110",
  2014=>"00000000",
  2015=>"11111111",
  2016=>"00000010",
  2017=>"00000000",
  2018=>"11111111",
  2019=>"00000010",
  2020=>"11111111",
  2021=>"00000001",
  2022=>"00000011",
  2023=>"11111110",
  2024=>"11111111",
  2025=>"00000000",
  2026=>"11111110",
  2027=>"00000001",
  2028=>"11111111",
  2029=>"00000010",
  2030=>"00000000",
  2031=>"11111110",
  2032=>"00000010",
  2033=>"11111111",
  2034=>"00000000",
  2035=>"11111110",
  2036=>"11111111",
  2037=>"00000001",
  2038=>"00000000",
  2039=>"11111111",
  2040=>"00000001",
  2041=>"00000001",
  2042=>"00000001",
  2043=>"11111110",
  2044=>"11111110",
  2045=>"11111111",
  2046=>"00000001",
  2047=>"00000010",
  2048=>"00000001",
  2049=>"00000000",
  2050=>"00000001",
  2051=>"11111110",
  2052=>"00000000",
  2053=>"00000001",
  2054=>"11111111",
  2055=>"00000000",
  2056=>"00000000",
  2057=>"00000000",
  2058=>"11111111",
  2059=>"00000000",
  2060=>"00000001",
  2061=>"00000000",
  2062=>"11111111",
  2063=>"00000001",
  2064=>"00000000",
  2065=>"11111111",
  2066=>"00000001",
  2067=>"00000000",
  2068=>"00000000",
  2069=>"11111111",
  2070=>"00000001",
  2071=>"11111111",
  2072=>"00000000",
  2073=>"11111111",
  2074=>"00000000",
  2075=>"11111110",
  2076=>"00000000",
  2077=>"00000000",
  2078=>"00000000",
  2079=>"00000000",
  2080=>"00000000",
  2081=>"00000000",
  2082=>"00000000",
  2083=>"11111111",
  2084=>"00000001",
  2085=>"11111111",
  2086=>"11111111",
  2087=>"00000000",
  2088=>"11111111",
  2089=>"00000000",
  2090=>"00000000",
  2091=>"00000000",
  2092=>"11111110",
  2093=>"00000000",
  2094=>"11111111",
  2095=>"00000001",
  2096=>"11111110",
  2097=>"11111110",
  2098=>"00000001",
  2099=>"00000001",
  2100=>"11111111",
  2101=>"00000000",
  2102=>"11111111",
  2103=>"00000000",
  2104=>"00000000",
  2105=>"00000001",
  2106=>"11111111",
  2107=>"11111111",
  2108=>"00000010",
  2109=>"00000000",
  2110=>"00000000",
  2111=>"00000000",
  2112=>"00000000",
  2113=>"00000000",
  2114=>"00000010",
  2115=>"11111111",
  2116=>"00000001",
  2117=>"11111111",
  2118=>"00000001",
  2119=>"00000000",
  2120=>"00000000",
  2121=>"00000000",
  2122=>"00000000",
  2123=>"00000011",
  2124=>"00000000",
  2125=>"00000001",
  2126=>"11111111",
  2127=>"00000000",
  2128=>"00000000",
  2129=>"00000000",
  2130=>"00000000",
  2131=>"00000000",
  2132=>"00000000",
  2133=>"00000000",
  2134=>"00000000",
  2135=>"00000001",
  2136=>"00000000",
  2137=>"00000000",
  2138=>"00000000",
  2139=>"00000000",
  2140=>"00000001",
  2141=>"00000000",
  2142=>"11111111",
  2143=>"00000000",
  2144=>"00000000",
  2145=>"11111111",
  2146=>"00000000",
  2147=>"11111111",
  2148=>"00000001",
  2149=>"00000000",
  2150=>"00000000",
  2151=>"00000000",
  2152=>"00000000",
  2153=>"00000000",
  2154=>"00000000",
  2155=>"00000000",
  2156=>"00000001",
  2157=>"00000000",
  2158=>"11111111",
  2159=>"00000000",
  2160=>"00000001",
  2161=>"00000000",
  2162=>"00000001",
  2163=>"00000000",
  2164=>"00000000",
  2165=>"00000000",
  2166=>"00000000",
  2167=>"00000000",
  2168=>"11111111",
  2169=>"00000000",
  2170=>"00000000",
  2171=>"00000000",
  2172=>"11111111",
  2173=>"00000000",
  2174=>"00000000",
  2175=>"00000000",
  2176=>"00000000",
  2177=>"00000000",
  2178=>"00000000",
  2179=>"00000000",
  2180=>"11111111",
  2181=>"11111111",
  2182=>"11111110",
  2183=>"00000000",
  2184=>"00000001",
  2185=>"00000001",
  2186=>"00000000",
  2187=>"00000000",
  2188=>"00000000",
  2189=>"00000000",
  2190=>"11111111",
  2191=>"11111111",
  2192=>"00000000",
  2193=>"00000000",
  2194=>"00000000",
  2195=>"11111111",
  2196=>"00000000",
  2197=>"00000000",
  2198=>"11111110",
  2199=>"00000000",
  2200=>"00000001",
  2201=>"00000000",
  2202=>"00000000",
  2203=>"00000000",
  2204=>"11111111",
  2205=>"00000000",
  2206=>"11111111",
  2207=>"00000000",
  2208=>"11111111",
  2209=>"00000000",
  2210=>"00000001",
  2211=>"00000000",
  2212=>"00000010",
  2213=>"00000000",
  2214=>"00000000",
  2215=>"11111111",
  2216=>"00000001",
  2217=>"00000000",
  2218=>"00000000",
  2219=>"00000000",
  2220=>"00000000",
  2221=>"00000000",
  2222=>"00000000",
  2223=>"11111110",
  2224=>"00000000",
  2225=>"00000000",
  2226=>"11111111",
  2227=>"00000000",
  2228=>"11111111",
  2229=>"00000000",
  2230=>"00000000",
  2231=>"00000000",
  2232=>"00000000",
  2233=>"00000000",
  2234=>"00000000",
  2235=>"00000000",
  2236=>"00000000",
  2237=>"00000000",
  2238=>"00000000",
  2239=>"00000001",
  2240=>"00000000",
  2241=>"00000000",
  2242=>"00000000",
  2243=>"00000000",
  2244=>"00000000",
  2245=>"00000000",
  2246=>"00000000",
  2247=>"11111110",
  2248=>"11111111",
  2249=>"00000000",
  2250=>"00000000",
  2251=>"00000000",
  2252=>"00000000",
  2253=>"00000000",
  2254=>"00000000",
  2255=>"00000000",
  2256=>"00000000",
  2257=>"00000001",
  2258=>"11111111",
  2259=>"11111111",
  2260=>"11111110",
  2261=>"00000000",
  2262=>"00000001",
  2263=>"00000000",
  2264=>"00000000",
  2265=>"11111110",
  2266=>"00000000",
  2267=>"00000000",
  2268=>"00000000",
  2269=>"00000000",
  2270=>"11111111",
  2271=>"00000000",
  2272=>"00000000",
  2273=>"00000000",
  2274=>"00000000",
  2275=>"00000000",
  2276=>"00000000",
  2277=>"00000000",
  2278=>"11111111",
  2279=>"00000000",
  2280=>"00000010",
  2281=>"11111111",
  2282=>"00000000",
  2283=>"00000010",
  2284=>"00000000",
  2285=>"00000000",
  2286=>"00000000",
  2287=>"11111010",
  2288=>"00000000",
  2289=>"00000000",
  2290=>"00000000",
  2291=>"00000001",
  2292=>"00000000",
  2293=>"00000000",
  2294=>"11111111",
  2295=>"00000000",
  2296=>"11111111",
  2297=>"11111101",
  2298=>"00000000",
  2299=>"00000001",
  2300=>"00000001",
  2301=>"00000000",
  2302=>"00000001",
  2303=>"00000000",
  2304=>"11111111",
  2305=>"00000000",
  2306=>"11111101",
  2307=>"00000000",
  2308=>"00000000",
  2309=>"00000000",
  2310=>"00000000",
  2311=>"00000000",
  2312=>"00000000",
  2313=>"00000000",
  2314=>"00000000",
  2315=>"00000000",
  2316=>"00000001",
  2317=>"00000000",
  2318=>"00000000",
  2319=>"00000000",
  2320=>"11111111",
  2321=>"00000000",
  2322=>"00000000",
  2323=>"00000000",
  2324=>"00000000",
  2325=>"00000000",
  2326=>"00000000",
  2327=>"00000000",
  2328=>"00000000",
  2329=>"11111111",
  2330=>"11111111",
  2331=>"00000000",
  2332=>"00000000",
  2333=>"00000001",
  2334=>"11111111",
  2335=>"00000000",
  2336=>"00000001",
  2337=>"00000010",
  2338=>"00000001",
  2339=>"00000000",
  2340=>"00000000",
  2341=>"00000000",
  2342=>"00000001",
  2343=>"00000000",
  2344=>"00000001",
  2345=>"11111111",
  2346=>"00000000",
  2347=>"00000000",
  2348=>"00000001",
  2349=>"11111101",
  2350=>"11111111",
  2351=>"11111111",
  2352=>"00000001",
  2353=>"00000000",
  2354=>"00000000",
  2355=>"11111111",
  2356=>"00000001",
  2357=>"00000000",
  2358=>"00000000",
  2359=>"11111111",
  2360=>"00000000",
  2361=>"00000000",
  2362=>"11111110",
  2363=>"11111111",
  2364=>"00000001",
  2365=>"00000010",
  2366=>"00000000",
  2367=>"00000000",
  2368=>"11111110",
  2369=>"00000001",
  2370=>"00000001",
  2371=>"11111111",
  2372=>"11111111",
  2373=>"00000000",
  2374=>"00000000",
  2375=>"00000001",
  2376=>"11111111",
  2377=>"00000000",
  2378=>"00000000",
  2379=>"00000001",
  2380=>"00000000",
  2381=>"00000010",
  2382=>"00000000",
  2383=>"00000000",
  2384=>"00000000",
  2385=>"00000000",
  2386=>"11111111",
  2387=>"00000000",
  2388=>"00000010",
  2389=>"00000001",
  2390=>"00000000",
  2391=>"11111111",
  2392=>"00000000",
  2393=>"00000000",
  2394=>"00000001",
  2395=>"00000000",
  2396=>"00000000",
  2397=>"00000000",
  2398=>"00000000",
  2399=>"11111111",
  2400=>"00000000",
  2401=>"11111111",
  2402=>"00000000",
  2403=>"00000000",
  2404=>"11111111",
  2405=>"00000000",
  2406=>"00000001",
  2407=>"00000001",
  2408=>"00000000",
  2409=>"00000000",
  2410=>"00000000",
  2411=>"00000010",
  2412=>"11111111",
  2413=>"00000000",
  2414=>"11111111",
  2415=>"00000000",
  2416=>"11111101",
  2417=>"00000000",
  2418=>"00000000",
  2419=>"11111111",
  2420=>"00000000",
  2421=>"00000001",
  2422=>"00000001",
  2423=>"00000000",
  2424=>"00000000",
  2425=>"00000000",
  2426=>"00000000",
  2427=>"11111111",
  2428=>"11111111",
  2429=>"11111111",
  2430=>"00000000",
  2431=>"00000000",
  2432=>"00000000",
  2433=>"00000000",
  2434=>"00000010",
  2435=>"00000000",
  2436=>"11111111",
  2437=>"00000001",
  2438=>"11111111",
  2439=>"11111111",
  2440=>"00000000",
  2441=>"00000000",
  2442=>"00000001",
  2443=>"00000001",
  2444=>"00000000",
  2445=>"00000010",
  2446=>"00000000",
  2447=>"00000000",
  2448=>"11111110",
  2449=>"00000000",
  2450=>"00000000",
  2451=>"00000000",
  2452=>"00000001",
  2453=>"00000000",
  2454=>"00000001",
  2455=>"00000000",
  2456=>"11111111",
  2457=>"00000000",
  2458=>"11111111",
  2459=>"00000000",
  2460=>"00000001",
  2461=>"11111111",
  2462=>"00000000",
  2463=>"00000000",
  2464=>"00000001",
  2465=>"11111111",
  2466=>"00000010",
  2467=>"00000001",
  2468=>"11111111",
  2469=>"00000001",
  2470=>"00000001",
  2471=>"00000000",
  2472=>"00000000",
  2473=>"00000000",
  2474=>"00000001",
  2475=>"11111111",
  2476=>"00000001",
  2477=>"00000000",
  2478=>"00000001",
  2479=>"00000000",
  2480=>"00000000",
  2481=>"00000000",
  2482=>"00000000",
  2483=>"00000001",
  2484=>"00000001",
  2485=>"00000000",
  2486=>"00000000",
  2487=>"11111111",
  2488=>"11111111",
  2489=>"00000001",
  2490=>"11111111",
  2491=>"00000000",
  2492=>"11111101",
  2493=>"00000001",
  2494=>"11111111",
  2495=>"11111111",
  2496=>"00000001",
  2497=>"00000000",
  2498=>"00000000",
  2499=>"00000000",
  2500=>"11111111",
  2501=>"00000000",
  2502=>"00000001",
  2503=>"00000000",
  2504=>"00000010",
  2505=>"00000000",
  2506=>"00000000",
  2507=>"00000000",
  2508=>"00000000",
  2509=>"11111111",
  2510=>"00000000",
  2511=>"00000000",
  2512=>"00000000",
  2513=>"00000000",
  2514=>"00000011",
  2515=>"00000001",
  2516=>"11111111",
  2517=>"00000001",
  2518=>"00000001",
  2519=>"11111110",
  2520=>"00000000",
  2521=>"00000000",
  2522=>"00000000",
  2523=>"11111111",
  2524=>"00000000",
  2525=>"11111111",
  2526=>"00000001",
  2527=>"00000000",
  2528=>"00000001",
  2529=>"00000000",
  2530=>"11111111",
  2531=>"00000001",
  2532=>"00000000",
  2533=>"00000000",
  2534=>"11111111",
  2535=>"11111110",
  2536=>"00000000",
  2537=>"00000000",
  2538=>"00000000",
  2539=>"00000001",
  2540=>"00000000",
  2541=>"00000000",
  2542=>"00000000",
  2543=>"00000000",
  2544=>"00000000",
  2545=>"00000000",
  2546=>"00000010",
  2547=>"00000001",
  2548=>"00000000",
  2549=>"00000000",
  2550=>"00000000",
  2551=>"00000000",
  2552=>"00000001",
  2553=>"00000000",
  2554=>"00000000",
  2555=>"00000000",
  2556=>"00000001",
  2557=>"00000000",
  2558=>"00000000",
  2559=>"00000001",
  2560=>"00000010",
  2561=>"11111111",
  2562=>"00000000",
  2563=>"00000000",
  2564=>"00000000",
  2565=>"00000001",
  2566=>"00000000",
  2567=>"00000000",
  2568=>"11111111",
  2569=>"00000000",
  2570=>"11111111",
  2571=>"00000001",
  2572=>"00000001",
  2573=>"00000000",
  2574=>"00000000",
  2575=>"11111111",
  2576=>"00000000",
  2577=>"00000000",
  2578=>"11111111",
  2579=>"00000000",
  2580=>"00000000",
  2581=>"11111110",
  2582=>"11111111",
  2583=>"00000000",
  2584=>"11111111",
  2585=>"00000000",
  2586=>"00000000",
  2587=>"00000000",
  2588=>"00000001",
  2589=>"00000001",
  2590=>"11111111",
  2591=>"00000000",
  2592=>"11111111",
  2593=>"00000001",
  2594=>"00000000",
  2595=>"11111111",
  2596=>"00000001",
  2597=>"00000000",
  2598=>"00000000",
  2599=>"00000000",
  2600=>"00000001",
  2601=>"11111110",
  2602=>"00000000",
  2603=>"11111111",
  2604=>"00000000",
  2605=>"11111111",
  2606=>"00000000",
  2607=>"00000000",
  2608=>"00000000",
  2609=>"00000001",
  2610=>"00000010",
  2611=>"00000000",
  2612=>"00000000",
  2613=>"00000000",
  2614=>"00000000",
  2615=>"00000001",
  2616=>"00000000",
  2617=>"00000000",
  2618=>"00000001",
  2619=>"00000000",
  2620=>"00000000",
  2621=>"11111110",
  2622=>"00000000",
  2623=>"00000000",
  2624=>"11111111",
  2625=>"00000000",
  2626=>"00000001",
  2627=>"00000001",
  2628=>"00000001",
  2629=>"11111111",
  2630=>"00000000",
  2631=>"00000000",
  2632=>"11111111",
  2633=>"11111111",
  2634=>"11111111",
  2635=>"00000000",
  2636=>"00000000",
  2637=>"11111111",
  2638=>"11111111",
  2639=>"00000000",
  2640=>"00000000",
  2641=>"00000000",
  2642=>"00000000",
  2643=>"00000010",
  2644=>"00000001",
  2645=>"00000000",
  2646=>"00000000",
  2647=>"00000000",
  2648=>"00000000",
  2649=>"00000000",
  2650=>"00000000",
  2651=>"11111111",
  2652=>"00000000",
  2653=>"00000001",
  2654=>"00000000",
  2655=>"00000000",
  2656=>"00000000",
  2657=>"11111111",
  2658=>"00000001",
  2659=>"00000000",
  2660=>"11111111",
  2661=>"00000000",
  2662=>"11111111",
  2663=>"11111110",
  2664=>"00000000",
  2665=>"00000001",
  2666=>"00000000",
  2667=>"11111111",
  2668=>"00000000",
  2669=>"00000000",
  2670=>"00000000",
  2671=>"00000000",
  2672=>"00000000",
  2673=>"00000000",
  2674=>"00000001",
  2675=>"00000000",
  2676=>"00000000",
  2677=>"00000000",
  2678=>"11111111",
  2679=>"00000000",
  2680=>"00000001",
  2681=>"00000000",
  2682=>"11111111",
  2683=>"00000000",
  2684=>"00000000",
  2685=>"00000000",
  2686=>"00000001",
  2687=>"11111111",
  2688=>"00000000",
  2689=>"00000000",
  2690=>"00000000",
  2691=>"00000000",
  2692=>"00000000",
  2693=>"00000000",
  2694=>"11111111",
  2695=>"00000000",
  2696=>"00000001",
  2697=>"00000000",
  2698=>"00000001",
  2699=>"11111111",
  2700=>"00000000",
  2701=>"00000000",
  2702=>"00000000",
  2703=>"00000001",
  2704=>"00000000",
  2705=>"00000000",
  2706=>"00000000",
  2707=>"11111111",
  2708=>"00000000",
  2709=>"00000000",
  2710=>"11111111",
  2711=>"00000001",
  2712=>"00000000",
  2713=>"00000000",
  2714=>"11111111",
  2715=>"00000001",
  2716=>"00000000",
  2717=>"00000000",
  2718=>"00000000",
  2719=>"00000000",
  2720=>"11111110",
  2721=>"00000000",
  2722=>"00000000",
  2723=>"00000000",
  2724=>"00000000",
  2725=>"00000000",
  2726=>"00000000",
  2727=>"00000000",
  2728=>"11111111",
  2729=>"00000000",
  2730=>"00000000",
  2731=>"00000000",
  2732=>"00000000",
  2733=>"00000000",
  2734=>"00000000",
  2735=>"00000000",
  2736=>"00000000",
  2737=>"11111111",
  2738=>"00000000",
  2739=>"00000000",
  2740=>"00000001",
  2741=>"11111111",
  2742=>"00000000",
  2743=>"00000001",
  2744=>"00000000",
  2745=>"11111101",
  2746=>"00000000",
  2747=>"00000000",
  2748=>"00000000",
  2749=>"00000001",
  2750=>"00000000",
  2751=>"11111111",
  2752=>"00000000",
  2753=>"00000001",
  2754=>"11111111",
  2755=>"00000000",
  2756=>"00000000",
  2757=>"11111111",
  2758=>"00000001",
  2759=>"00000000",
  2760=>"00000001",
  2761=>"00000000",
  2762=>"11111111",
  2763=>"00000000",
  2764=>"00000000",
  2765=>"00000001",
  2766=>"00000000",
  2767=>"00000000",
  2768=>"00000010",
  2769=>"00000001",
  2770=>"00000001",
  2771=>"00000001",
  2772=>"11111111",
  2773=>"00000000",
  2774=>"11111111",
  2775=>"11111111",
  2776=>"00000010",
  2777=>"11111111",
  2778=>"11111111",
  2779=>"00000000",
  2780=>"00000000",
  2781=>"11111111",
  2782=>"00000000",
  2783=>"00000000",
  2784=>"00000000",
  2785=>"00000000",
  2786=>"00000001",
  2787=>"00000000",
  2788=>"00000000",
  2789=>"00000000",
  2790=>"11111111",
  2791=>"11111111",
  2792=>"11111111",
  2793=>"00000000",
  2794=>"11111111",
  2795=>"00000000",
  2796=>"00000101",
  2797=>"00000001",
  2798=>"00000001",
  2799=>"00000000",
  2800=>"00000000",
  2801=>"00000001",
  2802=>"00000000",
  2803=>"00000000",
  2804=>"00000000",
  2805=>"00000000",
  2806=>"00000000",
  2807=>"00000000",
  2808=>"00000000",
  2809=>"00000000",
  2810=>"00000000",
  2811=>"00000000",
  2812=>"00000000",
  2813=>"00000000",
  2814=>"00000000",
  2815=>"00000000",
  2816=>"00000000",
  2817=>"00000000",
  2818=>"00000000",
  2819=>"00000001",
  2820=>"00000000",
  2821=>"11111111",
  2822=>"00000000",
  2823=>"00000001",
  2824=>"00000000",
  2825=>"00000010",
  2826=>"00000000",
  2827=>"00000000",
  2828=>"00000001",
  2829=>"00000000",
  2830=>"00000000",
  2831=>"00000000",
  2832=>"11111111",
  2833=>"00000001",
  2834=>"11111111",
  2835=>"00000000",
  2836=>"11111111",
  2837=>"00000001",
  2838=>"11111111",
  2839=>"00000001",
  2840=>"00000001",
  2841=>"11111111",
  2842=>"00000000",
  2843=>"00000000",
  2844=>"11111111",
  2845=>"00000000",
  2846=>"00000000",
  2847=>"00000000",
  2848=>"00000000",
  2849=>"00000000",
  2850=>"00000000",
  2851=>"00000000",
  2852=>"11111110",
  2853=>"00000000",
  2854=>"00000000",
  2855=>"00000000",
  2856=>"11111111",
  2857=>"00000000",
  2858=>"00000000",
  2859=>"00000000",
  2860=>"11111110",
  2861=>"00000000",
  2862=>"00000000",
  2863=>"00000000",
  2864=>"00000001",
  2865=>"00000001",
  2866=>"00000001",
  2867=>"00000000",
  2868=>"00000000",
  2869=>"00000000",
  2870=>"00000001",
  2871=>"00000000",
  2872=>"11111111",
  2873=>"00000000",
  2874=>"00000001",
  2875=>"00000001",
  2876=>"00000000",
  2877=>"00000000",
  2878=>"00000000",
  2879=>"00000010",
  2880=>"00000001",
  2881=>"00000001",
  2882=>"00000001",
  2883=>"00000000",
  2884=>"00000000",
  2885=>"00000000",
  2886=>"00000000",
  2887=>"00000000",
  2888=>"00000001",
  2889=>"00000001",
  2890=>"00000000",
  2891=>"00000001",
  2892=>"11111111",
  2893=>"00000000",
  2894=>"00000000",
  2895=>"00000001",
  2896=>"11111111",
  2897=>"11111111",
  2898=>"00000000",
  2899=>"00000000",
  2900=>"00000000",
  2901=>"11111111",
  2902=>"11111111",
  2903=>"00000000",
  2904=>"00000000",
  2905=>"00000000",
  2906=>"00000001",
  2907=>"00000000",
  2908=>"00000000",
  2909=>"00000000",
  2910=>"00000000",
  2911=>"00000000",
  2912=>"00000001",
  2913=>"00000000",
  2914=>"11111111",
  2915=>"00000001",
  2916=>"00000000",
  2917=>"00000000",
  2918=>"00000001",
  2919=>"11111111",
  2920=>"00000000",
  2921=>"00000000",
  2922=>"00000001",
  2923=>"00000000",
  2924=>"11111111",
  2925=>"00000000",
  2926=>"00000000",
  2927=>"00000000",
  2928=>"00000000",
  2929=>"11111111",
  2930=>"11111111",
  2931=>"00000000",
  2932=>"11111111",
  2933=>"00000000",
  2934=>"00000001",
  2935=>"00000100",
  2936=>"11111111",
  2937=>"00000000",
  2938=>"00000000",
  2939=>"00000000",
  2940=>"00000000",
  2941=>"00000000",
  2942=>"00000000",
  2943=>"00000000",
  2944=>"00000010",
  2945=>"00000000",
  2946=>"00000001",
  2947=>"00000000",
  2948=>"00000000",
  2949=>"11111111",
  2950=>"00000000",
  2951=>"00000000",
  2952=>"00000001",
  2953=>"00000001",
  2954=>"11111110",
  2955=>"00000010",
  2956=>"00000001",
  2957=>"00000001",
  2958=>"00000000",
  2959=>"11111111",
  2960=>"11111111",
  2961=>"00000000",
  2962=>"00000000",
  2963=>"11111111",
  2964=>"00000000",
  2965=>"00000001",
  2966=>"11111101",
  2967=>"11111111",
  2968=>"00000000",
  2969=>"00000000",
  2970=>"11111111",
  2971=>"00000001",
  2972=>"11111111",
  2973=>"00000000",
  2974=>"00000000",
  2975=>"00000001",
  2976=>"00000000",
  2977=>"00000010",
  2978=>"00000000",
  2979=>"00000000",
  2980=>"00000000",
  2981=>"00000000",
  2982=>"00000001",
  2983=>"00000000",
  2984=>"00000000",
  2985=>"00000000",
  2986=>"11111111",
  2987=>"11111111",
  2988=>"00000000",
  2989=>"00000000",
  2990=>"00000000",
  2991=>"00000000",
  2992=>"00000000",
  2993=>"11111111",
  2994=>"00000000",
  2995=>"11111111",
  2996=>"00000000",
  2997=>"00000000",
  2998=>"00000000",
  2999=>"00000000",
  3000=>"00000000",
  3001=>"00000000",
  3002=>"11111111",
  3003=>"00000000",
  3004=>"00000000",
  3005=>"00000000",
  3006=>"00000001",
  3007=>"11111110",
  3008=>"00000000",
  3009=>"00000001",
  3010=>"00000000",
  3011=>"00000000",
  3012=>"00000000",
  3013=>"00000000",
  3014=>"11111111",
  3015=>"11111101",
  3016=>"00000000",
  3017=>"00000000",
  3018=>"00000000",
  3019=>"00000000",
  3020=>"00000001",
  3021=>"00000000",
  3022=>"00000000",
  3023=>"00000001",
  3024=>"00000000",
  3025=>"00000000",
  3026=>"00000000",
  3027=>"00000001",
  3028=>"11111111",
  3029=>"00000000",
  3030=>"00000000",
  3031=>"00000001",
  3032=>"11111111",
  3033=>"00000000",
  3034=>"00000010",
  3035=>"00000001",
  3036=>"11111111",
  3037=>"00000000",
  3038=>"11111110",
  3039=>"00000000",
  3040=>"00000001",
  3041=>"00000000",
  3042=>"00000000",
  3043=>"11111110",
  3044=>"00000000",
  3045=>"00000000",
  3046=>"00000000",
  3047=>"00000000",
  3048=>"00000001",
  3049=>"00000001",
  3050=>"00000001",
  3051=>"00000000",
  3052=>"00000001",
  3053=>"11111111",
  3054=>"00000000",
  3055=>"00000001",
  3056=>"00000000",
  3057=>"00000000",
  3058=>"11111111",
  3059=>"00000000",
  3060=>"11111111",
  3061=>"00000000",
  3062=>"00000001",
  3063=>"00000000",
  3064=>"00000000",
  3065=>"00000000",
  3066=>"00000000",
  3067=>"00000000",
  3068=>"11111111",
  3069=>"00000000",
  3070=>"00000000",
  3071=>"11111111",
  3072=>"00000010",
  3073=>"00000001",
  3074=>"00000000",
  3075=>"11111111",
  3076=>"11111111",
  3077=>"00000000",
  3078=>"00000000",
  3079=>"11111111",
  3080=>"00000000",
  3081=>"00000000",
  3082=>"00000000",
  3083=>"00000000",
  3084=>"00000000",
  3085=>"00000000",
  3086=>"00000000",
  3087=>"00000001",
  3088=>"11111111",
  3089=>"00000000",
  3090=>"00000000",
  3091=>"00000000",
  3092=>"11111111",
  3093=>"11111111",
  3094=>"00000000",
  3095=>"00000000",
  3096=>"00000000",
  3097=>"11111111",
  3098=>"00000001",
  3099=>"00000010",
  3100=>"00000000",
  3101=>"00000000",
  3102=>"00000000",
  3103=>"00000000",
  3104=>"00000000",
  3105=>"00000000",
  3106=>"00000000",
  3107=>"11111111",
  3108=>"00000001",
  3109=>"00000000",
  3110=>"00000000",
  3111=>"00000000",
  3112=>"11111111",
  3113=>"00000000",
  3114=>"00000000",
  3115=>"00000000",
  3116=>"11111110",
  3117=>"00000000",
  3118=>"00000001",
  3119=>"11111111",
  3120=>"11111111",
  3121=>"11111110",
  3122=>"00000000",
  3123=>"11111111",
  3124=>"00000000",
  3125=>"00000001",
  3126=>"11111110",
  3127=>"00000001",
  3128=>"00000000",
  3129=>"00000001",
  3130=>"00000001",
  3131=>"00000001",
  3132=>"00000000",
  3133=>"00000000",
  3134=>"00000000",
  3135=>"00000000",
  3136=>"00000000",
  3137=>"00000000",
  3138=>"00000000",
  3139=>"00000000",
  3140=>"00000000",
  3141=>"00000001",
  3142=>"00000001",
  3143=>"00000001",
  3144=>"00000000",
  3145=>"00000000",
  3146=>"00000011",
  3147=>"11111111",
  3148=>"00000001",
  3149=>"00000001",
  3150=>"11111111",
  3151=>"00000000",
  3152=>"00000000",
  3153=>"00000001",
  3154=>"00000000",
  3155=>"00000000",
  3156=>"00000000",
  3157=>"11111111",
  3158=>"00000000",
  3159=>"00000000",
  3160=>"00000000",
  3161=>"00000001",
  3162=>"00000000",
  3163=>"00000000",
  3164=>"00000000",
  3165=>"00000001",
  3166=>"00000000",
  3167=>"00000000",
  3168=>"11111111",
  3169=>"00000000",
  3170=>"00000000",
  3171=>"11111111",
  3172=>"00000001",
  3173=>"11111111",
  3174=>"00000010",
  3175=>"11111111",
  3176=>"00000001",
  3177=>"00000001",
  3178=>"00000000",
  3179=>"00000001",
  3180=>"00000000",
  3181=>"00000000",
  3182=>"00000010",
  3183=>"00000000",
  3184=>"00000001",
  3185=>"00000000",
  3186=>"00000001",
  3187=>"00000000",
  3188=>"11111111",
  3189=>"00000001",
  3190=>"00000000",
  3191=>"00000000",
  3192=>"00000000",
  3193=>"00000000",
  3194=>"00000001",
  3195=>"00000000",
  3196=>"11111111",
  3197=>"00000001",
  3198=>"11111101",
  3199=>"00000000",
  3200=>"11111111",
  3201=>"00000000",
  3202=>"00000000",
  3203=>"00000000",
  3204=>"00000000",
  3205=>"11111111",
  3206=>"11111111",
  3207=>"00000000",
  3208=>"00000000",
  3209=>"00000000",
  3210=>"00000001",
  3211=>"00000000",
  3212=>"00000000",
  3213=>"00000001",
  3214=>"00000000",
  3215=>"00000000",
  3216=>"00000000",
  3217=>"00000000",
  3218=>"00000000",
  3219=>"00000000",
  3220=>"11111111",
  3221=>"00000000",
  3222=>"00000000",
  3223=>"11111111",
  3224=>"00000000",
  3225=>"00000000",
  3226=>"00000000",
  3227=>"00000001",
  3228=>"11111110",
  3229=>"00000001",
  3230=>"11111111",
  3231=>"00000000",
  3232=>"00000000",
  3233=>"00000000",
  3234=>"00000000",
  3235=>"00000001",
  3236=>"11111110",
  3237=>"00000000",
  3238=>"00000000",
  3239=>"00000000",
  3240=>"00000000",
  3241=>"00000000",
  3242=>"11111111",
  3243=>"00000000",
  3244=>"00000000",
  3245=>"00000000",
  3246=>"00000000",
  3247=>"00000001",
  3248=>"11111111",
  3249=>"11111111",
  3250=>"00000001",
  3251=>"00000001",
  3252=>"00000000",
  3253=>"00000000",
  3254=>"00000000",
  3255=>"00000001",
  3256=>"00000000",
  3257=>"00000000",
  3258=>"00000000",
  3259=>"00000001",
  3260=>"11111111",
  3261=>"11111110",
  3262=>"00000000",
  3263=>"00000000",
  3264=>"00000001",
  3265=>"00000000",
  3266=>"00000000",
  3267=>"00000000",
  3268=>"00000001",
  3269=>"00000000",
  3270=>"00000000",
  3271=>"00000001",
  3272=>"00000000",
  3273=>"11111111",
  3274=>"00000000",
  3275=>"00000000",
  3276=>"00000000",
  3277=>"00000000",
  3278=>"00000000",
  3279=>"00000000",
  3280=>"00000001",
  3281=>"00000000",
  3282=>"00000010",
  3283=>"11111110",
  3284=>"00000001",
  3285=>"00000000",
  3286=>"00000000",
  3287=>"00000000",
  3288=>"11111111",
  3289=>"00000001",
  3290=>"11111111",
  3291=>"00000000",
  3292=>"00000000",
  3293=>"00000000",
  3294=>"11111111",
  3295=>"00000001",
  3296=>"00000001",
  3297=>"00000000",
  3298=>"00000000",
  3299=>"00000001",
  3300=>"00000001",
  3301=>"00000001",
  3302=>"00000000",
  3303=>"00000000",
  3304=>"11111111",
  3305=>"11111111",
  3306=>"00000000",
  3307=>"00000000",
  3308=>"11111101",
  3309=>"00000000",
  3310=>"00000001",
  3311=>"11111100",
  3312=>"00000001",
  3313=>"00000001",
  3314=>"00000001",
  3315=>"00000000",
  3316=>"00000000",
  3317=>"00000001",
  3318=>"00000001",
  3319=>"11111111",
  3320=>"00000000",
  3321=>"00000100",
  3322=>"00000001",
  3323=>"00000000",
  3324=>"11111111",
  3325=>"00000000",
  3326=>"00000000",
  3327=>"11111111",
  3328=>"11111111",
  3329=>"00000000",
  3330=>"11111111",
  3331=>"00000000",
  3332=>"00000000",
  3333=>"00000001",
  3334=>"00000000",
  3335=>"00000000",
  3336=>"11111111",
  3337=>"00000000",
  3338=>"00000000",
  3339=>"11111111",
  3340=>"11111101",
  3341=>"00000000",
  3342=>"00000000",
  3343=>"00000000",
  3344=>"00000000",
  3345=>"00000000",
  3346=>"11111111",
  3347=>"00000001",
  3348=>"00000001",
  3349=>"00000001",
  3350=>"00000000",
  3351=>"00000001",
  3352=>"00000000",
  3353=>"00000001",
  3354=>"00000000",
  3355=>"11111110",
  3356=>"00000000",
  3357=>"00000001",
  3358=>"00000000",
  3359=>"00000000",
  3360=>"00000001",
  3361=>"11111110",
  3362=>"00000000",
  3363=>"00000000",
  3364=>"00000001",
  3365=>"00000001",
  3366=>"00000000",
  3367=>"00000000",
  3368=>"00000000",
  3369=>"00000000",
  3370=>"00000000",
  3371=>"00000001",
  3372=>"00000000",
  3373=>"11111111",
  3374=>"00000000",
  3375=>"00000000",
  3376=>"00000000",
  3377=>"00000001",
  3378=>"00000000",
  3379=>"00000000",
  3380=>"00000000",
  3381=>"00000000",
  3382=>"00000000",
  3383=>"00000000",
  3384=>"00000000",
  3385=>"00000000",
  3386=>"00000001",
  3387=>"11111111",
  3388=>"00000000",
  3389=>"00000000",
  3390=>"00000000",
  3391=>"11111110",
  3392=>"00000000",
  3393=>"00000000",
  3394=>"00000000",
  3395=>"00000000",
  3396=>"00000001",
  3397=>"00000000",
  3398=>"00000000",
  3399=>"11111111",
  3400=>"00000001",
  3401=>"00000000",
  3402=>"00000000",
  3403=>"11111111",
  3404=>"11111111",
  3405=>"00000000",
  3406=>"00000001",
  3407=>"00000000",
  3408=>"00000000",
  3409=>"00000000",
  3410=>"00000000",
  3411=>"00000000",
  3412=>"11111110",
  3413=>"00000000",
  3414=>"00000000",
  3415=>"00000000",
  3416=>"00000001",
  3417=>"00000000",
  3418=>"00000000",
  3419=>"11111111",
  3420=>"11111111",
  3421=>"11111111",
  3422=>"00000000",
  3423=>"00000000",
  3424=>"00000000",
  3425=>"11111111",
  3426=>"00000001",
  3427=>"11111111",
  3428=>"00000001",
  3429=>"00000000",
  3430=>"00000000",
  3431=>"00000000",
  3432=>"00000001",
  3433=>"00000000",
  3434=>"00000000",
  3435=>"00000000",
  3436=>"00000000",
  3437=>"00000000",
  3438=>"00000000",
  3439=>"00000000",
  3440=>"00000011",
  3441=>"00000000",
  3442=>"11111111",
  3443=>"00000000",
  3444=>"00000000",
  3445=>"00000000",
  3446=>"00000000",
  3447=>"00000000",
  3448=>"00000000",
  3449=>"00000000",
  3450=>"00000000",
  3451=>"00000000",
  3452=>"00000001",
  3453=>"00000000",
  3454=>"00000001",
  3455=>"00000000",
  3456=>"00000000",
  3457=>"00000000",
  3458=>"00000001",
  3459=>"00000001",
  3460=>"00000000",
  3461=>"00000000",
  3462=>"00000000",
  3463=>"00000010",
  3464=>"00000000",
  3465=>"00000010",
  3466=>"00000001",
  3467=>"00000000",
  3468=>"11111111",
  3469=>"00000000",
  3470=>"00000000",
  3471=>"00000000",
  3472=>"11111111",
  3473=>"00000000",
  3474=>"00000000",
  3475=>"00000001",
  3476=>"00000000",
  3477=>"00000001",
  3478=>"00000001",
  3479=>"00000000",
  3480=>"00000001",
  3481=>"00000000",
  3482=>"00000000",
  3483=>"00000000",
  3484=>"00000000",
  3485=>"00000001",
  3486=>"00000000",
  3487=>"00000000",
  3488=>"00000000",
  3489=>"00000000",
  3490=>"00000000",
  3491=>"00000000",
  3492=>"00000000",
  3493=>"00000001",
  3494=>"11111111",
  3495=>"00000000",
  3496=>"00000000",
  3497=>"00000001",
  3498=>"00000001",
  3499=>"00000000",
  3500=>"11111111",
  3501=>"00000001",
  3502=>"00000010",
  3503=>"00000000",
  3504=>"00000001",
  3505=>"00000000",
  3506=>"00000000",
  3507=>"00000000",
  3508=>"00000000",
  3509=>"00000000",
  3510=>"00000000",
  3511=>"00000000",
  3512=>"00000000",
  3513=>"00000001",
  3514=>"00000000",
  3515=>"00000000",
  3516=>"11111101",
  3517=>"00000001",
  3518=>"00000000",
  3519=>"11111111",
  3520=>"00000000",
  3521=>"00000000",
  3522=>"00000000",
  3523=>"00000001",
  3524=>"00000000",
  3525=>"00000000",
  3526=>"00000000",
  3527=>"00000000",
  3528=>"00000000",
  3529=>"00000000",
  3530=>"11111111",
  3531=>"00000000",
  3532=>"00000000",
  3533=>"11111110",
  3534=>"00000000",
  3535=>"00000000",
  3536=>"11111111",
  3537=>"11111110",
  3538=>"11111110",
  3539=>"00000001",
  3540=>"11111111",
  3541=>"00000001",
  3542=>"00000000",
  3543=>"00000000",
  3544=>"00000000",
  3545=>"00000000",
  3546=>"00000000",
  3547=>"00000000",
  3548=>"00000000",
  3549=>"00000010",
  3550=>"00000000",
  3551=>"00000001",
  3552=>"00000000",
  3553=>"00000000",
  3554=>"11111111",
  3555=>"00000001",
  3556=>"00000000",
  3557=>"00000000",
  3558=>"00000000",
  3559=>"00000010",
  3560=>"00000000",
  3561=>"00000000",
  3562=>"00000000",
  3563=>"00000000",
  3564=>"00000001",
  3565=>"00000000",
  3566=>"00000000",
  3567=>"00000000",
  3568=>"00000000",
  3569=>"00000000",
  3570=>"00000001",
  3571=>"00000000",
  3572=>"00000001",
  3573=>"00000000",
  3574=>"11111111",
  3575=>"00000000",
  3576=>"00000000",
  3577=>"00000000",
  3578=>"11111111",
  3579=>"00000000",
  3580=>"00000000",
  3581=>"00000001",
  3582=>"00000000",
  3583=>"11111111",
  3584=>"00000010",
  3585=>"00000000",
  3586=>"00000001",
  3587=>"00000000",
  3588=>"00000000",
  3589=>"00000000",
  3590=>"00000000",
  3591=>"11111111",
  3592=>"00000000",
  3593=>"00000000",
  3594=>"11111111",
  3595=>"11111111",
  3596=>"00000000",
  3597=>"11111111",
  3598=>"00000000",
  3599=>"00000000",
  3600=>"00000000",
  3601=>"00000000",
  3602=>"00000000",
  3603=>"00000000",
  3604=>"00000000",
  3605=>"00000001",
  3606=>"11111110",
  3607=>"00000000",
  3608=>"00000001",
  3609=>"00000000",
  3610=>"11111111",
  3611=>"00000000",
  3612=>"11111110",
  3613=>"00000000",
  3614=>"00000000",
  3615=>"11111111",
  3616=>"00000000",
  3617=>"00000000",
  3618=>"00000001",
  3619=>"11111111",
  3620=>"00000000",
  3621=>"11111111",
  3622=>"11111111",
  3623=>"00000000",
  3624=>"00000001",
  3625=>"11111111",
  3626=>"00000000",
  3627=>"00000000",
  3628=>"00000000",
  3629=>"00000000",
  3630=>"00000001",
  3631=>"00000000",
  3632=>"00000000",
  3633=>"11111111",
  3634=>"11111111",
  3635=>"00000001",
  3636=>"00000000",
  3637=>"11111111",
  3638=>"00000001",
  3639=>"00000000",
  3640=>"00000000",
  3641=>"00000000",
  3642=>"00000000",
  3643=>"00000000",
  3644=>"00000000",
  3645=>"00000000",
  3646=>"00000000",
  3647=>"00000000",
  3648=>"11111111",
  3649=>"00000000",
  3650=>"00000001",
  3651=>"00000001",
  3652=>"11111111",
  3653=>"11111110",
  3654=>"00000001",
  3655=>"00000000",
  3656=>"00000001",
  3657=>"00000000",
  3658=>"00000001",
  3659=>"00000000",
  3660=>"11111111",
  3661=>"00000000",
  3662=>"00000000",
  3663=>"00000000",
  3664=>"00000000",
  3665=>"00000000",
  3666=>"00000000",
  3667=>"00000000",
  3668=>"00000000",
  3669=>"00000000",
  3670=>"00000000",
  3671=>"00000000",
  3672=>"00000000",
  3673=>"11111111",
  3674=>"00000000",
  3675=>"11111111",
  3676=>"00000001",
  3677=>"11111111",
  3678=>"00000001",
  3679=>"00000000",
  3680=>"00000000",
  3681=>"00000000",
  3682=>"00000000",
  3683=>"00000001",
  3684=>"00000001",
  3685=>"11111111",
  3686=>"00000001",
  3687=>"00000000",
  3688=>"00000000",
  3689=>"00000010",
  3690=>"11111111",
  3691=>"11111101",
  3692=>"00000000",
  3693=>"00000000",
  3694=>"11111111",
  3695=>"00000000",
  3696=>"00000001",
  3697=>"11111111",
  3698=>"00000000",
  3699=>"00000000",
  3700=>"00000001",
  3701=>"00000000",
  3702=>"00000000",
  3703=>"00000000",
  3704=>"00000000",
  3705=>"00000000",
  3706=>"00000000",
  3707=>"00000000",
  3708=>"00000000",
  3709=>"00000000",
  3710=>"11111111",
  3711=>"00000001",
  3712=>"00000001",
  3713=>"00000000",
  3714=>"00000000",
  3715=>"00000000",
  3716=>"00000000",
  3717=>"00000000",
  3718=>"00000000",
  3719=>"00000000",
  3720=>"00000001",
  3721=>"11111111",
  3722=>"00000000",
  3723=>"00000000",
  3724=>"00000001",
  3725=>"00000000",
  3726=>"00000001",
  3727=>"00000001",
  3728=>"00000000",
  3729=>"00000000",
  3730=>"00000000",
  3731=>"11111101",
  3732=>"00000000",
  3733=>"00000000",
  3734=>"00000001",
  3735=>"00000000",
  3736=>"11111111",
  3737=>"00000000",
  3738=>"00000001",
  3739=>"00000000",
  3740=>"00000000",
  3741=>"00000000",
  3742=>"00000001",
  3743=>"00000001",
  3744=>"00000010",
  3745=>"00000000",
  3746=>"00000000",
  3747=>"00000001",
  3748=>"00000000",
  3749=>"00000000",
  3750=>"00000001",
  3751=>"00000001",
  3752=>"00000000",
  3753=>"11111111",
  3754=>"00000000",
  3755=>"00000000",
  3756=>"00000000",
  3757=>"00000000",
  3758=>"00000000",
  3759=>"00000000",
  3760=>"11111111",
  3761=>"11111111",
  3762=>"11111111",
  3763=>"00000000",
  3764=>"00000000",
  3765=>"00000000",
  3766=>"00000000",
  3767=>"00000001",
  3768=>"00000000",
  3769=>"00000001",
  3770=>"00000001",
  3771=>"00000000",
  3772=>"00000000",
  3773=>"00000000",
  3774=>"00000000",
  3775=>"00000000",
  3776=>"00000000",
  3777=>"00000000",
  3778=>"11111111",
  3779=>"00000000",
  3780=>"00000001",
  3781=>"00000000",
  3782=>"00000001",
  3783=>"00000000",
  3784=>"00000010",
  3785=>"11111111",
  3786=>"00000000",
  3787=>"11111111",
  3788=>"00000000",
  3789=>"00000001",
  3790=>"00000001",
  3791=>"00000000",
  3792=>"11111101",
  3793=>"00000000",
  3794=>"00000001",
  3795=>"00000001",
  3796=>"11111111",
  3797=>"00000000",
  3798=>"00000000",
  3799=>"11111111",
  3800=>"00000000",
  3801=>"11111111",
  3802=>"11111111",
  3803=>"00000000",
  3804=>"11111111",
  3805=>"00000000",
  3806=>"00000000",
  3807=>"00000000",
  3808=>"00000000",
  3809=>"00000001",
  3810=>"00000000",
  3811=>"00000000",
  3812=>"00000000",
  3813=>"11111111",
  3814=>"00000000",
  3815=>"00000001",
  3816=>"00000000",
  3817=>"00000000",
  3818=>"11111111",
  3819=>"11111111",
  3820=>"11111110",
  3821=>"00000000",
  3822=>"00000000",
  3823=>"00000000",
  3824=>"00000000",
  3825=>"00000000",
  3826=>"00000000",
  3827=>"00000000",
  3828=>"00000000",
  3829=>"00000000",
  3830=>"11111111",
  3831=>"11111111",
  3832=>"00000001",
  3833=>"11111111",
  3834=>"00000000",
  3835=>"00000000",
  3836=>"11111111",
  3837=>"00000000",
  3838=>"00000000",
  3839=>"00000000",
  3840=>"00000000",
  3841=>"00000001",
  3842=>"00000000",
  3843=>"00000000",
  3844=>"00000000",
  3845=>"00000001",
  3846=>"00000000",
  3847=>"00000000",
  3848=>"00000000",
  3849=>"00000000",
  3850=>"00000000",
  3851=>"00000000",
  3852=>"00000000",
  3853=>"11111111",
  3854=>"00000000",
  3855=>"11111101",
  3856=>"00000001",
  3857=>"11111111",
  3858=>"00000001",
  3859=>"00000000",
  3860=>"00000000",
  3861=>"00000001",
  3862=>"00000000",
  3863=>"00000000",
  3864=>"00000000",
  3865=>"00000000",
  3866=>"00000000",
  3867=>"00000000",
  3868=>"11111111",
  3869=>"00000000",
  3870=>"00000000",
  3871=>"00000000",
  3872=>"00000000",
  3873=>"00000001",
  3874=>"00000000",
  3875=>"00000000",
  3876=>"00000000",
  3877=>"00000000",
  3878=>"11111111",
  3879=>"11111111",
  3880=>"00000000",
  3881=>"00000000",
  3882=>"11111111",
  3883=>"00000000",
  3884=>"11111111",
  3885=>"00000000",
  3886=>"00000000",
  3887=>"00000001",
  3888=>"11111111",
  3889=>"00000001",
  3890=>"00000000",
  3891=>"00000000",
  3892=>"00000000",
  3893=>"00000000",
  3894=>"00000000",
  3895=>"00000000",
  3896=>"00000001",
  3897=>"11111111",
  3898=>"00000000",
  3899=>"00000000",
  3900=>"11111111",
  3901=>"00000001",
  3902=>"00000000",
  3903=>"00000000",
  3904=>"00000000",
  3905=>"11111111",
  3906=>"00000000",
  3907=>"00000000",
  3908=>"00000000",
  3909=>"00000000",
  3910=>"00000001",
  3911=>"00000000",
  3912=>"00000001",
  3913=>"00000000",
  3914=>"00000000",
  3915=>"00000000",
  3916=>"11111111",
  3917=>"00000000",
  3918=>"00000000",
  3919=>"00000000",
  3920=>"00000010",
  3921=>"11111111",
  3922=>"00000000",
  3923=>"11111111",
  3924=>"00000001",
  3925=>"00000000",
  3926=>"00000001",
  3927=>"00000000",
  3928=>"00000000",
  3929=>"00000001",
  3930=>"00000000",
  3931=>"00000000",
  3932=>"00000001",
  3933=>"00000000",
  3934=>"00000000",
  3935=>"00000000",
  3936=>"00000000",
  3937=>"00000000",
  3938=>"00000000",
  3939=>"00000000",
  3940=>"11111111",
  3941=>"00000000",
  3942=>"11111111",
  3943=>"00000000",
  3944=>"00000000",
  3945=>"00000001",
  3946=>"11111111",
  3947=>"00000001",
  3948=>"00000001",
  3949=>"00000000",
  3950=>"11111110",
  3951=>"00000000",
  3952=>"00000000",
  3953=>"00000000",
  3954=>"00000000",
  3955=>"00000000",
  3956=>"00000000",
  3957=>"00000000",
  3958=>"00000000",
  3959=>"11111110",
  3960=>"00000000",
  3961=>"00000001",
  3962=>"00000000",
  3963=>"00000001",
  3964=>"00000000",
  3965=>"00000000",
  3966=>"00000000",
  3967=>"00000000",
  3968=>"11111110",
  3969=>"00000000",
  3970=>"00000000",
  3971=>"00000000",
  3972=>"00000001",
  3973=>"00000000",
  3974=>"00000000",
  3975=>"00000000",
  3976=>"00000001",
  3977=>"11111111",
  3978=>"11111111",
  3979=>"00000001",
  3980=>"11111111",
  3981=>"11111111",
  3982=>"00000000",
  3983=>"11111111",
  3984=>"00000000",
  3985=>"00000000",
  3986=>"00000000",
  3987=>"00000000",
  3988=>"00000000",
  3989=>"00000000",
  3990=>"11111110",
  3991=>"00000000",
  3992=>"00000001",
  3993=>"00000000",
  3994=>"00000000",
  3995=>"00000000",
  3996=>"00000000",
  3997=>"00000000",
  3998=>"00000000",
  3999=>"00000001",
  4000=>"00000000",
  4001=>"00000001",
  4002=>"00000000",
  4003=>"00000000",
  4004=>"00000000",
  4005=>"00000001",
  4006=>"00000001",
  4007=>"00000000",
  4008=>"00000000",
  4009=>"00000000",
  4010=>"00000000",
  4011=>"00000000",
  4012=>"00000001",
  4013=>"11111111",
  4014=>"00000000",
  4015=>"11111111",
  4016=>"11111111",
  4017=>"00000000",
  4018=>"00000000",
  4019=>"00000001",
  4020=>"00000000",
  4021=>"00000000",
  4022=>"00000000",
  4023=>"11111111",
  4024=>"00000000",
  4025=>"00000000",
  4026=>"00000001",
  4027=>"11111111",
  4028=>"00000000",
  4029=>"00000000",
  4030=>"11111101",
  4031=>"00000000",
  4032=>"00000000",
  4033=>"00000000",
  4034=>"00000000",
  4035=>"00000000",
  4036=>"00000000",
  4037=>"00000000",
  4038=>"11111111",
  4039=>"11111100",
  4040=>"00000000",
  4041=>"00000000",
  4042=>"00000001",
  4043=>"00000000",
  4044=>"00000000",
  4045=>"00000000",
  4046=>"00000001",
  4047=>"00000000",
  4048=>"11111111",
  4049=>"00000000",
  4050=>"00000000",
  4051=>"00000000",
  4052=>"00000000",
  4053=>"00000000",
  4054=>"00000000",
  4055=>"00000001",
  4056=>"11111111",
  4057=>"00000000",
  4058=>"00000000",
  4059=>"00000001",
  4060=>"00000000",
  4061=>"00000000",
  4062=>"11111111",
  4063=>"00000001",
  4064=>"11111111",
  4065=>"00000001",
  4066=>"00000001",
  4067=>"00000001",
  4068=>"00000000",
  4069=>"00000000",
  4070=>"00000000",
  4071=>"00000000",
  4072=>"11111111",
  4073=>"00000000",
  4074=>"00000000",
  4075=>"00000000",
  4076=>"00000000",
  4077=>"00000001",
  4078=>"00000000",
  4079=>"00000000",
  4080=>"00000000",
  4081=>"00000010",
  4082=>"00000000",
  4083=>"00000001",
  4084=>"00000000",
  4085=>"00000000",
  4086=>"00000001",
  4087=>"00000000",
  4088=>"11111111",
  4089=>"11111111",
  4090=>"00000000",
  4091=>"00000000",
  4092=>"00000000",
  4093=>"00000000",
  4094=>"00000000",
  4095=>"00000000",
  4096=>"11111101",
  4097=>"00000000",
  4098=>"11111100",
  4099=>"11111110",
  4100=>"11111110",
  4101=>"00000010",
  4102=>"00000000",
  4103=>"00000010",
  4104=>"11111100",
  4105=>"00000001",
  4106=>"11111110",
  4107=>"11111111",
  4108=>"00000010",
  4109=>"11111111",
  4110=>"11111101",
  4111=>"00000001",
  4112=>"11111111",
  4113=>"11111011",
  4114=>"00000001",
  4115=>"11111110",
  4116=>"00000011",
  4117=>"11111110",
  4118=>"00000001",
  4119=>"11111110",
  4120=>"00000001",
  4121=>"11111110",
  4122=>"00000010",
  4123=>"11111011",
  4124=>"00000000",
  4125=>"11111101",
  4126=>"00000010",
  4127=>"11111101",
  4128=>"11111111",
  4129=>"11111110",
  4130=>"00000000",
  4131=>"11111111",
  4132=>"00000001",
  4133=>"11111110",
  4134=>"11111111",
  4135=>"11111001",
  4136=>"11111110",
  4137=>"00000001",
  4138=>"11111110",
  4139=>"11111110",
  4140=>"11111011",
  4141=>"00000001",
  4142=>"00000001",
  4143=>"11111111",
  4144=>"11111001",
  4145=>"00000000",
  4146=>"11111100",
  4147=>"00000010",
  4148=>"11111011",
  4149=>"11111010",
  4150=>"11111101",
  4151=>"00000011",
  4152=>"00000000",
  4153=>"11111111",
  4154=>"11111011",
  4155=>"00000000",
  4156=>"11111010",
  4157=>"00000000",
  4158=>"00000001",
  4159=>"11111101",
  4160=>"00000100",
  4161=>"11111110",
  4162=>"11111100",
  4163=>"11111110",
  4164=>"00000011",
  4165=>"00000001",
  4166=>"00000011",
  4167=>"11111110",
  4168=>"11111111",
  4169=>"00000000",
  4170=>"11111101",
  4171=>"11111010",
  4172=>"11111110",
  4173=>"11111111",
  4174=>"11111010",
  4175=>"11111011",
  4176=>"00000001",
  4177=>"00000001",
  4178=>"11111111",
  4179=>"00000000",
  4180=>"11111111",
  4181=>"11111100",
  4182=>"00000001",
  4183=>"11111011",
  4184=>"11111101",
  4185=>"00000000",
  4186=>"11111110",
  4187=>"00000001",
  4188=>"00000000",
  4189=>"11111111",
  4190=>"00000001",
  4191=>"00000001",
  4192=>"11111101",
  4193=>"00000001",
  4194=>"00000001",
  4195=>"11111100",
  4196=>"00000000",
  4197=>"11111100",
  4198=>"11111101",
  4199=>"11111101",
  4200=>"00000010",
  4201=>"00000001",
  4202=>"00000000",
  4203=>"00000100",
  4204=>"11111110",
  4205=>"11111111",
  4206=>"11111100",
  4207=>"11111111",
  4208=>"00000010",
  4209=>"00000000",
  4210=>"11111100",
  4211=>"11111110",
  4212=>"11111110",
  4213=>"00000100",
  4214=>"11111111",
  4215=>"11111101",
  4216=>"00000000",
  4217=>"11111011",
  4218=>"00000001",
  4219=>"00000000",
  4220=>"11111101",
  4221=>"00000001",
  4222=>"11111011",
  4223=>"00000010",
  4224=>"11111101",
  4225=>"00000000",
  4226=>"11111110",
  4227=>"00000000",
  4228=>"00000001",
  4229=>"11111110",
  4230=>"11111010",
  4231=>"00000000",
  4232=>"00000110",
  4233=>"00000000",
  4234=>"11111111",
  4235=>"11111110",
  4236=>"00000001",
  4237=>"11111100",
  4238=>"11111111",
  4239=>"11111110",
  4240=>"11111110",
  4241=>"00000001",
  4242=>"00000000",
  4243=>"00000001",
  4244=>"00000010",
  4245=>"11111111",
  4246=>"11111110",
  4247=>"11111101",
  4248=>"11111011",
  4249=>"00000001",
  4250=>"00000011",
  4251=>"00000001",
  4252=>"11111000",
  4253=>"00000010",
  4254=>"11111111",
  4255=>"11111110",
  4256=>"00000001",
  4257=>"00000010",
  4258=>"11111100",
  4259=>"00000001",
  4260=>"11111111",
  4261=>"11111111",
  4262=>"11111011",
  4263=>"11111100",
  4264=>"11111111",
  4265=>"11111100",
  4266=>"11111101",
  4267=>"11111110",
  4268=>"00000010",
  4269=>"00000000",
  4270=>"11111111",
  4271=>"11111011",
  4272=>"11111011",
  4273=>"11111101",
  4274=>"11111100",
  4275=>"00000011",
  4276=>"00000001",
  4277=>"00000000",
  4278=>"11111111",
  4279=>"11111111",
  4280=>"11111101",
  4281=>"11111110",
  4282=>"00000000",
  4283=>"11111110",
  4284=>"11111110",
  4285=>"11111110",
  4286=>"00000000",
  4287=>"00000100",
  4288=>"11111101",
  4289=>"00000001",
  4290=>"11111101",
  4291=>"00000011",
  4292=>"00000001",
  4293=>"11111111",
  4294=>"00000010",
  4295=>"11111100",
  4296=>"00000001",
  4297=>"11111101",
  4298=>"11111110",
  4299=>"11111101",
  4300=>"00000001",
  4301=>"00000010",
  4302=>"11111111",
  4303=>"11111111",
  4304=>"00000000",
  4305=>"00000011",
  4306=>"11111110",
  4307=>"11111100",
  4308=>"11111101",
  4309=>"11111110",
  4310=>"11111100",
  4311=>"00000001",
  4312=>"11111110",
  4313=>"11111111",
  4314=>"11111010",
  4315=>"00000011",
  4316=>"11111010",
  4317=>"11111110",
  4318=>"00000010",
  4319=>"00000000",
  4320=>"11111100",
  4321=>"11111101",
  4322=>"11111110",
  4323=>"11111101",
  4324=>"11111111",
  4325=>"11111110",
  4326=>"11111100",
  4327=>"00000011",
  4328=>"11111110",
  4329=>"11111110",
  4330=>"11111111",
  4331=>"11111001",
  4332=>"11111101",
  4333=>"11111111",
  4334=>"00000110",
  4335=>"11111010",
  4336=>"00000010",
  4337=>"00000001",
  4338=>"11111110",
  4339=>"00000001",
  4340=>"00000001",
  4341=>"00000000",
  4342=>"11111101",
  4343=>"11111110",
  4344=>"11111010",
  4345=>"11111011",
  4346=>"00000000",
  4347=>"11111010",
  4348=>"00000010",
  4349=>"11111101",
  4350=>"11111110",
  4351=>"11111100",
  4352=>"11111111",
  4353=>"00000000",
  4354=>"11111011",
  4355=>"00000100",
  4356=>"11111010",
  4357=>"11111111",
  4358=>"00000000",
  4359=>"00000000",
  4360=>"00000000",
  4361=>"11111101",
  4362=>"00000011",
  4363=>"11111111",
  4364=>"11111101",
  4365=>"00000010",
  4366=>"00000000",
  4367=>"00000000",
  4368=>"00000000",
  4369=>"00000001",
  4370=>"00000011",
  4371=>"11111111",
  4372=>"00000001",
  4373=>"11111101",
  4374=>"00000011",
  4375=>"00000000",
  4376=>"11111111",
  4377=>"11111101",
  4378=>"11111111",
  4379=>"11111100",
  4380=>"00000000",
  4381=>"11111110",
  4382=>"11111101",
  4383=>"00000000",
  4384=>"11111011",
  4385=>"11111111",
  4386=>"00000000",
  4387=>"11111101",
  4388=>"00000001",
  4389=>"11111111",
  4390=>"00000010",
  4391=>"00000000",
  4392=>"11111111",
  4393=>"00000001",
  4394=>"00000001",
  4395=>"11111110",
  4396=>"11111111",
  4397=>"11111100",
  4398=>"11111101",
  4399=>"11111100",
  4400=>"11111110",
  4401=>"11111101",
  4402=>"11111110",
  4403=>"11111100",
  4404=>"11111110",
  4405=>"11111101",
  4406=>"00000010",
  4407=>"11111110",
  4408=>"00000000",
  4409=>"11111101",
  4410=>"11111111",
  4411=>"11111011",
  4412=>"11111100",
  4413=>"00000101",
  4414=>"00000001",
  4415=>"11111011",
  4416=>"11111100",
  4417=>"11111111",
  4418=>"11111101",
  4419=>"00000010",
  4420=>"11111110",
  4421=>"00000000",
  4422=>"00000000",
  4423=>"11111001",
  4424=>"11111100",
  4425=>"00000000",
  4426=>"11111110",
  4427=>"11111111",
  4428=>"00000100",
  4429=>"00000101",
  4430=>"00000011",
  4431=>"00000000",
  4432=>"11111110",
  4433=>"11111111",
  4434=>"00000000",
  4435=>"00000010",
  4436=>"11111111",
  4437=>"11111101",
  4438=>"00000011",
  4439=>"00000001",
  4440=>"11111111",
  4441=>"00000000",
  4442=>"11111100",
  4443=>"00000001",
  4444=>"11111011",
  4445=>"11111111",
  4446=>"11111110",
  4447=>"11111101",
  4448=>"00000001",
  4449=>"11111000",
  4450=>"11111101",
  4451=>"11111101",
  4452=>"11111110",
  4453=>"11111111",
  4454=>"11111101",
  4455=>"11111111",
  4456=>"11111111",
  4457=>"11111111",
  4458=>"11111111",
  4459=>"00000001",
  4460=>"11111011",
  4461=>"11111110",
  4462=>"00000001",
  4463=>"00000000",
  4464=>"11111010",
  4465=>"00000000",
  4466=>"11111101",
  4467=>"11111111",
  4468=>"00000010",
  4469=>"11111110",
  4470=>"11111110",
  4471=>"11111001",
  4472=>"00000001",
  4473=>"11111110",
  4474=>"00000010",
  4475=>"11111101",
  4476=>"11111011",
  4477=>"11111100",
  4478=>"00000010",
  4479=>"00000011",
  4480=>"11111111",
  4481=>"00000001",
  4482=>"11111011",
  4483=>"00000010",
  4484=>"11111101",
  4485=>"00000001",
  4486=>"11111111",
  4487=>"11111111",
  4488=>"11111100",
  4489=>"11111011",
  4490=>"00000000",
  4491=>"11111000",
  4492=>"11111111",
  4493=>"11111111",
  4494=>"00000000",
  4495=>"11111110",
  4496=>"00000000",
  4497=>"00000010",
  4498=>"00000011",
  4499=>"11111110",
  4500=>"11111111",
  4501=>"11111110",
  4502=>"11111111",
  4503=>"00000001",
  4504=>"11111111",
  4505=>"11111101",
  4506=>"11111110",
  4507=>"11111111",
  4508=>"00000001",
  4509=>"11111100",
  4510=>"11111111",
  4511=>"11111110",
  4512=>"11111010",
  4513=>"00000010",
  4514=>"11111111",
  4515=>"00000011",
  4516=>"11111100",
  4517=>"00000010",
  4518=>"11111101",
  4519=>"11111101",
  4520=>"00000010",
  4521=>"00000001",
  4522=>"00000000",
  4523=>"11111100",
  4524=>"11111101",
  4525=>"11111110",
  4526=>"11111101",
  4527=>"11111100",
  4528=>"11111100",
  4529=>"11111111",
  4530=>"11111110",
  4531=>"11111011",
  4532=>"11111111",
  4533=>"11111111",
  4534=>"11111111",
  4535=>"00000000",
  4536=>"00000011",
  4537=>"11111011",
  4538=>"11111111",
  4539=>"00000000",
  4540=>"11111010",
  4541=>"11111111",
  4542=>"00000001",
  4543=>"11111100",
  4544=>"11111111",
  4545=>"00000001",
  4546=>"00000011",
  4547=>"00000010",
  4548=>"00000000",
  4549=>"00000001",
  4550=>"00000000",
  4551=>"00000000",
  4552=>"00000001",
  4553=>"00000000",
  4554=>"00000001",
  4555=>"00000001",
  4556=>"11111101",
  4557=>"11111100",
  4558=>"00000001",
  4559=>"11111100",
  4560=>"00000000",
  4561=>"11111011",
  4562=>"11111100",
  4563=>"11111110",
  4564=>"00000001",
  4565=>"11111111",
  4566=>"11111111",
  4567=>"00000000",
  4568=>"11111011",
  4569=>"00000000",
  4570=>"11111111",
  4571=>"11111101",
  4572=>"00000001",
  4573=>"11111100",
  4574=>"00000010",
  4575=>"00000001",
  4576=>"00000000",
  4577=>"00000000",
  4578=>"11111111",
  4579=>"11111110",
  4580=>"11111100",
  4581=>"00000000",
  4582=>"11111110",
  4583=>"11111001",
  4584=>"11111111",
  4585=>"00000000",
  4586=>"00000010",
  4587=>"00000011",
  4588=>"11111100",
  4589=>"00000010",
  4590=>"00000011",
  4591=>"00000001",
  4592=>"11111001",
  4593=>"11111101",
  4594=>"00000001",
  4595=>"11111111",
  4596=>"11111010",
  4597=>"11111111",
  4598=>"00000001",
  4599=>"11111110",
  4600=>"00000001",
  4601=>"00000000",
  4602=>"11111111",
  4603=>"11111111",
  4604=>"11111111",
  4605=>"11111110",
  4606=>"00000000",
  4607=>"00000101",
  4608=>"11111100",
  4609=>"11111111",
  4610=>"11111111",
  4611=>"00000011",
  4612=>"11111110",
  4613=>"11110111",
  4614=>"00000010",
  4615=>"00000000",
  4616=>"11111111",
  4617=>"00000001",
  4618=>"11111100",
  4619=>"11111101",
  4620=>"00000010",
  4621=>"11111001",
  4622=>"00000010",
  4623=>"00000000",
  4624=>"11111101",
  4625=>"00000011",
  4626=>"00000000",
  4627=>"11111101",
  4628=>"00000001",
  4629=>"11111111",
  4630=>"11111110",
  4631=>"11111110",
  4632=>"11111101",
  4633=>"11111100",
  4634=>"11111111",
  4635=>"00000000",
  4636=>"11111110",
  4637=>"00000001",
  4638=>"00000101",
  4639=>"00000010",
  4640=>"11111111",
  4641=>"00000001",
  4642=>"00000001",
  4643=>"11111110",
  4644=>"00000010",
  4645=>"11111111",
  4646=>"11111110",
  4647=>"00000010",
  4648=>"00000010",
  4649=>"11111111",
  4650=>"00000000",
  4651=>"00000010",
  4652=>"00000001",
  4653=>"11111111",
  4654=>"00000001",
  4655=>"00000001",
  4656=>"11111100",
  4657=>"11111110",
  4658=>"11111010",
  4659=>"11111110",
  4660=>"00000010",
  4661=>"11111111",
  4662=>"00000001",
  4663=>"11111110",
  4664=>"00000001",
  4665=>"00000000",
  4666=>"11111011",
  4667=>"11111101",
  4668=>"00000000",
  4669=>"11111100",
  4670=>"00000001",
  4671=>"00000000",
  4672=>"11111111",
  4673=>"11111111",
  4674=>"00000001",
  4675=>"00000001",
  4676=>"11111011",
  4677=>"11111111",
  4678=>"11111110",
  4679=>"11111110",
  4680=>"11111101",
  4681=>"11111000",
  4682=>"11111100",
  4683=>"00000000",
  4684=>"11111110",
  4685=>"11111111",
  4686=>"00000000",
  4687=>"11111001",
  4688=>"11111111",
  4689=>"00000011",
  4690=>"00000000",
  4691=>"11111110",
  4692=>"00000010",
  4693=>"11111111",
  4694=>"00000000",
  4695=>"11111110",
  4696=>"00000001",
  4697=>"00000001",
  4698=>"11111111",
  4699=>"00000001",
  4700=>"00000001",
  4701=>"11111100",
  4702=>"11111101",
  4703=>"11111101",
  4704=>"11111111",
  4705=>"00000011",
  4706=>"11111011",
  4707=>"11111111",
  4708=>"11111111",
  4709=>"11111100",
  4710=>"11111011",
  4711=>"00000000",
  4712=>"00000000",
  4713=>"00000000",
  4714=>"00000000",
  4715=>"11111011",
  4716=>"00000000",
  4717=>"00000000",
  4718=>"11111100",
  4719=>"11111110",
  4720=>"00000001",
  4721=>"00000010",
  4722=>"11111010",
  4723=>"11111101",
  4724=>"11111100",
  4725=>"00000001",
  4726=>"00000000",
  4727=>"11111111",
  4728=>"11111110",
  4729=>"11111101",
  4730=>"11111111",
  4731=>"11111101",
  4732=>"11111111",
  4733=>"00000010",
  4734=>"11111111",
  4735=>"00000001",
  4736=>"00000001",
  4737=>"00000001",
  4738=>"00000000",
  4739=>"11111110",
  4740=>"11111111",
  4741=>"00000000",
  4742=>"11111101",
  4743=>"00000011",
  4744=>"11111110",
  4745=>"11111010",
  4746=>"00000011",
  4747=>"00000001",
  4748=>"11111111",
  4749=>"11111100",
  4750=>"11111110",
  4751=>"11111011",
  4752=>"00000001",
  4753=>"11111111",
  4754=>"11111110",
  4755=>"11111010",
  4756=>"11111011",
  4757=>"00000001",
  4758=>"11111100",
  4759=>"00000001",
  4760=>"00000000",
  4761=>"00000001",
  4762=>"00000010",
  4763=>"00000000",
  4764=>"00000010",
  4765=>"00000011",
  4766=>"00000000",
  4767=>"11111101",
  4768=>"11111101",
  4769=>"00000001",
  4770=>"00000000",
  4771=>"00000001",
  4772=>"11111110",
  4773=>"00000011",
  4774=>"00000010",
  4775=>"11111100",
  4776=>"00000001",
  4777=>"11111111",
  4778=>"11111101",
  4779=>"11111110",
  4780=>"11111111",
  4781=>"00000010",
  4782=>"11111111",
  4783=>"11111111",
  4784=>"11111011",
  4785=>"00000001",
  4786=>"00000001",
  4787=>"11111110",
  4788=>"11111111",
  4789=>"11111101",
  4790=>"11111011",
  4791=>"00000001",
  4792=>"00000010",
  4793=>"00000100",
  4794=>"11111110",
  4795=>"11111101",
  4796=>"11111111",
  4797=>"11111111",
  4798=>"00000000",
  4799=>"11111111",
  4800=>"00000010",
  4801=>"11111100",
  4802=>"11111101",
  4803=>"00000001",
  4804=>"11111111",
  4805=>"11111001",
  4806=>"11111110",
  4807=>"11111110",
  4808=>"11111101",
  4809=>"00000010",
  4810=>"11111111",
  4811=>"00000001",
  4812=>"11111111",
  4813=>"00000000",
  4814=>"11111011",
  4815=>"00000001",
  4816=>"11111010",
  4817=>"00000010",
  4818=>"11111011",
  4819=>"00000010",
  4820=>"00000001",
  4821=>"11111110",
  4822=>"11111101",
  4823=>"11111111",
  4824=>"11111100",
  4825=>"00000001",
  4826=>"00000001",
  4827=>"00000001",
  4828=>"11111111",
  4829=>"11111110",
  4830=>"00000000",
  4831=>"11111110",
  4832=>"00000011",
  4833=>"00000010",
  4834=>"11111100",
  4835=>"11111011",
  4836=>"00000000",
  4837=>"00000000",
  4838=>"11111101",
  4839=>"11111100",
  4840=>"11111101",
  4841=>"00000000",
  4842=>"11111010",
  4843=>"00000011",
  4844=>"11111011",
  4845=>"11111110",
  4846=>"00000010",
  4847=>"11111111",
  4848=>"00000100",
  4849=>"11111010",
  4850=>"00000000",
  4851=>"11111111",
  4852=>"11111111",
  4853=>"11111110",
  4854=>"11111100",
  4855=>"00000000",
  4856=>"00000010",
  4857=>"11111110",
  4858=>"11111111",
  4859=>"00000000",
  4860=>"11111111",
  4861=>"00000010",
  4862=>"00000011",
  4863=>"00000000",
  4864=>"00000000",
  4865=>"00000100",
  4866=>"11111110",
  4867=>"00000011",
  4868=>"11111111",
  4869=>"11111000",
  4870=>"00000001",
  4871=>"00000110",
  4872=>"00000011",
  4873=>"11111011",
  4874=>"00000011",
  4875=>"11111101",
  4876=>"11111110",
  4877=>"00000001",
  4878=>"00000010",
  4879=>"11111011",
  4880=>"00000000",
  4881=>"11111110",
  4882=>"00000000",
  4883=>"11111011",
  4884=>"11111100",
  4885=>"11111111",
  4886=>"11111110",
  4887=>"11111011",
  4888=>"00000010",
  4889=>"11111111",
  4890=>"11111111",
  4891=>"11111111",
  4892=>"11111011",
  4893=>"11111111",
  4894=>"11111110",
  4895=>"00000000",
  4896=>"11111110",
  4897=>"00000001",
  4898=>"11111111",
  4899=>"00000001",
  4900=>"11111111",
  4901=>"00000000",
  4902=>"00000010",
  4903=>"11111111",
  4904=>"11111110",
  4905=>"00000001",
  4906=>"00000010",
  4907=>"00000010",
  4908=>"11111100",
  4909=>"00000000",
  4910=>"11111111",
  4911=>"11111100",
  4912=>"00000000",
  4913=>"00000001",
  4914=>"11111110",
  4915=>"11111110",
  4916=>"11111010",
  4917=>"00000011",
  4918=>"11111101",
  4919=>"00000000",
  4920=>"11111010",
  4921=>"11111101",
  4922=>"11111110",
  4923=>"11111110",
  4924=>"11111111",
  4925=>"11111101",
  4926=>"00000001",
  4927=>"11111011",
  4928=>"11111111",
  4929=>"11111110",
  4930=>"11111011",
  4931=>"00000001",
  4932=>"00000001",
  4933=>"00000010",
  4934=>"00000000",
  4935=>"00000001",
  4936=>"00000000",
  4937=>"00000001",
  4938=>"11111110",
  4939=>"11111011",
  4940=>"00000000",
  4941=>"11111011",
  4942=>"11111101",
  4943=>"11111011",
  4944=>"11111101",
  4945=>"00000000",
  4946=>"00000000",
  4947=>"00000000",
  4948=>"11111110",
  4949=>"00000000",
  4950=>"11111100",
  4951=>"00000000",
  4952=>"00000011",
  4953=>"00000010",
  4954=>"00000000",
  4955=>"00000001",
  4956=>"11111101",
  4957=>"11111111",
  4958=>"00000001",
  4959=>"00000000",
  4960=>"11111010",
  4961=>"00000000",
  4962=>"11111101",
  4963=>"11111101",
  4964=>"11111111",
  4965=>"00000001",
  4966=>"00000010",
  4967=>"11111110",
  4968=>"00000000",
  4969=>"00000001",
  4970=>"11111111",
  4971=>"00000011",
  4972=>"00000000",
  4973=>"11111110",
  4974=>"11111010",
  4975=>"11111111",
  4976=>"11111011",
  4977=>"11111101",
  4978=>"11111010",
  4979=>"00000000",
  4980=>"11111011",
  4981=>"00000000",
  4982=>"11111111",
  4983=>"11111011",
  4984=>"11111111",
  4985=>"11111100",
  4986=>"11111111",
  4987=>"00000001",
  4988=>"11111111",
  4989=>"11111111",
  4990=>"00000000",
  4991=>"00000001",
  4992=>"11111000",
  4993=>"00000010",
  4994=>"11111110",
  4995=>"00000000",
  4996=>"00000001",
  4997=>"11111100",
  4998=>"00000000",
  4999=>"11111110",
  5000=>"11111111",
  5001=>"11111110",
  5002=>"11111011",
  5003=>"11111011",
  5004=>"00000010",
  5005=>"11111101",
  5006=>"00000001",
  5007=>"11111111",
  5008=>"00000001",
  5009=>"00000010",
  5010=>"11111111",
  5011=>"11111100",
  5012=>"00000000",
  5013=>"00000001",
  5014=>"11111100",
  5015=>"11111110",
  5016=>"00000000",
  5017=>"00000001",
  5018=>"00000000",
  5019=>"00000001",
  5020=>"11111111",
  5021=>"11111011",
  5022=>"11111110",
  5023=>"11111111",
  5024=>"11111111",
  5025=>"11111101",
  5026=>"11111100",
  5027=>"11111010",
  5028=>"11111110",
  5029=>"11111100",
  5030=>"00000000",
  5031=>"00000001",
  5032=>"11111011",
  5033=>"11111110",
  5034=>"11111110",
  5035=>"11111010",
  5036=>"00000001",
  5037=>"11111101",
  5038=>"00000010",
  5039=>"11111111",
  5040=>"11111010",
  5041=>"11111100",
  5042=>"00000000",
  5043=>"11111110",
  5044=>"11111010",
  5045=>"11111011",
  5046=>"00000001",
  5047=>"11111010",
  5048=>"11111110",
  5049=>"11111100",
  5050=>"11111100",
  5051=>"11111111",
  5052=>"00000011",
  5053=>"11111111",
  5054=>"00000000",
  5055=>"11111011",
  5056=>"00000000",
  5057=>"00000010",
  5058=>"11111100",
  5059=>"11111100",
  5060=>"00000010",
  5061=>"11111111",
  5062=>"11111111",
  5063=>"11111010",
  5064=>"11111110",
  5065=>"11111100",
  5066=>"11111111",
  5067=>"00000001",
  5068=>"00000000",
  5069=>"11111110",
  5070=>"00000000",
  5071=>"11111101",
  5072=>"11111110",
  5073=>"00000010",
  5074=>"00000010",
  5075=>"00000011",
  5076=>"00000010",
  5077=>"00000001",
  5078=>"00000001",
  5079=>"00000001",
  5080=>"11111000",
  5081=>"11111110",
  5082=>"11111100",
  5083=>"00000001",
  5084=>"00000001",
  5085=>"00000000",
  5086=>"00000001",
  5087=>"00000011",
  5088=>"00000001",
  5089=>"11111101",
  5090=>"00000001",
  5091=>"11111100",
  5092=>"11111101",
  5093=>"11111011",
  5094=>"00000000",
  5095=>"00000001",
  5096=>"00000010",
  5097=>"11111010",
  5098=>"00000011",
  5099=>"00000010",
  5100=>"11111101",
  5101=>"11111110",
  5102=>"11111110",
  5103=>"00000010",
  5104=>"00000001",
  5105=>"11111011",
  5106=>"11111111",
  5107=>"00000001",
  5108=>"00000001",
  5109=>"11111111",
  5110=>"00000000",
  5111=>"00000000",
  5112=>"00000001",
  5113=>"00000000",
  5114=>"00000000",
  5115=>"00000010",
  5116=>"11111101",
  5117=>"11111111",
  5118=>"00000000",
  5119=>"11111111",
  5120=>"00000010",
  5121=>"11111101",
  5122=>"00000000",
  5123=>"11111110",
  5124=>"11111110",
  5125=>"00000011",
  5126=>"00000011",
  5127=>"11111100",
  5128=>"11111101",
  5129=>"11111111",
  5130=>"00000100",
  5131=>"11111111",
  5132=>"00000110",
  5133=>"11111110",
  5134=>"11111101",
  5135=>"00000010",
  5136=>"11111111",
  5137=>"00000001",
  5138=>"00000001",
  5139=>"11111110",
  5140=>"11111100",
  5141=>"00000101",
  5142=>"11111101",
  5143=>"00000001",
  5144=>"11111111",
  5145=>"00000011",
  5146=>"11111110",
  5147=>"00000000",
  5148=>"00000000",
  5149=>"00000000",
  5150=>"11111110",
  5151=>"11111110",
  5152=>"00000011",
  5153=>"11111111",
  5154=>"11111111",
  5155=>"11111111",
  5156=>"00000001",
  5157=>"00000000",
  5158=>"11111111",
  5159=>"00000000",
  5160=>"11111100",
  5161=>"11111111",
  5162=>"00000010",
  5163=>"00000010",
  5164=>"00000000",
  5165=>"00000010",
  5166=>"00000011",
  5167=>"00000110",
  5168=>"00000000",
  5169=>"00000000",
  5170=>"11111110",
  5171=>"11111111",
  5172=>"11111111",
  5173=>"11111111",
  5174=>"11111101",
  5175=>"00000100",
  5176=>"11111101",
  5177=>"00000000",
  5178=>"00000000",
  5179=>"00000011",
  5180=>"11111111",
  5181=>"00000011",
  5182=>"00000001",
  5183=>"11111101",
  5184=>"11111111",
  5185=>"11111110",
  5186=>"00000000",
  5187=>"00000100",
  5188=>"00000001",
  5189=>"11111100",
  5190=>"00000000",
  5191=>"00000000",
  5192=>"00000000",
  5193=>"11111110",
  5194=>"00000001",
  5195=>"11111110",
  5196=>"11111101",
  5197=>"00000001",
  5198=>"11111110",
  5199=>"00000000",
  5200=>"11111100",
  5201=>"11111110",
  5202=>"11111100",
  5203=>"00000000",
  5204=>"11111111",
  5205=>"11111110",
  5206=>"00000001",
  5207=>"00000010",
  5208=>"00000100",
  5209=>"11111101",
  5210=>"11111111",
  5211=>"00000011",
  5212=>"00000101",
  5213=>"11111110",
  5214=>"11111101",
  5215=>"00000000",
  5216=>"00000000",
  5217=>"00000001",
  5218=>"11111101",
  5219=>"00000001",
  5220=>"00000101",
  5221=>"00000010",
  5222=>"11111110",
  5223=>"11111110",
  5224=>"11111101",
  5225=>"00000100",
  5226=>"11111110",
  5227=>"11111100",
  5228=>"00000001",
  5229=>"11111101",
  5230=>"00000000",
  5231=>"00000011",
  5232=>"00000000",
  5233=>"00000001",
  5234=>"00000000",
  5235=>"11111101",
  5236=>"00000010",
  5237=>"11111110",
  5238=>"00000001",
  5239=>"00000010",
  5240=>"00000000",
  5241=>"11111101",
  5242=>"11111111",
  5243=>"00000001",
  5244=>"11111111",
  5245=>"00000001",
  5246=>"00000011",
  5247=>"00000001",
  5248=>"11111111",
  5249=>"11111100",
  5250=>"11111101",
  5251=>"11111101",
  5252=>"00000100",
  5253=>"11111110",
  5254=>"11111110",
  5255=>"11111100",
  5256=>"11111110",
  5257=>"00000000",
  5258=>"11111110",
  5259=>"00000010",
  5260=>"00000000",
  5261=>"00000010",
  5262=>"00000001",
  5263=>"11111101",
  5264=>"00000001",
  5265=>"00000001",
  5266=>"11111101",
  5267=>"11111111",
  5268=>"00000010",
  5269=>"00000010",
  5270=>"11111110",
  5271=>"11111111",
  5272=>"00000001",
  5273=>"00000011",
  5274=>"11111101",
  5275=>"11111101",
  5276=>"00000000",
  5277=>"00000010",
  5278=>"00000100",
  5279=>"00000001",
  5280=>"11111110",
  5281=>"11111100",
  5282=>"00000010",
  5283=>"11111101",
  5284=>"11111110",
  5285=>"00000011",
  5286=>"11111110",
  5287=>"00000000",
  5288=>"11111111",
  5289=>"11111110",
  5290=>"00000000",
  5291=>"11111101",
  5292=>"11111101",
  5293=>"11111110",
  5294=>"11111100",
  5295=>"11111110",
  5296=>"00000010",
  5297=>"11111110",
  5298=>"00000000",
  5299=>"00000101",
  5300=>"11111110",
  5301=>"00000001",
  5302=>"00000000",
  5303=>"11111100",
  5304=>"00000001",
  5305=>"11111111",
  5306=>"11111111",
  5307=>"11111101",
  5308=>"00000001",
  5309=>"11111110",
  5310=>"00000011",
  5311=>"00000001",
  5312=>"11111111",
  5313=>"00000010",
  5314=>"00000011",
  5315=>"00000000",
  5316=>"00000001",
  5317=>"11111100",
  5318=>"00000001",
  5319=>"11111101",
  5320=>"11111111",
  5321=>"00000001",
  5322=>"11111101",
  5323=>"00000010",
  5324=>"11111110",
  5325=>"11111111",
  5326=>"11111110",
  5327=>"11111110",
  5328=>"00000000",
  5329=>"00000000",
  5330=>"11111110",
  5331=>"00000100",
  5332=>"00000001",
  5333=>"11111111",
  5334=>"11111110",
  5335=>"11111110",
  5336=>"11111111",
  5337=>"11111110",
  5338=>"00000000",
  5339=>"00000001",
  5340=>"00000010",
  5341=>"11111111",
  5342=>"11111111",
  5343=>"11111101",
  5344=>"00000010",
  5345=>"11111110",
  5346=>"00000100",
  5347=>"00000000",
  5348=>"11111101",
  5349=>"11111101",
  5350=>"00000000",
  5351=>"00000000",
  5352=>"00000010",
  5353=>"00000001",
  5354=>"00000010",
  5355=>"11111110",
  5356=>"00000011",
  5357=>"00000000",
  5358=>"11111111",
  5359=>"00000001",
  5360=>"11111101",
  5361=>"00000010",
  5362=>"00000000",
  5363=>"00000110",
  5364=>"11111110",
  5365=>"00000010",
  5366=>"11111110",
  5367=>"00000001",
  5368=>"00000000",
  5369=>"11111111",
  5370=>"11111110",
  5371=>"00000011",
  5372=>"00000010",
  5373=>"00000010",
  5374=>"11111101",
  5375=>"00000001",
  5376=>"00000100",
  5377=>"00000000",
  5378=>"11111101",
  5379=>"00000001",
  5380=>"00000011",
  5381=>"00000001",
  5382=>"11111111",
  5383=>"00000110",
  5384=>"11111111",
  5385=>"11111110",
  5386=>"11111100",
  5387=>"11111111",
  5388=>"00000011",
  5389=>"11111111",
  5390=>"11111100",
  5391=>"11111100",
  5392=>"11111101",
  5393=>"00000000",
  5394=>"11111101",
  5395=>"00000000",
  5396=>"11111111",
  5397=>"11111111",
  5398=>"11111101",
  5399=>"00000010",
  5400=>"00000101",
  5401=>"11111111",
  5402=>"00000001",
  5403=>"00000000",
  5404=>"11111101",
  5405=>"00000111",
  5406=>"11111110",
  5407=>"00000101",
  5408=>"00000000",
  5409=>"11111110",
  5410=>"00000100",
  5411=>"00000000",
  5412=>"11111101",
  5413=>"11111110",
  5414=>"11111111",
  5415=>"11111111",
  5416=>"11111111",
  5417=>"11111110",
  5418=>"00001000",
  5419=>"11111110",
  5420=>"00000011",
  5421=>"11111101",
  5422=>"00000000",
  5423=>"11111101",
  5424=>"00000101",
  5425=>"00000001",
  5426=>"00000001",
  5427=>"11111110",
  5428=>"00000001",
  5429=>"00000001",
  5430=>"00000110",
  5431=>"11111111",
  5432=>"11111101",
  5433=>"00000001",
  5434=>"11111100",
  5435=>"11111111",
  5436=>"11111111",
  5437=>"11111101",
  5438=>"00000011",
  5439=>"11111101",
  5440=>"00000000",
  5441=>"00000001",
  5442=>"00000001",
  5443=>"00000000",
  5444=>"11111110",
  5445=>"00000010",
  5446=>"11111100",
  5447=>"00000000",
  5448=>"11111110",
  5449=>"00000101",
  5450=>"00000001",
  5451=>"11111111",
  5452=>"00000010",
  5453=>"00000010",
  5454=>"11111110",
  5455=>"00000001",
  5456=>"00000001",
  5457=>"00000100",
  5458=>"00000010",
  5459=>"00000001",
  5460=>"00000010",
  5461=>"00000010",
  5462=>"11111110",
  5463=>"00000010",
  5464=>"00000010",
  5465=>"11111101",
  5466=>"11111101",
  5467=>"00000010",
  5468=>"11111111",
  5469=>"00000010",
  5470=>"00000010",
  5471=>"00000010",
  5472=>"00000010",
  5473=>"00000000",
  5474=>"00000010",
  5475=>"00000010",
  5476=>"11111111",
  5477=>"00000001",
  5478=>"11111110",
  5479=>"00000011",
  5480=>"11111111",
  5481=>"11111110",
  5482=>"11111101",
  5483=>"00000000",
  5484=>"00000000",
  5485=>"11111111",
  5486=>"11111110",
  5487=>"11111111",
  5488=>"11111111",
  5489=>"11111110",
  5490=>"11111101",
  5491=>"11111101",
  5492=>"11111101",
  5493=>"11111110",
  5494=>"11111101",
  5495=>"00000001",
  5496=>"11111110",
  5497=>"11111100",
  5498=>"11111111",
  5499=>"00000000",
  5500=>"11111101",
  5501=>"00000000",
  5502=>"00000110",
  5503=>"00000001",
  5504=>"11111101",
  5505=>"11111110",
  5506=>"00000000",
  5507=>"00000010",
  5508=>"00000010",
  5509=>"00000000",
  5510=>"11111101",
  5511=>"11111111",
  5512=>"00000001",
  5513=>"11111111",
  5514=>"00000101",
  5515=>"11111110",
  5516=>"00000010",
  5517=>"11111110",
  5518=>"00000001",
  5519=>"11111101",
  5520=>"00000000",
  5521=>"00000010",
  5522=>"11111111",
  5523=>"00000001",
  5524=>"11111100",
  5525=>"11111111",
  5526=>"11111111",
  5527=>"11111111",
  5528=>"11111111",
  5529=>"00000010",
  5530=>"11111110",
  5531=>"00000011",
  5532=>"11111111",
  5533=>"11111110",
  5534=>"11111111",
  5535=>"00000000",
  5536=>"11111110",
  5537=>"00000001",
  5538=>"11111101",
  5539=>"11111101",
  5540=>"11111110",
  5541=>"11111101",
  5542=>"00000000",
  5543=>"11111110",
  5544=>"00000100",
  5545=>"00000010",
  5546=>"00000000",
  5547=>"00000000",
  5548=>"00000010",
  5549=>"11111101",
  5550=>"00000010",
  5551=>"11111101",
  5552=>"00000100",
  5553=>"11111110",
  5554=>"00000001",
  5555=>"00000010",
  5556=>"00000001",
  5557=>"00000011",
  5558=>"11111111",
  5559=>"11111101",
  5560=>"00000010",
  5561=>"00000001",
  5562=>"00000001",
  5563=>"11111100",
  5564=>"00000010",
  5565=>"11111101",
  5566=>"11111111",
  5567=>"00000100",
  5568=>"00000011",
  5569=>"00000011",
  5570=>"11111100",
  5571=>"11111110",
  5572=>"11111100",
  5573=>"00000000",
  5574=>"11111110",
  5575=>"00000001",
  5576=>"11111101",
  5577=>"00000000",
  5578=>"00000000",
  5579=>"00000011",
  5580=>"00000000",
  5581=>"00000000",
  5582=>"11111110",
  5583=>"00000000",
  5584=>"00000011",
  5585=>"00000000",
  5586=>"00000001",
  5587=>"00000000",
  5588=>"00000000",
  5589=>"00000001",
  5590=>"00000110",
  5591=>"11111101",
  5592=>"00000000",
  5593=>"00000011",
  5594=>"11111101",
  5595=>"11111101",
  5596=>"00000011",
  5597=>"00000001",
  5598=>"11111110",
  5599=>"11111111",
  5600=>"11111110",
  5601=>"11111110",
  5602=>"00000001",
  5603=>"00000000",
  5604=>"00000010",
  5605=>"00000010",
  5606=>"11111110",
  5607=>"00000010",
  5608=>"11111100",
  5609=>"00000010",
  5610=>"00000101",
  5611=>"00000010",
  5612=>"00000000",
  5613=>"00000011",
  5614=>"00000011",
  5615=>"11111110",
  5616=>"00000001",
  5617=>"00000010",
  5618=>"00000011",
  5619=>"11111100",
  5620=>"00000010",
  5621=>"00000010",
  5622=>"11111110",
  5623=>"00000000",
  5624=>"00000001",
  5625=>"11111110",
  5626=>"00000000",
  5627=>"11111111",
  5628=>"11111101",
  5629=>"00000000",
  5630=>"00000010",
  5631=>"00000000",
  5632=>"00000010",
  5633=>"11111111",
  5634=>"00000010",
  5635=>"00000001",
  5636=>"11111111",
  5637=>"11111110",
  5638=>"00000001",
  5639=>"11111111",
  5640=>"00000100",
  5641=>"00000000",
  5642=>"11111111",
  5643=>"11111111",
  5644=>"11111110",
  5645=>"00000001",
  5646=>"00000010",
  5647=>"00000011",
  5648=>"00000000",
  5649=>"00000101",
  5650=>"00000100",
  5651=>"11111110",
  5652=>"11111111",
  5653=>"11111101",
  5654=>"00000001",
  5655=>"11111110",
  5656=>"11111111",
  5657=>"11111110",
  5658=>"11111110",
  5659=>"00000000",
  5660=>"00000100",
  5661=>"11111101",
  5662=>"00000011",
  5663=>"00000001",
  5664=>"00000000",
  5665=>"00000010",
  5666=>"11111110",
  5667=>"00000001",
  5668=>"11111111",
  5669=>"11111100",
  5670=>"00000110",
  5671=>"11111111",
  5672=>"00000000",
  5673=>"11111101",
  5674=>"00000001",
  5675=>"00000100",
  5676=>"00000010",
  5677=>"11111111",
  5678=>"00000101",
  5679=>"11111110",
  5680=>"11111110",
  5681=>"00000100",
  5682=>"00000001",
  5683=>"00000010",
  5684=>"00000011",
  5685=>"11111110",
  5686=>"00000010",
  5687=>"11111110",
  5688=>"00000010",
  5689=>"11111111",
  5690=>"00000010",
  5691=>"11111111",
  5692=>"11111110",
  5693=>"11111111",
  5694=>"11111011",
  5695=>"00000010",
  5696=>"00000100",
  5697=>"11111110",
  5698=>"00000010",
  5699=>"11111111",
  5700=>"11111111",
  5701=>"00000000",
  5702=>"00000010",
  5703=>"00000100",
  5704=>"00000100",
  5705=>"00000001",
  5706=>"00000010",
  5707=>"11111111",
  5708=>"11111110",
  5709=>"00000011",
  5710=>"11111101",
  5711=>"00000000",
  5712=>"00000000",
  5713=>"00000001",
  5714=>"00000000",
  5715=>"00000001",
  5716=>"11111101",
  5717=>"11111110",
  5718=>"00000001",
  5719=>"00000010",
  5720=>"00000010",
  5721=>"00000000",
  5722=>"11111101",
  5723=>"11111110",
  5724=>"00000011",
  5725=>"11111101",
  5726=>"11111101",
  5727=>"00000010",
  5728=>"00000000",
  5729=>"00000010",
  5730=>"11111110",
  5731=>"00000101",
  5732=>"11111111",
  5733=>"11111111",
  5734=>"00000010",
  5735=>"11111110",
  5736=>"11111100",
  5737=>"00000011",
  5738=>"00000001",
  5739=>"11111111",
  5740=>"00000000",
  5741=>"00000001",
  5742=>"11111101",
  5743=>"11111110",
  5744=>"00000000",
  5745=>"00000000",
  5746=>"00000010",
  5747=>"00000001",
  5748=>"00000011",
  5749=>"00000001",
  5750=>"00000000",
  5751=>"11111111",
  5752=>"00000101",
  5753=>"00000011",
  5754=>"00000011",
  5755=>"00000011",
  5756=>"11111101",
  5757=>"00000001",
  5758=>"00000000",
  5759=>"00000011",
  5760=>"00000010",
  5761=>"11111101",
  5762=>"00000000",
  5763=>"00000001",
  5764=>"11111110",
  5765=>"00000000",
  5766=>"00000101",
  5767=>"11111110",
  5768=>"11111101",
  5769=>"00000010",
  5770=>"00000001",
  5771=>"00000100",
  5772=>"00000000",
  5773=>"00000001",
  5774=>"11111110",
  5775=>"11111111",
  5776=>"11111101",
  5777=>"11111100",
  5778=>"11111101",
  5779=>"11111110",
  5780=>"00000000",
  5781=>"00000010",
  5782=>"00000010",
  5783=>"00000010",
  5784=>"00000010",
  5785=>"11111110",
  5786=>"11111111",
  5787=>"00000010",
  5788=>"11111101",
  5789=>"11111101",
  5790=>"11111111",
  5791=>"00000000",
  5792=>"11111110",
  5793=>"00000011",
  5794=>"11111110",
  5795=>"00000001",
  5796=>"11111110",
  5797=>"11111111",
  5798=>"00000001",
  5799=>"11111111",
  5800=>"11111100",
  5801=>"00000001",
  5802=>"11111110",
  5803=>"00000000",
  5804=>"11111110",
  5805=>"00000000",
  5806=>"00000001",
  5807=>"00000001",
  5808=>"00000001",
  5809=>"11111101",
  5810=>"00000010",
  5811=>"11111100",
  5812=>"00000011",
  5813=>"00000010",
  5814=>"00000100",
  5815=>"00000001",
  5816=>"00000000",
  5817=>"11111101",
  5818=>"11111111",
  5819=>"00000010",
  5820=>"11111110",
  5821=>"00000001",
  5822=>"11111111",
  5823=>"00000000",
  5824=>"00000000",
  5825=>"00000001",
  5826=>"00000010",
  5827=>"00000010",
  5828=>"11111110",
  5829=>"00000001",
  5830=>"11111101",
  5831=>"11111101",
  5832=>"11111111",
  5833=>"11111110",
  5834=>"00000010",
  5835=>"11111111",
  5836=>"00000011",
  5837=>"00000000",
  5838=>"11111110",
  5839=>"11111110",
  5840=>"00000010",
  5841=>"00000011",
  5842=>"00000000",
  5843=>"00000001",
  5844=>"11111110",
  5845=>"11111111",
  5846=>"11111111",
  5847=>"11111110",
  5848=>"11111111",
  5849=>"00000100",
  5850=>"00000100",
  5851=>"00000010",
  5852=>"00000001",
  5853=>"11111110",
  5854=>"00000011",
  5855=>"11111111",
  5856=>"11111101",
  5857=>"00000010",
  5858=>"11111110",
  5859=>"11111110",
  5860=>"11111111",
  5861=>"11111101",
  5862=>"00000000",
  5863=>"00000000",
  5864=>"00000001",
  5865=>"11111111",
  5866=>"11111111",
  5867=>"11111111",
  5868=>"11111101",
  5869=>"00000010",
  5870=>"11111110",
  5871=>"00000011",
  5872=>"00000010",
  5873=>"00000010",
  5874=>"00000010",
  5875=>"00000011",
  5876=>"00000011",
  5877=>"11111111",
  5878=>"00000001",
  5879=>"11111111",
  5880=>"11111110",
  5881=>"00000001",
  5882=>"00000100",
  5883=>"00000001",
  5884=>"00000010",
  5885=>"00000011",
  5886=>"11111101",
  5887=>"11111110",
  5888=>"00000110",
  5889=>"11111111",
  5890=>"11111101",
  5891=>"11111101",
  5892=>"00000000",
  5893=>"00000010",
  5894=>"00000010",
  5895=>"11111101",
  5896=>"11111101",
  5897=>"11111101",
  5898=>"00000010",
  5899=>"11111110",
  5900=>"00000001",
  5901=>"00000010",
  5902=>"11111100",
  5903=>"11111101",
  5904=>"11111110",
  5905=>"00000100",
  5906=>"00000001",
  5907=>"11111110",
  5908=>"11111101",
  5909=>"00000000",
  5910=>"00000000",
  5911=>"11111110",
  5912=>"11111101",
  5913=>"00000000",
  5914=>"11111111",
  5915=>"11111110",
  5916=>"11111111",
  5917=>"00000000",
  5918=>"11111101",
  5919=>"11111100",
  5920=>"00000010",
  5921=>"00000001",
  5922=>"11111101",
  5923=>"11111110",
  5924=>"11111101",
  5925=>"11111100",
  5926=>"00000001",
  5927=>"11111101",
  5928=>"11111101",
  5929=>"11111100",
  5930=>"00000000",
  5931=>"00000011",
  5932=>"00000011",
  5933=>"00000000",
  5934=>"00000011",
  5935=>"11111110",
  5936=>"00000001",
  5937=>"11111111",
  5938=>"11111110",
  5939=>"00000001",
  5940=>"11111101",
  5941=>"00000000",
  5942=>"11111110",
  5943=>"11111110",
  5944=>"00000000",
  5945=>"00000001",
  5946=>"11111110",
  5947=>"00000001",
  5948=>"11111101",
  5949=>"11111111",
  5950=>"00000001",
  5951=>"11111101",
  5952=>"00000011",
  5953=>"00000001",
  5954=>"00000000",
  5955=>"00000011",
  5956=>"00000001",
  5957=>"11111101",
  5958=>"11111110",
  5959=>"11111101",
  5960=>"11111110",
  5961=>"00000010",
  5962=>"00000101",
  5963=>"11111110",
  5964=>"11111111",
  5965=>"00000001",
  5966=>"11111110",
  5967=>"00000011",
  5968=>"11111111",
  5969=>"00000000",
  5970=>"00000001",
  5971=>"11111101",
  5972=>"11111111",
  5973=>"00000011",
  5974=>"11111111",
  5975=>"11111101",
  5976=>"00000000",
  5977=>"00000010",
  5978=>"00000011",
  5979=>"11111110",
  5980=>"00000011",
  5981=>"11111111",
  5982=>"11111101",
  5983=>"00000010",
  5984=>"00000000",
  5985=>"00000011",
  5986=>"00000001",
  5987=>"11111110",
  5988=>"00000100",
  5989=>"00000001",
  5990=>"00000011",
  5991=>"11111100",
  5992=>"00000001",
  5993=>"00000010",
  5994=>"11111101",
  5995=>"11111101",
  5996=>"11111101",
  5997=>"11111101",
  5998=>"11111110",
  5999=>"11111111",
  6000=>"00000010",
  6001=>"00000000",
  6002=>"00000001",
  6003=>"11111110",
  6004=>"11111111",
  6005=>"11111101",
  6006=>"00000001",
  6007=>"00000010",
  6008=>"00000001",
  6009=>"11111101",
  6010=>"11111100",
  6011=>"11111111",
  6012=>"00000011",
  6013=>"11111101",
  6014=>"11111110",
  6015=>"11111101",
  6016=>"00000000",
  6017=>"11111100",
  6018=>"00000010",
  6019=>"11111101",
  6020=>"00000110",
  6021=>"00000000",
  6022=>"11111111",
  6023=>"00000000",
  6024=>"00000010",
  6025=>"00000000",
  6026=>"00000010",
  6027=>"11111110",
  6028=>"00000111",
  6029=>"00000000",
  6030=>"00000010",
  6031=>"00000000",
  6032=>"11111110",
  6033=>"11111100",
  6034=>"00000011",
  6035=>"00000010",
  6036=>"11111101",
  6037=>"11111101",
  6038=>"11111111",
  6039=>"00000000",
  6040=>"00000000",
  6041=>"00000010",
  6042=>"11111110",
  6043=>"11111110",
  6044=>"11111100",
  6045=>"00000000",
  6046=>"00000001",
  6047=>"11111111",
  6048=>"00000000",
  6049=>"11111110",
  6050=>"00000011",
  6051=>"00000001",
  6052=>"00000001",
  6053=>"11111110",
  6054=>"11111110",
  6055=>"00000001",
  6056=>"00000001",
  6057=>"00000100",
  6058=>"00000001",
  6059=>"11111111",
  6060=>"00000000",
  6061=>"11111110",
  6062=>"00000001",
  6063=>"00000011",
  6064=>"11111111",
  6065=>"11111111",
  6066=>"00000001",
  6067=>"11111111",
  6068=>"00000011",
  6069=>"11111110",
  6070=>"11111101",
  6071=>"00000000",
  6072=>"00000000",
  6073=>"00000000",
  6074=>"00000001",
  6075=>"00000011",
  6076=>"11111111",
  6077=>"00000010",
  6078=>"00000000",
  6079=>"00000001",
  6080=>"00000010",
  6081=>"11111101",
  6082=>"11111110",
  6083=>"11111110",
  6084=>"11111101",
  6085=>"00000001",
  6086=>"00000001",
  6087=>"00000010",
  6088=>"11111111",
  6089=>"11111111",
  6090=>"00000110",
  6091=>"11111101",
  6092=>"00000001",
  6093=>"00000010",
  6094=>"11111101",
  6095=>"00000100",
  6096=>"11111111",
  6097=>"00000101",
  6098=>"00000000",
  6099=>"11111101",
  6100=>"11111101",
  6101=>"11111111",
  6102=>"00000000",
  6103=>"11111110",
  6104=>"00000010",
  6105=>"11111111",
  6106=>"11111100",
  6107=>"00000011",
  6108=>"11111111",
  6109=>"11111111",
  6110=>"00000000",
  6111=>"11111100",
  6112=>"11111111",
  6113=>"00000100",
  6114=>"11111110",
  6115=>"00000001",
  6116=>"00000000",
  6117=>"11111101",
  6118=>"00000011",
  6119=>"00000011",
  6120=>"00000100",
  6121=>"00000001",
  6122=>"11111100",
  6123=>"11111111",
  6124=>"11111111",
  6125=>"11111101",
  6126=>"00000001",
  6127=>"00000000",
  6128=>"00000001",
  6129=>"00000001",
  6130=>"00000011",
  6131=>"11111100",
  6132=>"11111110",
  6133=>"00000000",
  6134=>"11111110",
  6135=>"11111100",
  6136=>"00000011",
  6137=>"11111101",
  6138=>"00000010",
  6139=>"11111101",
  6140=>"00000001",
  6141=>"11111110",
  6142=>"11111110",
  6143=>"11111101",
  6144=>"11111111",
  6145=>"00000000",
  6146=>"11111101",
  6147=>"00000010",
  6148=>"00000010",
  6149=>"00000010",
  6150=>"00000000",
  6151=>"11111110",
  6152=>"11111110",
  6153=>"00000000",
  6154=>"00000011",
  6155=>"00000011",
  6156=>"00000010",
  6157=>"11111110",
  6158=>"11111110",
  6159=>"00000000",
  6160=>"11111101",
  6161=>"11111110",
  6162=>"00000010",
  6163=>"11111111",
  6164=>"00000001",
  6165=>"00000011",
  6166=>"11111110",
  6167=>"11111111",
  6168=>"11111101",
  6169=>"11111110",
  6170=>"00000000",
  6171=>"00000011",
  6172=>"00000000",
  6173=>"00000011",
  6174=>"00000011",
  6175=>"00000100",
  6176=>"00000010",
  6177=>"00000011",
  6178=>"00000000",
  6179=>"11111110",
  6180=>"00000010",
  6181=>"11111101",
  6182=>"00000010",
  6183=>"11111110",
  6184=>"00000010",
  6185=>"00000001",
  6186=>"00000010",
  6187=>"11111110",
  6188=>"11111101",
  6189=>"11111100",
  6190=>"00000011",
  6191=>"11111101",
  6192=>"11111110",
  6193=>"00000001",
  6194=>"11111111",
  6195=>"00000011",
  6196=>"00000010",
  6197=>"00000001",
  6198=>"11111110",
  6199=>"00000101",
  6200=>"00000000",
  6201=>"00000011",
  6202=>"00000010",
  6203=>"11111110",
  6204=>"00000001",
  6205=>"00000001",
  6206=>"11111100",
  6207=>"00000000",
  6208=>"00000000",
  6209=>"00000000",
  6210=>"00000001",
  6211=>"11111110",
  6212=>"00000010",
  6213=>"00000000",
  6214=>"11111111",
  6215=>"11111110",
  6216=>"11111110",
  6217=>"00000110",
  6218=>"11111111",
  6219=>"11111111",
  6220=>"11111110",
  6221=>"11111111",
  6222=>"11111110",
  6223=>"11111111",
  6224=>"11111110",
  6225=>"00000000",
  6226=>"11111101",
  6227=>"11111100",
  6228=>"11111101",
  6229=>"11111110",
  6230=>"00000010",
  6231=>"00000010",
  6232=>"11111110",
  6233=>"11111111",
  6234=>"11111110",
  6235=>"00000010",
  6236=>"11111110",
  6237=>"11111101",
  6238=>"11111110",
  6239=>"00000000",
  6240=>"00000001",
  6241=>"00000010",
  6242=>"00000010",
  6243=>"11111110",
  6244=>"11111111",
  6245=>"11111110",
  6246=>"11111111",
  6247=>"11111111",
  6248=>"11111101",
  6249=>"00000110",
  6250=>"00000000",
  6251=>"11111111",
  6252=>"11111111",
  6253=>"00000111",
  6254=>"11111111",
  6255=>"00000010",
  6256=>"11111111",
  6257=>"00000000",
  6258=>"00000010",
  6259=>"00000010",
  6260=>"00000010",
  6261=>"00000000",
  6262=>"00000000",
  6263=>"00000011",
  6264=>"11111111",
  6265=>"00000010",
  6266=>"00000100",
  6267=>"00000000",
  6268=>"11111101",
  6269=>"00000010",
  6270=>"11111101",
  6271=>"00000000",
  6272=>"00000000",
  6273=>"00000111",
  6274=>"00000100",
  6275=>"00000011",
  6276=>"11111101",
  6277=>"11111110",
  6278=>"00000000",
  6279=>"11111110",
  6280=>"11111101",
  6281=>"11111101",
  6282=>"11111111",
  6283=>"00000000",
  6284=>"11111101",
  6285=>"00000010",
  6286=>"11111110",
  6287=>"00000000",
  6288=>"11111101",
  6289=>"00000011",
  6290=>"11111110",
  6291=>"00000100",
  6292=>"11111111",
  6293=>"11111110",
  6294=>"00000001",
  6295=>"00000011",
  6296=>"00000100",
  6297=>"11111111",
  6298=>"11111111",
  6299=>"11111100",
  6300=>"11111110",
  6301=>"11111111",
  6302=>"00000001",
  6303=>"00000001",
  6304=>"11111111",
  6305=>"00000011",
  6306=>"00000001",
  6307=>"00000001",
  6308=>"00000011",
  6309=>"11111110",
  6310=>"00000010",
  6311=>"00000011",
  6312=>"11111111",
  6313=>"11111110",
  6314=>"11111110",
  6315=>"00000000",
  6316=>"00000101",
  6317=>"00000010",
  6318=>"00000011",
  6319=>"11111110",
  6320=>"00000001",
  6321=>"11111111",
  6322=>"11111110",
  6323=>"11111111",
  6324=>"11111111",
  6325=>"00000011",
  6326=>"11111110",
  6327=>"11111111",
  6328=>"11111110",
  6329=>"00000001",
  6330=>"00000000",
  6331=>"11111110",
  6332=>"11111110",
  6333=>"11111110",
  6334=>"11111100",
  6335=>"00000000",
  6336=>"00000001",
  6337=>"00000001",
  6338=>"11111110",
  6339=>"11111111",
  6340=>"00000010",
  6341=>"11111101",
  6342=>"00000010",
  6343=>"11111101",
  6344=>"00000000",
  6345=>"11111101",
  6346=>"00000001",
  6347=>"11111101",
  6348=>"00000010",
  6349=>"11111111",
  6350=>"11111110",
  6351=>"00000001",
  6352=>"00000010",
  6353=>"11111110",
  6354=>"00000010",
  6355=>"00000010",
  6356=>"11111111",
  6357=>"11111110",
  6358=>"11111111",
  6359=>"11111111",
  6360=>"00000010",
  6361=>"00000001",
  6362=>"00000010",
  6363=>"11111111",
  6364=>"00000011",
  6365=>"00000001",
  6366=>"00000010",
  6367=>"00000001",
  6368=>"00000001",
  6369=>"11111111",
  6370=>"11111110",
  6371=>"11111111",
  6372=>"11111101",
  6373=>"00000001",
  6374=>"11111111",
  6375=>"11111111",
  6376=>"00000011",
  6377=>"00000010",
  6378=>"00000001",
  6379=>"00000001",
  6380=>"11111101",
  6381=>"11111100",
  6382=>"11111111",
  6383=>"00000000",
  6384=>"00000000",
  6385=>"11111101",
  6386=>"00000001",
  6387=>"00000101",
  6388=>"11111111",
  6389=>"00000011",
  6390=>"11111111",
  6391=>"11111110",
  6392=>"00000001",
  6393=>"11111110",
  6394=>"00000000",
  6395=>"00000000",
  6396=>"00000010",
  6397=>"11111111",
  6398=>"11111110",
  6399=>"00000000",
  6400=>"00000001",
  6401=>"11111110",
  6402=>"00000011",
  6403=>"00000101",
  6404=>"11111101",
  6405=>"11111110",
  6406=>"11111111",
  6407=>"11111100",
  6408=>"00000100",
  6409=>"11111110",
  6410=>"00000010",
  6411=>"11111100",
  6412=>"11111110",
  6413=>"00000101",
  6414=>"00000001",
  6415=>"00000010",
  6416=>"11111100",
  6417=>"11111100",
  6418=>"11111111",
  6419=>"11111110",
  6420=>"00000001",
  6421=>"00000010",
  6422=>"00000000",
  6423=>"11111111",
  6424=>"11111101",
  6425=>"11111101",
  6426=>"00000010",
  6427=>"11111100",
  6428=>"00000000",
  6429=>"11111101",
  6430=>"00000000",
  6431=>"11111111",
  6432=>"00000000",
  6433=>"11111110",
  6434=>"11111110",
  6435=>"11111111",
  6436=>"00000001",
  6437=>"00000001",
  6438=>"11111111",
  6439=>"00000000",
  6440=>"00000010",
  6441=>"11111100",
  6442=>"00000001",
  6443=>"00000101",
  6444=>"11111100",
  6445=>"11111101",
  6446=>"00000001",
  6447=>"11111101",
  6448=>"11111110",
  6449=>"11111110",
  6450=>"00000000",
  6451=>"11111101",
  6452=>"11111101",
  6453=>"11111011",
  6454=>"00000001",
  6455=>"11111110",
  6456=>"11111110",
  6457=>"00000011",
  6458=>"11111110",
  6459=>"00000000",
  6460=>"00000000",
  6461=>"00000000",
  6462=>"00000010",
  6463=>"00000011",
  6464=>"00000011",
  6465=>"11111101",
  6466=>"11111111",
  6467=>"11111110",
  6468=>"00000000",
  6469=>"00000010",
  6470=>"00000010",
  6471=>"00000000",
  6472=>"00000011",
  6473=>"00000000",
  6474=>"00000000",
  6475=>"00000010",
  6476=>"00000001",
  6477=>"11111101",
  6478=>"11111110",
  6479=>"00000001",
  6480=>"11111110",
  6481=>"11111111",
  6482=>"00000010",
  6483=>"00000000",
  6484=>"11111111",
  6485=>"00000000",
  6486=>"00000000",
  6487=>"00000000",
  6488=>"00000011",
  6489=>"00000001",
  6490=>"11111101",
  6491=>"11111111",
  6492=>"11111111",
  6493=>"00000011",
  6494=>"11111111",
  6495=>"11111110",
  6496=>"11111100",
  6497=>"00000001",
  6498=>"00000000",
  6499=>"00000010",
  6500=>"11111111",
  6501=>"00000000",
  6502=>"00000000",
  6503=>"11111110",
  6504=>"00000101",
  6505=>"00000001",
  6506=>"11111101",
  6507=>"00000000",
  6508=>"00000011",
  6509=>"11111111",
  6510=>"11111110",
  6511=>"11111101",
  6512=>"00000000",
  6513=>"00000011",
  6514=>"00000000",
  6515=>"00000100",
  6516=>"11111111",
  6517=>"11111110",
  6518=>"00000000",
  6519=>"11111110",
  6520=>"00000100",
  6521=>"00000010",
  6522=>"00000000",
  6523=>"00000000",
  6524=>"00000000",
  6525=>"11111110",
  6526=>"00000000",
  6527=>"00000100",
  6528=>"00000001",
  6529=>"00000011",
  6530=>"11111111",
  6531=>"11111101",
  6532=>"00000000",
  6533=>"00000100",
  6534=>"11111101",
  6535=>"11111111",
  6536=>"00000000",
  6537=>"11111111",
  6538=>"11111100",
  6539=>"11111110",
  6540=>"00000000",
  6541=>"11111110",
  6542=>"11111111",
  6543=>"11111110",
  6544=>"11111110",
  6545=>"11111100",
  6546=>"11111100",
  6547=>"00000000",
  6548=>"11111110",
  6549=>"00000001",
  6550=>"00000001",
  6551=>"11111100",
  6552=>"11111101",
  6553=>"11111110",
  6554=>"11111111",
  6555=>"00000010",
  6556=>"11111111",
  6557=>"00000000",
  6558=>"11111110",
  6559=>"11111101",
  6560=>"00000010",
  6561=>"00000000",
  6562=>"11111101",
  6563=>"11111110",
  6564=>"11111111",
  6565=>"00000000",
  6566=>"00000010",
  6567=>"00000010",
  6568=>"00000100",
  6569=>"11111111",
  6570=>"11111101",
  6571=>"11111111",
  6572=>"00000011",
  6573=>"00000000",
  6574=>"00000000",
  6575=>"11111101",
  6576=>"00000001",
  6577=>"00000010",
  6578=>"00000001",
  6579=>"00000010",
  6580=>"11111111",
  6581=>"11111111",
  6582=>"00000001",
  6583=>"11111111",
  6584=>"00000010",
  6585=>"11111101",
  6586=>"00000000",
  6587=>"11111101",
  6588=>"00000010",
  6589=>"00000011",
  6590=>"11111100",
  6591=>"00000000",
  6592=>"00000000",
  6593=>"11111110",
  6594=>"00000001",
  6595=>"11111100",
  6596=>"00000011",
  6597=>"11111111",
  6598=>"00000010",
  6599=>"00000011",
  6600=>"11111101",
  6601=>"00000010",
  6602=>"11111111",
  6603=>"00000010",
  6604=>"11111110",
  6605=>"00000001",
  6606=>"11111110",
  6607=>"00000011",
  6608=>"00000000",
  6609=>"00000000",
  6610=>"00000000",
  6611=>"00000011",
  6612=>"00000010",
  6613=>"11111111",
  6614=>"00000000",
  6615=>"00000010",
  6616=>"00000001",
  6617=>"00000010",
  6618=>"00000010",
  6619=>"11111111",
  6620=>"11111111",
  6621=>"00000011",
  6622=>"00000101",
  6623=>"11111101",
  6624=>"11111111",
  6625=>"00000001",
  6626=>"11111110",
  6627=>"00000000",
  6628=>"00000010",
  6629=>"00000110",
  6630=>"11111101",
  6631=>"00000010",
  6632=>"00000100",
  6633=>"11111111",
  6634=>"00000001",
  6635=>"11111101",
  6636=>"11111111",
  6637=>"00000111",
  6638=>"11111100",
  6639=>"00000010",
  6640=>"00000001",
  6641=>"00000001",
  6642=>"00000001",
  6643=>"11111110",
  6644=>"11111100",
  6645=>"11111100",
  6646=>"00000011",
  6647=>"00000001",
  6648=>"00000001",
  6649=>"00000001",
  6650=>"00000100",
  6651=>"11111110",
  6652=>"00000000",
  6653=>"00000001",
  6654=>"11111101",
  6655=>"00000010",
  6656=>"11111111",
  6657=>"11111111",
  6658=>"00000001",
  6659=>"11111101",
  6660=>"11111111",
  6661=>"00000001",
  6662=>"11111111",
  6663=>"11111110",
  6664=>"11111110",
  6665=>"11111101",
  6666=>"11111111",
  6667=>"00000000",
  6668=>"00000100",
  6669=>"00000000",
  6670=>"11111101",
  6671=>"11111110",
  6672=>"00000011",
  6673=>"00000011",
  6674=>"11111111",
  6675=>"00000011",
  6676=>"00000100",
  6677=>"11111110",
  6678=>"11111111",
  6679=>"00000010",
  6680=>"00000011",
  6681=>"00000000",
  6682=>"00000010",
  6683=>"00000000",
  6684=>"11111111",
  6685=>"00000101",
  6686=>"00000000",
  6687=>"00000010",
  6688=>"11111110",
  6689=>"00000010",
  6690=>"11111100",
  6691=>"00000001",
  6692=>"11111111",
  6693=>"11111110",
  6694=>"00000010",
  6695=>"00000001",
  6696=>"11111110",
  6697=>"11111101",
  6698=>"00000011",
  6699=>"11111101",
  6700=>"00000000",
  6701=>"11111111",
  6702=>"11111111",
  6703=>"00000001",
  6704=>"11111101",
  6705=>"00000010",
  6706=>"11111111",
  6707=>"11111110",
  6708=>"11111111",
  6709=>"00000001",
  6710=>"00000010",
  6711=>"00000000",
  6712=>"00000000",
  6713=>"00000010",
  6714=>"00000011",
  6715=>"00000101",
  6716=>"00000000",
  6717=>"00000000",
  6718=>"00000001",
  6719=>"00000010",
  6720=>"11111111",
  6721=>"00000001",
  6722=>"11111111",
  6723=>"00000010",
  6724=>"00000010",
  6725=>"11111110",
  6726=>"11111111",
  6727=>"11111110",
  6728=>"11111111",
  6729=>"00000000",
  6730=>"11111110",
  6731=>"00000010",
  6732=>"00000001",
  6733=>"00000001",
  6734=>"00000000",
  6735=>"00000010",
  6736=>"00000001",
  6737=>"00000000",
  6738=>"00000010",
  6739=>"11111101",
  6740=>"00000001",
  6741=>"00000101",
  6742=>"00000000",
  6743=>"11111111",
  6744=>"11111111",
  6745=>"11111111",
  6746=>"11111101",
  6747=>"00000010",
  6748=>"00000011",
  6749=>"00000011",
  6750=>"00000001",
  6751=>"11111110",
  6752=>"00000010",
  6753=>"11111110",
  6754=>"11111110",
  6755=>"00000000",
  6756=>"00000000",
  6757=>"00000000",
  6758=>"00000001",
  6759=>"00000011",
  6760=>"00000010",
  6761=>"00000010",
  6762=>"00000010",
  6763=>"00000000",
  6764=>"00000010",
  6765=>"11111101",
  6766=>"11111110",
  6767=>"11111110",
  6768=>"00000101",
  6769=>"11111101",
  6770=>"11111111",
  6771=>"11111111",
  6772=>"00000011",
  6773=>"00000101",
  6774=>"00000010",
  6775=>"11111111",
  6776=>"11111110",
  6777=>"00000011",
  6778=>"11111111",
  6779=>"11111101",
  6780=>"00000001",
  6781=>"11111101",
  6782=>"11111110",
  6783=>"00000000",
  6784=>"11111110",
  6785=>"11111111",
  6786=>"00000011",
  6787=>"00000010",
  6788=>"00000011",
  6789=>"00000000",
  6790=>"00000011",
  6791=>"00000010",
  6792=>"00000000",
  6793=>"00000001",
  6794=>"11111111",
  6795=>"11111110",
  6796=>"00000010",
  6797=>"11111111",
  6798=>"11111110",
  6799=>"00000001",
  6800=>"00000001",
  6801=>"00000010",
  6802=>"00000000",
  6803=>"00000000",
  6804=>"00000001",
  6805=>"11111110",
  6806=>"00000010",
  6807=>"00000011",
  6808=>"11111101",
  6809=>"11111101",
  6810=>"00000010",
  6811=>"00000010",
  6812=>"00000000",
  6813=>"11111111",
  6814=>"11111110",
  6815=>"00000000",
  6816=>"00000001",
  6817=>"11111101",
  6818=>"11111101",
  6819=>"00000001",
  6820=>"00000010",
  6821=>"11111110",
  6822=>"00000000",
  6823=>"11111101",
  6824=>"00000011",
  6825=>"11111111",
  6826=>"11111110",
  6827=>"00000001",
  6828=>"00000011",
  6829=>"00000000",
  6830=>"00000000",
  6831=>"00000001",
  6832=>"11111110",
  6833=>"00000010",
  6834=>"11111110",
  6835=>"00000001",
  6836=>"00000100",
  6837=>"11111110",
  6838=>"00000000",
  6839=>"11111100",
  6840=>"11111111",
  6841=>"00000001",
  6842=>"11111101",
  6843=>"00000001",
  6844=>"00000010",
  6845=>"11111111",
  6846=>"11111110",
  6847=>"00000000",
  6848=>"11111111",
  6849=>"00000001",
  6850=>"11111101",
  6851=>"00000010",
  6852=>"00000011",
  6853=>"00000000",
  6854=>"11111101",
  6855=>"00000001",
  6856=>"00000010",
  6857=>"11111110",
  6858=>"11111101",
  6859=>"00000010",
  6860=>"00000101",
  6861=>"00000000",
  6862=>"00000000",
  6863=>"00000100",
  6864=>"00000000",
  6865=>"00000011",
  6866=>"00000010",
  6867=>"11111111",
  6868=>"00000010",
  6869=>"11111111",
  6870=>"00000000",
  6871=>"11111101",
  6872=>"00000010",
  6873=>"00000000",
  6874=>"00000001",
  6875=>"00000001",
  6876=>"00000010",
  6877=>"11111101",
  6878=>"11111101",
  6879=>"11111101",
  6880=>"00000011",
  6881=>"11111101",
  6882=>"11111101",
  6883=>"00000000",
  6884=>"00000000",
  6885=>"11111110",
  6886=>"11111110",
  6887=>"11111111",
  6888=>"11111111",
  6889=>"00000010",
  6890=>"11111111",
  6891=>"00000010",
  6892=>"11111111",
  6893=>"00000011",
  6894=>"00000010",
  6895=>"00000101",
  6896=>"00000001",
  6897=>"00000001",
  6898=>"11111110",
  6899=>"00000000",
  6900=>"11111101",
  6901=>"00000001",
  6902=>"00000010",
  6903=>"11111100",
  6904=>"11111110",
  6905=>"00000000",
  6906=>"00000001",
  6907=>"11111101",
  6908=>"00000000",
  6909=>"00000011",
  6910=>"11111100",
  6911=>"00000000",
  6912=>"11111101",
  6913=>"11111110",
  6914=>"11111110",
  6915=>"00000000",
  6916=>"11111111",
  6917=>"11111111",
  6918=>"11111101",
  6919=>"11111111",
  6920=>"11111011",
  6921=>"00000000",
  6922=>"00000000",
  6923=>"11111110",
  6924=>"11111101",
  6925=>"11111111",
  6926=>"11111100",
  6927=>"00000010",
  6928=>"11111101",
  6929=>"11111111",
  6930=>"11111111",
  6931=>"11111111",
  6932=>"00000011",
  6933=>"11111101",
  6934=>"11111111",
  6935=>"11111111",
  6936=>"00000001",
  6937=>"11111100",
  6938=>"11111110",
  6939=>"11111111",
  6940=>"00000001",
  6941=>"11111110",
  6942=>"00000011",
  6943=>"00000110",
  6944=>"00000001",
  6945=>"00000011",
  6946=>"11111111",
  6947=>"00000101",
  6948=>"11111111",
  6949=>"00000001",
  6950=>"11111110",
  6951=>"11111101",
  6952=>"11111101",
  6953=>"00000011",
  6954=>"00000000",
  6955=>"00000001",
  6956=>"11111111",
  6957=>"00000011",
  6958=>"11111101",
  6959=>"11111111",
  6960=>"00000010",
  6961=>"00000001",
  6962=>"00000000",
  6963=>"00000010",
  6964=>"00000010",
  6965=>"11111011",
  6966=>"11111101",
  6967=>"00000001",
  6968=>"11111101",
  6969=>"11111111",
  6970=>"00000110",
  6971=>"00000010",
  6972=>"00000010",
  6973=>"00000001",
  6974=>"00000010",
  6975=>"00000000",
  6976=>"00000010",
  6977=>"00000000",
  6978=>"11111111",
  6979=>"11111100",
  6980=>"00000100",
  6981=>"00000001",
  6982=>"11111111",
  6983=>"00000011",
  6984=>"00000000",
  6985=>"11111101",
  6986=>"11111110",
  6987=>"00000010",
  6988=>"00000010",
  6989=>"00000000",
  6990=>"11111110",
  6991=>"00000001",
  6992=>"11111110",
  6993=>"00000011",
  6994=>"00000001",
  6995=>"11111100",
  6996=>"00000010",
  6997=>"00000011",
  6998=>"00000001",
  6999=>"00000011",
  7000=>"11111101",
  7001=>"00000001",
  7002=>"00000011",
  7003=>"00000100",
  7004=>"00000000",
  7005=>"00000001",
  7006=>"11111110",
  7007=>"11111101",
  7008=>"11111100",
  7009=>"00000001",
  7010=>"11111110",
  7011=>"00000100",
  7012=>"00000000",
  7013=>"00000011",
  7014=>"00000010",
  7015=>"00000100",
  7016=>"00000100",
  7017=>"11111101",
  7018=>"00000010",
  7019=>"11111111",
  7020=>"00000011",
  7021=>"11111110",
  7022=>"11111110",
  7023=>"00000010",
  7024=>"11111101",
  7025=>"00000011",
  7026=>"00000010",
  7027=>"11111100",
  7028=>"00000010",
  7029=>"00000000",
  7030=>"11111101",
  7031=>"00000001",
  7032=>"11111110",
  7033=>"00000101",
  7034=>"00000000",
  7035=>"11111111",
  7036=>"00000000",
  7037=>"11111100",
  7038=>"00000000",
  7039=>"00000001",
  7040=>"00000010",
  7041=>"11111101",
  7042=>"00000001",
  7043=>"11111101",
  7044=>"00000011",
  7045=>"00000000",
  7046=>"11111101",
  7047=>"11111111",
  7048=>"00000001",
  7049=>"00000011",
  7050=>"00000010",
  7051=>"11111111",
  7052=>"11111100",
  7053=>"11111110",
  7054=>"11111110",
  7055=>"11111101",
  7056=>"11111101",
  7057=>"11111110",
  7058=>"11111100",
  7059=>"00000001",
  7060=>"00000011",
  7061=>"11111101",
  7062=>"00000000",
  7063=>"11111101",
  7064=>"00000011",
  7065=>"00000010",
  7066=>"11111111",
  7067=>"00000001",
  7068=>"00000000",
  7069=>"00000000",
  7070=>"11111110",
  7071=>"11111111",
  7072=>"11111111",
  7073=>"00000010",
  7074=>"11111111",
  7075=>"11111110",
  7076=>"11111111",
  7077=>"00000010",
  7078=>"00000001",
  7079=>"11111011",
  7080=>"00000000",
  7081=>"00000001",
  7082=>"11111111",
  7083=>"00000000",
  7084=>"00000000",
  7085=>"00000001",
  7086=>"00000010",
  7087=>"00000011",
  7088=>"11111110",
  7089=>"00000010",
  7090=>"00000000",
  7091=>"11111100",
  7092=>"00000010",
  7093=>"11111110",
  7094=>"11111101",
  7095=>"00000100",
  7096=>"00000001",
  7097=>"00000010",
  7098=>"00000000",
  7099=>"00000011",
  7100=>"11111101",
  7101=>"00000001",
  7102=>"11111111",
  7103=>"00000001",
  7104=>"11111111",
  7105=>"00000001",
  7106=>"00000010",
  7107=>"00000010",
  7108=>"11111110",
  7109=>"11111111",
  7110=>"00000100",
  7111=>"00000001",
  7112=>"00000010",
  7113=>"11111111",
  7114=>"00000000",
  7115=>"00000001",
  7116=>"11111110",
  7117=>"11111101",
  7118=>"11111111",
  7119=>"11111111",
  7120=>"00000010",
  7121=>"00000110",
  7122=>"11111110",
  7123=>"00000011",
  7124=>"11111101",
  7125=>"11111111",
  7126=>"11111111",
  7127=>"00000000",
  7128=>"11111110",
  7129=>"11111011",
  7130=>"00000000",
  7131=>"11111110",
  7132=>"00000010",
  7133=>"00000010",
  7134=>"11111101",
  7135=>"00000000",
  7136=>"00000000",
  7137=>"00000010",
  7138=>"00000011",
  7139=>"00000001",
  7140=>"11111111",
  7141=>"00000110",
  7142=>"00000000",
  7143=>"11111101",
  7144=>"11111110",
  7145=>"00000010",
  7146=>"00000011",
  7147=>"11111111",
  7148=>"00000100",
  7149=>"11111110",
  7150=>"00000001",
  7151=>"00000001",
  7152=>"00000000",
  7153=>"11111101",
  7154=>"00000000",
  7155=>"11111111",
  7156=>"11111111",
  7157=>"11111101",
  7158=>"00000011",
  7159=>"00000011",
  7160=>"11111101",
  7161=>"11111111",
  7162=>"11111101",
  7163=>"00000100",
  7164=>"11111111",
  7165=>"11111110",
  7166=>"00000100",
  7167=>"00000100",
  7168=>"00000100",
  7169=>"00000010",
  7170=>"00000011",
  7171=>"11111110",
  7172=>"00000010",
  7173=>"11111101",
  7174=>"00000000",
  7175=>"00000100",
  7176=>"11111110",
  7177=>"11111101",
  7178=>"11111111",
  7179=>"11111110",
  7180=>"00000001",
  7181=>"00000110",
  7182=>"00000011",
  7183=>"00000000",
  7184=>"00000111",
  7185=>"00000000",
  7186=>"00000000",
  7187=>"11111110",
  7188=>"00000001",
  7189=>"00000010",
  7190=>"00000000",
  7191=>"00000010",
  7192=>"11111110",
  7193=>"11111101",
  7194=>"00000000",
  7195=>"00000011",
  7196=>"00000000",
  7197=>"11111111",
  7198=>"11111111",
  7199=>"00000011",
  7200=>"11111101",
  7201=>"11111111",
  7202=>"00000010",
  7203=>"11111100",
  7204=>"11111110",
  7205=>"11111101",
  7206=>"11111111",
  7207=>"00000001",
  7208=>"11111110",
  7209=>"11111110",
  7210=>"00000001",
  7211=>"00000000",
  7212=>"11111101",
  7213=>"00000010",
  7214=>"00000011",
  7215=>"11111110",
  7216=>"11111111",
  7217=>"00000010",
  7218=>"00000001",
  7219=>"00000000",
  7220=>"00000000",
  7221=>"00000011",
  7222=>"11111110",
  7223=>"00000011",
  7224=>"11111101",
  7225=>"00000010",
  7226=>"00000000",
  7227=>"00000001",
  7228=>"11111101",
  7229=>"11111101",
  7230=>"11111110",
  7231=>"11111110",
  7232=>"00000000",
  7233=>"00000100",
  7234=>"11111111",
  7235=>"00000010",
  7236=>"00000100",
  7237=>"11111111",
  7238=>"00000000",
  7239=>"11111101",
  7240=>"00000010",
  7241=>"11111101",
  7242=>"00000000",
  7243=>"00000011",
  7244=>"00000100",
  7245=>"11111111",
  7246=>"11111110",
  7247=>"00000001",
  7248=>"11111011",
  7249=>"00000011",
  7250=>"11111111",
  7251=>"11111111",
  7252=>"00000000",
  7253=>"00000010",
  7254=>"11111101",
  7255=>"00000011",
  7256=>"00000000",
  7257=>"00000011",
  7258=>"00000000",
  7259=>"00000000",
  7260=>"00000001",
  7261=>"00000010",
  7262=>"00000001",
  7263=>"00000100",
  7264=>"00000001",
  7265=>"11111100",
  7266=>"11111111",
  7267=>"11111111",
  7268=>"11111110",
  7269=>"00000011",
  7270=>"11111111",
  7271=>"11111101",
  7272=>"00000110",
  7273=>"00000010",
  7274=>"00000110",
  7275=>"00000001",
  7276=>"00000000",
  7277=>"11111100",
  7278=>"00000000",
  7279=>"00000001",
  7280=>"00000011",
  7281=>"00000101",
  7282=>"00000011",
  7283=>"00000001",
  7284=>"00000000",
  7285=>"00000101",
  7286=>"11111111",
  7287=>"00000010",
  7288=>"11111111",
  7289=>"00000001",
  7290=>"11111110",
  7291=>"00000101",
  7292=>"00000000",
  7293=>"00000011",
  7294=>"00000011",
  7295=>"11111101",
  7296=>"00000100",
  7297=>"11111100",
  7298=>"11111111",
  7299=>"11111110",
  7300=>"11111110",
  7301=>"11111101",
  7302=>"11111111",
  7303=>"11111100",
  7304=>"11111100",
  7305=>"00000000",
  7306=>"00000010",
  7307=>"11111110",
  7308=>"11111110",
  7309=>"11111110",
  7310=>"00000001",
  7311=>"11111111",
  7312=>"11111100",
  7313=>"00000001",
  7314=>"00000100",
  7315=>"00000001",
  7316=>"00000001",
  7317=>"11111111",
  7318=>"00000000",
  7319=>"00000000",
  7320=>"11111111",
  7321=>"00000100",
  7322=>"00000011",
  7323=>"00000000",
  7324=>"00000010",
  7325=>"11111110",
  7326=>"00000011",
  7327=>"11111111",
  7328=>"11111111",
  7329=>"00000001",
  7330=>"00000110",
  7331=>"11111111",
  7332=>"11111111",
  7333=>"11111111",
  7334=>"00000000",
  7335=>"11111111",
  7336=>"00000000",
  7337=>"11111111",
  7338=>"00000010",
  7339=>"00000011",
  7340=>"11111110",
  7341=>"11111110",
  7342=>"11111101",
  7343=>"00000001",
  7344=>"00000001",
  7345=>"11111101",
  7346=>"11111110",
  7347=>"11111110",
  7348=>"11111111",
  7349=>"11111111",
  7350=>"00000010",
  7351=>"00000000",
  7352=>"11111110",
  7353=>"11111110",
  7354=>"00000000",
  7355=>"00000011",
  7356=>"00000010",
  7357=>"11111110",
  7358=>"00000000",
  7359=>"00000010",
  7360=>"00000010",
  7361=>"00000000",
  7362=>"00000001",
  7363=>"11111100",
  7364=>"11111111",
  7365=>"00000100",
  7366=>"11111110",
  7367=>"00000011",
  7368=>"11111111",
  7369=>"11111101",
  7370=>"00000001",
  7371=>"00000010",
  7372=>"00000010",
  7373=>"00000101",
  7374=>"11111111",
  7375=>"00000000",
  7376=>"11111011",
  7377=>"11111101",
  7378=>"00000001",
  7379=>"00000000",
  7380=>"00000011",
  7381=>"11111110",
  7382=>"11111101",
  7383=>"11111101",
  7384=>"00000001",
  7385=>"00000001",
  7386=>"11111110",
  7387=>"00000000",
  7388=>"00000010",
  7389=>"00000000",
  7390=>"00000011",
  7391=>"11111111",
  7392=>"00000101",
  7393=>"00000000",
  7394=>"00000000",
  7395=>"00000001",
  7396=>"11111110",
  7397=>"00000011",
  7398=>"00000000",
  7399=>"11111111",
  7400=>"11111101",
  7401=>"00000000",
  7402=>"11111101",
  7403=>"00000001",
  7404=>"11111110",
  7405=>"00000001",
  7406=>"11111100",
  7407=>"11111110",
  7408=>"00000011",
  7409=>"00000100",
  7410=>"00000000",
  7411=>"00000001",
  7412=>"11111011",
  7413=>"00000001",
  7414=>"11111100",
  7415=>"11111111",
  7416=>"11111101",
  7417=>"11111110",
  7418=>"00000000",
  7419=>"00000011",
  7420=>"00000001",
  7421=>"11111111",
  7422=>"11111111",
  7423=>"00000001",
  7424=>"00000010",
  7425=>"00000000",
  7426=>"11111111",
  7427=>"00000000",
  7428=>"11111111",
  7429=>"00000000",
  7430=>"11111100",
  7431=>"00000000",
  7432=>"00000010",
  7433=>"00000000",
  7434=>"11111011",
  7435=>"00000100",
  7436=>"00000011",
  7437=>"11111110",
  7438=>"11111100",
  7439=>"00000000",
  7440=>"11111110",
  7441=>"00000000",
  7442=>"00000001",
  7443=>"11111100",
  7444=>"11111111",
  7445=>"00000011",
  7446=>"00000101",
  7447=>"00000001",
  7448=>"00000011",
  7449=>"11111101",
  7450=>"00000010",
  7451=>"00000010",
  7452=>"11111110",
  7453=>"00000100",
  7454=>"00000001",
  7455=>"00000111",
  7456=>"00000000",
  7457=>"00000000",
  7458=>"00000000",
  7459=>"00000011",
  7460=>"11111110",
  7461=>"00000001",
  7462=>"00000100",
  7463=>"00000011",
  7464=>"00000100",
  7465=>"00000001",
  7466=>"00000010",
  7467=>"00000001",
  7468=>"11111101",
  7469=>"11111101",
  7470=>"00000000",
  7471=>"11111110",
  7472=>"00000011",
  7473=>"00000101",
  7474=>"11111110",
  7475=>"00000000",
  7476=>"00000000",
  7477=>"11111011",
  7478=>"00000010",
  7479=>"11111111",
  7480=>"11111100",
  7481=>"11111111",
  7482=>"11111101",
  7483=>"00000001",
  7484=>"11111110",
  7485=>"11111111",
  7486=>"00000011",
  7487=>"00000001",
  7488=>"11111101",
  7489=>"11111111",
  7490=>"11111111",
  7491=>"11111111",
  7492=>"00000011",
  7493=>"00000101",
  7494=>"11111101",
  7495=>"00000100",
  7496=>"00000010",
  7497=>"11111110",
  7498=>"00000000",
  7499=>"00000101",
  7500=>"11111101",
  7501=>"11111100",
  7502=>"00000011",
  7503=>"00000100",
  7504=>"11111101",
  7505=>"11111110",
  7506=>"11111100",
  7507=>"00000011",
  7508=>"11111111",
  7509=>"00000100",
  7510=>"00000001",
  7511=>"00000010",
  7512=>"00000000",
  7513=>"11111111",
  7514=>"11111110",
  7515=>"11111111",
  7516=>"00000010",
  7517=>"00000011",
  7518=>"11111100",
  7519=>"00000011",
  7520=>"11111110",
  7521=>"00000001",
  7522=>"11111101",
  7523=>"11111111",
  7524=>"00000001",
  7525=>"00000000",
  7526=>"11111101",
  7527=>"11111111",
  7528=>"00000000",
  7529=>"00000100",
  7530=>"00000100",
  7531=>"00000010",
  7532=>"00000010",
  7533=>"00000011",
  7534=>"00000001",
  7535=>"11111101",
  7536=>"11111111",
  7537=>"11111111",
  7538=>"00000001",
  7539=>"00000000",
  7540=>"00000001",
  7541=>"00000000",
  7542=>"11111101",
  7543=>"00000010",
  7544=>"11111111",
  7545=>"11111100",
  7546=>"00000000",
  7547=>"11111101",
  7548=>"11111101",
  7549=>"00000000",
  7550=>"11111101",
  7551=>"11111101",
  7552=>"00000100",
  7553=>"11111101",
  7554=>"11111111",
  7555=>"11111111",
  7556=>"00000000",
  7557=>"11111111",
  7558=>"00000001",
  7559=>"11111101",
  7560=>"11111110",
  7561=>"00000011",
  7562=>"00000010",
  7563=>"11111100",
  7564=>"00000001",
  7565=>"11111111",
  7566=>"11111100",
  7567=>"00000011",
  7568=>"11111111",
  7569=>"00000111",
  7570=>"00000000",
  7571=>"00000010",
  7572=>"00000011",
  7573=>"11111110",
  7574=>"00000010",
  7575=>"11111111",
  7576=>"11111111",
  7577=>"11111101",
  7578=>"00000001",
  7579=>"00000000",
  7580=>"11111110",
  7581=>"00000010",
  7582=>"00000100",
  7583=>"11111111",
  7584=>"00000001",
  7585=>"11111100",
  7586=>"00000101",
  7587=>"11111110",
  7588=>"11111111",
  7589=>"00000010",
  7590=>"00000001",
  7591=>"00000010",
  7592=>"11111101",
  7593=>"00000011",
  7594=>"00000011",
  7595=>"00000010",
  7596=>"00000010",
  7597=>"00000010",
  7598=>"00000010",
  7599=>"11111110",
  7600=>"00000001",
  7601=>"11111100",
  7602=>"11111101",
  7603=>"00000010",
  7604=>"11111111",
  7605=>"00000011",
  7606=>"00000110",
  7607=>"00001000",
  7608=>"00000110",
  7609=>"11111111",
  7610=>"11111110",
  7611=>"11111110",
  7612=>"00000011",
  7613=>"11111101",
  7614=>"00000010",
  7615=>"00000001",
  7616=>"00000000",
  7617=>"11111110",
  7618=>"00000100",
  7619=>"00000001",
  7620=>"00000010",
  7621=>"11111110",
  7622=>"11111110",
  7623=>"11111101",
  7624=>"00000011",
  7625=>"00000101",
  7626=>"00000011",
  7627=>"00000010",
  7628=>"00000010",
  7629=>"00000000",
  7630=>"11111101",
  7631=>"11111101",
  7632=>"00000001",
  7633=>"11111111",
  7634=>"00000010",
  7635=>"00000100",
  7636=>"11111101",
  7637=>"00000001",
  7638=>"00000001",
  7639=>"11111101",
  7640=>"00000000",
  7641=>"00000001",
  7642=>"11111111",
  7643=>"00000001",
  7644=>"00000000",
  7645=>"00000100",
  7646=>"00000010",
  7647=>"00000001",
  7648=>"11111110",
  7649=>"00000100",
  7650=>"00000000",
  7651=>"11111111",
  7652=>"11111110",
  7653=>"11111111",
  7654=>"11111101",
  7655=>"11111110",
  7656=>"11111111",
  7657=>"11111111",
  7658=>"00000010",
  7659=>"00000111",
  7660=>"00000100",
  7661=>"00000001",
  7662=>"11111110",
  7663=>"11111101",
  7664=>"11111110",
  7665=>"11111101",
  7666=>"11111110",
  7667=>"11111101",
  7668=>"11111101",
  7669=>"11111100",
  7670=>"00000000",
  7671=>"11111110",
  7672=>"00000001",
  7673=>"00000011",
  7674=>"00000010",
  7675=>"00000100",
  7676=>"00000011",
  7677=>"00000001",
  7678=>"00000000",
  7679=>"00000110",
  7680=>"11111111",
  7681=>"00000011",
  7682=>"11111110",
  7683=>"00000000",
  7684=>"11111110",
  7685=>"00000001",
  7686=>"00000000",
  7687=>"00000101",
  7688=>"00000010",
  7689=>"00000001",
  7690=>"00000011",
  7691=>"00000000",
  7692=>"11111111",
  7693=>"11111111",
  7694=>"00000001",
  7695=>"00000010",
  7696=>"11111111",
  7697=>"11111100",
  7698=>"00000011",
  7699=>"11111101",
  7700=>"11111101",
  7701=>"11111110",
  7702=>"00000000",
  7703=>"11111111",
  7704=>"00000011",
  7705=>"00000001",
  7706=>"00000000",
  7707=>"00000010",
  7708=>"00000001",
  7709=>"11111100",
  7710=>"11111111",
  7711=>"00000101",
  7712=>"00000100",
  7713=>"00000010",
  7714=>"11111111",
  7715=>"00000000",
  7716=>"11111101",
  7717=>"11111101",
  7718=>"11111110",
  7719=>"00000001",
  7720=>"00000000",
  7721=>"11111101",
  7722=>"11111100",
  7723=>"00000010",
  7724=>"11111110",
  7725=>"11111101",
  7726=>"11111111",
  7727=>"11111110",
  7728=>"11111110",
  7729=>"00000000",
  7730=>"00000001",
  7731=>"11111110",
  7732=>"00000001",
  7733=>"00000000",
  7734=>"00000100",
  7735=>"11111111",
  7736=>"11111111",
  7737=>"11111111",
  7738=>"00000100",
  7739=>"11111101",
  7740=>"11111111",
  7741=>"11111111",
  7742=>"11111011",
  7743=>"11111110",
  7744=>"11111101",
  7745=>"00000010",
  7746=>"00000100",
  7747=>"11111110",
  7748=>"00000001",
  7749=>"11111101",
  7750=>"11111110",
  7751=>"11111111",
  7752=>"00000000",
  7753=>"00000001",
  7754=>"11111110",
  7755=>"00000001",
  7756=>"00000000",
  7757=>"00000010",
  7758=>"11111100",
  7759=>"00000011",
  7760=>"11111111",
  7761=>"00000011",
  7762=>"11111110",
  7763=>"00000011",
  7764=>"11111101",
  7765=>"11111100",
  7766=>"11111111",
  7767=>"11111111",
  7768=>"11111111",
  7769=>"11111111",
  7770=>"00000010",
  7771=>"00000010",
  7772=>"00000011",
  7773=>"00000010",
  7774=>"11111111",
  7775=>"00000100",
  7776=>"11111110",
  7777=>"00000101",
  7778=>"11111110",
  7779=>"00000101",
  7780=>"00000010",
  7781=>"11111111",
  7782=>"11111110",
  7783=>"00000000",
  7784=>"00000100",
  7785=>"00000010",
  7786=>"00000001",
  7787=>"00000010",
  7788=>"00000001",
  7789=>"00000011",
  7790=>"11111111",
  7791=>"00000010",
  7792=>"00000000",
  7793=>"00000001",
  7794=>"00000010",
  7795=>"00000001",
  7796=>"00000100",
  7797=>"11111011",
  7798=>"11111101",
  7799=>"11111100",
  7800=>"00000000",
  7801=>"00000001",
  7802=>"11111100",
  7803=>"11111100",
  7804=>"11111111",
  7805=>"11111101",
  7806=>"11111101",
  7807=>"00000000",
  7808=>"11111110",
  7809=>"11111101",
  7810=>"00000001",
  7811=>"11111110",
  7812=>"00000100",
  7813=>"00000110",
  7814=>"11111110",
  7815=>"00000100",
  7816=>"00000000",
  7817=>"11111110",
  7818=>"11111100",
  7819=>"00000101",
  7820=>"00000011",
  7821=>"00000001",
  7822=>"00000011",
  7823=>"11111111",
  7824=>"11111110",
  7825=>"11111111",
  7826=>"00000010",
  7827=>"11111110",
  7828=>"00000001",
  7829=>"00000001",
  7830=>"11111111",
  7831=>"00000010",
  7832=>"00000000",
  7833=>"00000000",
  7834=>"00000110",
  7835=>"00000011",
  7836=>"00000010",
  7837=>"00000010",
  7838=>"00000001",
  7839=>"00000010",
  7840=>"11111111",
  7841=>"00000111",
  7842=>"00000010",
  7843=>"11111100",
  7844=>"00000001",
  7845=>"11111110",
  7846=>"00000001",
  7847=>"11111111",
  7848=>"11111111",
  7849=>"00000011",
  7850=>"00000000",
  7851=>"11111110",
  7852=>"00000011",
  7853=>"00000101",
  7854=>"00000001",
  7855=>"00000110",
  7856=>"00000100",
  7857=>"11111110",
  7858=>"11111100",
  7859=>"11111111",
  7860=>"11111110",
  7861=>"00000000",
  7862=>"11111100",
  7863=>"11111111",
  7864=>"00000000",
  7865=>"00000100",
  7866=>"00000000",
  7867=>"11111111",
  7868=>"00000011",
  7869=>"00000001",
  7870=>"11111110",
  7871=>"11111110",
  7872=>"11111110",
  7873=>"11111110",
  7874=>"11111110",
  7875=>"11111100",
  7876=>"00000001",
  7877=>"11111101",
  7878=>"00000000",
  7879=>"00000011",
  7880=>"00000101",
  7881=>"11111110",
  7882=>"11111110",
  7883=>"00000001",
  7884=>"11111110",
  7885=>"00000010",
  7886=>"00000000",
  7887=>"11111110",
  7888=>"00000010",
  7889=>"00000000",
  7890=>"00000000",
  7891=>"11111100",
  7892=>"00000010",
  7893=>"00000000",
  7894=>"11111111",
  7895=>"00000001",
  7896=>"00000000",
  7897=>"00000011",
  7898=>"11111110",
  7899=>"11111100",
  7900=>"00000000",
  7901=>"11111110",
  7902=>"00000000",
  7903=>"11111101",
  7904=>"11111110",
  7905=>"00000000",
  7906=>"00000000",
  7907=>"00000010",
  7908=>"00000010",
  7909=>"00000001",
  7910=>"00000000",
  7911=>"00000010",
  7912=>"11111110",
  7913=>"00000000",
  7914=>"00000001",
  7915=>"00000001",
  7916=>"11111111",
  7917=>"00000001",
  7918=>"11111111",
  7919=>"11111101",
  7920=>"11111111",
  7921=>"00000011",
  7922=>"11111100",
  7923=>"00000000",
  7924=>"11111110",
  7925=>"00000010",
  7926=>"00000011",
  7927=>"00000010",
  7928=>"00000001",
  7929=>"11111111",
  7930=>"00000101",
  7931=>"11111101",
  7932=>"00000000",
  7933=>"11111110",
  7934=>"11111100",
  7935=>"00000010",
  7936=>"11111110",
  7937=>"00000010",
  7938=>"11111111",
  7939=>"00000001",
  7940=>"11111100",
  7941=>"11111101",
  7942=>"00000001",
  7943=>"11111101",
  7944=>"00000011",
  7945=>"11111110",
  7946=>"00000010",
  7947=>"00000011",
  7948=>"11111110",
  7949=>"00000011",
  7950=>"00000001",
  7951=>"00000001",
  7952=>"00000011",
  7953=>"00000111",
  7954=>"00000010",
  7955=>"11111110",
  7956=>"00000000",
  7957=>"00000101",
  7958=>"00000010",
  7959=>"11111110",
  7960=>"00000001",
  7961=>"00000010",
  7962=>"11111110",
  7963=>"11111101",
  7964=>"11111111",
  7965=>"00000000",
  7966=>"00000011",
  7967=>"11111110",
  7968=>"11111101",
  7969=>"11111110",
  7970=>"00000001",
  7971=>"11111110",
  7972=>"11111110",
  7973=>"11111110",
  7974=>"00000010",
  7975=>"11111101",
  7976=>"11111111",
  7977=>"11111101",
  7978=>"00000110",
  7979=>"00000010",
  7980=>"11111111",
  7981=>"00000001",
  7982=>"00000100",
  7983=>"11111100",
  7984=>"00000011",
  7985=>"11111111",
  7986=>"11111101",
  7987=>"11111110",
  7988=>"00000000",
  7989=>"11111110",
  7990=>"00000000",
  7991=>"11111111",
  7992=>"00000011",
  7993=>"00000011",
  7994=>"11111110",
  7995=>"00000001",
  7996=>"00000000",
  7997=>"11111111",
  7998=>"00000010",
  7999=>"11111111",
  8000=>"11111110",
  8001=>"11111101",
  8002=>"00000001",
  8003=>"00000000",
  8004=>"11111101",
  8005=>"11111110",
  8006=>"00000010",
  8007=>"00000001",
  8008=>"00000001",
  8009=>"00000010",
  8010=>"00000101",
  8011=>"00000010",
  8012=>"00000000",
  8013=>"00000010",
  8014=>"00000000",
  8015=>"11111111",
  8016=>"11111111",
  8017=>"00000110",
  8018=>"11111110",
  8019=>"00000011",
  8020=>"11111100",
  8021=>"00000010",
  8022=>"11111110",
  8023=>"00000010",
  8024=>"00000010",
  8025=>"11111111",
  8026=>"11111101",
  8027=>"00000100",
  8028=>"00000001",
  8029=>"00000000",
  8030=>"11111110",
  8031=>"00000101",
  8032=>"00000010",
  8033=>"00000001",
  8034=>"00000000",
  8035=>"00000101",
  8036=>"00000001",
  8037=>"11111110",
  8038=>"11111110",
  8039=>"11111101",
  8040=>"11111110",
  8041=>"11111101",
  8042=>"00000100",
  8043=>"00000100",
  8044=>"11111110",
  8045=>"00000001",
  8046=>"00000011",
  8047=>"00000000",
  8048=>"00000001",
  8049=>"11111111",
  8050=>"11111111",
  8051=>"00000001",
  8052=>"11111110",
  8053=>"11111110",
  8054=>"00000001",
  8055=>"00000010",
  8056=>"00000101",
  8057=>"00000100",
  8058=>"00000011",
  8059=>"11111101",
  8060=>"00000000",
  8061=>"11111100",
  8062=>"00000000",
  8063=>"11111110",
  8064=>"11111111",
  8065=>"00000010",
  8066=>"11111110",
  8067=>"00000011",
  8068=>"00000000",
  8069=>"00000001",
  8070=>"00000010",
  8071=>"00000010",
  8072=>"00000010",
  8073=>"00000010",
  8074=>"11111110",
  8075=>"11111101",
  8076=>"00000001",
  8077=>"11111110",
  8078=>"00000101",
  8079=>"11111110",
  8080=>"00000010",
  8081=>"00000001",
  8082=>"00000101",
  8083=>"00000010",
  8084=>"11111100",
  8085=>"00000000",
  8086=>"00000001",
  8087=>"00000011",
  8088=>"11111110",
  8089=>"00000000",
  8090=>"11111101",
  8091=>"00000011",
  8092=>"00000001",
  8093=>"00000000",
  8094=>"00000100",
  8095=>"00000010",
  8096=>"11111110",
  8097=>"11111101",
  8098=>"00000001",
  8099=>"00000001",
  8100=>"00000001",
  8101=>"11111110",
  8102=>"11111101",
  8103=>"00000000",
  8104=>"00000000",
  8105=>"11111110",
  8106=>"00000000",
  8107=>"00000011",
  8108=>"11111111",
  8109=>"11111101",
  8110=>"11111100",
  8111=>"11111101",
  8112=>"00000100",
  8113=>"00000011",
  8114=>"11111101",
  8115=>"11111101",
  8116=>"00000000",
  8117=>"00000011",
  8118=>"00000000",
  8119=>"00000001",
  8120=>"11111110",
  8121=>"11111111",
  8122=>"00000000",
  8123=>"00000010",
  8124=>"00000001",
  8125=>"00000000",
  8126=>"00000000",
  8127=>"11111111",
  8128=>"00000010",
  8129=>"00000001",
  8130=>"00000010",
  8131=>"11111101",
  8132=>"11111111",
  8133=>"00000001",
  8134=>"00000011",
  8135=>"00000010",
  8136=>"00000011",
  8137=>"11111101",
  8138=>"00000000",
  8139=>"11111110",
  8140=>"11111110",
  8141=>"00000001",
  8142=>"00000011",
  8143=>"11111111",
  8144=>"11111111",
  8145=>"00000010",
  8146=>"00000001",
  8147=>"11111100",
  8148=>"00000010",
  8149=>"00000100",
  8150=>"00000001",
  8151=>"00000010",
  8152=>"11111111",
  8153=>"11111101",
  8154=>"00000000",
  8155=>"11111110",
  8156=>"00000100",
  8157=>"11111110",
  8158=>"00000000",
  8159=>"11111111",
  8160=>"11111100",
  8161=>"11111101",
  8162=>"00000000",
  8163=>"00000001",
  8164=>"00000010",
  8165=>"00000000",
  8166=>"11111111",
  8167=>"00000010",
  8168=>"11111111",
  8169=>"00000001",
  8170=>"11111100",
  8171=>"00000011",
  8172=>"11111101",
  8173=>"00000010",
  8174=>"00000001",
  8175=>"00000100",
  8176=>"11111111",
  8177=>"11111110",
  8178=>"00000000",
  8179=>"11111100",
  8180=>"00000010",
  8181=>"00000000",
  8182=>"00000010",
  8183=>"11111100",
  8184=>"00000110",
  8185=>"11111111",
  8186=>"00000011",
  8187=>"00000011",
  8188=>"00000001",
  8189=>"00000111",
  8190=>"11111111",
  8191=>"00000000",
  8192=>"11111101",
  8193=>"00000001",
  8194=>"00000100",
  8195=>"00000010",
  8196=>"00000110",
  8197=>"11111100",
  8198=>"00000000",
  8199=>"11111111",
  8200=>"00000011",
  8201=>"00000000",
  8202=>"11111111",
  8203=>"00000010",
  8204=>"00000000",
  8205=>"00000001",
  8206=>"00000001",
  8207=>"11111100",
  8208=>"00000010",
  8209=>"11111110",
  8210=>"11111011",
  8211=>"11111111",
  8212=>"00000010",
  8213=>"00000010",
  8214=>"00000001",
  8215=>"00000000",
  8216=>"11111110",
  8217=>"11111110",
  8218=>"00000001",
  8219=>"00000001",
  8220=>"11111101",
  8221=>"00000001",
  8222=>"11111101",
  8223=>"11111110",
  8224=>"11111111",
  8225=>"11111110",
  8226=>"00000011",
  8227=>"11111110",
  8228=>"11111101",
  8229=>"11111111",
  8230=>"00000001",
  8231=>"00000000",
  8232=>"11111101",
  8233=>"00000011",
  8234=>"00000000",
  8235=>"00000001",
  8236=>"00000000",
  8237=>"00000011",
  8238=>"00000000",
  8239=>"11111111",
  8240=>"11111111",
  8241=>"00000010",
  8242=>"00000011",
  8243=>"00000010",
  8244=>"00000000",
  8245=>"00000010",
  8246=>"00000000",
  8247=>"00000011",
  8248=>"00000010",
  8249=>"00000010",
  8250=>"11111111",
  8251=>"00000100",
  8252=>"00000000",
  8253=>"00000001",
  8254=>"00000000",
  8255=>"00000100",
  8256=>"00000100",
  8257=>"00000011",
  8258=>"11111110",
  8259=>"00000011",
  8260=>"11111101",
  8261=>"00000001",
  8262=>"00000000",
  8263=>"11111111",
  8264=>"00000010",
  8265=>"11111100",
  8266=>"11111101",
  8267=>"00000001",
  8268=>"11111101",
  8269=>"00000101",
  8270=>"00000011",
  8271=>"11111101",
  8272=>"00000000",
  8273=>"00000010",
  8274=>"11111101",
  8275=>"11111101",
  8276=>"00000000",
  8277=>"00000001",
  8278=>"00000010",
  8279=>"00000000",
  8280=>"00000001",
  8281=>"00000000",
  8282=>"11111110",
  8283=>"11111101",
  8284=>"11111100",
  8285=>"00000010",
  8286=>"00000010",
  8287=>"00000001",
  8288=>"11111111",
  8289=>"11111101",
  8290=>"00000000",
  8291=>"00000010",
  8292=>"00000111",
  8293=>"11111110",
  8294=>"11111111",
  8295=>"00000010",
  8296=>"11111110",
  8297=>"00000010",
  8298=>"11111110",
  8299=>"11111100",
  8300=>"11111110",
  8301=>"11111101",
  8302=>"11111110",
  8303=>"00000010",
  8304=>"00000111",
  8305=>"00000000",
  8306=>"11111101",
  8307=>"00000001",
  8308=>"00000110",
  8309=>"11111100",
  8310=>"00000011",
  8311=>"11111111",
  8312=>"00000000",
  8313=>"11111110",
  8314=>"11111111",
  8315=>"00000001",
  8316=>"00000011",
  8317=>"00000010",
  8318=>"11111111",
  8319=>"00000100",
  8320=>"00000010",
  8321=>"00000011",
  8322=>"00000000",
  8323=>"00000001",
  8324=>"00000100",
  8325=>"00000100",
  8326=>"00000000",
  8327=>"11111100",
  8328=>"00000001",
  8329=>"00000101",
  8330=>"11111110",
  8331=>"00000100",
  8332=>"11111110",
  8333=>"00000000",
  8334=>"00000000",
  8335=>"11111100",
  8336=>"00000010",
  8337=>"00000011",
  8338=>"00000000",
  8339=>"00000100",
  8340=>"00000010",
  8341=>"11111110",
  8342=>"11111111",
  8343=>"11111110",
  8344=>"00000001",
  8345=>"00000100",
  8346=>"00000000",
  8347=>"11111100",
  8348=>"00000001",
  8349=>"00000110",
  8350=>"11111100",
  8351=>"00000000",
  8352=>"00000010",
  8353=>"00000001",
  8354=>"11111101",
  8355=>"11111111",
  8356=>"00000000",
  8357=>"00000011",
  8358=>"00000001",
  8359=>"11111101",
  8360=>"00000001",
  8361=>"00000001",
  8362=>"00000010",
  8363=>"00000010",
  8364=>"11111100",
  8365=>"00000001",
  8366=>"00000100",
  8367=>"11111110",
  8368=>"11111110",
  8369=>"11111111",
  8370=>"11111101",
  8371=>"00000110",
  8372=>"00000011",
  8373=>"00000000",
  8374=>"11111110",
  8375=>"11111110",
  8376=>"00000000",
  8377=>"00000001",
  8378=>"11111110",
  8379=>"11111110",
  8380=>"00000001",
  8381=>"00000000",
  8382=>"11111111",
  8383=>"11111111",
  8384=>"11111110",
  8385=>"11111111",
  8386=>"00000010",
  8387=>"00000010",
  8388=>"11111101",
  8389=>"00000010",
  8390=>"00000011",
  8391=>"00000001",
  8392=>"11111101",
  8393=>"00000000",
  8394=>"00000000",
  8395=>"00000000",
  8396=>"11111100",
  8397=>"11111100",
  8398=>"00000011",
  8399=>"11111110",
  8400=>"11111110",
  8401=>"00000001",
  8402=>"00000001",
  8403=>"11111101",
  8404=>"00000000",
  8405=>"11111111",
  8406=>"11111111",
  8407=>"00000000",
  8408=>"11111110",
  8409=>"00000000",
  8410=>"00000010",
  8411=>"00000001",
  8412=>"11111111",
  8413=>"11111111",
  8414=>"11111100",
  8415=>"11111111",
  8416=>"00000010",
  8417=>"11111101",
  8418=>"11111111",
  8419=>"00000010",
  8420=>"00000001",
  8421=>"11111101",
  8422=>"00000001",
  8423=>"00000011",
  8424=>"00000010",
  8425=>"00000011",
  8426=>"11111111",
  8427=>"00000010",
  8428=>"11111101",
  8429=>"11111101",
  8430=>"11111011",
  8431=>"11111110",
  8432=>"11111100",
  8433=>"11111111",
  8434=>"00000000",
  8435=>"00000000",
  8436=>"00000000",
  8437=>"00000011",
  8438=>"11111110",
  8439=>"00000001",
  8440=>"11111111",
  8441=>"11111101",
  8442=>"00000001",
  8443=>"00000000",
  8444=>"00000000",
  8445=>"11111111",
  8446=>"11111110",
  8447=>"11111110",
  8448=>"00000001",
  8449=>"11111110",
  8450=>"11111101",
  8451=>"11111111",
  8452=>"00000000",
  8453=>"00000000",
  8454=>"11111100",
  8455=>"11111101",
  8456=>"00000100",
  8457=>"11111111",
  8458=>"11111011",
  8459=>"00000000",
  8460=>"00000010",
  8461=>"11111100",
  8462=>"00000100",
  8463=>"00000001",
  8464=>"11111111",
  8465=>"11111110",
  8466=>"00000101",
  8467=>"00000011",
  8468=>"11111101",
  8469=>"11111101",
  8470=>"00000001",
  8471=>"00000000",
  8472=>"11111111",
  8473=>"11111101",
  8474=>"11111101",
  8475=>"00000001",
  8476=>"11111110",
  8477=>"11111101",
  8478=>"00000010",
  8479=>"11111110",
  8480=>"00000010",
  8481=>"00000011",
  8482=>"00000001",
  8483=>"11111111",
  8484=>"11111110",
  8485=>"11111110",
  8486=>"11111110",
  8487=>"11111100",
  8488=>"00000101",
  8489=>"11111111",
  8490=>"00000010",
  8491=>"00000001",
  8492=>"00000000",
  8493=>"00000000",
  8494=>"11111100",
  8495=>"00000000",
  8496=>"11111100",
  8497=>"11111101",
  8498=>"00000001",
  8499=>"11111110",
  8500=>"11111110",
  8501=>"11111110",
  8502=>"00000001",
  8503=>"11111110",
  8504=>"11111100",
  8505=>"00000010",
  8506=>"00000100",
  8507=>"00000010",
  8508=>"00000010",
  8509=>"00000001",
  8510=>"11111101",
  8511=>"00000001",
  8512=>"11111110",
  8513=>"00000000",
  8514=>"00000000",
  8515=>"00000011",
  8516=>"00000010",
  8517=>"00000001",
  8518=>"00000010",
  8519=>"00000000",
  8520=>"11111101",
  8521=>"11111111",
  8522=>"00000011",
  8523=>"11111111",
  8524=>"11111110",
  8525=>"00000101",
  8526=>"00000011",
  8527=>"11111110",
  8528=>"11111100",
  8529=>"00000001",
  8530=>"11111101",
  8531=>"11111110",
  8532=>"00000011",
  8533=>"00000011",
  8534=>"00000000",
  8535=>"11111101",
  8536=>"00000011",
  8537=>"11111111",
  8538=>"11111101",
  8539=>"11111111",
  8540=>"11111110",
  8541=>"11111110",
  8542=>"00000000",
  8543=>"00000000",
  8544=>"00000000",
  8545=>"00000001",
  8546=>"00000101",
  8547=>"11111111",
  8548=>"00000010",
  8549=>"00000001",
  8550=>"00000010",
  8551=>"00000000",
  8552=>"11111100",
  8553=>"00000011",
  8554=>"11111100",
  8555=>"11111110",
  8556=>"00000001",
  8557=>"11111110",
  8558=>"11111110",
  8559=>"00000010",
  8560=>"00000001",
  8561=>"00000011",
  8562=>"00000101",
  8563=>"11111111",
  8564=>"00000000",
  8565=>"11111111",
  8566=>"00000000",
  8567=>"11111111",
  8568=>"11111100",
  8569=>"00000010",
  8570=>"11111111",
  8571=>"11111100",
  8572=>"00000001",
  8573=>"11111111",
  8574=>"00000000",
  8575=>"00000000",
  8576=>"11111110",
  8577=>"11111111",
  8578=>"00000010",
  8579=>"00000101",
  8580=>"11111101",
  8581=>"11111111",
  8582=>"00000001",
  8583=>"11111110",
  8584=>"11111101",
  8585=>"00000100",
  8586=>"00000011",
  8587=>"00000011",
  8588=>"00000010",
  8589=>"00000100",
  8590=>"00000010",
  8591=>"11111110",
  8592=>"00000010",
  8593=>"11111111",
  8594=>"00000010",
  8595=>"00000000",
  8596=>"11111111",
  8597=>"11111111",
  8598=>"00000010",
  8599=>"11111110",
  8600=>"00000001",
  8601=>"11111101",
  8602=>"11111101",
  8603=>"00000001",
  8604=>"11111110",
  8605=>"00000000",
  8606=>"00000100",
  8607=>"00000000",
  8608=>"11111101",
  8609=>"11111111",
  8610=>"11111111",
  8611=>"11111101",
  8612=>"00000010",
  8613=>"11111011",
  8614=>"11111111",
  8615=>"11111101",
  8616=>"00000000",
  8617=>"00000011",
  8618=>"00000010",
  8619=>"11111110",
  8620=>"00000110",
  8621=>"00000010",
  8622=>"00000001",
  8623=>"00000000",
  8624=>"11111101",
  8625=>"00000010",
  8626=>"11111101",
  8627=>"11111101",
  8628=>"00000010",
  8629=>"11111100",
  8630=>"11111111",
  8631=>"00000001",
  8632=>"11111110",
  8633=>"11111111",
  8634=>"00000001",
  8635=>"11111110",
  8636=>"11111101",
  8637=>"00000000",
  8638=>"00000101",
  8639=>"11111101",
  8640=>"00000110",
  8641=>"11111110",
  8642=>"11111110",
  8643=>"00000101",
  8644=>"11111110",
  8645=>"11111111",
  8646=>"11111100",
  8647=>"11111100",
  8648=>"00000000",
  8649=>"00000100",
  8650=>"11111110",
  8651=>"11111111",
  8652=>"00000000",
  8653=>"11111110",
  8654=>"00000001",
  8655=>"00000010",
  8656=>"00000001",
  8657=>"11111111",
  8658=>"00000001",
  8659=>"11111111",
  8660=>"11111110",
  8661=>"00000011",
  8662=>"11111110",
  8663=>"11111111",
  8664=>"11111110",
  8665=>"11111111",
  8666=>"00000001",
  8667=>"11111101",
  8668=>"11111101",
  8669=>"00000011",
  8670=>"11111111",
  8671=>"00000110",
  8672=>"11111110",
  8673=>"00000000",
  8674=>"00000100",
  8675=>"00000001",
  8676=>"11111110",
  8677=>"00000001",
  8678=>"00000001",
  8679=>"00000011",
  8680=>"00000010",
  8681=>"11111101",
  8682=>"11111111",
  8683=>"00000010",
  8684=>"11111110",
  8685=>"00000010",
  8686=>"00000110",
  8687=>"00000000",
  8688=>"11111110",
  8689=>"00000001",
  8690=>"11111110",
  8691=>"00000000",
  8692=>"00000000",
  8693=>"00000000",
  8694=>"00000010",
  8695=>"00000011",
  8696=>"11111110",
  8697=>"00000000",
  8698=>"00000100",
  8699=>"11111110",
  8700=>"11111110",
  8701=>"11111111",
  8702=>"11111110",
  8703=>"00000000",
  8704=>"00000010",
  8705=>"11111101",
  8706=>"11111100",
  8707=>"11111101",
  8708=>"00000111",
  8709=>"00000001",
  8710=>"11111100",
  8711=>"00000011",
  8712=>"00000010",
  8713=>"00000000",
  8714=>"11111111",
  8715=>"00000011",
  8716=>"11111101",
  8717=>"11111111",
  8718=>"00000001",
  8719=>"11111110",
  8720=>"00000011",
  8721=>"00000001",
  8722=>"00000001",
  8723=>"11111110",
  8724=>"11111110",
  8725=>"00000000",
  8726=>"11111110",
  8727=>"11111111",
  8728=>"11111100",
  8729=>"11111101",
  8730=>"00000001",
  8731=>"11111110",
  8732=>"00000001",
  8733=>"00000011",
  8734=>"00000010",
  8735=>"11111110",
  8736=>"00000001",
  8737=>"00000100",
  8738=>"11111101",
  8739=>"00000011",
  8740=>"00000000",
  8741=>"11111111",
  8742=>"00000001",
  8743=>"11111101",
  8744=>"00000100",
  8745=>"00000100",
  8746=>"11111011",
  8747=>"11111101",
  8748=>"11111101",
  8749=>"00000001",
  8750=>"00000000",
  8751=>"00000001",
  8752=>"00000000",
  8753=>"00000000",
  8754=>"00000000",
  8755=>"00000011",
  8756=>"00000101",
  8757=>"11111111",
  8758=>"11111101",
  8759=>"00000001",
  8760=>"00000001",
  8761=>"00000011",
  8762=>"11111101",
  8763=>"00000010",
  8764=>"00000010",
  8765=>"00000010",
  8766=>"00000100",
  8767=>"00000001",
  8768=>"00000010",
  8769=>"11111111",
  8770=>"00000010",
  8771=>"11111101",
  8772=>"00000010",
  8773=>"00000000",
  8774=>"11111110",
  8775=>"00000001",
  8776=>"11111111",
  8777=>"00000000",
  8778=>"00000001",
  8779=>"11111111",
  8780=>"11111101",
  8781=>"11111111",
  8782=>"11111111",
  8783=>"00000001",
  8784=>"00000000",
  8785=>"00000000",
  8786=>"11111111",
  8787=>"11111111",
  8788=>"00000001",
  8789=>"00000000",
  8790=>"11111101",
  8791=>"11111111",
  8792=>"00000000",
  8793=>"11111110",
  8794=>"11111110",
  8795=>"00000000",
  8796=>"11111101",
  8797=>"11111101",
  8798=>"11111111",
  8799=>"00000001",
  8800=>"11111110",
  8801=>"00000100",
  8802=>"00000011",
  8803=>"11111101",
  8804=>"11111110",
  8805=>"11111101",
  8806=>"00000001",
  8807=>"00000010",
  8808=>"00000000",
  8809=>"00000001",
  8810=>"11111100",
  8811=>"00000011",
  8812=>"00000100",
  8813=>"11111111",
  8814=>"11111110",
  8815=>"00000001",
  8816=>"00000101",
  8817=>"00000100",
  8818=>"00000011",
  8819=>"00000011",
  8820=>"00000000",
  8821=>"11111010",
  8822=>"11111101",
  8823=>"11111100",
  8824=>"11111110",
  8825=>"11111111",
  8826=>"00000011",
  8827=>"11111110",
  8828=>"11111111",
  8829=>"00000011",
  8830=>"11111101",
  8831=>"00000001",
  8832=>"00000101",
  8833=>"00000001",
  8834=>"00000001",
  8835=>"11111110",
  8836=>"11111101",
  8837=>"00000000",
  8838=>"00000100",
  8839=>"00000010",
  8840=>"11111100",
  8841=>"00000011",
  8842=>"11111101",
  8843=>"11111101",
  8844=>"11111111",
  8845=>"00000010",
  8846=>"00000001",
  8847=>"11111111",
  8848=>"11111111",
  8849=>"11111111",
  8850=>"11111101",
  8851=>"00000010",
  8852=>"00000001",
  8853=>"11111111",
  8854=>"00000011",
  8855=>"00000100",
  8856=>"00000010",
  8857=>"00000001",
  8858=>"11111101",
  8859=>"00000100",
  8860=>"00000001",
  8861=>"11111100",
  8862=>"00000010",
  8863=>"00000000",
  8864=>"00000010",
  8865=>"00000000",
  8866=>"00000100",
  8867=>"00000100",
  8868=>"11111101",
  8869=>"00000101",
  8870=>"00000001",
  8871=>"11111111",
  8872=>"00000010",
  8873=>"00000011",
  8874=>"11111111",
  8875=>"00000010",
  8876=>"00000000",
  8877=>"00000010",
  8878=>"11111110",
  8879=>"00000100",
  8880=>"11111111",
  8881=>"11111111",
  8882=>"00000001",
  8883=>"00000100",
  8884=>"00000011",
  8885=>"00000011",
  8886=>"00000001",
  8887=>"11111110",
  8888=>"11111110",
  8889=>"00000000",
  8890=>"11111111",
  8891=>"11111101",
  8892=>"00000001",
  8893=>"11111101",
  8894=>"11111111",
  8895=>"00000000",
  8896=>"00000000",
  8897=>"11111111",
  8898=>"11111111",
  8899=>"00000000",
  8900=>"11111100",
  8901=>"11111101",
  8902=>"00000100",
  8903=>"00000001",
  8904=>"00000011",
  8905=>"11111110",
  8906=>"00000101",
  8907=>"00000000",
  8908=>"11111110",
  8909=>"00000010",
  8910=>"11111111",
  8911=>"11111111",
  8912=>"11111111",
  8913=>"11111101",
  8914=>"00000000",
  8915=>"11111111",
  8916=>"00000001",
  8917=>"11111101",
  8918=>"11111111",
  8919=>"11111101",
  8920=>"00000011",
  8921=>"00000010",
  8922=>"11111110",
  8923=>"00000001",
  8924=>"00000100",
  8925=>"00000010",
  8926=>"11111100",
  8927=>"11111111",
  8928=>"11111100",
  8929=>"00000001",
  8930=>"11111111",
  8931=>"11111110",
  8932=>"11111111",
  8933=>"11111110",
  8934=>"00000011",
  8935=>"00000000",
  8936=>"11111110",
  8937=>"00000011",
  8938=>"11111110",
  8939=>"11111111",
  8940=>"00000010",
  8941=>"00000000",
  8942=>"11111110",
  8943=>"11111101",
  8944=>"11111110",
  8945=>"00000001",
  8946=>"11111110",
  8947=>"11111101",
  8948=>"11111101",
  8949=>"00000000",
  8950=>"11111110",
  8951=>"11111100",
  8952=>"11111111",
  8953=>"11111110",
  8954=>"00000000",
  8955=>"11111110",
  8956=>"00000101",
  8957=>"00000101",
  8958=>"00000001",
  8959=>"11111101",
  8960=>"11111110",
  8961=>"11111101",
  8962=>"11111111",
  8963=>"11111101",
  8964=>"00000000",
  8965=>"11111110",
  8966=>"00000110",
  8967=>"11111111",
  8968=>"00000101",
  8969=>"11111101",
  8970=>"11111100",
  8971=>"00000001",
  8972=>"00000000",
  8973=>"11111110",
  8974=>"00000011",
  8975=>"00000001",
  8976=>"00000010",
  8977=>"00000010",
  8978=>"00000011",
  8979=>"11111101",
  8980=>"00000000",
  8981=>"11111110",
  8982=>"11111100",
  8983=>"11111100",
  8984=>"00000001",
  8985=>"00000000",
  8986=>"11111111",
  8987=>"11111111",
  8988=>"00000000",
  8989=>"11111111",
  8990=>"11111111",
  8991=>"11111100",
  8992=>"11111110",
  8993=>"00000000",
  8994=>"11111111",
  8995=>"00000000",
  8996=>"00000001",
  8997=>"11111111",
  8998=>"11111011",
  8999=>"00000011",
  9000=>"11111110",
  9001=>"11111110",
  9002=>"00000001",
  9003=>"00000011",
  9004=>"00000000",
  9005=>"00000000",
  9006=>"00000000",
  9007=>"11111111",
  9008=>"11111101",
  9009=>"00000000",
  9010=>"11111110",
  9011=>"00000010",
  9012=>"00000000",
  9013=>"11111111",
  9014=>"11111110",
  9015=>"00000011",
  9016=>"11111110",
  9017=>"00000010",
  9018=>"11111111",
  9019=>"00000001",
  9020=>"00000101",
  9021=>"00000010",
  9022=>"00000100",
  9023=>"11111111",
  9024=>"00000000",
  9025=>"00000000",
  9026=>"00000100",
  9027=>"11111111",
  9028=>"11111110",
  9029=>"00000100",
  9030=>"11111111",
  9031=>"00000010",
  9032=>"11111100",
  9033=>"00000110",
  9034=>"00000000",
  9035=>"00000001",
  9036=>"11111110",
  9037=>"00000001",
  9038=>"00000011",
  9039=>"00000000",
  9040=>"11111110",
  9041=>"11111111",
  9042=>"11111111",
  9043=>"00000000",
  9044=>"11111111",
  9045=>"11111111",
  9046=>"00000000",
  9047=>"00000000",
  9048=>"11111101",
  9049=>"00000101",
  9050=>"00000000",
  9051=>"11111100",
  9052=>"00000000",
  9053=>"11111100",
  9054=>"11111111",
  9055=>"11111110",
  9056=>"11111111",
  9057=>"11111110",
  9058=>"00000000",
  9059=>"00000001",
  9060=>"00000000",
  9061=>"00000010",
  9062=>"00000001",
  9063=>"11111110",
  9064=>"00000011",
  9065=>"00000011",
  9066=>"00000011",
  9067=>"11111101",
  9068=>"00000001",
  9069=>"00000000",
  9070=>"00000001",
  9071=>"00000001",
  9072=>"00000001",
  9073=>"11111110",
  9074=>"00000000",
  9075=>"11111110",
  9076=>"00000001",
  9077=>"00000010",
  9078=>"11111110",
  9079=>"00000101",
  9080=>"00000101",
  9081=>"00000000",
  9082=>"00000010",
  9083=>"11111111",
  9084=>"00000011",
  9085=>"11111110",
  9086=>"11111111",
  9087=>"11111101",
  9088=>"00000000",
  9089=>"11111101",
  9090=>"00000010",
  9091=>"00000010",
  9092=>"00000100",
  9093=>"11111110",
  9094=>"11111100",
  9095=>"00000001",
  9096=>"00000100",
  9097=>"00000110",
  9098=>"00000001",
  9099=>"11111111",
  9100=>"00000010",
  9101=>"11111111",
  9102=>"11111101",
  9103=>"11111110",
  9104=>"00000000",
  9105=>"00000000",
  9106=>"00000001",
  9107=>"11111110",
  9108=>"11111110",
  9109=>"00000001",
  9110=>"11111111",
  9111=>"11111101",
  9112=>"11111110",
  9113=>"11111110",
  9114=>"00000000",
  9115=>"11111101",
  9116=>"00000000",
  9117=>"11111111",
  9118=>"11111110",
  9119=>"11111100",
  9120=>"11111110",
  9121=>"00000101",
  9122=>"00000010",
  9123=>"11111110",
  9124=>"11111101",
  9125=>"00000100",
  9126=>"00000001",
  9127=>"11111011",
  9128=>"00000011",
  9129=>"00000001",
  9130=>"00000000",
  9131=>"11111111",
  9132=>"00000000",
  9133=>"00000001",
  9134=>"00000010",
  9135=>"11111101",
  9136=>"11111111",
  9137=>"11111111",
  9138=>"11111111",
  9139=>"00000001",
  9140=>"11111111",
  9141=>"00000011",
  9142=>"00000010",
  9143=>"00000000",
  9144=>"11111101",
  9145=>"00000000",
  9146=>"00000000",
  9147=>"00000010",
  9148=>"00000101",
  9149=>"00000001",
  9150=>"00000010",
  9151=>"11111101",
  9152=>"00000001",
  9153=>"00000000",
  9154=>"11111111",
  9155=>"00000010",
  9156=>"11111111",
  9157=>"00000100",
  9158=>"00000010",
  9159=>"11111111",
  9160=>"11111111",
  9161=>"11111111",
  9162=>"11111101",
  9163=>"00000011",
  9164=>"11111011",
  9165=>"00000001",
  9166=>"11111100",
  9167=>"11111101",
  9168=>"00000000",
  9169=>"00000010",
  9170=>"00000010",
  9171=>"00000011",
  9172=>"00000001",
  9173=>"11111111",
  9174=>"11111110",
  9175=>"00000011",
  9176=>"11111110",
  9177=>"00000010",
  9178=>"11111111",
  9179=>"00000110",
  9180=>"00000000",
  9181=>"00000100",
  9182=>"11111101",
  9183=>"11111110",
  9184=>"00000000",
  9185=>"11111100",
  9186=>"11111101",
  9187=>"00000010",
  9188=>"11111100",
  9189=>"11111100",
  9190=>"11111101",
  9191=>"00000010",
  9192=>"00000001",
  9193=>"00000001",
  9194=>"11111100",
  9195=>"11111111",
  9196=>"00000011",
  9197=>"11111111",
  9198=>"00000010",
  9199=>"00000001",
  9200=>"11111100",
  9201=>"11111110",
  9202=>"11111110",
  9203=>"00000011",
  9204=>"00000010",
  9205=>"00000001",
  9206=>"11111111",
  9207=>"00000001",
  9208=>"00000001",
  9209=>"00000010",
  9210=>"00000010",
  9211=>"11111100",
  9212=>"00000100",
  9213=>"00000011",
  9214=>"00000010",
  9215=>"11111110",
  9216=>"11111101",
  9217=>"00000101",
  9218=>"11111101",
  9219=>"11111110",
  9220=>"00000010",
  9221=>"11111100",
  9222=>"11111111",
  9223=>"00000101",
  9224=>"00000100",
  9225=>"00000010",
  9226=>"11111110",
  9227=>"00000001",
  9228=>"11111111",
  9229=>"00000110",
  9230=>"00000000",
  9231=>"11111111",
  9232=>"11111110",
  9233=>"00000001",
  9234=>"11111110",
  9235=>"00000100",
  9236=>"00000000",
  9237=>"00000001",
  9238=>"00000001",
  9239=>"00000011",
  9240=>"00000010",
  9241=>"00000101",
  9242=>"11111011",
  9243=>"00000000",
  9244=>"00000001",
  9245=>"00000000",
  9246=>"00000011",
  9247=>"00000011",
  9248=>"11111100",
  9249=>"00000100",
  9250=>"00000100",
  9251=>"00000011",
  9252=>"00000011",
  9253=>"00000000",
  9254=>"00000010",
  9255=>"00000010",
  9256=>"11111101",
  9257=>"11111101",
  9258=>"00000000",
  9259=>"11111110",
  9260=>"00000101",
  9261=>"00000001",
  9262=>"00000010",
  9263=>"11111101",
  9264=>"00000000",
  9265=>"00000100",
  9266=>"11111101",
  9267=>"00000100",
  9268=>"00000000",
  9269=>"00000100",
  9270=>"00000000",
  9271=>"11111100",
  9272=>"00000010",
  9273=>"00000010",
  9274=>"00000000",
  9275=>"00000010",
  9276=>"11111111",
  9277=>"11111100",
  9278=>"11111101",
  9279=>"11111111",
  9280=>"11111101",
  9281=>"00000010",
  9282=>"11111101",
  9283=>"00000100",
  9284=>"11111100",
  9285=>"00000011",
  9286=>"00000110",
  9287=>"00000000",
  9288=>"00000010",
  9289=>"11111110",
  9290=>"00000000",
  9291=>"00000010",
  9292=>"11111100",
  9293=>"11111110",
  9294=>"00000010",
  9295=>"00000000",
  9296=>"11111100",
  9297=>"00000101",
  9298=>"11111101",
  9299=>"00000100",
  9300=>"00000010",
  9301=>"00000011",
  9302=>"00000011",
  9303=>"00000001",
  9304=>"00000001",
  9305=>"00000100",
  9306=>"00000110",
  9307=>"00000111",
  9308=>"00000100",
  9309=>"11111100",
  9310=>"11111100",
  9311=>"00000011",
  9312=>"00000010",
  9313=>"11111100",
  9314=>"00000010",
  9315=>"11111101",
  9316=>"00000000",
  9317=>"00000000",
  9318=>"11111110",
  9319=>"00000010",
  9320=>"00000001",
  9321=>"11111010",
  9322=>"11111111",
  9323=>"00000011",
  9324=>"00000001",
  9325=>"00000000",
  9326=>"11111111",
  9327=>"11111111",
  9328=>"11111101",
  9329=>"00000001",
  9330=>"11111110",
  9331=>"11111101",
  9332=>"11111111",
  9333=>"00000000",
  9334=>"00000000",
  9335=>"11111010",
  9336=>"00000011",
  9337=>"00000011",
  9338=>"00000000",
  9339=>"11111110",
  9340=>"00000010",
  9341=>"00000011",
  9342=>"11111110",
  9343=>"00000001",
  9344=>"00000010",
  9345=>"11111100",
  9346=>"00000001",
  9347=>"11111111",
  9348=>"11111111",
  9349=>"00000101",
  9350=>"11111100",
  9351=>"00000001",
  9352=>"00000110",
  9353=>"11111110",
  9354=>"11111101",
  9355=>"11111111",
  9356=>"00000001",
  9357=>"00000000",
  9358=>"00000100",
  9359=>"00000010",
  9360=>"11111111",
  9361=>"00000001",
  9362=>"00000000",
  9363=>"00000000",
  9364=>"00000100",
  9365=>"11111111",
  9366=>"00000011",
  9367=>"00000001",
  9368=>"00000100",
  9369=>"11111111",
  9370=>"11111101",
  9371=>"00000010",
  9372=>"11111101",
  9373=>"00000001",
  9374=>"11111111",
  9375=>"00000011",
  9376=>"11111111",
  9377=>"00000010",
  9378=>"11111111",
  9379=>"11111101",
  9380=>"00000001",
  9381=>"11111110",
  9382=>"00000000",
  9383=>"00000011",
  9384=>"00000010",
  9385=>"00000010",
  9386=>"00000000",
  9387=>"11111011",
  9388=>"11111100",
  9389=>"11111010",
  9390=>"00000010",
  9391=>"11111101",
  9392=>"11111111",
  9393=>"11111101",
  9394=>"00000011",
  9395=>"11111100",
  9396=>"00000001",
  9397=>"11111110",
  9398=>"00000010",
  9399=>"11111111",
  9400=>"00000010",
  9401=>"00000110",
  9402=>"11111110",
  9403=>"00000011",
  9404=>"00000001",
  9405=>"11111111",
  9406=>"00000010",
  9407=>"00000110",
  9408=>"11111110",
  9409=>"00000100",
  9410=>"11111110",
  9411=>"00000101",
  9412=>"11111110",
  9413=>"11111111",
  9414=>"11111111",
  9415=>"00000100",
  9416=>"11111110",
  9417=>"00000100",
  9418=>"00000100",
  9419=>"11111111",
  9420=>"00000101",
  9421=>"11111111",
  9422=>"11111110",
  9423=>"11111011",
  9424=>"00000011",
  9425=>"11111101",
  9426=>"11111101",
  9427=>"11111111",
  9428=>"11111111",
  9429=>"00000110",
  9430=>"00000011",
  9431=>"11111111",
  9432=>"00000011",
  9433=>"00001001",
  9434=>"00000010",
  9435=>"11111100",
  9436=>"11111111",
  9437=>"11111110",
  9438=>"11111110",
  9439=>"11111110",
  9440=>"11111111",
  9441=>"00000000",
  9442=>"11111101",
  9443=>"00000001",
  9444=>"00000101",
  9445=>"00000011",
  9446=>"00000001",
  9447=>"11111100",
  9448=>"11111111",
  9449=>"11111111",
  9450=>"11111110",
  9451=>"11111110",
  9452=>"11111100",
  9453=>"00000001",
  9454=>"11111110",
  9455=>"00000010",
  9456=>"00000101",
  9457=>"00000001",
  9458=>"11111111",
  9459=>"11111101",
  9460=>"11111110",
  9461=>"11111101",
  9462=>"00000010",
  9463=>"11111111",
  9464=>"11111101",
  9465=>"11111111",
  9466=>"11111111",
  9467=>"11111110",
  9468=>"00000001",
  9469=>"00000010",
  9470=>"00000100",
  9471=>"11111101",
  9472=>"11111111",
  9473=>"00000100",
  9474=>"00000001",
  9475=>"11111101",
  9476=>"00000010",
  9477=>"11111111",
  9478=>"11111111",
  9479=>"11111101",
  9480=>"00000001",
  9481=>"00000010",
  9482=>"11111101",
  9483=>"00000011",
  9484=>"11111110",
  9485=>"00000000",
  9486=>"00000000",
  9487=>"00000011",
  9488=>"00000111",
  9489=>"00000001",
  9490=>"11111101",
  9491=>"11111110",
  9492=>"00000101",
  9493=>"00000010",
  9494=>"11111110",
  9495=>"00000011",
  9496=>"11111101",
  9497=>"11111100",
  9498=>"11111110",
  9499=>"00000011",
  9500=>"00000011",
  9501=>"11111101",
  9502=>"11111110",
  9503=>"11111110",
  9504=>"11111101",
  9505=>"00000011",
  9506=>"11111110",
  9507=>"00000010",
  9508=>"11111111",
  9509=>"00000011",
  9510=>"00000000",
  9511=>"00000100",
  9512=>"11111101",
  9513=>"00000111",
  9514=>"11111111",
  9515=>"11111110",
  9516=>"00000000",
  9517=>"00000011",
  9518=>"11111110",
  9519=>"11111110",
  9520=>"00000010",
  9521=>"00000001",
  9522=>"00000001",
  9523=>"00000010",
  9524=>"11111110",
  9525=>"00000101",
  9526=>"00000010",
  9527=>"00000000",
  9528=>"11111011",
  9529=>"00000011",
  9530=>"11111101",
  9531=>"00000101",
  9532=>"00000010",
  9533=>"11111110",
  9534=>"11111101",
  9535=>"00000011",
  9536=>"11111101",
  9537=>"00000001",
  9538=>"00000010",
  9539=>"11111110",
  9540=>"11111101",
  9541=>"11111111",
  9542=>"11111101",
  9543=>"00000001",
  9544=>"11111111",
  9545=>"00000000",
  9546=>"00000010",
  9547=>"00000010",
  9548=>"00000011",
  9549=>"11111101",
  9550=>"11111100",
  9551=>"00000000",
  9552=>"00000010",
  9553=>"00000000",
  9554=>"00000101",
  9555=>"11111101",
  9556=>"00000000",
  9557=>"00000000",
  9558=>"11111111",
  9559=>"00000001",
  9560=>"11111111",
  9561=>"00000010",
  9562=>"00000011",
  9563=>"11111101",
  9564=>"11111111",
  9565=>"00000010",
  9566=>"11111111",
  9567=>"00000000",
  9568=>"11111110",
  9569=>"00000100",
  9570=>"00000011",
  9571=>"00000010",
  9572=>"11111110",
  9573=>"11111110",
  9574=>"00000100",
  9575=>"00000001",
  9576=>"00000010",
  9577=>"00000001",
  9578=>"00000000",
  9579=>"11111111",
  9580=>"11111110",
  9581=>"00000001",
  9582=>"00000111",
  9583=>"00000011",
  9584=>"11111110",
  9585=>"00000100",
  9586=>"11111100",
  9587=>"00000010",
  9588=>"00000001",
  9589=>"00000001",
  9590=>"11111111",
  9591=>"00000010",
  9592=>"11111110",
  9593=>"00000011",
  9594=>"11111101",
  9595=>"00000010",
  9596=>"00000001",
  9597=>"11111111",
  9598=>"11111110",
  9599=>"11111110",
  9600=>"11111110",
  9601=>"00000011",
  9602=>"00000000",
  9603=>"11111110",
  9604=>"11111101",
  9605=>"00000011",
  9606=>"11111111",
  9607=>"11111101",
  9608=>"00000001",
  9609=>"00000010",
  9610=>"00000010",
  9611=>"00000001",
  9612=>"11111110",
  9613=>"11111111",
  9614=>"00000000",
  9615=>"00000000",
  9616=>"00000000",
  9617=>"11111110",
  9618=>"11111110",
  9619=>"00000101",
  9620=>"00000101",
  9621=>"00000000",
  9622=>"00000010",
  9623=>"11111110",
  9624=>"00000010",
  9625=>"00000001",
  9626=>"00000110",
  9627=>"11111011",
  9628=>"11111101",
  9629=>"00000011",
  9630=>"11111111",
  9631=>"00000000",
  9632=>"00000011",
  9633=>"00000111",
  9634=>"11111100",
  9635=>"11111110",
  9636=>"00000001",
  9637=>"11111100",
  9638=>"11111101",
  9639=>"00000101",
  9640=>"00000100",
  9641=>"00000000",
  9642=>"00000010",
  9643=>"00000001",
  9644=>"11111101",
  9645=>"00000000",
  9646=>"00000000",
  9647=>"00000001",
  9648=>"11111110",
  9649=>"00000011",
  9650=>"00000001",
  9651=>"11111110",
  9652=>"00000001",
  9653=>"11111111",
  9654=>"00000000",
  9655=>"00000101",
  9656=>"11111110",
  9657=>"00000000",
  9658=>"11111101",
  9659=>"00000100",
  9660=>"11111110",
  9661=>"11111111",
  9662=>"11111100",
  9663=>"11111101",
  9664=>"11111101",
  9665=>"11111101",
  9666=>"11111110",
  9667=>"00000011",
  9668=>"00000000",
  9669=>"00000000",
  9670=>"11111110",
  9671=>"11111110",
  9672=>"00000100",
  9673=>"11111110",
  9674=>"00000000",
  9675=>"11111110",
  9676=>"00000010",
  9677=>"00000000",
  9678=>"00000001",
  9679=>"11111100",
  9680=>"11111110",
  9681=>"11111111",
  9682=>"11111101",
  9683=>"00000001",
  9684=>"00000110",
  9685=>"00000000",
  9686=>"00000000",
  9687=>"00000000",
  9688=>"00000010",
  9689=>"00000011",
  9690=>"00000100",
  9691=>"11111110",
  9692=>"11111110",
  9693=>"11111110",
  9694=>"00000000",
  9695=>"00000000",
  9696=>"11111101",
  9697=>"11111111",
  9698=>"11111111",
  9699=>"00000010",
  9700=>"11111101",
  9701=>"00000011",
  9702=>"11111101",
  9703=>"11111101",
  9704=>"00000111",
  9705=>"00000011",
  9706=>"11111101",
  9707=>"00000010",
  9708=>"11111110",
  9709=>"11111011",
  9710=>"00000011",
  9711=>"11111111",
  9712=>"00000000",
  9713=>"00000110",
  9714=>"11111111",
  9715=>"11111110",
  9716=>"00000010",
  9717=>"00000101",
  9718=>"00000001",
  9719=>"00000001",
  9720=>"00000001",
  9721=>"00000001",
  9722=>"00000010",
  9723=>"00000011",
  9724=>"00000001",
  9725=>"11111100",
  9726=>"11111110",
  9727=>"11111100",
  9728=>"00000011",
  9729=>"11111111",
  9730=>"00000100",
  9731=>"00000101",
  9732=>"11111101",
  9733=>"00000011",
  9734=>"00000011",
  9735=>"11111101",
  9736=>"11111111",
  9737=>"11111101",
  9738=>"00000010",
  9739=>"00000000",
  9740=>"11111100",
  9741=>"00000001",
  9742=>"11111011",
  9743=>"00000000",
  9744=>"00000001",
  9745=>"11111100",
  9746=>"00000011",
  9747=>"11111110",
  9748=>"00000111",
  9749=>"00000000",
  9750=>"00000001",
  9751=>"00000000",
  9752=>"11111011",
  9753=>"00000001",
  9754=>"11111101",
  9755=>"00000010",
  9756=>"00000000",
  9757=>"11111100",
  9758=>"00000011",
  9759=>"11111101",
  9760=>"00000010",
  9761=>"00000000",
  9762=>"11111110",
  9763=>"00000001",
  9764=>"00000000",
  9765=>"11111101",
  9766=>"00000010",
  9767=>"00000011",
  9768=>"11111101",
  9769=>"00000000",
  9770=>"11111110",
  9771=>"00000000",
  9772=>"11111101",
  9773=>"00000001",
  9774=>"00000100",
  9775=>"00000110",
  9776=>"00000010",
  9777=>"00000000",
  9778=>"11111101",
  9779=>"00000010",
  9780=>"11111101",
  9781=>"00000011",
  9782=>"11111011",
  9783=>"00000000",
  9784=>"11111101",
  9785=>"11111111",
  9786=>"11111101",
  9787=>"00000011",
  9788=>"00000001",
  9789=>"00000101",
  9790=>"11111110",
  9791=>"11111110",
  9792=>"00000001",
  9793=>"00000000",
  9794=>"00000011",
  9795=>"00000110",
  9796=>"00000000",
  9797=>"00000010",
  9798=>"00000100",
  9799=>"00000000",
  9800=>"11111101",
  9801=>"00000001",
  9802=>"00000100",
  9803=>"11111111",
  9804=>"11111110",
  9805=>"00000001",
  9806=>"11111110",
  9807=>"00000010",
  9808=>"11111111",
  9809=>"11111101",
  9810=>"11111111",
  9811=>"00000001",
  9812=>"11111101",
  9813=>"00000000",
  9814=>"00000001",
  9815=>"11111111",
  9816=>"00000101",
  9817=>"00000011",
  9818=>"11111110",
  9819=>"11111111",
  9820=>"00000010",
  9821=>"11111111",
  9822=>"00000000",
  9823=>"00000000",
  9824=>"00000001",
  9825=>"00000000",
  9826=>"11111111",
  9827=>"11111110",
  9828=>"00000100",
  9829=>"00000000",
  9830=>"00000100",
  9831=>"00000011",
  9832=>"00000010",
  9833=>"00000010",
  9834=>"11111110",
  9835=>"00000010",
  9836=>"00000010",
  9837=>"11111110",
  9838=>"00000001",
  9839=>"00000010",
  9840=>"00000000",
  9841=>"11111100",
  9842=>"11111110",
  9843=>"00000010",
  9844=>"00000001",
  9845=>"11111101",
  9846=>"00000101",
  9847=>"00000001",
  9848=>"11111110",
  9849=>"11111101",
  9850=>"00000011",
  9851=>"11111100",
  9852=>"11111110",
  9853=>"00000010",
  9854=>"00000010",
  9855=>"11111100",
  9856=>"00000001",
  9857=>"00000010",
  9858=>"00000000",
  9859=>"00000001",
  9860=>"00000101",
  9861=>"00000000",
  9862=>"11111111",
  9863=>"11111111",
  9864=>"11111011",
  9865=>"00000000",
  9866=>"11111101",
  9867=>"00000011",
  9868=>"00000010",
  9869=>"00000100",
  9870=>"11111110",
  9871=>"11111111",
  9872=>"11111100",
  9873=>"00000011",
  9874=>"00000010",
  9875=>"00000010",
  9876=>"00000010",
  9877=>"00000001",
  9878=>"11111111",
  9879=>"00000110",
  9880=>"00000010",
  9881=>"11111100",
  9882=>"11111100",
  9883=>"11111101",
  9884=>"00000011",
  9885=>"11111111",
  9886=>"11111111",
  9887=>"00000001",
  9888=>"11111110",
  9889=>"00000011",
  9890=>"00000010",
  9891=>"11111111",
  9892=>"11111101",
  9893=>"11111111",
  9894=>"00000011",
  9895=>"11111110",
  9896=>"00000100",
  9897=>"11111101",
  9898=>"00000010",
  9899=>"00000010",
  9900=>"11111100",
  9901=>"11111100",
  9902=>"00000100",
  9903=>"11111110",
  9904=>"00000001",
  9905=>"00000011",
  9906=>"00000011",
  9907=>"00000001",
  9908=>"00000000",
  9909=>"11111101",
  9910=>"00000000",
  9911=>"11111110",
  9912=>"00000001",
  9913=>"00000000",
  9914=>"11111110",
  9915=>"11111100",
  9916=>"00000101",
  9917=>"11111111",
  9918=>"00000001",
  9919=>"11111110",
  9920=>"11111101",
  9921=>"00000000",
  9922=>"11111110",
  9923=>"11111011",
  9924=>"00000011",
  9925=>"00000000",
  9926=>"11111110",
  9927=>"00000010",
  9928=>"11111110",
  9929=>"11111011",
  9930=>"11111110",
  9931=>"11111111",
  9932=>"11111100",
  9933=>"11111110",
  9934=>"00000000",
  9935=>"00000100",
  9936=>"11111110",
  9937=>"11111111",
  9938=>"11111110",
  9939=>"11111111",
  9940=>"00000000",
  9941=>"00000100",
  9942=>"00000001",
  9943=>"00000100",
  9944=>"11111101",
  9945=>"00000010",
  9946=>"11111100",
  9947=>"11111101",
  9948=>"00000001",
  9949=>"00000000",
  9950=>"11111110",
  9951=>"00000011",
  9952=>"00000101",
  9953=>"00000001",
  9954=>"00000001",
  9955=>"00000010",
  9956=>"00000011",
  9957=>"11111100",
  9958=>"00000010",
  9959=>"00000100",
  9960=>"11111101",
  9961=>"11111111",
  9962=>"11111110",
  9963=>"11111110",
  9964=>"11111101",
  9965=>"00000000",
  9966=>"00000100",
  9967=>"11111110",
  9968=>"00000110",
  9969=>"00000011",
  9970=>"00000011",
  9971=>"11111111",
  9972=>"00000001",
  9973=>"00000010",
  9974=>"11111110",
  9975=>"00000010",
  9976=>"00000001",
  9977=>"00000000",
  9978=>"00000100",
  9979=>"00000101",
  9980=>"00000010",
  9981=>"11111011",
  9982=>"11111111",
  9983=>"00000100",
  9984=>"00000000",
  9985=>"11111110",
  9986=>"11111110",
  9987=>"11111101",
  9988=>"11111101",
  9989=>"00000010",
  9990=>"11111010",
  9991=>"00000000",
  9992=>"00000000",
  9993=>"11111100",
  9994=>"00000010",
  9995=>"00000011",
  9996=>"00000010",
  9997=>"11111101",
  9998=>"00000111",
  9999=>"11111111",
  10000=>"11111110",
  10001=>"00000011",
  10002=>"00000110",
  10003=>"00000011",
  10004=>"11111110",
  10005=>"11111111",
  10006=>"00000000",
  10007=>"00000100",
  10008=>"00000001",
  10009=>"00000000",
  10010=>"00000011",
  10011=>"11111111",
  10012=>"00000010",
  10013=>"11111101",
  10014=>"00000000",
  10015=>"11111100",
  10016=>"11111111",
  10017=>"00000010",
  10018=>"11111110",
  10019=>"00000001",
  10020=>"00000001",
  10021=>"00000000",
  10022=>"00000101",
  10023=>"11111111",
  10024=>"00000000",
  10025=>"00000000",
  10026=>"00000010",
  10027=>"11111011",
  10028=>"00000000",
  10029=>"00000001",
  10030=>"00000010",
  10031=>"00000100",
  10032=>"11111111",
  10033=>"11111111",
  10034=>"00000001",
  10035=>"00000100",
  10036=>"00000011",
  10037=>"11111110",
  10038=>"00000000",
  10039=>"00000000",
  10040=>"00000000",
  10041=>"11111100",
  10042=>"00000100",
  10043=>"00000011",
  10044=>"11111101",
  10045=>"11111110",
  10046=>"00000001",
  10047=>"11111110",
  10048=>"00000101",
  10049=>"11111101",
  10050=>"00000011",
  10051=>"00000001",
  10052=>"00000000",
  10053=>"00000010",
  10054=>"00000010",
  10055=>"00000010",
  10056=>"11111101",
  10057=>"00000001",
  10058=>"00000011",
  10059=>"00000001",
  10060=>"11111110",
  10061=>"00000000",
  10062=>"11111111",
  10063=>"00000010",
  10064=>"11111110",
  10065=>"11111111",
  10066=>"00000010",
  10067=>"00000011",
  10068=>"11111111",
  10069=>"11111100",
  10070=>"00000000",
  10071=>"00000011",
  10072=>"11111110",
  10073=>"11111101",
  10074=>"00000010",
  10075=>"11111110",
  10076=>"00000001",
  10077=>"00000000",
  10078=>"00000001",
  10079=>"00000000",
  10080=>"11111111",
  10081=>"00000000",
  10082=>"11111101",
  10083=>"00000010",
  10084=>"11111111",
  10085=>"00000010",
  10086=>"11111111",
  10087=>"11111111",
  10088=>"11111110",
  10089=>"11111111",
  10090=>"11111101",
  10091=>"00000001",
  10092=>"00000100",
  10093=>"00000001",
  10094=>"00000010",
  10095=>"00000101",
  10096=>"00000011",
  10097=>"00000000",
  10098=>"00000010",
  10099=>"00000100",
  10100=>"11111111",
  10101=>"11111100",
  10102=>"11111111",
  10103=>"11111110",
  10104=>"00000000",
  10105=>"00000001",
  10106=>"00000011",
  10107=>"11111100",
  10108=>"11111101",
  10109=>"11111101",
  10110=>"00000011",
  10111=>"00000000",
  10112=>"00000000",
  10113=>"00000101",
  10114=>"11111110",
  10115=>"00000110",
  10116=>"00000000",
  10117=>"00000011",
  10118=>"11111111",
  10119=>"00000100",
  10120=>"11111111",
  10121=>"11111111",
  10122=>"00000100",
  10123=>"11111110",
  10124=>"11111100",
  10125=>"00000001",
  10126=>"11111100",
  10127=>"00000100",
  10128=>"00000000",
  10129=>"00000101",
  10130=>"00000010",
  10131=>"11111101",
  10132=>"11111100",
  10133=>"11111100",
  10134=>"00000000",
  10135=>"00000000",
  10136=>"00000111",
  10137=>"11111100",
  10138=>"00000010",
  10139=>"00000011",
  10140=>"00000001",
  10141=>"11111110",
  10142=>"11111111",
  10143=>"11111110",
  10144=>"11111101",
  10145=>"11111111",
  10146=>"00000000",
  10147=>"00000001",
  10148=>"11111111",
  10149=>"00000000",
  10150=>"00000000",
  10151=>"11111110",
  10152=>"11111110",
  10153=>"00000000",
  10154=>"00000000",
  10155=>"11111111",
  10156=>"00000100",
  10157=>"00000000",
  10158=>"11111101",
  10159=>"00000010",
  10160=>"00000010",
  10161=>"00000011",
  10162=>"00000011",
  10163=>"00000100",
  10164=>"00000010",
  10165=>"00000000",
  10166=>"11111101",
  10167=>"00000100",
  10168=>"00000011",
  10169=>"00000001",
  10170=>"00000011",
  10171=>"11111110",
  10172=>"11111011",
  10173=>"11111101",
  10174=>"00000001",
  10175=>"11111101",
  10176=>"00000011",
  10177=>"00000011",
  10178=>"00000010",
  10179=>"11111111",
  10180=>"00000000",
  10181=>"11111111",
  10182=>"00000001",
  10183=>"00000001",
  10184=>"00000011",
  10185=>"11111110",
  10186=>"00000100",
  10187=>"00000010",
  10188=>"00000100",
  10189=>"11111011",
  10190=>"11111110",
  10191=>"11111111",
  10192=>"00000100",
  10193=>"11111100",
  10194=>"00000101",
  10195=>"00000011",
  10196=>"11111111",
  10197=>"00000100",
  10198=>"00000100",
  10199=>"11111101",
  10200=>"00000010",
  10201=>"00000001",
  10202=>"11111111",
  10203=>"00000001",
  10204=>"00000010",
  10205=>"00000101",
  10206=>"00000110",
  10207=>"00000101",
  10208=>"00000010",
  10209=>"00000001",
  10210=>"00000100",
  10211=>"11111111",
  10212=>"11111100",
  10213=>"00000001",
  10214=>"00000001",
  10215=>"00000101",
  10216=>"00000010",
  10217=>"00000011",
  10218=>"00000000",
  10219=>"00000100",
  10220=>"00000001",
  10221=>"00000011",
  10222=>"11111101",
  10223=>"00000001",
  10224=>"00000110",
  10225=>"00000010",
  10226=>"00000001",
  10227=>"11111111",
  10228=>"00000101",
  10229=>"00000000",
  10230=>"00000001",
  10231=>"00000100",
  10232=>"00000000",
  10233=>"00000010",
  10234=>"11111111",
  10235=>"11111101",
  10236=>"00000010",
  10237=>"00000000",
  10238=>"00000010",
  10239=>"00000010",
  10240=>"00000001",
  10241=>"00000001",
  10242=>"00000010",
  10243=>"11111100",
  10244=>"00000000",
  10245=>"00000010",
  10246=>"00000010",
  10247=>"11111110",
  10248=>"11111111",
  10249=>"11111111",
  10250=>"11111100",
  10251=>"11111110",
  10252=>"11111111",
  10253=>"11111101",
  10254=>"11111100",
  10255=>"11111111",
  10256=>"00000010",
  10257=>"00000100",
  10258=>"00000010",
  10259=>"00000100",
  10260=>"11111110",
  10261=>"00000000",
  10262=>"11111110",
  10263=>"11111111",
  10264=>"11111110",
  10265=>"00000001",
  10266=>"00000000",
  10267=>"11111110",
  10268=>"00000010",
  10269=>"11111111",
  10270=>"00000001",
  10271=>"00000001",
  10272=>"00000001",
  10273=>"00000001",
  10274=>"00000010",
  10275=>"00000001",
  10276=>"11111111",
  10277=>"00000100",
  10278=>"11111101",
  10279=>"11111100",
  10280=>"00000000",
  10281=>"11111110",
  10282=>"11111110",
  10283=>"11111101",
  10284=>"11111110",
  10285=>"11111111",
  10286=>"00000000",
  10287=>"11111110",
  10288=>"11111110",
  10289=>"00000000",
  10290=>"00000001",
  10291=>"00000000",
  10292=>"00000010",
  10293=>"11111110",
  10294=>"11111111",
  10295=>"11111110",
  10296=>"00000011",
  10297=>"00000010",
  10298=>"00000000",
  10299=>"00000010",
  10300=>"00000000",
  10301=>"00000001",
  10302=>"00000001",
  10303=>"00000011",
  10304=>"11111111",
  10305=>"11111110",
  10306=>"00000010",
  10307=>"11111100",
  10308=>"11111101",
  10309=>"11111101",
  10310=>"11111101",
  10311=>"00000100",
  10312=>"11111110",
  10313=>"11111110",
  10314=>"00000011",
  10315=>"00000000",
  10316=>"00000000",
  10317=>"00000000",
  10318=>"00000010",
  10319=>"00000001",
  10320=>"00000100",
  10321=>"00000001",
  10322=>"11111111",
  10323=>"00000000",
  10324=>"00000100",
  10325=>"00000000",
  10326=>"00000010",
  10327=>"00000001",
  10328=>"00000000",
  10329=>"11111111",
  10330=>"00000000",
  10331=>"11111101",
  10332=>"11111011",
  10333=>"11111110",
  10334=>"00000010",
  10335=>"11111111",
  10336=>"00000000",
  10337=>"00000010",
  10338=>"00000000",
  10339=>"00000100",
  10340=>"00000110",
  10341=>"00000000",
  10342=>"00000010",
  10343=>"11111110",
  10344=>"00000001",
  10345=>"00000010",
  10346=>"00000000",
  10347=>"11111111",
  10348=>"00000010",
  10349=>"11111110",
  10350=>"11111111",
  10351=>"00000001",
  10352=>"11111101",
  10353=>"00000010",
  10354=>"11111110",
  10355=>"11111111",
  10356=>"00000000",
  10357=>"11111110",
  10358=>"00000011",
  10359=>"00000100",
  10360=>"00000000",
  10361=>"11111111",
  10362=>"11111111",
  10363=>"00000000",
  10364=>"00000000",
  10365=>"00000011",
  10366=>"11111110",
  10367=>"11111110",
  10368=>"00000001",
  10369=>"00000010",
  10370=>"11111111",
  10371=>"00000000",
  10372=>"11111111",
  10373=>"11111110",
  10374=>"11111101",
  10375=>"11111110",
  10376=>"00000011",
  10377=>"00000001",
  10378=>"00000000",
  10379=>"00000001",
  10380=>"11111111",
  10381=>"11111101",
  10382=>"11111110",
  10383=>"11111111",
  10384=>"00000010",
  10385=>"00000000",
  10386=>"00000000",
  10387=>"11111111",
  10388=>"00000010",
  10389=>"00000001",
  10390=>"11111110",
  10391=>"00000000",
  10392=>"00000010",
  10393=>"11111110",
  10394=>"11111110",
  10395=>"00000001",
  10396=>"11111111",
  10397=>"00000100",
  10398=>"00000011",
  10399=>"11111111",
  10400=>"11111101",
  10401=>"11111101",
  10402=>"00000010",
  10403=>"11111111",
  10404=>"11111110",
  10405=>"11111101",
  10406=>"11111111",
  10407=>"00000010",
  10408=>"00000001",
  10409=>"11111100",
  10410=>"11111110",
  10411=>"11111100",
  10412=>"11111100",
  10413=>"00000001",
  10414=>"00000001",
  10415=>"00000010",
  10416=>"00000001",
  10417=>"11111110",
  10418=>"00000000",
  10419=>"00000000",
  10420=>"00000010",
  10421=>"00000000",
  10422=>"00000011",
  10423=>"00000000",
  10424=>"11111101",
  10425=>"11111101",
  10426=>"11111101",
  10427=>"11111111",
  10428=>"00000001",
  10429=>"00000010",
  10430=>"00000000",
  10431=>"00000101",
  10432=>"00000010",
  10433=>"00000000",
  10434=>"11111110",
  10435=>"11111110",
  10436=>"00000001",
  10437=>"00000001",
  10438=>"00000001",
  10439=>"11111111",
  10440=>"00000000",
  10441=>"11111101",
  10442=>"11111111",
  10443=>"00000011",
  10444=>"00000011",
  10445=>"11111101",
  10446=>"00000011",
  10447=>"00000000",
  10448=>"11111101",
  10449=>"11111101",
  10450=>"00000010",
  10451=>"00000001",
  10452=>"00000010",
  10453=>"00000001",
  10454=>"00000000",
  10455=>"11111100",
  10456=>"00000010",
  10457=>"00000000",
  10458=>"00000000",
  10459=>"00000100",
  10460=>"11111111",
  10461=>"11111110",
  10462=>"00000000",
  10463=>"11111111",
  10464=>"00000001",
  10465=>"00000001",
  10466=>"11111111",
  10467=>"11111111",
  10468=>"00000001",
  10469=>"11111110",
  10470=>"00000010",
  10471=>"00000000",
  10472=>"11111111",
  10473=>"11111110",
  10474=>"11111110",
  10475=>"11111111",
  10476=>"00000000",
  10477=>"11111101",
  10478=>"00000100",
  10479=>"00000001",
  10480=>"11111110",
  10481=>"00000000",
  10482=>"00000001",
  10483=>"11111111",
  10484=>"11111110",
  10485=>"11111110",
  10486=>"11111111",
  10487=>"11111111",
  10488=>"00000011",
  10489=>"00000011",
  10490=>"00000011",
  10491=>"11111110",
  10492=>"00000101",
  10493=>"11111111",
  10494=>"00000000",
  10495=>"00000000",
  10496=>"11111110",
  10497=>"00000011",
  10498=>"11111101",
  10499=>"00000100",
  10500=>"11111110",
  10501=>"00000100",
  10502=>"11111101",
  10503=>"00000000",
  10504=>"11111110",
  10505=>"00000000",
  10506=>"11111110",
  10507=>"00000000",
  10508=>"00000000",
  10509=>"11111100",
  10510=>"00000000",
  10511=>"11111100",
  10512=>"00000001",
  10513=>"11111110",
  10514=>"11111110",
  10515=>"11111101",
  10516=>"00000000",
  10517=>"00000001",
  10518=>"11111111",
  10519=>"11111110",
  10520=>"00000011",
  10521=>"11111110",
  10522=>"11111111",
  10523=>"00000000",
  10524=>"00000001",
  10525=>"00000011",
  10526=>"11111111",
  10527=>"11111101",
  10528=>"00000010",
  10529=>"11111111",
  10530=>"00000011",
  10531=>"11111101",
  10532=>"11111110",
  10533=>"00000010",
  10534=>"00000010",
  10535=>"00000000",
  10536=>"11111111",
  10537=>"00000100",
  10538=>"11111110",
  10539=>"00000100",
  10540=>"00000110",
  10541=>"00000001",
  10542=>"00000011",
  10543=>"00000010",
  10544=>"11111101",
  10545=>"11111111",
  10546=>"00000100",
  10547=>"00000000",
  10548=>"11111111",
  10549=>"11111110",
  10550=>"00000100",
  10551=>"11111101",
  10552=>"00000100",
  10553=>"11111111",
  10554=>"00000001",
  10555=>"00000000",
  10556=>"11111110",
  10557=>"11111101",
  10558=>"11111111",
  10559=>"11111110",
  10560=>"00000001",
  10561=>"11111110",
  10562=>"11111111",
  10563=>"00000001",
  10564=>"11111110",
  10565=>"11111110",
  10566=>"11111111",
  10567=>"00000000",
  10568=>"11111101",
  10569=>"00000001",
  10570=>"11111111",
  10571=>"11111101",
  10572=>"11111111",
  10573=>"00000010",
  10574=>"00000001",
  10575=>"00000000",
  10576=>"00000010",
  10577=>"00000001",
  10578=>"00000000",
  10579=>"11111111",
  10580=>"00000010",
  10581=>"11111110",
  10582=>"11111110",
  10583=>"00000001",
  10584=>"11111111",
  10585=>"11111101",
  10586=>"11111110",
  10587=>"00000010",
  10588=>"11111110",
  10589=>"11111111",
  10590=>"11111110",
  10591=>"00000000",
  10592=>"11111100",
  10593=>"11111111",
  10594=>"00000001",
  10595=>"11111110",
  10596=>"00000001",
  10597=>"11111110",
  10598=>"00000001",
  10599=>"00000001",
  10600=>"11111100",
  10601=>"11111110",
  10602=>"00000001",
  10603=>"00000000",
  10604=>"00000010",
  10605=>"00000001",
  10606=>"00000000",
  10607=>"00000010",
  10608=>"11111111",
  10609=>"00000011",
  10610=>"00000001",
  10611=>"11111101",
  10612=>"11111101",
  10613=>"11111101",
  10614=>"00000011",
  10615=>"00000001",
  10616=>"11111100",
  10617=>"11111100",
  10618=>"00000000",
  10619=>"11111101",
  10620=>"00000001",
  10621=>"00000000",
  10622=>"11111101",
  10623=>"00000010",
  10624=>"11111101",
  10625=>"00000000",
  10626=>"11111101",
  10627=>"00000010",
  10628=>"00000010",
  10629=>"00000010",
  10630=>"11111110",
  10631=>"00000011",
  10632=>"11111101",
  10633=>"11111110",
  10634=>"00000000",
  10635=>"00000010",
  10636=>"00000001",
  10637=>"11111110",
  10638=>"11111101",
  10639=>"00000010",
  10640=>"00000011",
  10641=>"11111101",
  10642=>"11111101",
  10643=>"00000010",
  10644=>"11111110",
  10645=>"11111101",
  10646=>"00000001",
  10647=>"11111110",
  10648=>"11111101",
  10649=>"11111101",
  10650=>"11111111",
  10651=>"00000101",
  10652=>"00000000",
  10653=>"11111111",
  10654=>"00000000",
  10655=>"00000010",
  10656=>"11111110",
  10657=>"00000100",
  10658=>"00000001",
  10659=>"11111110",
  10660=>"11111111",
  10661=>"11111100",
  10662=>"11111110",
  10663=>"00000000",
  10664=>"11111100",
  10665=>"00000001",
  10666=>"11111111",
  10667=>"00000011",
  10668=>"00000111",
  10669=>"00000100",
  10670=>"00000000",
  10671=>"00000001",
  10672=>"00000010",
  10673=>"00000011",
  10674=>"00000010",
  10675=>"11111110",
  10676=>"00000001",
  10677=>"11111110",
  10678=>"11111111",
  10679=>"00000001",
  10680=>"11111111",
  10681=>"00000010",
  10682=>"00000001",
  10683=>"11111111",
  10684=>"00000001",
  10685=>"11111111",
  10686=>"11111101",
  10687=>"00000001",
  10688=>"11111110",
  10689=>"00000100",
  10690=>"11111100",
  10691=>"00000011",
  10692=>"00000011",
  10693=>"11111111",
  10694=>"11111110",
  10695=>"11111101",
  10696=>"11111110",
  10697=>"00000001",
  10698=>"00000101",
  10699=>"11111110",
  10700=>"11111111",
  10701=>"00000000",
  10702=>"11111100",
  10703=>"00000000",
  10704=>"11111110",
  10705=>"00000001",
  10706=>"00000000",
  10707=>"11111101",
  10708=>"11111101",
  10709=>"00000100",
  10710=>"11111101",
  10711=>"00000001",
  10712=>"00000010",
  10713=>"00000001",
  10714=>"00000010",
  10715=>"11111110",
  10716=>"11111111",
  10717=>"11111110",
  10718=>"11111110",
  10719=>"00000000",
  10720=>"11111110",
  10721=>"11111101",
  10722=>"11111110",
  10723=>"11111110",
  10724=>"11111111",
  10725=>"00000010",
  10726=>"11111110",
  10727=>"00000001",
  10728=>"00000000",
  10729=>"00000010",
  10730=>"00000011",
  10731=>"11111101",
  10732=>"00000000",
  10733=>"00000100",
  10734=>"00000010",
  10735=>"00000001",
  10736=>"00000001",
  10737=>"11111110",
  10738=>"00000010",
  10739=>"00000010",
  10740=>"11111110",
  10741=>"11111111",
  10742=>"11111111",
  10743=>"11111100",
  10744=>"00000010",
  10745=>"11111110",
  10746=>"11111111",
  10747=>"11111110",
  10748=>"00000000",
  10749=>"00000001",
  10750=>"00000110",
  10751=>"00000001",
  10752=>"00000100",
  10753=>"11111110",
  10754=>"00000001",
  10755=>"00000000",
  10756=>"00001000",
  10757=>"00000010",
  10758=>"11111101",
  10759=>"00000000",
  10760=>"00000010",
  10761=>"11111100",
  10762=>"00000001",
  10763=>"11111111",
  10764=>"00000101",
  10765=>"11111111",
  10766=>"11111110",
  10767=>"00000000",
  10768=>"00000000",
  10769=>"11111111",
  10770=>"11111111",
  10771=>"00000001",
  10772=>"11111101",
  10773=>"00000010",
  10774=>"00000001",
  10775=>"11111110",
  10776=>"11111101",
  10777=>"11111110",
  10778=>"00000000",
  10779=>"00000001",
  10780=>"11111110",
  10781=>"11111110",
  10782=>"00000010",
  10783=>"11111100",
  10784=>"11111111",
  10785=>"00000000",
  10786=>"11111111",
  10787=>"00000010",
  10788=>"00000000",
  10789=>"00000010",
  10790=>"11111110",
  10791=>"11111111",
  10792=>"00000001",
  10793=>"00000011",
  10794=>"00000010",
  10795=>"00000000",
  10796=>"11111101",
  10797=>"11111101",
  10798=>"11111110",
  10799=>"00000010",
  10800=>"11111110",
  10801=>"00000000",
  10802=>"00000001",
  10803=>"00000000",
  10804=>"11111110",
  10805=>"00000000",
  10806=>"00000001",
  10807=>"00000011",
  10808=>"00000111",
  10809=>"11111110",
  10810=>"11111111",
  10811=>"11111100",
  10812=>"00000001",
  10813=>"11111101",
  10814=>"11111101",
  10815=>"11111110",
  10816=>"00000001",
  10817=>"11111111",
  10818=>"11111101",
  10819=>"11111110",
  10820=>"11111110",
  10821=>"11111110",
  10822=>"00000001",
  10823=>"00000001",
  10824=>"11111101",
  10825=>"11111110",
  10826=>"11111110",
  10827=>"11111110",
  10828=>"11111110",
  10829=>"11111101",
  10830=>"11111110",
  10831=>"00000000",
  10832=>"00000001",
  10833=>"11111101",
  10834=>"11111101",
  10835=>"11111110",
  10836=>"00000000",
  10837=>"11111100",
  10838=>"00000000",
  10839=>"00000001",
  10840=>"11111111",
  10841=>"00000011",
  10842=>"00000001",
  10843=>"11111110",
  10844=>"00000010",
  10845=>"00000001",
  10846=>"00000001",
  10847=>"00000000",
  10848=>"11111110",
  10849=>"00000001",
  10850=>"00000001",
  10851=>"11111111",
  10852=>"00000101",
  10853=>"11111110",
  10854=>"11111101",
  10855=>"11111101",
  10856=>"11111111",
  10857=>"11111110",
  10858=>"00000001",
  10859=>"00000010",
  10860=>"11111111",
  10861=>"00000001",
  10862=>"00000000",
  10863=>"11111111",
  10864=>"00000101",
  10865=>"00000100",
  10866=>"11111111",
  10867=>"11111111",
  10868=>"00000010",
  10869=>"00000010",
  10870=>"11111100",
  10871=>"11111110",
  10872=>"00000001",
  10873=>"00000001",
  10874=>"00000011",
  10875=>"00000001",
  10876=>"00000000",
  10877=>"00000001",
  10878=>"11111101",
  10879=>"00000001",
  10880=>"11111111",
  10881=>"00000001",
  10882=>"11111110",
  10883=>"11111110",
  10884=>"00000000",
  10885=>"11111110",
  10886=>"11111110",
  10887=>"11111110",
  10888=>"11111110",
  10889=>"00000001",
  10890=>"11111110",
  10891=>"11111100",
  10892=>"00000001",
  10893=>"00000010",
  10894=>"00000000",
  10895=>"00000001",
  10896=>"00000001",
  10897=>"00000001",
  10898=>"00000100",
  10899=>"00000001",
  10900=>"00000000",
  10901=>"00000010",
  10902=>"11111110",
  10903=>"11111101",
  10904=>"00000000",
  10905=>"00000010",
  10906=>"00000001",
  10907=>"11111100",
  10908=>"11111111",
  10909=>"00000001",
  10910=>"00000001",
  10911=>"00000001",
  10912=>"00000000",
  10913=>"00000010",
  10914=>"00000011",
  10915=>"11111111",
  10916=>"11111101",
  10917=>"11111110",
  10918=>"00000000",
  10919=>"00000000",
  10920=>"11111110",
  10921=>"00000101",
  10922=>"00000000",
  10923=>"00000010",
  10924=>"00000000",
  10925=>"11111101",
  10926=>"11111110",
  10927=>"00000000",
  10928=>"00000010",
  10929=>"11111110",
  10930=>"11111110",
  10931=>"00000001",
  10932=>"11111101",
  10933=>"00000001",
  10934=>"00000011",
  10935=>"00000011",
  10936=>"11111111",
  10937=>"00000000",
  10938=>"00000011",
  10939=>"00000100",
  10940=>"11111111",
  10941=>"00000001",
  10942=>"11111111",
  10943=>"11111101",
  10944=>"00000100",
  10945=>"11111111",
  10946=>"00000000",
  10947=>"00000010",
  10948=>"00000000",
  10949=>"11111101",
  10950=>"11111110",
  10951=>"00000000",
  10952=>"00000001",
  10953=>"00000110",
  10954=>"00000001",
  10955=>"00000001",
  10956=>"11111100",
  10957=>"00000000",
  10958=>"11111110",
  10959=>"00000010",
  10960=>"00000010",
  10961=>"11111111",
  10962=>"11111111",
  10963=>"11111101",
  10964=>"00000001",
  10965=>"11111101",
  10966=>"00000101",
  10967=>"11111110",
  10968=>"00000010",
  10969=>"00000010",
  10970=>"00000011",
  10971=>"11111111",
  10972=>"00000000",
  10973=>"00000000",
  10974=>"11111110",
  10975=>"11111110",
  10976=>"00000001",
  10977=>"00000101",
  10978=>"11111101",
  10979=>"11111111",
  10980=>"00000001",
  10981=>"11111110",
  10982=>"11111100",
  10983=>"00000000",
  10984=>"11111111",
  10985=>"11111111",
  10986=>"11111111",
  10987=>"11111111",
  10988=>"11111111",
  10989=>"00000010",
  10990=>"11111111",
  10991=>"11111101",
  10992=>"11111100",
  10993=>"00000001",
  10994=>"11111111",
  10995=>"00000010",
  10996=>"00000011",
  10997=>"11111110",
  10998=>"11111101",
  10999=>"00000001",
  11000=>"00000011",
  11001=>"11111110",
  11002=>"11111110",
  11003=>"11111111",
  11004=>"11111111",
  11005=>"00000000",
  11006=>"00000010",
  11007=>"11111110",
  11008=>"11111110",
  11009=>"00000010",
  11010=>"00000010",
  11011=>"11111101",
  11012=>"11111110",
  11013=>"00000001",
  11014=>"00000010",
  11015=>"11111111",
  11016=>"11111101",
  11017=>"11111110",
  11018=>"11111101",
  11019=>"11111110",
  11020=>"00000000",
  11021=>"00000000",
  11022=>"00000000",
  11023=>"00000001",
  11024=>"11111101",
  11025=>"11111111",
  11026=>"00000001",
  11027=>"11111110",
  11028=>"11111111",
  11029=>"00000000",
  11030=>"00000010",
  11031=>"00000000",
  11032=>"00000011",
  11033=>"11111100",
  11034=>"11111101",
  11035=>"11111110",
  11036=>"00000000",
  11037=>"11111100",
  11038=>"11111111",
  11039=>"00000011",
  11040=>"11111101",
  11041=>"11111111",
  11042=>"00000010",
  11043=>"11111110",
  11044=>"00000100",
  11045=>"00000010",
  11046=>"00000110",
  11047=>"11111101",
  11048=>"00000001",
  11049=>"11111100",
  11050=>"11111110",
  11051=>"11111111",
  11052=>"11111111",
  11053=>"00000000",
  11054=>"11111101",
  11055=>"00000000",
  11056=>"11111110",
  11057=>"00000011",
  11058=>"00000001",
  11059=>"00000001",
  11060=>"00000000",
  11061=>"00000001",
  11062=>"11111110",
  11063=>"11111110",
  11064=>"00000000",
  11065=>"00000000",
  11066=>"00000001",
  11067=>"11111101",
  11068=>"00000000",
  11069=>"11111101",
  11070=>"00000010",
  11071=>"00000001",
  11072=>"11111101",
  11073=>"00000010",
  11074=>"11111101",
  11075=>"11111101",
  11076=>"00000001",
  11077=>"11111101",
  11078=>"11111101",
  11079=>"11111111",
  11080=>"11111101",
  11081=>"00000000",
  11082=>"00000001",
  11083=>"11111111",
  11084=>"11111101",
  11085=>"00000010",
  11086=>"00000010",
  11087=>"11111110",
  11088=>"00000001",
  11089=>"00000000",
  11090=>"00000101",
  11091=>"11111110",
  11092=>"11111110",
  11093=>"11111110",
  11094=>"11111111",
  11095=>"00000100",
  11096=>"00000001",
  11097=>"00000101",
  11098=>"11111101",
  11099=>"11111110",
  11100=>"11111101",
  11101=>"00000010",
  11102=>"00000100",
  11103=>"11111110",
  11104=>"00000010",
  11105=>"11111100",
  11106=>"00000000",
  11107=>"11111101",
  11108=>"11111101",
  11109=>"00000001",
  11110=>"00000000",
  11111=>"11111101",
  11112=>"11111110",
  11113=>"00000011",
  11114=>"11111111",
  11115=>"11111111",
  11116=>"00000000",
  11117=>"11111111",
  11118=>"00000001",
  11119=>"11111110",
  11120=>"11111101",
  11121=>"00000000",
  11122=>"11111111",
  11123=>"11111110",
  11124=>"00000010",
  11125=>"00000010",
  11126=>"11111101",
  11127=>"00000001",
  11128=>"00000000",
  11129=>"11111110",
  11130=>"00000001",
  11131=>"00000010",
  11132=>"11111101",
  11133=>"00000010",
  11134=>"11111101",
  11135=>"11111100",
  11136=>"00000010",
  11137=>"00000000",
  11138=>"11111111",
  11139=>"00000101",
  11140=>"11111110",
  11141=>"00000010",
  11142=>"00000011",
  11143=>"00000001",
  11144=>"11111110",
  11145=>"00000001",
  11146=>"11111110",
  11147=>"00000001",
  11148=>"00000100",
  11149=>"00000010",
  11150=>"00000001",
  11151=>"11111101",
  11152=>"00000001",
  11153=>"11111101",
  11154=>"11111111",
  11155=>"00000010",
  11156=>"00000101",
  11157=>"11111111",
  11158=>"11111110",
  11159=>"00000000",
  11160=>"00000001",
  11161=>"11111111",
  11162=>"11111110",
  11163=>"11111101",
  11164=>"11111101",
  11165=>"00000000",
  11166=>"11111101",
  11167=>"11111100",
  11168=>"11111101",
  11169=>"11111111",
  11170=>"11111101",
  11171=>"00000000",
  11172=>"11111110",
  11173=>"11111101",
  11174=>"11111101",
  11175=>"00000011",
  11176=>"00000000",
  11177=>"11111111",
  11178=>"11111110",
  11179=>"11111111",
  11180=>"11111110",
  11181=>"11111101",
  11182=>"11111110",
  11183=>"11111100",
  11184=>"11111111",
  11185=>"00000000",
  11186=>"00000000",
  11187=>"00000000",
  11188=>"11111111",
  11189=>"00000010",
  11190=>"11111101",
  11191=>"11111111",
  11192=>"11111110",
  11193=>"00000000",
  11194=>"11111111",
  11195=>"00000001",
  11196=>"00001000",
  11197=>"00000000",
  11198=>"00000001",
  11199=>"11111110",
  11200=>"00000001",
  11201=>"00000010",
  11202=>"11111111",
  11203=>"11111110",
  11204=>"00000000",
  11205=>"00000000",
  11206=>"00000001",
  11207=>"11111110",
  11208=>"00000010",
  11209=>"00000000",
  11210=>"11111111",
  11211=>"11111111",
  11212=>"00000010",
  11213=>"00000100",
  11214=>"11111111",
  11215=>"00000001",
  11216=>"00000001",
  11217=>"11111100",
  11218=>"11111111",
  11219=>"11111110",
  11220=>"11111101",
  11221=>"11111101",
  11222=>"00000000",
  11223=>"11111111",
  11224=>"00000010",
  11225=>"00000011",
  11226=>"00000001",
  11227=>"00000010",
  11228=>"11111110",
  11229=>"11111110",
  11230=>"00000000",
  11231=>"11111101",
  11232=>"00000011",
  11233=>"11111111",
  11234=>"11111110",
  11235=>"11111110",
  11236=>"00000001",
  11237=>"11111110",
  11238=>"11111111",
  11239=>"00000001",
  11240=>"00000000",
  11241=>"11111101",
  11242=>"11111100",
  11243=>"00000011",
  11244=>"00000010",
  11245=>"11111111",
  11246=>"00000001",
  11247=>"00000000",
  11248=>"11111111",
  11249=>"00000001",
  11250=>"00000001",
  11251=>"00000000",
  11252=>"00000101",
  11253=>"11111111",
  11254=>"00000011",
  11255=>"00000001",
  11256=>"11111101",
  11257=>"00000000",
  11258=>"11111101",
  11259=>"00000001",
  11260=>"00000001",
  11261=>"00000001",
  11262=>"00000010",
  11263=>"00000000",
  11264=>"11111101",
  11265=>"11111111",
  11266=>"11111101",
  11267=>"00000100",
  11268=>"00000000",
  11269=>"00000001",
  11270=>"00000000",
  11271=>"11111011",
  11272=>"00000001",
  11273=>"00000010",
  11274=>"00000101",
  11275=>"00000000",
  11276=>"00000001",
  11277=>"00000000",
  11278=>"11111101",
  11279=>"11111111",
  11280=>"11111111",
  11281=>"11111101",
  11282=>"00000101",
  11283=>"11111110",
  11284=>"11111111",
  11285=>"00000011",
  11286=>"00000101",
  11287=>"00000011",
  11288=>"11111110",
  11289=>"11111110",
  11290=>"11111110",
  11291=>"11111100",
  11292=>"11111110",
  11293=>"11111110",
  11294=>"00000000",
  11295=>"11111101",
  11296=>"00000010",
  11297=>"00000001",
  11298=>"00000100",
  11299=>"11111101",
  11300=>"11111110",
  11301=>"11111111",
  11302=>"11111111",
  11303=>"00000100",
  11304=>"00000101",
  11305=>"11111110",
  11306=>"00000001",
  11307=>"00000000",
  11308=>"00000001",
  11309=>"00000001",
  11310=>"00000010",
  11311=>"11111110",
  11312=>"00000010",
  11313=>"00000011",
  11314=>"00000000",
  11315=>"11111111",
  11316=>"00000001",
  11317=>"00000000",
  11318=>"11111111",
  11319=>"00000001",
  11320=>"00000011",
  11321=>"00000000",
  11322=>"00000101",
  11323=>"00000011",
  11324=>"00000011",
  11325=>"00000000",
  11326=>"00000011",
  11327=>"00000001",
  11328=>"11111010",
  11329=>"00000011",
  11330=>"00000011",
  11331=>"11111111",
  11332=>"00000001",
  11333=>"11111101",
  11334=>"11111101",
  11335=>"00000011",
  11336=>"11111110",
  11337=>"00000001",
  11338=>"00000001",
  11339=>"00000010",
  11340=>"11111110",
  11341=>"11111111",
  11342=>"11111101",
  11343=>"11111101",
  11344=>"11111111",
  11345=>"11111111",
  11346=>"11111110",
  11347=>"00000100",
  11348=>"00000010",
  11349=>"00000000",
  11350=>"00000000",
  11351=>"11111111",
  11352=>"00000000",
  11353=>"00000001",
  11354=>"11111101",
  11355=>"11111100",
  11356=>"11111111",
  11357=>"11111111",
  11358=>"00000011",
  11359=>"11111110",
  11360=>"11111110",
  11361=>"00000100",
  11362=>"00000001",
  11363=>"00000001",
  11364=>"00000000",
  11365=>"00000011",
  11366=>"00000000",
  11367=>"11111101",
  11368=>"11111111",
  11369=>"00000001",
  11370=>"11111101",
  11371=>"00000000",
  11372=>"00000000",
  11373=>"11111100",
  11374=>"00000000",
  11375=>"00000010",
  11376=>"00000000",
  11377=>"00000100",
  11378=>"00000010",
  11379=>"11111101",
  11380=>"00000000",
  11381=>"11111110",
  11382=>"00000001",
  11383=>"00000010",
  11384=>"11111101",
  11385=>"11111101",
  11386=>"00000010",
  11387=>"11111101",
  11388=>"11111110",
  11389=>"00000010",
  11390=>"00000001",
  11391=>"00000000",
  11392=>"00000000",
  11393=>"11111110",
  11394=>"00000010",
  11395=>"11111110",
  11396=>"11111110",
  11397=>"11111110",
  11398=>"11111111",
  11399=>"00000001",
  11400=>"11111010",
  11401=>"00000000",
  11402=>"11111011",
  11403=>"00000000",
  11404=>"00000000",
  11405=>"00000000",
  11406=>"00000000",
  11407=>"11111011",
  11408=>"00000001",
  11409=>"11111100",
  11410=>"11111111",
  11411=>"00000101",
  11412=>"00000011",
  11413=>"11111101",
  11414=>"00000000",
  11415=>"00000011",
  11416=>"11111110",
  11417=>"11111111",
  11418=>"11111101",
  11419=>"00000010",
  11420=>"11111111",
  11421=>"11111110",
  11422=>"00000011",
  11423=>"00000000",
  11424=>"11111111",
  11425=>"00000101",
  11426=>"00000011",
  11427=>"00000010",
  11428=>"00000100",
  11429=>"11111101",
  11430=>"00000010",
  11431=>"11111111",
  11432=>"11111111",
  11433=>"00000110",
  11434=>"00000010",
  11435=>"00000011",
  11436=>"11111111",
  11437=>"11111110",
  11438=>"00000100",
  11439=>"11111110",
  11440=>"11111111",
  11441=>"00000000",
  11442=>"11111101",
  11443=>"11111101",
  11444=>"00000001",
  11445=>"00000011",
  11446=>"11111100",
  11447=>"11111111",
  11448=>"11111111",
  11449=>"00000001",
  11450=>"11111110",
  11451=>"11111111",
  11452=>"00000001",
  11453=>"11111111",
  11454=>"11111100",
  11455=>"00000100",
  11456=>"00000010",
  11457=>"00000010",
  11458=>"11111111",
  11459=>"00000101",
  11460=>"00000101",
  11461=>"00000001",
  11462=>"11111110",
  11463=>"11111111",
  11464=>"11111110",
  11465=>"00000001",
  11466=>"11111110",
  11467=>"00000100",
  11468=>"00000101",
  11469=>"00000000",
  11470=>"11111100",
  11471=>"11111101",
  11472=>"00000001",
  11473=>"11111100",
  11474=>"00000001",
  11475=>"11111101",
  11476=>"00000010",
  11477=>"00000001",
  11478=>"00000011",
  11479=>"11111011",
  11480=>"11111110",
  11481=>"11111100",
  11482=>"00000000",
  11483=>"00000100",
  11484=>"11111110",
  11485=>"00000000",
  11486=>"00000011",
  11487=>"11111110",
  11488=>"11111110",
  11489=>"11111101",
  11490=>"11111110",
  11491=>"11111110",
  11492=>"11111111",
  11493=>"11111101",
  11494=>"11111111",
  11495=>"00000010",
  11496=>"00000101",
  11497=>"11111100",
  11498=>"00000011",
  11499=>"00000011",
  11500=>"00000001",
  11501=>"00000100",
  11502=>"00000001",
  11503=>"11111110",
  11504=>"00000000",
  11505=>"00000011",
  11506=>"11111110",
  11507=>"00000011",
  11508=>"00000000",
  11509=>"11111011",
  11510=>"00000010",
  11511=>"00000100",
  11512=>"11111110",
  11513=>"11111111",
  11514=>"00000001",
  11515=>"00000000",
  11516=>"00000100",
  11517=>"00000010",
  11518=>"00000000",
  11519=>"11111111",
  11520=>"00000001",
  11521=>"00000001",
  11522=>"00000000",
  11523=>"00000101",
  11524=>"00000010",
  11525=>"11111110",
  11526=>"00000000",
  11527=>"00000011",
  11528=>"11111111",
  11529=>"00000000",
  11530=>"00000100",
  11531=>"00000011",
  11532=>"11111110",
  11533=>"11111101",
  11534=>"00000101",
  11535=>"11111100",
  11536=>"00000100",
  11537=>"11111101",
  11538=>"00000010",
  11539=>"00000000",
  11540=>"11111110",
  11541=>"00000000",
  11542=>"11111111",
  11543=>"00000001",
  11544=>"00000010",
  11545=>"11111111",
  11546=>"00000010",
  11547=>"00000100",
  11548=>"00000010",
  11549=>"11111110",
  11550=>"11111110",
  11551=>"11111100",
  11552=>"00000011",
  11553=>"00000011",
  11554=>"00000100",
  11555=>"00000010",
  11556=>"11111100",
  11557=>"00000001",
  11558=>"11111111",
  11559=>"00000001",
  11560=>"11111111",
  11561=>"11111100",
  11562=>"11111110",
  11563=>"00000001",
  11564=>"11111110",
  11565=>"11111101",
  11566=>"00000001",
  11567=>"00000000",
  11568=>"11111110",
  11569=>"11111110",
  11570=>"00000100",
  11571=>"00000001",
  11572=>"00000001",
  11573=>"00000000",
  11574=>"00000110",
  11575=>"00000001",
  11576=>"00000100",
  11577=>"00000001",
  11578=>"00000001",
  11579=>"11111110",
  11580=>"11111101",
  11581=>"00000001",
  11582=>"00000000",
  11583=>"00000011",
  11584=>"00000000",
  11585=>"11111101",
  11586=>"00000001",
  11587=>"00000000",
  11588=>"00000011",
  11589=>"11111011",
  11590=>"00000100",
  11591=>"11111111",
  11592=>"11111111",
  11593=>"11111101",
  11594=>"11111110",
  11595=>"00000000",
  11596=>"11111100",
  11597=>"00000101",
  11598=>"11111101",
  11599=>"11111111",
  11600=>"11111110",
  11601=>"00000100",
  11602=>"00000100",
  11603=>"00000011",
  11604=>"00000000",
  11605=>"00000101",
  11606=>"00000010",
  11607=>"11111100",
  11608=>"00000000",
  11609=>"11111101",
  11610=>"11111110",
  11611=>"00000001",
  11612=>"00000011",
  11613=>"00000000",
  11614=>"00000011",
  11615=>"11111101",
  11616=>"00000100",
  11617=>"00000000",
  11618=>"00000001",
  11619=>"00000010",
  11620=>"11111111",
  11621=>"00000000",
  11622=>"00000001",
  11623=>"11111111",
  11624=>"00000100",
  11625=>"11111011",
  11626=>"00000010",
  11627=>"00000000",
  11628=>"00000001",
  11629=>"00000001",
  11630=>"11111110",
  11631=>"11111101",
  11632=>"00000010",
  11633=>"00000000",
  11634=>"00000010",
  11635=>"11111111",
  11636=>"11111100",
  11637=>"11111111",
  11638=>"11111101",
  11639=>"00000011",
  11640=>"00000000",
  11641=>"11111110",
  11642=>"00000011",
  11643=>"11111110",
  11644=>"00000001",
  11645=>"00000000",
  11646=>"11111111",
  11647=>"00000010",
  11648=>"00000011",
  11649=>"11111110",
  11650=>"11111110",
  11651=>"11111110",
  11652=>"00000010",
  11653=>"00000011",
  11654=>"00000010",
  11655=>"00000010",
  11656=>"00000101",
  11657=>"11111110",
  11658=>"00000000",
  11659=>"00000101",
  11660=>"11111100",
  11661=>"00000100",
  11662=>"00000110",
  11663=>"00000011",
  11664=>"11111111",
  11665=>"00000110",
  11666=>"00000010",
  11667=>"11111111",
  11668=>"11111100",
  11669=>"00000010",
  11670=>"00000000",
  11671=>"00000010",
  11672=>"11111101",
  11673=>"11111111",
  11674=>"11111100",
  11675=>"00000110",
  11676=>"00000001",
  11677=>"11111111",
  11678=>"11111111",
  11679=>"11111111",
  11680=>"00000010",
  11681=>"00000010",
  11682=>"11111011",
  11683=>"11111111",
  11684=>"00000001",
  11685=>"11111111",
  11686=>"11111101",
  11687=>"00000000",
  11688=>"00000100",
  11689=>"00000000",
  11690=>"11111111",
  11691=>"00000101",
  11692=>"00000000",
  11693=>"11111101",
  11694=>"00000001",
  11695=>"00000010",
  11696=>"11111101",
  11697=>"00000010",
  11698=>"11111110",
  11699=>"11111111",
  11700=>"11111101",
  11701=>"00000011",
  11702=>"11111101",
  11703=>"11111110",
  11704=>"00000000",
  11705=>"11111101",
  11706=>"11111111",
  11707=>"00000010",
  11708=>"00000001",
  11709=>"00000001",
  11710=>"00000010",
  11711=>"11111111",
  11712=>"00000001",
  11713=>"00000101",
  11714=>"11111111",
  11715=>"00000100",
  11716=>"00000000",
  11717=>"00000010",
  11718=>"11111111",
  11719=>"00000000",
  11720=>"00000000",
  11721=>"00000010",
  11722=>"00000000",
  11723=>"11111110",
  11724=>"11111101",
  11725=>"00000011",
  11726=>"11111100",
  11727=>"11111110",
  11728=>"11111111",
  11729=>"00000001",
  11730=>"00000010",
  11731=>"11111110",
  11732=>"00000000",
  11733=>"00000001",
  11734=>"00000100",
  11735=>"00000000",
  11736=>"00000001",
  11737=>"00000010",
  11738=>"00000010",
  11739=>"11111110",
  11740=>"00000011",
  11741=>"00000001",
  11742=>"00000001",
  11743=>"11111110",
  11744=>"00000010",
  11745=>"11111011",
  11746=>"11111101",
  11747=>"11111111",
  11748=>"11111110",
  11749=>"00000010",
  11750=>"00000010",
  11751=>"00000000",
  11752=>"00000001",
  11753=>"00000001",
  11754=>"00000000",
  11755=>"11111111",
  11756=>"00000001",
  11757=>"00000010",
  11758=>"00000101",
  11759=>"00000000",
  11760=>"11111110",
  11761=>"00000000",
  11762=>"11111101",
  11763=>"00000000",
  11764=>"11111110",
  11765=>"00000000",
  11766=>"00000010",
  11767=>"00000100",
  11768=>"00000000",
  11769=>"00000001",
  11770=>"11111110",
  11771=>"00000010",
  11772=>"11111110",
  11773=>"00000010",
  11774=>"00000100",
  11775=>"11111100",
  11776=>"11111101",
  11777=>"00000010",
  11778=>"11111101",
  11779=>"11111100",
  11780=>"00000010",
  11781=>"00000011",
  11782=>"11111110",
  11783=>"00000011",
  11784=>"00000000",
  11785=>"11111100",
  11786=>"00000001",
  11787=>"00000101",
  11788=>"00000001",
  11789=>"00000001",
  11790=>"00000010",
  11791=>"00000011",
  11792=>"11111100",
  11793=>"00000011",
  11794=>"11111111",
  11795=>"11111101",
  11796=>"11111101",
  11797=>"00000000",
  11798=>"00000000",
  11799=>"00000100",
  11800=>"00000100",
  11801=>"00000000",
  11802=>"00000000",
  11803=>"11111111",
  11804=>"00000001",
  11805=>"00000100",
  11806=>"11111110",
  11807=>"11111110",
  11808=>"00000011",
  11809=>"00000000",
  11810=>"11111111",
  11811=>"11111111",
  11812=>"11111101",
  11813=>"00000011",
  11814=>"11111111",
  11815=>"00000011",
  11816=>"11111100",
  11817=>"00000100",
  11818=>"11111111",
  11819=>"00000101",
  11820=>"00000000",
  11821=>"11111110",
  11822=>"00000001",
  11823=>"00000010",
  11824=>"00000011",
  11825=>"11111111",
  11826=>"11111101",
  11827=>"11111111",
  11828=>"00000000",
  11829=>"11111110",
  11830=>"11111101",
  11831=>"00000010",
  11832=>"00000101",
  11833=>"00000011",
  11834=>"00000010",
  11835=>"11111110",
  11836=>"00000001",
  11837=>"11111110",
  11838=>"00000001",
  11839=>"00000001",
  11840=>"00000010",
  11841=>"11111011",
  11842=>"00000001",
  11843=>"00000000",
  11844=>"00000011",
  11845=>"00000011",
  11846=>"11111111",
  11847=>"00000001",
  11848=>"00000101",
  11849=>"00000100",
  11850=>"00000010",
  11851=>"00000000",
  11852=>"11111110",
  11853=>"00000001",
  11854=>"11111110",
  11855=>"11111101",
  11856=>"00000001",
  11857=>"11111100",
  11858=>"11111111",
  11859=>"11111110",
  11860=>"00000011",
  11861=>"00000000",
  11862=>"00000011",
  11863=>"00000001",
  11864=>"11111110",
  11865=>"00000000",
  11866=>"00000001",
  11867=>"11111111",
  11868=>"11111110",
  11869=>"11111110",
  11870=>"00000010",
  11871=>"11111111",
  11872=>"11111101",
  11873=>"00000001",
  11874=>"00000101",
  11875=>"11111100",
  11876=>"00000001",
  11877=>"11111110",
  11878=>"00000011",
  11879=>"00000000",
  11880=>"11111110",
  11881=>"00000001",
  11882=>"00000100",
  11883=>"11111111",
  11884=>"11111101",
  11885=>"11111100",
  11886=>"00000000",
  11887=>"00000010",
  11888=>"11111011",
  11889=>"00000100",
  11890=>"11111101",
  11891=>"00000010",
  11892=>"11111101",
  11893=>"00000011",
  11894=>"00000011",
  11895=>"11111101",
  11896=>"00000000",
  11897=>"00000001",
  11898=>"00000100",
  11899=>"00000011",
  11900=>"00000000",
  11901=>"00000010",
  11902=>"11111101",
  11903=>"00000001",
  11904=>"00000000",
  11905=>"00000101",
  11906=>"00000001",
  11907=>"11111101",
  11908=>"11111101",
  11909=>"00000001",
  11910=>"00000001",
  11911=>"11111111",
  11912=>"11111111",
  11913=>"00000000",
  11914=>"00000011",
  11915=>"00000001",
  11916=>"00000010",
  11917=>"00000000",
  11918=>"11111110",
  11919=>"00000010",
  11920=>"11111101",
  11921=>"11111111",
  11922=>"00000010",
  11923=>"11111111",
  11924=>"11111101",
  11925=>"00000000",
  11926=>"00000001",
  11927=>"11111101",
  11928=>"11111110",
  11929=>"11111101",
  11930=>"11111111",
  11931=>"00000010",
  11932=>"11111100",
  11933=>"11111101",
  11934=>"11111111",
  11935=>"00000010",
  11936=>"00000000",
  11937=>"11111101",
  11938=>"00000011",
  11939=>"00000000",
  11940=>"11111101",
  11941=>"11111100",
  11942=>"11111011",
  11943=>"00000000",
  11944=>"00000001",
  11945=>"00000110",
  11946=>"11111101",
  11947=>"11111111",
  11948=>"11111111",
  11949=>"11111110",
  11950=>"11111110",
  11951=>"11111101",
  11952=>"00000001",
  11953=>"00000001",
  11954=>"00000001",
  11955=>"00000011",
  11956=>"00000000",
  11957=>"11111100",
  11958=>"11111111",
  11959=>"00000000",
  11960=>"00000000",
  11961=>"00000000",
  11962=>"00000000",
  11963=>"00000010",
  11964=>"00000100",
  11965=>"00000010",
  11966=>"11111101",
  11967=>"00000000",
  11968=>"00000011",
  11969=>"00000010",
  11970=>"00000100",
  11971=>"00000110",
  11972=>"00000011",
  11973=>"11111101",
  11974=>"11111110",
  11975=>"11111110",
  11976=>"11111101",
  11977=>"00000000",
  11978=>"00000000",
  11979=>"11111110",
  11980=>"00000011",
  11981=>"00000010",
  11982=>"00000001",
  11983=>"00000000",
  11984=>"00000010",
  11985=>"11111110",
  11986=>"11111111",
  11987=>"11111011",
  11988=>"00000001",
  11989=>"00000010",
  11990=>"00000010",
  11991=>"11111100",
  11992=>"11111111",
  11993=>"00000001",
  11994=>"00000001",
  11995=>"11111111",
  11996=>"11111111",
  11997=>"00000010",
  11998=>"00000010",
  11999=>"00000000",
  12000=>"11111110",
  12001=>"00000010",
  12002=>"11111111",
  12003=>"00000011",
  12004=>"00000010",
  12005=>"00000001",
  12006=>"11111111",
  12007=>"00000011",
  12008=>"11111101",
  12009=>"00000100",
  12010=>"00000100",
  12011=>"00000101",
  12012=>"00000001",
  12013=>"00000001",
  12014=>"11111111",
  12015=>"11111111",
  12016=>"11111100",
  12017=>"00000001",
  12018=>"11111101",
  12019=>"00000001",
  12020=>"11111111",
  12021=>"00000000",
  12022=>"00000001",
  12023=>"00000011",
  12024=>"11111111",
  12025=>"11111110",
  12026=>"11111101",
  12027=>"00000011",
  12028=>"11111101",
  12029=>"00000011",
  12030=>"11111101",
  12031=>"11111111",
  12032=>"00000000",
  12033=>"00000010",
  12034=>"11111111",
  12035=>"00000110",
  12036=>"11111110",
  12037=>"00000010",
  12038=>"00000011",
  12039=>"11111011",
  12040=>"11111101",
  12041=>"00000001",
  12042=>"11111100",
  12043=>"11111100",
  12044=>"11111111",
  12045=>"00000001",
  12046=>"11111101",
  12047=>"00000000",
  12048=>"11111110",
  12049=>"11111111",
  12050=>"11111100",
  12051=>"00000001",
  12052=>"00000000",
  12053=>"00000010",
  12054=>"11111101",
  12055=>"00000011",
  12056=>"11111101",
  12057=>"11111101",
  12058=>"00000011",
  12059=>"11111111",
  12060=>"00000011",
  12061=>"00000101",
  12062=>"00000000",
  12063=>"00000010",
  12064=>"00000001",
  12065=>"00000100",
  12066=>"11111101",
  12067=>"00000001",
  12068=>"00000000",
  12069=>"00000100",
  12070=>"00000100",
  12071=>"00000100",
  12072=>"11111111",
  12073=>"00000100",
  12074=>"11111101",
  12075=>"00000001",
  12076=>"11111110",
  12077=>"11111110",
  12078=>"11111100",
  12079=>"11111111",
  12080=>"00000110",
  12081=>"00000000",
  12082=>"00000100",
  12083=>"11111101",
  12084=>"00000011",
  12085=>"11111011",
  12086=>"11111110",
  12087=>"11111101",
  12088=>"11111110",
  12089=>"00000101",
  12090=>"11111111",
  12091=>"11111110",
  12092=>"00000011",
  12093=>"00000011",
  12094=>"11111110",
  12095=>"11111111",
  12096=>"00000100",
  12097=>"00000000",
  12098=>"11111101",
  12099=>"00000000",
  12100=>"11111101",
  12101=>"00000011",
  12102=>"00000001",
  12103=>"11111110",
  12104=>"00000010",
  12105=>"11111111",
  12106=>"11111100",
  12107=>"11111110",
  12108=>"00000010",
  12109=>"11111101",
  12110=>"00000010",
  12111=>"00000000",
  12112=>"11111110",
  12113=>"11111111",
  12114=>"00000101",
  12115=>"11111101",
  12116=>"11111101",
  12117=>"00000101",
  12118=>"11111110",
  12119=>"11111111",
  12120=>"00000001",
  12121=>"11111101",
  12122=>"00000001",
  12123=>"00000001",
  12124=>"00000000",
  12125=>"00000011",
  12126=>"11111101",
  12127=>"11111111",
  12128=>"11111110",
  12129=>"11111101",
  12130=>"00000000",
  12131=>"11111100",
  12132=>"00000101",
  12133=>"00000011",
  12134=>"00000001",
  12135=>"00000100",
  12136=>"11111011",
  12137=>"00000000",
  12138=>"00000010",
  12139=>"00000010",
  12140=>"00000011",
  12141=>"11111110",
  12142=>"00000000",
  12143=>"00000011",
  12144=>"00000000",
  12145=>"00000001",
  12146=>"11111110",
  12147=>"00000100",
  12148=>"11111110",
  12149=>"11111111",
  12150=>"11111100",
  12151=>"11111110",
  12152=>"11111111",
  12153=>"00000010",
  12154=>"00000011",
  12155=>"11111110",
  12156=>"00000001",
  12157=>"00000101",
  12158=>"11111110",
  12159=>"00000000",
  12160=>"11111110",
  12161=>"00000000",
  12162=>"00000001",
  12163=>"00000101",
  12164=>"00000011",
  12165=>"11111110",
  12166=>"00000100",
  12167=>"00000010",
  12168=>"00000010",
  12169=>"00000011",
  12170=>"00000011",
  12171=>"00000010",
  12172=>"00000010",
  12173=>"11111111",
  12174=>"00000000",
  12175=>"11111111",
  12176=>"00000001",
  12177=>"11111111",
  12178=>"11111010",
  12179=>"00000100",
  12180=>"00000010",
  12181=>"11111111",
  12182=>"11111111",
  12183=>"11111111",
  12184=>"00000100",
  12185=>"11111111",
  12186=>"00000001",
  12187=>"11111111",
  12188=>"11111100",
  12189=>"00000001",
  12190=>"11111101",
  12191=>"11111110",
  12192=>"00000001",
  12193=>"00000011",
  12194=>"11111101",
  12195=>"11111101",
  12196=>"11111101",
  12197=>"00000011",
  12198=>"00000001",
  12199=>"00000110",
  12200=>"00000000",
  12201=>"11111110",
  12202=>"00000001",
  12203=>"11111111",
  12204=>"00000001",
  12205=>"00000110",
  12206=>"00000001",
  12207=>"11111110",
  12208=>"00000001",
  12209=>"00000010",
  12210=>"11111101",
  12211=>"11111111",
  12212=>"00000100",
  12213=>"00000000",
  12214=>"00000010",
  12215=>"00000011",
  12216=>"00000010",
  12217=>"11111111",
  12218=>"00000000",
  12219=>"00000010",
  12220=>"00000111",
  12221=>"00000000",
  12222=>"00000011",
  12223=>"00000000",
  12224=>"11111101",
  12225=>"00000101",
  12226=>"00000000",
  12227=>"11111111",
  12228=>"00000101",
  12229=>"11111101",
  12230=>"11111100",
  12231=>"11111111",
  12232=>"11111111",
  12233=>"00000011",
  12234=>"00000000",
  12235=>"11111101",
  12236=>"00000010",
  12237=>"11111110",
  12238=>"00000001",
  12239=>"11111101",
  12240=>"00000100",
  12241=>"00000010",
  12242=>"11111110",
  12243=>"00000010",
  12244=>"00000000",
  12245=>"11111110",
  12246=>"00000010",
  12247=>"00000100",
  12248=>"00000000",
  12249=>"00000110",
  12250=>"00000000",
  12251=>"11111110",
  12252=>"11111101",
  12253=>"11111110",
  12254=>"00000001",
  12255=>"00000001",
  12256=>"00000000",
  12257=>"11111110",
  12258=>"00000010",
  12259=>"11111111",
  12260=>"11111110",
  12261=>"11111100",
  12262=>"00000000",
  12263=>"11111101",
  12264=>"00000010",
  12265=>"11111111",
  12266=>"00000001",
  12267=>"00000010",
  12268=>"00000001",
  12269=>"00000100",
  12270=>"11111111",
  12271=>"11111110",
  12272=>"00000010",
  12273=>"00000001",
  12274=>"00000101",
  12275=>"11111101",
  12276=>"00000100",
  12277=>"00000000",
  12278=>"00000010",
  12279=>"11111101",
  12280=>"00000010",
  12281=>"00000000",
  12282=>"00000000",
  12283=>"00000101",
  12284=>"11111100",
  12285=>"11111101",
  12286=>"00000010",
  12287=>"11111111",
  12288=>"11111110",
  12289=>"00000000",
  12290=>"00000010",
  12291=>"00000001",
  12292=>"00000000",
  12293=>"00000001",
  12294=>"00000010",
  12295=>"11111110",
  12296=>"00000010",
  12297=>"11111110",
  12298=>"00000000",
  12299=>"11111101",
  12300=>"11111110",
  12301=>"11111110",
  12302=>"11111111",
  12303=>"00000100",
  12304=>"11111101",
  12305=>"11111110",
  12306=>"11111100",
  12307=>"00000010",
  12308=>"00000100",
  12309=>"00000011",
  12310=>"00000101",
  12311=>"11111111",
  12312=>"00000000",
  12313=>"00000000",
  12314=>"11111110",
  12315=>"11111111",
  12316=>"11111111",
  12317=>"00000010",
  12318=>"00000010",
  12319=>"00000001",
  12320=>"11111110",
  12321=>"00000001",
  12322=>"11111101",
  12323=>"00000100",
  12324=>"11111110",
  12325=>"11111101",
  12326=>"11111111",
  12327=>"00000011",
  12328=>"11111101",
  12329=>"00000101",
  12330=>"11111110",
  12331=>"11111111",
  12332=>"11111101",
  12333=>"11111111",
  12334=>"11111111",
  12335=>"11111101",
  12336=>"00000000",
  12337=>"11111111",
  12338=>"00000010",
  12339=>"11111111",
  12340=>"11111111",
  12341=>"00000010",
  12342=>"00000001",
  12343=>"00000011",
  12344=>"11111111",
  12345=>"11111101",
  12346=>"11111110",
  12347=>"00000000",
  12348=>"11111110",
  12349=>"11111110",
  12350=>"11111110",
  12351=>"11111111",
  12352=>"00000010",
  12353=>"00000000",
  12354=>"11111110",
  12355=>"11111111",
  12356=>"00000000",
  12357=>"11111110",
  12358=>"11111110",
  12359=>"00000001",
  12360=>"11111110",
  12361=>"11111110",
  12362=>"11111110",
  12363=>"11111110",
  12364=>"00000001",
  12365=>"11111111",
  12366=>"11111110",
  12367=>"11111111",
  12368=>"00000011",
  12369=>"11111110",
  12370=>"00000010",
  12371=>"00000010",
  12372=>"00000011",
  12373=>"00000001",
  12374=>"00000000",
  12375=>"11111110",
  12376=>"00000001",
  12377=>"00000011",
  12378=>"00000001",
  12379=>"00000010",
  12380=>"11111110",
  12381=>"11111101",
  12382=>"11111101",
  12383=>"11111101",
  12384=>"00000001",
  12385=>"11111111",
  12386=>"11111111",
  12387=>"11111110",
  12388=>"00000000",
  12389=>"00000000",
  12390=>"00000010",
  12391=>"00000011",
  12392=>"00000010",
  12393=>"00000001",
  12394=>"00000101",
  12395=>"11111111",
  12396=>"00000011",
  12397=>"11111101",
  12398=>"00000010",
  12399=>"11111110",
  12400=>"00000000",
  12401=>"00000001",
  12402=>"11111101",
  12403=>"11111110",
  12404=>"11111101",
  12405=>"00000011",
  12406=>"11111111",
  12407=>"00000001",
  12408=>"00000100",
  12409=>"11111111",
  12410=>"00000000",
  12411=>"00000001",
  12412=>"11111111",
  12413=>"11111111",
  12414=>"00000001",
  12415=>"00000010",
  12416=>"00000010",
  12417=>"11111101",
  12418=>"00000010",
  12419=>"00000000",
  12420=>"00000001",
  12421=>"00000001",
  12422=>"11111111",
  12423=>"00000010",
  12424=>"00000011",
  12425=>"11111110",
  12426=>"00000011",
  12427=>"11111101",
  12428=>"00000000",
  12429=>"00000010",
  12430=>"11111111",
  12431=>"00000011",
  12432=>"11111110",
  12433=>"11111111",
  12434=>"00000010",
  12435=>"00000000",
  12436=>"11111101",
  12437=>"11111110",
  12438=>"11111111",
  12439=>"00000001",
  12440=>"11111111",
  12441=>"00000110",
  12442=>"11111110",
  12443=>"00000000",
  12444=>"00000000",
  12445=>"11111110",
  12446=>"00000000",
  12447=>"11111111",
  12448=>"11111111",
  12449=>"00000000",
  12450=>"11111110",
  12451=>"11111110",
  12452=>"11111111",
  12453=>"00000001",
  12454=>"00000001",
  12455=>"11111111",
  12456=>"00000100",
  12457=>"11111111",
  12458=>"00000000",
  12459=>"11111101",
  12460=>"11111101",
  12461=>"00000011",
  12462=>"11111101",
  12463=>"00000001",
  12464=>"11111101",
  12465=>"00000011",
  12466=>"11111110",
  12467=>"11111110",
  12468=>"11111111",
  12469=>"00000000",
  12470=>"00000001",
  12471=>"00000011",
  12472=>"00000000",
  12473=>"11111111",
  12474=>"00000001",
  12475=>"11111110",
  12476=>"00000000",
  12477=>"00000010",
  12478=>"00000001",
  12479=>"00000101",
  12480=>"11111111",
  12481=>"00000000",
  12482=>"00000011",
  12483=>"00000010",
  12484=>"11111101",
  12485=>"00000000",
  12486=>"11111110",
  12487=>"00000010",
  12488=>"00000011",
  12489=>"00000000",
  12490=>"11111101",
  12491=>"11111111",
  12492=>"11111111",
  12493=>"11111110",
  12494=>"00000001",
  12495=>"11111111",
  12496=>"11111101",
  12497=>"00000010",
  12498=>"11111111",
  12499=>"11111111",
  12500=>"00000000",
  12501=>"11111110",
  12502=>"11111110",
  12503=>"11111101",
  12504=>"00000010",
  12505=>"00000000",
  12506=>"11111110",
  12507=>"11111110",
  12508=>"00000000",
  12509=>"00000111",
  12510=>"11111110",
  12511=>"00000011",
  12512=>"11111111",
  12513=>"11111111",
  12514=>"00000010",
  12515=>"00000000",
  12516=>"00000010",
  12517=>"00000011",
  12518=>"11111110",
  12519=>"00000000",
  12520=>"00000000",
  12521=>"11111111",
  12522=>"00000010",
  12523=>"00000001",
  12524=>"11111111",
  12525=>"00000100",
  12526=>"11111101",
  12527=>"11111111",
  12528=>"11111111",
  12529=>"00000000",
  12530=>"00000001",
  12531=>"11111101",
  12532=>"00000100",
  12533=>"00000100",
  12534=>"11111101",
  12535=>"00000010",
  12536=>"11111110",
  12537=>"11111110",
  12538=>"00000010",
  12539=>"00000010",
  12540=>"00000001",
  12541=>"11111111",
  12542=>"00000001",
  12543=>"00000000",
  12544=>"11111111",
  12545=>"00000100",
  12546=>"00000000",
  12547=>"11111101",
  12548=>"00000000",
  12549=>"11111101",
  12550=>"00000100",
  12551=>"00000010",
  12552=>"11111110",
  12553=>"00000000",
  12554=>"11111111",
  12555=>"00000001",
  12556=>"11111110",
  12557=>"00000101",
  12558=>"11111101",
  12559=>"00000000",
  12560=>"11111110",
  12561=>"00000101",
  12562=>"00000101",
  12563=>"11111111",
  12564=>"00000011",
  12565=>"00000011",
  12566=>"00000010",
  12567=>"11111101",
  12568=>"11111110",
  12569=>"00000100",
  12570=>"00000100",
  12571=>"11111101",
  12572=>"11111110",
  12573=>"00000010",
  12574=>"00000001",
  12575=>"00000010",
  12576=>"11111110",
  12577=>"11111110",
  12578=>"00000001",
  12579=>"00000000",
  12580=>"11111111",
  12581=>"00000000",
  12582=>"11111111",
  12583=>"00000001",
  12584=>"11111101",
  12585=>"00000010",
  12586=>"11111110",
  12587=>"11111111",
  12588=>"11111111",
  12589=>"11111111",
  12590=>"11111111",
  12591=>"00000010",
  12592=>"00000000",
  12593=>"11111110",
  12594=>"11111101",
  12595=>"00000010",
  12596=>"11111110",
  12597=>"00000101",
  12598=>"11111101",
  12599=>"11111110",
  12600=>"00000010",
  12601=>"00000011",
  12602=>"11111111",
  12603=>"11111110",
  12604=>"00000010",
  12605=>"11111101",
  12606=>"00000001",
  12607=>"00000010",
  12608=>"11111110",
  12609=>"00000000",
  12610=>"00000000",
  12611=>"00000000",
  12612=>"11111101",
  12613=>"00000100",
  12614=>"11111110",
  12615=>"11111110",
  12616=>"00000001",
  12617=>"11111110",
  12618=>"00000010",
  12619=>"11111111",
  12620=>"00000100",
  12621=>"00000010",
  12622=>"11111110",
  12623=>"11111111",
  12624=>"11111101",
  12625=>"11111110",
  12626=>"11111101",
  12627=>"00000000",
  12628=>"11111110",
  12629=>"11111101",
  12630=>"00000001",
  12631=>"11111110",
  12632=>"11111101",
  12633=>"11111110",
  12634=>"11111110",
  12635=>"00000011",
  12636=>"11111110",
  12637=>"00000011",
  12638=>"00000011",
  12639=>"11111111",
  12640=>"11111111",
  12641=>"00000011",
  12642=>"00000010",
  12643=>"00000001",
  12644=>"00000001",
  12645=>"11111110",
  12646=>"00000010",
  12647=>"00000000",
  12648=>"00000000",
  12649=>"00000001",
  12650=>"00000010",
  12651=>"11111111",
  12652=>"11111111",
  12653=>"11111101",
  12654=>"00000001",
  12655=>"00000000",
  12656=>"00000000",
  12657=>"00000000",
  12658=>"00000001",
  12659=>"00000001",
  12660=>"11111111",
  12661=>"00000001",
  12662=>"00000100",
  12663=>"00000000",
  12664=>"11111111",
  12665=>"11111101",
  12666=>"11111110",
  12667=>"00000000",
  12668=>"11111110",
  12669=>"00000001",
  12670=>"00000001",
  12671=>"00000000",
  12672=>"00000011",
  12673=>"00000001",
  12674=>"11111110",
  12675=>"11111110",
  12676=>"00000001",
  12677=>"11111101",
  12678=>"00000010",
  12679=>"11111111",
  12680=>"00000000",
  12681=>"00000001",
  12682=>"00000001",
  12683=>"11111101",
  12684=>"00000001",
  12685=>"11111110",
  12686=>"00000010",
  12687=>"11111111",
  12688=>"00000001",
  12689=>"11111111",
  12690=>"00000101",
  12691=>"11111111",
  12692=>"00000000",
  12693=>"00000010",
  12694=>"00000010",
  12695=>"11111101",
  12696=>"11111111",
  12697=>"11111101",
  12698=>"00000011",
  12699=>"11111111",
  12700=>"00000000",
  12701=>"11111111",
  12702=>"00000011",
  12703=>"11111110",
  12704=>"11111101",
  12705=>"11111110",
  12706=>"11111111",
  12707=>"11111101",
  12708=>"11111110",
  12709=>"11111101",
  12710=>"11111111",
  12711=>"00000010",
  12712=>"00000001",
  12713=>"11111111",
  12714=>"00000011",
  12715=>"00000011",
  12716=>"11111111",
  12717=>"00000000",
  12718=>"00000001",
  12719=>"11111110",
  12720=>"11111101",
  12721=>"00000010",
  12722=>"11111111",
  12723=>"00000010",
  12724=>"00000011",
  12725=>"11111110",
  12726=>"00000100",
  12727=>"00000010",
  12728=>"00000000",
  12729=>"00000001",
  12730=>"11111100",
  12731=>"11111100",
  12732=>"00000001",
  12733=>"11111101",
  12734=>"11111101",
  12735=>"11111101",
  12736=>"11111110",
  12737=>"00000001",
  12738=>"11111101",
  12739=>"00000000",
  12740=>"00000010",
  12741=>"00000010",
  12742=>"11111111",
  12743=>"11111111",
  12744=>"00000100",
  12745=>"11111111",
  12746=>"00000010",
  12747=>"11111110",
  12748=>"00000010",
  12749=>"00000001",
  12750=>"00000000",
  12751=>"00000010",
  12752=>"00000000",
  12753=>"00000010",
  12754=>"00000001",
  12755=>"00000000",
  12756=>"11111111",
  12757=>"00000010",
  12758=>"11111100",
  12759=>"00000011",
  12760=>"00000011",
  12761=>"11111101",
  12762=>"00000001",
  12763=>"00000001",
  12764=>"11111111",
  12765=>"00000010",
  12766=>"00000011",
  12767=>"11111110",
  12768=>"00000000",
  12769=>"00000011",
  12770=>"00000100",
  12771=>"11111110",
  12772=>"11111111",
  12773=>"11111100",
  12774=>"11111111",
  12775=>"11111110",
  12776=>"00000000",
  12777=>"00000000",
  12778=>"11111111",
  12779=>"11111111",
  12780=>"11111110",
  12781=>"00000000",
  12782=>"11111111",
  12783=>"00000010",
  12784=>"11111111",
  12785=>"00000011",
  12786=>"11111101",
  12787=>"00000011",
  12788=>"00000000",
  12789=>"11111101",
  12790=>"00000000",
  12791=>"00000000",
  12792=>"00000000",
  12793=>"11111101",
  12794=>"11111110",
  12795=>"11111110",
  12796=>"11111110",
  12797=>"11111101",
  12798=>"00000000",
  12799=>"00000001",
  12800=>"11111110",
  12801=>"00000000",
  12802=>"00000011",
  12803=>"00000010",
  12804=>"11111110",
  12805=>"11111110",
  12806=>"00000011",
  12807=>"00000010",
  12808=>"00000001",
  12809=>"11111101",
  12810=>"11111110",
  12811=>"11111101",
  12812=>"00000010",
  12813=>"11111111",
  12814=>"00000100",
  12815=>"00000000",
  12816=>"11111111",
  12817=>"00000010",
  12818=>"11111110",
  12819=>"00000011",
  12820=>"11111101",
  12821=>"00000000",
  12822=>"00000000",
  12823=>"11111110",
  12824=>"00000000",
  12825=>"00000011",
  12826=>"11111111",
  12827=>"00000100",
  12828=>"11111101",
  12829=>"11111100",
  12830=>"11111111",
  12831=>"00000000",
  12832=>"11111111",
  12833=>"11111110",
  12834=>"11111101",
  12835=>"00000001",
  12836=>"11111111",
  12837=>"11111101",
  12838=>"00000000",
  12839=>"11111110",
  12840=>"11111110",
  12841=>"00000000",
  12842=>"11111111",
  12843=>"11111110",
  12844=>"11111101",
  12845=>"00000000",
  12846=>"00000001",
  12847=>"00000000",
  12848=>"11111110",
  12849=>"00000001",
  12850=>"00000000",
  12851=>"11111110",
  12852=>"11111110",
  12853=>"00000010",
  12854=>"00000001",
  12855=>"00000010",
  12856=>"00000011",
  12857=>"00000010",
  12858=>"00000001",
  12859=>"00000010",
  12860=>"00000010",
  12861=>"11111110",
  12862=>"11111101",
  12863=>"11111111",
  12864=>"11111111",
  12865=>"00000010",
  12866=>"00000011",
  12867=>"00000010",
  12868=>"00000001",
  12869=>"11111111",
  12870=>"11111110",
  12871=>"00000001",
  12872=>"00000010",
  12873=>"11111110",
  12874=>"00000011",
  12875=>"00000010",
  12876=>"00000100",
  12877=>"00000000",
  12878=>"00000000",
  12879=>"00000010",
  12880=>"11111110",
  12881=>"00000101",
  12882=>"00000011",
  12883=>"11111111",
  12884=>"00000001",
  12885=>"11111110",
  12886=>"11111111",
  12887=>"00000001",
  12888=>"00000000",
  12889=>"00000011",
  12890=>"00000000",
  12891=>"11111110",
  12892=>"11111101",
  12893=>"00000001",
  12894=>"00000001",
  12895=>"00000000",
  12896=>"11111111",
  12897=>"11111111",
  12898=>"11111111",
  12899=>"00000101",
  12900=>"00000000",
  12901=>"00000001",
  12902=>"00000010",
  12903=>"00000000",
  12904=>"00000101",
  12905=>"00000010",
  12906=>"11111111",
  12907=>"11111111",
  12908=>"11111110",
  12909=>"00000011",
  12910=>"11111110",
  12911=>"11111110",
  12912=>"00000000",
  12913=>"11111101",
  12914=>"00000000",
  12915=>"11111111",
  12916=>"00000000",
  12917=>"00000001",
  12918=>"00000001",
  12919=>"00000100",
  12920=>"00000010",
  12921=>"00000000",
  12922=>"11111100",
  12923=>"00000010",
  12924=>"11111110",
  12925=>"11111111",
  12926=>"00000010",
  12927=>"00000000",
  12928=>"00000010",
  12929=>"00000011",
  12930=>"00000001",
  12931=>"11111110",
  12932=>"11111110",
  12933=>"00000000",
  12934=>"00000000",
  12935=>"11111100",
  12936=>"11111110",
  12937=>"11111101",
  12938=>"00000001",
  12939=>"00000000",
  12940=>"00000000",
  12941=>"00000010",
  12942=>"00000001",
  12943=>"11111110",
  12944=>"00000010",
  12945=>"11111111",
  12946=>"00000001",
  12947=>"11111111",
  12948=>"11111111",
  12949=>"00000000",
  12950=>"11111111",
  12951=>"00000101",
  12952=>"00000011",
  12953=>"11111101",
  12954=>"00000011",
  12955=>"11111101",
  12956=>"00000011",
  12957=>"00000001",
  12958=>"00000001",
  12959=>"11111110",
  12960=>"11111110",
  12961=>"11111111",
  12962=>"00000000",
  12963=>"00000000",
  12964=>"11111111",
  12965=>"11111111",
  12966=>"00000001",
  12967=>"00000010",
  12968=>"11111110",
  12969=>"11111110",
  12970=>"11111110",
  12971=>"11111111",
  12972=>"11111101",
  12973=>"00000101",
  12974=>"00000000",
  12975=>"11111101",
  12976=>"00000000",
  12977=>"11111100",
  12978=>"11111111",
  12979=>"00000000",
  12980=>"00000000",
  12981=>"00000011",
  12982=>"00000000",
  12983=>"11111111",
  12984=>"00000011",
  12985=>"11111111",
  12986=>"11111111",
  12987=>"00000000",
  12988=>"00000011",
  12989=>"00000100",
  12990=>"00000100",
  12991=>"11111110",
  12992=>"11111101",
  12993=>"00000001",
  12994=>"00000001",
  12995=>"11111111",
  12996=>"00000010",
  12997=>"00000001",
  12998=>"11111111",
  12999=>"11111110",
  13000=>"00000001",
  13001=>"00000000",
  13002=>"00000000",
  13003=>"00000010",
  13004=>"11111111",
  13005=>"00000100",
  13006=>"00000011",
  13007=>"00000010",
  13008=>"00000010",
  13009=>"00000000",
  13010=>"00000000",
  13011=>"00000011",
  13012=>"11111110",
  13013=>"11111101",
  13014=>"00000010",
  13015=>"11111110",
  13016=>"00000000",
  13017=>"00000000",
  13018=>"00000001",
  13019=>"11111111",
  13020=>"00000000",
  13021=>"00000000",
  13022=>"00000000",
  13023=>"00000000",
  13024=>"11111110",
  13025=>"11111111",
  13026=>"11111101",
  13027=>"11111111",
  13028=>"00000010",
  13029=>"11111111",
  13030=>"00000010",
  13031=>"00000000",
  13032=>"00000010",
  13033=>"11111101",
  13034=>"11111111",
  13035=>"11111111",
  13036=>"00000010",
  13037=>"11111110",
  13038=>"11111111",
  13039=>"00000011",
  13040=>"00000010",
  13041=>"00000001",
  13042=>"00000000",
  13043=>"00000010",
  13044=>"00000011",
  13045=>"00000000",
  13046=>"11111101",
  13047=>"11111101",
  13048=>"00000010",
  13049=>"00000001",
  13050=>"00000001",
  13051=>"11111110",
  13052=>"11111111",
  13053=>"11111101",
  13054=>"00000110",
  13055=>"00000000",
  13056=>"00000000",
  13057=>"00000011",
  13058=>"00000011",
  13059=>"11111110",
  13060=>"11111111",
  13061=>"11111111",
  13062=>"00000010",
  13063=>"11111110",
  13064=>"00000000",
  13065=>"11111110",
  13066=>"00000001",
  13067=>"11111111",
  13068=>"00000001",
  13069=>"00000010",
  13070=>"11111110",
  13071=>"11111110",
  13072=>"00000000",
  13073=>"00000000",
  13074=>"11111111",
  13075=>"00000100",
  13076=>"00000010",
  13077=>"11111111",
  13078=>"00000000",
  13079=>"00000011",
  13080=>"11111101",
  13081=>"00000011",
  13082=>"11111110",
  13083=>"00000001",
  13084=>"11111101",
  13085=>"00000001",
  13086=>"00000100",
  13087=>"00000001",
  13088=>"00000000",
  13089=>"00000001",
  13090=>"00000011",
  13091=>"00000011",
  13092=>"11111110",
  13093=>"00000001",
  13094=>"11111101",
  13095=>"00000000",
  13096=>"00000101",
  13097=>"11111111",
  13098=>"00000010",
  13099=>"11111111",
  13100=>"11111110",
  13101=>"00000001",
  13102=>"00000001",
  13103=>"00000001",
  13104=>"11111111",
  13105=>"11111100",
  13106=>"00000000",
  13107=>"11111111",
  13108=>"00000000",
  13109=>"00000001",
  13110=>"11111110",
  13111=>"00000001",
  13112=>"00000000",
  13113=>"11111110",
  13114=>"00000001",
  13115=>"00000011",
  13116=>"00000001",
  13117=>"00000010",
  13118=>"11111110",
  13119=>"00000001",
  13120=>"11111111",
  13121=>"11111110",
  13122=>"11111111",
  13123=>"00000000",
  13124=>"11111101",
  13125=>"00000000",
  13126=>"00000011",
  13127=>"11111101",
  13128=>"11111111",
  13129=>"00000000",
  13130=>"00000000",
  13131=>"11111111",
  13132=>"11111111",
  13133=>"11111110",
  13134=>"11111100",
  13135=>"00000001",
  13136=>"11111111",
  13137=>"00000000",
  13138=>"11111101",
  13139=>"00000000",
  13140=>"00000000",
  13141=>"11111110",
  13142=>"11111101",
  13143=>"11111111",
  13144=>"11111110",
  13145=>"00000010",
  13146=>"00000001",
  13147=>"11111110",
  13148=>"00000000",
  13149=>"11111111",
  13150=>"00000010",
  13151=>"11111101",
  13152=>"00000000",
  13153=>"11111110",
  13154=>"00000010",
  13155=>"11111110",
  13156=>"00000011",
  13157=>"00000000",
  13158=>"11111111",
  13159=>"11111101",
  13160=>"11111101",
  13161=>"00000001",
  13162=>"11111111",
  13163=>"00000001",
  13164=>"11111110",
  13165=>"00000000",
  13166=>"11111111",
  13167=>"00000000",
  13168=>"11111110",
  13169=>"00000000",
  13170=>"11111110",
  13171=>"00000000",
  13172=>"00000000",
  13173=>"11111111",
  13174=>"00000001",
  13175=>"00000001",
  13176=>"11111100",
  13177=>"11111111",
  13178=>"11111110",
  13179=>"00000010",
  13180=>"11111110",
  13181=>"11111101",
  13182=>"00000000",
  13183=>"00000001",
  13184=>"00000000",
  13185=>"11111111",
  13186=>"11111110",
  13187=>"00000000",
  13188=>"00000001",
  13189=>"00000001",
  13190=>"11111111",
  13191=>"00000011",
  13192=>"00000010",
  13193=>"11111101",
  13194=>"00000000",
  13195=>"00000010",
  13196=>"11111111",
  13197=>"00000011",
  13198=>"11111110",
  13199=>"00000010",
  13200=>"11111110",
  13201=>"00000000",
  13202=>"11111111",
  13203=>"00000001",
  13204=>"00000001",
  13205=>"00000100",
  13206=>"00000000",
  13207=>"00000001",
  13208=>"11111110",
  13209=>"00000001",
  13210=>"11111111",
  13211=>"00000010",
  13212=>"00000011",
  13213=>"00000010",
  13214=>"11111111",
  13215=>"00000000",
  13216=>"11111110",
  13217=>"11111111",
  13218=>"00000100",
  13219=>"00000011",
  13220=>"11111110",
  13221=>"11111111",
  13222=>"00000100",
  13223=>"00000001",
  13224=>"00000000",
  13225=>"00000000",
  13226=>"00000000",
  13227=>"11111110",
  13228=>"11111111",
  13229=>"00000010",
  13230=>"00000010",
  13231=>"11111111",
  13232=>"11111111",
  13233=>"00000011",
  13234=>"11111101",
  13235=>"11111110",
  13236=>"00000001",
  13237=>"00000011",
  13238=>"00000010",
  13239=>"11111110",
  13240=>"00000000",
  13241=>"11111101",
  13242=>"00000010",
  13243=>"11111110",
  13244=>"11111101",
  13245=>"11111110",
  13246=>"00000001",
  13247=>"11111110",
  13248=>"00000000",
  13249=>"00000000",
  13250=>"11111110",
  13251=>"00000000",
  13252=>"11111101",
  13253=>"11111101",
  13254=>"11111110",
  13255=>"00000000",
  13256=>"00000010",
  13257=>"00000000",
  13258=>"00000000",
  13259=>"00000010",
  13260=>"00000000",
  13261=>"11111110",
  13262=>"00000000",
  13263=>"00000100",
  13264=>"11111110",
  13265=>"00000000",
  13266=>"00000100",
  13267=>"11111101",
  13268=>"11111101",
  13269=>"00000010",
  13270=>"11111111",
  13271=>"00000000",
  13272=>"00000010",
  13273=>"11111101",
  13274=>"00000001",
  13275=>"11111100",
  13276=>"11111101",
  13277=>"00000000",
  13278=>"11111110",
  13279=>"00000000",
  13280=>"11111101",
  13281=>"11111110",
  13282=>"11111110",
  13283=>"11111101",
  13284=>"11111111",
  13285=>"11111111",
  13286=>"00000000",
  13287=>"00000011",
  13288=>"11111110",
  13289=>"11111110",
  13290=>"00000000",
  13291=>"00000100",
  13292=>"00000000",
  13293=>"11111110",
  13294=>"00000010",
  13295=>"00000011",
  13296=>"00000001",
  13297=>"00000001",
  13298=>"11111100",
  13299=>"00000101",
  13300=>"11111111",
  13301=>"00000000",
  13302=>"00000000",
  13303=>"00000000",
  13304=>"11111111",
  13305=>"11111111",
  13306=>"00000000",
  13307=>"00000000",
  13308=>"00000100",
  13309=>"00000001",
  13310=>"11111101",
  13311=>"11111101",
  13312=>"11111111",
  13313=>"00000010",
  13314=>"11111101",
  13315=>"11111111",
  13316=>"00000010",
  13317=>"00000001",
  13318=>"00000000",
  13319=>"11111101",
  13320=>"00000001",
  13321=>"11111101",
  13322=>"00000010",
  13323=>"00000000",
  13324=>"11111111",
  13325=>"00000000",
  13326=>"00000001",
  13327=>"11111101",
  13328=>"11111101",
  13329=>"11111111",
  13330=>"00000010",
  13331=>"00000000",
  13332=>"00000100",
  13333=>"11111111",
  13334=>"11111110",
  13335=>"11111110",
  13336=>"00000100",
  13337=>"00000010",
  13338=>"00000101",
  13339=>"00000010",
  13340=>"11111111",
  13341=>"00000110",
  13342=>"00000101",
  13343=>"11111111",
  13344=>"11111111",
  13345=>"11111101",
  13346=>"00000111",
  13347=>"11111111",
  13348=>"00000011",
  13349=>"11111110",
  13350=>"11111110",
  13351=>"00000000",
  13352=>"00000000",
  13353=>"11111100",
  13354=>"11111110",
  13355=>"00000101",
  13356=>"00000001",
  13357=>"00000000",
  13358=>"11111101",
  13359=>"00000010",
  13360=>"11111110",
  13361=>"11111100",
  13362=>"00000001",
  13363=>"00000100",
  13364=>"00000000",
  13365=>"00000000",
  13366=>"11111101",
  13367=>"11111110",
  13368=>"11111110",
  13369=>"00000011",
  13370=>"00000001",
  13371=>"00000001",
  13372=>"00000010",
  13373=>"11111110",
  13374=>"00000100",
  13375=>"11111110",
  13376=>"11111111",
  13377=>"00000001",
  13378=>"00000000",
  13379=>"11111101",
  13380=>"11111110",
  13381=>"00000001",
  13382=>"00000100",
  13383=>"00000000",
  13384=>"00000010",
  13385=>"11111101",
  13386=>"00000100",
  13387=>"11111101",
  13388=>"00000010",
  13389=>"00000010",
  13390=>"00000010",
  13391=>"00000100",
  13392=>"00000000",
  13393=>"11111110",
  13394=>"00000010",
  13395=>"00000000",
  13396=>"00000011",
  13397=>"11111101",
  13398=>"00000001",
  13399=>"11111111",
  13400=>"11111111",
  13401=>"11111011",
  13402=>"00000011",
  13403=>"11111101",
  13404=>"00000001",
  13405=>"00000000",
  13406=>"11111110",
  13407=>"00000011",
  13408=>"00000000",
  13409=>"00000001",
  13410=>"00000010",
  13411=>"11111111",
  13412=>"11111110",
  13413=>"11111111",
  13414=>"11111111",
  13415=>"00000010",
  13416=>"00000011",
  13417=>"00000100",
  13418=>"00000011",
  13419=>"11111101",
  13420=>"00000001",
  13421=>"00000010",
  13422=>"11111111",
  13423=>"11111101",
  13424=>"11111101",
  13425=>"00000000",
  13426=>"00000010",
  13427=>"11111101",
  13428=>"00000001",
  13429=>"11111111",
  13430=>"11111110",
  13431=>"00000001",
  13432=>"11111110",
  13433=>"11111111",
  13434=>"00000011",
  13435=>"00000000",
  13436=>"00000010",
  13437=>"11111011",
  13438=>"11111101",
  13439=>"11111110",
  13440=>"00000001",
  13441=>"00000001",
  13442=>"11111100",
  13443=>"00000101",
  13444=>"11111100",
  13445=>"00000001",
  13446=>"00000000",
  13447=>"00000011",
  13448=>"11111100",
  13449=>"11111111",
  13450=>"11111110",
  13451=>"00000000",
  13452=>"11111110",
  13453=>"00000001",
  13454=>"00000010",
  13455=>"11111111",
  13456=>"00000000",
  13457=>"11111110",
  13458=>"11111111",
  13459=>"11111110",
  13460=>"11111111",
  13461=>"00000011",
  13462=>"11111110",
  13463=>"00000001",
  13464=>"00000100",
  13465=>"00000001",
  13466=>"11111111",
  13467=>"00000010",
  13468=>"00000001",
  13469=>"11111101",
  13470=>"11111110",
  13471=>"00000011",
  13472=>"00000101",
  13473=>"11111110",
  13474=>"00000000",
  13475=>"00000011",
  13476=>"11111111",
  13477=>"11111100",
  13478=>"00000001",
  13479=>"00000000",
  13480=>"00000001",
  13481=>"00000000",
  13482=>"11111111",
  13483=>"00000001",
  13484=>"00000000",
  13485=>"11111101",
  13486=>"00000011",
  13487=>"00000010",
  13488=>"00000001",
  13489=>"00000000",
  13490=>"11111110",
  13491=>"11111111",
  13492=>"11111101",
  13493=>"11111110",
  13494=>"11111100",
  13495=>"00000100",
  13496=>"11111110",
  13497=>"00000000",
  13498=>"00000000",
  13499=>"11111111",
  13500=>"11111111",
  13501=>"00000011",
  13502=>"00000110",
  13503=>"11111110",
  13504=>"00000011",
  13505=>"11111111",
  13506=>"11111111",
  13507=>"11111110",
  13508=>"11111111",
  13509=>"00000001",
  13510=>"00000100",
  13511=>"00000010",
  13512=>"11111111",
  13513=>"11111101",
  13514=>"00000000",
  13515=>"00000000",
  13516=>"00000000",
  13517=>"00000000",
  13518=>"00000010",
  13519=>"11111100",
  13520=>"00000010",
  13521=>"00000100",
  13522=>"11111111",
  13523=>"00000000",
  13524=>"11111111",
  13525=>"00000000",
  13526=>"00000001",
  13527=>"00000000",
  13528=>"00000001",
  13529=>"11111101",
  13530=>"00000001",
  13531=>"11111011",
  13532=>"00000010",
  13533=>"00000000",
  13534=>"11111101",
  13535=>"00000100",
  13536=>"11111111",
  13537=>"00000000",
  13538=>"11111110",
  13539=>"00000011",
  13540=>"11111101",
  13541=>"11111111",
  13542=>"00000000",
  13543=>"00000110",
  13544=>"11111111",
  13545=>"00000010",
  13546=>"00000000",
  13547=>"00000010",
  13548=>"11111111",
  13549=>"11111100",
  13550=>"00000100",
  13551=>"00000010",
  13552=>"11111111",
  13553=>"11111111",
  13554=>"00000001",
  13555=>"00000010",
  13556=>"11111111",
  13557=>"11111101",
  13558=>"00000100",
  13559=>"11111111",
  13560=>"11111101",
  13561=>"00000011",
  13562=>"00000001",
  13563=>"11111101",
  13564=>"11111110",
  13565=>"00000010",
  13566=>"00000100",
  13567=>"00000101",
  13568=>"11111101",
  13569=>"11111101",
  13570=>"00000001",
  13571=>"00000010",
  13572=>"11111111",
  13573=>"11111101",
  13574=>"00000010",
  13575=>"00000011",
  13576=>"11111100",
  13577=>"00000100",
  13578=>"11111110",
  13579=>"11111111",
  13580=>"11111110",
  13581=>"11111111",
  13582=>"11111111",
  13583=>"11111101",
  13584=>"00000100",
  13585=>"00000100",
  13586=>"11111110",
  13587=>"00000000",
  13588=>"00000100",
  13589=>"00000000",
  13590=>"00000111",
  13591=>"11111111",
  13592=>"11111111",
  13593=>"00000000",
  13594=>"11111101",
  13595=>"11111101",
  13596=>"11111110",
  13597=>"11111101",
  13598=>"00000001",
  13599=>"11111101",
  13600=>"11111111",
  13601=>"00000000",
  13602=>"00000001",
  13603=>"00000000",
  13604=>"00000000",
  13605=>"11111110",
  13606=>"11111111",
  13607=>"00000011",
  13608=>"11111011",
  13609=>"00000100",
  13610=>"11111101",
  13611=>"11111101",
  13612=>"00000010",
  13613=>"11111111",
  13614=>"11111110",
  13615=>"00000000",
  13616=>"11111110",
  13617=>"00000001",
  13618=>"11111101",
  13619=>"11111110",
  13620=>"00000011",
  13621=>"11111101",
  13622=>"11111101",
  13623=>"11111100",
  13624=>"00000000",
  13625=>"11111111",
  13626=>"11111110",
  13627=>"00000000",
  13628=>"00000000",
  13629=>"00000110",
  13630=>"00000010",
  13631=>"00000001",
  13632=>"11111111",
  13633=>"11111111",
  13634=>"11111111",
  13635=>"00000101",
  13636=>"00000010",
  13637=>"00000000",
  13638=>"00000011",
  13639=>"00000000",
  13640=>"00000010",
  13641=>"00000100",
  13642=>"00000010",
  13643=>"11111110",
  13644=>"11111010",
  13645=>"00000001",
  13646=>"00000010",
  13647=>"11111111",
  13648=>"11111110",
  13649=>"00000001",
  13650=>"11111111",
  13651=>"11111110",
  13652=>"00000100",
  13653=>"00000000",
  13654=>"11111101",
  13655=>"11111111",
  13656=>"00000100",
  13657=>"11111101",
  13658=>"00000100",
  13659=>"11111111",
  13660=>"11111110",
  13661=>"00000000",
  13662=>"00000011",
  13663=>"00000001",
  13664=>"00000100",
  13665=>"11111110",
  13666=>"11111111",
  13667=>"00000000",
  13668=>"00000010",
  13669=>"11111110",
  13670=>"00000100",
  13671=>"00000001",
  13672=>"00000010",
  13673=>"00000000",
  13674=>"00000001",
  13675=>"00000011",
  13676=>"11111101",
  13677=>"11111110",
  13678=>"00000100",
  13679=>"00000000",
  13680=>"11111110",
  13681=>"00000010",
  13682=>"00000010",
  13683=>"11111110",
  13684=>"00000101",
  13685=>"00000100",
  13686=>"11111111",
  13687=>"00000010",
  13688=>"11111110",
  13689=>"00000001",
  13690=>"11111111",
  13691=>"00000000",
  13692=>"00000100",
  13693=>"11111110",
  13694=>"11111100",
  13695=>"00000100",
  13696=>"00000000",
  13697=>"00000000",
  13698=>"00000000",
  13699=>"00000001",
  13700=>"00000000",
  13701=>"11111111",
  13702=>"00000100",
  13703=>"11111110",
  13704=>"00000100",
  13705=>"11111111",
  13706=>"00000000",
  13707=>"11111100",
  13708=>"00000011",
  13709=>"00000011",
  13710=>"11111101",
  13711=>"11111100",
  13712=>"11111110",
  13713=>"00000000",
  13714=>"11111101",
  13715=>"11111101",
  13716=>"11111101",
  13717=>"00000100",
  13718=>"11111101",
  13719=>"11111110",
  13720=>"00000001",
  13721=>"11111110",
  13722=>"00000100",
  13723=>"11111100",
  13724=>"00000010",
  13725=>"00000001",
  13726=>"00000101",
  13727=>"11111100",
  13728=>"11111111",
  13729=>"11111110",
  13730=>"00000000",
  13731=>"00000000",
  13732=>"00000001",
  13733=>"11111011",
  13734=>"00000001",
  13735=>"00000000",
  13736=>"00000010",
  13737=>"00000000",
  13738=>"00000000",
  13739=>"11111110",
  13740=>"11111101",
  13741=>"11111101",
  13742=>"11111111",
  13743=>"00000011",
  13744=>"11111111",
  13745=>"00000000",
  13746=>"00000011",
  13747=>"11111111",
  13748=>"00000010",
  13749=>"00000100",
  13750=>"11111111",
  13751=>"00000010",
  13752=>"11111101",
  13753=>"11111101",
  13754=>"00000001",
  13755=>"00000010",
  13756=>"00000010",
  13757=>"00000001",
  13758=>"00000000",
  13759=>"11111101",
  13760=>"00000101",
  13761=>"11111100",
  13762=>"00000100",
  13763=>"11111111",
  13764=>"11111110",
  13765=>"00000010",
  13766=>"00000100",
  13767=>"00000101",
  13768=>"11111101",
  13769=>"00000000",
  13770=>"11111110",
  13771=>"00000001",
  13772=>"00000001",
  13773=>"00000001",
  13774=>"11111110",
  13775=>"00000000",
  13776=>"11111111",
  13777=>"11111101",
  13778=>"11111110",
  13779=>"00000010",
  13780=>"11111101",
  13781=>"00000000",
  13782=>"11111110",
  13783=>"11111110",
  13784=>"00000010",
  13785=>"00000110",
  13786=>"00000011",
  13787=>"00000001",
  13788=>"00000001",
  13789=>"00000010",
  13790=>"00000000",
  13791=>"11111111",
  13792=>"00000011",
  13793=>"00000011",
  13794=>"00000010",
  13795=>"11111101",
  13796=>"11111110",
  13797=>"11111111",
  13798=>"00000101",
  13799=>"11111111",
  13800=>"11111110",
  13801=>"11111101",
  13802=>"11111100",
  13803=>"00000001",
  13804=>"00000001",
  13805=>"11111111",
  13806=>"11111110",
  13807=>"00000101",
  13808=>"00000000",
  13809=>"00000000",
  13810=>"00000001",
  13811=>"00000000",
  13812=>"11111101",
  13813=>"00000010",
  13814=>"00000011",
  13815=>"00000001",
  13816=>"00000000",
  13817=>"00000010",
  13818=>"00000001",
  13819=>"11111011",
  13820=>"00000000",
  13821=>"11111111",
  13822=>"11111110",
  13823=>"11111101",
  13824=>"00000011",
  13825=>"11111111",
  13826=>"11111111",
  13827=>"11111010",
  13828=>"11111010",
  13829=>"00000010",
  13830=>"11111110",
  13831=>"11111110",
  13832=>"11111110",
  13833=>"00000011",
  13834=>"00000010",
  13835=>"00000001",
  13836=>"11111100",
  13837=>"00000000",
  13838=>"00000010",
  13839=>"11111111",
  13840=>"00000001",
  13841=>"11111011",
  13842=>"11111110",
  13843=>"00000100",
  13844=>"00000100",
  13845=>"00000010",
  13846=>"00000100",
  13847=>"00000011",
  13848=>"00000001",
  13849=>"00000001",
  13850=>"00000001",
  13851=>"00000010",
  13852=>"00000010",
  13853=>"00000100",
  13854=>"11111110",
  13855=>"00000100",
  13856=>"11111111",
  13857=>"00000000",
  13858=>"11111110",
  13859=>"11111110",
  13860=>"11111110",
  13861=>"00000000",
  13862=>"00000000",
  13863=>"11111111",
  13864=>"00000000",
  13865=>"00000000",
  13866=>"11111100",
  13867=>"11111101",
  13868=>"00000111",
  13869=>"00000010",
  13870=>"00000000",
  13871=>"00000101",
  13872=>"00000101",
  13873=>"00000001",
  13874=>"00000010",
  13875=>"00000001",
  13876=>"00000001",
  13877=>"00000011",
  13878=>"11111101",
  13879=>"11111101",
  13880=>"11111111",
  13881=>"00000011",
  13882=>"11111101",
  13883=>"11111110",
  13884=>"00000001",
  13885=>"11111111",
  13886=>"00000100",
  13887=>"00000100",
  13888=>"00000000",
  13889=>"11111011",
  13890=>"00000100",
  13891=>"11111111",
  13892=>"00000001",
  13893=>"00000000",
  13894=>"11111101",
  13895=>"00000010",
  13896=>"11111101",
  13897=>"11111101",
  13898=>"00000001",
  13899=>"00000011",
  13900=>"00000001",
  13901=>"00000010",
  13902=>"00000100",
  13903=>"00000010",
  13904=>"00000011",
  13905=>"00000010",
  13906=>"11111111",
  13907=>"00000011",
  13908=>"11111101",
  13909=>"00000100",
  13910=>"11111101",
  13911=>"00000000",
  13912=>"11111111",
  13913=>"11111111",
  13914=>"00000010",
  13915=>"00000101",
  13916=>"00000000",
  13917=>"00000000",
  13918=>"00000010",
  13919=>"00000001",
  13920=>"00000010",
  13921=>"00000010",
  13922=>"00000000",
  13923=>"11111011",
  13924=>"11111101",
  13925=>"00000001",
  13926=>"00000010",
  13927=>"11111110",
  13928=>"00000001",
  13929=>"00000001",
  13930=>"11111110",
  13931=>"00000001",
  13932=>"11111110",
  13933=>"00000010",
  13934=>"00000000",
  13935=>"00000000",
  13936=>"00000000",
  13937=>"00000010",
  13938=>"00000010",
  13939=>"00000100",
  13940=>"11111111",
  13941=>"00000011",
  13942=>"11111111",
  13943=>"00000100",
  13944=>"00000010",
  13945=>"00000010",
  13946=>"00000010",
  13947=>"00000000",
  13948=>"00000000",
  13949=>"11111111",
  13950=>"11111100",
  13951=>"00000011",
  13952=>"11111110",
  13953=>"00000001",
  13954=>"11111110",
  13955=>"11111111",
  13956=>"11111111",
  13957=>"00000010",
  13958=>"00000011",
  13959=>"11111001",
  13960=>"00000100",
  13961=>"00000010",
  13962=>"00000010",
  13963=>"11111110",
  13964=>"00000001",
  13965=>"00000011",
  13966=>"00000010",
  13967=>"11111110",
  13968=>"00000010",
  13969=>"00000000",
  13970=>"11111101",
  13971=>"11111110",
  13972=>"11111111",
  13973=>"00000011",
  13974=>"11111101",
  13975=>"11111110",
  13976=>"11111100",
  13977=>"00000110",
  13978=>"11111111",
  13979=>"00000000",
  13980=>"11111101",
  13981=>"00000001",
  13982=>"11111111",
  13983=>"00000001",
  13984=>"11111111",
  13985=>"00000000",
  13986=>"00000100",
  13987=>"00000000",
  13988=>"00000000",
  13989=>"00000001",
  13990=>"00000001",
  13991=>"00000001",
  13992=>"11111101",
  13993=>"11111101",
  13994=>"00000000",
  13995=>"00000010",
  13996=>"00000010",
  13997=>"11111101",
  13998=>"11111101",
  13999=>"11111111",
  14000=>"00000001",
  14001=>"11111100",
  14002=>"00000011",
  14003=>"00000101",
  14004=>"00000000",
  14005=>"00000010",
  14006=>"11111110",
  14007=>"00000010",
  14008=>"00000000",
  14009=>"00000010",
  14010=>"11111111",
  14011=>"00000011",
  14012=>"11111111",
  14013=>"00000010",
  14014=>"00000001",
  14015=>"00000010",
  14016=>"00000001",
  14017=>"11111110",
  14018=>"11111110",
  14019=>"11111100",
  14020=>"00000010",
  14021=>"00000010",
  14022=>"11111111",
  14023=>"00000100",
  14024=>"00000100",
  14025=>"00000011",
  14026=>"00000010",
  14027=>"00000011",
  14028=>"00000011",
  14029=>"00000000",
  14030=>"00000000",
  14031=>"00000001",
  14032=>"00000001",
  14033=>"11111100",
  14034=>"00000010",
  14035=>"11111101",
  14036=>"00000010",
  14037=>"00000001",
  14038=>"00000010",
  14039=>"00000000",
  14040=>"00000001",
  14041=>"00000010",
  14042=>"11111111",
  14043=>"11111011",
  14044=>"00000011",
  14045=>"00000001",
  14046=>"00000001",
  14047=>"11111111",
  14048=>"00000101",
  14049=>"00000100",
  14050=>"11111111",
  14051=>"00000000",
  14052=>"00000010",
  14053=>"00000001",
  14054=>"00000000",
  14055=>"00000010",
  14056=>"00000001",
  14057=>"00000011",
  14058=>"11111110",
  14059=>"11111110",
  14060=>"11111111",
  14061=>"00000100",
  14062=>"11111110",
  14063=>"11111110",
  14064=>"00001000",
  14065=>"00000001",
  14066=>"11111110",
  14067=>"00000001",
  14068=>"00000000",
  14069=>"11111100",
  14070=>"11111111",
  14071=>"11111110",
  14072=>"00000110",
  14073=>"11111111",
  14074=>"11111110",
  14075=>"00000011",
  14076=>"11111101",
  14077=>"00000011",
  14078=>"00000001",
  14079=>"00000011",
  14080=>"00000110",
  14081=>"11111111",
  14082=>"00000010",
  14083=>"00000010",
  14084=>"11111111",
  14085=>"00000001",
  14086=>"11111101",
  14087=>"00000100",
  14088=>"00000000",
  14089=>"00000010",
  14090=>"11111111",
  14091=>"11111101",
  14092=>"00000001",
  14093=>"11111110",
  14094=>"11111110",
  14095=>"00000000",
  14096=>"00000000",
  14097=>"00000001",
  14098=>"11111101",
  14099=>"00000010",
  14100=>"00000001",
  14101=>"00000000",
  14102=>"00000011",
  14103=>"00000000",
  14104=>"00000011",
  14105=>"11111111",
  14106=>"11111111",
  14107=>"00000111",
  14108=>"11111110",
  14109=>"00000000",
  14110=>"00000010",
  14111=>"11111101",
  14112=>"00000011",
  14113=>"11111101",
  14114=>"00000001",
  14115=>"00000000",
  14116=>"11111110",
  14117=>"11111100",
  14118=>"11111111",
  14119=>"00000010",
  14120=>"00000100",
  14121=>"00000011",
  14122=>"00000010",
  14123=>"11111111",
  14124=>"00000010",
  14125=>"11111101",
  14126=>"00000100",
  14127=>"11111101",
  14128=>"11111111",
  14129=>"00000110",
  14130=>"00000011",
  14131=>"11111110",
  14132=>"11111110",
  14133=>"00000011",
  14134=>"00000011",
  14135=>"11111100",
  14136=>"00000010",
  14137=>"11111100",
  14138=>"11111101",
  14139=>"11111101",
  14140=>"11111110",
  14141=>"00000010",
  14142=>"11111101",
  14143=>"00000100",
  14144=>"11111101",
  14145=>"00000010",
  14146=>"00000000",
  14147=>"00000000",
  14148=>"00000100",
  14149=>"00000011",
  14150=>"11111111",
  14151=>"00000011",
  14152=>"11111111",
  14153=>"00000010",
  14154=>"11111101",
  14155=>"11111101",
  14156=>"00000100",
  14157=>"00000100",
  14158=>"11111111",
  14159=>"00000011",
  14160=>"00000010",
  14161=>"00000010",
  14162=>"00000001",
  14163=>"11111110",
  14164=>"00000010",
  14165=>"11111111",
  14166=>"00000000",
  14167=>"11111111",
  14168=>"00000100",
  14169=>"11111111",
  14170=>"00000000",
  14171=>"11111100",
  14172=>"00000000",
  14173=>"00000001",
  14174=>"00000110",
  14175=>"00000100",
  14176=>"00000010",
  14177=>"11111110",
  14178=>"11111101",
  14179=>"00000101",
  14180=>"11111101",
  14181=>"11111111",
  14182=>"11111110",
  14183=>"11111110",
  14184=>"11111100",
  14185=>"00000000",
  14186=>"00000010",
  14187=>"11111100",
  14188=>"11111101",
  14189=>"00000001",
  14190=>"00000010",
  14191=>"00000101",
  14192=>"00000010",
  14193=>"00000010",
  14194=>"11111110",
  14195=>"11111111",
  14196=>"11111110",
  14197=>"00000001",
  14198=>"00000011",
  14199=>"00000011",
  14200=>"00000010",
  14201=>"00000001",
  14202=>"11111110",
  14203=>"11111111",
  14204=>"11111111",
  14205=>"00000101",
  14206=>"00000011",
  14207=>"00000100",
  14208=>"11111110",
  14209=>"00000100",
  14210=>"00000001",
  14211=>"00000000",
  14212=>"11111100",
  14213=>"00000100",
  14214=>"00000010",
  14215=>"00000000",
  14216=>"11111101",
  14217=>"11111110",
  14218=>"00000000",
  14219=>"00000000",
  14220=>"11111101",
  14221=>"11111101",
  14222=>"00000000",
  14223=>"00000101",
  14224=>"00000001",
  14225=>"00000011",
  14226=>"00000011",
  14227=>"00000001",
  14228=>"00000010",
  14229=>"00000000",
  14230=>"00000011",
  14231=>"00000011",
  14232=>"00000011",
  14233=>"00000001",
  14234=>"00000100",
  14235=>"11111110",
  14236=>"00000010",
  14237=>"00000011",
  14238=>"11111101",
  14239=>"00000101",
  14240=>"00000001",
  14241=>"00000001",
  14242=>"11111110",
  14243=>"00000000",
  14244=>"00000000",
  14245=>"00000010",
  14246=>"00000011",
  14247=>"11111110",
  14248=>"11111110",
  14249=>"11111101",
  14250=>"00000001",
  14251=>"00000000",
  14252=>"00000000",
  14253=>"11111101",
  14254=>"11111111",
  14255=>"00000100",
  14256=>"00000000",
  14257=>"00000101",
  14258=>"00000001",
  14259=>"00000001",
  14260=>"11111110",
  14261=>"00000010",
  14262=>"00000000",
  14263=>"11111110",
  14264=>"11111111",
  14265=>"11111110",
  14266=>"00000010",
  14267=>"11111101",
  14268=>"11111011",
  14269=>"00000001",
  14270=>"11111101",
  14271=>"00000001",
  14272=>"11111111",
  14273=>"11111101",
  14274=>"11111101",
  14275=>"11111111",
  14276=>"11111101",
  14277=>"11111101",
  14278=>"11111110",
  14279=>"11111111",
  14280=>"00000000",
  14281=>"00000010",
  14282=>"00000110",
  14283=>"00000000",
  14284=>"00000101",
  14285=>"11111111",
  14286=>"00000010",
  14287=>"00000000",
  14288=>"11111110",
  14289=>"11111101",
  14290=>"11111100",
  14291=>"00000001",
  14292=>"00000010",
  14293=>"00000000",
  14294=>"00000011",
  14295=>"11111110",
  14296=>"00000011",
  14297=>"00000000",
  14298=>"00000011",
  14299=>"00000010",
  14300=>"00000011",
  14301=>"00000100",
  14302=>"00000001",
  14303=>"11111110",
  14304=>"00000010",
  14305=>"00000010",
  14306=>"00000000",
  14307=>"11111110",
  14308=>"00000100",
  14309=>"00000010",
  14310=>"00000000",
  14311=>"11111100",
  14312=>"00000001",
  14313=>"00000010",
  14314=>"00000110",
  14315=>"11111101",
  14316=>"11111111",
  14317=>"11111110",
  14318=>"00000001",
  14319=>"11111110",
  14320=>"00000010",
  14321=>"00000010",
  14322=>"00000000",
  14323=>"00000010",
  14324=>"11111111",
  14325=>"00000000",
  14326=>"00000001",
  14327=>"11111111",
  14328=>"00000011",
  14329=>"11111111",
  14330=>"11111111",
  14331=>"00000001",
  14332=>"00000011",
  14333=>"00000001",
  14334=>"00000011",
  14335=>"00000010",
  14336=>"00000000",
  14337=>"11111110",
  14338=>"00000011",
  14339=>"00000001",
  14340=>"00000001",
  14341=>"11111111",
  14342=>"00000100",
  14343=>"11111111",
  14344=>"11111100",
  14345=>"00000011",
  14346=>"11111111",
  14347=>"11111101",
  14348=>"11111110",
  14349=>"11111100",
  14350=>"00000000",
  14351=>"00000010",
  14352=>"00000110",
  14353=>"11111111",
  14354=>"11111111",
  14355=>"11111110",
  14356=>"11111101",
  14357=>"11111110",
  14358=>"00000100",
  14359=>"00000001",
  14360=>"00000000",
  14361=>"00000010",
  14362=>"11111111",
  14363=>"00000001",
  14364=>"00000101",
  14365=>"11111111",
  14366=>"11111110",
  14367=>"11111110",
  14368=>"11111111",
  14369=>"11111101",
  14370=>"00000100",
  14371=>"11111111",
  14372=>"00000010",
  14373=>"00000001",
  14374=>"00000000",
  14375=>"00000011",
  14376=>"00000010",
  14377=>"11111101",
  14378=>"11111110",
  14379=>"00000001",
  14380=>"11111110",
  14381=>"00000010",
  14382=>"00000010",
  14383=>"00000001",
  14384=>"11111111",
  14385=>"11111110",
  14386=>"11111110",
  14387=>"11111111",
  14388=>"00000000",
  14389=>"00000010",
  14390=>"11111110",
  14391=>"11111101",
  14392=>"00000001",
  14393=>"00000000",
  14394=>"00000000",
  14395=>"00000000",
  14396=>"00000011",
  14397=>"11111110",
  14398=>"11111101",
  14399=>"00000000",
  14400=>"11111111",
  14401=>"00000010",
  14402=>"11111101",
  14403=>"11111101",
  14404=>"00000001",
  14405=>"00000001",
  14406=>"11111100",
  14407=>"11111110",
  14408=>"00000010",
  14409=>"11111111",
  14410=>"00000010",
  14411=>"00000001",
  14412=>"11111101",
  14413=>"00000000",
  14414=>"00000001",
  14415=>"00000000",
  14416=>"00001000",
  14417=>"11111101",
  14418=>"00000100",
  14419=>"11111110",
  14420=>"00000011",
  14421=>"00000001",
  14422=>"00000000",
  14423=>"00000010",
  14424=>"11111110",
  14425=>"11111101",
  14426=>"00000000",
  14427=>"11111110",
  14428=>"11111101",
  14429=>"00000010",
  14430=>"00000100",
  14431=>"11111110",
  14432=>"00000000",
  14433=>"00000100",
  14434=>"11111111",
  14435=>"11111101",
  14436=>"11111111",
  14437=>"00000001",
  14438=>"11111111",
  14439=>"11111111",
  14440=>"00000011",
  14441=>"11111101",
  14442=>"11111110",
  14443=>"11111111",
  14444=>"00000001",
  14445=>"00000001",
  14446=>"00000000",
  14447=>"00000001",
  14448=>"00000100",
  14449=>"11111101",
  14450=>"11111110",
  14451=>"00000001",
  14452=>"00000100",
  14453=>"00000001",
  14454=>"00000101",
  14455=>"11111100",
  14456=>"00000000",
  14457=>"00000000",
  14458=>"11111111",
  14459=>"00000100",
  14460=>"11111110",
  14461=>"11111111",
  14462=>"00000000",
  14463=>"00000101",
  14464=>"11111111",
  14465=>"00000011",
  14466=>"00000010",
  14467=>"00000010",
  14468=>"11111111",
  14469=>"11111111",
  14470=>"11111110",
  14471=>"11111110",
  14472=>"00000000",
  14473=>"11111111",
  14474=>"11111110",
  14475=>"11111110",
  14476=>"11111101",
  14477=>"00000010",
  14478=>"11111101",
  14479=>"00000011",
  14480=>"00000100",
  14481=>"11111101",
  14482=>"00000101",
  14483=>"00000001",
  14484=>"00000100",
  14485=>"00000001",
  14486=>"11111111",
  14487=>"00000001",
  14488=>"11111101",
  14489=>"00000001",
  14490=>"00000100",
  14491=>"11111101",
  14492=>"11111101",
  14493=>"11111100",
  14494=>"11111101",
  14495=>"11111110",
  14496=>"00000001",
  14497=>"00000010",
  14498=>"11111100",
  14499=>"00000000",
  14500=>"11111110",
  14501=>"11111110",
  14502=>"00000001",
  14503=>"00000001",
  14504=>"11111111",
  14505=>"11111110",
  14506=>"11111110",
  14507=>"00000000",
  14508=>"00000000",
  14509=>"11111101",
  14510=>"11111110",
  14511=>"11111110",
  14512=>"00000000",
  14513=>"11111111",
  14514=>"00000010",
  14515=>"11111110",
  14516=>"11111100",
  14517=>"11111101",
  14518=>"11111101",
  14519=>"11111110",
  14520=>"00000011",
  14521=>"00000000",
  14522=>"00000001",
  14523=>"00000001",
  14524=>"00000001",
  14525=>"00000000",
  14526=>"11111110",
  14527=>"00000000",
  14528=>"00000000",
  14529=>"11111110",
  14530=>"11111111",
  14531=>"00000001",
  14532=>"11111111",
  14533=>"11111100",
  14534=>"11111101",
  14535=>"00000000",
  14536=>"11111111",
  14537=>"11111111",
  14538=>"11111101",
  14539=>"11111111",
  14540=>"11111111",
  14541=>"00000000",
  14542=>"00000001",
  14543=>"00000011",
  14544=>"00000001",
  14545=>"00000011",
  14546=>"11111111",
  14547=>"00000001",
  14548=>"00000000",
  14549=>"11111111",
  14550=>"11111101",
  14551=>"00000001",
  14552=>"11111101",
  14553=>"11111111",
  14554=>"11111111",
  14555=>"00000010",
  14556=>"11111101",
  14557=>"00000001",
  14558=>"00000000",
  14559=>"11111111",
  14560=>"00000001",
  14561=>"00000000",
  14562=>"11111101",
  14563=>"11111101",
  14564=>"00000000",
  14565=>"11111110",
  14566=>"00000001",
  14567=>"11111110",
  14568=>"00000000",
  14569=>"00000001",
  14570=>"11111111",
  14571=>"11111110",
  14572=>"00000000",
  14573=>"00000011",
  14574=>"11111101",
  14575=>"11111111",
  14576=>"00000000",
  14577=>"00000001",
  14578=>"11111110",
  14579=>"00000001",
  14580=>"00000010",
  14581=>"11111110",
  14582=>"11111111",
  14583=>"00000001",
  14584=>"00000010",
  14585=>"00000001",
  14586=>"00000001",
  14587=>"00000010",
  14588=>"11111110",
  14589=>"00000010",
  14590=>"11111111",
  14591=>"11111101",
  14592=>"00000001",
  14593=>"00000000",
  14594=>"00000000",
  14595=>"11111110",
  14596=>"00000010",
  14597=>"11111101",
  14598=>"00000001",
  14599=>"11111111",
  14600=>"11111110",
  14601=>"00000001",
  14602=>"00000001",
  14603=>"00000001",
  14604=>"00000010",
  14605=>"00000011",
  14606=>"00000100",
  14607=>"11111111",
  14608=>"11111100",
  14609=>"11111101",
  14610=>"11111100",
  14611=>"00000010",
  14612=>"11111111",
  14613=>"11111111",
  14614=>"00000000",
  14615=>"11111101",
  14616=>"11111100",
  14617=>"11111101",
  14618=>"00000010",
  14619=>"11111111",
  14620=>"00000011",
  14621=>"11111111",
  14622=>"11111111",
  14623=>"00000000",
  14624=>"00000010",
  14625=>"00000010",
  14626=>"00000100",
  14627=>"00000001",
  14628=>"11111100",
  14629=>"11111110",
  14630=>"11111111",
  14631=>"11111110",
  14632=>"00000000",
  14633=>"00000001",
  14634=>"00000001",
  14635=>"11111110",
  14636=>"11111111",
  14637=>"00000011",
  14638=>"11111111",
  14639=>"11111110",
  14640=>"11111111",
  14641=>"00000000",
  14642=>"11111101",
  14643=>"11111111",
  14644=>"00000001",
  14645=>"00000010",
  14646=>"00000000",
  14647=>"00000011",
  14648=>"00000000",
  14649=>"00000001",
  14650=>"00000000",
  14651=>"00000001",
  14652=>"00000010",
  14653=>"00000001",
  14654=>"11111110",
  14655=>"00000010",
  14656=>"00000001",
  14657=>"11111110",
  14658=>"11111111",
  14659=>"00000001",
  14660=>"00000000",
  14661=>"11111111",
  14662=>"00000100",
  14663=>"00000010",
  14664=>"00000001",
  14665=>"00000001",
  14666=>"11111100",
  14667=>"00000010",
  14668=>"00000000",
  14669=>"11111111",
  14670=>"11111101",
  14671=>"00000000",
  14672=>"00000101",
  14673=>"11111111",
  14674=>"11111100",
  14675=>"00000011",
  14676=>"00000010",
  14677=>"00000001",
  14678=>"00000100",
  14679=>"00000000",
  14680=>"11111101",
  14681=>"11111111",
  14682=>"11111110",
  14683=>"11111101",
  14684=>"11111101",
  14685=>"00000001",
  14686=>"00000010",
  14687=>"00000010",
  14688=>"00000010",
  14689=>"00000000",
  14690=>"11111110",
  14691=>"11111110",
  14692=>"00000100",
  14693=>"11111110",
  14694=>"11111111",
  14695=>"00000000",
  14696=>"00000000",
  14697=>"11111111",
  14698=>"11111110",
  14699=>"00000001",
  14700=>"00000001",
  14701=>"11111101",
  14702=>"11111011",
  14703=>"00000010",
  14704=>"11111111",
  14705=>"11111101",
  14706=>"00000000",
  14707=>"11111101",
  14708=>"00000000",
  14709=>"11111111",
  14710=>"00000001",
  14711=>"00000010",
  14712=>"00000000",
  14713=>"00000010",
  14714=>"00000001",
  14715=>"00000010",
  14716=>"00000000",
  14717=>"00000001",
  14718=>"11111111",
  14719=>"11111101",
  14720=>"00000010",
  14721=>"00000001",
  14722=>"00000011",
  14723=>"00000001",
  14724=>"00000010",
  14725=>"00000010",
  14726=>"11111101",
  14727=>"00000000",
  14728=>"11111110",
  14729=>"11111110",
  14730=>"00000101",
  14731=>"00000011",
  14732=>"00000000",
  14733=>"11111101",
  14734=>"00000000",
  14735=>"11111111",
  14736=>"11111110",
  14737=>"11111110",
  14738=>"00000010",
  14739=>"00000001",
  14740=>"00000011",
  14741=>"00000000",
  14742=>"11111111",
  14743=>"00000010",
  14744=>"11111110",
  14745=>"00000000",
  14746=>"11111110",
  14747=>"00000011",
  14748=>"00000101",
  14749=>"00000010",
  14750=>"11111111",
  14751=>"00000100",
  14752=>"11111111",
  14753=>"11111100",
  14754=>"00000010",
  14755=>"11111110",
  14756=>"00000100",
  14757=>"00000001",
  14758=>"00000010",
  14759=>"11111101",
  14760=>"00000001",
  14761=>"00000011",
  14762=>"11111110",
  14763=>"11111110",
  14764=>"00000001",
  14765=>"00000010",
  14766=>"00000010",
  14767=>"00000010",
  14768=>"11111101",
  14769=>"11111111",
  14770=>"00000000",
  14771=>"00000010",
  14772=>"00000011",
  14773=>"11111100",
  14774=>"11111110",
  14775=>"11111111",
  14776=>"11111111",
  14777=>"00000000",
  14778=>"11111100",
  14779=>"11111101",
  14780=>"11111110",
  14781=>"00000001",
  14782=>"00001001",
  14783=>"00000001",
  14784=>"11111110",
  14785=>"00000010",
  14786=>"00000001",
  14787=>"11111110",
  14788=>"11111111",
  14789=>"11111111",
  14790=>"00000000",
  14791=>"11111111",
  14792=>"11111110",
  14793=>"00000001",
  14794=>"11111111",
  14795=>"11111100",
  14796=>"00000001",
  14797=>"11111111",
  14798=>"00000100",
  14799=>"11111111",
  14800=>"00000011",
  14801=>"00000001",
  14802=>"11111111",
  14803=>"00000011",
  14804=>"11111111",
  14805=>"00000001",
  14806=>"11111101",
  14807=>"00000001",
  14808=>"11111111",
  14809=>"11111110",
  14810=>"00000001",
  14811=>"00000000",
  14812=>"00000001",
  14813=>"00000011",
  14814=>"11111101",
  14815=>"11111111",
  14816=>"11111111",
  14817=>"11111110",
  14818=>"00000001",
  14819=>"00000001",
  14820=>"00000010",
  14821=>"11111110",
  14822=>"11111100",
  14823=>"00000011",
  14824=>"11111101",
  14825=>"00000001",
  14826=>"00000010",
  14827=>"00000001",
  14828=>"00000011",
  14829=>"00000000",
  14830=>"11111110",
  14831=>"00000011",
  14832=>"11111110",
  14833=>"00000001",
  14834=>"00000010",
  14835=>"11111111",
  14836=>"00000001",
  14837=>"00000010",
  14838=>"11111111",
  14839=>"00000011",
  14840=>"11111110",
  14841=>"11111111",
  14842=>"00000000",
  14843=>"11111100",
  14844=>"11111111",
  14845=>"00000101",
  14846=>"11111110",
  14847=>"00000100",
  14848=>"11111101",
  14849=>"11111110",
  14850=>"11111111",
  14851=>"00000000",
  14852=>"11111111",
  14853=>"11111110",
  14854=>"11111111",
  14855=>"00000010",
  14856=>"11111110",
  14857=>"00000001",
  14858=>"00000000",
  14859=>"11111110",
  14860=>"11111110",
  14861=>"11111101",
  14862=>"11111110",
  14863=>"00000001",
  14864=>"00000001",
  14865=>"00000010",
  14866=>"11111101",
  14867=>"00000000",
  14868=>"00000000",
  14869=>"00000000",
  14870=>"00000000",
  14871=>"00000100",
  14872=>"00000011",
  14873=>"11111110",
  14874=>"00000111",
  14875=>"11111110",
  14876=>"11111101",
  14877=>"11111110",
  14878=>"11111101",
  14879=>"11111101",
  14880=>"11111111",
  14881=>"00000000",
  14882=>"00000110",
  14883=>"11111101",
  14884=>"11111111",
  14885=>"00000000",
  14886=>"00000001",
  14887=>"00000000",
  14888=>"11111101",
  14889=>"11111111",
  14890=>"00000101",
  14891=>"00000000",
  14892=>"11111110",
  14893=>"00000011",
  14894=>"11111101",
  14895=>"11111110",
  14896=>"00000000",
  14897=>"11111111",
  14898=>"00000011",
  14899=>"00000000",
  14900=>"11111100",
  14901=>"11111101",
  14902=>"11111111",
  14903=>"11111101",
  14904=>"11111110",
  14905=>"11111101",
  14906=>"00000000",
  14907=>"00000000",
  14908=>"00000101",
  14909=>"11111111",
  14910=>"00000000",
  14911=>"11111101",
  14912=>"11111101",
  14913=>"00000011",
  14914=>"11111101",
  14915=>"00000001",
  14916=>"11111101",
  14917=>"00000010",
  14918=>"11111101",
  14919=>"11111110",
  14920=>"11111111",
  14921=>"00000000",
  14922=>"00000001",
  14923=>"00000010",
  14924=>"00000000",
  14925=>"11111101",
  14926=>"11111101",
  14927=>"11111111",
  14928=>"00000000",
  14929=>"00000011",
  14930=>"00000110",
  14931=>"00000001",
  14932=>"00000000",
  14933=>"11111101",
  14934=>"00000010",
  14935=>"00000011",
  14936=>"11111111",
  14937=>"11111100",
  14938=>"00000000",
  14939=>"00000000",
  14940=>"00000000",
  14941=>"11111110",
  14942=>"11111111",
  14943=>"00000000",
  14944=>"00000001",
  14945=>"00000000",
  14946=>"11111110",
  14947=>"00000010",
  14948=>"00000000",
  14949=>"11111110",
  14950=>"11111110",
  14951=>"00000011",
  14952=>"00000111",
  14953=>"11111101",
  14954=>"00000010",
  14955=>"00000001",
  14956=>"11111110",
  14957=>"00000100",
  14958=>"00000010",
  14959=>"00000010",
  14960=>"00000000",
  14961=>"00000001",
  14962=>"00000000",
  14963=>"11111110",
  14964=>"00000010",
  14965=>"11111111",
  14966=>"11111101",
  14967=>"11111110",
  14968=>"11111111",
  14969=>"00000001",
  14970=>"00000001",
  14971=>"00000010",
  14972=>"00000010",
  14973=>"11111101",
  14974=>"00000000",
  14975=>"00000000",
  14976=>"00000010",
  14977=>"00000010",
  14978=>"00000000",
  14979=>"11111111",
  14980=>"00000010",
  14981=>"11111111",
  14982=>"11111101",
  14983=>"00000100",
  14984=>"00000001",
  14985=>"11111101",
  14986=>"11111111",
  14987=>"00000011",
  14988=>"00000011",
  14989=>"11111111",
  14990=>"00000010",
  14991=>"00000011",
  14992=>"11111111",
  14993=>"11111111",
  14994=>"11111101",
  14995=>"11111111",
  14996=>"00000010",
  14997=>"11111110",
  14998=>"00000010",
  14999=>"11111110",
  15000=>"00000100",
  15001=>"00000001",
  15002=>"11111100",
  15003=>"00000010",
  15004=>"00000000",
  15005=>"00000000",
  15006=>"11111110",
  15007=>"11111110",
  15008=>"00000000",
  15009=>"00000011",
  15010=>"00000000",
  15011=>"11111110",
  15012=>"11111111",
  15013=>"00000100",
  15014=>"11111100",
  15015=>"11111100",
  15016=>"11111101",
  15017=>"00000001",
  15018=>"11111101",
  15019=>"11111101",
  15020=>"11111110",
  15021=>"00000100",
  15022=>"00000010",
  15023=>"11111110",
  15024=>"11111111",
  15025=>"00000110",
  15026=>"00000001",
  15027=>"11111101",
  15028=>"11111101",
  15029=>"11111111",
  15030=>"11111110",
  15031=>"11111110",
  15032=>"00000011",
  15033=>"00000000",
  15034=>"00000011",
  15035=>"00000000",
  15036=>"11111101",
  15037=>"11111110",
  15038=>"00000110",
  15039=>"11111111",
  15040=>"11111110",
  15041=>"00000010",
  15042=>"00000011",
  15043=>"00000000",
  15044=>"00000011",
  15045=>"11111101",
  15046=>"00000000",
  15047=>"00000010",
  15048=>"00000010",
  15049=>"11111111",
  15050=>"00000000",
  15051=>"11111101",
  15052=>"11111110",
  15053=>"00000001",
  15054=>"00000000",
  15055=>"00000010",
  15056=>"00000000",
  15057=>"11111101",
  15058=>"00000001",
  15059=>"00000001",
  15060=>"00000001",
  15061=>"11111100",
  15062=>"00000010",
  15063=>"00000000",
  15064=>"11111111",
  15065=>"00000010",
  15066=>"11111110",
  15067=>"00000000",
  15068=>"11111100",
  15069=>"11111110",
  15070=>"00000100",
  15071=>"11111110",
  15072=>"00000100",
  15073=>"00000001",
  15074=>"00000001",
  15075=>"11111111",
  15076=>"11111101",
  15077=>"11111110",
  15078=>"11111110",
  15079=>"00000010",
  15080=>"00000011",
  15081=>"00000010",
  15082=>"00000010",
  15083=>"11111111",
  15084=>"00000000",
  15085=>"11111111",
  15086=>"11111101",
  15087=>"11111100",
  15088=>"00000000",
  15089=>"00000011",
  15090=>"00000001",
  15091=>"11111111",
  15092=>"00000101",
  15093=>"00000000",
  15094=>"11111101",
  15095=>"00000000",
  15096=>"00000000",
  15097=>"11111111",
  15098=>"00000010",
  15099=>"00000000",
  15100=>"00000000",
  15101=>"00000011",
  15102=>"00000101",
  15103=>"11111111",
  15104=>"00000000",
  15105=>"00000010",
  15106=>"11111110",
  15107=>"00000011",
  15108=>"11111100",
  15109=>"11111111",
  15110=>"11111111",
  15111=>"00000010",
  15112=>"11111101",
  15113=>"00000000",
  15114=>"11111111",
  15115=>"00000001",
  15116=>"00001000",
  15117=>"11111110",
  15118=>"00000001",
  15119=>"00000010",
  15120=>"11111110",
  15121=>"00000000",
  15122=>"11111101",
  15123=>"11111110",
  15124=>"11111111",
  15125=>"11111110",
  15126=>"00000010",
  15127=>"00000000",
  15128=>"00000000",
  15129=>"00000010",
  15130=>"11111110",
  15131=>"11111101",
  15132=>"11111110",
  15133=>"00000001",
  15134=>"00000000",
  15135=>"00000000",
  15136=>"00000011",
  15137=>"11111111",
  15138=>"00000001",
  15139=>"11111011",
  15140=>"00000010",
  15141=>"11111100",
  15142=>"11111100",
  15143=>"11111100",
  15144=>"00000000",
  15145=>"11111111",
  15146=>"00000010",
  15147=>"11111111",
  15148=>"00000001",
  15149=>"00000001",
  15150=>"11111101",
  15151=>"11111101",
  15152=>"11111110",
  15153=>"11111110",
  15154=>"00000000",
  15155=>"11111110",
  15156=>"00000000",
  15157=>"00000101",
  15158=>"11111101",
  15159=>"11111101",
  15160=>"11111110",
  15161=>"11111110",
  15162=>"11111101",
  15163=>"11111110",
  15164=>"00000000",
  15165=>"00000100",
  15166=>"11111110",
  15167=>"00000001",
  15168=>"11111110",
  15169=>"00000000",
  15170=>"00000001",
  15171=>"11111101",
  15172=>"00000000",
  15173=>"00000010",
  15174=>"00000000",
  15175=>"11111110",
  15176=>"11111110",
  15177=>"11111101",
  15178=>"00000001",
  15179=>"00000011",
  15180=>"00000001",
  15181=>"00000001",
  15182=>"00000001",
  15183=>"00000011",
  15184=>"11111110",
  15185=>"11111111",
  15186=>"11111110",
  15187=>"00000000",
  15188=>"11111110",
  15189=>"11111110",
  15190=>"00000001",
  15191=>"11111101",
  15192=>"00000001",
  15193=>"00000011",
  15194=>"00000000",
  15195=>"00000000",
  15196=>"00000001",
  15197=>"00000010",
  15198=>"00000010",
  15199=>"11111110",
  15200=>"11111111",
  15201=>"11111111",
  15202=>"00000000",
  15203=>"00000000",
  15204=>"11111101",
  15205=>"00000010",
  15206=>"11111101",
  15207=>"11111110",
  15208=>"11111110",
  15209=>"00000000",
  15210=>"11111101",
  15211=>"11111101",
  15212=>"00000000",
  15213=>"00000100",
  15214=>"00000100",
  15215=>"00000000",
  15216=>"11111110",
  15217=>"11111110",
  15218=>"11111110",
  15219=>"11111101",
  15220=>"00000000",
  15221=>"00000110",
  15222=>"11111111",
  15223=>"11111110",
  15224=>"00000010",
  15225=>"11111101",
  15226=>"00000000",
  15227=>"00000000",
  15228=>"00000011",
  15229=>"11111111",
  15230=>"00000011",
  15231=>"11111101",
  15232=>"00000011",
  15233=>"11111111",
  15234=>"11111101",
  15235=>"11111100",
  15236=>"11111110",
  15237=>"11111101",
  15238=>"11111110",
  15239=>"00000010",
  15240=>"00000001",
  15241=>"11111110",
  15242=>"00000000",
  15243=>"11111110",
  15244=>"11111110",
  15245=>"00000000",
  15246=>"00000010",
  15247=>"11111111",
  15248=>"00000011",
  15249=>"11111100",
  15250=>"00000000",
  15251=>"11111110",
  15252=>"11111100",
  15253=>"11111100",
  15254=>"00000000",
  15255=>"00000110",
  15256=>"11111100",
  15257=>"11111101",
  15258=>"00000000",
  15259=>"00000011",
  15260=>"00000000",
  15261=>"11111111",
  15262=>"00000100",
  15263=>"11111110",
  15264=>"00000001",
  15265=>"11111101",
  15266=>"11111111",
  15267=>"00000011",
  15268=>"11111101",
  15269=>"00000000",
  15270=>"11111111",
  15271=>"00000010",
  15272=>"11111101",
  15273=>"11111100",
  15274=>"00000001",
  15275=>"00000000",
  15276=>"11111111",
  15277=>"00000011",
  15278=>"00000100",
  15279=>"11111110",
  15280=>"00000010",
  15281=>"11111110",
  15282=>"00000101",
  15283=>"00000011",
  15284=>"00000000",
  15285=>"11111110",
  15286=>"00000011",
  15287=>"00000000",
  15288=>"11111111",
  15289=>"11111111",
  15290=>"00000000",
  15291=>"00000001",
  15292=>"00000010",
  15293=>"11111111",
  15294=>"11111110",
  15295=>"00000000",
  15296=>"00000000",
  15297=>"00000001",
  15298=>"11111111",
  15299=>"00000001",
  15300=>"00000000",
  15301=>"00000011",
  15302=>"11111110",
  15303=>"00000000",
  15304=>"00000001",
  15305=>"11111101",
  15306=>"00000010",
  15307=>"11111111",
  15308=>"11111100",
  15309=>"00000001",
  15310=>"00000001",
  15311=>"00000001",
  15312=>"11111111",
  15313=>"11111110",
  15314=>"00000100",
  15315=>"00000100",
  15316=>"00000011",
  15317=>"00000000",
  15318=>"00000000",
  15319=>"11111110",
  15320=>"11111101",
  15321=>"11111011",
  15322=>"11111101",
  15323=>"00000001",
  15324=>"00000001",
  15325=>"11111110",
  15326=>"11111101",
  15327=>"11111101",
  15328=>"00000010",
  15329=>"00000000",
  15330=>"00000000",
  15331=>"11111111",
  15332=>"11111110",
  15333=>"00000011",
  15334=>"00000100",
  15335=>"11111101",
  15336=>"11111101",
  15337=>"00000010",
  15338=>"11111110",
  15339=>"11111101",
  15340=>"00000000",
  15341=>"11111111",
  15342=>"11111111",
  15343=>"00000100",
  15344=>"00000000",
  15345=>"00000100",
  15346=>"00000001",
  15347=>"00000000",
  15348=>"11111111",
  15349=>"11111111",
  15350=>"11111111",
  15351=>"00000000",
  15352=>"11111111",
  15353=>"11111111",
  15354=>"00000000",
  15355=>"00000011",
  15356=>"00000001",
  15357=>"00000000",
  15358=>"00000001",
  15359=>"00000001",
  15360=>"11111101",
  15361=>"00000000",
  15362=>"11111110",
  15363=>"11111110",
  15364=>"11111111",
  15365=>"00000010",
  15366=>"00000000",
  15367=>"00000101",
  15368=>"00000010",
  15369=>"11111101",
  15370=>"00000010",
  15371=>"11111110",
  15372=>"11111110",
  15373=>"11111110",
  15374=>"11111110",
  15375=>"00000001",
  15376=>"11111101",
  15377=>"11111110",
  15378=>"11111101",
  15379=>"00000001",
  15380=>"11111111",
  15381=>"00000000",
  15382=>"11111111",
  15383=>"00000010",
  15384=>"11111100",
  15385=>"00000010",
  15386=>"00000100",
  15387=>"00000010",
  15388=>"11111111",
  15389=>"00000100",
  15390=>"00000001",
  15391=>"00000000",
  15392=>"11111110",
  15393=>"11111111",
  15394=>"00000011",
  15395=>"00000010",
  15396=>"11111111",
  15397=>"11111111",
  15398=>"11111111",
  15399=>"11111101",
  15400=>"11111111",
  15401=>"00000000",
  15402=>"11111111",
  15403=>"00000110",
  15404=>"00000010",
  15405=>"00000000",
  15406=>"00000000",
  15407=>"00000010",
  15408=>"00000001",
  15409=>"00000001",
  15410=>"11111111",
  15411=>"11111111",
  15412=>"11111111",
  15413=>"00000010",
  15414=>"11111111",
  15415=>"11111101",
  15416=>"00000001",
  15417=>"11111110",
  15418=>"11111101",
  15419=>"11111110",
  15420=>"11111110",
  15421=>"00000000",
  15422=>"00000000",
  15423=>"11111111",
  15424=>"00000011",
  15425=>"11111110",
  15426=>"11111111",
  15427=>"11111111",
  15428=>"00000001",
  15429=>"00000011",
  15430=>"11111111",
  15431=>"11111101",
  15432=>"11111111",
  15433=>"00000000",
  15434=>"00000010",
  15435=>"11111110",
  15436=>"11111111",
  15437=>"11111111",
  15438=>"00000001",
  15439=>"11111110",
  15440=>"11111101",
  15441=>"11111111",
  15442=>"11111111",
  15443=>"00000000",
  15444=>"11111110",
  15445=>"00000001",
  15446=>"00000101",
  15447=>"00000010",
  15448=>"11111101",
  15449=>"00000001",
  15450=>"11111110",
  15451=>"11111110",
  15452=>"11111111",
  15453=>"00000000",
  15454=>"00000000",
  15455=>"00000000",
  15456=>"00000011",
  15457=>"11111101",
  15458=>"00000010",
  15459=>"00000000",
  15460=>"00000101",
  15461=>"11111101",
  15462=>"00000001",
  15463=>"11111110",
  15464=>"00000001",
  15465=>"11111111",
  15466=>"11111111",
  15467=>"11111101",
  15468=>"00000010",
  15469=>"00000000",
  15470=>"11111111",
  15471=>"11111100",
  15472=>"11111111",
  15473=>"00000001",
  15474=>"00000001",
  15475=>"00000001",
  15476=>"00000001",
  15477=>"11111110",
  15478=>"00000000",
  15479=>"00000000",
  15480=>"11111101",
  15481=>"00000001",
  15482=>"00000010",
  15483=>"00000000",
  15484=>"11111111",
  15485=>"11111110",
  15486=>"00000010",
  15487=>"11111111",
  15488=>"11111111",
  15489=>"00000001",
  15490=>"11111101",
  15491=>"11111111",
  15492=>"00000001",
  15493=>"00000010",
  15494=>"00000001",
  15495=>"00000000",
  15496=>"11111111",
  15497=>"11111110",
  15498=>"00000010",
  15499=>"00000000",
  15500=>"11111111",
  15501=>"11111110",
  15502=>"11111111",
  15503=>"00000011",
  15504=>"00000010",
  15505=>"00000011",
  15506=>"00000001",
  15507=>"11111111",
  15508=>"11111110",
  15509=>"11111111",
  15510=>"11111111",
  15511=>"00000001",
  15512=>"11111110",
  15513=>"00000001",
  15514=>"11111110",
  15515=>"00000000",
  15516=>"11111110",
  15517=>"11111101",
  15518=>"00000010",
  15519=>"00000001",
  15520=>"00000100",
  15521=>"11111110",
  15522=>"11111110",
  15523=>"00000000",
  15524=>"00000010",
  15525=>"00000010",
  15526=>"11111110",
  15527=>"11111111",
  15528=>"11111101",
  15529=>"11111110",
  15530=>"00000010",
  15531=>"11111111",
  15532=>"11111111",
  15533=>"11111101",
  15534=>"00000000",
  15535=>"11111110",
  15536=>"11111110",
  15537=>"11111110",
  15538=>"00000000",
  15539=>"00000000",
  15540=>"11111111",
  15541=>"00000001",
  15542=>"11111101",
  15543=>"00000001",
  15544=>"00000000",
  15545=>"11111111",
  15546=>"11111110",
  15547=>"00000010",
  15548=>"11111111",
  15549=>"11111111",
  15550=>"00000010",
  15551=>"11111100",
  15552=>"11111111",
  15553=>"00000010",
  15554=>"00000000",
  15555=>"11111110",
  15556=>"00000000",
  15557=>"00000010",
  15558=>"00000001",
  15559=>"00000001",
  15560=>"11111100",
  15561=>"00000000",
  15562=>"11111101",
  15563=>"11111110",
  15564=>"00000001",
  15565=>"00000001",
  15566=>"00000000",
  15567=>"00000101",
  15568=>"00000000",
  15569=>"11111111",
  15570=>"11111110",
  15571=>"11111111",
  15572=>"11111101",
  15573=>"00000000",
  15574=>"11111101",
  15575=>"00000010",
  15576=>"00000000",
  15577=>"11111111",
  15578=>"00000000",
  15579=>"00000001",
  15580=>"00000000",
  15581=>"11111110",
  15582=>"00000001",
  15583=>"00000101",
  15584=>"00000010",
  15585=>"00000000",
  15586=>"11111110",
  15587=>"11111111",
  15588=>"11111111",
  15589=>"00000011",
  15590=>"11111101",
  15591=>"00000011",
  15592=>"11111111",
  15593=>"11111110",
  15594=>"00000010",
  15595=>"00000011",
  15596=>"00000001",
  15597=>"11111110",
  15598=>"00000010",
  15599=>"11111111",
  15600=>"00000011",
  15601=>"11111110",
  15602=>"00000011",
  15603=>"00000001",
  15604=>"00000000",
  15605=>"00000011",
  15606=>"11111111",
  15607=>"11111101",
  15608=>"11111110",
  15609=>"00000011",
  15610=>"11111101",
  15611=>"00000001",
  15612=>"11111101",
  15613=>"00000010",
  15614=>"00000010",
  15615=>"00000011",
  15616=>"11111111",
  15617=>"00000100",
  15618=>"11111110",
  15619=>"11111101",
  15620=>"00000010",
  15621=>"11111111",
  15622=>"00000000",
  15623=>"11111101",
  15624=>"11111111",
  15625=>"11111111",
  15626=>"00000010",
  15627=>"11111111",
  15628=>"00000001",
  15629=>"00000010",
  15630=>"00000011",
  15631=>"11111111",
  15632=>"00000101",
  15633=>"00000100",
  15634=>"00000011",
  15635=>"11111111",
  15636=>"00000001",
  15637=>"11111110",
  15638=>"00000010",
  15639=>"11111100",
  15640=>"11111101",
  15641=>"00000010",
  15642=>"00000001",
  15643=>"11111101",
  15644=>"00000010",
  15645=>"00000001",
  15646=>"11111101",
  15647=>"11111110",
  15648=>"00000000",
  15649=>"11111111",
  15650=>"11111110",
  15651=>"00000000",
  15652=>"00000011",
  15653=>"00000001",
  15654=>"00000000",
  15655=>"00000000",
  15656=>"11111110",
  15657=>"00000000",
  15658=>"00000001",
  15659=>"11111101",
  15660=>"11111111",
  15661=>"00000000",
  15662=>"11111111",
  15663=>"11111101",
  15664=>"11111110",
  15665=>"00000000",
  15666=>"00000001",
  15667=>"11111110",
  15668=>"00000100",
  15669=>"11111111",
  15670=>"11111101",
  15671=>"00000001",
  15672=>"11111110",
  15673=>"11111100",
  15674=>"00000001",
  15675=>"11111101",
  15676=>"00000000",
  15677=>"00000011",
  15678=>"11111111",
  15679=>"11111111",
  15680=>"11111111",
  15681=>"00000001",
  15682=>"00000001",
  15683=>"11111101",
  15684=>"00000000",
  15685=>"11111101",
  15686=>"00000000",
  15687=>"00000011",
  15688=>"00000000",
  15689=>"11111110",
  15690=>"11111111",
  15691=>"00000010",
  15692=>"00000010",
  15693=>"00000001",
  15694=>"11111110",
  15695=>"11111110",
  15696=>"11111110",
  15697=>"00000010",
  15698=>"11111110",
  15699=>"11111101",
  15700=>"00000000",
  15701=>"11111111",
  15702=>"00000001",
  15703=>"00000000",
  15704=>"00000000",
  15705=>"00000011",
  15706=>"00000001",
  15707=>"11111110",
  15708=>"00000010",
  15709=>"11111101",
  15710=>"11111110",
  15711=>"11111110",
  15712=>"00000100",
  15713=>"11111110",
  15714=>"11111110",
  15715=>"00000000",
  15716=>"11111110",
  15717=>"00000011",
  15718=>"11111111",
  15719=>"11111101",
  15720=>"00000100",
  15721=>"00000000",
  15722=>"00000011",
  15723=>"00000001",
  15724=>"11111110",
  15725=>"11111110",
  15726=>"00000010",
  15727=>"00000000",
  15728=>"11111110",
  15729=>"11111110",
  15730=>"00000010",
  15731=>"00000000",
  15732=>"00000000",
  15733=>"00000000",
  15734=>"11111110",
  15735=>"11111110",
  15736=>"00000000",
  15737=>"00000011",
  15738=>"11111111",
  15739=>"00000000",
  15740=>"11111110",
  15741=>"00000000",
  15742=>"11111111",
  15743=>"11111110",
  15744=>"00000000",
  15745=>"00000010",
  15746=>"00000000",
  15747=>"00000100",
  15748=>"00000000",
  15749=>"11111110",
  15750=>"00000110",
  15751=>"00000000",
  15752=>"00000001",
  15753=>"00000010",
  15754=>"11111110",
  15755=>"11111110",
  15756=>"11111110",
  15757=>"11111110",
  15758=>"00000001",
  15759=>"00000000",
  15760=>"11111101",
  15761=>"11111110",
  15762=>"11111111",
  15763=>"00000000",
  15764=>"00000010",
  15765=>"00000010",
  15766=>"00000000",
  15767=>"11111101",
  15768=>"00000011",
  15769=>"00000010",
  15770=>"00000000",
  15771=>"00000010",
  15772=>"11111111",
  15773=>"00000010",
  15774=>"00000010",
  15775=>"11111101",
  15776=>"00000010",
  15777=>"11111110",
  15778=>"11111101",
  15779=>"11111111",
  15780=>"11111111",
  15781=>"11111100",
  15782=>"00000011",
  15783=>"11111110",
  15784=>"00000100",
  15785=>"11111101",
  15786=>"11111110",
  15787=>"11111101",
  15788=>"11111100",
  15789=>"00000001",
  15790=>"11111111",
  15791=>"11111110",
  15792=>"11111110",
  15793=>"00000010",
  15794=>"00000101",
  15795=>"00000001",
  15796=>"00000000",
  15797=>"00000000",
  15798=>"00000010",
  15799=>"11111101",
  15800=>"11111111",
  15801=>"11111111",
  15802=>"00000100",
  15803=>"11111101",
  15804=>"11111111",
  15805=>"00000001",
  15806=>"11111110",
  15807=>"11111101",
  15808=>"11111110",
  15809=>"11111110",
  15810=>"00000001",
  15811=>"00000001",
  15812=>"11111110",
  15813=>"11111110",
  15814=>"00000100",
  15815=>"11111110",
  15816=>"11111111",
  15817=>"00000001",
  15818=>"11111110",
  15819=>"00000000",
  15820=>"00000001",
  15821=>"11111111",
  15822=>"00000010",
  15823=>"00000001",
  15824=>"11111111",
  15825=>"00000001",
  15826=>"00000001",
  15827=>"00000011",
  15828=>"00000000",
  15829=>"11111111",
  15830=>"11111110",
  15831=>"11111101",
  15832=>"11111101",
  15833=>"11111101",
  15834=>"11111101",
  15835=>"11111111",
  15836=>"00000010",
  15837=>"11111110",
  15838=>"11111111",
  15839=>"00000011",
  15840=>"00000000",
  15841=>"00000110",
  15842=>"11111111",
  15843=>"00000001",
  15844=>"11111111",
  15845=>"11111101",
  15846=>"00000010",
  15847=>"00000001",
  15848=>"11111101",
  15849=>"11111101",
  15850=>"11111110",
  15851=>"00000001",
  15852=>"00000000",
  15853=>"11111101",
  15854=>"00000000",
  15855=>"00000010",
  15856=>"00000001",
  15857=>"11111101",
  15858=>"00000010",
  15859=>"11111111",
  15860=>"00000000",
  15861=>"00000100",
  15862=>"11111110",
  15863=>"00000010",
  15864=>"11111101",
  15865=>"11111110",
  15866=>"11111110",
  15867=>"00000011",
  15868=>"00000000",
  15869=>"00000000",
  15870=>"00000010",
  15871=>"11111100",
  15872=>"00000000",
  15873=>"11111110",
  15874=>"00000001",
  15875=>"00000000",
  15876=>"11111111",
  15877=>"00000010",
  15878=>"11111111",
  15879=>"11111111",
  15880=>"00000000",
  15881=>"00000000",
  15882=>"11111110",
  15883=>"11111110",
  15884=>"00000010",
  15885=>"00000001",
  15886=>"11111111",
  15887=>"00000001",
  15888=>"00000010",
  15889=>"11111100",
  15890=>"00000011",
  15891=>"00000010",
  15892=>"00000110",
  15893=>"11111110",
  15894=>"11111111",
  15895=>"11111110",
  15896=>"00000010",
  15897=>"11111110",
  15898=>"11111100",
  15899=>"11111110",
  15900=>"00000010",
  15901=>"00000011",
  15902=>"11111110",
  15903=>"00000000",
  15904=>"11111110",
  15905=>"00000011",
  15906=>"11111111",
  15907=>"00000001",
  15908=>"11111111",
  15909=>"00000010",
  15910=>"11111110",
  15911=>"11111101",
  15912=>"00000001",
  15913=>"11111110",
  15914=>"11111110",
  15915=>"00000000",
  15916=>"11111111",
  15917=>"11111111",
  15918=>"11111110",
  15919=>"00000010",
  15920=>"00000000",
  15921=>"11111110",
  15922=>"00000001",
  15923=>"11111110",
  15924=>"11111111",
  15925=>"00000101",
  15926=>"11111111",
  15927=>"11111101",
  15928=>"11111111",
  15929=>"11111111",
  15930=>"00000000",
  15931=>"11111110",
  15932=>"11111111",
  15933=>"00000010",
  15934=>"00000010",
  15935=>"00000001",
  15936=>"00000000",
  15937=>"11111101",
  15938=>"11111110",
  15939=>"11111101",
  15940=>"00000001",
  15941=>"11111110",
  15942=>"11111101",
  15943=>"11111111",
  15944=>"00000000",
  15945=>"11111110",
  15946=>"00000100",
  15947=>"00000001",
  15948=>"00000000",
  15949=>"11111101",
  15950=>"00000001",
  15951=>"00000010",
  15952=>"11111111",
  15953=>"11111110",
  15954=>"11111101",
  15955=>"00000010",
  15956=>"11111110",
  15957=>"00000001",
  15958=>"11111101",
  15959=>"00000001",
  15960=>"11111110",
  15961=>"11111111",
  15962=>"00000011",
  15963=>"11111110",
  15964=>"11111101",
  15965=>"00000001",
  15966=>"00000001",
  15967=>"00000001",
  15968=>"00000011",
  15969=>"00000010",
  15970=>"00000001",
  15971=>"00000001",
  15972=>"11111101",
  15973=>"00000001",
  15974=>"11111110",
  15975=>"00000001",
  15976=>"11111101",
  15977=>"11111110",
  15978=>"11111111",
  15979=>"00000000",
  15980=>"11111111",
  15981=>"11111101",
  15982=>"00000000",
  15983=>"00000001",
  15984=>"11111110",
  15985=>"00000000",
  15986=>"00000010",
  15987=>"00000001",
  15988=>"11111111",
  15989=>"00000001",
  15990=>"11111110",
  15991=>"00000001",
  15992=>"11111110",
  15993=>"11111101",
  15994=>"00000000",
  15995=>"11111110",
  15996=>"00000010",
  15997=>"11111111",
  15998=>"00000011",
  15999=>"00000001",
  16000=>"11111111",
  16001=>"00000001",
  16002=>"00000000",
  16003=>"00000000",
  16004=>"11111110",
  16005=>"00000000",
  16006=>"11111101",
  16007=>"11111111",
  16008=>"00000011",
  16009=>"00000001",
  16010=>"11111100",
  16011=>"11111110",
  16012=>"00000001",
  16013=>"00000001",
  16014=>"00000001",
  16015=>"11111110",
  16016=>"00000001",
  16017=>"11111111",
  16018=>"00000001",
  16019=>"00000000",
  16020=>"11111101",
  16021=>"00000010",
  16022=>"00000001",
  16023=>"11111101",
  16024=>"00000010",
  16025=>"00000001",
  16026=>"11111111",
  16027=>"00000001",
  16028=>"11111101",
  16029=>"11111101",
  16030=>"11111111",
  16031=>"11111111",
  16032=>"00000010",
  16033=>"00000001",
  16034=>"11111101",
  16035=>"00000000",
  16036=>"00000000",
  16037=>"00000001",
  16038=>"00000001",
  16039=>"11111101",
  16040=>"11111111",
  16041=>"00000001",
  16042=>"11111110",
  16043=>"11111110",
  16044=>"11111111",
  16045=>"11111101",
  16046=>"00000000",
  16047=>"11111111",
  16048=>"11111111",
  16049=>"11111100",
  16050=>"11111101",
  16051=>"11111111",
  16052=>"00000001",
  16053=>"00000001",
  16054=>"00000000",
  16055=>"00000010",
  16056=>"00000010",
  16057=>"00000001",
  16058=>"11111111",
  16059=>"11111110",
  16060=>"11111110",
  16061=>"00000001",
  16062=>"11111101",
  16063=>"00000011",
  16064=>"11111111",
  16065=>"11111111",
  16066=>"11111111",
  16067=>"00000000",
  16068=>"00000010",
  16069=>"11111110",
  16070=>"00000010",
  16071=>"11111110",
  16072=>"11111101",
  16073=>"00000000",
  16074=>"11111111",
  16075=>"00000010",
  16076=>"11111110",
  16077=>"00000001",
  16078=>"00000010",
  16079=>"00000010",
  16080=>"00000010",
  16081=>"11111101",
  16082=>"00000000",
  16083=>"00000001",
  16084=>"00000010",
  16085=>"00000100",
  16086=>"11111110",
  16087=>"11111110",
  16088=>"00000001",
  16089=>"00000000",
  16090=>"00000001",
  16091=>"00000011",
  16092=>"11111111",
  16093=>"00000010",
  16094=>"00000010",
  16095=>"00000010",
  16096=>"11111101",
  16097=>"11111100",
  16098=>"00000000",
  16099=>"00000001",
  16100=>"11111110",
  16101=>"11111111",
  16102=>"11111101",
  16103=>"11111110",
  16104=>"00000001",
  16105=>"00000000",
  16106=>"00000001",
  16107=>"00000011",
  16108=>"11111111",
  16109=>"00000000",
  16110=>"00000001",
  16111=>"11111101",
  16112=>"00000001",
  16113=>"00000010",
  16114=>"00000100",
  16115=>"00000001",
  16116=>"11111111",
  16117=>"11111101",
  16118=>"00000010",
  16119=>"11111101",
  16120=>"00000010",
  16121=>"00000001",
  16122=>"00000010",
  16123=>"00000010",
  16124=>"00000001",
  16125=>"00000000",
  16126=>"00000000",
  16127=>"00000000",
  16128=>"00000001",
  16129=>"11111101",
  16130=>"11111111",
  16131=>"00000010",
  16132=>"00000010",
  16133=>"00000000",
  16134=>"11111111",
  16135=>"00000100",
  16136=>"11111110",
  16137=>"00000010",
  16138=>"11111111",
  16139=>"00000000",
  16140=>"11111111",
  16141=>"11111100",
  16142=>"00000010",
  16143=>"11111111",
  16144=>"00000011",
  16145=>"11111111",
  16146=>"00000010",
  16147=>"11111111",
  16148=>"00000000",
  16149=>"00000010",
  16150=>"00000000",
  16151=>"11111110",
  16152=>"11111111",
  16153=>"00000000",
  16154=>"11111101",
  16155=>"00000100",
  16156=>"11111110",
  16157=>"00000001",
  16158=>"00000001",
  16159=>"00000010",
  16160=>"00000011",
  16161=>"00000001",
  16162=>"00000001",
  16163=>"11111111",
  16164=>"00000000",
  16165=>"00000010",
  16166=>"11111101",
  16167=>"00000100",
  16168=>"00000010",
  16169=>"00000000",
  16170=>"11111111",
  16171=>"11111110",
  16172=>"00000000",
  16173=>"00000001",
  16174=>"00000001",
  16175=>"11111111",
  16176=>"11111110",
  16177=>"00000001",
  16178=>"00000010",
  16179=>"00000010",
  16180=>"11111111",
  16181=>"00000001",
  16182=>"00000011",
  16183=>"00000001",
  16184=>"11111110",
  16185=>"11111101",
  16186=>"00000010",
  16187=>"11111110",
  16188=>"00000100",
  16189=>"11111110",
  16190=>"11111110",
  16191=>"00000001",
  16192=>"11111110",
  16193=>"00000101",
  16194=>"11111111",
  16195=>"00000010",
  16196=>"00000101",
  16197=>"11111111",
  16198=>"00000010",
  16199=>"00000001",
  16200=>"00000010",
  16201=>"00000001",
  16202=>"11111110",
  16203=>"11111111",
  16204=>"00000000",
  16205=>"00000011",
  16206=>"00000100",
  16207=>"00000001",
  16208=>"00000000",
  16209=>"00000001",
  16210=>"00000001",
  16211=>"00000100",
  16212=>"00000001",
  16213=>"00000000",
  16214=>"00000001",
  16215=>"00000000",
  16216=>"00000001",
  16217=>"11111111",
  16218=>"00000010",
  16219=>"11111110",
  16220=>"00000001",
  16221=>"11111101",
  16222=>"00000011",
  16223=>"11111111",
  16224=>"00000100",
  16225=>"11111110",
  16226=>"11111100",
  16227=>"00000110",
  16228=>"00000000",
  16229=>"00000010",
  16230=>"00000000",
  16231=>"11111110",
  16232=>"11111101",
  16233=>"11111101",
  16234=>"00000001",
  16235=>"00000001",
  16236=>"11111101",
  16237=>"00000010",
  16238=>"00000001",
  16239=>"00000001",
  16240=>"00000000",
  16241=>"00000000",
  16242=>"11111111",
  16243=>"11111111",
  16244=>"00000010",
  16245=>"11111101",
  16246=>"00000001",
  16247=>"00000001",
  16248=>"00000000",
  16249=>"00000001",
  16250=>"00000011",
  16251=>"11111111",
  16252=>"00000000",
  16253=>"00000011",
  16254=>"00000000",
  16255=>"00000011",
  16256=>"11111110",
  16257=>"00000001",
  16258=>"00000001",
  16259=>"00000001",
  16260=>"11111110",
  16261=>"11111111",
  16262=>"00000010",
  16263=>"11111111",
  16264=>"11111111",
  16265=>"00000001",
  16266=>"00000000",
  16267=>"11111111",
  16268=>"11111110",
  16269=>"11111110",
  16270=>"00000010",
  16271=>"11111101",
  16272=>"00000000",
  16273=>"00000010",
  16274=>"11111110",
  16275=>"11111111",
  16276=>"00000001",
  16277=>"11111101",
  16278=>"11111110",
  16279=>"11111110",
  16280=>"00000001",
  16281=>"11111101",
  16282=>"00000011",
  16283=>"11111110",
  16284=>"11111101",
  16285=>"11111111",
  16286=>"11111101",
  16287=>"11111110",
  16288=>"11111110",
  16289=>"00000001",
  16290=>"00000010",
  16291=>"11111111",
  16292=>"11111110",
  16293=>"11111111",
  16294=>"00000011",
  16295=>"00000000",
  16296=>"11111110",
  16297=>"11111111",
  16298=>"00000011",
  16299=>"00000000",
  16300=>"00000000",
  16301=>"00000010",
  16302=>"00000000",
  16303=>"11111111",
  16304=>"11111111",
  16305=>"00000101",
  16306=>"00000000",
  16307=>"00000010",
  16308=>"00000010",
  16309=>"00000001",
  16310=>"00000000",
  16311=>"00000000",
  16312=>"11111011",
  16313=>"00000011",
  16314=>"00000010",
  16315=>"11111101",
  16316=>"11111110",
  16317=>"11111101",
  16318=>"11111110",
  16319=>"11111111",
  16320=>"00000010",
  16321=>"00000001",
  16322=>"00000000",
  16323=>"00000100",
  16324=>"11111111",
  16325=>"00000001",
  16326=>"00000000",
  16327=>"00000000",
  16328=>"11111101",
  16329=>"00000001",
  16330=>"11111110",
  16331=>"00000001",
  16332=>"00000000",
  16333=>"00000001",
  16334=>"00000001",
  16335=>"00000010",
  16336=>"00000001",
  16337=>"00000001",
  16338=>"00000000",
  16339=>"00000001",
  16340=>"00000000",
  16341=>"00000110",
  16342=>"11111110",
  16343=>"00000000",
  16344=>"00000010",
  16345=>"11111111",
  16346=>"00000001",
  16347=>"11111110",
  16348=>"11111110",
  16349=>"00000100",
  16350=>"00000001",
  16351=>"11111110",
  16352=>"00000001",
  16353=>"11111110",
  16354=>"11111110",
  16355=>"11111110",
  16356=>"00000010",
  16357=>"00000000",
  16358=>"00000001",
  16359=>"11111110",
  16360=>"00000011",
  16361=>"11111101",
  16362=>"00000100",
  16363=>"11111111",
  16364=>"00000101",
  16365=>"00000001",
  16366=>"11111110",
  16367=>"00000000",
  16368=>"00000000",
  16369=>"11111110",
  16370=>"11111110",
  16371=>"00000010",
  16372=>"11111100",
  16373=>"00000000",
  16374=>"11111110",
  16375=>"00000011",
  16376=>"00000001",
  16377=>"00000010",
  16378=>"11111110",
  16379=>"00000010",
  16380=>"00000001",
  16381=>"00000001",
  16382=>"11111101",
  16383=>"00000000",
  16384=>"11111100",
  16385=>"11111101",
  16386=>"00000001",
  16387=>"00000011",
  16388=>"00000000",
  16389=>"00000001",
  16390=>"11111101",
  16391=>"11111111",
  16392=>"11111111",
  16393=>"00000101",
  16394=>"00000010",
  16395=>"11111110",
  16396=>"00000000",
  16397=>"11111111",
  16398=>"00000011",
  16399=>"00000101",
  16400=>"11111101",
  16401=>"11111111",
  16402=>"00000001",
  16403=>"11111110",
  16404=>"00000100",
  16405=>"11111110",
  16406=>"11111111",
  16407=>"00000001",
  16408=>"11111101",
  16409=>"11111111",
  16410=>"00000001",
  16411=>"00000010",
  16412=>"11111101",
  16413=>"00000001",
  16414=>"11111110",
  16415=>"11111111",
  16416=>"00000001",
  16417=>"00000010",
  16418=>"11111010",
  16419=>"11111111",
  16420=>"11111101",
  16421=>"11111101",
  16422=>"00000010",
  16423=>"00000000",
  16424=>"00000100",
  16425=>"00000100",
  16426=>"00000010",
  16427=>"00000001",
  16428=>"11111110",
  16429=>"00000010",
  16430=>"00000000",
  16431=>"11111111",
  16432=>"11111110",
  16433=>"11111111",
  16434=>"00000000",
  16435=>"11111101",
  16436=>"00000000",
  16437=>"00000001",
  16438=>"00000001",
  16439=>"00000001",
  16440=>"11111101",
  16441=>"00000010",
  16442=>"00000000",
  16443=>"11111100",
  16444=>"11111110",
  16445=>"00000001",
  16446=>"11111100",
  16447=>"00000011",
  16448=>"00000000",
  16449=>"11111110",
  16450=>"11111110",
  16451=>"00000001",
  16452=>"11111101",
  16453=>"11111101",
  16454=>"11111111",
  16455=>"11111101",
  16456=>"00000010",
  16457=>"11111110",
  16458=>"00000001",
  16459=>"00000010",
  16460=>"00000100",
  16461=>"11111101",
  16462=>"11111110",
  16463=>"00000011",
  16464=>"00000000",
  16465=>"00000001",
  16466=>"00001000",
  16467=>"11111110",
  16468=>"00000001",
  16469=>"00000010",
  16470=>"00000010",
  16471=>"00000000",
  16472=>"11111100",
  16473=>"00000000",
  16474=>"00000000",
  16475=>"11111101",
  16476=>"11111110",
  16477=>"11111111",
  16478=>"00000011",
  16479=>"00000010",
  16480=>"00000001",
  16481=>"11111110",
  16482=>"00000000",
  16483=>"00000010",
  16484=>"11111100",
  16485=>"00000010",
  16486=>"11111101",
  16487=>"00000011",
  16488=>"00000001",
  16489=>"00000010",
  16490=>"00000110",
  16491=>"00000001",
  16492=>"11111111",
  16493=>"11111110",
  16494=>"00000001",
  16495=>"00000101",
  16496=>"11111100",
  16497=>"00000001",
  16498=>"11111110",
  16499=>"00000000",
  16500=>"11111110",
  16501=>"00000001",
  16502=>"11111100",
  16503=>"11111110",
  16504=>"00000010",
  16505=>"00000001",
  16506=>"11111111",
  16507=>"00000010",
  16508=>"11111111",
  16509=>"00000000",
  16510=>"00000000",
  16511=>"11111101",
  16512=>"00000000",
  16513=>"11111100",
  16514=>"11111110",
  16515=>"00000000",
  16516=>"00000001",
  16517=>"11111111",
  16518=>"00000000",
  16519=>"00000001",
  16520=>"11111110",
  16521=>"11111111",
  16522=>"11111110",
  16523=>"00000001",
  16524=>"11111111",
  16525=>"11111101",
  16526=>"00000000",
  16527=>"00000010",
  16528=>"00000010",
  16529=>"00000011",
  16530=>"11111101",
  16531=>"11111101",
  16532=>"00000010",
  16533=>"11111110",
  16534=>"11111111",
  16535=>"00000000",
  16536=>"11111101",
  16537=>"00000011",
  16538=>"11111110",
  16539=>"11111111",
  16540=>"11111110",
  16541=>"00000001",
  16542=>"00000000",
  16543=>"11111111",
  16544=>"00000010",
  16545=>"00000010",
  16546=>"11111110",
  16547=>"00000001",
  16548=>"11111111",
  16549=>"00000000",
  16550=>"11111110",
  16551=>"00000001",
  16552=>"00000010",
  16553=>"00000010",
  16554=>"11111111",
  16555=>"00000010",
  16556=>"00000010",
  16557=>"00000010",
  16558=>"00000011",
  16559=>"00000000",
  16560=>"11111111",
  16561=>"11111110",
  16562=>"00000000",
  16563=>"00000000",
  16564=>"11111111",
  16565=>"11111100",
  16566=>"00000011",
  16567=>"11111110",
  16568=>"00000011",
  16569=>"11111110",
  16570=>"00000010",
  16571=>"11111110",
  16572=>"11111101",
  16573=>"00000000",
  16574=>"00000000",
  16575=>"00000100",
  16576=>"00000000",
  16577=>"00000010",
  16578=>"11111111",
  16579=>"00000011",
  16580=>"11111110",
  16581=>"00000010",
  16582=>"11111111",
  16583=>"11111101",
  16584=>"00000100",
  16585=>"00000010",
  16586=>"00000000",
  16587=>"00000000",
  16588=>"11111111",
  16589=>"00000000",
  16590=>"11111100",
  16591=>"00000100",
  16592=>"00000000",
  16593=>"00000010",
  16594=>"11111111",
  16595=>"00000010",
  16596=>"00000010",
  16597=>"11111111",
  16598=>"11111111",
  16599=>"00000011",
  16600=>"00000001",
  16601=>"11111101",
  16602=>"00000001",
  16603=>"00000001",
  16604=>"00000010",
  16605=>"11111111",
  16606=>"11111111",
  16607=>"11111110",
  16608=>"11111101",
  16609=>"00000011",
  16610=>"11111100",
  16611=>"11111110",
  16612=>"00000010",
  16613=>"00000000",
  16614=>"11111110",
  16615=>"11111111",
  16616=>"11111111",
  16617=>"00000100",
  16618=>"00000011",
  16619=>"00000001",
  16620=>"11111111",
  16621=>"11111100",
  16622=>"00000000",
  16623=>"11111101",
  16624=>"00000100",
  16625=>"11111101",
  16626=>"00000010",
  16627=>"00000000",
  16628=>"00000000",
  16629=>"00000011",
  16630=>"11111111",
  16631=>"11111110",
  16632=>"11111111",
  16633=>"11111100",
  16634=>"00000001",
  16635=>"11111101",
  16636=>"11111111",
  16637=>"00000000",
  16638=>"11111111",
  16639=>"11111111",
  16640=>"11111100",
  16641=>"11111111",
  16642=>"00000000",
  16643=>"00000001",
  16644=>"00000010",
  16645=>"00000010",
  16646=>"00000001",
  16647=>"11111110",
  16648=>"00000010",
  16649=>"11111111",
  16650=>"11111010",
  16651=>"11111101",
  16652=>"00000000",
  16653=>"00000010",
  16654=>"11111101",
  16655=>"11111110",
  16656=>"00000011",
  16657=>"11111101",
  16658=>"00000011",
  16659=>"00000000",
  16660=>"11111110",
  16661=>"11111111",
  16662=>"00000000",
  16663=>"00000001",
  16664=>"11111110",
  16665=>"00000000",
  16666=>"00000010",
  16667=>"00000000",
  16668=>"00000000",
  16669=>"11111101",
  16670=>"00000011",
  16671=>"00000000",
  16672=>"11111110",
  16673=>"00000000",
  16674=>"00000001",
  16675=>"11111110",
  16676=>"11111111",
  16677=>"11111111",
  16678=>"00000000",
  16679=>"11111101",
  16680=>"00000010",
  16681=>"11111111",
  16682=>"11111110",
  16683=>"11111111",
  16684=>"11111110",
  16685=>"11111111",
  16686=>"00000000",
  16687=>"11111100",
  16688=>"00000001",
  16689=>"00000000",
  16690=>"00000000",
  16691=>"11111110",
  16692=>"00000010",
  16693=>"00000001",
  16694=>"00000001",
  16695=>"11111100",
  16696=>"00000011",
  16697=>"00000001",
  16698=>"00000001",
  16699=>"11111111",
  16700=>"00000100",
  16701=>"11111111",
  16702=>"11111110",
  16703=>"11111110",
  16704=>"11111101",
  16705=>"00000101",
  16706=>"00000000",
  16707=>"11111110",
  16708=>"11111101",
  16709=>"00000010",
  16710=>"00000001",
  16711=>"00000001",
  16712=>"11111111",
  16713=>"00000011",
  16714=>"00000011",
  16715=>"00000000",
  16716=>"00000001",
  16717=>"11111111",
  16718=>"00000010",
  16719=>"00000001",
  16720=>"11111011",
  16721=>"11111111",
  16722=>"11111110",
  16723=>"00000101",
  16724=>"00000011",
  16725=>"11111101",
  16726=>"00000100",
  16727=>"00000111",
  16728=>"00000001",
  16729=>"11111111",
  16730=>"11111111",
  16731=>"00000001",
  16732=>"11111101",
  16733=>"11111111",
  16734=>"00000010",
  16735=>"11111101",
  16736=>"00000000",
  16737=>"11111110",
  16738=>"00000000",
  16739=>"00000001",
  16740=>"00000010",
  16741=>"11111110",
  16742=>"00000000",
  16743=>"11111110",
  16744=>"00000000",
  16745=>"11111110",
  16746=>"00000001",
  16747=>"00000100",
  16748=>"00000011",
  16749=>"00000000",
  16750=>"00000011",
  16751=>"00000001",
  16752=>"11111101",
  16753=>"11111101",
  16754=>"00000001",
  16755=>"11111101",
  16756=>"11111100",
  16757=>"00000000",
  16758=>"00000011",
  16759=>"00000010",
  16760=>"00000101",
  16761=>"11111110",
  16762=>"11111110",
  16763=>"00000011",
  16764=>"00000001",
  16765=>"00000011",
  16766=>"11111011",
  16767=>"11111101",
  16768=>"11111100",
  16769=>"00000010",
  16770=>"00000000",
  16771=>"00000010",
  16772=>"00000010",
  16773=>"00000010",
  16774=>"11111101",
  16775=>"00000010",
  16776=>"11111101",
  16777=>"00000001",
  16778=>"00000000",
  16779=>"00000001",
  16780=>"11111110",
  16781=>"11111111",
  16782=>"00000010",
  16783=>"00000000",
  16784=>"00000000",
  16785=>"11111111",
  16786=>"11111111",
  16787=>"00000000",
  16788=>"00000110",
  16789=>"00000000",
  16790=>"11111111",
  16791=>"00000111",
  16792=>"00000000",
  16793=>"00000010",
  16794=>"00000011",
  16795=>"00000100",
  16796=>"00000011",
  16797=>"00000011",
  16798=>"00000011",
  16799=>"00000000",
  16800=>"11111111",
  16801=>"11111111",
  16802=>"00000000",
  16803=>"11111101",
  16804=>"11111110",
  16805=>"00000100",
  16806=>"11111101",
  16807=>"00000001",
  16808=>"00000000",
  16809=>"00000010",
  16810=>"11111111",
  16811=>"00000010",
  16812=>"11111101",
  16813=>"11111110",
  16814=>"11111110",
  16815=>"00000001",
  16816=>"00000000",
  16817=>"11111111",
  16818=>"11111110",
  16819=>"00000001",
  16820=>"00000010",
  16821=>"00000001",
  16822=>"00000001",
  16823=>"00000011",
  16824=>"11111111",
  16825=>"11111111",
  16826=>"00000011",
  16827=>"11111101",
  16828=>"11111110",
  16829=>"00000010",
  16830=>"00000011",
  16831=>"00000000",
  16832=>"11111111",
  16833=>"00000001",
  16834=>"00000101",
  16835=>"00000001",
  16836=>"11111101",
  16837=>"00000100",
  16838=>"11111110",
  16839=>"00000100",
  16840=>"00000001",
  16841=>"00000000",
  16842=>"00000000",
  16843=>"00000010",
  16844=>"00000010",
  16845=>"00000001",
  16846=>"00000001",
  16847=>"11111111",
  16848=>"11111110",
  16849=>"00000001",
  16850=>"11111110",
  16851=>"00000001",
  16852=>"11111111",
  16853=>"00000000",
  16854=>"00000010",
  16855=>"00000001",
  16856=>"00000010",
  16857=>"00000010",
  16858=>"00000010",
  16859=>"11111101",
  16860=>"00000000",
  16861=>"00000000",
  16862=>"00000001",
  16863=>"11111100",
  16864=>"11111110",
  16865=>"00000001",
  16866=>"00000001",
  16867=>"11111111",
  16868=>"00000001",
  16869=>"00000101",
  16870=>"11111101",
  16871=>"11111110",
  16872=>"00000100",
  16873=>"00000001",
  16874=>"11111110",
  16875=>"11111111",
  16876=>"11111111",
  16877=>"00000000",
  16878=>"00000000",
  16879=>"00000000",
  16880=>"11111111",
  16881=>"00000010",
  16882=>"11111110",
  16883=>"00000010",
  16884=>"11111111",
  16885=>"11111101",
  16886=>"11111111",
  16887=>"11111111",
  16888=>"00000001",
  16889=>"11111110",
  16890=>"00000000",
  16891=>"11111111",
  16892=>"00000100",
  16893=>"11111101",
  16894=>"11111110",
  16895=>"11111110",
  16896=>"00000001",
  16897=>"11111100",
  16898=>"00000001",
  16899=>"11111110",
  16900=>"11111100",
  16901=>"00000000",
  16902=>"11111111",
  16903=>"00000000",
  16904=>"11111101",
  16905=>"11111110",
  16906=>"00000001",
  16907=>"11111111",
  16908=>"11111101",
  16909=>"00000000",
  16910=>"00000011",
  16911=>"00000000",
  16912=>"11111110",
  16913=>"11111100",
  16914=>"11111110",
  16915=>"00000011",
  16916=>"11111100",
  16917=>"00000000",
  16918=>"11111101",
  16919=>"00000010",
  16920=>"00000011",
  16921=>"11111111",
  16922=>"11111110",
  16923=>"00000010",
  16924=>"00000000",
  16925=>"00000001",
  16926=>"00000001",
  16927=>"11111111",
  16928=>"00000010",
  16929=>"11111110",
  16930=>"00000001",
  16931=>"00000011",
  16932=>"00000010",
  16933=>"11111110",
  16934=>"11111111",
  16935=>"00000010",
  16936=>"00000001",
  16937=>"11111101",
  16938=>"11111111",
  16939=>"00000000",
  16940=>"00000011",
  16941=>"00000011",
  16942=>"11111110",
  16943=>"00000011",
  16944=>"00000011",
  16945=>"11111110",
  16946=>"00000001",
  16947=>"11111101",
  16948=>"11111101",
  16949=>"00000000",
  16950=>"00000101",
  16951=>"00000001",
  16952=>"11111111",
  16953=>"11111101",
  16954=>"00000010",
  16955=>"00000011",
  16956=>"00000010",
  16957=>"00000001",
  16958=>"11111110",
  16959=>"11111111",
  16960=>"11111110",
  16961=>"00000101",
  16962=>"11111101",
  16963=>"00000010",
  16964=>"11111110",
  16965=>"11111111",
  16966=>"00000001",
  16967=>"00000001",
  16968=>"00000000",
  16969=>"00000011",
  16970=>"00000001",
  16971=>"11111110",
  16972=>"00000011",
  16973=>"00000010",
  16974=>"11111110",
  16975=>"00000010",
  16976=>"11111110",
  16977=>"00000011",
  16978=>"00000011",
  16979=>"11111111",
  16980=>"00000000",
  16981=>"00000011",
  16982=>"11111111",
  16983=>"11111111",
  16984=>"00000011",
  16985=>"11111101",
  16986=>"11111111",
  16987=>"00000001",
  16988=>"11111101",
  16989=>"00000000",
  16990=>"11111110",
  16991=>"11111110",
  16992=>"00000001",
  16993=>"11111111",
  16994=>"00000011",
  16995=>"00000001",
  16996=>"00000001",
  16997=>"00000001",
  16998=>"00000001",
  16999=>"00000000",
  17000=>"11111111",
  17001=>"11111110",
  17002=>"00000000",
  17003=>"11111110",
  17004=>"11111100",
  17005=>"00000110",
  17006=>"11111101",
  17007=>"00000000",
  17008=>"00000010",
  17009=>"11111101",
  17010=>"00000010",
  17011=>"11111101",
  17012=>"00000011",
  17013=>"11111110",
  17014=>"00000010",
  17015=>"00000111",
  17016=>"11111111",
  17017=>"11111110",
  17018=>"11111111",
  17019=>"00000000",
  17020=>"00000010",
  17021=>"00000000",
  17022=>"00000100",
  17023=>"11111110",
  17024=>"11111100",
  17025=>"00000000",
  17026=>"11111100",
  17027=>"00000011",
  17028=>"11111110",
  17029=>"00000100",
  17030=>"11111110",
  17031=>"00000011",
  17032=>"00000011",
  17033=>"11111101",
  17034=>"11111101",
  17035=>"11111111",
  17036=>"00000010",
  17037=>"11111111",
  17038=>"00000010",
  17039=>"00000001",
  17040=>"11111110",
  17041=>"00000010",
  17042=>"00000001",
  17043=>"11111111",
  17044=>"11111110",
  17045=>"00000010",
  17046=>"11111110",
  17047=>"00000001",
  17048=>"00000011",
  17049=>"00000011",
  17050=>"11111110",
  17051=>"00000000",
  17052=>"00000000",
  17053=>"00000010",
  17054=>"00000100",
  17055=>"11111110",
  17056=>"00000001",
  17057=>"11111101",
  17058=>"11111110",
  17059=>"00000010",
  17060=>"00000010",
  17061=>"00000001",
  17062=>"00000010",
  17063=>"00000010",
  17064=>"00000001",
  17065=>"11111101",
  17066=>"00000100",
  17067=>"00000000",
  17068=>"00000000",
  17069=>"00000010",
  17070=>"11111101",
  17071=>"00000110",
  17072=>"00000000",
  17073=>"00000011",
  17074=>"11111110",
  17075=>"00000001",
  17076=>"11111110",
  17077=>"11111111",
  17078=>"11111110",
  17079=>"11111101",
  17080=>"11111101",
  17081=>"00000000",
  17082=>"00000010",
  17083=>"11111111",
  17084=>"00000000",
  17085=>"00000001",
  17086=>"00000010",
  17087=>"11111110",
  17088=>"00000010",
  17089=>"11111111",
  17090=>"11111101",
  17091=>"00000001",
  17092=>"00000001",
  17093=>"00000010",
  17094=>"11111111",
  17095=>"11111111",
  17096=>"00000010",
  17097=>"11111110",
  17098=>"00000011",
  17099=>"11111111",
  17100=>"11111100",
  17101=>"00000011",
  17102=>"11111111",
  17103=>"11111111",
  17104=>"00000000",
  17105=>"00000000",
  17106=>"11111110",
  17107=>"00000111",
  17108=>"11111110",
  17109=>"00000001",
  17110=>"11111100",
  17111=>"11111111",
  17112=>"11111110",
  17113=>"00000010",
  17114=>"00000001",
  17115=>"00000000",
  17116=>"11111111",
  17117=>"00000000",
  17118=>"00000010",
  17119=>"11111110",
  17120=>"00000011",
  17121=>"00000010",
  17122=>"00000011",
  17123=>"00000000",
  17124=>"00000010",
  17125=>"11111110",
  17126=>"00000100",
  17127=>"00000010",
  17128=>"00000000",
  17129=>"00000010",
  17130=>"11111110",
  17131=>"11111111",
  17132=>"00000001",
  17133=>"00000000",
  17134=>"11111101",
  17135=>"00000001",
  17136=>"11111101",
  17137=>"11111110",
  17138=>"11111110",
  17139=>"11111110",
  17140=>"00000011",
  17141=>"11111110",
  17142=>"00000000",
  17143=>"00000011",
  17144=>"00000011",
  17145=>"11111111",
  17146=>"11111111",
  17147=>"11111111",
  17148=>"00000100",
  17149=>"11111101",
  17150=>"00000010",
  17151=>"00000011",
  17152=>"11111110",
  17153=>"00000000",
  17154=>"00000001",
  17155=>"11111101",
  17156=>"00000001",
  17157=>"11111111",
  17158=>"00000010",
  17159=>"11111101",
  17160=>"11111110",
  17161=>"11111110",
  17162=>"00000001",
  17163=>"00000100",
  17164=>"00000010",
  17165=>"11111111",
  17166=>"11111100",
  17167=>"00000010",
  17168=>"00000001",
  17169=>"11111111",
  17170=>"11111100",
  17171=>"11111110",
  17172=>"00000000",
  17173=>"00000000",
  17174=>"11111111",
  17175=>"00000001",
  17176=>"00000001",
  17177=>"00000100",
  17178=>"00000100",
  17179=>"00000010",
  17180=>"11111110",
  17181=>"00000010",
  17182=>"00000000",
  17183=>"11111111",
  17184=>"11111110",
  17185=>"11111100",
  17186=>"00000001",
  17187=>"00000101",
  17188=>"11111111",
  17189=>"00000000",
  17190=>"00000001",
  17191=>"00000010",
  17192=>"00000010",
  17193=>"11111110",
  17194=>"00000000",
  17195=>"00000000",
  17196=>"00000001",
  17197=>"00000011",
  17198=>"11111101",
  17199=>"11111111",
  17200=>"11111101",
  17201=>"11111111",
  17202=>"00000001",
  17203=>"00000001",
  17204=>"00000010",
  17205=>"11111101",
  17206=>"11111101",
  17207=>"00000010",
  17208=>"00000001",
  17209=>"11111100",
  17210=>"11111111",
  17211=>"00000011",
  17212=>"00000010",
  17213=>"00000100",
  17214=>"11111111",
  17215=>"00000010",
  17216=>"11111101",
  17217=>"11111100",
  17218=>"00000001",
  17219=>"00000001",
  17220=>"00000000",
  17221=>"11111111",
  17222=>"11111101",
  17223=>"11111110",
  17224=>"00000001",
  17225=>"00000001",
  17226=>"00000011",
  17227=>"11111110",
  17228=>"11111111",
  17229=>"11111110",
  17230=>"00000001",
  17231=>"00000000",
  17232=>"11111110",
  17233=>"11111111",
  17234=>"11111101",
  17235=>"11111101",
  17236=>"11111111",
  17237=>"11111110",
  17238=>"00000001",
  17239=>"11111110",
  17240=>"11111110",
  17241=>"11111101",
  17242=>"11111111",
  17243=>"00000100",
  17244=>"11111101",
  17245=>"00000010",
  17246=>"00000010",
  17247=>"11111110",
  17248=>"00000001",
  17249=>"11111110",
  17250=>"00000000",
  17251=>"11111111",
  17252=>"11111111",
  17253=>"00000001",
  17254=>"00000000",
  17255=>"11111101",
  17256=>"00000000",
  17257=>"11111110",
  17258=>"11111111",
  17259=>"00000101",
  17260=>"00000000",
  17261=>"11111110",
  17262=>"11111111",
  17263=>"00000010",
  17264=>"00000001",
  17265=>"11111110",
  17266=>"00000011",
  17267=>"11111101",
  17268=>"00000000",
  17269=>"00000010",
  17270=>"11111110",
  17271=>"00000001",
  17272=>"00000011",
  17273=>"00000000",
  17274=>"00000010",
  17275=>"11111110",
  17276=>"11111011",
  17277=>"11111111",
  17278=>"11111101",
  17279=>"00000011",
  17280=>"00000001",
  17281=>"00000001",
  17282=>"00000011",
  17283=>"11111101",
  17284=>"00000000",
  17285=>"00000000",
  17286=>"11111110",
  17287=>"11111110",
  17288=>"00000011",
  17289=>"00000011",
  17290=>"11111101",
  17291=>"00000001",
  17292=>"00000001",
  17293=>"00000001",
  17294=>"11111110",
  17295=>"11111111",
  17296=>"00000100",
  17297=>"11111101",
  17298=>"00000010",
  17299=>"11111111",
  17300=>"00000010",
  17301=>"00000001",
  17302=>"11111110",
  17303=>"00000000",
  17304=>"11111111",
  17305=>"00000100",
  17306=>"00000010",
  17307=>"00000011",
  17308=>"11111101",
  17309=>"11111101",
  17310=>"11111110",
  17311=>"00000011",
  17312=>"00000011",
  17313=>"11111101",
  17314=>"11111110",
  17315=>"00000001",
  17316=>"00000001",
  17317=>"11111111",
  17318=>"00000010",
  17319=>"00000000",
  17320=>"11111110",
  17321=>"00000011",
  17322=>"11111101",
  17323=>"11111101",
  17324=>"00000000",
  17325=>"11111110",
  17326=>"00000000",
  17327=>"11111111",
  17328=>"11111110",
  17329=>"11111110",
  17330=>"00000011",
  17331=>"11111101",
  17332=>"00000001",
  17333=>"11111101",
  17334=>"00000010",
  17335=>"11111110",
  17336=>"11111101",
  17337=>"00000001",
  17338=>"11111111",
  17339=>"11111101",
  17340=>"00000000",
  17341=>"00000001",
  17342=>"11111101",
  17343=>"00000010",
  17344=>"00000100",
  17345=>"11111100",
  17346=>"11111110",
  17347=>"00000001",
  17348=>"00000000",
  17349=>"11111110",
  17350=>"11111111",
  17351=>"00000000",
  17352=>"11111110",
  17353=>"11111111",
  17354=>"00000010",
  17355=>"11111111",
  17356=>"11111111",
  17357=>"11111111",
  17358=>"00000010",
  17359=>"00000011",
  17360=>"11111111",
  17361=>"00000001",
  17362=>"11111100",
  17363=>"11111110",
  17364=>"00000010",
  17365=>"00000011",
  17366=>"11111110",
  17367=>"11111101",
  17368=>"00000000",
  17369=>"00000001",
  17370=>"11111110",
  17371=>"11111110",
  17372=>"11111110",
  17373=>"11111110",
  17374=>"11111100",
  17375=>"11111100",
  17376=>"11111111",
  17377=>"11111110",
  17378=>"00000000",
  17379=>"00000010",
  17380=>"00000000",
  17381=>"00000101",
  17382=>"00000001",
  17383=>"11111111",
  17384=>"11111101",
  17385=>"11111111",
  17386=>"11111100",
  17387=>"00000100",
  17388=>"00000001",
  17389=>"00000011",
  17390=>"00000000",
  17391=>"11111110",
  17392=>"00000001",
  17393=>"00000000",
  17394=>"11111110",
  17395=>"00000100",
  17396=>"11111110",
  17397=>"00000001",
  17398=>"00000000",
  17399=>"11111110",
  17400=>"11111101",
  17401=>"00000001",
  17402=>"00000001",
  17403=>"00000000",
  17404=>"11111110",
  17405=>"11111111",
  17406=>"00000000",
  17407=>"00000000",
  17408=>"00000010",
  17409=>"11111110",
  17410=>"00000000",
  17411=>"11111101",
  17412=>"11111101",
  17413=>"00000010",
  17414=>"00000001",
  17415=>"11111101",
  17416=>"11111110",
  17417=>"00000001",
  17418=>"00000011",
  17419=>"11111101",
  17420=>"00000000",
  17421=>"00000000",
  17422=>"11111110",
  17423=>"00000000",
  17424=>"11111110",
  17425=>"00000010",
  17426=>"00000101",
  17427=>"00000000",
  17428=>"11111110",
  17429=>"00000000",
  17430=>"00000010",
  17431=>"00000001",
  17432=>"00000000",
  17433=>"11111101",
  17434=>"11111101",
  17435=>"00000001",
  17436=>"00000010",
  17437=>"00000000",
  17438=>"11111111",
  17439=>"11111110",
  17440=>"00000100",
  17441=>"00000010",
  17442=>"11111101",
  17443=>"11111100",
  17444=>"00000000",
  17445=>"00000010",
  17446=>"11111111",
  17447=>"00000010",
  17448=>"00000001",
  17449=>"11111111",
  17450=>"11111101",
  17451=>"11111101",
  17452=>"00000001",
  17453=>"11111111",
  17454=>"11111111",
  17455=>"11111110",
  17456=>"11111101",
  17457=>"11111111",
  17458=>"00000001",
  17459=>"11111110",
  17460=>"11111101",
  17461=>"11111111",
  17462=>"00000010",
  17463=>"00000001",
  17464=>"00000000",
  17465=>"00000001",
  17466=>"11111110",
  17467=>"11111100",
  17468=>"00000000",
  17469=>"00000000",
  17470=>"11111110",
  17471=>"00000000",
  17472=>"00000001",
  17473=>"00000000",
  17474=>"00000000",
  17475=>"11111101",
  17476=>"00000001",
  17477=>"00000010",
  17478=>"00000010",
  17479=>"11111110",
  17480=>"11111101",
  17481=>"00000000",
  17482=>"11111111",
  17483=>"11111101",
  17484=>"11111111",
  17485=>"00000010",
  17486=>"11111110",
  17487=>"00000000",
  17488=>"11111111",
  17489=>"00000010",
  17490=>"00000001",
  17491=>"11111110",
  17492=>"11111110",
  17493=>"00000001",
  17494=>"00000001",
  17495=>"00000010",
  17496=>"11111110",
  17497=>"11111101",
  17498=>"00000010",
  17499=>"11111100",
  17500=>"00000001",
  17501=>"11111101",
  17502=>"11111111",
  17503=>"11111110",
  17504=>"00000000",
  17505=>"11111110",
  17506=>"11111110",
  17507=>"11111101",
  17508=>"00000001",
  17509=>"11111111",
  17510=>"11111111",
  17511=>"11111110",
  17512=>"11111111",
  17513=>"00000000",
  17514=>"11111111",
  17515=>"00000101",
  17516=>"11111111",
  17517=>"00000000",
  17518=>"11111101",
  17519=>"00000010",
  17520=>"11111111",
  17521=>"00000000",
  17522=>"00000001",
  17523=>"00000001",
  17524=>"11111110",
  17525=>"00000010",
  17526=>"11111111",
  17527=>"00000100",
  17528=>"00000011",
  17529=>"11111110",
  17530=>"11111111",
  17531=>"00000011",
  17532=>"11111111",
  17533=>"11111110",
  17534=>"11111110",
  17535=>"11111111",
  17536=>"11111110",
  17537=>"00000001",
  17538=>"11111110",
  17539=>"11111111",
  17540=>"00000011",
  17541=>"00000001",
  17542=>"00000000",
  17543=>"11111111",
  17544=>"11111110",
  17545=>"00000001",
  17546=>"00000011",
  17547=>"00000010",
  17548=>"00000010",
  17549=>"11111101",
  17550=>"11111111",
  17551=>"11111101",
  17552=>"00000010",
  17553=>"11111110",
  17554=>"00000001",
  17555=>"00000100",
  17556=>"11111100",
  17557=>"00000011",
  17558=>"00000000",
  17559=>"11111101",
  17560=>"11111110",
  17561=>"11111110",
  17562=>"00000100",
  17563=>"00000010",
  17564=>"11111111",
  17565=>"11111101",
  17566=>"00000001",
  17567=>"00000000",
  17568=>"11111111",
  17569=>"11111100",
  17570=>"00000010",
  17571=>"11111111",
  17572=>"00000001",
  17573=>"11111111",
  17574=>"00000001",
  17575=>"11111101",
  17576=>"11111101",
  17577=>"00000000",
  17578=>"00000010",
  17579=>"11111100",
  17580=>"00000011",
  17581=>"11111111",
  17582=>"11111101",
  17583=>"00000000",
  17584=>"00000001",
  17585=>"00000001",
  17586=>"00000000",
  17587=>"00000000",
  17588=>"00000001",
  17589=>"11111110",
  17590=>"00000000",
  17591=>"11111110",
  17592=>"11111110",
  17593=>"00000000",
  17594=>"00000000",
  17595=>"00000001",
  17596=>"00000011",
  17597=>"11111111",
  17598=>"11111111",
  17599=>"11111110",
  17600=>"00000000",
  17601=>"11111111",
  17602=>"00000010",
  17603=>"11111101",
  17604=>"00000001",
  17605=>"11111111",
  17606=>"11111101",
  17607=>"00000010",
  17608=>"11111111",
  17609=>"11111101",
  17610=>"00000011",
  17611=>"00000011",
  17612=>"11111101",
  17613=>"11111101",
  17614=>"00000000",
  17615=>"00000010",
  17616=>"00000100",
  17617=>"00000110",
  17618=>"11111110",
  17619=>"00000010",
  17620=>"00000010",
  17621=>"00000111",
  17622=>"00000001",
  17623=>"11111110",
  17624=>"00000000",
  17625=>"11111111",
  17626=>"00000011",
  17627=>"11111111",
  17628=>"00000001",
  17629=>"11111110",
  17630=>"00000011",
  17631=>"11111110",
  17632=>"00000001",
  17633=>"11111110",
  17634=>"00000001",
  17635=>"11111111",
  17636=>"00000001",
  17637=>"00000000",
  17638=>"11111111",
  17639=>"11111101",
  17640=>"00000001",
  17641=>"11111110",
  17642=>"00000010",
  17643=>"00000010",
  17644=>"00000000",
  17645=>"11111101",
  17646=>"00000001",
  17647=>"00000000",
  17648=>"11111101",
  17649=>"11111101",
  17650=>"11111110",
  17651=>"11111100",
  17652=>"11111101",
  17653=>"11111101",
  17654=>"11111111",
  17655=>"00000001",
  17656=>"00000000",
  17657=>"11111111",
  17658=>"00000001",
  17659=>"11111111",
  17660=>"00000000",
  17661=>"11111110",
  17662=>"00000000",
  17663=>"11111101",
  17664=>"00000000",
  17665=>"11111101",
  17666=>"00000010",
  17667=>"11111110",
  17668=>"00000001",
  17669=>"00000010",
  17670=>"00000010",
  17671=>"00000001",
  17672=>"11111101",
  17673=>"00000000",
  17674=>"00000101",
  17675=>"00000000",
  17676=>"00000010",
  17677=>"00000000",
  17678=>"11111100",
  17679=>"00000110",
  17680=>"11111111",
  17681=>"11111110",
  17682=>"11111100",
  17683=>"00000010",
  17684=>"11111110",
  17685=>"11111101",
  17686=>"11111100",
  17687=>"00000000",
  17688=>"11111111",
  17689=>"00000100",
  17690=>"11111101",
  17691=>"11111101",
  17692=>"11111101",
  17693=>"00000001",
  17694=>"11111110",
  17695=>"00000001",
  17696=>"00000010",
  17697=>"00000000",
  17698=>"11111110",
  17699=>"00000010",
  17700=>"11111111",
  17701=>"00000001",
  17702=>"00000000",
  17703=>"11111111",
  17704=>"11111100",
  17705=>"11111110",
  17706=>"11111101",
  17707=>"00000011",
  17708=>"11111111",
  17709=>"11111101",
  17710=>"00000011",
  17711=>"00000100",
  17712=>"11111111",
  17713=>"11111101",
  17714=>"11111111",
  17715=>"00000000",
  17716=>"11111111",
  17717=>"11111111",
  17718=>"11111110",
  17719=>"00000100",
  17720=>"11111110",
  17721=>"11111101",
  17722=>"00000100",
  17723=>"11111111",
  17724=>"00000010",
  17725=>"11111101",
  17726=>"11111101",
  17727=>"00000001",
  17728=>"00000000",
  17729=>"00000000",
  17730=>"11111111",
  17731=>"11111101",
  17732=>"00000010",
  17733=>"00000010",
  17734=>"00000011",
  17735=>"11111110",
  17736=>"00000010",
  17737=>"00000100",
  17738=>"11111011",
  17739=>"11111111",
  17740=>"00000010",
  17741=>"00000010",
  17742=>"11111110",
  17743=>"11111101",
  17744=>"00000110",
  17745=>"00000011",
  17746=>"00000000",
  17747=>"11111110",
  17748=>"11111111",
  17749=>"00000011",
  17750=>"11111111",
  17751=>"00000011",
  17752=>"11111110",
  17753=>"11111110",
  17754=>"00000010",
  17755=>"11111101",
  17756=>"11111111",
  17757=>"00000011",
  17758=>"00000010",
  17759=>"00000011",
  17760=>"11111101",
  17761=>"11111111",
  17762=>"11111101",
  17763=>"11111100",
  17764=>"11111111",
  17765=>"00000000",
  17766=>"11111110",
  17767=>"11111110",
  17768=>"11111110",
  17769=>"11111101",
  17770=>"00000001",
  17771=>"00000100",
  17772=>"11111110",
  17773=>"11111110",
  17774=>"11111101",
  17775=>"11111101",
  17776=>"00000010",
  17777=>"00000000",
  17778=>"11111111",
  17779=>"11111110",
  17780=>"00000011",
  17781=>"00000000",
  17782=>"00000011",
  17783=>"00000010",
  17784=>"11111101",
  17785=>"00000101",
  17786=>"11111110",
  17787=>"11111111",
  17788=>"00000001",
  17789=>"11111110",
  17790=>"11111111",
  17791=>"00000100",
  17792=>"00000000",
  17793=>"11111110",
  17794=>"00000010",
  17795=>"00000001",
  17796=>"11111101",
  17797=>"11111101",
  17798=>"11111100",
  17799=>"11111111",
  17800=>"11111101",
  17801=>"00000001",
  17802=>"11111111",
  17803=>"11111111",
  17804=>"00000011",
  17805=>"11111110",
  17806=>"11111110",
  17807=>"00000000",
  17808=>"11111101",
  17809=>"00000001",
  17810=>"11111110",
  17811=>"00000000",
  17812=>"11111111",
  17813=>"00000001",
  17814=>"00000000",
  17815=>"11111111",
  17816=>"00000000",
  17817=>"00000101",
  17818=>"00000001",
  17819=>"11111110",
  17820=>"00000111",
  17821=>"11111111",
  17822=>"11111101",
  17823=>"00000000",
  17824=>"00000010",
  17825=>"11111101",
  17826=>"11111110",
  17827=>"00000000",
  17828=>"00000000",
  17829=>"00000011",
  17830=>"11111110",
  17831=>"11111111",
  17832=>"11111101",
  17833=>"00000000",
  17834=>"00000000",
  17835=>"00000001",
  17836=>"00000000",
  17837=>"00000011",
  17838=>"00000001",
  17839=>"00000000",
  17840=>"00000000",
  17841=>"00000000",
  17842=>"11111111",
  17843=>"11111101",
  17844=>"11111111",
  17845=>"00000111",
  17846=>"00000000",
  17847=>"11111101",
  17848=>"00000001",
  17849=>"00000000",
  17850=>"00000001",
  17851=>"11111111",
  17852=>"00000010",
  17853=>"00000011",
  17854=>"00000100",
  17855=>"00000001",
  17856=>"11111110",
  17857=>"11111111",
  17858=>"00000010",
  17859=>"11111111",
  17860=>"00000000",
  17861=>"00000000",
  17862=>"00000100",
  17863=>"00000000",
  17864=>"00000001",
  17865=>"00000000",
  17866=>"00000000",
  17867=>"00000000",
  17868=>"11111110",
  17869=>"11111111",
  17870=>"11111110",
  17871=>"00000010",
  17872=>"11111110",
  17873=>"00000000",
  17874=>"00000001",
  17875=>"00000001",
  17876=>"11111111",
  17877=>"11111111",
  17878=>"00000011",
  17879=>"11111110",
  17880=>"00000010",
  17881=>"11111111",
  17882=>"00000000",
  17883=>"00000011",
  17884=>"11111110",
  17885=>"00000001",
  17886=>"11111111",
  17887=>"00000001",
  17888=>"00000000",
  17889=>"00000000",
  17890=>"11111101",
  17891=>"11111110",
  17892=>"11111110",
  17893=>"00000110",
  17894=>"00000001",
  17895=>"11111110",
  17896=>"11111111",
  17897=>"00000000",
  17898=>"00000010",
  17899=>"00000000",
  17900=>"00000010",
  17901=>"00000011",
  17902=>"11111111",
  17903=>"00000101",
  17904=>"00000000",
  17905=>"11111110",
  17906=>"00000000",
  17907=>"11111100",
  17908=>"00000010",
  17909=>"11111110",
  17910=>"11111110",
  17911=>"00000000",
  17912=>"00000001",
  17913=>"00000011",
  17914=>"00000000",
  17915=>"11111100",
  17916=>"11111111",
  17917=>"00000110",
  17918=>"00000001",
  17919=>"00000101",
  17920=>"00000001",
  17921=>"00000010",
  17922=>"11111101",
  17923=>"11111101",
  17924=>"00000010",
  17925=>"11111100",
  17926=>"11111111",
  17927=>"11111110",
  17928=>"00000000",
  17929=>"00000110",
  17930=>"00000010",
  17931=>"11111110",
  17932=>"00000011",
  17933=>"00000000",
  17934=>"11111101",
  17935=>"11111111",
  17936=>"00000011",
  17937=>"00000011",
  17938=>"11111110",
  17939=>"00000010",
  17940=>"00000001",
  17941=>"00000001",
  17942=>"00000000",
  17943=>"00000001",
  17944=>"11111111",
  17945=>"11111100",
  17946=>"00000011",
  17947=>"00000000",
  17948=>"11111100",
  17949=>"00000001",
  17950=>"00000000",
  17951=>"00000001",
  17952=>"11111111",
  17953=>"00000000",
  17954=>"00000001",
  17955=>"11111111",
  17956=>"00000100",
  17957=>"11111101",
  17958=>"00000001",
  17959=>"11111110",
  17960=>"00000010",
  17961=>"00000001",
  17962=>"00000100",
  17963=>"00000000",
  17964=>"11111101",
  17965=>"00000010",
  17966=>"11111100",
  17967=>"11111100",
  17968=>"11111110",
  17969=>"11111111",
  17970=>"00000001",
  17971=>"11111101",
  17972=>"00000011",
  17973=>"00000000",
  17974=>"00000010",
  17975=>"11111110",
  17976=>"11111110",
  17977=>"11111111",
  17978=>"00000010",
  17979=>"11111110",
  17980=>"00000011",
  17981=>"00000000",
  17982=>"11111110",
  17983=>"11111110",
  17984=>"11111101",
  17985=>"00000101",
  17986=>"00000000",
  17987=>"00000010",
  17988=>"00000010",
  17989=>"11111111",
  17990=>"11111101",
  17991=>"00000001",
  17992=>"11111101",
  17993=>"00000010",
  17994=>"11111111",
  17995=>"11111111",
  17996=>"00000000",
  17997=>"11111111",
  17998=>"11111110",
  17999=>"11111111",
  18000=>"11111110",
  18001=>"11111101",
  18002=>"00000000",
  18003=>"00000010",
  18004=>"11111110",
  18005=>"11111101",
  18006=>"11111110",
  18007=>"00000000",
  18008=>"11111111",
  18009=>"11111101",
  18010=>"00000001",
  18011=>"11111110",
  18012=>"11111111",
  18013=>"00000010",
  18014=>"00000001",
  18015=>"00000000",
  18016=>"00000000",
  18017=>"00000000",
  18018=>"11111110",
  18019=>"11111111",
  18020=>"11111110",
  18021=>"11111111",
  18022=>"11111110",
  18023=>"11111110",
  18024=>"11111011",
  18025=>"00000000",
  18026=>"00000000",
  18027=>"11111111",
  18028=>"11111110",
  18029=>"00000011",
  18030=>"00000010",
  18031=>"11111101",
  18032=>"00000001",
  18033=>"11111111",
  18034=>"11111110",
  18035=>"11111100",
  18036=>"00000000",
  18037=>"11111110",
  18038=>"11111111",
  18039=>"11111101",
  18040=>"11111111",
  18041=>"11111110",
  18042=>"11111110",
  18043=>"00000010",
  18044=>"00000011",
  18045=>"11111101",
  18046=>"11111110",
  18047=>"00000000",
  18048=>"00000001",
  18049=>"11111111",
  18050=>"00000101",
  18051=>"00000001",
  18052=>"00000001",
  18053=>"11111101",
  18054=>"00000101",
  18055=>"00000110",
  18056=>"00000001",
  18057=>"11111111",
  18058=>"11111101",
  18059=>"00000001",
  18060=>"11111101",
  18061=>"11111110",
  18062=>"11111110",
  18063=>"11111110",
  18064=>"00000011",
  18065=>"00000000",
  18066=>"11111101",
  18067=>"11111110",
  18068=>"00000010",
  18069=>"00000000",
  18070=>"11111111",
  18071=>"11111101",
  18072=>"00000010",
  18073=>"11111111",
  18074=>"11111111",
  18075=>"00000001",
  18076=>"00000000",
  18077=>"11111111",
  18078=>"11111111",
  18079=>"11111110",
  18080=>"00000010",
  18081=>"11111111",
  18082=>"00000011",
  18083=>"00000000",
  18084=>"00000000",
  18085=>"00000010",
  18086=>"00000000",
  18087=>"11111111",
  18088=>"00000000",
  18089=>"00000001",
  18090=>"11111101",
  18091=>"11111111",
  18092=>"11111101",
  18093=>"00000000",
  18094=>"11111111",
  18095=>"00000010",
  18096=>"00000001",
  18097=>"00000010",
  18098=>"00000010",
  18099=>"00000001",
  18100=>"11111110",
  18101=>"11111110",
  18102=>"00000010",
  18103=>"00000011",
  18104=>"00000000",
  18105=>"11111110",
  18106=>"00000001",
  18107=>"11111111",
  18108=>"11111111",
  18109=>"11111110",
  18110=>"11111111",
  18111=>"11111110",
  18112=>"00000000",
  18113=>"11111111",
  18114=>"00000010",
  18115=>"00000110",
  18116=>"11111110",
  18117=>"11111111",
  18118=>"00000000",
  18119=>"11111111",
  18120=>"11111111",
  18121=>"11111110",
  18122=>"00000001",
  18123=>"11111111",
  18124=>"00000011",
  18125=>"00000000",
  18126=>"00000010",
  18127=>"11111111",
  18128=>"11111101",
  18129=>"00000001",
  18130=>"11111111",
  18131=>"11111111",
  18132=>"00000010",
  18133=>"11111110",
  18134=>"11111101",
  18135=>"00000000",
  18136=>"11111111",
  18137=>"00000011",
  18138=>"00000010",
  18139=>"00000010",
  18140=>"11111110",
  18141=>"11111110",
  18142=>"00000110",
  18143=>"11111111",
  18144=>"00000001",
  18145=>"00000000",
  18146=>"00000001",
  18147=>"00000001",
  18148=>"11111110",
  18149=>"00000101",
  18150=>"11111110",
  18151=>"00000000",
  18152=>"11111110",
  18153=>"11111110",
  18154=>"00000010",
  18155=>"11111101",
  18156=>"00000000",
  18157=>"00000010",
  18158=>"00000000",
  18159=>"00000010",
  18160=>"00000000",
  18161=>"00000011",
  18162=>"00000001",
  18163=>"00000001",
  18164=>"11111110",
  18165=>"00000011",
  18166=>"11111110",
  18167=>"00000010",
  18168=>"00000010",
  18169=>"00000010",
  18170=>"11111111",
  18171=>"00000011",
  18172=>"00000011",
  18173=>"00000010",
  18174=>"00000011",
  18175=>"00000000",
  18176=>"11111101",
  18177=>"11111110",
  18178=>"11111111",
  18179=>"00000000",
  18180=>"11111110",
  18181=>"11111111",
  18182=>"11111101",
  18183=>"11111110",
  18184=>"00000000",
  18185=>"00000001",
  18186=>"11111111",
  18187=>"11111110",
  18188=>"00000001",
  18189=>"00000010",
  18190=>"00000010",
  18191=>"00000000",
  18192=>"00000010",
  18193=>"00000000",
  18194=>"11111101",
  18195=>"11111110",
  18196=>"00000000",
  18197=>"11111110",
  18198=>"00000100",
  18199=>"11111110",
  18200=>"11111101",
  18201=>"00000000",
  18202=>"11111110",
  18203=>"11111101",
  18204=>"00000001",
  18205=>"00000110",
  18206=>"00000001",
  18207=>"11111110",
  18208=>"11111101",
  18209=>"00000010",
  18210=>"00000001",
  18211=>"11111101",
  18212=>"11111111",
  18213=>"00000001",
  18214=>"11111111",
  18215=>"00000001",
  18216=>"00000000",
  18217=>"00000011",
  18218=>"11111111",
  18219=>"11111111",
  18220=>"00000010",
  18221=>"00000011",
  18222=>"00000010",
  18223=>"00000001",
  18224=>"00000001",
  18225=>"00000001",
  18226=>"00000100",
  18227=>"11111101",
  18228=>"11111110",
  18229=>"00000011",
  18230=>"11111111",
  18231=>"11111110",
  18232=>"00000000",
  18233=>"00000001",
  18234=>"11111111",
  18235=>"11111101",
  18236=>"00000010",
  18237=>"00000010",
  18238=>"11111111",
  18239=>"00000010",
  18240=>"00000011",
  18241=>"11111101",
  18242=>"11111101",
  18243=>"11111110",
  18244=>"00000001",
  18245=>"00000001",
  18246=>"11111101",
  18247=>"11111110",
  18248=>"11111111",
  18249=>"11111111",
  18250=>"00000000",
  18251=>"11111110",
  18252=>"11111111",
  18253=>"00000000",
  18254=>"00000001",
  18255=>"00000010",
  18256=>"00000000",
  18257=>"00000011",
  18258=>"00000001",
  18259=>"00000001",
  18260=>"00000000",
  18261=>"11111111",
  18262=>"11111101",
  18263=>"00000011",
  18264=>"11111110",
  18265=>"11111111",
  18266=>"11111101",
  18267=>"00000100",
  18268=>"11111111",
  18269=>"00000000",
  18270=>"00000001",
  18271=>"11111110",
  18272=>"00000000",
  18273=>"00000101",
  18274=>"11111111",
  18275=>"11111111",
  18276=>"00000000",
  18277=>"11111111",
  18278=>"00000001",
  18279=>"00000010",
  18280=>"00000111",
  18281=>"11111110",
  18282=>"11111101",
  18283=>"11111111",
  18284=>"11111101",
  18285=>"00000010",
  18286=>"11111110",
  18287=>"00000000",
  18288=>"00000000",
  18289=>"11111101",
  18290=>"11111111",
  18291=>"11111110",
  18292=>"11111111",
  18293=>"11111110",
  18294=>"00000000",
  18295=>"11111111",
  18296=>"00000001",
  18297=>"00000000",
  18298=>"11111111",
  18299=>"11111110",
  18300=>"11111110",
  18301=>"11111110",
  18302=>"11111111",
  18303=>"11111111",
  18304=>"00000010",
  18305=>"00000000",
  18306=>"11111101",
  18307=>"11111101",
  18308=>"11111100",
  18309=>"00000001",
  18310=>"11111111",
  18311=>"00000001",
  18312=>"11111101",
  18313=>"11111111",
  18314=>"11111101",
  18315=>"11111110",
  18316=>"00000000",
  18317=>"11111101",
  18318=>"00000101",
  18319=>"11111110",
  18320=>"11111110",
  18321=>"11111101",
  18322=>"00000001",
  18323=>"00000000",
  18324=>"00000000",
  18325=>"00000011",
  18326=>"11111101",
  18327=>"11111111",
  18328=>"11111101",
  18329=>"11111111",
  18330=>"11111110",
  18331=>"00000001",
  18332=>"11111111",
  18333=>"00000000",
  18334=>"00000100",
  18335=>"11111110",
  18336=>"11111100",
  18337=>"00000010",
  18338=>"00000000",
  18339=>"11111110",
  18340=>"00000010",
  18341=>"00000100",
  18342=>"11111110",
  18343=>"00000100",
  18344=>"11111111",
  18345=>"11111101",
  18346=>"11111110",
  18347=>"00000001",
  18348=>"11111110",
  18349=>"11111110",
  18350=>"00000011",
  18351=>"11111111",
  18352=>"11111110",
  18353=>"11111110",
  18354=>"00001000",
  18355=>"00000010",
  18356=>"11111110",
  18357=>"11111110",
  18358=>"11111101",
  18359=>"11111110",
  18360=>"11111110",
  18361=>"11111111",
  18362=>"00000000",
  18363=>"00000010",
  18364=>"00000010",
  18365=>"11111111",
  18366=>"11111101",
  18367=>"00000010",
  18368=>"00000001",
  18369=>"00000001",
  18370=>"11111101",
  18371=>"11111101",
  18372=>"00000000",
  18373=>"11111101",
  18374=>"00000100",
  18375=>"11111101",
  18376=>"11111110",
  18377=>"11111100",
  18378=>"00000011",
  18379=>"00000010",
  18380=>"11111101",
  18381=>"00000001",
  18382=>"00000001",
  18383=>"11111111",
  18384=>"00000010",
  18385=>"00000010",
  18386=>"11111011",
  18387=>"11111101",
  18388=>"00000011",
  18389=>"11111100",
  18390=>"11111110",
  18391=>"11111110",
  18392=>"00000000",
  18393=>"00000011",
  18394=>"11111101",
  18395=>"11111111",
  18396=>"11111101",
  18397=>"11111101",
  18398=>"11111110",
  18399=>"00000011",
  18400=>"00000001",
  18401=>"11111110",
  18402=>"00000000",
  18403=>"11111111",
  18404=>"11111111",
  18405=>"00000010",
  18406=>"11111111",
  18407=>"00000000",
  18408=>"00000000",
  18409=>"11111111",
  18410=>"11111101",
  18411=>"00000001",
  18412=>"00000001",
  18413=>"00000011",
  18414=>"11111101",
  18415=>"00000101",
  18416=>"00000010",
  18417=>"11111111",
  18418=>"00000011",
  18419=>"00000001",
  18420=>"11111110",
  18421=>"11111111",
  18422=>"00000010",
  18423=>"00000010",
  18424=>"11111101",
  18425=>"00000011",
  18426=>"11111101",
  18427=>"00000000",
  18428=>"11111101",
  18429=>"11111110",
  18430=>"11111101",
  18431=>"00000010",
  18432=>"11111111",
  18433=>"00000001",
  18434=>"11111110",
  18435=>"11111100",
  18436=>"11111110",
  18437=>"00000001",
  18438=>"00000000",
  18439=>"11111101",
  18440=>"11111100",
  18441=>"00000010",
  18442=>"11111101",
  18443=>"00000100",
  18444=>"00000000",
  18445=>"11111101",
  18446=>"00000010",
  18447=>"11111110",
  18448=>"11111111",
  18449=>"00000001",
  18450=>"00000110",
  18451=>"00000001",
  18452=>"11111110",
  18453=>"00000010",
  18454=>"11111110",
  18455=>"11111111",
  18456=>"00000001",
  18457=>"11111110",
  18458=>"00000000",
  18459=>"00000011",
  18460=>"00000001",
  18461=>"00000010",
  18462=>"00000010",
  18463=>"11111110",
  18464=>"00000010",
  18465=>"11111100",
  18466=>"11111110",
  18467=>"11111110",
  18468=>"00000010",
  18469=>"00000010",
  18470=>"11111111",
  18471=>"00000001",
  18472=>"00000000",
  18473=>"00000000",
  18474=>"00000001",
  18475=>"11111100",
  18476=>"00000000",
  18477=>"00000001",
  18478=>"11111111",
  18479=>"11111100",
  18480=>"00000010",
  18481=>"11111111",
  18482=>"00000001",
  18483=>"00000011",
  18484=>"11111110",
  18485=>"11111101",
  18486=>"00000000",
  18487=>"11111110",
  18488=>"11111111",
  18489=>"11111110",
  18490=>"00000100",
  18491=>"11111100",
  18492=>"11111110",
  18493=>"00000010",
  18494=>"11111111",
  18495=>"11111101",
  18496=>"00000001",
  18497=>"00000010",
  18498=>"11111111",
  18499=>"00000000",
  18500=>"00000010",
  18501=>"00000010",
  18502=>"11111111",
  18503=>"11111110",
  18504=>"11111111",
  18505=>"11111111",
  18506=>"11111101",
  18507=>"00000011",
  18508=>"00000011",
  18509=>"00000000",
  18510=>"00000010",
  18511=>"00000001",
  18512=>"00000010",
  18513=>"00000000",
  18514=>"00000000",
  18515=>"11111110",
  18516=>"00000001",
  18517=>"11111101",
  18518=>"11111110",
  18519=>"11111101",
  18520=>"11111110",
  18521=>"00000001",
  18522=>"11111110",
  18523=>"00000000",
  18524=>"00000101",
  18525=>"11111111",
  18526=>"11111111",
  18527=>"00000000",
  18528=>"00000000",
  18529=>"00000011",
  18530=>"11111110",
  18531=>"11111101",
  18532=>"00000001",
  18533=>"00000001",
  18534=>"11111110",
  18535=>"00000010",
  18536=>"00000001",
  18537=>"00000000",
  18538=>"00000001",
  18539=>"00000110",
  18540=>"11111101",
  18541=>"00000110",
  18542=>"00000001",
  18543=>"11111110",
  18544=>"11111111",
  18545=>"11111110",
  18546=>"11111110",
  18547=>"11111101",
  18548=>"11111111",
  18549=>"11111111",
  18550=>"11111101",
  18551=>"00000011",
  18552=>"00000001",
  18553=>"11111110",
  18554=>"11111101",
  18555=>"00000011",
  18556=>"11111100",
  18557=>"00000010",
  18558=>"11111111",
  18559=>"11111110",
  18560=>"00000000",
  18561=>"00000010",
  18562=>"00000010",
  18563=>"11111101",
  18564=>"00000001",
  18565=>"00000000",
  18566=>"11111110",
  18567=>"00000000",
  18568=>"11111110",
  18569=>"11111101",
  18570=>"00000001",
  18571=>"00000000",
  18572=>"00000010",
  18573=>"11111110",
  18574=>"00000000",
  18575=>"11111110",
  18576=>"11111111",
  18577=>"00000010",
  18578=>"00000000",
  18579=>"00000001",
  18580=>"11111110",
  18581=>"00000010",
  18582=>"11111110",
  18583=>"00000011",
  18584=>"11111110",
  18585=>"11111110",
  18586=>"00000001",
  18587=>"11111100",
  18588=>"11111101",
  18589=>"11111101",
  18590=>"00000001",
  18591=>"00000000",
  18592=>"11111101",
  18593=>"11111100",
  18594=>"00000000",
  18595=>"00000010",
  18596=>"00000010",
  18597=>"00000001",
  18598=>"11111111",
  18599=>"00000011",
  18600=>"00000001",
  18601=>"00000010",
  18602=>"11111111",
  18603=>"00000011",
  18604=>"00000101",
  18605=>"00000100",
  18606=>"11111100",
  18607=>"11111111",
  18608=>"00000001",
  18609=>"00000001",
  18610=>"11111101",
  18611=>"00000010",
  18612=>"00000001",
  18613=>"00000000",
  18614=>"00000001",
  18615=>"00000001",
  18616=>"00000010",
  18617=>"11111110",
  18618=>"00000011",
  18619=>"00000001",
  18620=>"00000000",
  18621=>"00000000",
  18622=>"00000000",
  18623=>"00000010",
  18624=>"11111111",
  18625=>"11111110",
  18626=>"00000001",
  18627=>"11111110",
  18628=>"11111101",
  18629=>"00000001",
  18630=>"11111110",
  18631=>"00000011",
  18632=>"00000011",
  18633=>"00000010",
  18634=>"00000010",
  18635=>"11111111",
  18636=>"11111111",
  18637=>"00000100",
  18638=>"11111100",
  18639=>"11111100",
  18640=>"00000011",
  18641=>"11111100",
  18642=>"00000010",
  18643=>"00000010",
  18644=>"00000001",
  18645=>"00000000",
  18646=>"00000000",
  18647=>"00000000",
  18648=>"11111101",
  18649=>"11111110",
  18650=>"11111111",
  18651=>"00000011",
  18652=>"00000010",
  18653=>"11111101",
  18654=>"00000001",
  18655=>"11111110",
  18656=>"11111111",
  18657=>"11111110",
  18658=>"00000000",
  18659=>"11111111",
  18660=>"11111100",
  18661=>"00000001",
  18662=>"11111101",
  18663=>"00000001",
  18664=>"11111111",
  18665=>"00000010",
  18666=>"00000000",
  18667=>"00000010",
  18668=>"11111111",
  18669=>"00000001",
  18670=>"00000010",
  18671=>"00000010",
  18672=>"00000000",
  18673=>"00000001",
  18674=>"00000001",
  18675=>"11111011",
  18676=>"11111110",
  18677=>"11111110",
  18678=>"00000000",
  18679=>"00000000",
  18680=>"00000100",
  18681=>"11111100",
  18682=>"00000000",
  18683=>"00000010",
  18684=>"11111110",
  18685=>"11111110",
  18686=>"11111101",
  18687=>"11111111",
  18688=>"11111111",
  18689=>"00000000",
  18690=>"00000001",
  18691=>"11111111",
  18692=>"00000000",
  18693=>"00000001",
  18694=>"11111101",
  18695=>"11111101",
  18696=>"00000011",
  18697=>"00000010",
  18698=>"00000101",
  18699=>"11111110",
  18700=>"11111110",
  18701=>"00000001",
  18702=>"00000101",
  18703=>"00000010",
  18704=>"11111111",
  18705=>"00000001",
  18706=>"11111101",
  18707=>"00000011",
  18708=>"11111101",
  18709=>"00000000",
  18710=>"11111110",
  18711=>"00000001",
  18712=>"00000000",
  18713=>"00000001",
  18714=>"00000010",
  18715=>"00000010",
  18716=>"00000101",
  18717=>"00000001",
  18718=>"11111101",
  18719=>"11111101",
  18720=>"00000001",
  18721=>"00000001",
  18722=>"00000000",
  18723=>"11111110",
  18724=>"00000010",
  18725=>"00000101",
  18726=>"11111110",
  18727=>"11111110",
  18728=>"00000001",
  18729=>"11111101",
  18730=>"11111111",
  18731=>"00000100",
  18732=>"00000010",
  18733=>"11111111",
  18734=>"00000000",
  18735=>"11111111",
  18736=>"11111101",
  18737=>"00000001",
  18738=>"11111110",
  18739=>"11111110",
  18740=>"11111111",
  18741=>"00000001",
  18742=>"11111101",
  18743=>"11111111",
  18744=>"00000010",
  18745=>"00000011",
  18746=>"00000011",
  18747=>"11111110",
  18748=>"00000001",
  18749=>"11111101",
  18750=>"11111111",
  18751=>"00000000",
  18752=>"00000100",
  18753=>"11111100",
  18754=>"00000001",
  18755=>"00000000",
  18756=>"00000010",
  18757=>"00000001",
  18758=>"11111100",
  18759=>"00000000",
  18760=>"11111110",
  18761=>"00000001",
  18762=>"11111101",
  18763=>"11111101",
  18764=>"00000101",
  18765=>"00000010",
  18766=>"00000000",
  18767=>"11111101",
  18768=>"00000001",
  18769=>"00000001",
  18770=>"00000000",
  18771=>"11111101",
  18772=>"11111110",
  18773=>"11111110",
  18774=>"11111110",
  18775=>"00000001",
  18776=>"11111110",
  18777=>"11111101",
  18778=>"11111110",
  18779=>"11111101",
  18780=>"11111110",
  18781=>"11111111",
  18782=>"00000001",
  18783=>"11111101",
  18784=>"11111111",
  18785=>"11111101",
  18786=>"00000001",
  18787=>"11111111",
  18788=>"11111110",
  18789=>"00000000",
  18790=>"00000001",
  18791=>"11111111",
  18792=>"11111110",
  18793=>"00000010",
  18794=>"11111110",
  18795=>"11111100",
  18796=>"00000011",
  18797=>"00000011",
  18798=>"11111101",
  18799=>"11111111",
  18800=>"00000000",
  18801=>"11111110",
  18802=>"11111111",
  18803=>"00000001",
  18804=>"00000000",
  18805=>"00000000",
  18806=>"00000001",
  18807=>"11111101",
  18808=>"00000011",
  18809=>"00000100",
  18810=>"11111101",
  18811=>"00000011",
  18812=>"11111111",
  18813=>"00000001",
  18814=>"00000001",
  18815=>"00000100",
  18816=>"11111100",
  18817=>"00000001",
  18818=>"11111110",
  18819=>"11111101",
  18820=>"11111111",
  18821=>"00000101",
  18822=>"11111111",
  18823=>"00000000",
  18824=>"00000011",
  18825=>"00000001",
  18826=>"00000000",
  18827=>"11111111",
  18828=>"00000000",
  18829=>"00000001",
  18830=>"11111100",
  18831=>"11111110",
  18832=>"11111110",
  18833=>"00000000",
  18834=>"11111100",
  18835=>"00000010",
  18836=>"11111101",
  18837=>"00000001",
  18838=>"00000011",
  18839=>"00000110",
  18840=>"11111111",
  18841=>"11111101",
  18842=>"00000001",
  18843=>"00000001",
  18844=>"00000000",
  18845=>"00000001",
  18846=>"11111111",
  18847=>"00000001",
  18848=>"00000000",
  18849=>"00000001",
  18850=>"11111101",
  18851=>"00000010",
  18852=>"00000000",
  18853=>"00000011",
  18854=>"00000000",
  18855=>"11111110",
  18856=>"00000001",
  18857=>"11111101",
  18858=>"00000010",
  18859=>"11111101",
  18860=>"00000010",
  18861=>"00000011",
  18862=>"11111111",
  18863=>"11111101",
  18864=>"11111111",
  18865=>"11111101",
  18866=>"00000001",
  18867=>"00000000",
  18868=>"11111100",
  18869=>"00000010",
  18870=>"11111110",
  18871=>"11111110",
  18872=>"00000010",
  18873=>"11111101",
  18874=>"11111111",
  18875=>"00000010",
  18876=>"00000011",
  18877=>"00000001",
  18878=>"11111110",
  18879=>"11111111",
  18880=>"11111110",
  18881=>"11111111",
  18882=>"11111101",
  18883=>"00000100",
  18884=>"11111110",
  18885=>"00000010",
  18886=>"11111110",
  18887=>"00000000",
  18888=>"00000010",
  18889=>"11111101",
  18890=>"00000010",
  18891=>"00000011",
  18892=>"11111101",
  18893=>"11111111",
  18894=>"00000010",
  18895=>"11111110",
  18896=>"00000001",
  18897=>"00000010",
  18898=>"00000011",
  18899=>"00000001",
  18900=>"00000001",
  18901=>"11111110",
  18902=>"11111100",
  18903=>"00000010",
  18904=>"11111111",
  18905=>"00000000",
  18906=>"00000000",
  18907=>"11111111",
  18908=>"11111101",
  18909=>"11111101",
  18910=>"00000010",
  18911=>"00000000",
  18912=>"00000001",
  18913=>"11111100",
  18914=>"00000000",
  18915=>"11111101",
  18916=>"00000001",
  18917=>"00000001",
  18918=>"00000000",
  18919=>"00000001",
  18920=>"00000011",
  18921=>"00000001",
  18922=>"00000000",
  18923=>"00000001",
  18924=>"11111101",
  18925=>"11111111",
  18926=>"11111111",
  18927=>"00000001",
  18928=>"11111110",
  18929=>"11111110",
  18930=>"11111111",
  18931=>"11111101",
  18932=>"11111111",
  18933=>"11111111",
  18934=>"00000001",
  18935=>"00000010",
  18936=>"00000010",
  18937=>"11111111",
  18938=>"11111110",
  18939=>"00000111",
  18940=>"11111110",
  18941=>"11111100",
  18942=>"11111111",
  18943=>"11111101",
  18944=>"11111101",
  18945=>"00000100",
  18946=>"11111111",
  18947=>"00000010",
  18948=>"00000001",
  18949=>"00000100",
  18950=>"00000000",
  18951=>"11111111",
  18952=>"00000001",
  18953=>"11111011",
  18954=>"11111111",
  18955=>"00000001",
  18956=>"00000010",
  18957=>"00000001",
  18958=>"11111111",
  18959=>"00000001",
  18960=>"00000011",
  18961=>"00000100",
  18962=>"00000010",
  18963=>"00000000",
  18964=>"11111101",
  18965=>"00000000",
  18966=>"11111110",
  18967=>"11111100",
  18968=>"00000011",
  18969=>"00000001",
  18970=>"11111100",
  18971=>"11111101",
  18972=>"00000001",
  18973=>"00000011",
  18974=>"11111110",
  18975=>"00000010",
  18976=>"00000001",
  18977=>"11111110",
  18978=>"00000010",
  18979=>"11111111",
  18980=>"11111110",
  18981=>"11111111",
  18982=>"00000010",
  18983=>"00000000",
  18984=>"11111111",
  18985=>"11111111",
  18986=>"00000100",
  18987=>"11111110",
  18988=>"11111100",
  18989=>"11111101",
  18990=>"00000011",
  18991=>"00000011",
  18992=>"11111101",
  18993=>"11111111",
  18994=>"11111111",
  18995=>"00000000",
  18996=>"11111101",
  18997=>"00000001",
  18998=>"11111111",
  18999=>"00000100",
  19000=>"11111111",
  19001=>"00000010",
  19002=>"11111101",
  19003=>"11111101",
  19004=>"11111110",
  19005=>"11111110",
  19006=>"00000110",
  19007=>"00000010",
  19008=>"00000010",
  19009=>"00000001",
  19010=>"11111101",
  19011=>"11111101",
  19012=>"11111110",
  19013=>"11111101",
  19014=>"11111101",
  19015=>"00000001",
  19016=>"11111111",
  19017=>"00000010",
  19018=>"00000001",
  19019=>"00000010",
  19020=>"11111101",
  19021=>"00000000",
  19022=>"00000000",
  19023=>"11111110",
  19024=>"11111100",
  19025=>"00000000",
  19026=>"00000000",
  19027=>"11111110",
  19028=>"00000011",
  19029=>"00000101",
  19030=>"11111110",
  19031=>"00000011",
  19032=>"00000000",
  19033=>"11111111",
  19034=>"11111101",
  19035=>"00000010",
  19036=>"00000000",
  19037=>"00000011",
  19038=>"00000001",
  19039=>"11111110",
  19040=>"00000010",
  19041=>"00000001",
  19042=>"11111110",
  19043=>"00000010",
  19044=>"00000010",
  19045=>"11111111",
  19046=>"00000000",
  19047=>"11111110",
  19048=>"11111110",
  19049=>"11111111",
  19050=>"00000001",
  19051=>"11111110",
  19052=>"00000101",
  19053=>"11111100",
  19054=>"00000000",
  19055=>"11111101",
  19056=>"00000010",
  19057=>"11111111",
  19058=>"11111111",
  19059=>"11111101",
  19060=>"11111110",
  19061=>"00000001",
  19062=>"11111110",
  19063=>"00000001",
  19064=>"00000001",
  19065=>"11111101",
  19066=>"11111111",
  19067=>"11111111",
  19068=>"11111110",
  19069=>"11111110",
  19070=>"00000000",
  19071=>"00000100",
  19072=>"11111101",
  19073=>"00000010",
  19074=>"00000010",
  19075=>"11111101",
  19076=>"11111110",
  19077=>"11111111",
  19078=>"11111110",
  19079=>"11111111",
  19080=>"00000010",
  19081=>"11111110",
  19082=>"00000100",
  19083=>"00000010",
  19084=>"11111101",
  19085=>"11111111",
  19086=>"00000010",
  19087=>"00000010",
  19088=>"00000010",
  19089=>"00000000",
  19090=>"11111110",
  19091=>"00000010",
  19092=>"00000010",
  19093=>"11111110",
  19094=>"00000001",
  19095=>"00000001",
  19096=>"11111111",
  19097=>"11111100",
  19098=>"00000010",
  19099=>"00000000",
  19100=>"11111101",
  19101=>"11111111",
  19102=>"00000000",
  19103=>"00000001",
  19104=>"11111111",
  19105=>"11111110",
  19106=>"00000001",
  19107=>"11111111",
  19108=>"00000000",
  19109=>"11111101",
  19110=>"00000011",
  19111=>"00000001",
  19112=>"11111110",
  19113=>"00000011",
  19114=>"00000000",
  19115=>"00000000",
  19116=>"11111111",
  19117=>"11111110",
  19118=>"11111111",
  19119=>"11111100",
  19120=>"00000000",
  19121=>"11111111",
  19122=>"00000010",
  19123=>"00000000",
  19124=>"00000010",
  19125=>"00000000",
  19126=>"11111110",
  19127=>"11111101",
  19128=>"00000001",
  19129=>"11111111",
  19130=>"00000001",
  19131=>"11111101",
  19132=>"00000010",
  19133=>"11111111",
  19134=>"00000000",
  19135=>"00000010",
  19136=>"00000010",
  19137=>"11111101",
  19138=>"11111111",
  19139=>"00000010",
  19140=>"11111110",
  19141=>"11111110",
  19142=>"11111101",
  19143=>"11111110",
  19144=>"00000001",
  19145=>"11111111",
  19146=>"00000000",
  19147=>"11111101",
  19148=>"00000101",
  19149=>"11111101",
  19150=>"11111110",
  19151=>"00000001",
  19152=>"00000000",
  19153=>"11111110",
  19154=>"11111110",
  19155=>"11111101",
  19156=>"00000010",
  19157=>"00000000",
  19158=>"11111111",
  19159=>"00000010",
  19160=>"00000001",
  19161=>"11111111",
  19162=>"00000000",
  19163=>"11111111",
  19164=>"00000001",
  19165=>"11111101",
  19166=>"11111111",
  19167=>"00000000",
  19168=>"11111011",
  19169=>"00000010",
  19170=>"00000001",
  19171=>"11111110",
  19172=>"00000010",
  19173=>"00000110",
  19174=>"00000000",
  19175=>"00000001",
  19176=>"00000001",
  19177=>"11111111",
  19178=>"11111101",
  19179=>"11111111",
  19180=>"00000000",
  19181=>"11111101",
  19182=>"11111101",
  19183=>"11111101",
  19184=>"11111111",
  19185=>"11111111",
  19186=>"11111111",
  19187=>"00000000",
  19188=>"00000000",
  19189=>"00000010",
  19190=>"00000011",
  19191=>"11111111",
  19192=>"11111101",
  19193=>"11111111",
  19194=>"00000010",
  19195=>"00000100",
  19196=>"00000000",
  19197=>"00000000",
  19198=>"11111110",
  19199=>"00000001",
  19200=>"00000010",
  19201=>"11111110",
  19202=>"00000110",
  19203=>"00000011",
  19204=>"11111101",
  19205=>"00000010",
  19206=>"00000000",
  19207=>"00000000",
  19208=>"11111100",
  19209=>"00000001",
  19210=>"11111101",
  19211=>"00000000",
  19212=>"00000001",
  19213=>"11111110",
  19214=>"00000010",
  19215=>"11111111",
  19216=>"11111111",
  19217=>"11111101",
  19218=>"00000000",
  19219=>"11111101",
  19220=>"00000010",
  19221=>"00000000",
  19222=>"00000000",
  19223=>"11111101",
  19224=>"11111101",
  19225=>"11111110",
  19226=>"11111100",
  19227=>"11111111",
  19228=>"00000001",
  19229=>"11111100",
  19230=>"11111101",
  19231=>"00000101",
  19232=>"11111111",
  19233=>"11111111",
  19234=>"00000000",
  19235=>"00000010",
  19236=>"00000011",
  19237=>"00000000",
  19238=>"11111101",
  19239=>"11111100",
  19240=>"00000010",
  19241=>"11111101",
  19242=>"00000001",
  19243=>"00000101",
  19244=>"11111111",
  19245=>"11111111",
  19246=>"11111111",
  19247=>"00000001",
  19248=>"00000000",
  19249=>"11111101",
  19250=>"00000001",
  19251=>"11111111",
  19252=>"11111101",
  19253=>"11111101",
  19254=>"11111111",
  19255=>"11111101",
  19256=>"00000001",
  19257=>"00000000",
  19258=>"00000000",
  19259=>"11111111",
  19260=>"00000010",
  19261=>"11111101",
  19262=>"11111110",
  19263=>"11111111",
  19264=>"11111110",
  19265=>"00000001",
  19266=>"00000011",
  19267=>"11111110",
  19268=>"11111100",
  19269=>"11111110",
  19270=>"00000000",
  19271=>"00000001",
  19272=>"00000000",
  19273=>"11111110",
  19274=>"00000010",
  19275=>"00000011",
  19276=>"00000011",
  19277=>"11111111",
  19278=>"00000001",
  19279=>"11111111",
  19280=>"00000001",
  19281=>"00000000",
  19282=>"00000011",
  19283=>"00000001",
  19284=>"00000010",
  19285=>"00000001",
  19286=>"00000001",
  19287=>"11111111",
  19288=>"11111101",
  19289=>"00000001",
  19290=>"11111110",
  19291=>"00000100",
  19292=>"00000000",
  19293=>"11111110",
  19294=>"11111101",
  19295=>"11111101",
  19296=>"11111101",
  19297=>"11111110",
  19298=>"11111111",
  19299=>"11111111",
  19300=>"11111111",
  19301=>"00000010",
  19302=>"11111110",
  19303=>"00000101",
  19304=>"11111110",
  19305=>"11111101",
  19306=>"00000000",
  19307=>"00000010",
  19308=>"00000000",
  19309=>"00000000",
  19310=>"11111110",
  19311=>"11111100",
  19312=>"00000001",
  19313=>"11111111",
  19314=>"00000001",
  19315=>"00000001",
  19316=>"00000001",
  19317=>"00000000",
  19318=>"11111110",
  19319=>"00000000",
  19320=>"11111110",
  19321=>"00000000",
  19322=>"00000001",
  19323=>"00000100",
  19324=>"00000001",
  19325=>"00000101",
  19326=>"00000010",
  19327=>"00000010",
  19328=>"11111110",
  19329=>"11111110",
  19330=>"11111110",
  19331=>"00000001",
  19332=>"11111100",
  19333=>"11111110",
  19334=>"11111111",
  19335=>"11111101",
  19336=>"11111101",
  19337=>"11111100",
  19338=>"11111110",
  19339=>"00000000",
  19340=>"11111110",
  19341=>"11111111",
  19342=>"00000000",
  19343=>"11111101",
  19344=>"00000010",
  19345=>"11111110",
  19346=>"11111110",
  19347=>"00000001",
  19348=>"11111100",
  19349=>"00000000",
  19350=>"11111110",
  19351=>"11111110",
  19352=>"11111111",
  19353=>"00000100",
  19354=>"11111110",
  19355=>"00000011",
  19356=>"00000010",
  19357=>"11111110",
  19358=>"00000010",
  19359=>"11111101",
  19360=>"00000001",
  19361=>"00000010",
  19362=>"00000000",
  19363=>"00000001",
  19364=>"11111110",
  19365=>"11111101",
  19366=>"00000011",
  19367=>"11111101",
  19368=>"11111101",
  19369=>"11111110",
  19370=>"00000001",
  19371=>"11111111",
  19372=>"00000001",
  19373=>"11111111",
  19374=>"11111111",
  19375=>"00000001",
  19376=>"00000001",
  19377=>"00000011",
  19378=>"00000010",
  19379=>"00000001",
  19380=>"00000001",
  19381=>"11111110",
  19382=>"11111101",
  19383=>"00000010",
  19384=>"11111101",
  19385=>"11111111",
  19386=>"00000010",
  19387=>"00000001",
  19388=>"11111111",
  19389=>"00000011",
  19390=>"00000011",
  19391=>"11111101",
  19392=>"11111111",
  19393=>"11111111",
  19394=>"00000011",
  19395=>"00000001",
  19396=>"00000000",
  19397=>"00000010",
  19398=>"00000110",
  19399=>"00000000",
  19400=>"00000010",
  19401=>"11111111",
  19402=>"00000011",
  19403=>"11111111",
  19404=>"00000101",
  19405=>"11111111",
  19406=>"00000010",
  19407=>"00000001",
  19408=>"11111111",
  19409=>"00000100",
  19410=>"11111111",
  19411=>"11111101",
  19412=>"11111100",
  19413=>"00000010",
  19414=>"00000011",
  19415=>"11111110",
  19416=>"11111110",
  19417=>"00000101",
  19418=>"00000001",
  19419=>"00000000",
  19420=>"00000010",
  19421=>"00000000",
  19422=>"00000001",
  19423=>"11111101",
  19424=>"11111110",
  19425=>"11111111",
  19426=>"00000010",
  19427=>"00000001",
  19428=>"11111111",
  19429=>"00000010",
  19430=>"11111110",
  19431=>"11111110",
  19432=>"11111111",
  19433=>"11111110",
  19434=>"00000110",
  19435=>"11111110",
  19436=>"00000000",
  19437=>"00000000",
  19438=>"11111101",
  19439=>"00000010",
  19440=>"00000010",
  19441=>"00000000",
  19442=>"00000100",
  19443=>"00000000",
  19444=>"11111110",
  19445=>"00000001",
  19446=>"00000010",
  19447=>"00000001",
  19448=>"00000000",
  19449=>"00000001",
  19450=>"00000100",
  19451=>"11111111",
  19452=>"11111110",
  19453=>"00000000",
  19454=>"11111111",
  19455=>"00000001",
  19456=>"00000001",
  19457=>"11111110",
  19458=>"11111110",
  19459=>"00000011",
  19460=>"11111111",
  19461=>"00000011",
  19462=>"00000001",
  19463=>"00000000",
  19464=>"00000100",
  19465=>"00000011",
  19466=>"00000100",
  19467=>"00000000",
  19468=>"11111111",
  19469=>"00000101",
  19470=>"00000001",
  19471=>"00000011",
  19472=>"00000000",
  19473=>"11111111",
  19474=>"00000100",
  19475=>"00000100",
  19476=>"11111110",
  19477=>"11111110",
  19478=>"11111101",
  19479=>"00000101",
  19480=>"00000100",
  19481=>"00000001",
  19482=>"00000010",
  19483=>"11111111",
  19484=>"11111101",
  19485=>"00000010",
  19486=>"11111111",
  19487=>"11111111",
  19488=>"11111101",
  19489=>"00000101",
  19490=>"00000011",
  19491=>"00000000",
  19492=>"11111111",
  19493=>"00000011",
  19494=>"00000000",
  19495=>"11111110",
  19496=>"11111111",
  19497=>"00000001",
  19498=>"00000100",
  19499=>"00000001",
  19500=>"00000001",
  19501=>"11111110",
  19502=>"00000000",
  19503=>"00000001",
  19504=>"11111111",
  19505=>"11111110",
  19506=>"00000010",
  19507=>"00000100",
  19508=>"00000010",
  19509=>"11111110",
  19510=>"00000011",
  19511=>"11111100",
  19512=>"00000001",
  19513=>"11111110",
  19514=>"11111111",
  19515=>"11111111",
  19516=>"00000001",
  19517=>"11111111",
  19518=>"00000111",
  19519=>"00000011",
  19520=>"00000000",
  19521=>"00000011",
  19522=>"11111110",
  19523=>"00000001",
  19524=>"00000000",
  19525=>"00000100",
  19526=>"00000010",
  19527=>"00000001",
  19528=>"11111101",
  19529=>"00000011",
  19530=>"00000000",
  19531=>"11111110",
  19532=>"11111101",
  19533=>"11111011",
  19534=>"11111111",
  19535=>"00000000",
  19536=>"00000001",
  19537=>"00000000",
  19538=>"00000010",
  19539=>"00000010",
  19540=>"11111111",
  19541=>"11111110",
  19542=>"00000010",
  19543=>"00000011",
  19544=>"11111110",
  19545=>"11111110",
  19546=>"00000001",
  19547=>"11111100",
  19548=>"11111110",
  19549=>"00000010",
  19550=>"11111100",
  19551=>"11111111",
  19552=>"11111111",
  19553=>"00000000",
  19554=>"00000110",
  19555=>"11111110",
  19556=>"00000001",
  19557=>"00000010",
  19558=>"00000001",
  19559=>"00000100",
  19560=>"11111110",
  19561=>"00000010",
  19562=>"11111011",
  19563=>"00000101",
  19564=>"00000010",
  19565=>"00000001",
  19566=>"00000000",
  19567=>"00000100",
  19568=>"00000011",
  19569=>"00000011",
  19570=>"00000001",
  19571=>"11111100",
  19572=>"11111110",
  19573=>"00000000",
  19574=>"00000101",
  19575=>"00000010",
  19576=>"11111111",
  19577=>"00000000",
  19578=>"00000100",
  19579=>"00000010",
  19580=>"00000000",
  19581=>"00000100",
  19582=>"00000100",
  19583=>"00000100",
  19584=>"00000010",
  19585=>"00000001",
  19586=>"00000100",
  19587=>"00000011",
  19588=>"00000010",
  19589=>"11111101",
  19590=>"00000010",
  19591=>"11111110",
  19592=>"00000101",
  19593=>"00000001",
  19594=>"00000010",
  19595=>"00000001",
  19596=>"11111110",
  19597=>"11111100",
  19598=>"00000000",
  19599=>"00000100",
  19600=>"00000010",
  19601=>"00000101",
  19602=>"00000100",
  19603=>"00000010",
  19604=>"11111101",
  19605=>"00000100",
  19606=>"00000000",
  19607=>"00000100",
  19608=>"11111111",
  19609=>"00000010",
  19610=>"11111111",
  19611=>"00000100",
  19612=>"00000000",
  19613=>"00000100",
  19614=>"00000001",
  19615=>"00000000",
  19616=>"11111110",
  19617=>"11111100",
  19618=>"11111101",
  19619=>"00000111",
  19620=>"11111100",
  19621=>"00000010",
  19622=>"11111110",
  19623=>"11111101",
  19624=>"11111110",
  19625=>"00000110",
  19626=>"00000001",
  19627=>"00000100",
  19628=>"00000100",
  19629=>"00000101",
  19630=>"00000010",
  19631=>"00000100",
  19632=>"00000011",
  19633=>"00000100",
  19634=>"00000000",
  19635=>"11111101",
  19636=>"00000001",
  19637=>"00000100",
  19638=>"11111110",
  19639=>"00000100",
  19640=>"11111111",
  19641=>"00000011",
  19642=>"00000010",
  19643=>"00000101",
  19644=>"11111101",
  19645=>"11111101",
  19646=>"11111110",
  19647=>"11111110",
  19648=>"00000000",
  19649=>"00000000",
  19650=>"00000000",
  19651=>"00000101",
  19652=>"00000000",
  19653=>"00000100",
  19654=>"00000010",
  19655=>"00000000",
  19656=>"00000010",
  19657=>"00000000",
  19658=>"00000010",
  19659=>"00000011",
  19660=>"11111110",
  19661=>"00000000",
  19662=>"11111111",
  19663=>"00000000",
  19664=>"00000110",
  19665=>"00000100",
  19666=>"00000000",
  19667=>"00000000",
  19668=>"11111111",
  19669=>"00000010",
  19670=>"11111101",
  19671=>"00000101",
  19672=>"11111111",
  19673=>"00000010",
  19674=>"00000010",
  19675=>"00000010",
  19676=>"11111110",
  19677=>"11111110",
  19678=>"11111110",
  19679=>"00000001",
  19680=>"00000011",
  19681=>"00000001",
  19682=>"11111111",
  19683=>"11111101",
  19684=>"00000001",
  19685=>"11111100",
  19686=>"00000110",
  19687=>"11111110",
  19688=>"00000000",
  19689=>"00000010",
  19690=>"00000010",
  19691=>"00000010",
  19692=>"00000011",
  19693=>"11111111",
  19694=>"11111101",
  19695=>"00000100",
  19696=>"00000100",
  19697=>"00000010",
  19698=>"11111110",
  19699=>"11111111",
  19700=>"00000010",
  19701=>"00000001",
  19702=>"11111101",
  19703=>"00000011",
  19704=>"00000001",
  19705=>"00000011",
  19706=>"00000000",
  19707=>"00000000",
  19708=>"11111011",
  19709=>"00000000",
  19710=>"11111101",
  19711=>"00000001",
  19712=>"00000001",
  19713=>"11111111",
  19714=>"00000011",
  19715=>"11111100",
  19716=>"00000001",
  19717=>"00000100",
  19718=>"11111111",
  19719=>"00000001",
  19720=>"00000001",
  19721=>"11111110",
  19722=>"00000111",
  19723=>"11111111",
  19724=>"11111110",
  19725=>"11111110",
  19726=>"11111101",
  19727=>"00000001",
  19728=>"11111100",
  19729=>"00000000",
  19730=>"00000010",
  19731=>"00000010",
  19732=>"11111100",
  19733=>"00000011",
  19734=>"00000010",
  19735=>"00000010",
  19736=>"00000010",
  19737=>"11111111",
  19738=>"11111101",
  19739=>"00000010",
  19740=>"00000100",
  19741=>"11111101",
  19742=>"00000001",
  19743=>"00000010",
  19744=>"00000000",
  19745=>"00000000",
  19746=>"11111111",
  19747=>"00000001",
  19748=>"00000100",
  19749=>"00000010",
  19750=>"00000101",
  19751=>"00000110",
  19752=>"00000100",
  19753=>"00000011",
  19754=>"11111111",
  19755=>"11111111",
  19756=>"11111101",
  19757=>"00000010",
  19758=>"00000010",
  19759=>"11111101",
  19760=>"11111101",
  19761=>"11111111",
  19762=>"00000011",
  19763=>"11111110",
  19764=>"11111101",
  19765=>"00000001",
  19766=>"00000000",
  19767=>"00000011",
  19768=>"00000010",
  19769=>"00000010",
  19770=>"00000100",
  19771=>"00000000",
  19772=>"00000010",
  19773=>"11111100",
  19774=>"00000010",
  19775=>"11111101",
  19776=>"00000110",
  19777=>"11111110",
  19778=>"11111110",
  19779=>"11111111",
  19780=>"00000011",
  19781=>"00000111",
  19782=>"00000000",
  19783=>"11111111",
  19784=>"00000010",
  19785=>"00000011",
  19786=>"00000001",
  19787=>"00000010",
  19788=>"00000010",
  19789=>"11111001",
  19790=>"00000110",
  19791=>"00000000",
  19792=>"11111111",
  19793=>"00000001",
  19794=>"00000010",
  19795=>"11111111",
  19796=>"11111101",
  19797=>"11111111",
  19798=>"11111100",
  19799=>"00000000",
  19800=>"00000011",
  19801=>"00000100",
  19802=>"00000010",
  19803=>"00000100",
  19804=>"11111101",
  19805=>"00000001",
  19806=>"11111101",
  19807=>"11111101",
  19808=>"00000000",
  19809=>"11111111",
  19810=>"00000000",
  19811=>"11111110",
  19812=>"11111101",
  19813=>"11111101",
  19814=>"00000001",
  19815=>"00000100",
  19816=>"00000101",
  19817=>"00000000",
  19818=>"00000010",
  19819=>"00000000",
  19820=>"00000011",
  19821=>"00000100",
  19822=>"00000011",
  19823=>"11111100",
  19824=>"00000000",
  19825=>"11111101",
  19826=>"11111111",
  19827=>"00000001",
  19828=>"00000001",
  19829=>"00000000",
  19830=>"11111101",
  19831=>"00000001",
  19832=>"11111100",
  19833=>"00000100",
  19834=>"11111110",
  19835=>"00000000",
  19836=>"11111110",
  19837=>"11111111",
  19838=>"00000010",
  19839=>"00000001",
  19840=>"00000001",
  19841=>"11111101",
  19842=>"11111101",
  19843=>"11111111",
  19844=>"11111111",
  19845=>"00000011",
  19846=>"00000010",
  19847=>"00000000",
  19848=>"11111110",
  19849=>"11111111",
  19850=>"11111111",
  19851=>"00000110",
  19852=>"11111101",
  19853=>"11111110",
  19854=>"00000110",
  19855=>"00000001",
  19856=>"00000101",
  19857=>"00000011",
  19858=>"11111011",
  19859=>"11111111",
  19860=>"00000101",
  19861=>"11111101",
  19862=>"00000001",
  19863=>"11111111",
  19864=>"11111110",
  19865=>"11111101",
  19866=>"00000010",
  19867=>"11111111",
  19868=>"11111110",
  19869=>"11111110",
  19870=>"11111111",
  19871=>"00000011",
  19872=>"11111110",
  19873=>"11111100",
  19874=>"00000010",
  19875=>"00000001",
  19876=>"00000011",
  19877=>"00000001",
  19878=>"00000001",
  19879=>"11111111",
  19880=>"11111110",
  19881=>"11111110",
  19882=>"11111110",
  19883=>"11111100",
  19884=>"00000001",
  19885=>"11111111",
  19886=>"00000011",
  19887=>"00000001",
  19888=>"00000011",
  19889=>"00000010",
  19890=>"00000100",
  19891=>"11111111",
  19892=>"11111100",
  19893=>"00000100",
  19894=>"00000001",
  19895=>"11111101",
  19896=>"00000110",
  19897=>"00000001",
  19898=>"00000000",
  19899=>"00000001",
  19900=>"00000001",
  19901=>"11111111",
  19902=>"00000101",
  19903=>"11111110",
  19904=>"00000010",
  19905=>"11111101",
  19906=>"00000010",
  19907=>"11111110",
  19908=>"00000100",
  19909=>"00000000",
  19910=>"11111111",
  19911=>"00000101",
  19912=>"11111111",
  19913=>"11111111",
  19914=>"00000101",
  19915=>"11111111",
  19916=>"00000011",
  19917=>"00000000",
  19918=>"00000011",
  19919=>"00000001",
  19920=>"11111110",
  19921=>"00000011",
  19922=>"00000000",
  19923=>"00000000",
  19924=>"00000000",
  19925=>"00000000",
  19926=>"00000001",
  19927=>"00000001",
  19928=>"11111110",
  19929=>"00000010",
  19930=>"00000100",
  19931=>"00000110",
  19932=>"11111011",
  19933=>"00000000",
  19934=>"00000100",
  19935=>"00000001",
  19936=>"00000000",
  19937=>"00000010",
  19938=>"00000000",
  19939=>"11111110",
  19940=>"00000100",
  19941=>"11111111",
  19942=>"11111101",
  19943=>"00000001",
  19944=>"00000100",
  19945=>"00000010",
  19946=>"00000011",
  19947=>"00000101",
  19948=>"11111111",
  19949=>"00000001",
  19950=>"11111101",
  19951=>"00000010",
  19952=>"11111111",
  19953=>"00000100",
  19954=>"00000000",
  19955=>"00000010",
  19956=>"00000000",
  19957=>"00000100",
  19958=>"00000000",
  19959=>"00000001",
  19960=>"11111110",
  19961=>"11111101",
  19962=>"00000001",
  19963=>"00000001",
  19964=>"00000001",
  19965=>"00000001",
  19966=>"00000100",
  19967=>"11111010",
  19968=>"11111110",
  19969=>"00000001",
  19970=>"11111101",
  19971=>"00000001",
  19972=>"11111101",
  19973=>"00000000",
  19974=>"00000100",
  19975=>"00000010",
  19976=>"11111110",
  19977=>"11111111",
  19978=>"00000001",
  19979=>"00000001",
  19980=>"11111101",
  19981=>"00000001",
  19982=>"11111111",
  19983=>"00000000",
  19984=>"00000010",
  19985=>"00000010",
  19986=>"11111111",
  19987=>"00000000",
  19988=>"00000011",
  19989=>"00000010",
  19990=>"11111110",
  19991=>"00000001",
  19992=>"00000000",
  19993=>"00000000",
  19994=>"00000010",
  19995=>"11111110",
  19996=>"11111111",
  19997=>"00000000",
  19998=>"11111101",
  19999=>"00000000",
  20000=>"11111111",
  20001=>"11111111",
  20002=>"00000011",
  20003=>"11111111",
  20004=>"00000101",
  20005=>"00000010",
  20006=>"11111111",
  20007=>"11111110",
  20008=>"11111101",
  20009=>"00000100",
  20010=>"00000011",
  20011=>"11111100",
  20012=>"00000001",
  20013=>"00000000",
  20014=>"00000011",
  20015=>"00000001",
  20016=>"11111111",
  20017=>"00000011",
  20018=>"00000001",
  20019=>"00000010",
  20020=>"00000000",
  20021=>"00000101",
  20022=>"00000001",
  20023=>"11111100",
  20024=>"00000010",
  20025=>"00000100",
  20026=>"11111110",
  20027=>"00000010",
  20028=>"11111111",
  20029=>"00000000",
  20030=>"00000001",
  20031=>"00000000",
  20032=>"11111101",
  20033=>"11111110",
  20034=>"00000011",
  20035=>"00000100",
  20036=>"00000001",
  20037=>"11111111",
  20038=>"11111110",
  20039=>"00000100",
  20040=>"11111110",
  20041=>"00000011",
  20042=>"00000100",
  20043=>"00000010",
  20044=>"00000000",
  20045=>"00000000",
  20046=>"11111110",
  20047=>"11111110",
  20048=>"11111111",
  20049=>"11111101",
  20050=>"00000001",
  20051=>"00000001",
  20052=>"00000100",
  20053=>"11111110",
  20054=>"00000011",
  20055=>"00000011",
  20056=>"11111101",
  20057=>"00000011",
  20058=>"11111111",
  20059=>"00000011",
  20060=>"00000001",
  20061=>"00000100",
  20062=>"00000001",
  20063=>"00000000",
  20064=>"00000011",
  20065=>"11111110",
  20066=>"00000000",
  20067=>"00000001",
  20068=>"11111111",
  20069=>"11111111",
  20070=>"11111111",
  20071=>"00000010",
  20072=>"11111110",
  20073=>"11111110",
  20074=>"11111101",
  20075=>"11111101",
  20076=>"00000010",
  20077=>"11111110",
  20078=>"11111111",
  20079=>"00000100",
  20080=>"00000001",
  20081=>"11111100",
  20082=>"00000001",
  20083=>"00000001",
  20084=>"00000000",
  20085=>"00000010",
  20086=>"00000011",
  20087=>"00000001",
  20088=>"00000000",
  20089=>"00000001",
  20090=>"00000000",
  20091=>"00000011",
  20092=>"11111111",
  20093=>"00000010",
  20094=>"11111111",
  20095=>"11111101",
  20096=>"11111101",
  20097=>"00000001",
  20098=>"11111111",
  20099=>"00000001",
  20100=>"00000100",
  20101=>"00000101",
  20102=>"00000011",
  20103=>"11111110",
  20104=>"00000010",
  20105=>"11111110",
  20106=>"11111110",
  20107=>"11111110",
  20108=>"11111111",
  20109=>"00000010",
  20110=>"11111111",
  20111=>"00000000",
  20112=>"00000110",
  20113=>"11111100",
  20114=>"00000100",
  20115=>"00000000",
  20116=>"11111110",
  20117=>"00000010",
  20118=>"11111100",
  20119=>"00000010",
  20120=>"11111011",
  20121=>"00000001",
  20122=>"00000001",
  20123=>"11111011",
  20124=>"00000010",
  20125=>"00000101",
  20126=>"11111101",
  20127=>"11111111",
  20128=>"11111111",
  20129=>"00000010",
  20130=>"00000000",
  20131=>"00000001",
  20132=>"00000001",
  20133=>"00000011",
  20134=>"00000011",
  20135=>"00000000",
  20136=>"00000101",
  20137=>"00000100",
  20138=>"00000000",
  20139=>"11111110",
  20140=>"00000011",
  20141=>"11111101",
  20142=>"00000010",
  20143=>"00000001",
  20144=>"11111101",
  20145=>"00000010",
  20146=>"11111011",
  20147=>"00000010",
  20148=>"11111110",
  20149=>"11111111",
  20150=>"11111110",
  20151=>"00000001",
  20152=>"00000110",
  20153=>"00000111",
  20154=>"00000010",
  20155=>"11111111",
  20156=>"00000010",
  20157=>"00000010",
  20158=>"00000000",
  20159=>"11111111",
  20160=>"11111111",
  20161=>"00000011",
  20162=>"00000001",
  20163=>"00000101",
  20164=>"11111111",
  20165=>"11111100",
  20166=>"00000100",
  20167=>"11111111",
  20168=>"11111101",
  20169=>"00000001",
  20170=>"00000010",
  20171=>"00000100",
  20172=>"00000011",
  20173=>"11111110",
  20174=>"11111111",
  20175=>"00000011",
  20176=>"00000010",
  20177=>"00000011",
  20178=>"11111111",
  20179=>"11111110",
  20180=>"00000011",
  20181=>"00000010",
  20182=>"00000101",
  20183=>"00000100",
  20184=>"00000000",
  20185=>"11111111",
  20186=>"11111110",
  20187=>"11111110",
  20188=>"11111100",
  20189=>"00000001",
  20190=>"11111111",
  20191=>"00000010",
  20192=>"00000001",
  20193=>"00000100",
  20194=>"11111111",
  20195=>"00000001",
  20196=>"11111011",
  20197=>"11111111",
  20198=>"11111101",
  20199=>"11111101",
  20200=>"00000011",
  20201=>"00000000",
  20202=>"00000100",
  20203=>"00000010",
  20204=>"00000001",
  20205=>"11111111",
  20206=>"00000000",
  20207=>"00000011",
  20208=>"11111100",
  20209=>"00000000",
  20210=>"11111111",
  20211=>"11111100",
  20212=>"00000001",
  20213=>"11111110",
  20214=>"00000101",
  20215=>"00000010",
  20216=>"00000000",
  20217=>"00000111",
  20218=>"11111101",
  20219=>"00000011",
  20220=>"00000010",
  20221=>"00000001",
  20222=>"11111001",
  20223=>"11111011",
  20224=>"00000000",
  20225=>"11111110",
  20226=>"00000101",
  20227=>"00000001",
  20228=>"00000010",
  20229=>"00000100",
  20230=>"00000011",
  20231=>"00000000",
  20232=>"00000010",
  20233=>"00000010",
  20234=>"11111100",
  20235=>"11111110",
  20236=>"11111100",
  20237=>"00000000",
  20238=>"11111111",
  20239=>"11111110",
  20240=>"00000000",
  20241=>"11111100",
  20242=>"00000000",
  20243=>"00000011",
  20244=>"00000001",
  20245=>"11111101",
  20246=>"00000000",
  20247=>"00000001",
  20248=>"11111110",
  20249=>"00000010",
  20250=>"00000001",
  20251=>"00000010",
  20252=>"11111111",
  20253=>"00000011",
  20254=>"00000100",
  20255=>"00000011",
  20256=>"00000101",
  20257=>"00000100",
  20258=>"11111110",
  20259=>"00000001",
  20260=>"00000101",
  20261=>"00000100",
  20262=>"00000011",
  20263=>"00000000",
  20264=>"11111111",
  20265=>"00000100",
  20266=>"00000011",
  20267=>"00000010",
  20268=>"00000000",
  20269=>"00000100",
  20270=>"00000000",
  20271=>"00000001",
  20272=>"11111011",
  20273=>"00000011",
  20274=>"00000001",
  20275=>"00000000",
  20276=>"11111101",
  20277=>"00000100",
  20278=>"11111111",
  20279=>"11111110",
  20280=>"00000001",
  20281=>"00000001",
  20282=>"11111101",
  20283=>"00000010",
  20284=>"11111110",
  20285=>"11111101",
  20286=>"00000001",
  20287=>"11111101",
  20288=>"00000100",
  20289=>"00000000",
  20290=>"00000000",
  20291=>"00000100",
  20292=>"00000000",
  20293=>"11111111",
  20294=>"11111101",
  20295=>"00000011",
  20296=>"11111110",
  20297=>"00000101",
  20298=>"11111111",
  20299=>"11111101",
  20300=>"00000010",
  20301=>"11111101",
  20302=>"00000001",
  20303=>"00000011",
  20304=>"11111110",
  20305=>"11111011",
  20306=>"00000001",
  20307=>"11111110",
  20308=>"00000011",
  20309=>"00000011",
  20310=>"11111111",
  20311=>"00000010",
  20312=>"00000001",
  20313=>"11111110",
  20314=>"11111111",
  20315=>"00000001",
  20316=>"00000001",
  20317=>"00000001",
  20318=>"00000000",
  20319=>"00000000",
  20320=>"11111111",
  20321=>"11111111",
  20322=>"11111111",
  20323=>"00000001",
  20324=>"11111111",
  20325=>"11111110",
  20326=>"00000011",
  20327=>"00000011",
  20328=>"00000010",
  20329=>"11111110",
  20330=>"00000001",
  20331=>"11111111",
  20332=>"00000000",
  20333=>"00000011",
  20334=>"11111111",
  20335=>"11111111",
  20336=>"00000001",
  20337=>"11111111",
  20338=>"00000001",
  20339=>"00000011",
  20340=>"11111110",
  20341=>"00000010",
  20342=>"11111110",
  20343=>"11111111",
  20344=>"00000001",
  20345=>"00000000",
  20346=>"11111101",
  20347=>"00000111",
  20348=>"00000000",
  20349=>"00000110",
  20350=>"11111111",
  20351=>"00000010",
  20352=>"11111111",
  20353=>"11111110",
  20354=>"00000000",
  20355=>"00000101",
  20356=>"00000101",
  20357=>"11111110",
  20358=>"00000010",
  20359=>"11111110",
  20360=>"00000000",
  20361=>"00000000",
  20362=>"00000000",
  20363=>"00000001",
  20364=>"11111110",
  20365=>"00000010",
  20366=>"11111100",
  20367=>"00000100",
  20368=>"11111101",
  20369=>"00000100",
  20370=>"11111111",
  20371=>"11111111",
  20372=>"00000000",
  20373=>"00000100",
  20374=>"00000011",
  20375=>"00000100",
  20376=>"11111101",
  20377=>"00000110",
  20378=>"00000011",
  20379=>"11111111",
  20380=>"00000110",
  20381=>"00000100",
  20382=>"00000000",
  20383=>"11111101",
  20384=>"11111111",
  20385=>"11111111",
  20386=>"11111110",
  20387=>"11111110",
  20388=>"00000101",
  20389=>"00000100",
  20390=>"11111111",
  20391=>"00000000",
  20392=>"11111110",
  20393=>"11111101",
  20394=>"11111110",
  20395=>"11111110",
  20396=>"00000011",
  20397=>"11111111",
  20398=>"11111110",
  20399=>"00000010",
  20400=>"11111101",
  20401=>"00000010",
  20402=>"11111011",
  20403=>"00000000",
  20404=>"00000001",
  20405=>"00000010",
  20406=>"00000001",
  20407=>"00000001",
  20408=>"00000100",
  20409=>"11111110",
  20410=>"11111111",
  20411=>"00000010",
  20412=>"00000000",
  20413=>"00000000",
  20414=>"11111100",
  20415=>"00000010",
  20416=>"11111100",
  20417=>"11111101",
  20418=>"00000011",
  20419=>"11111100",
  20420=>"11111101",
  20421=>"11111111",
  20422=>"00000001",
  20423=>"11111110",
  20424=>"00000000",
  20425=>"00000001",
  20426=>"00000000",
  20427=>"00000000",
  20428=>"11111101",
  20429=>"00000010",
  20430=>"00000001",
  20431=>"11111110",
  20432=>"00000001",
  20433=>"00000011",
  20434=>"00000011",
  20435=>"11111110",
  20436=>"00000100",
  20437=>"11111101",
  20438=>"00000101",
  20439=>"00000000",
  20440=>"00000000",
  20441=>"00000000",
  20442=>"11111110",
  20443=>"00000010",
  20444=>"00000011",
  20445=>"11111101",
  20446=>"11111110",
  20447=>"00000011",
  20448=>"11111111",
  20449=>"11111111",
  20450=>"00000100",
  20451=>"00000000",
  20452=>"00000010",
  20453=>"00000000",
  20454=>"00000011",
  20455=>"00000010",
  20456=>"11111010",
  20457=>"11111110",
  20458=>"00000010",
  20459=>"11111101",
  20460=>"11111011",
  20461=>"00000010",
  20462=>"11111111",
  20463=>"00000001",
  20464=>"00000011",
  20465=>"00000011",
  20466=>"00000101",
  20467=>"11111101",
  20468=>"11111110",
  20469=>"00000010",
  20470=>"00000010",
  20471=>"00000001",
  20472=>"11111010",
  20473=>"00000001",
  20474=>"11111111",
  20475=>"00000011",
  20476=>"00000011",
  20477=>"00000010",
  20478=>"00000001",
  20479=>"00000000",
  20480=>"00000011",
  20481=>"11111111",
  20482=>"00000001",
  20483=>"00000000",
  20484=>"00000010",
  20485=>"11111110",
  20486=>"11111111",
  20487=>"11111110",
  20488=>"00000011",
  20489=>"11111111",
  20490=>"11111101",
  20491=>"00000011",
  20492=>"11111101",
  20493=>"11111110",
  20494=>"00000001",
  20495=>"00000000",
  20496=>"11111110",
  20497=>"00000000",
  20498=>"00000010",
  20499=>"00000000",
  20500=>"11111111",
  20501=>"11111111",
  20502=>"11111101",
  20503=>"11111110",
  20504=>"00000111",
  20505=>"00000000",
  20506=>"00000011",
  20507=>"00000001",
  20508=>"11111110",
  20509=>"00000000",
  20510=>"00000011",
  20511=>"11111110",
  20512=>"00000100",
  20513=>"00000010",
  20514=>"00000001",
  20515=>"00000100",
  20516=>"11111111",
  20517=>"11111110",
  20518=>"00000010",
  20519=>"00000010",
  20520=>"00000000",
  20521=>"00000101",
  20522=>"00000000",
  20523=>"00000010",
  20524=>"11111111",
  20525=>"11111101",
  20526=>"11111110",
  20527=>"00000000",
  20528=>"00000010",
  20529=>"11111101",
  20530=>"00000100",
  20531=>"00000001",
  20532=>"00000000",
  20533=>"11111110",
  20534=>"00000101",
  20535=>"11111111",
  20536=>"00000001",
  20537=>"00000010",
  20538=>"11111101",
  20539=>"00000100",
  20540=>"11111111",
  20541=>"11111110",
  20542=>"11111110",
  20543=>"11111111",
  20544=>"00000110",
  20545=>"00000011",
  20546=>"11111110",
  20547=>"00000010",
  20548=>"11111101",
  20549=>"00000010",
  20550=>"11111110",
  20551=>"00000100",
  20552=>"00000100",
  20553=>"11111100",
  20554=>"11111110",
  20555=>"11111111",
  20556=>"11111111",
  20557=>"00000001",
  20558=>"00000100",
  20559=>"00000010",
  20560=>"00000000",
  20561=>"00000001",
  20562=>"11111110",
  20563=>"00000011",
  20564=>"00000100",
  20565=>"11111111",
  20566=>"11111101",
  20567=>"00000000",
  20568=>"11111110",
  20569=>"11111111",
  20570=>"00000001",
  20571=>"00000010",
  20572=>"11111101",
  20573=>"00000011",
  20574=>"00000100",
  20575=>"00000010",
  20576=>"00000010",
  20577=>"11111100",
  20578=>"00000001",
  20579=>"00000001",
  20580=>"11111011",
  20581=>"11111101",
  20582=>"11111101",
  20583=>"00000110",
  20584=>"11111101",
  20585=>"11111110",
  20586=>"11111101",
  20587=>"11111110",
  20588=>"00000001",
  20589=>"11111110",
  20590=>"00000100",
  20591=>"11111101",
  20592=>"00000011",
  20593=>"11111111",
  20594=>"11111111",
  20595=>"00000011",
  20596=>"00000011",
  20597=>"11111101",
  20598=>"11111110",
  20599=>"11111101",
  20600=>"11111110",
  20601=>"00000110",
  20602=>"00000010",
  20603=>"11111110",
  20604=>"11111110",
  20605=>"00000001",
  20606=>"11111111",
  20607=>"00000000",
  20608=>"00000001",
  20609=>"00000100",
  20610=>"00000000",
  20611=>"00000000",
  20612=>"11111101",
  20613=>"00000000",
  20614=>"00000011",
  20615=>"11111110",
  20616=>"00000010",
  20617=>"00000010",
  20618=>"00000001",
  20619=>"11111111",
  20620=>"00000111",
  20621=>"00000000",
  20622=>"00000010",
  20623=>"00000001",
  20624=>"00000010",
  20625=>"00000001",
  20626=>"00000010",
  20627=>"00000001",
  20628=>"00000101",
  20629=>"11111100",
  20630=>"00000011",
  20631=>"11111110",
  20632=>"00000011",
  20633=>"11111110",
  20634=>"00000100",
  20635=>"11111110",
  20636=>"00000100",
  20637=>"11111011",
  20638=>"11111110",
  20639=>"11111111",
  20640=>"00000010",
  20641=>"00000001",
  20642=>"11111110",
  20643=>"11111011",
  20644=>"00000101",
  20645=>"00000010",
  20646=>"11111110",
  20647=>"00000001",
  20648=>"00000010",
  20649=>"00000001",
  20650=>"11111101",
  20651=>"00000001",
  20652=>"00000000",
  20653=>"00000100",
  20654=>"11111111",
  20655=>"11111101",
  20656=>"00000001",
  20657=>"11111110",
  20658=>"00000100",
  20659=>"11111110",
  20660=>"11111101",
  20661=>"00000001",
  20662=>"00000001",
  20663=>"11111111",
  20664=>"00000011",
  20665=>"11111111",
  20666=>"00000000",
  20667=>"00000010",
  20668=>"11111101",
  20669=>"00000001",
  20670=>"11111110",
  20671=>"11111010",
  20672=>"11111110",
  20673=>"00000000",
  20674=>"11111111",
  20675=>"11111100",
  20676=>"11111111",
  20677=>"11111111",
  20678=>"00000011",
  20679=>"00000010",
  20680=>"11111101",
  20681=>"00000011",
  20682=>"00000000",
  20683=>"11111111",
  20684=>"11111111",
  20685=>"00000000",
  20686=>"00000000",
  20687=>"11111101",
  20688=>"00000011",
  20689=>"11111101",
  20690=>"11111111",
  20691=>"00000011",
  20692=>"00000011",
  20693=>"00000011",
  20694=>"00000101",
  20695=>"00000010",
  20696=>"11111101",
  20697=>"00000001",
  20698=>"00000001",
  20699=>"11111100",
  20700=>"11111110",
  20701=>"11111110",
  20702=>"11111111",
  20703=>"11111101",
  20704=>"00000011",
  20705=>"00000010",
  20706=>"11111111",
  20707=>"00000011",
  20708=>"00000011",
  20709=>"11111111",
  20710=>"00000001",
  20711=>"11111100",
  20712=>"11111110",
  20713=>"00000011",
  20714=>"00000001",
  20715=>"00000010",
  20716=>"11111110",
  20717=>"00000100",
  20718=>"00000010",
  20719=>"00000011",
  20720=>"11111110",
  20721=>"11111110",
  20722=>"00000010",
  20723=>"00000011",
  20724=>"00000100",
  20725=>"00000000",
  20726=>"00000001",
  20727=>"00000010",
  20728=>"11111110",
  20729=>"00000000",
  20730=>"11111110",
  20731=>"11111110",
  20732=>"00000000",
  20733=>"00000000",
  20734=>"11111111",
  20735=>"00000001",
  20736=>"11111100",
  20737=>"00000011",
  20738=>"11111111",
  20739=>"11111101",
  20740=>"00000011",
  20741=>"00000010",
  20742=>"11111101",
  20743=>"11111101",
  20744=>"00000010",
  20745=>"00000000",
  20746=>"00000010",
  20747=>"00000101",
  20748=>"00000000",
  20749=>"00000001",
  20750=>"00000001",
  20751=>"00000001",
  20752=>"00000000",
  20753=>"00000000",
  20754=>"00000011",
  20755=>"00000001",
  20756=>"00000101",
  20757=>"11111111",
  20758=>"11111111",
  20759=>"11111100",
  20760=>"00000010",
  20761=>"00000001",
  20762=>"11111110",
  20763=>"00000001",
  20764=>"11111101",
  20765=>"11111111",
  20766=>"11111101",
  20767=>"11111111",
  20768=>"11111110",
  20769=>"00000000",
  20770=>"00000000",
  20771=>"11111101",
  20772=>"00000000",
  20773=>"00000010",
  20774=>"11111100",
  20775=>"11111101",
  20776=>"11111111",
  20777=>"00000101",
  20778=>"11111100",
  20779=>"11111100",
  20780=>"11111110",
  20781=>"00000010",
  20782=>"00000001",
  20783=>"00000100",
  20784=>"11111101",
  20785=>"11111111",
  20786=>"00000001",
  20787=>"11111110",
  20788=>"00000000",
  20789=>"11111110",
  20790=>"11111100",
  20791=>"00000010",
  20792=>"00000010",
  20793=>"11111110",
  20794=>"11111110",
  20795=>"00000011",
  20796=>"00000010",
  20797=>"11111111",
  20798=>"11111111",
  20799=>"00000010",
  20800=>"00000001",
  20801=>"00000011",
  20802=>"00000010",
  20803=>"00000100",
  20804=>"00000010",
  20805=>"00000010",
  20806=>"11111100",
  20807=>"11111111",
  20808=>"00000011",
  20809=>"11111101",
  20810=>"00000001",
  20811=>"11111101",
  20812=>"00000110",
  20813=>"00000011",
  20814=>"11111100",
  20815=>"11111101",
  20816=>"11111110",
  20817=>"00000000",
  20818=>"11111110",
  20819=>"00000001",
  20820=>"00000000",
  20821=>"11111110",
  20822=>"00000001",
  20823=>"11111101",
  20824=>"00000001",
  20825=>"00000010",
  20826=>"11111110",
  20827=>"11111110",
  20828=>"00000001",
  20829=>"00000001",
  20830=>"11111110",
  20831=>"11111110",
  20832=>"11111111",
  20833=>"11111101",
  20834=>"11111110",
  20835=>"00000000",
  20836=>"00000100",
  20837=>"11111111",
  20838=>"11111111",
  20839=>"00000001",
  20840=>"11111111",
  20841=>"00000101",
  20842=>"00000010",
  20843=>"11111110",
  20844=>"00000010",
  20845=>"00000001",
  20846=>"11111101",
  20847=>"11111110",
  20848=>"11111111",
  20849=>"11111111",
  20850=>"00000001",
  20851=>"00000100",
  20852=>"00000011",
  20853=>"00000000",
  20854=>"11111101",
  20855=>"11111111",
  20856=>"00000111",
  20857=>"11111110",
  20858=>"00000100",
  20859=>"00000001",
  20860=>"00000010",
  20861=>"00000001",
  20862=>"00000011",
  20863=>"11111101",
  20864=>"00000001",
  20865=>"11111101",
  20866=>"00000000",
  20867=>"00000010",
  20868=>"11111111",
  20869=>"11111100",
  20870=>"00000001",
  20871=>"00000011",
  20872=>"00000011",
  20873=>"00000000",
  20874=>"00000001",
  20875=>"00000000",
  20876=>"11111101",
  20877=>"11111101",
  20878=>"00000011",
  20879=>"11111110",
  20880=>"00000000",
  20881=>"00000001",
  20882=>"11111111",
  20883=>"11111110",
  20884=>"11111101",
  20885=>"11111110",
  20886=>"00000001",
  20887=>"11111100",
  20888=>"00000000",
  20889=>"11111110",
  20890=>"00000000",
  20891=>"11111011",
  20892=>"11111100",
  20893=>"00000001",
  20894=>"11111110",
  20895=>"00000100",
  20896=>"00000010",
  20897=>"00000101",
  20898=>"00000001",
  20899=>"00000101",
  20900=>"00000010",
  20901=>"00000001",
  20902=>"00000010",
  20903=>"00000011",
  20904=>"00000000",
  20905=>"11111111",
  20906=>"11111111",
  20907=>"00000100",
  20908=>"00000001",
  20909=>"11111101",
  20910=>"11111110",
  20911=>"00000101",
  20912=>"00000010",
  20913=>"00000001",
  20914=>"11111110",
  20915=>"00000010",
  20916=>"00000001",
  20917=>"11111111",
  20918=>"00000100",
  20919=>"11111010",
  20920=>"00000010",
  20921=>"00000100",
  20922=>"11111110",
  20923=>"00000010",
  20924=>"11111101",
  20925=>"11111111",
  20926=>"00000000",
  20927=>"00000010",
  20928=>"11111101",
  20929=>"00000001",
  20930=>"11111110",
  20931=>"11111100",
  20932=>"00000101",
  20933=>"11111111",
  20934=>"00000100",
  20935=>"00000100",
  20936=>"00000010",
  20937=>"11111100",
  20938=>"00000001",
  20939=>"11111111",
  20940=>"11111101",
  20941=>"00000100",
  20942=>"11111110",
  20943=>"00000101",
  20944=>"00000001",
  20945=>"00000000",
  20946=>"00000001",
  20947=>"11111100",
  20948=>"00000101",
  20949=>"00000011",
  20950=>"11111100",
  20951=>"00000010",
  20952=>"11111111",
  20953=>"11111100",
  20954=>"00000000",
  20955=>"11111110",
  20956=>"00000001",
  20957=>"11111110",
  20958=>"11111110",
  20959=>"00000010",
  20960=>"00000100",
  20961=>"00000101",
  20962=>"00000100",
  20963=>"00000010",
  20964=>"11111110",
  20965=>"00000000",
  20966=>"00000000",
  20967=>"11111110",
  20968=>"11111110",
  20969=>"11111110",
  20970=>"11111110",
  20971=>"00000010",
  20972=>"11111110",
  20973=>"00000001",
  20974=>"11111101",
  20975=>"00000000",
  20976=>"11111101",
  20977=>"11111101",
  20978=>"11111111",
  20979=>"11111011",
  20980=>"00000100",
  20981=>"11111110",
  20982=>"00000010",
  20983=>"11111100",
  20984=>"00000010",
  20985=>"11111111",
  20986=>"11111111",
  20987=>"11111101",
  20988=>"11111111",
  20989=>"00000001",
  20990=>"11111101",
  20991=>"11111101",
  20992=>"00000000",
  20993=>"00000011",
  20994=>"00000011",
  20995=>"00000110",
  20996=>"11111111",
  20997=>"00000000",
  20998=>"00000101",
  20999=>"00000001",
  21000=>"00000000",
  21001=>"11111111",
  21002=>"00000001",
  21003=>"00000001",
  21004=>"00000101",
  21005=>"11111110",
  21006=>"11111101",
  21007=>"11111101",
  21008=>"11111110",
  21009=>"00000011",
  21010=>"11111101",
  21011=>"11111110",
  21012=>"11111011",
  21013=>"00000100",
  21014=>"11111110",
  21015=>"00000011",
  21016=>"11111111",
  21017=>"00000100",
  21018=>"11111100",
  21019=>"00000001",
  21020=>"11111111",
  21021=>"11111100",
  21022=>"00000101",
  21023=>"00000010",
  21024=>"00000010",
  21025=>"00000010",
  21026=>"00000101",
  21027=>"11111110",
  21028=>"00000000",
  21029=>"00000000",
  21030=>"11111110",
  21031=>"00000101",
  21032=>"00000001",
  21033=>"00000010",
  21034=>"00000011",
  21035=>"00000001",
  21036=>"00000110",
  21037=>"00000010",
  21038=>"00000011",
  21039=>"11111101",
  21040=>"11111111",
  21041=>"00000010",
  21042=>"00000000",
  21043=>"00000001",
  21044=>"00000101",
  21045=>"11111111",
  21046=>"11111111",
  21047=>"11111111",
  21048=>"11111110",
  21049=>"11111110",
  21050=>"00000011",
  21051=>"00000011",
  21052=>"00000000",
  21053=>"00000001",
  21054=>"00000101",
  21055=>"00000000",
  21056=>"00000000",
  21057=>"00000000",
  21058=>"00000000",
  21059=>"00000010",
  21060=>"11111110",
  21061=>"00000100",
  21062=>"00000000",
  21063=>"00000010",
  21064=>"00000000",
  21065=>"00000000",
  21066=>"11111111",
  21067=>"11111110",
  21068=>"11111110",
  21069=>"11111111",
  21070=>"00000010",
  21071=>"00000001",
  21072=>"11111110",
  21073=>"00000100",
  21074=>"11111100",
  21075=>"11111101",
  21076=>"00000010",
  21077=>"00000011",
  21078=>"00000000",
  21079=>"11111101",
  21080=>"00000100",
  21081=>"11111110",
  21082=>"00000011",
  21083=>"11111111",
  21084=>"00000011",
  21085=>"00000010",
  21086=>"00000010",
  21087=>"11111111",
  21088=>"00000000",
  21089=>"11111100",
  21090=>"11111101",
  21091=>"00000001",
  21092=>"00000100",
  21093=>"00000011",
  21094=>"00000001",
  21095=>"11111110",
  21096=>"11111110",
  21097=>"00000011",
  21098=>"00000001",
  21099=>"11111110",
  21100=>"11111111",
  21101=>"11111101",
  21102=>"00000011",
  21103=>"00000010",
  21104=>"11111011",
  21105=>"00000100",
  21106=>"00000010",
  21107=>"00000010",
  21108=>"11111111",
  21109=>"11111100",
  21110=>"00000100",
  21111=>"00000000",
  21112=>"11111101",
  21113=>"00000011",
  21114=>"00000001",
  21115=>"11111110",
  21116=>"11111111",
  21117=>"00000001",
  21118=>"11111111",
  21119=>"00000001",
  21120=>"00000001",
  21121=>"11111111",
  21122=>"11111111",
  21123=>"00000010",
  21124=>"00000000",
  21125=>"00000000",
  21126=>"00000100",
  21127=>"00000010",
  21128=>"00000100",
  21129=>"00000000",
  21130=>"00000100",
  21131=>"11111110",
  21132=>"00000010",
  21133=>"00000001",
  21134=>"00000010",
  21135=>"00000010",
  21136=>"00000001",
  21137=>"00000001",
  21138=>"11111111",
  21139=>"11111101",
  21140=>"00000011",
  21141=>"11111101",
  21142=>"11111111",
  21143=>"00000010",
  21144=>"00000010",
  21145=>"11111101",
  21146=>"00000011",
  21147=>"11111101",
  21148=>"00000100",
  21149=>"11111111",
  21150=>"11111101",
  21151=>"11111111",
  21152=>"00000100",
  21153=>"11111111",
  21154=>"11111101",
  21155=>"11111110",
  21156=>"00000000",
  21157=>"11111100",
  21158=>"00000101",
  21159=>"11111110",
  21160=>"00000010",
  21161=>"11111111",
  21162=>"11111111",
  21163=>"11111111",
  21164=>"00000000",
  21165=>"11111101",
  21166=>"11111101",
  21167=>"00000011",
  21168=>"00000010",
  21169=>"11111111",
  21170=>"00000011",
  21171=>"11111111",
  21172=>"00000000",
  21173=>"11111110",
  21174=>"00000001",
  21175=>"11111100",
  21176=>"11111111",
  21177=>"11111110",
  21178=>"11111111",
  21179=>"11111111",
  21180=>"00000001",
  21181=>"00000000",
  21182=>"00000101",
  21183=>"00000000",
  21184=>"11111100",
  21185=>"11111110",
  21186=>"00000010",
  21187=>"11111110",
  21188=>"11111101",
  21189=>"00000100",
  21190=>"00000001",
  21191=>"00000011",
  21192=>"00000000",
  21193=>"11111100",
  21194=>"11111101",
  21195=>"00000010",
  21196=>"11111101",
  21197=>"11111110",
  21198=>"00000010",
  21199=>"00000010",
  21200=>"00000000",
  21201=>"00000011",
  21202=>"00000000",
  21203=>"00000011",
  21204=>"00000010",
  21205=>"00000000",
  21206=>"11111110",
  21207=>"00000001",
  21208=>"11111110",
  21209=>"11111111",
  21210=>"11111100",
  21211=>"00000100",
  21212=>"00000101",
  21213=>"00000101",
  21214=>"11111101",
  21215=>"11111101",
  21216=>"11111100",
  21217=>"11111101",
  21218=>"11111111",
  21219=>"11111111",
  21220=>"11111101",
  21221=>"11111110",
  21222=>"11111110",
  21223=>"00000001",
  21224=>"11111110",
  21225=>"11111110",
  21226=>"11111111",
  21227=>"11111111",
  21228=>"00000000",
  21229=>"11111101",
  21230=>"11111111",
  21231=>"11111101",
  21232=>"00000010",
  21233=>"00000001",
  21234=>"11111101",
  21235=>"00000011",
  21236=>"00000000",
  21237=>"11111111",
  21238=>"11111111",
  21239=>"00000011",
  21240=>"00000010",
  21241=>"11111111",
  21242=>"11111111",
  21243=>"00000011",
  21244=>"11111111",
  21245=>"11111011",
  21246=>"00000100",
  21247=>"00000011",
  21248=>"11111111",
  21249=>"00000000",
  21250=>"00000100",
  21251=>"11111101",
  21252=>"11111110",
  21253=>"00000011",
  21254=>"00000011",
  21255=>"00000001",
  21256=>"11111110",
  21257=>"11111110",
  21258=>"00000010",
  21259=>"00000110",
  21260=>"11111110",
  21261=>"00000011",
  21262=>"11111011",
  21263=>"11111110",
  21264=>"00000000",
  21265=>"11111110",
  21266=>"00000100",
  21267=>"11111110",
  21268=>"00000000",
  21269=>"00000000",
  21270=>"00000011",
  21271=>"11111101",
  21272=>"00000000",
  21273=>"11111111",
  21274=>"00000010",
  21275=>"11111100",
  21276=>"00000010",
  21277=>"00000010",
  21278=>"00000010",
  21279=>"00000010",
  21280=>"00000100",
  21281=>"00000000",
  21282=>"11111110",
  21283=>"11111110",
  21284=>"11111111",
  21285=>"11111100",
  21286=>"00000001",
  21287=>"00000010",
  21288=>"11111111",
  21289=>"11111110",
  21290=>"00000000",
  21291=>"00000011",
  21292=>"11111110",
  21293=>"00000010",
  21294=>"00000010",
  21295=>"00000011",
  21296=>"00000011",
  21297=>"00000010",
  21298=>"00000011",
  21299=>"00000000",
  21300=>"00000000",
  21301=>"00000100",
  21302=>"00000010",
  21303=>"00000110",
  21304=>"11111110",
  21305=>"00000000",
  21306=>"11111111",
  21307=>"00000001",
  21308=>"11111101",
  21309=>"00000001",
  21310=>"00000001",
  21311=>"11111101",
  21312=>"11111110",
  21313=>"00000000",
  21314=>"11111111",
  21315=>"00000110",
  21316=>"00000011",
  21317=>"00000010",
  21318=>"11111111",
  21319=>"00000101",
  21320=>"11111110",
  21321=>"11111100",
  21322=>"00000001",
  21323=>"00000000",
  21324=>"00000010",
  21325=>"00000001",
  21326=>"00000100",
  21327=>"00000001",
  21328=>"00000000",
  21329=>"00000010",
  21330=>"11111101",
  21331=>"00000110",
  21332=>"00000001",
  21333=>"00000000",
  21334=>"00000010",
  21335=>"00000001",
  21336=>"11111101",
  21337=>"00000001",
  21338=>"11111111",
  21339=>"11111110",
  21340=>"00000001",
  21341=>"00000011",
  21342=>"11111110",
  21343=>"00000001",
  21344=>"11111110",
  21345=>"00000001",
  21346=>"00000010",
  21347=>"00000011",
  21348=>"00000000",
  21349=>"00000100",
  21350=>"00000100",
  21351=>"00000000",
  21352=>"00000111",
  21353=>"11111110",
  21354=>"00000100",
  21355=>"00000011",
  21356=>"11111101",
  21357=>"00000010",
  21358=>"11111111",
  21359=>"11111111",
  21360=>"00000000",
  21361=>"11111110",
  21362=>"00000000",
  21363=>"11111100",
  21364=>"00000100",
  21365=>"11111100",
  21366=>"00000101",
  21367=>"11111101",
  21368=>"00000001",
  21369=>"11111111",
  21370=>"00000000",
  21371=>"00000000",
  21372=>"11111110",
  21373=>"00000110",
  21374=>"11111111",
  21375=>"00000010",
  21376=>"00000001",
  21377=>"00000001",
  21378=>"00000000",
  21379=>"11111100",
  21380=>"00000000",
  21381=>"11111111",
  21382=>"00000000",
  21383=>"00000000",
  21384=>"00000010",
  21385=>"11111110",
  21386=>"11111110",
  21387=>"00000011",
  21388=>"11111100",
  21389=>"00000000",
  21390=>"00000000",
  21391=>"00000001",
  21392=>"00000001",
  21393=>"00000101",
  21394=>"11111111",
  21395=>"00000011",
  21396=>"00000100",
  21397=>"00000001",
  21398=>"00000101",
  21399=>"00000100",
  21400=>"00000001",
  21401=>"11111111",
  21402=>"00000001",
  21403=>"00000001",
  21404=>"11111110",
  21405=>"00000001",
  21406=>"00000000",
  21407=>"00000101",
  21408=>"00000010",
  21409=>"00000011",
  21410=>"11111101",
  21411=>"00000000",
  21412=>"11111110",
  21413=>"00000100",
  21414=>"11111110",
  21415=>"11111011",
  21416=>"11111111",
  21417=>"00000000",
  21418=>"00000100",
  21419=>"11111110",
  21420=>"00000011",
  21421=>"00000000",
  21422=>"00000011",
  21423=>"00000010",
  21424=>"11111110",
  21425=>"11111100",
  21426=>"11111110",
  21427=>"11111101",
  21428=>"00000000",
  21429=>"11111110",
  21430=>"00000110",
  21431=>"11111110",
  21432=>"00000011",
  21433=>"00000010",
  21434=>"11111100",
  21435=>"11111101",
  21436=>"11111110",
  21437=>"11111101",
  21438=>"00000011",
  21439=>"11111110",
  21440=>"11111101",
  21441=>"00000100",
  21442=>"00000010",
  21443=>"00000000",
  21444=>"00000011",
  21445=>"00000101",
  21446=>"11111110",
  21447=>"00000001",
  21448=>"11111101",
  21449=>"00000001",
  21450=>"00000001",
  21451=>"00000010",
  21452=>"00000011",
  21453=>"00000000",
  21454=>"00000000",
  21455=>"11111101",
  21456=>"00000001",
  21457=>"11111100",
  21458=>"11111101",
  21459=>"11111100",
  21460=>"11111110",
  21461=>"11111100",
  21462=>"11111111",
  21463=>"11111110",
  21464=>"00000000",
  21465=>"11111110",
  21466=>"11111101",
  21467=>"00000011",
  21468=>"00000010",
  21469=>"11111110",
  21470=>"11111111",
  21471=>"11111110",
  21472=>"00000110",
  21473=>"00000011",
  21474=>"00000000",
  21475=>"00000010",
  21476=>"00000001",
  21477=>"11111100",
  21478=>"00000000",
  21479=>"00000100",
  21480=>"11111110",
  21481=>"11111110",
  21482=>"00000011",
  21483=>"11111110",
  21484=>"00000010",
  21485=>"11111111",
  21486=>"11111110",
  21487=>"11111110",
  21488=>"11111111",
  21489=>"00000000",
  21490=>"00000011",
  21491=>"00000010",
  21492=>"00000001",
  21493=>"00000010",
  21494=>"00000011",
  21495=>"11111100",
  21496=>"11111110",
  21497=>"00000011",
  21498=>"11111110",
  21499=>"00000010",
  21500=>"00000000",
  21501=>"11111111",
  21502=>"00000101",
  21503=>"00000010",
  21504=>"11111110",
  21505=>"11111111",
  21506=>"11111111",
  21507=>"00000010",
  21508=>"11111111",
  21509=>"00000010",
  21510=>"11111110",
  21511=>"11111100",
  21512=>"11111101",
  21513=>"11111101",
  21514=>"11111111",
  21515=>"00000010",
  21516=>"11111111",
  21517=>"00000000",
  21518=>"11111110",
  21519=>"00000010",
  21520=>"00000000",
  21521=>"00000010",
  21522=>"11111101",
  21523=>"00000010",
  21524=>"11111111",
  21525=>"11111101",
  21526=>"11111110",
  21527=>"00000000",
  21528=>"00000001",
  21529=>"11111101",
  21530=>"00000000",
  21531=>"11111111",
  21532=>"00000000",
  21533=>"00000000",
  21534=>"11111111",
  21535=>"00000001",
  21536=>"00000100",
  21537=>"00000011",
  21538=>"11111110",
  21539=>"00000000",
  21540=>"00000001",
  21541=>"00000000",
  21542=>"00000011",
  21543=>"00000010",
  21544=>"00000000",
  21545=>"00000000",
  21546=>"00000001",
  21547=>"11111100",
  21548=>"11111111",
  21549=>"00000100",
  21550=>"00000010",
  21551=>"00000011",
  21552=>"00000000",
  21553=>"11111101",
  21554=>"00000000",
  21555=>"11111101",
  21556=>"11111110",
  21557=>"00000000",
  21558=>"00000001",
  21559=>"00000011",
  21560=>"00000011",
  21561=>"00000000",
  21562=>"11111111",
  21563=>"11111110",
  21564=>"00000011",
  21565=>"00000011",
  21566=>"00000000",
  21567=>"00000010",
  21568=>"00000001",
  21569=>"11111101",
  21570=>"00000000",
  21571=>"11111111",
  21572=>"00000100",
  21573=>"00000001",
  21574=>"11111110",
  21575=>"11111110",
  21576=>"00000000",
  21577=>"00000111",
  21578=>"11111111",
  21579=>"00000011",
  21580=>"00000101",
  21581=>"11111101",
  21582=>"00000001",
  21583=>"00000000",
  21584=>"11111110",
  21585=>"11111110",
  21586=>"00000011",
  21587=>"11111111",
  21588=>"00000010",
  21589=>"00000010",
  21590=>"00000000",
  21591=>"00000000",
  21592=>"11111110",
  21593=>"11111101",
  21594=>"00000001",
  21595=>"11111101",
  21596=>"11111101",
  21597=>"00000000",
  21598=>"00000101",
  21599=>"00000010",
  21600=>"00000000",
  21601=>"11111101",
  21602=>"11111110",
  21603=>"11111111",
  21604=>"11111100",
  21605=>"00000001",
  21606=>"00000010",
  21607=>"11111111",
  21608=>"00000001",
  21609=>"11111101",
  21610=>"00000010",
  21611=>"11111110",
  21612=>"11111101",
  21613=>"11111110",
  21614=>"00000101",
  21615=>"00000001",
  21616=>"11111111",
  21617=>"00000000",
  21618=>"11111110",
  21619=>"00000000",
  21620=>"11111110",
  21621=>"00000011",
  21622=>"00000011",
  21623=>"11111111",
  21624=>"00000001",
  21625=>"11111111",
  21626=>"11111110",
  21627=>"00000100",
  21628=>"11111110",
  21629=>"11111101",
  21630=>"11111111",
  21631=>"00000011",
  21632=>"00000000",
  21633=>"00000010",
  21634=>"11111100",
  21635=>"00000011",
  21636=>"00000000",
  21637=>"00000010",
  21638=>"11111111",
  21639=>"00000100",
  21640=>"11111101",
  21641=>"00000010",
  21642=>"00000001",
  21643=>"11111111",
  21644=>"11111101",
  21645=>"11111111",
  21646=>"11111101",
  21647=>"00000001",
  21648=>"00000100",
  21649=>"11111101",
  21650=>"00000010",
  21651=>"11111110",
  21652=>"00000010",
  21653=>"11111110",
  21654=>"00000000",
  21655=>"11111111",
  21656=>"00000001",
  21657=>"11111101",
  21658=>"11111100",
  21659=>"00000001",
  21660=>"11111111",
  21661=>"11111110",
  21662=>"00000000",
  21663=>"11111101",
  21664=>"11111101",
  21665=>"00000011",
  21666=>"00000010",
  21667=>"11111111",
  21668=>"00000001",
  21669=>"11111110",
  21670=>"11111110",
  21671=>"00000001",
  21672=>"11111100",
  21673=>"11111111",
  21674=>"11111111",
  21675=>"11111110",
  21676=>"00000100",
  21677=>"11111110",
  21678=>"00000000",
  21679=>"00000011",
  21680=>"00000001",
  21681=>"11111110",
  21682=>"11111110",
  21683=>"00000000",
  21684=>"11111111",
  21685=>"00000100",
  21686=>"00000010",
  21687=>"11111101",
  21688=>"00000010",
  21689=>"00000001",
  21690=>"00000001",
  21691=>"11111110",
  21692=>"11111111",
  21693=>"11111111",
  21694=>"11111110",
  21695=>"11111111",
  21696=>"00000010",
  21697=>"11111110",
  21698=>"00000010",
  21699=>"11111111",
  21700=>"11111111",
  21701=>"11111110",
  21702=>"11111101",
  21703=>"11111111",
  21704=>"00000101",
  21705=>"11111111",
  21706=>"00000000",
  21707=>"00000001",
  21708=>"00000001",
  21709=>"11111110",
  21710=>"00000100",
  21711=>"00000001",
  21712=>"11111110",
  21713=>"00000110",
  21714=>"00000001",
  21715=>"00000011",
  21716=>"00000001",
  21717=>"00000000",
  21718=>"11111110",
  21719=>"00000011",
  21720=>"00000001",
  21721=>"00000010",
  21722=>"00000011",
  21723=>"00000010",
  21724=>"11111110",
  21725=>"11111110",
  21726=>"00000001",
  21727=>"11111100",
  21728=>"11111111",
  21729=>"11111111",
  21730=>"00000010",
  21731=>"00000010",
  21732=>"00000001",
  21733=>"00000000",
  21734=>"11111111",
  21735=>"00000001",
  21736=>"00000011",
  21737=>"00000001",
  21738=>"00000001",
  21739=>"00000001",
  21740=>"00000011",
  21741=>"11111111",
  21742=>"11111101",
  21743=>"00000000",
  21744=>"11111111",
  21745=>"00000000",
  21746=>"11111111",
  21747=>"11111101",
  21748=>"11111111",
  21749=>"11111111",
  21750=>"00000000",
  21751=>"11111100",
  21752=>"00000000",
  21753=>"00000000",
  21754=>"11111101",
  21755=>"00000001",
  21756=>"00000010",
  21757=>"11111111",
  21758=>"00000000",
  21759=>"11111110",
  21760=>"00000100",
  21761=>"11111101",
  21762=>"11111110",
  21763=>"00000000",
  21764=>"00000010",
  21765=>"11111110",
  21766=>"11111111",
  21767=>"00000001",
  21768=>"11111100",
  21769=>"11111110",
  21770=>"00000010",
  21771=>"11111101",
  21772=>"00000010",
  21773=>"11111110",
  21774=>"00000011",
  21775=>"00000110",
  21776=>"11111101",
  21777=>"00000011",
  21778=>"11111011",
  21779=>"00000011",
  21780=>"11111110",
  21781=>"00000011",
  21782=>"00000001",
  21783=>"00000010",
  21784=>"00000000",
  21785=>"00000011",
  21786=>"00000001",
  21787=>"11111111",
  21788=>"11111110",
  21789=>"11111101",
  21790=>"00000010",
  21791=>"11111101",
  21792=>"11111111",
  21793=>"00000010",
  21794=>"00000011",
  21795=>"11111100",
  21796=>"11111101",
  21797=>"11111111",
  21798=>"00000010",
  21799=>"11111110",
  21800=>"00000000",
  21801=>"11111100",
  21802=>"11111111",
  21803=>"11111101",
  21804=>"00000000",
  21805=>"00000011",
  21806=>"11111110",
  21807=>"00000101",
  21808=>"00000101",
  21809=>"11111110",
  21810=>"00000000",
  21811=>"11111110",
  21812=>"11111110",
  21813=>"11111111",
  21814=>"11111110",
  21815=>"00000001",
  21816=>"11111110",
  21817=>"00000010",
  21818=>"11111101",
  21819=>"00000000",
  21820=>"00000001",
  21821=>"00000000",
  21822=>"00000000",
  21823=>"11111110",
  21824=>"00000001",
  21825=>"00000011",
  21826=>"11111110",
  21827=>"00000010",
  21828=>"11111110",
  21829=>"00000011",
  21830=>"11111101",
  21831=>"00000001",
  21832=>"11111110",
  21833=>"11111101",
  21834=>"00000011",
  21835=>"00000010",
  21836=>"11111101",
  21837=>"11111100",
  21838=>"11111111",
  21839=>"11111110",
  21840=>"00000001",
  21841=>"11111100",
  21842=>"00000000",
  21843=>"11111111",
  21844=>"00000000",
  21845=>"00000100",
  21846=>"11111101",
  21847=>"00000010",
  21848=>"00000000",
  21849=>"00000001",
  21850=>"11111110",
  21851=>"00000001",
  21852=>"11111110",
  21853=>"00000011",
  21854=>"00000001",
  21855=>"00000010",
  21856=>"00000000",
  21857=>"11111100",
  21858=>"00000000",
  21859=>"00000001",
  21860=>"00000011",
  21861=>"00000001",
  21862=>"00000000",
  21863=>"11111101",
  21864=>"00000010",
  21865=>"00000001",
  21866=>"00000010",
  21867=>"11111110",
  21868=>"00000000",
  21869=>"11111101",
  21870=>"00000010",
  21871=>"00000011",
  21872=>"11111110",
  21873=>"11111110",
  21874=>"00000000",
  21875=>"00000000",
  21876=>"00000110",
  21877=>"00000000",
  21878=>"00000000",
  21879=>"00000000",
  21880=>"00000101",
  21881=>"00000000",
  21882=>"11111110",
  21883=>"11111110",
  21884=>"00000000",
  21885=>"11111110",
  21886=>"00000101",
  21887=>"11111101",
  21888=>"11111110",
  21889=>"11111110",
  21890=>"11111110",
  21891=>"11111100",
  21892=>"00000011",
  21893=>"00000000",
  21894=>"11111100",
  21895=>"00000001",
  21896=>"11111111",
  21897=>"00000001",
  21898=>"11111110",
  21899=>"11111110",
  21900=>"00000110",
  21901=>"00000001",
  21902=>"00000100",
  21903=>"11111110",
  21904=>"00000001",
  21905=>"11111110",
  21906=>"00000111",
  21907=>"00000001",
  21908=>"11111101",
  21909=>"11111110",
  21910=>"00000000",
  21911=>"00000110",
  21912=>"00000001",
  21913=>"00000010",
  21914=>"11111100",
  21915=>"11111110",
  21916=>"00000101",
  21917=>"00000011",
  21918=>"00000010",
  21919=>"00000011",
  21920=>"11111101",
  21921=>"00000001",
  21922=>"00000101",
  21923=>"00000010",
  21924=>"00000010",
  21925=>"00000110",
  21926=>"00000011",
  21927=>"11111101",
  21928=>"00000000",
  21929=>"00000010",
  21930=>"11111110",
  21931=>"00000000",
  21932=>"00000000",
  21933=>"11111101",
  21934=>"00000010",
  21935=>"11111110",
  21936=>"00000000",
  21937=>"00000000",
  21938=>"11111100",
  21939=>"00000001",
  21940=>"11111101",
  21941=>"00000000",
  21942=>"00000000",
  21943=>"00000101",
  21944=>"00000000",
  21945=>"00000000",
  21946=>"11111110",
  21947=>"11111101",
  21948=>"00000001",
  21949=>"00000001",
  21950=>"00000011",
  21951=>"00000010",
  21952=>"00000000",
  21953=>"00000100",
  21954=>"00000000",
  21955=>"11111110",
  21956=>"00000001",
  21957=>"11111101",
  21958=>"11111111",
  21959=>"11111110",
  21960=>"00000100",
  21961=>"00000100",
  21962=>"11111101",
  21963=>"11111111",
  21964=>"00000100",
  21965=>"11111101",
  21966=>"00000001",
  21967=>"11111110",
  21968=>"00000010",
  21969=>"00000001",
  21970=>"11111101",
  21971=>"00000001",
  21972=>"11111111",
  21973=>"00000000",
  21974=>"00000100",
  21975=>"00000000",
  21976=>"11111111",
  21977=>"11111100",
  21978=>"00000000",
  21979=>"00000110",
  21980=>"11111100",
  21981=>"11111111",
  21982=>"11111111",
  21983=>"00000001",
  21984=>"11111111",
  21985=>"00000010",
  21986=>"11111101",
  21987=>"11111101",
  21988=>"00000011",
  21989=>"11111110",
  21990=>"00000001",
  21991=>"00000010",
  21992=>"11111100",
  21993=>"00000010",
  21994=>"11111110",
  21995=>"11111100",
  21996=>"00000000",
  21997=>"11111100",
  21998=>"11111111",
  21999=>"00000001",
  22000=>"00000100",
  22001=>"00000000",
  22002=>"00000000",
  22003=>"11111110",
  22004=>"11111111",
  22005=>"11111111",
  22006=>"00000010",
  22007=>"00000001",
  22008=>"00000001",
  22009=>"00000001",
  22010=>"00000000",
  22011=>"11111111",
  22012=>"11111110",
  22013=>"00000001",
  22014=>"11111101",
  22015=>"00000011",
  22016=>"00000010",
  22017=>"11111101",
  22018=>"11111111",
  22019=>"00000000",
  22020=>"00000001",
  22021=>"11111110",
  22022=>"00000010",
  22023=>"00000100",
  22024=>"00000001",
  22025=>"00001000",
  22026=>"00000100",
  22027=>"11111111",
  22028=>"11111101",
  22029=>"00000000",
  22030=>"00000011",
  22031=>"00000100",
  22032=>"00000101",
  22033=>"11111111",
  22034=>"11111110",
  22035=>"11111101",
  22036=>"00000001",
  22037=>"00000011",
  22038=>"00000011",
  22039=>"11111101",
  22040=>"11111111",
  22041=>"11111110",
  22042=>"00000000",
  22043=>"00000000",
  22044=>"11111110",
  22045=>"00000010",
  22046=>"00000011",
  22047=>"00000101",
  22048=>"00000001",
  22049=>"00000001",
  22050=>"11111111",
  22051=>"11111111",
  22052=>"00000001",
  22053=>"11111111",
  22054=>"11111111",
  22055=>"11111111",
  22056=>"11111111",
  22057=>"11111110",
  22058=>"00000010",
  22059=>"11111111",
  22060=>"00000000",
  22061=>"00000010",
  22062=>"11111101",
  22063=>"11111111",
  22064=>"11111110",
  22065=>"11111111",
  22066=>"00000001",
  22067=>"00000010",
  22068=>"11111111",
  22069=>"00000001",
  22070=>"00000000",
  22071=>"00000001",
  22072=>"11111100",
  22073=>"00000001",
  22074=>"11111110",
  22075=>"11111110",
  22076=>"11111101",
  22077=>"11111110",
  22078=>"11111100",
  22079=>"11111101",
  22080=>"00000010",
  22081=>"00000101",
  22082=>"00000000",
  22083=>"00000001",
  22084=>"11111110",
  22085=>"11111101",
  22086=>"00000001",
  22087=>"00000000",
  22088=>"11111111",
  22089=>"00000001",
  22090=>"00000010",
  22091=>"00000010",
  22092=>"00000011",
  22093=>"11111110",
  22094=>"11111111",
  22095=>"00000001",
  22096=>"00000011",
  22097=>"11111110",
  22098=>"00000101",
  22099=>"00000010",
  22100=>"00000011",
  22101=>"00000001",
  22102=>"00000001",
  22103=>"00000011",
  22104=>"11111111",
  22105=>"00000100",
  22106=>"11111110",
  22107=>"00000100",
  22108=>"11111111",
  22109=>"11111111",
  22110=>"00000010",
  22111=>"00000010",
  22112=>"11111101",
  22113=>"00000001",
  22114=>"11111111",
  22115=>"11111111",
  22116=>"00000000",
  22117=>"11111110",
  22118=>"00000010",
  22119=>"00000010",
  22120=>"00000110",
  22121=>"00000010",
  22122=>"00000001",
  22123=>"00000010",
  22124=>"11111101",
  22125=>"00000000",
  22126=>"11111111",
  22127=>"00000001",
  22128=>"11111110",
  22129=>"11111101",
  22130=>"00000001",
  22131=>"11111101",
  22132=>"11111101",
  22133=>"11111111",
  22134=>"11111101",
  22135=>"11111111",
  22136=>"11111111",
  22137=>"11111101",
  22138=>"11111110",
  22139=>"11111111",
  22140=>"00000001",
  22141=>"11111110",
  22142=>"11111111",
  22143=>"00000001",
  22144=>"00000001",
  22145=>"00000000",
  22146=>"11111100",
  22147=>"11111110",
  22148=>"00000010",
  22149=>"11111100",
  22150=>"11111011",
  22151=>"00000101",
  22152=>"00000011",
  22153=>"00000001",
  22154=>"00000000",
  22155=>"11111100",
  22156=>"00000001",
  22157=>"00000010",
  22158=>"00000010",
  22159=>"11111101",
  22160=>"11111101",
  22161=>"00000011",
  22162=>"11111101",
  22163=>"11111111",
  22164=>"11111101",
  22165=>"11111101",
  22166=>"00000001",
  22167=>"11111110",
  22168=>"11111110",
  22169=>"00000110",
  22170=>"00000011",
  22171=>"00000011",
  22172=>"11111101",
  22173=>"11111101",
  22174=>"00000010",
  22175=>"00000010",
  22176=>"00000010",
  22177=>"11111111",
  22178=>"11111100",
  22179=>"00000000",
  22180=>"00000011",
  22181=>"11111100",
  22182=>"11111111",
  22183=>"11111111",
  22184=>"00000000",
  22185=>"00000010",
  22186=>"00000001",
  22187=>"00000000",
  22188=>"00000011",
  22189=>"00000001",
  22190=>"11111111",
  22191=>"00000010",
  22192=>"11111110",
  22193=>"00000001",
  22194=>"00000101",
  22195=>"11111101",
  22196=>"00000010",
  22197=>"11111111",
  22198=>"00000000",
  22199=>"11111111",
  22200=>"11111110",
  22201=>"11111110",
  22202=>"11111101",
  22203=>"00000010",
  22204=>"00000000",
  22205=>"11111111",
  22206=>"11111110",
  22207=>"11111110",
  22208=>"00000010",
  22209=>"11111110",
  22210=>"00000011",
  22211=>"11111111",
  22212=>"11111110",
  22213=>"00000001",
  22214=>"11111110",
  22215=>"00000011",
  22216=>"11111111",
  22217=>"00000001",
  22218=>"11111111",
  22219=>"11111100",
  22220=>"11111110",
  22221=>"00000101",
  22222=>"00000001",
  22223=>"00000000",
  22224=>"00000001",
  22225=>"00000001",
  22226=>"00000001",
  22227=>"00000001",
  22228=>"00000101",
  22229=>"11111100",
  22230=>"00000010",
  22231=>"11111111",
  22232=>"00000011",
  22233=>"00000001",
  22234=>"00000100",
  22235=>"00000001",
  22236=>"11111101",
  22237=>"11111110",
  22238=>"11111101",
  22239=>"11111110",
  22240=>"11111111",
  22241=>"00000001",
  22242=>"00000010",
  22243=>"00000001",
  22244=>"00000000",
  22245=>"00000010",
  22246=>"00000000",
  22247=>"00000001",
  22248=>"00000000",
  22249=>"11111101",
  22250=>"00000000",
  22251=>"00000010",
  22252=>"00000011",
  22253=>"11111111",
  22254=>"11111110",
  22255=>"00000010",
  22256=>"11111011",
  22257=>"00000011",
  22258=>"11111100",
  22259=>"11111101",
  22260=>"11111011",
  22261=>"00000010",
  22262=>"11111110",
  22263=>"11111110",
  22264=>"11111110",
  22265=>"11111111",
  22266=>"11111110",
  22267=>"00000000",
  22268=>"00000000",
  22269=>"11111100",
  22270=>"00000011",
  22271=>"00000000",
  22272=>"11111110",
  22273=>"00000001",
  22274=>"11111100",
  22275=>"00000010",
  22276=>"11111111",
  22277=>"00000001",
  22278=>"11111111",
  22279=>"11111101",
  22280=>"00000010",
  22281=>"11111110",
  22282=>"00000100",
  22283=>"00000001",
  22284=>"00000010",
  22285=>"11111101",
  22286=>"11111111",
  22287=>"00000010",
  22288=>"11111110",
  22289=>"11111111",
  22290=>"00000000",
  22291=>"11111110",
  22292=>"11111110",
  22293=>"11111101",
  22294=>"00000000",
  22295=>"00000001",
  22296=>"11111110",
  22297=>"00000001",
  22298=>"11111111",
  22299=>"00000000",
  22300=>"11111101",
  22301=>"11111100",
  22302=>"11111100",
  22303=>"11111101",
  22304=>"00000010",
  22305=>"11111110",
  22306=>"00000011",
  22307=>"11111110",
  22308=>"11111110",
  22309=>"11111110",
  22310=>"11111110",
  22311=>"11111101",
  22312=>"00000000",
  22313=>"11111100",
  22314=>"11111100",
  22315=>"11111100",
  22316=>"11111111",
  22317=>"11111111",
  22318=>"00000010",
  22319=>"00000000",
  22320=>"00000101",
  22321=>"11111110",
  22322=>"00000010",
  22323=>"11111110",
  22324=>"00000001",
  22325=>"11111100",
  22326=>"00000010",
  22327=>"00000001",
  22328=>"00000010",
  22329=>"00000001",
  22330=>"11111111",
  22331=>"00000010",
  22332=>"00000001",
  22333=>"00000000",
  22334=>"11111110",
  22335=>"00000000",
  22336=>"00000010",
  22337=>"11111101",
  22338=>"00000001",
  22339=>"00000011",
  22340=>"11111111",
  22341=>"11111110",
  22342=>"11111100",
  22343=>"00000010",
  22344=>"00000001",
  22345=>"11111100",
  22346=>"11111101",
  22347=>"00000001",
  22348=>"00000000",
  22349=>"00000011",
  22350=>"11111101",
  22351=>"00000000",
  22352=>"00000001",
  22353=>"00000011",
  22354=>"11111111",
  22355=>"11111101",
  22356=>"00000011",
  22357=>"00000000",
  22358=>"00000010",
  22359=>"00000010",
  22360=>"11111100",
  22361=>"11111101",
  22362=>"00000001",
  22363=>"00000011",
  22364=>"11111111",
  22365=>"00000100",
  22366=>"11111101",
  22367=>"11111100",
  22368=>"00000010",
  22369=>"00000010",
  22370=>"11111101",
  22371=>"11111111",
  22372=>"11111111",
  22373=>"11111101",
  22374=>"11111110",
  22375=>"00000000",
  22376=>"11111101",
  22377=>"00000010",
  22378=>"00000001",
  22379=>"00000000",
  22380=>"11111111",
  22381=>"00000001",
  22382=>"11111110",
  22383=>"11111011",
  22384=>"11111111",
  22385=>"00000010",
  22386=>"11111101",
  22387=>"11111111",
  22388=>"00000010",
  22389=>"00000101",
  22390=>"11111110",
  22391=>"00000001",
  22392=>"11111100",
  22393=>"00000010",
  22394=>"00000001",
  22395=>"00000000",
  22396=>"00000100",
  22397=>"11111100",
  22398=>"00000100",
  22399=>"00000000",
  22400=>"11111111",
  22401=>"00000101",
  22402=>"11111110",
  22403=>"00000001",
  22404=>"00000010",
  22405=>"00000000",
  22406=>"00000010",
  22407=>"11111101",
  22408=>"00000011",
  22409=>"11111101",
  22410=>"00000001",
  22411=>"00000000",
  22412=>"00000001",
  22413=>"00000110",
  22414=>"00000001",
  22415=>"11111110",
  22416=>"00000011",
  22417=>"00000000",
  22418=>"00000001",
  22419=>"00000000",
  22420=>"11111111",
  22421=>"00000010",
  22422=>"00000000",
  22423=>"00000000",
  22424=>"00000000",
  22425=>"11111100",
  22426=>"00000010",
  22427=>"11111111",
  22428=>"11111100",
  22429=>"00000001",
  22430=>"11111101",
  22431=>"11111110",
  22432=>"11111111",
  22433=>"11111110",
  22434=>"11111101",
  22435=>"00000000",
  22436=>"00000011",
  22437=>"00000000",
  22438=>"00000001",
  22439=>"00000011",
  22440=>"00000001",
  22441=>"11111111",
  22442=>"11111110",
  22443=>"00000000",
  22444=>"11111111",
  22445=>"00000011",
  22446=>"11111110",
  22447=>"11111110",
  22448=>"11111111",
  22449=>"11111100",
  22450=>"00000110",
  22451=>"00000011",
  22452=>"00000001",
  22453=>"11111111",
  22454=>"11111110",
  22455=>"00000000",
  22456=>"11111101",
  22457=>"11111111",
  22458=>"11111101",
  22459=>"11111111",
  22460=>"11111011",
  22461=>"11111111",
  22462=>"00000000",
  22463=>"00000000",
  22464=>"00000101",
  22465=>"00000010",
  22466=>"11111100",
  22467=>"00000000",
  22468=>"11111111",
  22469=>"00000001",
  22470=>"11111111",
  22471=>"11111110",
  22472=>"11111101",
  22473=>"00000000",
  22474=>"11111110",
  22475=>"11111110",
  22476=>"11111111",
  22477=>"00000011",
  22478=>"00000110",
  22479=>"00000010",
  22480=>"00000010",
  22481=>"11111110",
  22482=>"00000001",
  22483=>"00000011",
  22484=>"00000011",
  22485=>"00000100",
  22486=>"11111110",
  22487=>"11111110",
  22488=>"11111110",
  22489=>"00000000",
  22490=>"11111111",
  22491=>"11111110",
  22492=>"00000000",
  22493=>"11111101",
  22494=>"00000100",
  22495=>"00000000",
  22496=>"00000001",
  22497=>"00000010",
  22498=>"00000010",
  22499=>"11111111",
  22500=>"00000010",
  22501=>"11111110",
  22502=>"11111101",
  22503=>"11111111",
  22504=>"00000010",
  22505=>"00000000",
  22506=>"00000001",
  22507=>"11111101",
  22508=>"11111111",
  22509=>"00000010",
  22510=>"11111101",
  22511=>"00000001",
  22512=>"11111101",
  22513=>"00000001",
  22514=>"11111101",
  22515=>"11111100",
  22516=>"00000000",
  22517=>"00000010",
  22518=>"11111101",
  22519=>"00000010",
  22520=>"00000010",
  22521=>"00000000",
  22522=>"11111101",
  22523=>"00000000",
  22524=>"11111111",
  22525=>"00000010",
  22526=>"11111101",
  22527=>"11111110",
  22528=>"00000001",
  22529=>"11111111",
  22530=>"11111111",
  22531=>"11111110",
  22532=>"11111110",
  22533=>"00000001",
  22534=>"00000001",
  22535=>"11111111",
  22536=>"11111110",
  22537=>"00000000",
  22538=>"11111111",
  22539=>"00000000",
  22540=>"11111110",
  22541=>"00000000",
  22542=>"11111101",
  22543=>"11111111",
  22544=>"11111110",
  22545=>"11111110",
  22546=>"11111111",
  22547=>"00000001",
  22548=>"00000000",
  22549=>"00000001",
  22550=>"00000001",
  22551=>"00000001",
  22552=>"11111110",
  22553=>"00000010",
  22554=>"00000000",
  22555=>"00000000",
  22556=>"00000001",
  22557=>"00000000",
  22558=>"00000011",
  22559=>"00000001",
  22560=>"00000000",
  22561=>"11111110",
  22562=>"11111101",
  22563=>"00000011",
  22564=>"00000011",
  22565=>"00000001",
  22566=>"11111101",
  22567=>"11111110",
  22568=>"11111111",
  22569=>"11111111",
  22570=>"00000001",
  22571=>"00000001",
  22572=>"00000010",
  22573=>"00000001",
  22574=>"11111110",
  22575=>"11111110",
  22576=>"00000010",
  22577=>"00000001",
  22578=>"11111101",
  22579=>"00000000",
  22580=>"11111111",
  22581=>"00000001",
  22582=>"11111111",
  22583=>"11111111",
  22584=>"00000000",
  22585=>"00000000",
  22586=>"11111110",
  22587=>"00000000",
  22588=>"11111111",
  22589=>"00000010",
  22590=>"00000000",
  22591=>"00000001",
  22592=>"11111110",
  22593=>"11111111",
  22594=>"00000000",
  22595=>"11111110",
  22596=>"11111101",
  22597=>"00000001",
  22598=>"11111111",
  22599=>"00000001",
  22600=>"11111111",
  22601=>"11111101",
  22602=>"11111111",
  22603=>"11111101",
  22604=>"00000010",
  22605=>"00000000",
  22606=>"11111110",
  22607=>"00000001",
  22608=>"11111110",
  22609=>"11111110",
  22610=>"11111111",
  22611=>"11111111",
  22612=>"00000011",
  22613=>"00000001",
  22614=>"00000011",
  22615=>"00000001",
  22616=>"00000000",
  22617=>"11111101",
  22618=>"00000000",
  22619=>"00000000",
  22620=>"11111101",
  22621=>"00000001",
  22622=>"00000000",
  22623=>"00000000",
  22624=>"11111110",
  22625=>"00000011",
  22626=>"00000011",
  22627=>"00000000",
  22628=>"11111111",
  22629=>"00000010",
  22630=>"00000010",
  22631=>"00000001",
  22632=>"11111111",
  22633=>"11111110",
  22634=>"00000001",
  22635=>"00000010",
  22636=>"00000001",
  22637=>"00000001",
  22638=>"00000001",
  22639=>"00000000",
  22640=>"11111101",
  22641=>"11111110",
  22642=>"11111110",
  22643=>"11111101",
  22644=>"11111100",
  22645=>"11111110",
  22646=>"00000000",
  22647=>"11111111",
  22648=>"11111111",
  22649=>"11111101",
  22650=>"11111101",
  22651=>"11111110",
  22652=>"00000010",
  22653=>"11111110",
  22654=>"00000010",
  22655=>"11111101",
  22656=>"11111111",
  22657=>"11111111",
  22658=>"11111110",
  22659=>"00000001",
  22660=>"11111111",
  22661=>"11111110",
  22662=>"00000001",
  22663=>"00000000",
  22664=>"11111111",
  22665=>"11111111",
  22666=>"00000000",
  22667=>"11111100",
  22668=>"11111110",
  22669=>"11111111",
  22670=>"00000011",
  22671=>"11111111",
  22672=>"00000000",
  22673=>"11111101",
  22674=>"11111110",
  22675=>"00000000",
  22676=>"11111110",
  22677=>"00000010",
  22678=>"11111101",
  22679=>"00000001",
  22680=>"11111101",
  22681=>"11111101",
  22682=>"11111110",
  22683=>"11111101",
  22684=>"11111111",
  22685=>"11111110",
  22686=>"11111110",
  22687=>"00000001",
  22688=>"00000011",
  22689=>"11111111",
  22690=>"00000000",
  22691=>"00000011",
  22692=>"00000010",
  22693=>"11111111",
  22694=>"00000010",
  22695=>"11111111",
  22696=>"00000010",
  22697=>"11111100",
  22698=>"11111111",
  22699=>"00000001",
  22700=>"11111111",
  22701=>"11111101",
  22702=>"11111101",
  22703=>"00000010",
  22704=>"11111111",
  22705=>"11111110",
  22706=>"00000000",
  22707=>"00000100",
  22708=>"11111110",
  22709=>"11111111",
  22710=>"00000010",
  22711=>"11111111",
  22712=>"00000000",
  22713=>"00000010",
  22714=>"11111111",
  22715=>"00000010",
  22716=>"00000011",
  22717=>"00000000",
  22718=>"00000010",
  22719=>"11111111",
  22720=>"00000010",
  22721=>"00000000",
  22722=>"11111111",
  22723=>"00000000",
  22724=>"00000011",
  22725=>"00000011",
  22726=>"00000100",
  22727=>"00000000",
  22728=>"00000001",
  22729=>"11111110",
  22730=>"11111110",
  22731=>"11111110",
  22732=>"00000000",
  22733=>"00000000",
  22734=>"11111111",
  22735=>"00000100",
  22736=>"11111111",
  22737=>"00000001",
  22738=>"00000001",
  22739=>"00000001",
  22740=>"11111111",
  22741=>"11111110",
  22742=>"11111111",
  22743=>"00000001",
  22744=>"11111110",
  22745=>"00000000",
  22746=>"00000001",
  22747=>"11111100",
  22748=>"00000010",
  22749=>"00000010",
  22750=>"11111111",
  22751=>"00000111",
  22752=>"00000010",
  22753=>"00000010",
  22754=>"00000000",
  22755=>"00000010",
  22756=>"00000001",
  22757=>"00000010",
  22758=>"11111110",
  22759=>"00000010",
  22760=>"00000001",
  22761=>"00000000",
  22762=>"00000010",
  22763=>"11111111",
  22764=>"00000001",
  22765=>"11111110",
  22766=>"11111111",
  22767=>"11111111",
  22768=>"00000000",
  22769=>"00000000",
  22770=>"11111110",
  22771=>"00000100",
  22772=>"00000101",
  22773=>"11111110",
  22774=>"00000010",
  22775=>"11111101",
  22776=>"00000001",
  22777=>"00000001",
  22778=>"11111101",
  22779=>"00000001",
  22780=>"11111101",
  22781=>"00000010",
  22782=>"00000001",
  22783=>"00000010",
  22784=>"00000000",
  22785=>"11111110",
  22786=>"00000000",
  22787=>"00000000",
  22788=>"00000001",
  22789=>"00000101",
  22790=>"11111110",
  22791=>"00000010",
  22792=>"11111110",
  22793=>"11111101",
  22794=>"00000001",
  22795=>"00000100",
  22796=>"11111110",
  22797=>"00000010",
  22798=>"11111111",
  22799=>"00000001",
  22800=>"00000000",
  22801=>"00000011",
  22802=>"00000101",
  22803=>"00000000",
  22804=>"00000100",
  22805=>"00000000",
  22806=>"00000001",
  22807=>"00000010",
  22808=>"11111101",
  22809=>"00000000",
  22810=>"11111110",
  22811=>"11111101",
  22812=>"11111110",
  22813=>"00000010",
  22814=>"00000011",
  22815=>"00000000",
  22816=>"11111101",
  22817=>"00000001",
  22818=>"11111101",
  22819=>"00000010",
  22820=>"00000001",
  22821=>"11111110",
  22822=>"11111111",
  22823=>"00000011",
  22824=>"11111110",
  22825=>"11111110",
  22826=>"00000001",
  22827=>"11111110",
  22828=>"11111111",
  22829=>"00000011",
  22830=>"11111110",
  22831=>"00000001",
  22832=>"11111111",
  22833=>"11111101",
  22834=>"11111111",
  22835=>"11111110",
  22836=>"00000010",
  22837=>"00000010",
  22838=>"00000000",
  22839=>"00000000",
  22840=>"00000000",
  22841=>"00000001",
  22842=>"00000000",
  22843=>"00000001",
  22844=>"00000010",
  22845=>"00000001",
  22846=>"11111111",
  22847=>"00000011",
  22848=>"11111111",
  22849=>"11111111",
  22850=>"00000010",
  22851=>"00000010",
  22852=>"00000001",
  22853=>"11111110",
  22854=>"00000001",
  22855=>"00000010",
  22856=>"00000000",
  22857=>"11111101",
  22858=>"00000001",
  22859=>"00000010",
  22860=>"11111100",
  22861=>"00000010",
  22862=>"00000000",
  22863=>"00000000",
  22864=>"00000000",
  22865=>"00000010",
  22866=>"00000001",
  22867=>"11111101",
  22868=>"00000001",
  22869=>"11111111",
  22870=>"00000001",
  22871=>"11111101",
  22872=>"11111110",
  22873=>"00000000",
  22874=>"00000010",
  22875=>"00000001",
  22876=>"11111110",
  22877=>"11111111",
  22878=>"11111110",
  22879=>"11111111",
  22880=>"00000011",
  22881=>"11111101",
  22882=>"11111110",
  22883=>"00000001",
  22884=>"00000000",
  22885=>"00000000",
  22886=>"00000001",
  22887=>"11111110",
  22888=>"00000001",
  22889=>"00000011",
  22890=>"11111101",
  22891=>"00000001",
  22892=>"00000000",
  22893=>"00000000",
  22894=>"11111110",
  22895=>"11111110",
  22896=>"00000001",
  22897=>"11111110",
  22898=>"11111111",
  22899=>"00000001",
  22900=>"00000000",
  22901=>"00000010",
  22902=>"00000001",
  22903=>"00000001",
  22904=>"11111111",
  22905=>"11111111",
  22906=>"11111101",
  22907=>"11111111",
  22908=>"11111110",
  22909=>"11111110",
  22910=>"00000001",
  22911=>"11111101",
  22912=>"11111111",
  22913=>"00000011",
  22914=>"00000001",
  22915=>"00000011",
  22916=>"00000000",
  22917=>"11111111",
  22918=>"00000010",
  22919=>"11111111",
  22920=>"11111111",
  22921=>"00000001",
  22922=>"11111101",
  22923=>"00000001",
  22924=>"00000000",
  22925=>"00000001",
  22926=>"00000010",
  22927=>"00000000",
  22928=>"00000000",
  22929=>"11111101",
  22930=>"00000001",
  22931=>"00000010",
  22932=>"11111101",
  22933=>"00000000",
  22934=>"00000010",
  22935=>"11111111",
  22936=>"00000001",
  22937=>"00000011",
  22938=>"00000010",
  22939=>"00000101",
  22940=>"11111100",
  22941=>"00000001",
  22942=>"11111100",
  22943=>"11111110",
  22944=>"00000010",
  22945=>"00000001",
  22946=>"00000010",
  22947=>"00000001",
  22948=>"11111101",
  22949=>"00000001",
  22950=>"11111111",
  22951=>"00000000",
  22952=>"00000001",
  22953=>"00000000",
  22954=>"11111111",
  22955=>"11111101",
  22956=>"11111110",
  22957=>"11111110",
  22958=>"11111110",
  22959=>"00000010",
  22960=>"11111111",
  22961=>"00000010",
  22962=>"00000000",
  22963=>"00000000",
  22964=>"11111110",
  22965=>"11111110",
  22966=>"00000011",
  22967=>"11111101",
  22968=>"11111110",
  22969=>"00000010",
  22970=>"00000010",
  22971=>"00000000",
  22972=>"00000001",
  22973=>"11111101",
  22974=>"11111111",
  22975=>"00000000",
  22976=>"00000001",
  22977=>"11111111",
  22978=>"00000010",
  22979=>"11111101",
  22980=>"11111110",
  22981=>"00000001",
  22982=>"00000010",
  22983=>"00000010",
  22984=>"11111110",
  22985=>"11111101",
  22986=>"00000011",
  22987=>"11111111",
  22988=>"11111111",
  22989=>"11111110",
  22990=>"00000001",
  22991=>"00000011",
  22992=>"11111101",
  22993=>"11111111",
  22994=>"00000000",
  22995=>"11111101",
  22996=>"00000001",
  22997=>"11111111",
  22998=>"11111101",
  22999=>"00000010",
  23000=>"00000000",
  23001=>"11111101",
  23002=>"11111101",
  23003=>"11111101",
  23004=>"00000000",
  23005=>"11111111",
  23006=>"00000001",
  23007=>"00000001",
  23008=>"00000100",
  23009=>"00000010",
  23010=>"00000010",
  23011=>"11111101",
  23012=>"11111111",
  23013=>"11111111",
  23014=>"00000100",
  23015=>"00000000",
  23016=>"11111111",
  23017=>"00000000",
  23018=>"00000001",
  23019=>"11111100",
  23020=>"00000010",
  23021=>"00000001",
  23022=>"00000001",
  23023=>"00000010",
  23024=>"11111110",
  23025=>"11111110",
  23026=>"00000011",
  23027=>"00000011",
  23028=>"00000001",
  23029=>"11111110",
  23030=>"00000000",
  23031=>"00000011",
  23032=>"11111110",
  23033=>"00000001",
  23034=>"11111101",
  23035=>"11111110",
  23036=>"11111110",
  23037=>"00000011",
  23038=>"11111110",
  23039=>"11111101",
  23040=>"00000001",
  23041=>"11111111",
  23042=>"11111101",
  23043=>"00000001",
  23044=>"00000000",
  23045=>"00000001",
  23046=>"11111110",
  23047=>"11111111",
  23048=>"00000000",
  23049=>"00000000",
  23050=>"11111111",
  23051=>"00000000",
  23052=>"00000100",
  23053=>"11111111",
  23054=>"11111111",
  23055=>"11111101",
  23056=>"00000000",
  23057=>"11111110",
  23058=>"00000011",
  23059=>"11111110",
  23060=>"00000001",
  23061=>"00000000",
  23062=>"11111101",
  23063=>"00000000",
  23064=>"11111111",
  23065=>"11111110",
  23066=>"00000010",
  23067=>"00000000",
  23068=>"11111110",
  23069=>"11111110",
  23070=>"00000001",
  23071=>"00000000",
  23072=>"11111111",
  23073=>"00000001",
  23074=>"00000000",
  23075=>"11111101",
  23076=>"00000011",
  23077=>"00000011",
  23078=>"11111111",
  23079=>"11111101",
  23080=>"11111111",
  23081=>"00000010",
  23082=>"00000000",
  23083=>"11111110",
  23084=>"00000110",
  23085=>"11111110",
  23086=>"11111101",
  23087=>"00000000",
  23088=>"00000000",
  23089=>"11111101",
  23090=>"00000001",
  23091=>"00000001",
  23092=>"00000000",
  23093=>"00000011",
  23094=>"11111111",
  23095=>"00000010",
  23096=>"11111101",
  23097=>"00000000",
  23098=>"00000000",
  23099=>"11111110",
  23100=>"00000001",
  23101=>"11111101",
  23102=>"00000011",
  23103=>"11111110",
  23104=>"00000010",
  23105=>"11111101",
  23106=>"11111110",
  23107=>"00000000",
  23108=>"11111111",
  23109=>"00000000",
  23110=>"00000001",
  23111=>"11111111",
  23112=>"11111111",
  23113=>"11111110",
  23114=>"00000010",
  23115=>"11111110",
  23116=>"00000000",
  23117=>"00000010",
  23118=>"00000010",
  23119=>"00000010",
  23120=>"00000010",
  23121=>"00000000",
  23122=>"00000001",
  23123=>"00000001",
  23124=>"11111110",
  23125=>"11111110",
  23126=>"11111111",
  23127=>"11111101",
  23128=>"00000001",
  23129=>"00000010",
  23130=>"11111111",
  23131=>"11111111",
  23132=>"11111110",
  23133=>"11111100",
  23134=>"00000000",
  23135=>"00000010",
  23136=>"11111111",
  23137=>"00000010",
  23138=>"00000000",
  23139=>"11111111",
  23140=>"11111111",
  23141=>"11111110",
  23142=>"11111110",
  23143=>"00000000",
  23144=>"00000000",
  23145=>"00000001",
  23146=>"00000010",
  23147=>"11111110",
  23148=>"11111111",
  23149=>"00000001",
  23150=>"11111101",
  23151=>"11111111",
  23152=>"11111110",
  23153=>"00000001",
  23154=>"00000001",
  23155=>"00000001",
  23156=>"11111110",
  23157=>"00000000",
  23158=>"00000011",
  23159=>"00000010",
  23160=>"11111110",
  23161=>"11111101",
  23162=>"11111111",
  23163=>"11111110",
  23164=>"11111110",
  23165=>"11111110",
  23166=>"11111110",
  23167=>"11111111",
  23168=>"00000001",
  23169=>"00000001",
  23170=>"11111101",
  23171=>"11111110",
  23172=>"00000001",
  23173=>"11111101",
  23174=>"00000001",
  23175=>"11111110",
  23176=>"00000001",
  23177=>"00000001",
  23178=>"00000001",
  23179=>"11111110",
  23180=>"00000000",
  23181=>"00000000",
  23182=>"00000000",
  23183=>"00000010",
  23184=>"11111111",
  23185=>"11111111",
  23186=>"11111111",
  23187=>"11111111",
  23188=>"00000000",
  23189=>"11111101",
  23190=>"11111111",
  23191=>"11111111",
  23192=>"11111101",
  23193=>"00000001",
  23194=>"00000001",
  23195=>"11111111",
  23196=>"00000001",
  23197=>"00000100",
  23198=>"00000000",
  23199=>"00000000",
  23200=>"11111111",
  23201=>"00000000",
  23202=>"00000000",
  23203=>"11111101",
  23204=>"00000010",
  23205=>"00000010",
  23206=>"11111110",
  23207=>"00000000",
  23208=>"11111110",
  23209=>"00000010",
  23210=>"00000010",
  23211=>"00000010",
  23212=>"11111110",
  23213=>"11111111",
  23214=>"00000001",
  23215=>"00000000",
  23216=>"00000010",
  23217=>"11111101",
  23218=>"00000011",
  23219=>"11111110",
  23220=>"11111111",
  23221=>"11111111",
  23222=>"11111101",
  23223=>"00000001",
  23224=>"00000011",
  23225=>"00000001",
  23226=>"00000000",
  23227=>"00000000",
  23228=>"00000000",
  23229=>"11111110",
  23230=>"11111110",
  23231=>"00000100",
  23232=>"00000010",
  23233=>"11111101",
  23234=>"11111101",
  23235=>"11111111",
  23236=>"00000000",
  23237=>"11111111",
  23238=>"11111110",
  23239=>"00000011",
  23240=>"11111111",
  23241=>"00000100",
  23242=>"00000010",
  23243=>"00000010",
  23244=>"11111110",
  23245=>"00000000",
  23246=>"11111111",
  23247=>"11111101",
  23248=>"00000001",
  23249=>"11111110",
  23250=>"00000001",
  23251=>"00000100",
  23252=>"11111111",
  23253=>"00000001",
  23254=>"11111110",
  23255=>"11111110",
  23256=>"11111111",
  23257=>"00000000",
  23258=>"11111101",
  23259=>"00000100",
  23260=>"00000001",
  23261=>"00000000",
  23262=>"00000100",
  23263=>"00000000",
  23264=>"11111110",
  23265=>"11111101",
  23266=>"11111101",
  23267=>"00000010",
  23268=>"00000000",
  23269=>"11111101",
  23270=>"00000100",
  23271=>"00000001",
  23272=>"11111101",
  23273=>"00000001",
  23274=>"00000001",
  23275=>"11111111",
  23276=>"11111111",
  23277=>"00000010",
  23278=>"00000001",
  23279=>"00000010",
  23280=>"11111111",
  23281=>"11111110",
  23282=>"00000100",
  23283=>"00000000",
  23284=>"00000001",
  23285=>"11111101",
  23286=>"00000001",
  23287=>"00000011",
  23288=>"00000001",
  23289=>"00000001",
  23290=>"00000010",
  23291=>"00000001",
  23292=>"11111110",
  23293=>"00000001",
  23294=>"00001000",
  23295=>"00000001",
  23296=>"00000010",
  23297=>"11111101",
  23298=>"11111110",
  23299=>"00000000",
  23300=>"11111101",
  23301=>"11111110",
  23302=>"11111101",
  23303=>"00000000",
  23304=>"00000111",
  23305=>"00000100",
  23306=>"00000000",
  23307=>"11111110",
  23308=>"11111111",
  23309=>"11111101",
  23310=>"11111101",
  23311=>"00000001",
  23312=>"11111101",
  23313=>"11111110",
  23314=>"11111110",
  23315=>"00000010",
  23316=>"11111110",
  23317=>"00000010",
  23318=>"00000001",
  23319=>"00000011",
  23320=>"00000011",
  23321=>"00000000",
  23322=>"00000000",
  23323=>"11111101",
  23324=>"00000000",
  23325=>"11111111",
  23326=>"00000001",
  23327=>"11111111",
  23328=>"00000000",
  23329=>"11111101",
  23330=>"00000010",
  23331=>"00000001",
  23332=>"11111111",
  23333=>"11111101",
  23334=>"00000010",
  23335=>"00000001",
  23336=>"00000010",
  23337=>"11111110",
  23338=>"11111111",
  23339=>"11111111",
  23340=>"11111111",
  23341=>"11111111",
  23342=>"11111110",
  23343=>"00000000",
  23344=>"00000000",
  23345=>"00000001",
  23346=>"11111110",
  23347=>"00000010",
  23348=>"11111111",
  23349=>"11111101",
  23350=>"00000001",
  23351=>"11111110",
  23352=>"00000001",
  23353=>"11111110",
  23354=>"11111110",
  23355=>"11111111",
  23356=>"00000000",
  23357=>"00000000",
  23358=>"00000010",
  23359=>"00000000",
  23360=>"00000010",
  23361=>"00000010",
  23362=>"00000001",
  23363=>"11111101",
  23364=>"11111110",
  23365=>"00000001",
  23366=>"00000001",
  23367=>"11111101",
  23368=>"11111110",
  23369=>"00000000",
  23370=>"00000000",
  23371=>"11111111",
  23372=>"11111110",
  23373=>"00000010",
  23374=>"00000011",
  23375=>"00000001",
  23376=>"11111111",
  23377=>"11111111",
  23378=>"11111111",
  23379=>"00000000",
  23380=>"00000000",
  23381=>"11111110",
  23382=>"00000001",
  23383=>"11111101",
  23384=>"11111111",
  23385=>"00000001",
  23386=>"11111111",
  23387=>"11111110",
  23388=>"00000001",
  23389=>"11111110",
  23390=>"00000001",
  23391=>"00000000",
  23392=>"11111110",
  23393=>"11111111",
  23394=>"00000000",
  23395=>"11111110",
  23396=>"11111110",
  23397=>"00000010",
  23398=>"11111110",
  23399=>"11111110",
  23400=>"11111111",
  23401=>"11111101",
  23402=>"00000010",
  23403=>"00000000",
  23404=>"00000010",
  23405=>"00000000",
  23406=>"11111111",
  23407=>"11111110",
  23408=>"11111101",
  23409=>"00000010",
  23410=>"00000001",
  23411=>"11111111",
  23412=>"11111110",
  23413=>"11111111",
  23414=>"11111111",
  23415=>"00000001",
  23416=>"11111111",
  23417=>"00000000",
  23418=>"00000001",
  23419=>"11111101",
  23420=>"00000010",
  23421=>"11111111",
  23422=>"00000000",
  23423=>"11111101",
  23424=>"11111101",
  23425=>"11111110",
  23426=>"11111111",
  23427=>"11111110",
  23428=>"00000001",
  23429=>"00000001",
  23430=>"00000000",
  23431=>"11111110",
  23432=>"00000001",
  23433=>"11111110",
  23434=>"00000100",
  23435=>"00000001",
  23436=>"11111101",
  23437=>"11111110",
  23438=>"00000001",
  23439=>"11111101",
  23440=>"11111110",
  23441=>"00000001",
  23442=>"11111110",
  23443=>"11111110",
  23444=>"00000101",
  23445=>"00000101",
  23446=>"00000010",
  23447=>"11111110",
  23448=>"11111110",
  23449=>"00000001",
  23450=>"00000001",
  23451=>"11111110",
  23452=>"11111111",
  23453=>"00000001",
  23454=>"11111111",
  23455=>"00000001",
  23456=>"00000100",
  23457=>"00000010",
  23458=>"00000001",
  23459=>"00000000",
  23460=>"11111111",
  23461=>"11111101",
  23462=>"00000011",
  23463=>"11111111",
  23464=>"11111111",
  23465=>"00000011",
  23466=>"00000011",
  23467=>"00000000",
  23468=>"11111111",
  23469=>"11111111",
  23470=>"00000000",
  23471=>"00000000",
  23472=>"00000001",
  23473=>"00000001",
  23474=>"00000000",
  23475=>"00000001",
  23476=>"00000000",
  23477=>"00000000",
  23478=>"00000010",
  23479=>"00000001",
  23480=>"00000000",
  23481=>"11111110",
  23482=>"11111110",
  23483=>"00000000",
  23484=>"00000010",
  23485=>"11111111",
  23486=>"11111110",
  23487=>"00000000",
  23488=>"11111110",
  23489=>"00000001",
  23490=>"11111101",
  23491=>"00000000",
  23492=>"00000011",
  23493=>"11111101",
  23494=>"00000000",
  23495=>"11111110",
  23496=>"00000010",
  23497=>"00000001",
  23498=>"00000001",
  23499=>"11111110",
  23500=>"00000010",
  23501=>"11111101",
  23502=>"00000000",
  23503=>"00000000",
  23504=>"00000010",
  23505=>"11111101",
  23506=>"11111110",
  23507=>"11111111",
  23508=>"00000001",
  23509=>"11111110",
  23510=>"11111110",
  23511=>"11111110",
  23512=>"11111111",
  23513=>"11111111",
  23514=>"00000101",
  23515=>"11111110",
  23516=>"00000010",
  23517=>"11111100",
  23518=>"00000000",
  23519=>"11111101",
  23520=>"00000001",
  23521=>"00000011",
  23522=>"00000010",
  23523=>"00000001",
  23524=>"00000001",
  23525=>"11111111",
  23526=>"00000001",
  23527=>"00000000",
  23528=>"00000101",
  23529=>"00000000",
  23530=>"00000101",
  23531=>"00000001",
  23532=>"00000000",
  23533=>"11111111",
  23534=>"11111110",
  23535=>"11111111",
  23536=>"00000000",
  23537=>"00000000",
  23538=>"00000010",
  23539=>"11111111",
  23540=>"00000000",
  23541=>"11111101",
  23542=>"00000000",
  23543=>"11111100",
  23544=>"11111110",
  23545=>"00000000",
  23546=>"11111101",
  23547=>"11111101",
  23548=>"00000000",
  23549=>"00000000",
  23550=>"11111111",
  23551=>"00000000",
  23552=>"11111111",
  23553=>"11111101",
  23554=>"00000010",
  23555=>"11111110",
  23556=>"00000000",
  23557=>"00000010",
  23558=>"00000010",
  23559=>"11111110",
  23560=>"11111110",
  23561=>"00000000",
  23562=>"11111101",
  23563=>"00000011",
  23564=>"11111110",
  23565=>"11111111",
  23566=>"11111111",
  23567=>"00000010",
  23568=>"11111101",
  23569=>"11111101",
  23570=>"11111101",
  23571=>"00000010",
  23572=>"11111111",
  23573=>"11111101",
  23574=>"00000011",
  23575=>"00000000",
  23576=>"00000001",
  23577=>"00000001",
  23578=>"00000001",
  23579=>"11111101",
  23580=>"00000000",
  23581=>"11111101",
  23582=>"00000000",
  23583=>"11111100",
  23584=>"11111101",
  23585=>"11111111",
  23586=>"11111101",
  23587=>"00000000",
  23588=>"00000000",
  23589=>"11111101",
  23590=>"11111101",
  23591=>"00000000",
  23592=>"00000010",
  23593=>"11111110",
  23594=>"00000000",
  23595=>"11111100",
  23596=>"00000001",
  23597=>"00000001",
  23598=>"00000010",
  23599=>"00000000",
  23600=>"11111101",
  23601=>"11111110",
  23602=>"00000000",
  23603=>"11111110",
  23604=>"00000000",
  23605=>"11111110",
  23606=>"00000010",
  23607=>"00000011",
  23608=>"11111110",
  23609=>"11111111",
  23610=>"11111110",
  23611=>"00000001",
  23612=>"00000001",
  23613=>"00000010",
  23614=>"00000001",
  23615=>"00000001",
  23616=>"11111110",
  23617=>"00000010",
  23618=>"00000000",
  23619=>"00000001",
  23620=>"00000010",
  23621=>"11111111",
  23622=>"11111111",
  23623=>"00000011",
  23624=>"00000001",
  23625=>"00000010",
  23626=>"00000010",
  23627=>"11111111",
  23628=>"00000001",
  23629=>"00000011",
  23630=>"00000010",
  23631=>"00000001",
  23632=>"11111101",
  23633=>"11111110",
  23634=>"11111100",
  23635=>"00000000",
  23636=>"11111111",
  23637=>"00000010",
  23638=>"11111111",
  23639=>"00000000",
  23640=>"11111110",
  23641=>"00000000",
  23642=>"11111110",
  23643=>"11111110",
  23644=>"11111111",
  23645=>"00000011",
  23646=>"00000010",
  23647=>"00000000",
  23648=>"00000001",
  23649=>"11111111",
  23650=>"11111111",
  23651=>"00000010",
  23652=>"00000011",
  23653=>"00000010",
  23654=>"11111110",
  23655=>"00000000",
  23656=>"00000010",
  23657=>"00000100",
  23658=>"00000001",
  23659=>"11111111",
  23660=>"00000010",
  23661=>"00000100",
  23662=>"11111110",
  23663=>"00000000",
  23664=>"11111110",
  23665=>"11111110",
  23666=>"11111101",
  23667=>"00000001",
  23668=>"11111101",
  23669=>"11111111",
  23670=>"11111111",
  23671=>"11111111",
  23672=>"11111110",
  23673=>"11111111",
  23674=>"00000010",
  23675=>"11111111",
  23676=>"11111111",
  23677=>"11111111",
  23678=>"11111111",
  23679=>"00000100",
  23680=>"00000010",
  23681=>"00000001",
  23682=>"00000001",
  23683=>"00000000",
  23684=>"00000000",
  23685=>"00000001",
  23686=>"00000000",
  23687=>"11111111",
  23688=>"00000011",
  23689=>"11111111",
  23690=>"00000011",
  23691=>"00000000",
  23692=>"11111111",
  23693=>"11111101",
  23694=>"11111110",
  23695=>"11111111",
  23696=>"11111110",
  23697=>"11111110",
  23698=>"11111101",
  23699=>"11111111",
  23700=>"00000000",
  23701=>"11111111",
  23702=>"00000001",
  23703=>"00000010",
  23704=>"00000001",
  23705=>"11111111",
  23706=>"00000001",
  23707=>"00000011",
  23708=>"00000010",
  23709=>"00000100",
  23710=>"00000001",
  23711=>"00000011",
  23712=>"11111111",
  23713=>"11111111",
  23714=>"11111111",
  23715=>"11111101",
  23716=>"11111110",
  23717=>"00000010",
  23718=>"11111111",
  23719=>"00000010",
  23720=>"11111110",
  23721=>"11111101",
  23722=>"11111110",
  23723=>"11111111",
  23724=>"11111101",
  23725=>"00000010",
  23726=>"00000101",
  23727=>"00000000",
  23728=>"00000001",
  23729=>"00000011",
  23730=>"00000100",
  23731=>"11111110",
  23732=>"11111111",
  23733=>"00000001",
  23734=>"11111111",
  23735=>"00001000",
  23736=>"11111110",
  23737=>"00000001",
  23738=>"00000001",
  23739=>"11111101",
  23740=>"00000001",
  23741=>"00000001",
  23742=>"00000010",
  23743=>"11111111",
  23744=>"11111101",
  23745=>"11111111",
  23746=>"11111111",
  23747=>"11111101",
  23748=>"11111110",
  23749=>"00000011",
  23750=>"11111101",
  23751=>"00000000",
  23752=>"11111110",
  23753=>"11111110",
  23754=>"11111101",
  23755=>"11111110",
  23756=>"00000001",
  23757=>"11111101",
  23758=>"00000001",
  23759=>"11111111",
  23760=>"11111100",
  23761=>"00000000",
  23762=>"00000011",
  23763=>"11111111",
  23764=>"11111111",
  23765=>"11111110",
  23766=>"11111110",
  23767=>"00000000",
  23768=>"11111110",
  23769=>"11111101",
  23770=>"00000000",
  23771=>"00000111",
  23772=>"00000001",
  23773=>"11111111",
  23774=>"11111111",
  23775=>"00000000",
  23776=>"00000010",
  23777=>"00000010",
  23778=>"00000010",
  23779=>"00000011",
  23780=>"00000011",
  23781=>"00000010",
  23782=>"00000001",
  23783=>"00000001",
  23784=>"11111111",
  23785=>"00000000",
  23786=>"11111101",
  23787=>"00000011",
  23788=>"00000001",
  23789=>"00000011",
  23790=>"00000000",
  23791=>"00000000",
  23792=>"00000000",
  23793=>"11111110",
  23794=>"00000010",
  23795=>"11111011",
  23796=>"00000001",
  23797=>"11111101",
  23798=>"00000000",
  23799=>"00000011",
  23800=>"11111110",
  23801=>"11111110",
  23802=>"00000011",
  23803=>"00000011",
  23804=>"00000010",
  23805=>"11111110",
  23806=>"00000001",
  23807=>"11111111",
  23808=>"00000010",
  23809=>"00000001",
  23810=>"11111110",
  23811=>"00000010",
  23812=>"00000000",
  23813=>"00000010",
  23814=>"11111111",
  23815=>"00000011",
  23816=>"00000000",
  23817=>"11111111",
  23818=>"00000010",
  23819=>"11111101",
  23820=>"11111111",
  23821=>"11111110",
  23822=>"00000001",
  23823=>"00000011",
  23824=>"00000000",
  23825=>"11111111",
  23826=>"00000101",
  23827=>"11111111",
  23828=>"00000001",
  23829=>"11111111",
  23830=>"11111110",
  23831=>"00000011",
  23832=>"00000001",
  23833=>"11111101",
  23834=>"00000011",
  23835=>"11111110",
  23836=>"11111111",
  23837=>"00000010",
  23838=>"00000000",
  23839=>"11111110",
  23840=>"11111111",
  23841=>"00000001",
  23842=>"00000010",
  23843=>"00000011",
  23844=>"00000000",
  23845=>"11111110",
  23846=>"00000001",
  23847=>"00000010",
  23848=>"00000011",
  23849=>"00000000",
  23850=>"11111100",
  23851=>"00000100",
  23852=>"00000100",
  23853=>"00000000",
  23854=>"00000010",
  23855=>"00000000",
  23856=>"11111111",
  23857=>"00000010",
  23858=>"00000001",
  23859=>"11111110",
  23860=>"11111110",
  23861=>"11111101",
  23862=>"11111101",
  23863=>"00000010",
  23864=>"11111111",
  23865=>"11111101",
  23866=>"11111101",
  23867=>"11111111",
  23868=>"00000000",
  23869=>"00000011",
  23870=>"00000000",
  23871=>"11111110",
  23872=>"11111110",
  23873=>"00000000",
  23874=>"11111110",
  23875=>"00000010",
  23876=>"00000001",
  23877=>"00000001",
  23878=>"00000000",
  23879=>"11111111",
  23880=>"00000000",
  23881=>"00000000",
  23882=>"11111111",
  23883=>"00000000",
  23884=>"11111111",
  23885=>"11111111",
  23886=>"11111101",
  23887=>"00000010",
  23888=>"00000000",
  23889=>"00000011",
  23890=>"11111101",
  23891=>"11111111",
  23892=>"11111101",
  23893=>"11111110",
  23894=>"00000000",
  23895=>"11111101",
  23896=>"11111110",
  23897=>"00000000",
  23898=>"00000000",
  23899=>"11111101",
  23900=>"11111110",
  23901=>"11111110",
  23902=>"11111110",
  23903=>"00000001",
  23904=>"00000010",
  23905=>"11111110",
  23906=>"11111111",
  23907=>"00000000",
  23908=>"11111101",
  23909=>"00000011",
  23910=>"11111101",
  23911=>"00000000",
  23912=>"00000000",
  23913=>"11111111",
  23914=>"11111110",
  23915=>"11111101",
  23916=>"00000001",
  23917=>"11111110",
  23918=>"11111101",
  23919=>"00000011",
  23920=>"11111110",
  23921=>"11111101",
  23922=>"11111111",
  23923=>"11111110",
  23924=>"11111110",
  23925=>"00000011",
  23926=>"00000000",
  23927=>"00000000",
  23928=>"00000000",
  23929=>"11111110",
  23930=>"00000000",
  23931=>"00000010",
  23932=>"00000000",
  23933=>"00000001",
  23934=>"11111110",
  23935=>"11111110",
  23936=>"11111101",
  23937=>"00000000",
  23938=>"11111101",
  23939=>"11111101",
  23940=>"00000001",
  23941=>"11111101",
  23942=>"00000000",
  23943=>"11111110",
  23944=>"00000000",
  23945=>"00000001",
  23946=>"11111111",
  23947=>"11111111",
  23948=>"11111110",
  23949=>"00000000",
  23950=>"11111110",
  23951=>"11111111",
  23952=>"00000000",
  23953=>"00000000",
  23954=>"00000001",
  23955=>"00000011",
  23956=>"00000001",
  23957=>"11111110",
  23958=>"00000000",
  23959=>"11111110",
  23960=>"11111111",
  23961=>"11111111",
  23962=>"11111101",
  23963=>"11111011",
  23964=>"11111101",
  23965=>"11111111",
  23966=>"11111111",
  23967=>"11111101",
  23968=>"11111110",
  23969=>"11111111",
  23970=>"11111110",
  23971=>"00000000",
  23972=>"00000000",
  23973=>"00000010",
  23974=>"00000010",
  23975=>"11111101",
  23976=>"00000001",
  23977=>"11111111",
  23978=>"11111111",
  23979=>"00000010",
  23980=>"00000011",
  23981=>"00000100",
  23982=>"11111111",
  23983=>"11111111",
  23984=>"11111111",
  23985=>"11111101",
  23986=>"00000000",
  23987=>"11111110",
  23988=>"11111111",
  23989=>"00000001",
  23990=>"00000000",
  23991=>"00000000",
  23992=>"11111101",
  23993=>"00000000",
  23994=>"00000101",
  23995=>"11111101",
  23996=>"11111101",
  23997=>"11111110",
  23998=>"11111101",
  23999=>"11111110",
  24000=>"00000001",
  24001=>"11111110",
  24002=>"00000001",
  24003=>"11111110",
  24004=>"11111110",
  24005=>"00000010",
  24006=>"11111101",
  24007=>"11111100",
  24008=>"11111110",
  24009=>"00000000",
  24010=>"11111100",
  24011=>"11111101",
  24012=>"11111110",
  24013=>"11111111",
  24014=>"11111111",
  24015=>"00000100",
  24016=>"00000000",
  24017=>"00000011",
  24018=>"00000010",
  24019=>"00000001",
  24020=>"00000010",
  24021=>"00000001",
  24022=>"00000000",
  24023=>"11111101",
  24024=>"00000010",
  24025=>"11111110",
  24026=>"11111101",
  24027=>"11111101",
  24028=>"00000000",
  24029=>"00000000",
  24030=>"11111110",
  24031=>"11111111",
  24032=>"00000010",
  24033=>"11111100",
  24034=>"00000000",
  24035=>"11111111",
  24036=>"00000001",
  24037=>"00000000",
  24038=>"00000000",
  24039=>"11111110",
  24040=>"11111111",
  24041=>"11111111",
  24042=>"11111110",
  24043=>"00000000",
  24044=>"00000001",
  24045=>"00000010",
  24046=>"00000000",
  24047=>"11111110",
  24048=>"00000010",
  24049=>"11111110",
  24050=>"11111101",
  24051=>"00000011",
  24052=>"00000001",
  24053=>"00000000",
  24054=>"00000001",
  24055=>"00000001",
  24056=>"11111101",
  24057=>"00000011",
  24058=>"00000001",
  24059=>"00000001",
  24060=>"11111111",
  24061=>"00000100",
  24062=>"11111110",
  24063=>"00000000",
  24064=>"00000010",
  24065=>"00000000",
  24066=>"00000000",
  24067=>"00000000",
  24068=>"11111111",
  24069=>"11111011",
  24070=>"00000100",
  24071=>"00000010",
  24072=>"00000000",
  24073=>"00000010",
  24074=>"11111111",
  24075=>"11111110",
  24076=>"00000001",
  24077=>"00000010",
  24078=>"00000000",
  24079=>"11111111",
  24080=>"11111111",
  24081=>"11111111",
  24082=>"00000101",
  24083=>"11111101",
  24084=>"11111101",
  24085=>"00000000",
  24086=>"00000010",
  24087=>"11111110",
  24088=>"00000001",
  24089=>"00000000",
  24090=>"11111100",
  24091=>"11111101",
  24092=>"00000000",
  24093=>"11111101",
  24094=>"11111110",
  24095=>"11111110",
  24096=>"00000010",
  24097=>"00000010",
  24098=>"11111101",
  24099=>"11111101",
  24100=>"11111100",
  24101=>"00000101",
  24102=>"00000010",
  24103=>"00000001",
  24104=>"00000101",
  24105=>"11111111",
  24106=>"00000001",
  24107=>"00000000",
  24108=>"11111110",
  24109=>"11111110",
  24110=>"00000011",
  24111=>"00000000",
  24112=>"00000001",
  24113=>"00000011",
  24114=>"00000010",
  24115=>"11111100",
  24116=>"00000000",
  24117=>"00000000",
  24118=>"11111110",
  24119=>"11111110",
  24120=>"11111100",
  24121=>"11111101",
  24122=>"11111101",
  24123=>"00000001",
  24124=>"11111111",
  24125=>"11111111",
  24126=>"00000001",
  24127=>"11111101",
  24128=>"11111111",
  24129=>"11111101",
  24130=>"11111101",
  24131=>"00000000",
  24132=>"00000010",
  24133=>"11111101",
  24134=>"00000011",
  24135=>"00000011",
  24136=>"11111111",
  24137=>"00000001",
  24138=>"11111110",
  24139=>"00000010",
  24140=>"11111100",
  24141=>"11111101",
  24142=>"00000000",
  24143=>"00000010",
  24144=>"11111100",
  24145=>"11111111",
  24146=>"00000010",
  24147=>"00000000",
  24148=>"11111101",
  24149=>"11111101",
  24150=>"00000001",
  24151=>"11111101",
  24152=>"11111110",
  24153=>"00000011",
  24154=>"00000001",
  24155=>"00000001",
  24156=>"11111110",
  24157=>"00000000",
  24158=>"00000010",
  24159=>"00000010",
  24160=>"00000010",
  24161=>"11111101",
  24162=>"11111110",
  24163=>"00000001",
  24164=>"11111110",
  24165=>"11111111",
  24166=>"00000000",
  24167=>"00000010",
  24168=>"11111100",
  24169=>"11111101",
  24170=>"00000001",
  24171=>"11111101",
  24172=>"11111110",
  24173=>"00000000",
  24174=>"00000010",
  24175=>"11111110",
  24176=>"00000101",
  24177=>"00000000",
  24178=>"00000010",
  24179=>"00000010",
  24180=>"00000001",
  24181=>"00000010",
  24182=>"11111110",
  24183=>"11111101",
  24184=>"11111111",
  24185=>"11111100",
  24186=>"00000011",
  24187=>"00000010",
  24188=>"00000010",
  24189=>"00000011",
  24190=>"11111111",
  24191=>"00000001",
  24192=>"11111101",
  24193=>"00000001",
  24194=>"00000000",
  24195=>"11111111",
  24196=>"00000100",
  24197=>"11111110",
  24198=>"11111110",
  24199=>"00000011",
  24200=>"11111101",
  24201=>"11111110",
  24202=>"00000011",
  24203=>"11111111",
  24204=>"00000010",
  24205=>"00000001",
  24206=>"00000010",
  24207=>"00000001",
  24208=>"00000000",
  24209=>"00000000",
  24210=>"00000001",
  24211=>"11111110",
  24212=>"11111101",
  24213=>"00000001",
  24214=>"00000000",
  24215=>"11111111",
  24216=>"00000011",
  24217=>"00000001",
  24218=>"11111110",
  24219=>"00000011",
  24220=>"11111110",
  24221=>"00000000",
  24222=>"11111111",
  24223=>"00000000",
  24224=>"11111110",
  24225=>"00000001",
  24226=>"00000101",
  24227=>"11111111",
  24228=>"11111110",
  24229=>"11111110",
  24230=>"11111101",
  24231=>"00000001",
  24232=>"00000001",
  24233=>"11111101",
  24234=>"00000001",
  24235=>"11111111",
  24236=>"00000001",
  24237=>"00000000",
  24238=>"11111100",
  24239=>"11111111",
  24240=>"11111110",
  24241=>"00000010",
  24242=>"00000010",
  24243=>"11111110",
  24244=>"00000001",
  24245=>"11111101",
  24246=>"00000001",
  24247=>"00000000",
  24248=>"00000000",
  24249=>"00000000",
  24250=>"11111110",
  24251=>"00000011",
  24252=>"11111111",
  24253=>"00000000",
  24254=>"11111110",
  24255=>"11111111",
  24256=>"00000011",
  24257=>"11111110",
  24258=>"00000000",
  24259=>"00000011",
  24260=>"00000001",
  24261=>"00000001",
  24262=>"11111110",
  24263=>"11111110",
  24264=>"00000010",
  24265=>"00000100",
  24266=>"00000001",
  24267=>"00000010",
  24268=>"11111111",
  24269=>"00000010",
  24270=>"11111111",
  24271=>"00000010",
  24272=>"00000000",
  24273=>"11111100",
  24274=>"00000001",
  24275=>"11111101",
  24276=>"11111110",
  24277=>"00000000",
  24278=>"00000000",
  24279=>"00000001",
  24280=>"11111110",
  24281=>"00000010",
  24282=>"00000010",
  24283=>"11111111",
  24284=>"00000000",
  24285=>"11111110",
  24286=>"00000011",
  24287=>"11111100",
  24288=>"11111111",
  24289=>"00000000",
  24290=>"00000010",
  24291=>"11111101",
  24292=>"11111110",
  24293=>"00000101",
  24294=>"11111111",
  24295=>"11111110",
  24296=>"00000010",
  24297=>"11111110",
  24298=>"11111101",
  24299=>"11111111",
  24300=>"00000010",
  24301=>"00000000",
  24302=>"00000011",
  24303=>"11111110",
  24304=>"11111111",
  24305=>"00000001",
  24306=>"00000000",
  24307=>"00000010",
  24308=>"11111110",
  24309=>"11111101",
  24310=>"00000001",
  24311=>"00000000",
  24312=>"00000010",
  24313=>"00000000",
  24314=>"00000001",
  24315=>"11111111",
  24316=>"00000000",
  24317=>"00000011",
  24318=>"11111111",
  24319=>"11111101",
  24320=>"11111101",
  24321=>"11111110",
  24322=>"11111100",
  24323=>"00000000",
  24324=>"11111111",
  24325=>"00000000",
  24326=>"00000010",
  24327=>"00000010",
  24328=>"11111111",
  24329=>"00000001",
  24330=>"11111110",
  24331=>"11111111",
  24332=>"11111110",
  24333=>"11111110",
  24334=>"00000100",
  24335=>"00000010",
  24336=>"11111101",
  24337=>"11111111",
  24338=>"00000001",
  24339=>"11111110",
  24340=>"11111111",
  24341=>"00000000",
  24342=>"00000000",
  24343=>"00000000",
  24344=>"00000000",
  24345=>"11111111",
  24346=>"00000100",
  24347=>"00000001",
  24348=>"11111101",
  24349=>"11111110",
  24350=>"00000001",
  24351=>"11111101",
  24352=>"11111111",
  24353=>"00000100",
  24354=>"00000010",
  24355=>"00000000",
  24356=>"00000000",
  24357=>"11111111",
  24358=>"00000000",
  24359=>"11111101",
  24360=>"11111101",
  24361=>"00000010",
  24362=>"00000000",
  24363=>"11111111",
  24364=>"11111110",
  24365=>"11111111",
  24366=>"11111110",
  24367=>"11111110",
  24368=>"00000010",
  24369=>"11111110",
  24370=>"11111101",
  24371=>"11111110",
  24372=>"00000001",
  24373=>"00000101",
  24374=>"00000001",
  24375=>"00000010",
  24376=>"11111111",
  24377=>"00000000",
  24378=>"00000000",
  24379=>"11111111",
  24380=>"11111100",
  24381=>"11111111",
  24382=>"00000001",
  24383=>"00000000",
  24384=>"11111111",
  24385=>"11111110",
  24386=>"11111110",
  24387=>"00000001",
  24388=>"00000000",
  24389=>"00000010",
  24390=>"00000011",
  24391=>"00000000",
  24392=>"00000001",
  24393=>"00000000",
  24394=>"11111101",
  24395=>"00000001",
  24396=>"00000011",
  24397=>"11111111",
  24398=>"00000001",
  24399=>"00000010",
  24400=>"00000001",
  24401=>"11111101",
  24402=>"00000010",
  24403=>"00000000",
  24404=>"11111101",
  24405=>"00000001",
  24406=>"11111111",
  24407=>"11111111",
  24408=>"11111111",
  24409=>"00000100",
  24410=>"00000010",
  24411=>"11111110",
  24412=>"11111110",
  24413=>"00000000",
  24414=>"00000101",
  24415=>"00000000",
  24416=>"00000011",
  24417=>"11111110",
  24418=>"00000001",
  24419=>"11111110",
  24420=>"11111101",
  24421=>"11111111",
  24422=>"00000101",
  24423=>"00000010",
  24424=>"11111100",
  24425=>"00000111",
  24426=>"11111110",
  24427=>"00000010",
  24428=>"11111110",
  24429=>"11111110",
  24430=>"00000001",
  24431=>"11111100",
  24432=>"00000000",
  24433=>"00000001",
  24434=>"11111111",
  24435=>"00000010",
  24436=>"11111111",
  24437=>"00000010",
  24438=>"11111110",
  24439=>"00000010",
  24440=>"00000000",
  24441=>"11111110",
  24442=>"11111101",
  24443=>"11111101",
  24444=>"00000001",
  24445=>"11111100",
  24446=>"00000000",
  24447=>"11111111",
  24448=>"11111110",
  24449=>"11111110",
  24450=>"00000001",
  24451=>"11111110",
  24452=>"00000001",
  24453=>"00000001",
  24454=>"00000110",
  24455=>"00000010",
  24456=>"00000000",
  24457=>"11111110",
  24458=>"00000001",
  24459=>"11111101",
  24460=>"00000011",
  24461=>"11111111",
  24462=>"11111101",
  24463=>"11111101",
  24464=>"11111110",
  24465=>"11111111",
  24466=>"00000000",
  24467=>"00000000",
  24468=>"00000000",
  24469=>"00000010",
  24470=>"11111110",
  24471=>"00000010",
  24472=>"00000101",
  24473=>"11111110",
  24474=>"00000011",
  24475=>"00000000",
  24476=>"11111111",
  24477=>"00000001",
  24478=>"11111111",
  24479=>"00000000",
  24480=>"00000011",
  24481=>"00000100",
  24482=>"00000001",
  24483=>"00000001",
  24484=>"00000000",
  24485=>"00000000",
  24486=>"00000000",
  24487=>"11111111",
  24488=>"11111110",
  24489=>"00000001",
  24490=>"11111111",
  24491=>"00000010",
  24492=>"00000010",
  24493=>"11111111",
  24494=>"00000011",
  24495=>"11111101",
  24496=>"11111101",
  24497=>"00000001",
  24498=>"00000000",
  24499=>"11111101",
  24500=>"00000000",
  24501=>"00000010",
  24502=>"11111110",
  24503=>"00000000",
  24504=>"11111101",
  24505=>"11111111",
  24506=>"11111110",
  24507=>"00000000",
  24508=>"00000100",
  24509=>"11111110",
  24510=>"00000010",
  24511=>"00000010",
  24512=>"11111110",
  24513=>"00000100",
  24514=>"00000010",
  24515=>"11111110",
  24516=>"00000000",
  24517=>"11111111",
  24518=>"11111111",
  24519=>"00000000",
  24520=>"00000011",
  24521=>"00000011",
  24522=>"11111110",
  24523=>"00000100",
  24524=>"11111110",
  24525=>"00000000",
  24526=>"00000001",
  24527=>"11111111",
  24528=>"00000010",
  24529=>"11111110",
  24530=>"11111111",
  24531=>"00000000",
  24532=>"11111101",
  24533=>"00000010",
  24534=>"11111101",
  24535=>"11111111",
  24536=>"11111110",
  24537=>"11111110",
  24538=>"00000000",
  24539=>"11111111",
  24540=>"00000000",
  24541=>"11111111",
  24542=>"11111101",
  24543=>"11111100",
  24544=>"11111110",
  24545=>"00000011",
  24546=>"11111101",
  24547=>"00000000",
  24548=>"11111111",
  24549=>"11111111",
  24550=>"00000100",
  24551=>"11111100",
  24552=>"11111111",
  24553=>"11111110",
  24554=>"00000001",
  24555=>"00000011",
  24556=>"00000000",
  24557=>"00000000",
  24558=>"11111101",
  24559=>"00000000",
  24560=>"11111100",
  24561=>"00000001",
  24562=>"00000010",
  24563=>"11111101",
  24564=>"00000011",
  24565=>"00000011",
  24566=>"00000000",
  24567=>"00000010",
  24568=>"11111101",
  24569=>"11111101",
  24570=>"00000100",
  24571=>"00000010",
  24572=>"00000000",
  24573=>"11111101",
  24574=>"00000001",
  24575=>"00000001",
  24576=>"00000011",
  24577=>"00000111",
  24578=>"11111111",
  24579=>"11111110",
  24580=>"00000000",
  24581=>"00000000",
  24582=>"11111110",
  24583=>"00000111",
  24584=>"00000010",
  24585=>"00000011",
  24586=>"00000001",
  24587=>"11111101",
  24588=>"11111111",
  24589=>"00000010",
  24590=>"00000010",
  24591=>"00000000",
  24592=>"00000000",
  24593=>"00000001",
  24594=>"00000010",
  24595=>"00000000",
  24596=>"00000010",
  24597=>"11111110",
  24598=>"11111101",
  24599=>"00000000",
  24600=>"00000001",
  24601=>"11111110",
  24602=>"11111111",
  24603=>"11111110",
  24604=>"11111101",
  24605=>"11111110",
  24606=>"00000110",
  24607=>"11111101",
  24608=>"11111110",
  24609=>"11111110",
  24610=>"11111101",
  24611=>"00000010",
  24612=>"00000010",
  24613=>"00000000",
  24614=>"00000001",
  24615=>"11111111",
  24616=>"11111111",
  24617=>"00000000",
  24618=>"00000011",
  24619=>"00000011",
  24620=>"11111111",
  24621=>"11111101",
  24622=>"00000000",
  24623=>"00000011",
  24624=>"00000000",
  24625=>"11111111",
  24626=>"11111111",
  24627=>"11111100",
  24628=>"00000000",
  24629=>"11111111",
  24630=>"00000001",
  24631=>"00000011",
  24632=>"00000000",
  24633=>"11111110",
  24634=>"11111110",
  24635=>"11111111",
  24636=>"00000000",
  24637=>"11111101",
  24638=>"00000000",
  24639=>"00000011",
  24640=>"11111101",
  24641=>"00000000",
  24642=>"00000010",
  24643=>"00000010",
  24644=>"11111101",
  24645=>"00000001",
  24646=>"00000000",
  24647=>"00000001",
  24648=>"11111100",
  24649=>"00000000",
  24650=>"00000000",
  24651=>"00000000",
  24652=>"00000001",
  24653=>"00000100",
  24654=>"00000000",
  24655=>"11111111",
  24656=>"11111111",
  24657=>"11111111",
  24658=>"11111111",
  24659=>"00000010",
  24660=>"00000001",
  24661=>"00000010",
  24662=>"00000010",
  24663=>"11111110",
  24664=>"11111111",
  24665=>"00000001",
  24666=>"00000001",
  24667=>"00000010",
  24668=>"00000001",
  24669=>"00000100",
  24670=>"00000001",
  24671=>"11111110",
  24672=>"00000001",
  24673=>"00000000",
  24674=>"11111110",
  24675=>"00000001",
  24676=>"00000011",
  24677=>"11111111",
  24678=>"11111110",
  24679=>"11111101",
  24680=>"11111110",
  24681=>"11111111",
  24682=>"11111111",
  24683=>"00000001",
  24684=>"00000000",
  24685=>"00000000",
  24686=>"11111110",
  24687=>"00000000",
  24688=>"11111101",
  24689=>"11111111",
  24690=>"00000000",
  24691=>"00000011",
  24692=>"11111110",
  24693=>"11111101",
  24694=>"11111101",
  24695=>"00000000",
  24696=>"11111110",
  24697=>"00000000",
  24698=>"11111110",
  24699=>"11111101",
  24700=>"11111111",
  24701=>"11111100",
  24702=>"11111111",
  24703=>"00000001",
  24704=>"00000000",
  24705=>"00000001",
  24706=>"00000001",
  24707=>"00000010",
  24708=>"11111110",
  24709=>"00000001",
  24710=>"11111111",
  24711=>"11111111",
  24712=>"00000000",
  24713=>"00000001",
  24714=>"11111111",
  24715=>"00000001",
  24716=>"00000011",
  24717=>"00000001",
  24718=>"00000000",
  24719=>"00000011",
  24720=>"00000011",
  24721=>"00000010",
  24722=>"00000001",
  24723=>"11111111",
  24724=>"11111101",
  24725=>"00000100",
  24726=>"00000010",
  24727=>"11111111",
  24728=>"11111111",
  24729=>"11111111",
  24730=>"00000001",
  24731=>"00000011",
  24732=>"00000000",
  24733=>"11111100",
  24734=>"00000000",
  24735=>"00000100",
  24736=>"00000011",
  24737=>"11111110",
  24738=>"11111111",
  24739=>"00000100",
  24740=>"00000011",
  24741=>"00000001",
  24742=>"00000001",
  24743=>"11111110",
  24744=>"00000000",
  24745=>"00000001",
  24746=>"00000001",
  24747=>"11111110",
  24748=>"11111100",
  24749=>"11111110",
  24750=>"11111100",
  24751=>"11111111",
  24752=>"11111101",
  24753=>"00000010",
  24754=>"00000001",
  24755=>"11111111",
  24756=>"00000011",
  24757=>"00000001",
  24758=>"00000101",
  24759=>"11111100",
  24760=>"00000010",
  24761=>"00000010",
  24762=>"00000001",
  24763=>"00000000",
  24764=>"11111111",
  24765=>"11111111",
  24766=>"11111111",
  24767=>"11111111",
  24768=>"00000001",
  24769=>"11111111",
  24770=>"11111101",
  24771=>"00000010",
  24772=>"11111111",
  24773=>"11111110",
  24774=>"00000101",
  24775=>"00000010",
  24776=>"11111101",
  24777=>"00000011",
  24778=>"11111100",
  24779=>"00000000",
  24780=>"11111101",
  24781=>"11111100",
  24782=>"00000001",
  24783=>"11111111",
  24784=>"00000010",
  24785=>"11111101",
  24786=>"00000000",
  24787=>"00000010",
  24788=>"00000001",
  24789=>"11111110",
  24790=>"00000011",
  24791=>"00000010",
  24792=>"00000011",
  24793=>"00000000",
  24794=>"11111110",
  24795=>"11111110",
  24796=>"00000010",
  24797=>"11111111",
  24798=>"11111111",
  24799=>"11111111",
  24800=>"11111110",
  24801=>"00000000",
  24802=>"11111110",
  24803=>"11111111",
  24804=>"00000101",
  24805=>"00000100",
  24806=>"11111110",
  24807=>"11111101",
  24808=>"00000010",
  24809=>"11111110",
  24810=>"00000001",
  24811=>"00000001",
  24812=>"11111111",
  24813=>"11111110",
  24814=>"00000110",
  24815=>"11111111",
  24816=>"11111101",
  24817=>"00000010",
  24818=>"00000101",
  24819=>"11111110",
  24820=>"00001000",
  24821=>"00000000",
  24822=>"00000100",
  24823=>"00000010",
  24824=>"11111110",
  24825=>"11111111",
  24826=>"00000010",
  24827=>"11111101",
  24828=>"00000010",
  24829=>"11111110",
  24830=>"00000000",
  24831=>"00000001",
  24832=>"00000001",
  24833=>"00000001",
  24834=>"11111110",
  24835=>"00000001",
  24836=>"00000001",
  24837=>"11111110",
  24838=>"00000101",
  24839=>"00000000",
  24840=>"11111110",
  24841=>"11111111",
  24842=>"11111101",
  24843=>"00000001",
  24844=>"11111110",
  24845=>"11111110",
  24846=>"11111100",
  24847=>"00000000",
  24848=>"00000001",
  24849=>"00000011",
  24850=>"00000000",
  24851=>"00000010",
  24852=>"00000001",
  24853=>"00000010",
  24854=>"11111111",
  24855=>"00000011",
  24856=>"00000010",
  24857=>"11111111",
  24858=>"00000001",
  24859=>"00000000",
  24860=>"00000001",
  24861=>"11111111",
  24862=>"11111111",
  24863=>"00000001",
  24864=>"11111101",
  24865=>"11111111",
  24866=>"11111101",
  24867=>"00000001",
  24868=>"11111111",
  24869=>"11111110",
  24870=>"11111101",
  24871=>"11111100",
  24872=>"11111101",
  24873=>"11111101",
  24874=>"00000011",
  24875=>"11111111",
  24876=>"11111110",
  24877=>"00000011",
  24878=>"11111110",
  24879=>"00000100",
  24880=>"00000010",
  24881=>"11111110",
  24882=>"00000000",
  24883=>"00000000",
  24884=>"00000101",
  24885=>"11111101",
  24886=>"11111111",
  24887=>"00000010",
  24888=>"11111111",
  24889=>"00000010",
  24890=>"00000000",
  24891=>"11111111",
  24892=>"11111111",
  24893=>"00000101",
  24894=>"00000110",
  24895=>"11111111",
  24896=>"11111110",
  24897=>"11111110",
  24898=>"00000011",
  24899=>"00000011",
  24900=>"11111110",
  24901=>"11111100",
  24902=>"00000001",
  24903=>"00000001",
  24904=>"11111110",
  24905=>"00000000",
  24906=>"11111110",
  24907=>"00000000",
  24908=>"11111110",
  24909=>"00000000",
  24910=>"00000001",
  24911=>"11111101",
  24912=>"00000001",
  24913=>"11111110",
  24914=>"00000010",
  24915=>"00000000",
  24916=>"11111110",
  24917=>"00000000",
  24918=>"11111111",
  24919=>"00000001",
  24920=>"00000001",
  24921=>"00000100",
  24922=>"00000101",
  24923=>"00000110",
  24924=>"00000011",
  24925=>"00000010",
  24926=>"11111110",
  24927=>"00000011",
  24928=>"00000101",
  24929=>"11111111",
  24930=>"00000100",
  24931=>"11111101",
  24932=>"11111110",
  24933=>"00000001",
  24934=>"00000010",
  24935=>"11111111",
  24936=>"11111101",
  24937=>"11111100",
  24938=>"00000010",
  24939=>"11111111",
  24940=>"00000001",
  24941=>"11111111",
  24942=>"11111111",
  24943=>"11111111",
  24944=>"00000001",
  24945=>"00000100",
  24946=>"00000101",
  24947=>"00000010",
  24948=>"00000001",
  24949=>"11111111",
  24950=>"11111111",
  24951=>"11111110",
  24952=>"11111110",
  24953=>"11111101",
  24954=>"11111111",
  24955=>"11111110",
  24956=>"11111111",
  24957=>"00000001",
  24958=>"11111110",
  24959=>"11111100",
  24960=>"00000001",
  24961=>"00000110",
  24962=>"11111111",
  24963=>"11111110",
  24964=>"00000010",
  24965=>"11111101",
  24966=>"00000001",
  24967=>"00000010",
  24968=>"11111110",
  24969=>"00000000",
  24970=>"00000001",
  24971=>"00000010",
  24972=>"00000011",
  24973=>"00000001",
  24974=>"11111110",
  24975=>"00000001",
  24976=>"11111110",
  24977=>"11111110",
  24978=>"11111101",
  24979=>"00000100",
  24980=>"00000001",
  24981=>"00000001",
  24982=>"11111110",
  24983=>"11111110",
  24984=>"00000100",
  24985=>"11111111",
  24986=>"11111110",
  24987=>"11111011",
  24988=>"00000010",
  24989=>"00000001",
  24990=>"11111110",
  24991=>"00000010",
  24992=>"11111111",
  24993=>"00000001",
  24994=>"00000010",
  24995=>"00000111",
  24996=>"11111111",
  24997=>"11111111",
  24998=>"11111111",
  24999=>"00000011",
  25000=>"11111100",
  25001=>"11111110",
  25002=>"00000011",
  25003=>"11111110",
  25004=>"00000000",
  25005=>"11111101",
  25006=>"00000010",
  25007=>"11111101",
  25008=>"00000000",
  25009=>"00000010",
  25010=>"00000110",
  25011=>"00000000",
  25012=>"00000000",
  25013=>"11111101",
  25014=>"00000000",
  25015=>"11111111",
  25016=>"11111111",
  25017=>"00000101",
  25018=>"11111111",
  25019=>"00000010",
  25020=>"11111111",
  25021=>"00000001",
  25022=>"11111110",
  25023=>"00000010",
  25024=>"11111101",
  25025=>"11111111",
  25026=>"00000010",
  25027=>"00000001",
  25028=>"00000001",
  25029=>"11111110",
  25030=>"00000001",
  25031=>"11111100",
  25032=>"00000000",
  25033=>"00000000",
  25034=>"11111110",
  25035=>"11111111",
  25036=>"00000010",
  25037=>"00000010",
  25038=>"11111110",
  25039=>"11111110",
  25040=>"11111111",
  25041=>"11111111",
  25042=>"00000010",
  25043=>"00000001",
  25044=>"00000000",
  25045=>"11111101",
  25046=>"11111100",
  25047=>"11111101",
  25048=>"11111111",
  25049=>"00000001",
  25050=>"00000000",
  25051=>"00000001",
  25052=>"00000101",
  25053=>"11111101",
  25054=>"00000000",
  25055=>"11111110",
  25056=>"11111111",
  25057=>"11111110",
  25058=>"00000001",
  25059=>"00000000",
  25060=>"00000000",
  25061=>"11111111",
  25062=>"00000001",
  25063=>"00000000",
  25064=>"11111101",
  25065=>"00000001",
  25066=>"00000011",
  25067=>"00000001",
  25068=>"11111111",
  25069=>"11111100",
  25070=>"11111111",
  25071=>"00000000",
  25072=>"00000000",
  25073=>"00000100",
  25074=>"00000000",
  25075=>"00000110",
  25076=>"11111110",
  25077=>"00000000",
  25078=>"11111101",
  25079=>"11111110",
  25080=>"00000010",
  25081=>"00000000",
  25082=>"00000010",
  25083=>"00000010",
  25084=>"00000010",
  25085=>"00000000",
  25086=>"00000100",
  25087=>"11111110",
  25088=>"00000010",
  25089=>"00000010",
  25090=>"00000001",
  25091=>"00000011",
  25092=>"11111110",
  25093=>"11111110",
  25094=>"00000010",
  25095=>"11111111",
  25096=>"00000010",
  25097=>"00000000",
  25098=>"11111111",
  25099=>"11111110",
  25100=>"00000001",
  25101=>"00000001",
  25102=>"00000100",
  25103=>"11111110",
  25104=>"00000001",
  25105=>"11111111",
  25106=>"11111101",
  25107=>"00000001",
  25108=>"00000011",
  25109=>"11111110",
  25110=>"00000011",
  25111=>"00000000",
  25112=>"00000010",
  25113=>"00000001",
  25114=>"11111111",
  25115=>"00000001",
  25116=>"11111111",
  25117=>"11111111",
  25118=>"00000011",
  25119=>"11111110",
  25120=>"11111110",
  25121=>"11111111",
  25122=>"00000010",
  25123=>"00000001",
  25124=>"00000001",
  25125=>"00000001",
  25126=>"11111110",
  25127=>"11111111",
  25128=>"00000001",
  25129=>"00000000",
  25130=>"11111110",
  25131=>"00000100",
  25132=>"11111100",
  25133=>"11111110",
  25134=>"11111101",
  25135=>"00000001",
  25136=>"00000001",
  25137=>"11111110",
  25138=>"11111111",
  25139=>"11111110",
  25140=>"11111111",
  25141=>"11111101",
  25142=>"00000000",
  25143=>"11111110",
  25144=>"00000001",
  25145=>"11111110",
  25146=>"00000001",
  25147=>"11111111",
  25148=>"00000000",
  25149=>"00000011",
  25150=>"00000000",
  25151=>"00000101",
  25152=>"11111101",
  25153=>"11111101",
  25154=>"00000000",
  25155=>"00000000",
  25156=>"00000001",
  25157=>"00000011",
  25158=>"00000111",
  25159=>"00000010",
  25160=>"11111111",
  25161=>"11111111",
  25162=>"00000011",
  25163=>"00000000",
  25164=>"00000000",
  25165=>"00000110",
  25166=>"11111101",
  25167=>"11111101",
  25168=>"11111101",
  25169=>"00000000",
  25170=>"11111111",
  25171=>"00000000",
  25172=>"11111110",
  25173=>"11111101",
  25174=>"00000010",
  25175=>"11111110",
  25176=>"00000001",
  25177=>"00000000",
  25178=>"00000010",
  25179=>"11111101",
  25180=>"11111101",
  25181=>"11111101",
  25182=>"11111110",
  25183=>"11111101",
  25184=>"11111110",
  25185=>"00000001",
  25186=>"00000010",
  25187=>"00000011",
  25188=>"00000011",
  25189=>"00000001",
  25190=>"00000001",
  25191=>"11111110",
  25192=>"11111100",
  25193=>"00000001",
  25194=>"00000010",
  25195=>"00000001",
  25196=>"00000001",
  25197=>"00000001",
  25198=>"00000110",
  25199=>"00000100",
  25200=>"11111100",
  25201=>"11111111",
  25202=>"11111110",
  25203=>"00000000",
  25204=>"00000000",
  25205=>"11111110",
  25206=>"11111101",
  25207=>"00000100",
  25208=>"00000000",
  25209=>"00000001",
  25210=>"11111101",
  25211=>"00000001",
  25212=>"00000001",
  25213=>"11111111",
  25214=>"00000001",
  25215=>"00000001",
  25216=>"11111101",
  25217=>"11111111",
  25218=>"00000001",
  25219=>"00000100",
  25220=>"11111100",
  25221=>"11111111",
  25222=>"00000001",
  25223=>"11111100",
  25224=>"11111111",
  25225=>"00000000",
  25226=>"00000111",
  25227=>"00000011",
  25228=>"11111101",
  25229=>"00000010",
  25230=>"00000001",
  25231=>"11111110",
  25232=>"11111101",
  25233=>"11111100",
  25234=>"00000001",
  25235=>"00000000",
  25236=>"11111101",
  25237=>"00000011",
  25238=>"00000001",
  25239=>"00000000",
  25240=>"11111111",
  25241=>"00000001",
  25242=>"11111110",
  25243=>"11111110",
  25244=>"11111101",
  25245=>"00000111",
  25246=>"00000010",
  25247=>"11111111",
  25248=>"00000000",
  25249=>"00000001",
  25250=>"00000011",
  25251=>"00000001",
  25252=>"11111101",
  25253=>"00000001",
  25254=>"00000000",
  25255=>"11111110",
  25256=>"00000000",
  25257=>"11111110",
  25258=>"11111110",
  25259=>"00000001",
  25260=>"11111101",
  25261=>"00000001",
  25262=>"00000011",
  25263=>"11111101",
  25264=>"00000011",
  25265=>"00000001",
  25266=>"00000010",
  25267=>"11111100",
  25268=>"11111111",
  25269=>"00000000",
  25270=>"00000001",
  25271=>"00000001",
  25272=>"11111110",
  25273=>"11111101",
  25274=>"00000001",
  25275=>"11111101",
  25276=>"11111100",
  25277=>"00000011",
  25278=>"11111101",
  25279=>"00000000",
  25280=>"11111111",
  25281=>"00000010",
  25282=>"00000010",
  25283=>"00000000",
  25284=>"11111111",
  25285=>"11111110",
  25286=>"00000011",
  25287=>"11111111",
  25288=>"00000000",
  25289=>"00000110",
  25290=>"11111100",
  25291=>"11111111",
  25292=>"00000001",
  25293=>"00000011",
  25294=>"00000010",
  25295=>"00000000",
  25296=>"00000000",
  25297=>"00000100",
  25298=>"00000011",
  25299=>"00000010",
  25300=>"00000010",
  25301=>"00000000",
  25302=>"00000001",
  25303=>"11111110",
  25304=>"00000000",
  25305=>"00000000",
  25306=>"11111110",
  25307=>"00000010",
  25308=>"00000000",
  25309=>"00000000",
  25310=>"00000001",
  25311=>"00000011",
  25312=>"00000001",
  25313=>"00000010",
  25314=>"11111111",
  25315=>"00000101",
  25316=>"00000101",
  25317=>"11111110",
  25318=>"11111101",
  25319=>"11111111",
  25320=>"11111111",
  25321=>"11111110",
  25322=>"00000011",
  25323=>"11111110",
  25324=>"11111110",
  25325=>"00000010",
  25326=>"00000011",
  25327=>"00000000",
  25328=>"11111110",
  25329=>"00000000",
  25330=>"00000001",
  25331=>"11111110",
  25332=>"11111100",
  25333=>"11111111",
  25334=>"11111111",
  25335=>"00000000",
  25336=>"00000001",
  25337=>"11111111",
  25338=>"11111110",
  25339=>"11111100",
  25340=>"11111101",
  25341=>"11111011",
  25342=>"00000011",
  25343=>"11111111",
  25344=>"00000100",
  25345=>"11111110",
  25346=>"11111111",
  25347=>"00000001",
  25348=>"00000100",
  25349=>"00000010",
  25350=>"00000010",
  25351=>"00000110",
  25352=>"00000101",
  25353=>"00000100",
  25354=>"11111110",
  25355=>"11111110",
  25356=>"00000000",
  25357=>"00000101",
  25358=>"00000011",
  25359=>"00000001",
  25360=>"00000001",
  25361=>"11111111",
  25362=>"00000100",
  25363=>"00000000",
  25364=>"00000010",
  25365=>"11111110",
  25366=>"11111100",
  25367=>"00000000",
  25368=>"00000011",
  25369=>"11111110",
  25370=>"00000000",
  25371=>"00000010",
  25372=>"11111110",
  25373=>"11111111",
  25374=>"11111110",
  25375=>"11111011",
  25376=>"00000010",
  25377=>"00000100",
  25378=>"00000010",
  25379=>"00000000",
  25380=>"00000000",
  25381=>"00000000",
  25382=>"00000000",
  25383=>"11111110",
  25384=>"11111111",
  25385=>"00000001",
  25386=>"11111111",
  25387=>"11111011",
  25388=>"00000001",
  25389=>"11111101",
  25390=>"00000011",
  25391=>"11111110",
  25392=>"00000000",
  25393=>"00000000",
  25394=>"00000000",
  25395=>"00000011",
  25396=>"00000010",
  25397=>"00000000",
  25398=>"00000000",
  25399=>"00000001",
  25400=>"00000010",
  25401=>"00000010",
  25402=>"00000000",
  25403=>"00000010",
  25404=>"11111110",
  25405=>"00000000",
  25406=>"11111101",
  25407=>"11111110",
  25408=>"11111111",
  25409=>"00000010",
  25410=>"00000001",
  25411=>"00000000",
  25412=>"11111110",
  25413=>"11111111",
  25414=>"11111101",
  25415=>"00000010",
  25416=>"11111110",
  25417=>"11111111",
  25418=>"00000001",
  25419=>"00000000",
  25420=>"00000000",
  25421=>"00000000",
  25422=>"00000010",
  25423=>"00000010",
  25424=>"11111111",
  25425=>"11111110",
  25426=>"00000110",
  25427=>"11111110",
  25428=>"00000011",
  25429=>"11111110",
  25430=>"00000001",
  25431=>"00000001",
  25432=>"11111110",
  25433=>"00000011",
  25434=>"00000000",
  25435=>"11111111",
  25436=>"00000000",
  25437=>"11111111",
  25438=>"00000010",
  25439=>"00000011",
  25440=>"11111110",
  25441=>"11111111",
  25442=>"00000011",
  25443=>"11111111",
  25444=>"00000010",
  25445=>"00000001",
  25446=>"11111110",
  25447=>"00000110",
  25448=>"11111100",
  25449=>"11111100",
  25450=>"00000000",
  25451=>"00000000",
  25452=>"00000001",
  25453=>"11111111",
  25454=>"00000001",
  25455=>"00000011",
  25456=>"00000010",
  25457=>"00000001",
  25458=>"00000011",
  25459=>"00000001",
  25460=>"00000011",
  25461=>"00000001",
  25462=>"00000110",
  25463=>"00000100",
  25464=>"00000000",
  25465=>"11111111",
  25466=>"00000000",
  25467=>"00000011",
  25468=>"00000001",
  25469=>"11111011",
  25470=>"00000011",
  25471=>"00000101",
  25472=>"11111111",
  25473=>"00000000",
  25474=>"11111111",
  25475=>"11111100",
  25476=>"11111100",
  25477=>"00000001",
  25478=>"11111110",
  25479=>"11111110",
  25480=>"00000001",
  25481=>"00000001",
  25482=>"00000001",
  25483=>"11111111",
  25484=>"11111110",
  25485=>"11111111",
  25486=>"11111101",
  25487=>"00000001",
  25488=>"11111100",
  25489=>"11111110",
  25490=>"11111110",
  25491=>"00000011",
  25492=>"00000010",
  25493=>"11111100",
  25494=>"00000010",
  25495=>"11111101",
  25496=>"11111111",
  25497=>"11111101",
  25498=>"11111100",
  25499=>"11111110",
  25500=>"00000000",
  25501=>"00000010",
  25502=>"11111110",
  25503=>"00000001",
  25504=>"00000001",
  25505=>"00000000",
  25506=>"00000010",
  25507=>"11111111",
  25508=>"00000000",
  25509=>"11111101",
  25510=>"00000000",
  25511=>"00000010",
  25512=>"00000010",
  25513=>"00000000",
  25514=>"11111110",
  25515=>"00000011",
  25516=>"00000001",
  25517=>"11111111",
  25518=>"00000001",
  25519=>"00000011",
  25520=>"00000001",
  25521=>"00000010",
  25522=>"00000001",
  25523=>"11111101",
  25524=>"00000010",
  25525=>"00000001",
  25526=>"11111101",
  25527=>"11111111",
  25528=>"00000110",
  25529=>"11111111",
  25530=>"00000001",
  25531=>"11111110",
  25532=>"11111101",
  25533=>"00000100",
  25534=>"00000001",
  25535=>"00000010",
  25536=>"00000000",
  25537=>"11111111",
  25538=>"11111101",
  25539=>"00000010",
  25540=>"00000011",
  25541=>"00000001",
  25542=>"00000010",
  25543=>"00000001",
  25544=>"11111110",
  25545=>"00000101",
  25546=>"11111111",
  25547=>"11111110",
  25548=>"11111101",
  25549=>"11111110",
  25550=>"11111101",
  25551=>"00000001",
  25552=>"11111110",
  25553=>"00000001",
  25554=>"00000011",
  25555=>"11111100",
  25556=>"11111111",
  25557=>"00000011",
  25558=>"00000000",
  25559=>"11111111",
  25560=>"11111110",
  25561=>"11111101",
  25562=>"00000001",
  25563=>"00000000",
  25564=>"00000110",
  25565=>"11111110",
  25566=>"11111111",
  25567=>"00000001",
  25568=>"00000100",
  25569=>"11111111",
  25570=>"00000000",
  25571=>"00000001",
  25572=>"11111110",
  25573=>"11111100",
  25574=>"11111110",
  25575=>"11111110",
  25576=>"00000011",
  25577=>"00000010",
  25578=>"11111110",
  25579=>"11111101",
  25580=>"00000011",
  25581=>"11111111",
  25582=>"00000001",
  25583=>"11111101",
  25584=>"11111101",
  25585=>"00000000",
  25586=>"11111100",
  25587=>"00000010",
  25588=>"00000000",
  25589=>"00000000",
  25590=>"11111110",
  25591=>"00000000",
  25592=>"00000010",
  25593=>"00000100",
  25594=>"11111110",
  25595=>"11111111",
  25596=>"11111110",
  25597=>"00000000",
  25598=>"11111100",
  25599=>"11111101",
  25600=>"00000001",
  25601=>"11111111",
  25602=>"00000001",
  25603=>"00000011",
  25604=>"00000000",
  25605=>"11111111",
  25606=>"11111111",
  25607=>"11111111",
  25608=>"00000000",
  25609=>"00000000",
  25610=>"00000000",
  25611=>"00000001",
  25612=>"00000001",
  25613=>"11111111",
  25614=>"00000001",
  25615=>"11111111",
  25616=>"00000010",
  25617=>"00000010",
  25618=>"00000010",
  25619=>"11111110",
  25620=>"00000000",
  25621=>"11111110",
  25622=>"00000001",
  25623=>"00000001",
  25624=>"00000001",
  25625=>"00000001",
  25626=>"11111111",
  25627=>"00000001",
  25628=>"11111111",
  25629=>"11111111",
  25630=>"00000010",
  25631=>"11111110",
  25632=>"00000001",
  25633=>"00000000",
  25634=>"00000001",
  25635=>"11111110",
  25636=>"00000010",
  25637=>"11111111",
  25638=>"00000000",
  25639=>"00000000",
  25640=>"00000001",
  25641=>"00000001",
  25642=>"00000000",
  25643=>"00000000",
  25644=>"11111111",
  25645=>"11111101",
  25646=>"00000010",
  25647=>"00000001",
  25648=>"00000001",
  25649=>"00000001",
  25650=>"00000001",
  25651=>"00000000",
  25652=>"00000001",
  25653=>"00000000",
  25654=>"11111111",
  25655=>"00000010",
  25656=>"11111111",
  25657=>"00000000",
  25658=>"00000001",
  25659=>"00000000",
  25660=>"11111111",
  25661=>"00000001",
  25662=>"00000001",
  25663=>"11111110",
  25664=>"11111111",
  25665=>"00000000",
  25666=>"11111111",
  25667=>"11111111",
  25668=>"00000001",
  25669=>"00000001",
  25670=>"00000001",
  25671=>"00000000",
  25672=>"00000001",
  25673=>"00000010",
  25674=>"00000001",
  25675=>"00000001",
  25676=>"11111110",
  25677=>"00000000",
  25678=>"00000001",
  25679=>"00000010",
  25680=>"00000001",
  25681=>"00000000",
  25682=>"11111110",
  25683=>"00000000",
  25684=>"00000010",
  25685=>"00000000",
  25686=>"11111110",
  25687=>"11111111",
  25688=>"11111111",
  25689=>"00000000",
  25690=>"00000000",
  25691=>"00000000",
  25692=>"11111111",
  25693=>"11111110",
  25694=>"00000001",
  25695=>"00000000",
  25696=>"00000000",
  25697=>"11111111",
  25698=>"00000010",
  25699=>"11111111",
  25700=>"00000001",
  25701=>"00000000",
  25702=>"00000000",
  25703=>"00000000",
  25704=>"00000000",
  25705=>"00000000",
  25706=>"00000000",
  25707=>"00000000",
  25708=>"11111110",
  25709=>"11111111",
  25710=>"11111111",
  25711=>"00000001",
  25712=>"00000000",
  25713=>"00000010",
  25714=>"00000010",
  25715=>"00000000",
  25716=>"00000000",
  25717=>"11111110",
  25718=>"00000001",
  25719=>"00000000",
  25720=>"00000010",
  25721=>"00000000",
  25722=>"11111111",
  25723=>"00000000",
  25724=>"00000000",
  25725=>"00000011",
  25726=>"00000010",
  25727=>"00000000",
  25728=>"00000010",
  25729=>"00000001",
  25730=>"00000001",
  25731=>"00000001",
  25732=>"00000001",
  25733=>"11111110",
  25734=>"11111111",
  25735=>"11111110",
  25736=>"11111111",
  25737=>"00000010",
  25738=>"00000000",
  25739=>"00000001",
  25740=>"00000011",
  25741=>"11111111",
  25742=>"11111110",
  25743=>"00000000",
  25744=>"11111111",
  25745=>"11111111",
  25746=>"11111110",
  25747=>"00000001",
  25748=>"11111111",
  25749=>"00000000",
  25750=>"11111111",
  25751=>"11111111",
  25752=>"11111111",
  25753=>"00000000",
  25754=>"11111111",
  25755=>"00000001",
  25756=>"00000000",
  25757=>"11111111",
  25758=>"11111110",
  25759=>"00000001",
  25760=>"11111110",
  25761=>"00000001",
  25762=>"00000000",
  25763=>"00000001",
  25764=>"00000001",
  25765=>"00000001",
  25766=>"00000010",
  25767=>"11111111",
  25768=>"00000001",
  25769=>"00000000",
  25770=>"11111110",
  25771=>"00000001",
  25772=>"00000001",
  25773=>"00000001",
  25774=>"11111111",
  25775=>"11111110",
  25776=>"00000000",
  25777=>"11111111",
  25778=>"00000000",
  25779=>"00000010",
  25780=>"11111110",
  25781=>"11111101",
  25782=>"11111110",
  25783=>"11111111",
  25784=>"00000001",
  25785=>"11111111",
  25786=>"00000001",
  25787=>"00000000",
  25788=>"00000000",
  25789=>"00000010",
  25790=>"11111111",
  25791=>"00000001",
  25792=>"00000000",
  25793=>"00000000",
  25794=>"00000001",
  25795=>"00000000",
  25796=>"11111111",
  25797=>"00000000",
  25798=>"00000000",
  25799=>"11111110",
  25800=>"11111111",
  25801=>"00000001",
  25802=>"00000001",
  25803=>"11111101",
  25804=>"11111111",
  25805=>"11111111",
  25806=>"11111110",
  25807=>"00000001",
  25808=>"00000000",
  25809=>"00000010",
  25810=>"00000001",
  25811=>"00000000",
  25812=>"00000001",
  25813=>"00000000",
  25814=>"00000001",
  25815=>"11111111",
  25816=>"00000000",
  25817=>"00000001",
  25818=>"00000001",
  25819=>"00000011",
  25820=>"00000000",
  25821=>"00000010",
  25822=>"00000001",
  25823=>"11111110",
  25824=>"11111111",
  25825=>"00000000",
  25826=>"00000000",
  25827=>"00000001",
  25828=>"11111101",
  25829=>"11111110",
  25830=>"00000011",
  25831=>"11111110",
  25832=>"11111110",
  25833=>"00000001",
  25834=>"11111110",
  25835=>"11111111",
  25836=>"11111111",
  25837=>"11111110",
  25838=>"00000000",
  25839=>"00000001",
  25840=>"00000010",
  25841=>"11111110",
  25842=>"11111111",
  25843=>"00000000",
  25844=>"00000010",
  25845=>"11111101",
  25846=>"11111101",
  25847=>"11111110",
  25848=>"00000000",
  25849=>"00000010",
  25850=>"00000001",
  25851=>"11111111",
  25852=>"00000001",
  25853=>"00000001",
  25854=>"00000000",
  25855=>"11111110",
  25856=>"11111111",
  25857=>"00000001",
  25858=>"00000001",
  25859=>"11111110",
  25860=>"11111110",
  25861=>"00000000",
  25862=>"00000001",
  25863=>"11111111",
  25864=>"00000000",
  25865=>"00000001",
  25866=>"11111111",
  25867=>"00000001",
  25868=>"00000010",
  25869=>"00000010",
  25870=>"00000000",
  25871=>"00000001",
  25872=>"00000000",
  25873=>"00000001",
  25874=>"00000001",
  25875=>"00000000",
  25876=>"00000010",
  25877=>"00000000",
  25878=>"00000001",
  25879=>"00000000",
  25880=>"00000000",
  25881=>"00000001",
  25882=>"00000010",
  25883=>"11111110",
  25884=>"11111111",
  25885=>"00000010",
  25886=>"11111111",
  25887=>"00000000",
  25888=>"00000001",
  25889=>"11111110",
  25890=>"00000000",
  25891=>"00000001",
  25892=>"00000001",
  25893=>"11111111",
  25894=>"00000010",
  25895=>"00000010",
  25896=>"00000001",
  25897=>"11111111",
  25898=>"00000000",
  25899=>"00000001",
  25900=>"00000010",
  25901=>"00000011",
  25902=>"00000000",
  25903=>"00000001",
  25904=>"00000001",
  25905=>"00000001",
  25906=>"11111111",
  25907=>"00000000",
  25908=>"00000000",
  25909=>"00000010",
  25910=>"11111110",
  25911=>"00000011",
  25912=>"00000000",
  25913=>"00000000",
  25914=>"11111111",
  25915=>"00000001",
  25916=>"00000001",
  25917=>"00000000",
  25918=>"11111110",
  25919=>"11111111",
  25920=>"00000001",
  25921=>"00000001",
  25922=>"00000011",
  25923=>"00000001",
  25924=>"11111011",
  25925=>"00000010",
  25926=>"11111111",
  25927=>"00000001",
  25928=>"11111110",
  25929=>"00000001",
  25930=>"00000000",
  25931=>"11111110",
  25932=>"00000000",
  25933=>"00000000",
  25934=>"00000000",
  25935=>"11111111",
  25936=>"00000001",
  25937=>"00000001",
  25938=>"00000001",
  25939=>"11111111",
  25940=>"00000010",
  25941=>"00000010",
  25942=>"11111110",
  25943=>"11111110",
  25944=>"00000000",
  25945=>"00000000",
  25946=>"00000010",
  25947=>"11111110",
  25948=>"00000010",
  25949=>"11111111",
  25950=>"00000000",
  25951=>"00000000",
  25952=>"11111111",
  25953=>"11111111",
  25954=>"11111111",
  25955=>"11111110",
  25956=>"11111111",
  25957=>"00000000",
  25958=>"00000010",
  25959=>"11111111",
  25960=>"11111110",
  25961=>"00000000",
  25962=>"11111110",
  25963=>"00000001",
  25964=>"11111101",
  25965=>"00000001",
  25966=>"11111111",
  25967=>"00000001",
  25968=>"00000010",
  25969=>"00000010",
  25970=>"11111111",
  25971=>"00000001",
  25972=>"00000001",
  25973=>"11111110",
  25974=>"00000010",
  25975=>"11111111",
  25976=>"00000001",
  25977=>"00000010",
  25978=>"00000000",
  25979=>"11111111",
  25980=>"11111110",
  25981=>"00000000",
  25982=>"11111111",
  25983=>"11111111",
  25984=>"11111111",
  25985=>"00000001",
  25986=>"11111111",
  25987=>"00000000",
  25988=>"00000001",
  25989=>"11111111",
  25990=>"00000001",
  25991=>"11111110",
  25992=>"00000001",
  25993=>"00000010",
  25994=>"00000010",
  25995=>"00000010",
  25996=>"00000001",
  25997=>"00000010",
  25998=>"00000001",
  25999=>"00000001",
  26000=>"00000001",
  26001=>"00000001",
  26002=>"00000000",
  26003=>"00000000",
  26004=>"00000001",
  26005=>"00000000",
  26006=>"00000001",
  26007=>"00000001",
  26008=>"11111111",
  26009=>"11111111",
  26010=>"00000001",
  26011=>"11111111",
  26012=>"00000010",
  26013=>"11111110",
  26014=>"00000000",
  26015=>"11111111",
  26016=>"00000000",
  26017=>"00000001",
  26018=>"11111111",
  26019=>"11111111",
  26020=>"11111111",
  26021=>"11111110",
  26022=>"11111111",
  26023=>"00000001",
  26024=>"11111110",
  26025=>"11111111",
  26026=>"00000000",
  26027=>"00000000",
  26028=>"11111101",
  26029=>"11111110",
  26030=>"00000000",
  26031=>"00000001",
  26032=>"00000001",
  26033=>"11111110",
  26034=>"11111111",
  26035=>"00000001",
  26036=>"11111110",
  26037=>"00000010",
  26038=>"11111111",
  26039=>"00000001",
  26040=>"11111110",
  26041=>"00000010",
  26042=>"00000010",
  26043=>"11111101",
  26044=>"00000010",
  26045=>"11111111",
  26046=>"00000000",
  26047=>"11111110",
  26048=>"11111111",
  26049=>"00000001",
  26050=>"00000001",
  26051=>"11111110",
  26052=>"00000010",
  26053=>"00000010",
  26054=>"00000010",
  26055=>"00000010",
  26056=>"11111110",
  26057=>"00000000",
  26058=>"00000001",
  26059=>"11111111",
  26060=>"00000001",
  26061=>"11111111",
  26062=>"00000001",
  26063=>"11111111",
  26064=>"00000000",
  26065=>"11111111",
  26066=>"00000001",
  26067=>"00000010",
  26068=>"00000001",
  26069=>"00000001",
  26070=>"00000000",
  26071=>"11111110",
  26072=>"00000001",
  26073=>"00000000",
  26074=>"11111110",
  26075=>"00000001",
  26076=>"00000010",
  26077=>"11111111",
  26078=>"00000001",
  26079=>"11111110",
  26080=>"11111111",
  26081=>"00000000",
  26082=>"00000000",
  26083=>"00000010",
  26084=>"00000000",
  26085=>"11111110",
  26086=>"00000010",
  26087=>"00000001",
  26088=>"00000001",
  26089=>"00000001",
  26090=>"00000010",
  26091=>"11111111",
  26092=>"11111111",
  26093=>"00000001",
  26094=>"00000001",
  26095=>"00000010",
  26096=>"00000001",
  26097=>"00000001",
  26098=>"00000001",
  26099=>"00000011",
  26100=>"00000000",
  26101=>"11111111",
  26102=>"00000001",
  26103=>"00000000",
  26104=>"00000010",
  26105=>"11111110",
  26106=>"11111111",
  26107=>"00000000",
  26108=>"00000000",
  26109=>"11111111",
  26110=>"00000001",
  26111=>"11111111",
  26112=>"00000000",
  26113=>"00000000",
  26114=>"00000000",
  26115=>"11111110",
  26116=>"00000000",
  26117=>"11111111",
  26118=>"00000010",
  26119=>"00000000",
  26120=>"11111111",
  26121=>"00000010",
  26122=>"00000010",
  26123=>"00000000",
  26124=>"00000001",
  26125=>"00000001",
  26126=>"00000000",
  26127=>"00000000",
  26128=>"11111111",
  26129=>"11111111",
  26130=>"00000001",
  26131=>"00000010",
  26132=>"00000000",
  26133=>"00000000",
  26134=>"00000001",
  26135=>"11111111",
  26136=>"00000000",
  26137=>"00000001",
  26138=>"11111110",
  26139=>"00000000",
  26140=>"00000000",
  26141=>"11111110",
  26142=>"11111111",
  26143=>"11111111",
  26144=>"00000000",
  26145=>"11111111",
  26146=>"00000000",
  26147=>"00000010",
  26148=>"00000000",
  26149=>"00000000",
  26150=>"00000000",
  26151=>"00000001",
  26152=>"11111111",
  26153=>"00000000",
  26154=>"11111110",
  26155=>"00000010",
  26156=>"11111111",
  26157=>"00000001",
  26158=>"00000001",
  26159=>"00000001",
  26160=>"00000001",
  26161=>"11111110",
  26162=>"00000000",
  26163=>"11111111",
  26164=>"00000000",
  26165=>"00000010",
  26166=>"00000001",
  26167=>"00000001",
  26168=>"00000000",
  26169=>"11111101",
  26170=>"00000000",
  26171=>"11111111",
  26172=>"11111110",
  26173=>"00000000",
  26174=>"11111111",
  26175=>"11111111",
  26176=>"11111111",
  26177=>"00000001",
  26178=>"11111111",
  26179=>"00000001",
  26180=>"11111110",
  26181=>"00000001",
  26182=>"00000001",
  26183=>"00000000",
  26184=>"11111111",
  26185=>"00000000",
  26186=>"11111111",
  26187=>"00000001",
  26188=>"11111110",
  26189=>"00000001",
  26190=>"00000000",
  26191=>"11111111",
  26192=>"00000010",
  26193=>"00000000",
  26194=>"00000000",
  26195=>"11111111",
  26196=>"00000001",
  26197=>"00000000",
  26198=>"00000001",
  26199=>"11111110",
  26200=>"00000000",
  26201=>"11111111",
  26202=>"11111111",
  26203=>"00000000",
  26204=>"00000011",
  26205=>"11111111",
  26206=>"00000001",
  26207=>"11111111",
  26208=>"11111111",
  26209=>"11111111",
  26210=>"00000010",
  26211=>"11111111",
  26212=>"11111101",
  26213=>"11111111",
  26214=>"00000010",
  26215=>"00000000",
  26216=>"11111111",
  26217=>"11111111",
  26218=>"00000010",
  26219=>"00000000",
  26220=>"11111111",
  26221=>"11111111",
  26222=>"00000000",
  26223=>"00000010",
  26224=>"00000001",
  26225=>"11111111",
  26226=>"11111111",
  26227=>"11111111",
  26228=>"00000000",
  26229=>"00000001",
  26230=>"00000000",
  26231=>"00000001",
  26232=>"00000010",
  26233=>"00000000",
  26234=>"11111111",
  26235=>"00000001",
  26236=>"11111110",
  26237=>"00000011",
  26238=>"00000001",
  26239=>"11111110",
  26240=>"11111111",
  26241=>"00000010",
  26242=>"00000001",
  26243=>"11111110",
  26244=>"11111111",
  26245=>"00000000",
  26246=>"00000000",
  26247=>"11111110",
  26248=>"00000000",
  26249=>"11111111",
  26250=>"00000000",
  26251=>"00000000",
  26252=>"11111111",
  26253=>"11111111",
  26254=>"00000001",
  26255=>"11111111",
  26256=>"00000000",
  26257=>"11111111",
  26258=>"00000001",
  26259=>"00000000",
  26260=>"00000010",
  26261=>"11111111",
  26262=>"11111111",
  26263=>"00000011",
  26264=>"00000001",
  26265=>"00000010",
  26266=>"00000001",
  26267=>"00000000",
  26268=>"00000000",
  26269=>"00000010",
  26270=>"00000010",
  26271=>"00000001",
  26272=>"00000001",
  26273=>"00000000",
  26274=>"00000011",
  26275=>"00000001",
  26276=>"11111110",
  26277=>"11111111",
  26278=>"11111101",
  26279=>"00000001",
  26280=>"00000001",
  26281=>"00000000",
  26282=>"00000000",
  26283=>"00000001",
  26284=>"11111110",
  26285=>"11111110",
  26286=>"00000001",
  26287=>"11111111",
  26288=>"11111110",
  26289=>"11111111",
  26290=>"11111111",
  26291=>"11111101",
  26292=>"11111111",
  26293=>"00000001",
  26294=>"00000001",
  26295=>"00000001",
  26296=>"11111111",
  26297=>"00000001",
  26298=>"00000000",
  26299=>"00000001",
  26300=>"00000000",
  26301=>"00000000",
  26302=>"00000000",
  26303=>"11111111",
  26304=>"11111111",
  26305=>"00000000",
  26306=>"11111110",
  26307=>"11111110",
  26308=>"00000001",
  26309=>"11111111",
  26310=>"00000001",
  26311=>"00000001",
  26312=>"11111101",
  26313=>"11111111",
  26314=>"11111111",
  26315=>"11111111",
  26316=>"11111111",
  26317=>"00000001",
  26318=>"11111111",
  26319=>"00000000",
  26320=>"11111110",
  26321=>"00000001",
  26322=>"00000001",
  26323=>"00000000",
  26324=>"11111110",
  26325=>"11111111",
  26326=>"11111111",
  26327=>"11111111",
  26328=>"11111111",
  26329=>"11111111",
  26330=>"00000000",
  26331=>"00000001",
  26332=>"00000001",
  26333=>"00000010",
  26334=>"11111110",
  26335=>"00000001",
  26336=>"00000000",
  26337=>"11111110",
  26338=>"00000010",
  26339=>"00000001",
  26340=>"11111111",
  26341=>"00000001",
  26342=>"00000000",
  26343=>"00000000",
  26344=>"00000001",
  26345=>"11111111",
  26346=>"00000000",
  26347=>"11111111",
  26348=>"11111111",
  26349=>"00000001",
  26350=>"00000001",
  26351=>"00000000",
  26352=>"00000000",
  26353=>"11111111",
  26354=>"00000011",
  26355=>"00000000",
  26356=>"00000000",
  26357=>"00000001",
  26358=>"00000001",
  26359=>"00000001",
  26360=>"00000001",
  26361=>"11111110",
  26362=>"00000001",
  26363=>"11111111",
  26364=>"00000011",
  26365=>"00000010",
  26366=>"11111110",
  26367=>"00000000",
  26368=>"00000001",
  26369=>"00000010",
  26370=>"00000001",
  26371=>"11111111",
  26372=>"00000001",
  26373=>"11111110",
  26374=>"00000001",
  26375=>"00000000",
  26376=>"00000000",
  26377=>"11111110",
  26378=>"00000001",
  26379=>"00000000",
  26380=>"11111110",
  26381=>"11111111",
  26382=>"11111111",
  26383=>"00000000",
  26384=>"00000000",
  26385=>"11111111",
  26386=>"11111111",
  26387=>"11111110",
  26388=>"00000001",
  26389=>"00000001",
  26390=>"11111111",
  26391=>"00000000",
  26392=>"00000010",
  26393=>"00000010",
  26394=>"00000000",
  26395=>"00000010",
  26396=>"00000000",
  26397=>"00000001",
  26398=>"11111110",
  26399=>"00000000",
  26400=>"00000000",
  26401=>"11111110",
  26402=>"00000001",
  26403=>"11111111",
  26404=>"11111111",
  26405=>"00000001",
  26406=>"00000001",
  26407=>"00000000",
  26408=>"00000001",
  26409=>"00000000",
  26410=>"00000001",
  26411=>"00000001",
  26412=>"00000000",
  26413=>"11111101",
  26414=>"11111111",
  26415=>"11111110",
  26416=>"11111111",
  26417=>"00000000",
  26418=>"11111111",
  26419=>"11111111",
  26420=>"11111111",
  26421=>"11111111",
  26422=>"00000001",
  26423=>"11111111",
  26424=>"00000010",
  26425=>"00000001",
  26426=>"11111111",
  26427=>"00000001",
  26428=>"00000000",
  26429=>"11111111",
  26430=>"11111110",
  26431=>"11111110",
  26432=>"00000001",
  26433=>"00000010",
  26434=>"00000001",
  26435=>"00000000",
  26436=>"11111111",
  26437=>"00000001",
  26438=>"00000000",
  26439=>"00000010",
  26440=>"11111111",
  26441=>"11111111",
  26442=>"00000000",
  26443=>"00000001",
  26444=>"00000000",
  26445=>"00000010",
  26446=>"00000001",
  26447=>"00000001",
  26448=>"11111111",
  26449=>"00000001",
  26450=>"11111111",
  26451=>"00000010",
  26452=>"11111111",
  26453=>"11111110",
  26454=>"11111110",
  26455=>"00000010",
  26456=>"00000001",
  26457=>"11111110",
  26458=>"11111111",
  26459=>"11111110",
  26460=>"00000000",
  26461=>"00000000",
  26462=>"11111111",
  26463=>"00000001",
  26464=>"11111110",
  26465=>"00000001",
  26466=>"00000000",
  26467=>"00000000",
  26468=>"00000000",
  26469=>"11111111",
  26470=>"00000000",
  26471=>"00000001",
  26472=>"00000001",
  26473=>"11111110",
  26474=>"11111111",
  26475=>"00000001",
  26476=>"11111111",
  26477=>"00000000",
  26478=>"00000000",
  26479=>"11111111",
  26480=>"11111110",
  26481=>"00000010",
  26482=>"11111101",
  26483=>"11111111",
  26484=>"00000010",
  26485=>"11111111",
  26486=>"11111110",
  26487=>"00000000",
  26488=>"00000000",
  26489=>"00000001",
  26490=>"00000010",
  26491=>"00000000",
  26492=>"11111111",
  26493=>"11111111",
  26494=>"00000000",
  26495=>"00000001",
  26496=>"00000001",
  26497=>"11111111",
  26498=>"11111110",
  26499=>"11111111",
  26500=>"11111111",
  26501=>"00000001",
  26502=>"11111111",
  26503=>"11111111",
  26504=>"00000001",
  26505=>"00000001",
  26506=>"00000011",
  26507=>"00000010",
  26508=>"11111110",
  26509=>"00000000",
  26510=>"11111111",
  26511=>"00000000",
  26512=>"00000001",
  26513=>"11111111",
  26514=>"00000000",
  26515=>"00000001",
  26516=>"00000001",
  26517=>"00000000",
  26518=>"11111111",
  26519=>"00000010",
  26520=>"00000000",
  26521=>"11111111",
  26522=>"00000000",
  26523=>"11111111",
  26524=>"00000000",
  26525=>"11111110",
  26526=>"11111111",
  26527=>"11111110",
  26528=>"00000000",
  26529=>"11111111",
  26530=>"00000000",
  26531=>"00000010",
  26532=>"00000011",
  26533=>"00000010",
  26534=>"11111101",
  26535=>"00000000",
  26536=>"00000001",
  26537=>"00000011",
  26538=>"00000000",
  26539=>"00000010",
  26540=>"00000001",
  26541=>"11111111",
  26542=>"11111111",
  26543=>"00000000",
  26544=>"00000000",
  26545=>"00000001",
  26546=>"00000000",
  26547=>"11111110",
  26548=>"11111111",
  26549=>"00000000",
  26550=>"00000001",
  26551=>"00000001",
  26552=>"00000000",
  26553=>"00000000",
  26554=>"11111110",
  26555=>"00000010",
  26556=>"00000001",
  26557=>"11111111",
  26558=>"11111110",
  26559=>"11111110",
  26560=>"11111111",
  26561=>"00000001",
  26562=>"11111111",
  26563=>"11111111",
  26564=>"00000000",
  26565=>"11111110",
  26566=>"11111111",
  26567=>"11111111",
  26568=>"11111111",
  26569=>"11111101",
  26570=>"11111111",
  26571=>"00000010",
  26572=>"11111110",
  26573=>"00000001",
  26574=>"11111111",
  26575=>"00000001",
  26576=>"00000000",
  26577=>"00000000",
  26578=>"00000010",
  26579=>"00000010",
  26580=>"00000010",
  26581=>"00000010",
  26582=>"00000000",
  26583=>"00000000",
  26584=>"11111111",
  26585=>"00000000",
  26586=>"11111111",
  26587=>"11111110",
  26588=>"00000010",
  26589=>"00000000",
  26590=>"00000000",
  26591=>"00000000",
  26592=>"11111110",
  26593=>"00000000",
  26594=>"00000001",
  26595=>"00000010",
  26596=>"00000001",
  26597=>"00000011",
  26598=>"00000000",
  26599=>"11111111",
  26600=>"00000001",
  26601=>"00000000",
  26602=>"00000000",
  26603=>"11111111",
  26604=>"11111110",
  26605=>"11111111",
  26606=>"00000001",
  26607=>"00000000",
  26608=>"11111110",
  26609=>"00000000",
  26610=>"11111110",
  26611=>"00000000",
  26612=>"11111111",
  26613=>"00000010",
  26614=>"11111111",
  26615=>"00000001",
  26616=>"00000001",
  26617=>"00000010",
  26618=>"00000010",
  26619=>"00000010",
  26620=>"00000000",
  26621=>"11111111",
  26622=>"00000010",
  26623=>"00000000",
  26624=>"00000010",
  26625=>"00000010",
  26626=>"11111111",
  26627=>"00000000",
  26628=>"00000001",
  26629=>"00000000",
  26630=>"00000010",
  26631=>"11111111",
  26632=>"00000001",
  26633=>"00000011",
  26634=>"00000001",
  26635=>"00000010",
  26636=>"00000000",
  26637=>"00000000",
  26638=>"00000000",
  26639=>"00000001",
  26640=>"00000010",
  26641=>"00000001",
  26642=>"11111111",
  26643=>"11111110",
  26644=>"00000001",
  26645=>"00000010",
  26646=>"00000001",
  26647=>"11111111",
  26648=>"00000001",
  26649=>"00000000",
  26650=>"00000011",
  26651=>"11111111",
  26652=>"00000000",
  26653=>"00000001",
  26654=>"00000000",
  26655=>"11111111",
  26656=>"00000000",
  26657=>"00000001",
  26658=>"11111101",
  26659=>"11111101",
  26660=>"11111111",
  26661=>"00000001",
  26662=>"00000010",
  26663=>"11111110",
  26664=>"00000001",
  26665=>"11111110",
  26666=>"11111111",
  26667=>"11111111",
  26668=>"00000000",
  26669=>"11111111",
  26670=>"00000010",
  26671=>"00000000",
  26672=>"11111111",
  26673=>"00000000",
  26674=>"00000001",
  26675=>"00000001",
  26676=>"11111110",
  26677=>"00000001",
  26678=>"11111110",
  26679=>"11111110",
  26680=>"11111111",
  26681=>"00000010",
  26682=>"11111111",
  26683=>"00000001",
  26684=>"00000001",
  26685=>"00000001",
  26686=>"11111110",
  26687=>"11111111",
  26688=>"00000001",
  26689=>"11111110",
  26690=>"11111111",
  26691=>"00000010",
  26692=>"00000010",
  26693=>"00000010",
  26694=>"11111111",
  26695=>"00000001",
  26696=>"11111110",
  26697=>"11111110",
  26698=>"11111110",
  26699=>"11111110",
  26700=>"00000000",
  26701=>"11111110",
  26702=>"00000000",
  26703=>"00000001",
  26704=>"00000000",
  26705=>"00000000",
  26706=>"00000000",
  26707=>"00000001",
  26708=>"00000011",
  26709=>"00000001",
  26710=>"00000001",
  26711=>"11111110",
  26712=>"00000001",
  26713=>"11111111",
  26714=>"00000001",
  26715=>"00000000",
  26716=>"11111110",
  26717=>"00000011",
  26718=>"00000001",
  26719=>"00000001",
  26720=>"11111111",
  26721=>"00000001",
  26722=>"00000001",
  26723=>"11111110",
  26724=>"00000000",
  26725=>"00000001",
  26726=>"00000001",
  26727=>"11111110",
  26728=>"00000010",
  26729=>"11111110",
  26730=>"11111111",
  26731=>"11111111",
  26732=>"11111110",
  26733=>"00000001",
  26734=>"11111110",
  26735=>"00000001",
  26736=>"11111110",
  26737=>"00000000",
  26738=>"00000000",
  26739=>"11111110",
  26740=>"11111110",
  26741=>"11111111",
  26742=>"11111111",
  26743=>"00000010",
  26744=>"00000000",
  26745=>"11111110",
  26746=>"11111111",
  26747=>"00000000",
  26748=>"00000010",
  26749=>"00000000",
  26750=>"11111111",
  26751=>"11111111",
  26752=>"00000000",
  26753=>"11111111",
  26754=>"11111110",
  26755=>"11111111",
  26756=>"00000010",
  26757=>"11111110",
  26758=>"11111110",
  26759=>"00000010",
  26760=>"00000000",
  26761=>"11111111",
  26762=>"00000010",
  26763=>"11111111",
  26764=>"00000001",
  26765=>"11111100",
  26766=>"00000010",
  26767=>"00000010",
  26768=>"00000001",
  26769=>"11111111",
  26770=>"00000110",
  26771=>"00000001",
  26772=>"00000000",
  26773=>"11111110",
  26774=>"00000000",
  26775=>"11111111",
  26776=>"11111110",
  26777=>"00000000",
  26778=>"00000001",
  26779=>"11111110",
  26780=>"11111111",
  26781=>"11111110",
  26782=>"11111110",
  26783=>"00000001",
  26784=>"11111111",
  26785=>"00000000",
  26786=>"00000001",
  26787=>"00000010",
  26788=>"00000000",
  26789=>"11111110",
  26790=>"00000000",
  26791=>"00000000",
  26792=>"11111110",
  26793=>"00000000",
  26794=>"00000001",
  26795=>"11111111",
  26796=>"11111111",
  26797=>"00000000",
  26798=>"11111110",
  26799=>"11111110",
  26800=>"00000001",
  26801=>"11111110",
  26802=>"00000001",
  26803=>"00000000",
  26804=>"11111110",
  26805=>"11111110",
  26806=>"00000000",
  26807=>"11111111",
  26808=>"00000001",
  26809=>"11111110",
  26810=>"11111111",
  26811=>"11111111",
  26812=>"11111111",
  26813=>"00000000",
  26814=>"00000001",
  26815=>"00000000",
  26816=>"00000001",
  26817=>"00000001",
  26818=>"11111111",
  26819=>"00000000",
  26820=>"00000001",
  26821=>"00000010",
  26822=>"00000010",
  26823=>"11111110",
  26824=>"11111111",
  26825=>"00000001",
  26826=>"11111111",
  26827=>"00000011",
  26828=>"11111111",
  26829=>"11111111",
  26830=>"11111101",
  26831=>"11111110",
  26832=>"00000000",
  26833=>"00000010",
  26834=>"00000000",
  26835=>"00000001",
  26836=>"11111110",
  26837=>"11111111",
  26838=>"00000010",
  26839=>"00000001",
  26840=>"00000000",
  26841=>"00000001",
  26842=>"11111110",
  26843=>"00000010",
  26844=>"11111101",
  26845=>"00000011",
  26846=>"00000000",
  26847=>"00000001",
  26848=>"00000010",
  26849=>"00000010",
  26850=>"11111111",
  26851=>"00000000",
  26852=>"00000001",
  26853=>"11111111",
  26854=>"00000001",
  26855=>"11111111",
  26856=>"00000010",
  26857=>"00000001",
  26858=>"11111111",
  26859=>"00000010",
  26860=>"11111111",
  26861=>"11111111",
  26862=>"00000010",
  26863=>"00000001",
  26864=>"11111110",
  26865=>"11111111",
  26866=>"11111111",
  26867=>"00000000",
  26868=>"00000000",
  26869=>"00000001",
  26870=>"11111110",
  26871=>"00000001",
  26872=>"00000010",
  26873=>"11111111",
  26874=>"00000001",
  26875=>"00000001",
  26876=>"11111111",
  26877=>"11111111",
  26878=>"00000001",
  26879=>"00000010",
  26880=>"11111110",
  26881=>"11111111",
  26882=>"00000000",
  26883=>"00000001",
  26884=>"11111110",
  26885=>"00000000",
  26886=>"11111110",
  26887=>"00000010",
  26888=>"11111111",
  26889=>"11111111",
  26890=>"00000001",
  26891=>"00000001",
  26892=>"00000000",
  26893=>"00000011",
  26894=>"00000000",
  26895=>"00000000",
  26896=>"11111111",
  26897=>"00000001",
  26898=>"00000001",
  26899=>"00000000",
  26900=>"11111111",
  26901=>"00000000",
  26902=>"00000001",
  26903=>"11111110",
  26904=>"11111111",
  26905=>"00000001",
  26906=>"11111110",
  26907=>"11111110",
  26908=>"00000001",
  26909=>"00000001",
  26910=>"11111110",
  26911=>"00000001",
  26912=>"00000001",
  26913=>"11111111",
  26914=>"00000001",
  26915=>"11111110",
  26916=>"00000010",
  26917=>"00000001",
  26918=>"11111110",
  26919=>"00000001",
  26920=>"00000010",
  26921=>"00000010",
  26922=>"11111111",
  26923=>"11111111",
  26924=>"00000001",
  26925=>"00000010",
  26926=>"11111101",
  26927=>"00000010",
  26928=>"00000001",
  26929=>"00000001",
  26930=>"11111111",
  26931=>"11111110",
  26932=>"00000001",
  26933=>"11111111",
  26934=>"00000000",
  26935=>"00000001",
  26936=>"00000000",
  26937=>"00000000",
  26938=>"11111101",
  26939=>"00000000",
  26940=>"00000000",
  26941=>"11111101",
  26942=>"11111111",
  26943=>"11111111",
  26944=>"11111111",
  26945=>"00000000",
  26946=>"11111111",
  26947=>"11111111",
  26948=>"11111111",
  26949=>"00000000",
  26950=>"00000001",
  26951=>"11111111",
  26952=>"00000000",
  26953=>"11111111",
  26954=>"00000001",
  26955=>"00000010",
  26956=>"00000010",
  26957=>"00000001",
  26958=>"00000001",
  26959=>"00000000",
  26960=>"00000001",
  26961=>"11111111",
  26962=>"00000010",
  26963=>"11111111",
  26964=>"11111111",
  26965=>"00000001",
  26966=>"11111110",
  26967=>"00000000",
  26968=>"00000010",
  26969=>"11111101",
  26970=>"00000001",
  26971=>"11111110",
  26972=>"11111111",
  26973=>"00000010",
  26974=>"11111111",
  26975=>"00000000",
  26976=>"00000000",
  26977=>"00000010",
  26978=>"00000001",
  26979=>"00000010",
  26980=>"11111111",
  26981=>"00000000",
  26982=>"11111111",
  26983=>"11111110",
  26984=>"00000000",
  26985=>"00000010",
  26986=>"11111110",
  26987=>"00000001",
  26988=>"00000001",
  26989=>"11111110",
  26990=>"00000000",
  26991=>"00000001",
  26992=>"00000000",
  26993=>"00000000",
  26994=>"00000001",
  26995=>"11111111",
  26996=>"00000001",
  26997=>"00000001",
  26998=>"11111110",
  26999=>"00000001",
  27000=>"00000010",
  27001=>"11111111",
  27002=>"00000001",
  27003=>"11111110",
  27004=>"11111110",
  27005=>"11111111",
  27006=>"00000000",
  27007=>"00000001",
  27008=>"00000001",
  27009=>"00000000",
  27010=>"00000000",
  27011=>"11111110",
  27012=>"00000011",
  27013=>"00000001",
  27014=>"00000001",
  27015=>"00000001",
  27016=>"00000000",
  27017=>"00000010",
  27018=>"00000000",
  27019=>"00000001",
  27020=>"11111110",
  27021=>"00000010",
  27022=>"00000011",
  27023=>"00000001",
  27024=>"11111111",
  27025=>"11111111",
  27026=>"00000001",
  27027=>"11111111",
  27028=>"00000001",
  27029=>"00000010",
  27030=>"00000001",
  27031=>"00000000",
  27032=>"11111111",
  27033=>"00000001",
  27034=>"00000001",
  27035=>"11111101",
  27036=>"00000010",
  27037=>"11111110",
  27038=>"00000001",
  27039=>"00000001",
  27040=>"00000000",
  27041=>"11111111",
  27042=>"00000001",
  27043=>"00000000",
  27044=>"00000010",
  27045=>"00000000",
  27046=>"11111110",
  27047=>"00000000",
  27048=>"00000000",
  27049=>"00000001",
  27050=>"00000010",
  27051=>"11111111",
  27052=>"00000001",
  27053=>"00000000",
  27054=>"00000001",
  27055=>"11111111",
  27056=>"11111111",
  27057=>"11111111",
  27058=>"11111111",
  27059=>"00000001",
  27060=>"11111111",
  27061=>"11111110",
  27062=>"11111110",
  27063=>"11111111",
  27064=>"00000001",
  27065=>"00000001",
  27066=>"00000001",
  27067=>"00000011",
  27068=>"11111101",
  27069=>"11111111",
  27070=>"00000000",
  27071=>"00000000",
  27072=>"00000000",
  27073=>"00000000",
  27074=>"11111111",
  27075=>"00000000",
  27076=>"00000001",
  27077=>"11111111",
  27078=>"11111111",
  27079=>"11111111",
  27080=>"11111110",
  27081=>"11111111",
  27082=>"00000000",
  27083=>"00000001",
  27084=>"00000001",
  27085=>"11111111",
  27086=>"00000001",
  27087=>"00000001",
  27088=>"00000000",
  27089=>"11111111",
  27090=>"11111101",
  27091=>"00000001",
  27092=>"00000000",
  27093=>"00000000",
  27094=>"11111110",
  27095=>"11111111",
  27096=>"11111110",
  27097=>"11111111",
  27098=>"11111101",
  27099=>"00000000",
  27100=>"00000001",
  27101=>"00000001",
  27102=>"00000001",
  27103=>"11111111",
  27104=>"11111110",
  27105=>"00000001",
  27106=>"00000011",
  27107=>"11111110",
  27108=>"11111101",
  27109=>"11111111",
  27110=>"00000001",
  27111=>"11111110",
  27112=>"11111111",
  27113=>"00000001",
  27114=>"00000001",
  27115=>"11111111",
  27116=>"11111110",
  27117=>"11111111",
  27118=>"11111111",
  27119=>"00000001",
  27120=>"00000000",
  27121=>"00000001",
  27122=>"00000000",
  27123=>"00000001",
  27124=>"00000000",
  27125=>"00000010",
  27126=>"11111101",
  27127=>"00000001",
  27128=>"11111111",
  27129=>"11111111",
  27130=>"11111110",
  27131=>"00000010",
  27132=>"00000010",
  27133=>"00000001",
  27134=>"00000010",
  27135=>"11111111",
  27136=>"00000000",
  27137=>"00000001",
  27138=>"00000001",
  27139=>"00000001",
  27140=>"00000010",
  27141=>"00000010",
  27142=>"00000000",
  27143=>"11111111",
  27144=>"00000001",
  27145=>"00000000",
  27146=>"00000000",
  27147=>"00000010",
  27148=>"00000001",
  27149=>"00000001",
  27150=>"00000000",
  27151=>"11111111",
  27152=>"11111111",
  27153=>"11111110",
  27154=>"11111110",
  27155=>"00000010",
  27156=>"00000001",
  27157=>"11111110",
  27158=>"00000001",
  27159=>"00000010",
  27160=>"11111110",
  27161=>"00000010",
  27162=>"00000001",
  27163=>"11111110",
  27164=>"00000000",
  27165=>"11111111",
  27166=>"00000000",
  27167=>"00000001",
  27168=>"00000000",
  27169=>"00000011",
  27170=>"00000000",
  27171=>"11111110",
  27172=>"00000001",
  27173=>"11111110",
  27174=>"00000000",
  27175=>"00000010",
  27176=>"00000000",
  27177=>"00000001",
  27178=>"00000010",
  27179=>"00000000",
  27180=>"00000000",
  27181=>"00000000",
  27182=>"00000010",
  27183=>"00000000",
  27184=>"00000000",
  27185=>"00000010",
  27186=>"11111111",
  27187=>"11111111",
  27188=>"11111111",
  27189=>"11111110",
  27190=>"11111111",
  27191=>"00000000",
  27192=>"00000001",
  27193=>"00000001",
  27194=>"11111111",
  27195=>"11111111",
  27196=>"11111111",
  27197=>"00000010",
  27198=>"11111111",
  27199=>"00000000",
  27200=>"00000001",
  27201=>"11111111",
  27202=>"00000000",
  27203=>"00000001",
  27204=>"00000000",
  27205=>"00000001",
  27206=>"00000000",
  27207=>"11111111",
  27208=>"00000000",
  27209=>"00000000",
  27210=>"00000000",
  27211=>"11111111",
  27212=>"11111111",
  27213=>"11111110",
  27214=>"00000001",
  27215=>"00000001",
  27216=>"11111111",
  27217=>"11111111",
  27218=>"11111110",
  27219=>"11111111",
  27220=>"11111111",
  27221=>"11111110",
  27222=>"00000000",
  27223=>"00000001",
  27224=>"11111111",
  27225=>"11111111",
  27226=>"11111111",
  27227=>"11111111",
  27228=>"11111110",
  27229=>"11111110",
  27230=>"00000000",
  27231=>"00000001",
  27232=>"00000000",
  27233=>"11111110",
  27234=>"00000000",
  27235=>"00000000",
  27236=>"11111110",
  27237=>"11111110",
  27238=>"00000000",
  27239=>"00000001",
  27240=>"11111111",
  27241=>"00000010",
  27242=>"00000001",
  27243=>"00000000",
  27244=>"11111111",
  27245=>"11111111",
  27246=>"00000000",
  27247=>"11111110",
  27248=>"11111111",
  27249=>"11111111",
  27250=>"11111111",
  27251=>"00000000",
  27252=>"00000001",
  27253=>"00000000",
  27254=>"00000000",
  27255=>"00000010",
  27256=>"11111110",
  27257=>"00000000",
  27258=>"11111110",
  27259=>"11111111",
  27260=>"11111110",
  27261=>"00000000",
  27262=>"11111111",
  27263=>"00000001",
  27264=>"00000000",
  27265=>"00000001",
  27266=>"11111111",
  27267=>"00000000",
  27268=>"00000001",
  27269=>"00000001",
  27270=>"11111110",
  27271=>"00000010",
  27272=>"00000010",
  27273=>"00000000",
  27274=>"11111111",
  27275=>"00000001",
  27276=>"00000010",
  27277=>"00000001",
  27278=>"00000010",
  27279=>"11111111",
  27280=>"11111110",
  27281=>"11111111",
  27282=>"00000000",
  27283=>"00000000",
  27284=>"11111110",
  27285=>"11111111",
  27286=>"00000000",
  27287=>"00000000",
  27288=>"00000001",
  27289=>"00000001",
  27290=>"00000000",
  27291=>"00000010",
  27292=>"00000001",
  27293=>"11111111",
  27294=>"00000001",
  27295=>"11111110",
  27296=>"11111111",
  27297=>"11111111",
  27298=>"00000001",
  27299=>"00000001",
  27300=>"00000001",
  27301=>"00000000",
  27302=>"00000001",
  27303=>"00000010",
  27304=>"00000000",
  27305=>"00000000",
  27306=>"00000000",
  27307=>"11111111",
  27308=>"11111111",
  27309=>"00000000",
  27310=>"00000000",
  27311=>"11111110",
  27312=>"00000001",
  27313=>"11111111",
  27314=>"00000011",
  27315=>"00000001",
  27316=>"00000000",
  27317=>"11111111",
  27318=>"11111111",
  27319=>"11111110",
  27320=>"11111111",
  27321=>"00000000",
  27322=>"11111110",
  27323=>"00000000",
  27324=>"11111111",
  27325=>"11111110",
  27326=>"00000000",
  27327=>"11111111",
  27328=>"11111110",
  27329=>"11111111",
  27330=>"11111111",
  27331=>"11111111",
  27332=>"11111111",
  27333=>"00000000",
  27334=>"00000010",
  27335=>"11111100",
  27336=>"00000000",
  27337=>"00000001",
  27338=>"11111110",
  27339=>"00000001",
  27340=>"11111110",
  27341=>"00000001",
  27342=>"00000001",
  27343=>"00000001",
  27344=>"00000010",
  27345=>"00000000",
  27346=>"00000001",
  27347=>"00000000",
  27348=>"11111111",
  27349=>"11111100",
  27350=>"00000001",
  27351=>"00000001",
  27352=>"00000001",
  27353=>"11111110",
  27354=>"00000010",
  27355=>"00000001",
  27356=>"11111111",
  27357=>"11111111",
  27358=>"11111110",
  27359=>"00000000",
  27360=>"00000000",
  27361=>"00000001",
  27362=>"00000000",
  27363=>"11111111",
  27364=>"00000011",
  27365=>"00000000",
  27366=>"00000000",
  27367=>"00000001",
  27368=>"00000001",
  27369=>"00000001",
  27370=>"00000000",
  27371=>"00000010",
  27372=>"00000000",
  27373=>"11111111",
  27374=>"00000010",
  27375=>"00000000",
  27376=>"11111111",
  27377=>"00000000",
  27378=>"00000010",
  27379=>"00000000",
  27380=>"00000001",
  27381=>"00000001",
  27382=>"00000000",
  27383=>"11111101",
  27384=>"00000000",
  27385=>"00000011",
  27386=>"00000000",
  27387=>"00000001",
  27388=>"11111111",
  27389=>"00000010",
  27390=>"11111110",
  27391=>"00000001",
  27392=>"11111111",
  27393=>"00000000",
  27394=>"11111111",
  27395=>"11111110",
  27396=>"00000001",
  27397=>"00000001",
  27398=>"00000010",
  27399=>"00000010",
  27400=>"11111111",
  27401=>"00000000",
  27402=>"00000000",
  27403=>"00000001",
  27404=>"00000000",
  27405=>"00000000",
  27406=>"00000000",
  27407=>"00000001",
  27408=>"00000001",
  27409=>"11111101",
  27410=>"11111111",
  27411=>"00000010",
  27412=>"00000010",
  27413=>"11111111",
  27414=>"00000010",
  27415=>"00000000",
  27416=>"11111111",
  27417=>"11111111",
  27418=>"11111111",
  27419=>"00000000",
  27420=>"00000010",
  27421=>"00000000",
  27422=>"11111111",
  27423=>"11111111",
  27424=>"11111101",
  27425=>"00000000",
  27426=>"00000001",
  27427=>"00000100",
  27428=>"11111101",
  27429=>"00000000",
  27430=>"00000000",
  27431=>"11111111",
  27432=>"00000011",
  27433=>"00000000",
  27434=>"00000001",
  27435=>"00000000",
  27436=>"00000001",
  27437=>"11111111",
  27438=>"11111110",
  27439=>"00000001",
  27440=>"00000000",
  27441=>"00000000",
  27442=>"00000001",
  27443=>"11111110",
  27444=>"00000001",
  27445=>"00000000",
  27446=>"00000001",
  27447=>"00000010",
  27448=>"00000001",
  27449=>"00000010",
  27450=>"00000010",
  27451=>"00000001",
  27452=>"00000000",
  27453=>"00000010",
  27454=>"00000010",
  27455=>"11111111",
  27456=>"00000000",
  27457=>"00000000",
  27458=>"11111110",
  27459=>"11111111",
  27460=>"00000000",
  27461=>"11111101",
  27462=>"00000001",
  27463=>"11111111",
  27464=>"00000000",
  27465=>"00000010",
  27466=>"00000001",
  27467=>"11111110",
  27468=>"00000010",
  27469=>"00000001",
  27470=>"11111110",
  27471=>"11111110",
  27472=>"00000000",
  27473=>"11111111",
  27474=>"11111111",
  27475=>"11111111",
  27476=>"00000001",
  27477=>"00000001",
  27478=>"11111100",
  27479=>"11111111",
  27480=>"00000010",
  27481=>"00000000",
  27482=>"11111111",
  27483=>"00000000",
  27484=>"00000001",
  27485=>"11111110",
  27486=>"00000001",
  27487=>"00000010",
  27488=>"00000000",
  27489=>"00000000",
  27490=>"00000000",
  27491=>"00000010",
  27492=>"11111111",
  27493=>"11111101",
  27494=>"11111111",
  27495=>"00000001",
  27496=>"00000001",
  27497=>"00000000",
  27498=>"11111111",
  27499=>"00000000",
  27500=>"00000010",
  27501=>"11111111",
  27502=>"00000000",
  27503=>"11111111",
  27504=>"00000000",
  27505=>"11111110",
  27506=>"11111111",
  27507=>"00000000",
  27508=>"11111110",
  27509=>"00000000",
  27510=>"00000010",
  27511=>"00000010",
  27512=>"00000001",
  27513=>"00000001",
  27514=>"00000000",
  27515=>"00000000",
  27516=>"00000001",
  27517=>"11111110",
  27518=>"11111111",
  27519=>"00000000",
  27520=>"11111111",
  27521=>"00000001",
  27522=>"00000000",
  27523=>"00000010",
  27524=>"11111110",
  27525=>"00000000",
  27526=>"00000001",
  27527=>"00000010",
  27528=>"00000000",
  27529=>"00000000",
  27530=>"00000001",
  27531=>"00000000",
  27532=>"11111110",
  27533=>"11111111",
  27534=>"00000001",
  27535=>"00000001",
  27536=>"11111111",
  27537=>"11111111",
  27538=>"11111111",
  27539=>"00000001",
  27540=>"11111111",
  27541=>"00000010",
  27542=>"00000000",
  27543=>"11111111",
  27544=>"00000001",
  27545=>"00000010",
  27546=>"00000001",
  27547=>"00000001",
  27548=>"00000000",
  27549=>"00000000",
  27550=>"00000000",
  27551=>"00000001",
  27552=>"00000000",
  27553=>"00000010",
  27554=>"00000000",
  27555=>"00000000",
  27556=>"00000011",
  27557=>"00000010",
  27558=>"00000000",
  27559=>"00000000",
  27560=>"00000001",
  27561=>"00000000",
  27562=>"00000001",
  27563=>"00000001",
  27564=>"00000000",
  27565=>"00000000",
  27566=>"00000000",
  27567=>"00000000",
  27568=>"00000000",
  27569=>"11111111",
  27570=>"11111110",
  27571=>"00000011",
  27572=>"11111111",
  27573=>"00000000",
  27574=>"11111110",
  27575=>"00000011",
  27576=>"00000001",
  27577=>"11111111",
  27578=>"00000000",
  27579=>"00000001",
  27580=>"00000001",
  27581=>"11111110",
  27582=>"11111110",
  27583=>"11111111",
  27584=>"00000010",
  27585=>"00000000",
  27586=>"00000001",
  27587=>"00000000",
  27588=>"11111110",
  27589=>"11111111",
  27590=>"11111111",
  27591=>"00000010",
  27592=>"00000001",
  27593=>"00000011",
  27594=>"00000001",
  27595=>"00000000",
  27596=>"11111101",
  27597=>"00000010",
  27598=>"00000011",
  27599=>"00000001",
  27600=>"11111111",
  27601=>"00000010",
  27602=>"00000001",
  27603=>"11111110",
  27604=>"00000000",
  27605=>"11111111",
  27606=>"00000000",
  27607=>"11111110",
  27608=>"11111111",
  27609=>"11111111",
  27610=>"00000001",
  27611=>"11111111",
  27612=>"11111110",
  27613=>"00000000",
  27614=>"00000001",
  27615=>"11111111",
  27616=>"00000010",
  27617=>"00000000",
  27618=>"00000010",
  27619=>"11111111",
  27620=>"00000010",
  27621=>"00000010",
  27622=>"11111110",
  27623=>"00000010",
  27624=>"00000001",
  27625=>"00000000",
  27626=>"11111110",
  27627=>"00000011",
  27628=>"00000000",
  27629=>"11111111",
  27630=>"00000001",
  27631=>"00000001",
  27632=>"11111110",
  27633=>"11111111",
  27634=>"00000010",
  27635=>"11111111",
  27636=>"11111111",
  27637=>"00000000",
  27638=>"00000001",
  27639=>"11111110",
  27640=>"11111111",
  27641=>"00000000",
  27642=>"00000001",
  27643=>"11111111",
  27644=>"00000001",
  27645=>"00000001",
  27646=>"00000000",
  27647=>"00000011",
  27648=>"00000000",
  27649=>"11111111",
  27650=>"00000000",
  27651=>"11111111",
  27652=>"00000000",
  27653=>"00000000",
  27654=>"00000000",
  27655=>"00000000",
  27656=>"00000000",
  27657=>"00000000",
  27658=>"00000001",
  27659=>"00000000",
  27660=>"11111111",
  27661=>"00000000",
  27662=>"00000001",
  27663=>"00000000",
  27664=>"00000000",
  27665=>"00000001",
  27666=>"00000000",
  27667=>"00000001",
  27668=>"00000000",
  27669=>"00000000",
  27670=>"00000000",
  27671=>"00000000",
  27672=>"00000000",
  27673=>"00000000",
  27674=>"11111111",
  27675=>"00000000",
  27676=>"00000000",
  27677=>"11111111",
  27678=>"00000000",
  27679=>"00000000",
  27680=>"00000000",
  27681=>"00000000",
  27682=>"00000000",
  27683=>"00000000",
  27684=>"00000000",
  27685=>"00000000",
  27686=>"00000000",
  27687=>"00000000",
  27688=>"00000001",
  27689=>"00000000",
  27690=>"00000000",
  27691=>"00000000",
  27692=>"00000000",
  27693=>"00000000",
  27694=>"00000001",
  27695=>"00000000",
  27696=>"00000000",
  27697=>"00000000",
  27698=>"00000000",
  27699=>"00000000",
  27700=>"00000000",
  27701=>"00000000",
  27702=>"00000010",
  27703=>"11111111",
  27704=>"00000001",
  27705=>"00000000",
  27706=>"00000000",
  27707=>"00000000",
  27708=>"00000001",
  27709=>"11111111",
  27710=>"00000000",
  27711=>"00000000",
  27712=>"00000000",
  27713=>"00000000",
  27714=>"00000000",
  27715=>"00000000",
  27716=>"00000000",
  27717=>"00000000",
  27718=>"00000000",
  27719=>"11111111",
  27720=>"00000000",
  27721=>"00000000",
  27722=>"11111111",
  27723=>"00000001",
  27724=>"00000000",
  27725=>"00000000",
  27726=>"00000000",
  27727=>"00000000",
  27728=>"00000000",
  27729=>"00000000",
  27730=>"00000000",
  27731=>"00000000",
  27732=>"00000000",
  27733=>"00000001",
  27734=>"00000000",
  27735=>"00000000",
  27736=>"00000000",
  27737=>"00000000",
  27738=>"00000001",
  27739=>"11111111",
  27740=>"00000000",
  27741=>"00000000",
  27742=>"00000000",
  27743=>"00000000",
  27744=>"00000001",
  27745=>"00000000",
  27746=>"00000000",
  27747=>"00000000",
  27748=>"00000000",
  27749=>"00000000",
  27750=>"11111111",
  27751=>"00000001",
  27752=>"00000000",
  27753=>"00000000",
  27754=>"00000000",
  27755=>"11111101",
  27756=>"00000000",
  27757=>"00000000",
  27758=>"00000000",
  27759=>"00000000",
  27760=>"00000000",
  27761=>"11111111",
  27762=>"00000000",
  27763=>"00000000",
  27764=>"00000000",
  27765=>"00000000",
  27766=>"00000000",
  27767=>"00000000",
  27768=>"00000000",
  27769=>"00000000",
  27770=>"00000000",
  27771=>"00000000",
  27772=>"00000000",
  27773=>"11111111",
  27774=>"00000001",
  27775=>"00000000",
  27776=>"00000000",
  27777=>"00000000",
  27778=>"00000001",
  27779=>"00000000",
  27780=>"00000000",
  27781=>"11111111",
  27782=>"00000000",
  27783=>"00000000",
  27784=>"11111111",
  27785=>"00000001",
  27786=>"11111111",
  27787=>"00000000",
  27788=>"00000000",
  27789=>"11111111",
  27790=>"00000000",
  27791=>"00000000",
  27792=>"00000000",
  27793=>"00000001",
  27794=>"00000000",
  27795=>"00000000",
  27796=>"00000000",
  27797=>"00000000",
  27798=>"00000000",
  27799=>"00000001",
  27800=>"00000000",
  27801=>"00000000",
  27802=>"00000000",
  27803=>"00000000",
  27804=>"00000010",
  27805=>"11111111",
  27806=>"00000000",
  27807=>"00000000",
  27808=>"00000000",
  27809=>"00000000",
  27810=>"00000001",
  27811=>"00000000",
  27812=>"00000010",
  27813=>"00000000",
  27814=>"00000001",
  27815=>"00000001",
  27816=>"00000000",
  27817=>"00000001",
  27818=>"00000001",
  27819=>"00000000",
  27820=>"11111111",
  27821=>"00000000",
  27822=>"00000000",
  27823=>"00000000",
  27824=>"00000000",
  27825=>"00000000",
  27826=>"00000000",
  27827=>"00000000",
  27828=>"00000000",
  27829=>"00000000",
  27830=>"00000000",
  27831=>"00000000",
  27832=>"00000000",
  27833=>"00000000",
  27834=>"00000000",
  27835=>"00000000",
  27836=>"00000000",
  27837=>"11111111",
  27838=>"00000000",
  27839=>"00000000",
  27840=>"00000001",
  27841=>"11111111",
  27842=>"00000000",
  27843=>"00000000",
  27844=>"11111111",
  27845=>"00000000",
  27846=>"00000000",
  27847=>"00000001",
  27848=>"00000000",
  27849=>"00000001",
  27850=>"00000000",
  27851=>"00000000",
  27852=>"00000000",
  27853=>"00000000",
  27854=>"11111111",
  27855=>"00000000",
  27856=>"00000000",
  27857=>"00000000",
  27858=>"11111101",
  27859=>"00000001",
  27860=>"00000000",
  27861=>"00000000",
  27862=>"00000001",
  27863=>"00000000",
  27864=>"00000000",
  27865=>"00000000",
  27866=>"11111111",
  27867=>"00000000",
  27868=>"00000000",
  27869=>"00000000",
  27870=>"11111111",
  27871=>"00000000",
  27872=>"00000000",
  27873=>"00000000",
  27874=>"00000000",
  27875=>"00000000",
  27876=>"00000000",
  27877=>"00000000",
  27878=>"00000000",
  27879=>"00000000",
  27880=>"00000000",
  27881=>"00000000",
  27882=>"00000000",
  27883=>"00000001",
  27884=>"00000001",
  27885=>"00000000",
  27886=>"11111111",
  27887=>"11111111",
  27888=>"00000000",
  27889=>"00000000",
  27890=>"00000000",
  27891=>"00000000",
  27892=>"00000000",
  27893=>"00000000",
  27894=>"11111111",
  27895=>"00000000",
  27896=>"00000000",
  27897=>"11111111",
  27898=>"00000000",
  27899=>"00000000",
  27900=>"00000000",
  27901=>"00000000",
  27902=>"00000000",
  27903=>"00000001",
  27904=>"00000000",
  27905=>"00000000",
  27906=>"00000000",
  27907=>"00000000",
  27908=>"00000000",
  27909=>"00000000",
  27910=>"11111111",
  27911=>"00000000",
  27912=>"00000000",
  27913=>"00000000",
  27914=>"00000000",
  27915=>"00000000",
  27916=>"00000000",
  27917=>"00000000",
  27918=>"00000000",
  27919=>"00000000",
  27920=>"00000000",
  27921=>"00000000",
  27922=>"11111111",
  27923=>"00000000",
  27924=>"11111111",
  27925=>"00000000",
  27926=>"00000000",
  27927=>"00000000",
  27928=>"00000000",
  27929=>"00000000",
  27930=>"00000000",
  27931=>"00000000",
  27932=>"11111111",
  27933=>"00000000",
  27934=>"00000001",
  27935=>"00000000",
  27936=>"00000000",
  27937=>"00000000",
  27938=>"00000010",
  27939=>"00000000",
  27940=>"00000000",
  27941=>"00000000",
  27942=>"00000000",
  27943=>"00000000",
  27944=>"00000000",
  27945=>"11111111",
  27946=>"00000000",
  27947=>"00000000",
  27948=>"00000000",
  27949=>"11111101",
  27950=>"00000000",
  27951=>"00000001",
  27952=>"00000000",
  27953=>"00000000",
  27954=>"00000000",
  27955=>"00000000",
  27956=>"00000001",
  27957=>"00000000",
  27958=>"00000000",
  27959=>"00000000",
  27960=>"00000000",
  27961=>"00000001",
  27962=>"11111111",
  27963=>"00000000",
  27964=>"11111111",
  27965=>"00000000",
  27966=>"00000000",
  27967=>"00000001",
  27968=>"11111101",
  27969=>"00000000",
  27970=>"00000000",
  27971=>"11111111",
  27972=>"11111110",
  27973=>"00000000",
  27974=>"00000000",
  27975=>"00000001",
  27976=>"00000000",
  27977=>"00000000",
  27978=>"00000000",
  27979=>"00000000",
  27980=>"00000000",
  27981=>"00000000",
  27982=>"11111111",
  27983=>"00000000",
  27984=>"00000000",
  27985=>"00000000",
  27986=>"00000000",
  27987=>"00000000",
  27988=>"00000000",
  27989=>"00000000",
  27990=>"11111111",
  27991=>"00000000",
  27992=>"00000000",
  27993=>"00000000",
  27994=>"00000000",
  27995=>"00000000",
  27996=>"00000001",
  27997=>"00000000",
  27998=>"00000000",
  27999=>"00000000",
  28000=>"00000000",
  28001=>"00000000",
  28002=>"00000000",
  28003=>"00000000",
  28004=>"11111111",
  28005=>"00000000",
  28006=>"00000000",
  28007=>"00000000",
  28008=>"00000000",
  28009=>"00000000",
  28010=>"11111111",
  28011=>"00000000",
  28012=>"00000000",
  28013=>"00000000",
  28014=>"00000000",
  28015=>"00000000",
  28016=>"11111110",
  28017=>"00000000",
  28018=>"00000000",
  28019=>"00000000",
  28020=>"00000000",
  28021=>"00000000",
  28022=>"00000000",
  28023=>"00000000",
  28024=>"00000000",
  28025=>"00000000",
  28026=>"00000000",
  28027=>"00000000",
  28028=>"00000000",
  28029=>"00000000",
  28030=>"11111111",
  28031=>"00000000",
  28032=>"00000000",
  28033=>"11111111",
  28034=>"00000000",
  28035=>"11111111",
  28036=>"11111111",
  28037=>"00000000",
  28038=>"00000000",
  28039=>"11111111",
  28040=>"00000000",
  28041=>"00000000",
  28042=>"00000000",
  28043=>"00000000",
  28044=>"00000000",
  28045=>"00000001",
  28046=>"00000000",
  28047=>"00000000",
  28048=>"00000001",
  28049=>"11111111",
  28050=>"00000000",
  28051=>"00000000",
  28052=>"00000000",
  28053=>"00000000",
  28054=>"11111111",
  28055=>"00000000",
  28056=>"00000000",
  28057=>"00000000",
  28058=>"00000000",
  28059=>"00000001",
  28060=>"00000000",
  28061=>"00000000",
  28062=>"00000000",
  28063=>"00000000",
  28064=>"00000000",
  28065=>"00000000",
  28066=>"00000001",
  28067=>"00000000",
  28068=>"00000000",
  28069=>"00000000",
  28070=>"00000000",
  28071=>"00000000",
  28072=>"11111111",
  28073=>"00000000",
  28074=>"00000000",
  28075=>"00000000",
  28076=>"00000000",
  28077=>"00000000",
  28078=>"00000000",
  28079=>"00000000",
  28080=>"00000000",
  28081=>"00000000",
  28082=>"00000000",
  28083=>"00000001",
  28084=>"00000000",
  28085=>"00000000",
  28086=>"00000001",
  28087=>"00000000",
  28088=>"00000000",
  28089=>"00000000",
  28090=>"00000000",
  28091=>"00000000",
  28092=>"00000000",
  28093=>"11111111",
  28094=>"00000000",
  28095=>"00000000",
  28096=>"00000000",
  28097=>"00000000",
  28098=>"00000000",
  28099=>"00000000",
  28100=>"00000000",
  28101=>"00000000",
  28102=>"00000000",
  28103=>"00000000",
  28104=>"00000000",
  28105=>"00000000",
  28106=>"00000000",
  28107=>"00000000",
  28108=>"00000000",
  28109=>"00000000",
  28110=>"00000001",
  28111=>"00000000",
  28112=>"00000000",
  28113=>"00000001",
  28114=>"00000000",
  28115=>"00000000",
  28116=>"00000000",
  28117=>"00000000",
  28118=>"00000000",
  28119=>"00000000",
  28120=>"00000000",
  28121=>"00000000",
  28122=>"00000000",
  28123=>"00000000",
  28124=>"00000000",
  28125=>"11111111",
  28126=>"00000000",
  28127=>"00000000",
  28128=>"00000000",
  28129=>"00000000",
  28130=>"00000000",
  28131=>"11111111",
  28132=>"11111111",
  28133=>"00000000",
  28134=>"00000000",
  28135=>"00000000",
  28136=>"00000000",
  28137=>"00000000",
  28138=>"00000000",
  28139=>"00000000",
  28140=>"00000000",
  28141=>"00000000",
  28142=>"00000000",
  28143=>"00000000",
  28144=>"00000000",
  28145=>"00000001",
  28146=>"00000000",
  28147=>"00000000",
  28148=>"00000000",
  28149=>"00000000",
  28150=>"00000000",
  28151=>"00000001",
  28152=>"00000000",
  28153=>"00000000",
  28154=>"00000000",
  28155=>"00000000",
  28156=>"00000000",
  28157=>"00000001",
  28158=>"00000000",
  28159=>"00000000",
  28160=>"00000000",
  28161=>"00000000",
  28162=>"00000000",
  28163=>"11111111",
  28164=>"00000000",
  28165=>"00000001",
  28166=>"00000000",
  28167=>"00000000",
  28168=>"00000000",
  28169=>"00000000",
  28170=>"00000000",
  28171=>"00000001",
  28172=>"11111111",
  28173=>"00000001",
  28174=>"00000000",
  28175=>"00000000",
  28176=>"00000000",
  28177=>"00000000",
  28178=>"00000000",
  28179=>"00000000",
  28180=>"00000000",
  28181=>"11111111",
  28182=>"00000000",
  28183=>"00000000",
  28184=>"00000000",
  28185=>"00000000",
  28186=>"00000000",
  28187=>"00000000",
  28188=>"00000000",
  28189=>"00000000",
  28190=>"11111111",
  28191=>"00000000",
  28192=>"00000001",
  28193=>"00000000",
  28194=>"11111111",
  28195=>"00000000",
  28196=>"00000000",
  28197=>"00000000",
  28198=>"00000000",
  28199=>"00000001",
  28200=>"00000000",
  28201=>"00000000",
  28202=>"00000000",
  28203=>"00000000",
  28204=>"00000000",
  28205=>"00000000",
  28206=>"00000000",
  28207=>"00000000",
  28208=>"00000000",
  28209=>"00000000",
  28210=>"00000000",
  28211=>"00000000",
  28212=>"00000000",
  28213=>"00000000",
  28214=>"00000000",
  28215=>"00000000",
  28216=>"00000000",
  28217=>"00000000",
  28218=>"00000000",
  28219=>"00000000",
  28220=>"00000000",
  28221=>"00000000",
  28222=>"11111111",
  28223=>"00000000",
  28224=>"00000001",
  28225=>"00000000",
  28226=>"00000000",
  28227=>"11111111",
  28228=>"00000000",
  28229=>"00000000",
  28230=>"00000000",
  28231=>"00000000",
  28232=>"00000000",
  28233=>"00000000",
  28234=>"00000000",
  28235=>"00000000",
  28236=>"00000000",
  28237=>"00000000",
  28238=>"00000000",
  28239=>"00000000",
  28240=>"11111111",
  28241=>"00000000",
  28242=>"00000000",
  28243=>"00000000",
  28244=>"00000000",
  28245=>"11111111",
  28246=>"00000000",
  28247=>"00000000",
  28248=>"00000000",
  28249=>"00000000",
  28250=>"00000000",
  28251=>"00000000",
  28252=>"00000000",
  28253=>"00000000",
  28254=>"00000000",
  28255=>"00000000",
  28256=>"00000000",
  28257=>"11111111",
  28258=>"00000000",
  28259=>"00000000",
  28260=>"00000000",
  28261=>"00000000",
  28262=>"00000000",
  28263=>"00000000",
  28264=>"00000000",
  28265=>"00000001",
  28266=>"00000000",
  28267=>"00000000",
  28268=>"00000000",
  28269=>"00000000",
  28270=>"00000000",
  28271=>"00000000",
  28272=>"00000000",
  28273=>"00000000",
  28274=>"00000001",
  28275=>"00000000",
  28276=>"00000001",
  28277=>"00000000",
  28278=>"00000000",
  28279=>"00000000",
  28280=>"00000000",
  28281=>"11111111",
  28282=>"11111111",
  28283=>"00000001",
  28284=>"11111111",
  28285=>"11111110",
  28286=>"00000000",
  28287=>"00000000",
  28288=>"11111111",
  28289=>"00000000",
  28290=>"00000000",
  28291=>"00000000",
  28292=>"00000000",
  28293=>"00000000",
  28294=>"00000000",
  28295=>"11111111",
  28296=>"00000000",
  28297=>"00000001",
  28298=>"00000000",
  28299=>"00000000",
  28300=>"11111111",
  28301=>"00000000",
  28302=>"11111110",
  28303=>"00000000",
  28304=>"00000000",
  28305=>"00000000",
  28306=>"00000000",
  28307=>"00000001",
  28308=>"00000000",
  28309=>"00000000",
  28310=>"11111111",
  28311=>"00000000",
  28312=>"00000000",
  28313=>"00000000",
  28314=>"00000000",
  28315=>"00000000",
  28316=>"00000000",
  28317=>"00000000",
  28318=>"00000000",
  28319=>"00000000",
  28320=>"11111110",
  28321=>"00000000",
  28322=>"00000000",
  28323=>"00000001",
  28324=>"11111111",
  28325=>"11111111",
  28326=>"00000000",
  28327=>"00000000",
  28328=>"00000000",
  28329=>"00000000",
  28330=>"00000000",
  28331=>"00000001",
  28332=>"11111111",
  28333=>"00000000",
  28334=>"00000000",
  28335=>"00000001",
  28336=>"00000001",
  28337=>"00000000",
  28338=>"00000000",
  28339=>"00000000",
  28340=>"11111111",
  28341=>"00000000",
  28342=>"00000000",
  28343=>"00000000",
  28344=>"00000000",
  28345=>"00000000",
  28346=>"11111111",
  28347=>"00000000",
  28348=>"00000000",
  28349=>"00000001",
  28350=>"00000001",
  28351=>"00000000",
  28352=>"00000000",
  28353=>"00000001",
  28354=>"00000001",
  28355=>"00000000",
  28356=>"00000000",
  28357=>"00000001",
  28358=>"00000000",
  28359=>"11111111",
  28360=>"11111111",
  28361=>"00000000",
  28362=>"00000000",
  28363=>"00000000",
  28364=>"11111111",
  28365=>"00000000",
  28366=>"00000000",
  28367=>"00000000",
  28368=>"00000010",
  28369=>"00000000",
  28370=>"00000001",
  28371=>"00000000",
  28372=>"00000000",
  28373=>"00000000",
  28374=>"00000000",
  28375=>"00000000",
  28376=>"00000000",
  28377=>"00000001",
  28378=>"00000000",
  28379=>"00000000",
  28380=>"00000000",
  28381=>"00000000",
  28382=>"00000000",
  28383=>"00000000",
  28384=>"00000000",
  28385=>"00000000",
  28386=>"00000001",
  28387=>"00000000",
  28388=>"00000000",
  28389=>"00000000",
  28390=>"00000000",
  28391=>"00000000",
  28392=>"00000000",
  28393=>"00000000",
  28394=>"00000000",
  28395=>"00000000",
  28396=>"00000010",
  28397=>"00000000",
  28398=>"00000000",
  28399=>"00000000",
  28400=>"00000000",
  28401=>"00000000",
  28402=>"00000000",
  28403=>"00000001",
  28404=>"00000000",
  28405=>"00000000",
  28406=>"00000000",
  28407=>"00000000",
  28408=>"00000000",
  28409=>"00000000",
  28410=>"11111111",
  28411=>"00000000",
  28412=>"00000000",
  28413=>"00000000",
  28414=>"00000000",
  28415=>"11111111",
  28416=>"00000000",
  28417=>"00000000",
  28418=>"00000000",
  28419=>"00000000",
  28420=>"00000000",
  28421=>"00000000",
  28422=>"11111111",
  28423=>"11111111",
  28424=>"00000000",
  28425=>"00000000",
  28426=>"11111111",
  28427=>"00000000",
  28428=>"00000000",
  28429=>"00000000",
  28430=>"00000000",
  28431=>"00000001",
  28432=>"00000000",
  28433=>"00000000",
  28434=>"11111111",
  28435=>"00000000",
  28436=>"00000000",
  28437=>"00000001",
  28438=>"00000000",
  28439=>"00000000",
  28440=>"00000000",
  28441=>"00000000",
  28442=>"00000000",
  28443=>"00000000",
  28444=>"00000001",
  28445=>"00000000",
  28446=>"00000000",
  28447=>"00000000",
  28448=>"00000000",
  28449=>"00000000",
  28450=>"00000000",
  28451=>"00000000",
  28452=>"00000001",
  28453=>"00000000",
  28454=>"00000000",
  28455=>"00000001",
  28456=>"00000000",
  28457=>"00000000",
  28458=>"00000000",
  28459=>"11111111",
  28460=>"00000000",
  28461=>"00000000",
  28462=>"00000000",
  28463=>"00000000",
  28464=>"00000000",
  28465=>"00000000",
  28466=>"00000000",
  28467=>"00000000",
  28468=>"00000000",
  28469=>"00000000",
  28470=>"00000000",
  28471=>"00000000",
  28472=>"00000000",
  28473=>"00000001",
  28474=>"00000001",
  28475=>"00000000",
  28476=>"00000000",
  28477=>"11111111",
  28478=>"00000001",
  28479=>"00000001",
  28480=>"00000000",
  28481=>"00000000",
  28482=>"00000000",
  28483=>"00000000",
  28484=>"00000000",
  28485=>"00000000",
  28486=>"00000000",
  28487=>"11111111",
  28488=>"00000000",
  28489=>"00000000",
  28490=>"00000000",
  28491=>"00000001",
  28492=>"00000001",
  28493=>"00000000",
  28494=>"00000000",
  28495=>"00000000",
  28496=>"11111111",
  28497=>"11111111",
  28498=>"00000000",
  28499=>"00000000",
  28500=>"00000000",
  28501=>"00000000",
  28502=>"00000000",
  28503=>"00000000",
  28504=>"00000000",
  28505=>"00000000",
  28506=>"00000000",
  28507=>"00000000",
  28508=>"11111111",
  28509=>"00000000",
  28510=>"00000000",
  28511=>"00000000",
  28512=>"00000001",
  28513=>"00000000",
  28514=>"00000000",
  28515=>"00000000",
  28516=>"00000000",
  28517=>"00000000",
  28518=>"00000000",
  28519=>"00000000",
  28520=>"00000000",
  28521=>"00000000",
  28522=>"00000001",
  28523=>"00000000",
  28524=>"11111111",
  28525=>"00000000",
  28526=>"00000000",
  28527=>"00000000",
  28528=>"00000000",
  28529=>"00000000",
  28530=>"11111111",
  28531=>"00000000",
  28532=>"00000000",
  28533=>"00000000",
  28534=>"00000000",
  28535=>"00000001",
  28536=>"00000000",
  28537=>"11111111",
  28538=>"00000000",
  28539=>"11111111",
  28540=>"00000000",
  28541=>"00000001",
  28542=>"00000000",
  28543=>"00000000",
  28544=>"00000001",
  28545=>"00000000",
  28546=>"00000001",
  28547=>"00000000",
  28548=>"00000000",
  28549=>"00000000",
  28550=>"00000000",
  28551=>"00000000",
  28552=>"00000000",
  28553=>"00000000",
  28554=>"00000000",
  28555=>"00000001",
  28556=>"00000000",
  28557=>"00000000",
  28558=>"00000000",
  28559=>"00000000",
  28560=>"00000001",
  28561=>"00000000",
  28562=>"00000000",
  28563=>"11111110",
  28564=>"00000000",
  28565=>"00000000",
  28566=>"00000010",
  28567=>"00000000",
  28568=>"00000000",
  28569=>"00000000",
  28570=>"11111111",
  28571=>"00000000",
  28572=>"00000000",
  28573=>"00000000",
  28574=>"00000000",
  28575=>"00000000",
  28576=>"00000000",
  28577=>"00000000",
  28578=>"00000000",
  28579=>"00000000",
  28580=>"00000000",
  28581=>"00000000",
  28582=>"00000000",
  28583=>"00000000",
  28584=>"00000000",
  28585=>"00000000",
  28586=>"00000000",
  28587=>"00000000",
  28588=>"11111111",
  28589=>"00000001",
  28590=>"00000000",
  28591=>"00000000",
  28592=>"00000001",
  28593=>"00000000",
  28594=>"00000000",
  28595=>"11111111",
  28596=>"00000000",
  28597=>"00000000",
  28598=>"00000000",
  28599=>"00000000",
  28600=>"00000000",
  28601=>"00000000",
  28602=>"00000001",
  28603=>"00000000",
  28604=>"00000000",
  28605=>"00000000",
  28606=>"00000000",
  28607=>"00000000",
  28608=>"00000000",
  28609=>"11111111",
  28610=>"00000000",
  28611=>"11111111",
  28612=>"00000000",
  28613=>"00000000",
  28614=>"00000000",
  28615=>"00000001",
  28616=>"00000000",
  28617=>"00000000",
  28618=>"00000000",
  28619=>"00000000",
  28620=>"00000000",
  28621=>"00000000",
  28622=>"00000000",
  28623=>"00000000",
  28624=>"00000001",
  28625=>"00000000",
  28626=>"00000000",
  28627=>"11111111",
  28628=>"11111111",
  28629=>"00000000",
  28630=>"00000000",
  28631=>"00000000",
  28632=>"00000000",
  28633=>"00000000",
  28634=>"00000000",
  28635=>"00000000",
  28636=>"00000000",
  28637=>"00000001",
  28638=>"00000001",
  28639=>"00000000",
  28640=>"00000001",
  28641=>"00000000",
  28642=>"11111111",
  28643=>"00000000",
  28644=>"00000000",
  28645=>"00000000",
  28646=>"00000000",
  28647=>"00000001",
  28648=>"00000000",
  28649=>"00000000",
  28650=>"00000000",
  28651=>"11111111",
  28652=>"00000001",
  28653=>"00000000",
  28654=>"00000000",
  28655=>"00000000",
  28656=>"00000000",
  28657=>"00000000",
  28658=>"00000000",
  28659=>"11111111",
  28660=>"00000000",
  28661=>"00000001",
  28662=>"00000000",
  28663=>"00000000",
  28664=>"00000000",
  28665=>"00000000",
  28666=>"00000000",
  28667=>"11111111",
  28668=>"00000000",
  28669=>"00000000",
  28670=>"00000000",
  28671=>"00000000",
  28672=>"00000000",
  28673=>"00000000",
  28674=>"00000000",
  28675=>"00000000",
  28676=>"00000000",
  28677=>"00000000",
  28678=>"00000000",
  28679=>"00000000",
  28680=>"00000000",
  28681=>"00000000",
  28682=>"00000000",
  28683=>"00000000",
  28684=>"00000000",
  28685=>"00000001",
  28686=>"00000000",
  28687=>"00000000",
  28688=>"00000000",
  28689=>"00000000",
  28690=>"00000000",
  28691=>"00000000",
  28692=>"00000000",
  28693=>"00000001",
  28694=>"00000000",
  28695=>"00000000",
  28696=>"00000000",
  28697=>"00000000",
  28698=>"00000000",
  28699=>"00000001",
  28700=>"11111111",
  28701=>"00000000",
  28702=>"00000000",
  28703=>"00000000",
  28704=>"00000000",
  28705=>"00000000",
  28706=>"11111111",
  28707=>"00000000",
  28708=>"00000000",
  28709=>"00000000",
  28710=>"00000000",
  28711=>"00000000",
  28712=>"00000000",
  28713=>"00000000",
  28714=>"00000000",
  28715=>"00000000",
  28716=>"00000000",
  28717=>"00000000",
  28718=>"11111111",
  28719=>"11111111",
  28720=>"00000000",
  28721=>"00000001",
  28722=>"00000000",
  28723=>"11111111",
  28724=>"00000000",
  28725=>"00000000",
  28726=>"11111110",
  28727=>"00000000",
  28728=>"00000000",
  28729=>"00000000",
  28730=>"00000001",
  28731=>"00000000",
  28732=>"00000000",
  28733=>"00000000",
  28734=>"00000000",
  28735=>"00000000",
  28736=>"00000000",
  28737=>"00000000",
  28738=>"11111111",
  28739=>"00000000",
  28740=>"00000000",
  28741=>"00000001",
  28742=>"00000000",
  28743=>"00000000",
  28744=>"00000000",
  28745=>"00000000",
  28746=>"00000000",
  28747=>"11111110",
  28748=>"00000000",
  28749=>"00000000",
  28750=>"00000000",
  28751=>"11111111",
  28752=>"00000000",
  28753=>"00000000",
  28754=>"00000000",
  28755=>"00000000",
  28756=>"00000000",
  28757=>"00000000",
  28758=>"00000000",
  28759=>"00000001",
  28760=>"00000000",
  28761=>"00000000",
  28762=>"00000000",
  28763=>"00000000",
  28764=>"00000000",
  28765=>"00000000",
  28766=>"00000000",
  28767=>"00000000",
  28768=>"00000000",
  28769=>"00000000",
  28770=>"00000000",
  28771=>"00000000",
  28772=>"00000000",
  28773=>"00000000",
  28774=>"00000000",
  28775=>"00000000",
  28776=>"00000000",
  28777=>"00000000",
  28778=>"00000000",
  28779=>"00000000",
  28780=>"00000000",
  28781=>"00000000",
  28782=>"00000000",
  28783=>"00000000",
  28784=>"00000000",
  28785=>"00000000",
  28786=>"00000000",
  28787=>"00000000",
  28788=>"00000000",
  28789=>"00000000",
  28790=>"00000000",
  28791=>"00000000",
  28792=>"00000000",
  28793=>"00000000",
  28794=>"00000000",
  28795=>"00000000",
  28796=>"00000000",
  28797=>"00000000",
  28798=>"00000000",
  28799=>"00000000",
  28800=>"00000000",
  28801=>"00000000",
  28802=>"00000000",
  28803=>"00000000",
  28804=>"00000000",
  28805=>"00000001",
  28806=>"00000000",
  28807=>"00000000",
  28808=>"11111111",
  28809=>"11111111",
  28810=>"00000000",
  28811=>"00000000",
  28812=>"00000000",
  28813=>"00000000",
  28814=>"00000000",
  28815=>"00000000",
  28816=>"00000000",
  28817=>"00000000",
  28818=>"11111110",
  28819=>"00000000",
  28820=>"00000000",
  28821=>"00000000",
  28822=>"00000000",
  28823=>"00000000",
  28824=>"00000000",
  28825=>"00000000",
  28826=>"00000000",
  28827=>"00000000",
  28828=>"11111111",
  28829=>"00000000",
  28830=>"00000000",
  28831=>"00000000",
  28832=>"00000000",
  28833=>"00000000",
  28834=>"00000000",
  28835=>"00000000",
  28836=>"11111111",
  28837=>"00000000",
  28838=>"00000000",
  28839=>"00000000",
  28840=>"00000000",
  28841=>"00000000",
  28842=>"00000000",
  28843=>"00000000",
  28844=>"00000000",
  28845=>"00000000",
  28846=>"00000000",
  28847=>"00000000",
  28848=>"00000000",
  28849=>"00000000",
  28850=>"00000010",
  28851=>"00000000",
  28852=>"00000000",
  28853=>"00000000",
  28854=>"00000000",
  28855=>"00000000",
  28856=>"00000000",
  28857=>"00000000",
  28858=>"00000000",
  28859=>"00000000",
  28860=>"00000000",
  28861=>"11111100",
  28862=>"00000000",
  28863=>"11111111",
  28864=>"00000000",
  28865=>"11111111",
  28866=>"00000001",
  28867=>"00000000",
  28868=>"00000000",
  28869=>"00000000",
  28870=>"00000000",
  28871=>"00000000",
  28872=>"00000000",
  28873=>"00000001",
  28874=>"00000000",
  28875=>"00000000",
  28876=>"00000000",
  28877=>"00000000",
  28878=>"11111111",
  28879=>"00000000",
  28880=>"00000000",
  28881=>"00000000",
  28882=>"00000001",
  28883=>"00000000",
  28884=>"00000000",
  28885=>"00000000",
  28886=>"00000000",
  28887=>"00000000",
  28888=>"00000001",
  28889=>"00000000",
  28890=>"00000001",
  28891=>"00000000",
  28892=>"00000000",
  28893=>"00000000",
  28894=>"00000000",
  28895=>"00000000",
  28896=>"00000000",
  28897=>"00000000",
  28898=>"00000000",
  28899=>"00000000",
  28900=>"00000000",
  28901=>"00000000",
  28902=>"00000001",
  28903=>"00000000",
  28904=>"00000000",
  28905=>"00000000",
  28906=>"00000000",
  28907=>"11111111",
  28908=>"00000000",
  28909=>"00000000",
  28910=>"00000000",
  28911=>"00000010",
  28912=>"00000000",
  28913=>"00000000",
  28914=>"00000000",
  28915=>"00000000",
  28916=>"11111111",
  28917=>"00000000",
  28918=>"00000000",
  28919=>"00000000",
  28920=>"00000000",
  28921=>"00000000",
  28922=>"00000000",
  28923=>"00000000",
  28924=>"11111111",
  28925=>"00000000",
  28926=>"00000000",
  28927=>"00000000",
  28928=>"11111111",
  28929=>"00000000",
  28930=>"00000000",
  28931=>"00000001",
  28932=>"11111110",
  28933=>"00000000",
  28934=>"00000000",
  28935=>"00000000",
  28936=>"11111111",
  28937=>"00000001",
  28938=>"00000000",
  28939=>"00000000",
  28940=>"11111111",
  28941=>"00000000",
  28942=>"00000000",
  28943=>"00000000",
  28944=>"00000000",
  28945=>"00000000",
  28946=>"00000000",
  28947=>"00000000",
  28948=>"00000000",
  28949=>"00000001",
  28950=>"11111111",
  28951=>"11111111",
  28952=>"00000001",
  28953=>"00000000",
  28954=>"00000000",
  28955=>"00000000",
  28956=>"00000000",
  28957=>"00000000",
  28958=>"00000000",
  28959=>"00000000",
  28960=>"00000000",
  28961=>"00000000",
  28962=>"11111011",
  28963=>"00000000",
  28964=>"00000000",
  28965=>"00000000",
  28966=>"00000000",
  28967=>"00000000",
  28968=>"00000000",
  28969=>"00000000",
  28970=>"00000000",
  28971=>"00000000",
  28972=>"00000000",
  28973=>"00000010",
  28974=>"00000000",
  28975=>"00000000",
  28976=>"00000000",
  28977=>"00000000",
  28978=>"00000000",
  28979=>"00000000",
  28980=>"00000000",
  28981=>"00000000",
  28982=>"00000000",
  28983=>"00000000",
  28984=>"00000000",
  28985=>"00000000",
  28986=>"00000000",
  28987=>"00000011",
  28988=>"00000000",
  28989=>"11111111",
  28990=>"00000000",
  28991=>"00000001",
  28992=>"00000001",
  28993=>"00000000",
  28994=>"00000000",
  28995=>"00000000",
  28996=>"00000000",
  28997=>"00000000",
  28998=>"00000000",
  28999=>"00000001",
  29000=>"00000001",
  29001=>"00000000",
  29002=>"00000000",
  29003=>"11111111",
  29004=>"00000000",
  29005=>"11111111",
  29006=>"00000000",
  29007=>"00000000",
  29008=>"00000000",
  29009=>"00000000",
  29010=>"00000000",
  29011=>"00000000",
  29012=>"11111110",
  29013=>"00000000",
  29014=>"00000000",
  29015=>"00000000",
  29016=>"00000000",
  29017=>"00000000",
  29018=>"11111111",
  29019=>"00000000",
  29020=>"00000000",
  29021=>"11111110",
  29022=>"00000000",
  29023=>"00000000",
  29024=>"00000000",
  29025=>"00000000",
  29026=>"00000000",
  29027=>"00000000",
  29028=>"00000000",
  29029=>"00000000",
  29030=>"00000000",
  29031=>"00000000",
  29032=>"00000000",
  29033=>"00000000",
  29034=>"00000000",
  29035=>"00000000",
  29036=>"00000000",
  29037=>"00000000",
  29038=>"00000000",
  29039=>"00000000",
  29040=>"00000001",
  29041=>"00000000",
  29042=>"00000001",
  29043=>"00000000",
  29044=>"00000000",
  29045=>"00000000",
  29046=>"00000000",
  29047=>"00000000",
  29048=>"00000000",
  29049=>"00000000",
  29050=>"00000000",
  29051=>"00000000",
  29052=>"00000000",
  29053=>"00000000",
  29054=>"00000000",
  29055=>"00000000",
  29056=>"00000000",
  29057=>"11111111",
  29058=>"00000000",
  29059=>"00000000",
  29060=>"00000000",
  29061=>"11111111",
  29062=>"00000000",
  29063=>"00000000",
  29064=>"00000000",
  29065=>"00000001",
  29066=>"00000000",
  29067=>"00000000",
  29068=>"00000000",
  29069=>"11111111",
  29070=>"00000000",
  29071=>"00000000",
  29072=>"00000000",
  29073=>"00000000",
  29074=>"00000000",
  29075=>"00000000",
  29076=>"00000000",
  29077=>"11111111",
  29078=>"11111111",
  29079=>"00000000",
  29080=>"00000000",
  29081=>"00000001",
  29082=>"00000000",
  29083=>"11111111",
  29084=>"00000000",
  29085=>"00000000",
  29086=>"00000000",
  29087=>"00000000",
  29088=>"00000000",
  29089=>"00000000",
  29090=>"00000000",
  29091=>"00000000",
  29092=>"00000000",
  29093=>"00000000",
  29094=>"00000000",
  29095=>"00000000",
  29096=>"00000000",
  29097=>"00000000",
  29098=>"00000000",
  29099=>"00000000",
  29100=>"00000000",
  29101=>"00000000",
  29102=>"00000000",
  29103=>"00000000",
  29104=>"00000000",
  29105=>"00000000",
  29106=>"00000000",
  29107=>"00000000",
  29108=>"00000000",
  29109=>"00000000",
  29110=>"00000000",
  29111=>"00000000",
  29112=>"00000000",
  29113=>"00000000",
  29114=>"00000000",
  29115=>"00000000",
  29116=>"00000000",
  29117=>"00000001",
  29118=>"00000000",
  29119=>"00000000",
  29120=>"00000000",
  29121=>"00000000",
  29122=>"00000000",
  29123=>"00000000",
  29124=>"00000000",
  29125=>"00000000",
  29126=>"00000000",
  29127=>"00000000",
  29128=>"00000000",
  29129=>"00000000",
  29130=>"00000000",
  29131=>"00000000",
  29132=>"00000000",
  29133=>"00000001",
  29134=>"00000000",
  29135=>"00000000",
  29136=>"00000000",
  29137=>"00000000",
  29138=>"00000000",
  29139=>"00000000",
  29140=>"00000000",
  29141=>"11111111",
  29142=>"00000000",
  29143=>"00000000",
  29144=>"00000000",
  29145=>"00000000",
  29146=>"00000000",
  29147=>"00000000",
  29148=>"00000000",
  29149=>"00000001",
  29150=>"00000000",
  29151=>"00000000",
  29152=>"00000001",
  29153=>"00000000",
  29154=>"00000000",
  29155=>"00000000",
  29156=>"11111111",
  29157=>"00000000",
  29158=>"00000000",
  29159=>"00000001",
  29160=>"00000000",
  29161=>"00000000",
  29162=>"00000001",
  29163=>"00000000",
  29164=>"11111111",
  29165=>"00000000",
  29166=>"00000000",
  29167=>"00000000",
  29168=>"00000001",
  29169=>"00000000",
  29170=>"00000000",
  29171=>"00000000",
  29172=>"00000001",
  29173=>"00000000",
  29174=>"00000000",
  29175=>"00000000",
  29176=>"00000000",
  29177=>"00000001",
  29178=>"00000000",
  29179=>"11111111",
  29180=>"00000010",
  29181=>"00000000",
  29182=>"00000000",
  29183=>"11111110",
  29184=>"11111111",
  29185=>"00000000",
  29186=>"00000000",
  29187=>"00000000",
  29188=>"00000000",
  29189=>"00000000",
  29190=>"00000000",
  29191=>"11111111",
  29192=>"00000000",
  29193=>"00000000",
  29194=>"00000001",
  29195=>"11111111",
  29196=>"00000000",
  29197=>"00000001",
  29198=>"00000000",
  29199=>"00000000",
  29200=>"00000000",
  29201=>"00000000",
  29202=>"00000000",
  29203=>"00000000",
  29204=>"00000000",
  29205=>"00000000",
  29206=>"00000001",
  29207=>"00000000",
  29208=>"00000000",
  29209=>"00000000",
  29210=>"00000000",
  29211=>"00000000",
  29212=>"11111111",
  29213=>"00000000",
  29214=>"11111111",
  29215=>"00000000",
  29216=>"00000000",
  29217=>"00000000",
  29218=>"00000000",
  29219=>"00000000",
  29220=>"00000000",
  29221=>"00000000",
  29222=>"00000000",
  29223=>"00000000",
  29224=>"11111111",
  29225=>"00000001",
  29226=>"00000000",
  29227=>"00000000",
  29228=>"00000000",
  29229=>"00000000",
  29230=>"00000000",
  29231=>"00000000",
  29232=>"00000001",
  29233=>"00000000",
  29234=>"00000000",
  29235=>"00000001",
  29236=>"00000000",
  29237=>"00000000",
  29238=>"00000000",
  29239=>"00000000",
  29240=>"11111111",
  29241=>"00000000",
  29242=>"00000000",
  29243=>"00000001",
  29244=>"00000000",
  29245=>"00000001",
  29246=>"00000000",
  29247=>"00000000",
  29248=>"00000000",
  29249=>"00000000",
  29250=>"11111111",
  29251=>"00000000",
  29252=>"00000001",
  29253=>"00000010",
  29254=>"00000000",
  29255=>"00000000",
  29256=>"00000001",
  29257=>"00000000",
  29258=>"00000000",
  29259=>"00000000",
  29260=>"00000000",
  29261=>"00000000",
  29262=>"00000000",
  29263=>"00000000",
  29264=>"00000000",
  29265=>"00000000",
  29266=>"00000000",
  29267=>"00000000",
  29268=>"00000000",
  29269=>"00000000",
  29270=>"00000000",
  29271=>"00000000",
  29272=>"00000000",
  29273=>"00000000",
  29274=>"00000000",
  29275=>"00000000",
  29276=>"00000000",
  29277=>"00000000",
  29278=>"00000000",
  29279=>"00000000",
  29280=>"00000000",
  29281=>"00000000",
  29282=>"00000000",
  29283=>"00000000",
  29284=>"00000001",
  29285=>"00000001",
  29286=>"00000001",
  29287=>"00000000",
  29288=>"00000000",
  29289=>"00000000",
  29290=>"11111111",
  29291=>"00000000",
  29292=>"00000000",
  29293=>"00000000",
  29294=>"00000000",
  29295=>"00000000",
  29296=>"00000000",
  29297=>"00000000",
  29298=>"00000001",
  29299=>"00000000",
  29300=>"00000000",
  29301=>"00000000",
  29302=>"00000000",
  29303=>"00000000",
  29304=>"00000000",
  29305=>"00000000",
  29306=>"00000000",
  29307=>"00000000",
  29308=>"00000001",
  29309=>"00000000",
  29310=>"00000000",
  29311=>"00000000",
  29312=>"11111111",
  29313=>"00000000",
  29314=>"00000000",
  29315=>"00000000",
  29316=>"00000000",
  29317=>"00000000",
  29318=>"00000000",
  29319=>"00000000",
  29320=>"00000000",
  29321=>"00000000",
  29322=>"00000000",
  29323=>"00000000",
  29324=>"00000000",
  29325=>"11111111",
  29326=>"00000000",
  29327=>"00000000",
  29328=>"00000000",
  29329=>"00000000",
  29330=>"00000000",
  29331=>"11111110",
  29332=>"00000000",
  29333=>"00000000",
  29334=>"00000001",
  29335=>"00000000",
  29336=>"00000000",
  29337=>"00000000",
  29338=>"00000000",
  29339=>"00000000",
  29340=>"00000000",
  29341=>"00000000",
  29342=>"00000000",
  29343=>"00000000",
  29344=>"00000001",
  29345=>"00000000",
  29346=>"00000000",
  29347=>"00000000",
  29348=>"00000000",
  29349=>"11111111",
  29350=>"00000000",
  29351=>"00000000",
  29352=>"00000000",
  29353=>"00000000",
  29354=>"00000000",
  29355=>"00000000",
  29356=>"00000000",
  29357=>"00000000",
  29358=>"00000000",
  29359=>"00000000",
  29360=>"00000000",
  29361=>"00000000",
  29362=>"11111111",
  29363=>"00000000",
  29364=>"11111111",
  29365=>"00000000",
  29366=>"00000000",
  29367=>"00000000",
  29368=>"00000000",
  29369=>"00000001",
  29370=>"00000000",
  29371=>"00000000",
  29372=>"00000000",
  29373=>"00000000",
  29374=>"00000000",
  29375=>"00000000",
  29376=>"00000000",
  29377=>"00000000",
  29378=>"00000001",
  29379=>"00000000",
  29380=>"00000000",
  29381=>"00000000",
  29382=>"00000000",
  29383=>"00000000",
  29384=>"00000000",
  29385=>"00000000",
  29386=>"00000000",
  29387=>"00000000",
  29388=>"00000001",
  29389=>"00000000",
  29390=>"00000000",
  29391=>"00000000",
  29392=>"11111110",
  29393=>"00000000",
  29394=>"00000000",
  29395=>"00000000",
  29396=>"11111111",
  29397=>"00000000",
  29398=>"00000000",
  29399=>"00000000",
  29400=>"00000000",
  29401=>"00000001",
  29402=>"00000000",
  29403=>"00000000",
  29404=>"00000000",
  29405=>"00000000",
  29406=>"11111111",
  29407=>"00000000",
  29408=>"00000000",
  29409=>"00000000",
  29410=>"00000000",
  29411=>"00000000",
  29412=>"00000000",
  29413=>"00000000",
  29414=>"00000000",
  29415=>"00000000",
  29416=>"00000000",
  29417=>"00000000",
  29418=>"00000000",
  29419=>"00000000",
  29420=>"11111110",
  29421=>"00000000",
  29422=>"00000000",
  29423=>"00000000",
  29424=>"00000000",
  29425=>"00000000",
  29426=>"11111111",
  29427=>"00000000",
  29428=>"00000000",
  29429=>"00000000",
  29430=>"00000000",
  29431=>"00000000",
  29432=>"00000000",
  29433=>"00000000",
  29434=>"00000000",
  29435=>"00000000",
  29436=>"00000000",
  29437=>"11111111",
  29438=>"00000000",
  29439=>"00000000",
  29440=>"00000000",
  29441=>"11111111",
  29442=>"00000000",
  29443=>"11111111",
  29444=>"00000000",
  29445=>"00000011",
  29446=>"00000000",
  29447=>"11111111",
  29448=>"00000000",
  29449=>"00000000",
  29450=>"00000000",
  29451=>"11111111",
  29452=>"00000000",
  29453=>"00000000",
  29454=>"00000000",
  29455=>"11111111",
  29456=>"00000000",
  29457=>"11111111",
  29458=>"00000000",
  29459=>"00000000",
  29460=>"00000000",
  29461=>"00000000",
  29462=>"00000000",
  29463=>"00000000",
  29464=>"00000000",
  29465=>"00000000",
  29466=>"00000000",
  29467=>"00000000",
  29468=>"00000000",
  29469=>"00000000",
  29470=>"00000000",
  29471=>"00000000",
  29472=>"00000000",
  29473=>"00000000",
  29474=>"00000000",
  29475=>"11111111",
  29476=>"00000000",
  29477=>"00000000",
  29478=>"00000000",
  29479=>"00000000",
  29480=>"00000000",
  29481=>"00000000",
  29482=>"00000000",
  29483=>"00000000",
  29484=>"00000000",
  29485=>"00000000",
  29486=>"00000000",
  29487=>"00000000",
  29488=>"00000000",
  29489=>"00000000",
  29490=>"00000000",
  29491=>"00000000",
  29492=>"00000001",
  29493=>"11111111",
  29494=>"00000000",
  29495=>"00000000",
  29496=>"00000001",
  29497=>"11111110",
  29498=>"00000000",
  29499=>"00000000",
  29500=>"00000000",
  29501=>"00000000",
  29502=>"11111111",
  29503=>"00000000",
  29504=>"00000000",
  29505=>"00000000",
  29506=>"00000000",
  29507=>"00000000",
  29508=>"00000000",
  29509=>"00000000",
  29510=>"00000000",
  29511=>"00000000",
  29512=>"00000000",
  29513=>"00000000",
  29514=>"00000000",
  29515=>"00000000",
  29516=>"00000000",
  29517=>"11111111",
  29518=>"00000000",
  29519=>"00000000",
  29520=>"00000000",
  29521=>"00000000",
  29522=>"00000000",
  29523=>"00000000",
  29524=>"00000000",
  29525=>"00000000",
  29526=>"11111111",
  29527=>"00000000",
  29528=>"00000000",
  29529=>"00000000",
  29530=>"11111111",
  29531=>"00000000",
  29532=>"00000001",
  29533=>"00000000",
  29534=>"00000000",
  29535=>"00000000",
  29536=>"00000000",
  29537=>"00000000",
  29538=>"00000000",
  29539=>"00000000",
  29540=>"00000000",
  29541=>"00000000",
  29542=>"00000000",
  29543=>"00000000",
  29544=>"00000000",
  29545=>"00000000",
  29546=>"11111111",
  29547=>"00000000",
  29548=>"00000001",
  29549=>"00000000",
  29550=>"00000001",
  29551=>"00000000",
  29552=>"00000000",
  29553=>"00000000",
  29554=>"11111111",
  29555=>"00000000",
  29556=>"00000000",
  29557=>"00000000",
  29558=>"00000000",
  29559=>"11111111",
  29560=>"00000000",
  29561=>"00000001",
  29562=>"00000001",
  29563=>"00000000",
  29564=>"00000000",
  29565=>"11111111",
  29566=>"00000000",
  29567=>"00000000",
  29568=>"11111111",
  29569=>"00000000",
  29570=>"00000001",
  29571=>"00000000",
  29572=>"00000000",
  29573=>"00000001",
  29574=>"00000000",
  29575=>"00000000",
  29576=>"00000000",
  29577=>"00000001",
  29578=>"00000000",
  29579=>"00000000",
  29580=>"00000000",
  29581=>"00000000",
  29582=>"00000000",
  29583=>"11111111",
  29584=>"11111111",
  29585=>"00000000",
  29586=>"00000000",
  29587=>"00000001",
  29588=>"00000000",
  29589=>"00000000",
  29590=>"00000000",
  29591=>"00000000",
  29592=>"00000000",
  29593=>"00000000",
  29594=>"00000001",
  29595=>"00000000",
  29596=>"00000000",
  29597=>"00000000",
  29598=>"00000000",
  29599=>"11111111",
  29600=>"00000000",
  29601=>"11111110",
  29602=>"00000000",
  29603=>"00000000",
  29604=>"00000000",
  29605=>"00000000",
  29606=>"00000000",
  29607=>"00000000",
  29608=>"00000001",
  29609=>"00000001",
  29610=>"00000000",
  29611=>"00000001",
  29612=>"00000000",
  29613=>"00000000",
  29614=>"00000000",
  29615=>"00000000",
  29616=>"00000000",
  29617=>"00000000",
  29618=>"00000000",
  29619=>"00000000",
  29620=>"00000000",
  29621=>"00000000",
  29622=>"00000000",
  29623=>"00000001",
  29624=>"00000000",
  29625=>"00000000",
  29626=>"00000000",
  29627=>"00000000",
  29628=>"00000000",
  29629=>"00000000",
  29630=>"00000000",
  29631=>"00000000",
  29632=>"00000000",
  29633=>"00000000",
  29634=>"00000001",
  29635=>"00000000",
  29636=>"00000000",
  29637=>"00000000",
  29638=>"00000000",
  29639=>"11111111",
  29640=>"00000000",
  29641=>"00000001",
  29642=>"00000000",
  29643=>"00000000",
  29644=>"00000000",
  29645=>"00000000",
  29646=>"00000000",
  29647=>"00000000",
  29648=>"00000000",
  29649=>"00000000",
  29650=>"00000000",
  29651=>"00000000",
  29652=>"00000000",
  29653=>"00000000",
  29654=>"00000000",
  29655=>"00000000",
  29656=>"00000000",
  29657=>"00000000",
  29658=>"00000000",
  29659=>"00000000",
  29660=>"00000000",
  29661=>"00000000",
  29662=>"00000001",
  29663=>"00000000",
  29664=>"00000001",
  29665=>"00000000",
  29666=>"00000000",
  29667=>"00000000",
  29668=>"00000000",
  29669=>"00000000",
  29670=>"00000000",
  29671=>"00000000",
  29672=>"11111111",
  29673=>"00000000",
  29674=>"00000000",
  29675=>"00000000",
  29676=>"11111111",
  29677=>"00000000",
  29678=>"00000000",
  29679=>"00000000",
  29680=>"00000000",
  29681=>"00000000",
  29682=>"00000000",
  29683=>"00000000",
  29684=>"00000000",
  29685=>"00000000",
  29686=>"00000000",
  29687=>"00000000",
  29688=>"00000000",
  29689=>"00000000",
  29690=>"00000000",
  29691=>"00000000",
  29692=>"00000000",
  29693=>"00000000",
  29694=>"11111111",
  29695=>"00000000",
  29696=>"00000000",
  29697=>"11111101",
  29698=>"11111010",
  29699=>"11111100",
  29700=>"00000001",
  29701=>"00000001",
  29702=>"11111100",
  29703=>"00000001",
  29704=>"00000001",
  29705=>"11111111",
  29706=>"11111100",
  29707=>"11111011",
  29708=>"11111110",
  29709=>"11111111",
  29710=>"00000101",
  29711=>"00000000",
  29712=>"11111111",
  29713=>"00000101",
  29714=>"00000011",
  29715=>"00000010",
  29716=>"00000011",
  29717=>"11111000",
  29718=>"00000100",
  29719=>"11111111",
  29720=>"00000001",
  29721=>"11111111",
  29722=>"00000001",
  29723=>"00000000",
  29724=>"11111011",
  29725=>"00000011",
  29726=>"11111111",
  29727=>"00000000",
  29728=>"11111111",
  29729=>"11111111",
  29730=>"11111110",
  29731=>"11111110",
  29732=>"11111101",
  29733=>"11111101",
  29734=>"00000000",
  29735=>"11111001",
  29736=>"11111011",
  29737=>"00000001",
  29738=>"00000000",
  29739=>"11111111",
  29740=>"00000100",
  29741=>"11111011",
  29742=>"11111011",
  29743=>"11111111",
  29744=>"11111001",
  29745=>"11111011",
  29746=>"11111101",
  29747=>"11111010",
  29748=>"11111010",
  29749=>"00000001",
  29750=>"11111010",
  29751=>"00000001",
  29752=>"00000001",
  29753=>"00000000",
  29754=>"00000010",
  29755=>"00000010",
  29756=>"11111011",
  29757=>"11111000",
  29758=>"00000010",
  29759=>"11111110",
  29760=>"00000010",
  29761=>"11111000",
  29762=>"00000001",
  29763=>"11110010",
  29764=>"00000010",
  29765=>"11111100",
  29766=>"00000010",
  29767=>"00000110",
  29768=>"11111100",
  29769=>"00000011",
  29770=>"00000000",
  29771=>"11111001",
  29772=>"00000010",
  29773=>"00000000",
  29774=>"11111111",
  29775=>"11110111",
  29776=>"00000100",
  29777=>"11111111",
  29778=>"11111110",
  29779=>"11111101",
  29780=>"11111110",
  29781=>"00000000",
  29782=>"11111111",
  29783=>"11111001",
  29784=>"00000100",
  29785=>"00000010",
  29786=>"11111011",
  29787=>"11111110",
  29788=>"00000001",
  29789=>"00000010",
  29790=>"11111110",
  29791=>"11111111",
  29792=>"00000011",
  29793=>"11111110",
  29794=>"00000001",
  29795=>"00000000",
  29796=>"00000010",
  29797=>"11110111",
  29798=>"00000001",
  29799=>"00000010",
  29800=>"00000101",
  29801=>"00000010",
  29802=>"00000010",
  29803=>"00000010",
  29804=>"00000001",
  29805=>"00000000",
  29806=>"00000000",
  29807=>"00000001",
  29808=>"00000010",
  29809=>"11111010",
  29810=>"00000001",
  29811=>"11111110",
  29812=>"00000010",
  29813=>"00000000",
  29814=>"00000000",
  29815=>"00000000",
  29816=>"00000000",
  29817=>"00000000",
  29818=>"00000011",
  29819=>"11111111",
  29820=>"00000010",
  29821=>"11111111",
  29822=>"11111010",
  29823=>"11111111",
  29824=>"11111110",
  29825=>"00000010",
  29826=>"00000000",
  29827=>"00000000",
  29828=>"00000001",
  29829=>"00000001",
  29830=>"11111001",
  29831=>"11111111",
  29832=>"00000101",
  29833=>"11111101",
  29834=>"11111110",
  29835=>"00000000",
  29836=>"00000011",
  29837=>"11111110",
  29838=>"11111100",
  29839=>"11111111",
  29840=>"11111110",
  29841=>"00000001",
  29842=>"11111100",
  29843=>"11111100",
  29844=>"11111111",
  29845=>"00000001",
  29846=>"00000001",
  29847=>"11111010",
  29848=>"00000000",
  29849=>"00000001",
  29850=>"00000010",
  29851=>"00000000",
  29852=>"11111000",
  29853=>"11111110",
  29854=>"11110101",
  29855=>"00000011",
  29856=>"00000011",
  29857=>"11111110",
  29858=>"00000000",
  29859=>"00000001",
  29860=>"11111010",
  29861=>"00000010",
  29862=>"00000000",
  29863=>"11111001",
  29864=>"00000001",
  29865=>"11111110",
  29866=>"00000000",
  29867=>"00000000",
  29868=>"00000010",
  29869=>"00000001",
  29870=>"00000011",
  29871=>"00000100",
  29872=>"00000001",
  29873=>"11111010",
  29874=>"00001000",
  29875=>"11111111",
  29876=>"00000000",
  29877=>"00000011",
  29878=>"11111111",
  29879=>"00000000",
  29880=>"00000000",
  29881=>"00000001",
  29882=>"11111101",
  29883=>"00000000",
  29884=>"11111111",
  29885=>"11111000",
  29886=>"11111110",
  29887=>"11111111",
  29888=>"11111011",
  29889=>"00000000",
  29890=>"11111000",
  29891=>"00000001",
  29892=>"11111111",
  29893=>"00000010",
  29894=>"00000000",
  29895=>"11111011",
  29896=>"11111011",
  29897=>"00000010",
  29898=>"00000010",
  29899=>"11111111",
  29900=>"00000001",
  29901=>"11111111",
  29902=>"11111101",
  29903=>"11111110",
  29904=>"11111111",
  29905=>"00000000",
  29906=>"11111100",
  29907=>"11111011",
  29908=>"11111001",
  29909=>"00000001",
  29910=>"11110101",
  29911=>"00000001",
  29912=>"11111010",
  29913=>"11111011",
  29914=>"11111010",
  29915=>"00000010",
  29916=>"11111101",
  29917=>"00000010",
  29918=>"11111111",
  29919=>"00000000",
  29920=>"11111101",
  29921=>"00000001",
  29922=>"11111111",
  29923=>"00000001",
  29924=>"11111111",
  29925=>"00000001",
  29926=>"11111110",
  29927=>"00000000",
  29928=>"11111001",
  29929=>"11111111",
  29930=>"11111100",
  29931=>"11111101",
  29932=>"11110110",
  29933=>"11111111",
  29934=>"00000101",
  29935=>"11111011",
  29936=>"00000001",
  29937=>"00000010",
  29938=>"00000010",
  29939=>"00000001",
  29940=>"11111101",
  29941=>"00000000",
  29942=>"11111011",
  29943=>"11111101",
  29944=>"11111101",
  29945=>"00000001",
  29946=>"00000001",
  29947=>"11111001",
  29948=>"11111100",
  29949=>"00000001",
  29950=>"11111011",
  29951=>"00000000",
  29952=>"11111000",
  29953=>"11111111",
  29954=>"00000000",
  29955=>"00000110",
  29956=>"11110111",
  29957=>"00000011",
  29958=>"11111111",
  29959=>"11111111",
  29960=>"11111011",
  29961=>"00000001",
  29962=>"00000010",
  29963=>"11111110",
  29964=>"11111001",
  29965=>"00000011",
  29966=>"00000001",
  29967=>"00000010",
  29968=>"11111111",
  29969=>"00000000",
  29970=>"00000001",
  29971=>"00000000",
  29972=>"00000010",
  29973=>"00000011",
  29974=>"00000100",
  29975=>"00000010",
  29976=>"00000011",
  29977=>"11111111",
  29978=>"11111000",
  29979=>"11111011",
  29980=>"11111110",
  29981=>"11111011",
  29982=>"11111101",
  29983=>"00000000",
  29984=>"00000000",
  29985=>"00000011",
  29986=>"11111111",
  29987=>"00000000",
  29988=>"00000001",
  29989=>"00000010",
  29990=>"11111110",
  29991=>"11111111",
  29992=>"00000010",
  29993=>"11111101",
  29994=>"11111111",
  29995=>"00000000",
  29996=>"00000001",
  29997=>"11111000",
  29998=>"11111101",
  29999=>"11111110",
  30000=>"00000000",
  30001=>"11111000",
  30002=>"00000010",
  30003=>"00000010",
  30004=>"00000000",
  30005=>"11111111",
  30006=>"11111111",
  30007=>"11111110",
  30008=>"11111111",
  30009=>"11111111",
  30010=>"11111101",
  30011=>"00001001",
  30012=>"11111110",
  30013=>"00000000",
  30014=>"11111110",
  30015=>"11111010",
  30016=>"11110111",
  30017=>"11111111",
  30018=>"11110111",
  30019=>"00000000",
  30020=>"11111011",
  30021=>"11111110",
  30022=>"11111111",
  30023=>"11111110",
  30024=>"11111111",
  30025=>"00000000",
  30026=>"11111110",
  30027=>"11111011",
  30028=>"00000010",
  30029=>"00000001",
  30030=>"11111111",
  30031=>"00000010",
  30032=>"00000001",
  30033=>"11111110",
  30034=>"11111111",
  30035=>"11111101",
  30036=>"00000001",
  30037=>"00000010",
  30038=>"00000001",
  30039=>"11111111",
  30040=>"11111110",
  30041=>"00000100",
  30042=>"11110111",
  30043=>"00000001",
  30044=>"11111100",
  30045=>"11110110",
  30046=>"00000011",
  30047=>"00000000",
  30048=>"00000000",
  30049=>"00000001",
  30050=>"11111001",
  30051=>"00000000",
  30052=>"11111001",
  30053=>"00000000",
  30054=>"11110111",
  30055=>"11111110",
  30056=>"00000000",
  30057=>"11111101",
  30058=>"11111110",
  30059=>"00000001",
  30060=>"00000011",
  30061=>"00000000",
  30062=>"11111111",
  30063=>"11111111",
  30064=>"11111001",
  30065=>"00000011",
  30066=>"00000101",
  30067=>"00000001",
  30068=>"00000001",
  30069=>"00000001",
  30070=>"11111101",
  30071=>"11110101",
  30072=>"00000010",
  30073=>"11111111",
  30074=>"00000010",
  30075=>"11111101",
  30076=>"11111110",
  30077=>"11111111",
  30078=>"00000000",
  30079=>"00000000",
  30080=>"00000000",
  30081=>"11111111",
  30082=>"11111110",
  30083=>"00000001",
  30084=>"11111010",
  30085=>"00000001",
  30086=>"11111100",
  30087=>"00000000",
  30088=>"11111011",
  30089=>"00000001",
  30090=>"00000000",
  30091=>"11111001",
  30092=>"11111111",
  30093=>"00000011",
  30094=>"11111111",
  30095=>"00000000",
  30096=>"11111010",
  30097=>"00000000",
  30098=>"00000001",
  30099=>"11111001",
  30100=>"00000000",
  30101=>"00000100",
  30102=>"11111011",
  30103=>"00000000",
  30104=>"11111101",
  30105=>"00000010",
  30106=>"11111101",
  30107=>"00000101",
  30108=>"00000000",
  30109=>"00000010",
  30110=>"00000000",
  30111=>"11111111",
  30112=>"00000000",
  30113=>"11111101",
  30114=>"00000011",
  30115=>"00000001",
  30116=>"11111100",
  30117=>"00000010",
  30118=>"11111111",
  30119=>"11111110",
  30120=>"00000001",
  30121=>"00000011",
  30122=>"11111100",
  30123=>"11111011",
  30124=>"11111111",
  30125=>"00000010",
  30126=>"00000000",
  30127=>"00000010",
  30128=>"11111111",
  30129=>"11111111",
  30130=>"11111101",
  30131=>"00000010",
  30132=>"11111110",
  30133=>"11111111",
  30134=>"11111101",
  30135=>"11111111",
  30136=>"11111110",
  30137=>"11111111",
  30138=>"00000000",
  30139=>"00000010",
  30140=>"11111011",
  30141=>"00000000",
  30142=>"00000000",
  30143=>"11111000",
  30144=>"00000001",
  30145=>"00000010",
  30146=>"00000001",
  30147=>"00000011",
  30148=>"00000001",
  30149=>"11111111",
  30150=>"00000000",
  30151=>"11111110",
  30152=>"00000001",
  30153=>"11111110",
  30154=>"11111110",
  30155=>"11111111",
  30156=>"11111111",
  30157=>"11110111",
  30158=>"11111111",
  30159=>"11111100",
  30160=>"11111100",
  30161=>"11111100",
  30162=>"00000001",
  30163=>"00000011",
  30164=>"00000000",
  30165=>"00000011",
  30166=>"00000000",
  30167=>"00000010",
  30168=>"11111010",
  30169=>"00000000",
  30170=>"11111110",
  30171=>"11111110",
  30172=>"00000001",
  30173=>"11111111",
  30174=>"11111111",
  30175=>"11111111",
  30176=>"00000010",
  30177=>"00000001",
  30178=>"00000000",
  30179=>"11111010",
  30180=>"11111001",
  30181=>"00000000",
  30182=>"11111111",
  30183=>"11111010",
  30184=>"00000001",
  30185=>"00000001",
  30186=>"00000001",
  30187=>"00000011",
  30188=>"11110111",
  30189=>"11111111",
  30190=>"00000101",
  30191=>"00000010",
  30192=>"11111101",
  30193=>"00000000",
  30194=>"11111011",
  30195=>"00000000",
  30196=>"11111011",
  30197=>"00000100",
  30198=>"11111100",
  30199=>"11111110",
  30200=>"00000110",
  30201=>"00000001",
  30202=>"11111110",
  30203=>"11111111",
  30204=>"11111110",
  30205=>"00000010",
  30206=>"00000001",
  30207=>"00000100",
  30208=>"11111011",
  30209=>"11111110",
  30210=>"00000010",
  30211=>"00000001",
  30212=>"11111111",
  30213=>"11110111",
  30214=>"00000010",
  30215=>"11111001",
  30216=>"11110111",
  30217=>"00000011",
  30218=>"11111110",
  30219=>"11111010",
  30220=>"00000010",
  30221=>"11111011",
  30222=>"00000000",
  30223=>"00000001",
  30224=>"00000000",
  30225=>"00000010",
  30226=>"00000001",
  30227=>"11111111",
  30228=>"00000001",
  30229=>"11110110",
  30230=>"11111110",
  30231=>"00000001",
  30232=>"00000000",
  30233=>"00000000",
  30234=>"11111110",
  30235=>"11110110",
  30236=>"00000011",
  30237=>"00000010",
  30238=>"00000000",
  30239=>"11111110",
  30240=>"11111110",
  30241=>"00000000",
  30242=>"00000000",
  30243=>"11111110",
  30244=>"00000000",
  30245=>"11111111",
  30246=>"11111011",
  30247=>"00000010",
  30248=>"00000010",
  30249=>"11111000",
  30250=>"00000001",
  30251=>"00000000",
  30252=>"00000000",
  30253=>"11111111",
  30254=>"11111110",
  30255=>"11111110",
  30256=>"11111111",
  30257=>"11111101",
  30258=>"11111001",
  30259=>"00000100",
  30260=>"11111101",
  30261=>"11111111",
  30262=>"00000000",
  30263=>"00000001",
  30264=>"00000000",
  30265=>"00000000",
  30266=>"11111001",
  30267=>"00000011",
  30268=>"00000010",
  30269=>"00000011",
  30270=>"11111100",
  30271=>"11111110",
  30272=>"11111110",
  30273=>"11111111",
  30274=>"00000110",
  30275=>"00001000",
  30276=>"00000101",
  30277=>"11111110",
  30278=>"11111110",
  30279=>"00000010",
  30280=>"11111111",
  30281=>"11111010",
  30282=>"00000000",
  30283=>"00000001",
  30284=>"11111110",
  30285=>"00000000",
  30286=>"00000100",
  30287=>"11111111",
  30288=>"11111101",
  30289=>"00000011",
  30290=>"00000000",
  30291=>"11111100",
  30292=>"00000100",
  30293=>"11111110",
  30294=>"11111101",
  30295=>"11111100",
  30296=>"00000000",
  30297=>"11111101",
  30298=>"11110111",
  30299=>"11111011",
  30300=>"00000001",
  30301=>"11111000",
  30302=>"11111111",
  30303=>"11110110",
  30304=>"00000000",
  30305=>"00000000",
  30306=>"11111110",
  30307=>"00000001",
  30308=>"00000010",
  30309=>"11111000",
  30310=>"11110111",
  30311=>"11111011",
  30312=>"11111111",
  30313=>"00000100",
  30314=>"11111000",
  30315=>"00000000",
  30316=>"00000001",
  30317=>"00000010",
  30318=>"11111111",
  30319=>"00000010",
  30320=>"00000011",
  30321=>"11111001",
  30322=>"11111000",
  30323=>"11111111",
  30324=>"11111010",
  30325=>"11111101",
  30326=>"11111111",
  30327=>"00000000",
  30328=>"00000000",
  30329=>"11111111",
  30330=>"00000000",
  30331=>"11111101",
  30332=>"00000000",
  30333=>"11111111",
  30334=>"00000000",
  30335=>"11111100",
  30336=>"11110111",
  30337=>"11111110",
  30338=>"11111110",
  30339=>"11111101",
  30340=>"00000000",
  30341=>"00000010",
  30342=>"11111111",
  30343=>"00000001",
  30344=>"00000010",
  30345=>"11111010",
  30346=>"00000001",
  30347=>"11111111",
  30348=>"11111001",
  30349=>"11111011",
  30350=>"11111100",
  30351=>"00000001",
  30352=>"11111110",
  30353=>"00000000",
  30354=>"11111110",
  30355=>"11111000",
  30356=>"00000001",
  30357=>"00000101",
  30358=>"11111010",
  30359=>"00000010",
  30360=>"11111011",
  30361=>"00000001",
  30362=>"11111111",
  30363=>"00000000",
  30364=>"11111111",
  30365=>"00000001",
  30366=>"00000100",
  30367=>"11111111",
  30368=>"11111011",
  30369=>"00000001",
  30370=>"11111101",
  30371=>"00000001",
  30372=>"11111111",
  30373=>"00000000",
  30374=>"00000001",
  30375=>"11111110",
  30376=>"11111111",
  30377=>"11111110",
  30378=>"00000000",
  30379=>"11111011",
  30380=>"11111111",
  30381=>"00000001",
  30382=>"11111101",
  30383=>"00000010",
  30384=>"11111000",
  30385=>"00000000",
  30386=>"00000011",
  30387=>"11111110",
  30388=>"11111010",
  30389=>"00000001",
  30390=>"11111110",
  30391=>"11111111",
  30392=>"11111111",
  30393=>"11111001",
  30394=>"11111010",
  30395=>"11111110",
  30396=>"00000010",
  30397=>"11111010",
  30398=>"00000000",
  30399=>"11111000",
  30400=>"00000001",
  30401=>"00000001",
  30402=>"11111011",
  30403=>"11111111",
  30404=>"00000000",
  30405=>"00000000",
  30406=>"11111111",
  30407=>"00000010",
  30408=>"11111011",
  30409=>"00000000",
  30410=>"11111111",
  30411=>"00000000",
  30412=>"11111111",
  30413=>"00000010",
  30414=>"11111001",
  30415=>"11111110",
  30416=>"11111010",
  30417=>"11111111",
  30418=>"00000001",
  30419=>"00000001",
  30420=>"11111011",
  30421=>"11111110",
  30422=>"11111001",
  30423=>"11111100",
  30424=>"11111111",
  30425=>"11111011",
  30426=>"11111010",
  30427=>"11111110",
  30428=>"00000000",
  30429=>"00000000",
  30430=>"00000010",
  30431=>"11111110",
  30432=>"00000001",
  30433=>"00000001",
  30434=>"11111100",
  30435=>"11111101",
  30436=>"11111111",
  30437=>"00000010",
  30438=>"00000010",
  30439=>"11111100",
  30440=>"11111000",
  30441=>"11111111",
  30442=>"00000011",
  30443=>"11111101",
  30444=>"00000001",
  30445=>"11111101",
  30446=>"00000001",
  30447=>"00000000",
  30448=>"00000000",
  30449=>"11111011",
  30450=>"00000000",
  30451=>"11111111",
  30452=>"00000001",
  30453=>"11111111",
  30454=>"11111101",
  30455=>"00000000",
  30456=>"11111110",
  30457=>"00000000",
  30458=>"11111110",
  30459=>"00000010",
  30460=>"11111111",
  30461=>"00000010",
  30462=>"00000010",
  30463=>"11111100",
  30464=>"00000001",
  30465=>"00001000",
  30466=>"11111110",
  30467=>"00000001",
  30468=>"00000000",
  30469=>"11111010",
  30470=>"11111111",
  30471=>"00000010",
  30472=>"00000000",
  30473=>"00000001",
  30474=>"11111001",
  30475=>"11111111",
  30476=>"11111111",
  30477=>"00000000",
  30478=>"11111110",
  30479=>"11111110",
  30480=>"00000001",
  30481=>"00000001",
  30482=>"00000001",
  30483=>"11111110",
  30484=>"11111111",
  30485=>"11111110",
  30486=>"00000001",
  30487=>"11111110",
  30488=>"00000010",
  30489=>"00000001",
  30490=>"11111111",
  30491=>"00000000",
  30492=>"00000010",
  30493=>"00000010",
  30494=>"00000001",
  30495=>"11111101",
  30496=>"00000000",
  30497=>"00000010",
  30498=>"11111010",
  30499=>"11111110",
  30500=>"00000011",
  30501=>"00000001",
  30502=>"11111111",
  30503=>"00000001",
  30504=>"00000001",
  30505=>"00000000",
  30506=>"11111101",
  30507=>"00000001",
  30508=>"11111000",
  30509=>"11111111",
  30510=>"11111101",
  30511=>"00000100",
  30512=>"11111101",
  30513=>"00000011",
  30514=>"11111111",
  30515=>"00000000",
  30516=>"11111000",
  30517=>"00000001",
  30518=>"11111100",
  30519=>"11111001",
  30520=>"00000010",
  30521=>"11111000",
  30522=>"00000001",
  30523=>"00000000",
  30524=>"00000001",
  30525=>"11111010",
  30526=>"11111111",
  30527=>"00000100",
  30528=>"00000010",
  30529=>"00000001",
  30530=>"00000001",
  30531=>"00000001",
  30532=>"00000011",
  30533=>"11111100",
  30534=>"00000001",
  30535=>"11111111",
  30536=>"00000010",
  30537=>"00000000",
  30538=>"00000000",
  30539=>"00000001",
  30540=>"11111001",
  30541=>"11111001",
  30542=>"00000000",
  30543=>"11111100",
  30544=>"11111001",
  30545=>"11111010",
  30546=>"00000001",
  30547=>"11111101",
  30548=>"11111100",
  30549=>"11111001",
  30550=>"11111011",
  30551=>"00000001",
  30552=>"11111111",
  30553=>"00000001",
  30554=>"11110101",
  30555=>"11111110",
  30556=>"00000010",
  30557=>"00000001",
  30558=>"00000000",
  30559=>"00000000",
  30560=>"00000010",
  30561=>"00000000",
  30562=>"00000010",
  30563=>"00000000",
  30564=>"11111001",
  30565=>"11111100",
  30566=>"11111011",
  30567=>"00000000",
  30568=>"00000000",
  30569=>"00000100",
  30570=>"11111110",
  30571=>"00000010",
  30572=>"00000000",
  30573=>"11111100",
  30574=>"00000100",
  30575=>"11111110",
  30576=>"11111001",
  30577=>"00000000",
  30578=>"11111000",
  30579=>"00000000",
  30580=>"11111111",
  30581=>"00000001",
  30582=>"00000001",
  30583=>"11111011",
  30584=>"11111111",
  30585=>"00000100",
  30586=>"11111110",
  30587=>"00000001",
  30588=>"00000001",
  30589=>"11111101",
  30590=>"00000000",
  30591=>"11111100",
  30592=>"11111101",
  30593=>"00000010",
  30594=>"11110111",
  30595=>"00000000",
  30596=>"00000001",
  30597=>"11111010",
  30598=>"00000000",
  30599=>"00000000",
  30600=>"11111110",
  30601=>"00000010",
  30602=>"11111100",
  30603=>"00000001",
  30604=>"00000010",
  30605=>"11111101",
  30606=>"00000000",
  30607=>"11110111",
  30608=>"11111011",
  30609=>"00000000",
  30610=>"11111111",
  30611=>"11111000",
  30612=>"11111111",
  30613=>"11111111",
  30614=>"11111011",
  30615=>"11111101",
  30616=>"11111110",
  30617=>"11111110",
  30618=>"00000001",
  30619=>"00000010",
  30620=>"00000000",
  30621=>"11111111",
  30622=>"00000100",
  30623=>"11111101",
  30624=>"00000010",
  30625=>"11111000",
  30626=>"00000010",
  30627=>"11111001",
  30628=>"11111101",
  30629=>"11111111",
  30630=>"00000011",
  30631=>"00000001",
  30632=>"11110111",
  30633=>"11111110",
  30634=>"00000011",
  30635=>"11111001",
  30636=>"00000001",
  30637=>"11111010",
  30638=>"11111101",
  30639=>"11111001",
  30640=>"00000111",
  30641=>"11111101",
  30642=>"00000000",
  30643=>"11111111",
  30644=>"11111010",
  30645=>"11111111",
  30646=>"00000000",
  30647=>"00000000",
  30648=>"00000001",
  30649=>"11111000",
  30650=>"11111111",
  30651=>"00000000",
  30652=>"00000000",
  30653=>"00000001",
  30654=>"11111010",
  30655=>"11111010",
  30656=>"11111110",
  30657=>"00000011",
  30658=>"00000000",
  30659=>"11111111",
  30660=>"11111110",
  30661=>"11111110",
  30662=>"11111110",
  30663=>"11111011",
  30664=>"00000010",
  30665=>"00000000",
  30666=>"00000010",
  30667=>"00000001",
  30668=>"00000001",
  30669=>"00000000",
  30670=>"00000000",
  30671=>"00000000",
  30672=>"11111011",
  30673=>"11111110",
  30674=>"00000000",
  30675=>"00000000",
  30676=>"11111100",
  30677=>"00000011",
  30678=>"00000000",
  30679=>"00000001",
  30680=>"11111000",
  30681=>"00000000",
  30682=>"00000101",
  30683=>"00000001",
  30684=>"11111110",
  30685=>"00000010",
  30686=>"11111100",
  30687=>"00000001",
  30688=>"00000110",
  30689=>"11111110",
  30690=>"11111101",
  30691=>"11111001",
  30692=>"11111011",
  30693=>"11111101",
  30694=>"00000000",
  30695=>"00000010",
  30696=>"11111110",
  30697=>"11111010",
  30698=>"00000100",
  30699=>"00000000",
  30700=>"00000011",
  30701=>"11111111",
  30702=>"11111101",
  30703=>"11111101",
  30704=>"11111111",
  30705=>"11111110",
  30706=>"11111111",
  30707=>"00000111",
  30708=>"00000000",
  30709=>"00000111",
  30710=>"00000011",
  30711=>"11111110",
  30712=>"00000000",
  30713=>"00000000",
  30714=>"11111111",
  30715=>"11111110",
  30716=>"11111110",
  30717=>"11111110",
  30718=>"00000000",
  30719=>"00000001",
  30720=>"00000001",
  30721=>"11111111",
  30722=>"00000001",
  30723=>"00000010",
  30724=>"11111100",
  30725=>"00000000",
  30726=>"00000001",
  30727=>"11111111",
  30728=>"00000001",
  30729=>"11111110",
  30730=>"00000010",
  30731=>"00000001",
  30732=>"00000100",
  30733=>"00000010",
  30734=>"00000011",
  30735=>"00000000",
  30736=>"11111111",
  30737=>"00000000",
  30738=>"00000001",
  30739=>"00000001",
  30740=>"11111111",
  30741=>"00000010",
  30742=>"11111100",
  30743=>"11111110",
  30744=>"11111111",
  30745=>"11111110",
  30746=>"11111110",
  30747=>"00000001",
  30748=>"11111111",
  30749=>"11111110",
  30750=>"11111111",
  30751=>"11111111",
  30752=>"00000001",
  30753=>"11111101",
  30754=>"11111101",
  30755=>"00000001",
  30756=>"00000010",
  30757=>"00000011",
  30758=>"11111111",
  30759=>"00000000",
  30760=>"11111110",
  30761=>"11111101",
  30762=>"11111110",
  30763=>"11111110",
  30764=>"11111101",
  30765=>"00000010",
  30766=>"00000010",
  30767=>"00000010",
  30768=>"00000000",
  30769=>"00000000",
  30770=>"11111101",
  30771=>"00000001",
  30772=>"11111110",
  30773=>"11111101",
  30774=>"11111101",
  30775=>"00000000",
  30776=>"11111110",
  30777=>"11111110",
  30778=>"11111110",
  30779=>"00000100",
  30780=>"00000000",
  30781=>"00000011",
  30782=>"11111110",
  30783=>"11111110",
  30784=>"11111101",
  30785=>"11111110",
  30786=>"11111101",
  30787=>"00000010",
  30788=>"11111101",
  30789=>"11111110",
  30790=>"11111110",
  30791=>"11111101",
  30792=>"11111111",
  30793=>"11111111",
  30794=>"11111110",
  30795=>"00000000",
  30796=>"11111110",
  30797=>"11111111",
  30798=>"00000011",
  30799=>"00000001",
  30800=>"00000001",
  30801=>"00000010",
  30802=>"11111111",
  30803=>"00000000",
  30804=>"11111101",
  30805=>"00000001",
  30806=>"11111101",
  30807=>"00000000",
  30808=>"00000110",
  30809=>"11111101",
  30810=>"11111111",
  30811=>"11111111",
  30812=>"00000000",
  30813=>"00000001",
  30814=>"00000000",
  30815=>"00000000",
  30816=>"00000011",
  30817=>"00000000",
  30818=>"11111101",
  30819=>"00000100",
  30820=>"00000110",
  30821=>"11111111",
  30822=>"11111110",
  30823=>"11111111",
  30824=>"00000010",
  30825=>"00000010",
  30826=>"00000010",
  30827=>"11111101",
  30828=>"00000010",
  30829=>"00000000",
  30830=>"00000001",
  30831=>"00000010",
  30832=>"00000001",
  30833=>"00000000",
  30834=>"11111101",
  30835=>"00000000",
  30836=>"11111101",
  30837=>"11111110",
  30838=>"11111101",
  30839=>"00000101",
  30840=>"00000000",
  30841=>"11111110",
  30842=>"11111111",
  30843=>"00000010",
  30844=>"00000011",
  30845=>"11111110",
  30846=>"00000011",
  30847=>"00000001",
  30848=>"00000000",
  30849=>"11111101",
  30850=>"00000001",
  30851=>"00000000",
  30852=>"00000001",
  30853=>"00000010",
  30854=>"11111110",
  30855=>"11111110",
  30856=>"11111111",
  30857=>"00000010",
  30858=>"11111111",
  30859=>"11111101",
  30860=>"11111111",
  30861=>"11111110",
  30862=>"00000000",
  30863=>"11111101",
  30864=>"00000001",
  30865=>"00000001",
  30866=>"00000001",
  30867=>"00000000",
  30868=>"00000001",
  30869=>"00000001",
  30870=>"00000000",
  30871=>"11111110",
  30872=>"11111100",
  30873=>"00000100",
  30874=>"11111100",
  30875=>"00000010",
  30876=>"11111110",
  30877=>"11111100",
  30878=>"00000010",
  30879=>"00000001",
  30880=>"11111110",
  30881=>"00000000",
  30882=>"00000000",
  30883=>"11111111",
  30884=>"11111111",
  30885=>"11111111",
  30886=>"00000001",
  30887=>"00000010",
  30888=>"11111110",
  30889=>"11111101",
  30890=>"11111110",
  30891=>"00000010",
  30892=>"11111110",
  30893=>"00000001",
  30894=>"00000011",
  30895=>"00000010",
  30896=>"00000000",
  30897=>"00000000",
  30898=>"00000000",
  30899=>"00000000",
  30900=>"11111110",
  30901=>"11111110",
  30902=>"00000000",
  30903=>"11111110",
  30904=>"11111111",
  30905=>"00000000",
  30906=>"11111110",
  30907=>"11111110",
  30908=>"00000010",
  30909=>"00000010",
  30910=>"11111110",
  30911=>"00000011",
  30912=>"00000000",
  30913=>"00000000",
  30914=>"11111111",
  30915=>"11111110",
  30916=>"00000010",
  30917=>"11111110",
  30918=>"00000110",
  30919=>"11111110",
  30920=>"11111101",
  30921=>"11111101",
  30922=>"00000011",
  30923=>"11111111",
  30924=>"00000000",
  30925=>"00000001",
  30926=>"00000000",
  30927=>"11111111",
  30928=>"00000000",
  30929=>"11111100",
  30930=>"00000000",
  30931=>"00000010",
  30932=>"11111111",
  30933=>"11111100",
  30934=>"00000010",
  30935=>"00000000",
  30936=>"00000001",
  30937=>"11111110",
  30938=>"00000010",
  30939=>"11111111",
  30940=>"11111111",
  30941=>"00000011",
  30942=>"00000010",
  30943=>"00000000",
  30944=>"11111111",
  30945=>"11111110",
  30946=>"00000011",
  30947=>"11111110",
  30948=>"11111110",
  30949=>"00000001",
  30950=>"11111110",
  30951=>"11111111",
  30952=>"00000010",
  30953=>"11111110",
  30954=>"00000011",
  30955=>"00000001",
  30956=>"11111110",
  30957=>"11111101",
  30958=>"11111100",
  30959=>"00000001",
  30960=>"11111101",
  30961=>"00000010",
  30962=>"11111111",
  30963=>"00000010",
  30964=>"00000000",
  30965=>"00000000",
  30966=>"11111101",
  30967=>"11111110",
  30968=>"00000010",
  30969=>"11111101",
  30970=>"11111111",
  30971=>"00000010",
  30972=>"11111101",
  30973=>"00000010",
  30974=>"00000000",
  30975=>"00000001",
  30976=>"00000011",
  30977=>"11111110",
  30978=>"11111111",
  30979=>"11111101",
  30980=>"11111110",
  30981=>"00000011",
  30982=>"11111110",
  30983=>"00000110",
  30984=>"11111110",
  30985=>"11111101",
  30986=>"00000000",
  30987=>"11111110",
  30988=>"11111111",
  30989=>"11111111",
  30990=>"11111100",
  30991=>"11111101",
  30992=>"11111101",
  30993=>"11111111",
  30994=>"00000001",
  30995=>"00000001",
  30996=>"00000001",
  30997=>"00000100",
  30998=>"00000010",
  30999=>"00000001",
  31000=>"00001000",
  31001=>"11111111",
  31002=>"11111111",
  31003=>"00000010",
  31004=>"00000011",
  31005=>"00000110",
  31006=>"11111111",
  31007=>"00000100",
  31008=>"11111110",
  31009=>"11111100",
  31010=>"00000010",
  31011=>"11111110",
  31012=>"00000001",
  31013=>"11111100",
  31014=>"11111111",
  31015=>"11111101",
  31016=>"11111111",
  31017=>"00000000",
  31018=>"00000100",
  31019=>"11111101",
  31020=>"11111111",
  31021=>"00000000",
  31022=>"00000000",
  31023=>"00000000",
  31024=>"00000110",
  31025=>"11111111",
  31026=>"00000001",
  31027=>"00000001",
  31028=>"11111101",
  31029=>"11111110",
  31030=>"00000010",
  31031=>"11111101",
  31032=>"00000001",
  31033=>"00000000",
  31034=>"11111101",
  31035=>"00000000",
  31036=>"11111111",
  31037=>"11111111",
  31038=>"11111111",
  31039=>"00000001",
  31040=>"00000000",
  31041=>"00000001",
  31042=>"00000011",
  31043=>"11111111",
  31044=>"00000001",
  31045=>"11111110",
  31046=>"00000000",
  31047=>"00000010",
  31048=>"11111101",
  31049=>"00000101",
  31050=>"11111111",
  31051=>"00000000",
  31052=>"11111110",
  31053=>"00000011",
  31054=>"11111101",
  31055=>"11111110",
  31056=>"11111110",
  31057=>"11111111",
  31058=>"11111101",
  31059=>"11111111",
  31060=>"00000001",
  31061=>"11111110",
  31062=>"00000000",
  31063=>"11111111",
  31064=>"00000100",
  31065=>"00000000",
  31066=>"00000001",
  31067=>"11111110",
  31068=>"11111110",
  31069=>"11111110",
  31070=>"11111101",
  31071=>"00000000",
  31072=>"00000010",
  31073=>"11111101",
  31074=>"00000100",
  31075=>"00000010",
  31076=>"11111110",
  31077=>"00000000",
  31078=>"00000000",
  31079=>"11111111",
  31080=>"11111110",
  31081=>"11111101",
  31082=>"00000001",
  31083=>"00000000",
  31084=>"00000001",
  31085=>"00000010",
  31086=>"00000010",
  31087=>"11111110",
  31088=>"11111110",
  31089=>"00000010",
  31090=>"00000000",
  31091=>"00000000",
  31092=>"11111101",
  31093=>"11111110",
  31094=>"11111110",
  31095=>"11111110",
  31096=>"00000001",
  31097=>"00000001",
  31098=>"11111110",
  31099=>"00000001",
  31100=>"00000010",
  31101=>"11111110",
  31102=>"00000010",
  31103=>"00000001",
  31104=>"11111110",
  31105=>"11111111",
  31106=>"00000000",
  31107=>"00000010",
  31108=>"00000010",
  31109=>"11111110",
  31110=>"00000001",
  31111=>"11111101",
  31112=>"11111110",
  31113=>"11111111",
  31114=>"00000100",
  31115=>"11111110",
  31116=>"11111111",
  31117=>"00000001",
  31118=>"11111111",
  31119=>"11111110",
  31120=>"00000001",
  31121=>"11111110",
  31122=>"11111101",
  31123=>"00000011",
  31124=>"11111110",
  31125=>"11111101",
  31126=>"00000010",
  31127=>"11111101",
  31128=>"00000010",
  31129=>"00000000",
  31130=>"11111101",
  31131=>"00000110",
  31132=>"11111111",
  31133=>"00000001",
  31134=>"00000010",
  31135=>"00000010",
  31136=>"11111100",
  31137=>"00000000",
  31138=>"11111111",
  31139=>"00000001",
  31140=>"00000000",
  31141=>"11111101",
  31142=>"11111101",
  31143=>"00000011",
  31144=>"00000011",
  31145=>"00000011",
  31146=>"11111110",
  31147=>"00000000",
  31148=>"00000001",
  31149=>"00000000",
  31150=>"11111101",
  31151=>"11111101",
  31152=>"00000001",
  31153=>"11111101",
  31154=>"00000011",
  31155=>"11111101",
  31156=>"11111101",
  31157=>"00000010",
  31158=>"11111110",
  31159=>"11111110",
  31160=>"00000101",
  31161=>"00000000",
  31162=>"11111101",
  31163=>"11111111",
  31164=>"11111111",
  31165=>"00000001",
  31166=>"11111111",
  31167=>"00000000",
  31168=>"00000000",
  31169=>"00000100",
  31170=>"11111110",
  31171=>"00000010",
  31172=>"11111100",
  31173=>"11111110",
  31174=>"00000001",
  31175=>"00000001",
  31176=>"11111101",
  31177=>"11111111",
  31178=>"00000001",
  31179=>"00000000",
  31180=>"00000000",
  31181=>"00000000",
  31182=>"00000100",
  31183=>"11111111",
  31184=>"00000001",
  31185=>"00000001",
  31186=>"11111111",
  31187=>"00000001",
  31188=>"00000000",
  31189=>"00000000",
  31190=>"00000111",
  31191=>"11111111",
  31192=>"11111110",
  31193=>"00000110",
  31194=>"00000001",
  31195=>"00000000",
  31196=>"00000010",
  31197=>"11111110",
  31198=>"00000000",
  31199=>"11111101",
  31200=>"00000010",
  31201=>"00000001",
  31202=>"11111110",
  31203=>"00000010",
  31204=>"11111110",
  31205=>"00000011",
  31206=>"00000001",
  31207=>"11111110",
  31208=>"00000001",
  31209=>"11111101",
  31210=>"00000101",
  31211=>"00000001",
  31212=>"00000001",
  31213=>"00000001",
  31214=>"00000100",
  31215=>"11111101",
  31216=>"11111110",
  31217=>"11111110",
  31218=>"00000010",
  31219=>"00000000",
  31220=>"00000011",
  31221=>"00000001",
  31222=>"00000001",
  31223=>"00000011",
  31224=>"00000001",
  31225=>"00000000",
  31226=>"11111101",
  31227=>"00000010",
  31228=>"00000000",
  31229=>"00000001",
  31230=>"00000011",
  31231=>"00000001",
  31232=>"00000000",
  31233=>"00000010",
  31234=>"00000000",
  31235=>"00000000",
  31236=>"00000101",
  31237=>"00000011",
  31238=>"00000001",
  31239=>"00000010",
  31240=>"11111110",
  31241=>"00000001",
  31242=>"00000000",
  31243=>"00000001",
  31244=>"11111101",
  31245=>"11111111",
  31246=>"00000011",
  31247=>"11111111",
  31248=>"00000000",
  31249=>"00000110",
  31250=>"00000011",
  31251=>"11111110",
  31252=>"00000000",
  31253=>"00000000",
  31254=>"11111110",
  31255=>"00000001",
  31256=>"11111101",
  31257=>"11111110",
  31258=>"11111111",
  31259=>"00000001",
  31260=>"00000100",
  31261=>"00000001",
  31262=>"11111111",
  31263=>"11111111",
  31264=>"00000001",
  31265=>"00000001",
  31266=>"11111101",
  31267=>"00000011",
  31268=>"11111111",
  31269=>"11111100",
  31270=>"00000011",
  31271=>"11111111",
  31272=>"00000000",
  31273=>"11111110",
  31274=>"11111111",
  31275=>"00000010",
  31276=>"00000001",
  31277=>"11111101",
  31278=>"00000101",
  31279=>"00000001",
  31280=>"11111101",
  31281=>"00000011",
  31282=>"11111110",
  31283=>"00000010",
  31284=>"11111111",
  31285=>"11111101",
  31286=>"11111111",
  31287=>"11111111",
  31288=>"00000001",
  31289=>"11111110",
  31290=>"00000011",
  31291=>"00000000",
  31292=>"11111101",
  31293=>"11111101",
  31294=>"00000001",
  31295=>"11111100",
  31296=>"00000001",
  31297=>"11111110",
  31298=>"00000100",
  31299=>"11111101",
  31300=>"11111110",
  31301=>"00000000",
  31302=>"00000001",
  31303=>"00000101",
  31304=>"00000100",
  31305=>"11111101",
  31306=>"11111111",
  31307=>"11111110",
  31308=>"11111110",
  31309=>"00000000",
  31310=>"11111101",
  31311=>"11111111",
  31312=>"00000010",
  31313=>"11111110",
  31314=>"00000100",
  31315=>"11111111",
  31316=>"11111110",
  31317=>"11111101",
  31318=>"11111111",
  31319=>"00000010",
  31320=>"00000001",
  31321=>"11111111",
  31322=>"11111111",
  31323=>"00000000",
  31324=>"11111111",
  31325=>"11111110",
  31326=>"00000000",
  31327=>"11111101",
  31328=>"00000001",
  31329=>"00000001",
  31330=>"11111111",
  31331=>"00000011",
  31332=>"11111101",
  31333=>"11111110",
  31334=>"11111111",
  31335=>"00000011",
  31336=>"11111101",
  31337=>"00000101",
  31338=>"11111101",
  31339=>"11111111",
  31340=>"11111101",
  31341=>"11111101",
  31342=>"11111111",
  31343=>"11111101",
  31344=>"11111110",
  31345=>"00000000",
  31346=>"11111111",
  31347=>"00000001",
  31348=>"00000010",
  31349=>"00000001",
  31350=>"00000001",
  31351=>"11111101",
  31352=>"00000101",
  31353=>"00000011",
  31354=>"00000101",
  31355=>"00000001",
  31356=>"11111110",
  31357=>"11111111",
  31358=>"11111110",
  31359=>"00000010",
  31360=>"00000011",
  31361=>"00000000",
  31362=>"11111110",
  31363=>"11111101",
  31364=>"00000000",
  31365=>"00000001",
  31366=>"00000100",
  31367=>"00000001",
  31368=>"11111111",
  31369=>"00000010",
  31370=>"11111101",
  31371=>"00000001",
  31372=>"11111110",
  31373=>"00000001",
  31374=>"00000010",
  31375=>"00000000",
  31376=>"11111110",
  31377=>"11111110",
  31378=>"11111110",
  31379=>"00000011",
  31380=>"11111100",
  31381=>"11111101",
  31382=>"11111110",
  31383=>"00000110",
  31384=>"00000011",
  31385=>"00000011",
  31386=>"11111111",
  31387=>"11111111",
  31388=>"11111110",
  31389=>"00000000",
  31390=>"00000010",
  31391=>"11111110",
  31392=>"11111110",
  31393=>"00000000",
  31394=>"11111111",
  31395=>"00000100",
  31396=>"00000001",
  31397=>"11111111",
  31398=>"00000000",
  31399=>"11111111",
  31400=>"11111101",
  31401=>"00000001",
  31402=>"11111100",
  31403=>"11111110",
  31404=>"00000000",
  31405=>"11111110",
  31406=>"00000001",
  31407=>"00000011",
  31408=>"11111111",
  31409=>"11111110",
  31410=>"00000010",
  31411=>"11111110",
  31412=>"11111111",
  31413=>"00000110",
  31414=>"00000001",
  31415=>"11111110",
  31416=>"00000001",
  31417=>"00000000",
  31418=>"11111111",
  31419=>"11111110",
  31420=>"11111110",
  31421=>"11111110",
  31422=>"11111110",
  31423=>"00000001",
  31424=>"11111111",
  31425=>"00000000",
  31426=>"00000000",
  31427=>"00000101",
  31428=>"00000010",
  31429=>"11111101",
  31430=>"11111110",
  31431=>"11111100",
  31432=>"00000001",
  31433=>"11111101",
  31434=>"00000000",
  31435=>"11111110",
  31436=>"11111110",
  31437=>"11111110",
  31438=>"11111110",
  31439=>"00000000",
  31440=>"11111111",
  31441=>"11111110",
  31442=>"11111101",
  31443=>"11111111",
  31444=>"00000010",
  31445=>"11111111",
  31446=>"00000010",
  31447=>"00000000",
  31448=>"11111101",
  31449=>"11111101",
  31450=>"00000001",
  31451=>"00000000",
  31452=>"11111111",
  31453=>"11111101",
  31454=>"00000011",
  31455=>"11111111",
  31456=>"00000000",
  31457=>"11111111",
  31458=>"00000000",
  31459=>"00000001",
  31460=>"11111111",
  31461=>"00000000",
  31462=>"00000000",
  31463=>"11111101",
  31464=>"00000011",
  31465=>"00000011",
  31466=>"00000001",
  31467=>"11111110",
  31468=>"11111110",
  31469=>"00000101",
  31470=>"00000010",
  31471=>"00000000",
  31472=>"00000100",
  31473=>"00000010",
  31474=>"00000010",
  31475=>"00000010",
  31476=>"00000000",
  31477=>"00000000",
  31478=>"00000000",
  31479=>"11111111",
  31480=>"11111111",
  31481=>"11111110",
  31482=>"00000011",
  31483=>"00000000",
  31484=>"11111111",
  31485=>"00000010",
  31486=>"11111101",
  31487=>"00000010",
  31488=>"00000111",
  31489=>"00000001",
  31490=>"00000000",
  31491=>"11111110",
  31492=>"11111110",
  31493=>"11111110",
  31494=>"00000000",
  31495=>"11111101",
  31496=>"11111101",
  31497=>"11111101",
  31498=>"00000000",
  31499=>"11111101",
  31500=>"00000010",
  31501=>"00000000",
  31502=>"11111111",
  31503=>"00000001",
  31504=>"11111110",
  31505=>"00000010",
  31506=>"11111111",
  31507=>"00000000",
  31508=>"11111101",
  31509=>"00000010",
  31510=>"11111101",
  31511=>"00000000",
  31512=>"11111101",
  31513=>"00000010",
  31514=>"00000001",
  31515=>"11111111",
  31516=>"00000000",
  31517=>"00000001",
  31518=>"11111110",
  31519=>"00000000",
  31520=>"11111111",
  31521=>"00000100",
  31522=>"00000001",
  31523=>"11111111",
  31524=>"11111110",
  31525=>"11111101",
  31526=>"00000100",
  31527=>"11111101",
  31528=>"11111110",
  31529=>"11111101",
  31530=>"11111111",
  31531=>"11111111",
  31532=>"00000000",
  31533=>"11111110",
  31534=>"00000100",
  31535=>"00000001",
  31536=>"00000010",
  31537=>"11111110",
  31538=>"11111110",
  31539=>"00000000",
  31540=>"11111111",
  31541=>"11111110",
  31542=>"11111111",
  31543=>"00000000",
  31544=>"11111110",
  31545=>"00000010",
  31546=>"00000010",
  31547=>"00000001",
  31548=>"11111110",
  31549=>"11111110",
  31550=>"11111110",
  31551=>"11111111",
  31552=>"00000001",
  31553=>"00000001",
  31554=>"11111101",
  31555=>"00000000",
  31556=>"11111100",
  31557=>"00000001",
  31558=>"00000000",
  31559=>"11111111",
  31560=>"11111110",
  31561=>"11111111",
  31562=>"00000010",
  31563=>"11111111",
  31564=>"11111111",
  31565=>"00000000",
  31566=>"11111110",
  31567=>"00000010",
  31568=>"00000001",
  31569=>"00000001",
  31570=>"11111111",
  31571=>"11111101",
  31572=>"00000000",
  31573=>"00000010",
  31574=>"00000001",
  31575=>"00000010",
  31576=>"00000000",
  31577=>"00000000",
  31578=>"00000001",
  31579=>"00000000",
  31580=>"00000010",
  31581=>"00000000",
  31582=>"11111100",
  31583=>"11111110",
  31584=>"00000001",
  31585=>"11111110",
  31586=>"00000000",
  31587=>"11111110",
  31588=>"11111111",
  31589=>"11111110",
  31590=>"00000100",
  31591=>"11111100",
  31592=>"00000011",
  31593=>"00000011",
  31594=>"00000000",
  31595=>"00000010",
  31596=>"11111101",
  31597=>"00000000",
  31598=>"00000010",
  31599=>"00000010",
  31600=>"11111110",
  31601=>"11111110",
  31602=>"11111110",
  31603=>"11111101",
  31604=>"11111110",
  31605=>"00000001",
  31606=>"00000000",
  31607=>"00000001",
  31608=>"11111111",
  31609=>"00000000",
  31610=>"11111100",
  31611=>"11111101",
  31612=>"00000001",
  31613=>"11111101",
  31614=>"11111110",
  31615=>"00000001",
  31616=>"11111111",
  31617=>"11111101",
  31618=>"00000000",
  31619=>"11111110",
  31620=>"00000011",
  31621=>"00000000",
  31622=>"11111111",
  31623=>"11111110",
  31624=>"00000010",
  31625=>"00000100",
  31626=>"11111111",
  31627=>"11111101",
  31628=>"00000110",
  31629=>"11111101",
  31630=>"00000011",
  31631=>"00000010",
  31632=>"00000000",
  31633=>"11111100",
  31634=>"11111111",
  31635=>"00000000",
  31636=>"00000000",
  31637=>"11111111",
  31638=>"00000011",
  31639=>"00000010",
  31640=>"11111101",
  31641=>"00000100",
  31642=>"11111101",
  31643=>"00000000",
  31644=>"11111101",
  31645=>"00000000",
  31646=>"00000001",
  31647=>"11111110",
  31648=>"11111111",
  31649=>"11111110",
  31650=>"00000010",
  31651=>"11111110",
  31652=>"00000001",
  31653=>"00000011",
  31654=>"11111110",
  31655=>"00000011",
  31656=>"00000011",
  31657=>"00000010",
  31658=>"00000001",
  31659=>"00000001",
  31660=>"00000000",
  31661=>"00000001",
  31662=>"00000000",
  31663=>"11111101",
  31664=>"00000001",
  31665=>"00000000",
  31666=>"00000000",
  31667=>"00000000",
  31668=>"11111110",
  31669=>"11111111",
  31670=>"11111111",
  31671=>"00000000",
  31672=>"11111111",
  31673=>"00000001",
  31674=>"11111101",
  31675=>"00000000",
  31676=>"00000101",
  31677=>"00000100",
  31678=>"00000001",
  31679=>"00000000",
  31680=>"00000100",
  31681=>"11111111",
  31682=>"00000000",
  31683=>"00000000",
  31684=>"11111111",
  31685=>"00000010",
  31686=>"11111110",
  31687=>"11111111",
  31688=>"11111111",
  31689=>"11111101",
  31690=>"00000100",
  31691=>"11111101",
  31692=>"00000010",
  31693=>"00000000",
  31694=>"11111110",
  31695=>"00000001",
  31696=>"00000001",
  31697=>"00000011",
  31698=>"00000101",
  31699=>"11111101",
  31700=>"11111110",
  31701=>"11111111",
  31702=>"11111110",
  31703=>"00000000",
  31704=>"00000011",
  31705=>"11111111",
  31706=>"11111101",
  31707=>"00000101",
  31708=>"11111101",
  31709=>"00000011",
  31710=>"00000000",
  31711=>"11111100",
  31712=>"11111110",
  31713=>"00000101",
  31714=>"00000001",
  31715=>"00000001",
  31716=>"00000010",
  31717=>"11111110",
  31718=>"00000110",
  31719=>"11111110",
  31720=>"00000001",
  31721=>"00000001",
  31722=>"11111101",
  31723=>"11111110",
  31724=>"00000010",
  31725=>"11111110",
  31726=>"00000011",
  31727=>"00000010",
  31728=>"11111101",
  31729=>"00000001",
  31730=>"00000100",
  31731=>"11111110",
  31732=>"11111101",
  31733=>"11111111",
  31734=>"00000001",
  31735=>"11111100",
  31736=>"00000001",
  31737=>"11111101",
  31738=>"11111101",
  31739=>"00000001",
  31740=>"00000011",
  31741=>"11111111",
  31742=>"00000100",
  31743=>"11111110",
  31744=>"00000000",
  31745=>"00000000",
  31746=>"00000010",
  31747=>"11111110",
  31748=>"00000100",
  31749=>"00000010",
  31750=>"11111111",
  31751=>"11111101",
  31752=>"00000000",
  31753=>"00000000",
  31754=>"11111111",
  31755=>"00000010",
  31756=>"00000010",
  31757=>"11111100",
  31758=>"00000001",
  31759=>"11111100",
  31760=>"00000000",
  31761=>"00000001",
  31762=>"11111111",
  31763=>"00000010",
  31764=>"00000100",
  31765=>"11111111",
  31766=>"00000010",
  31767=>"11111111",
  31768=>"11111111",
  31769=>"00000011",
  31770=>"11111100",
  31771=>"11111110",
  31772=>"11111111",
  31773=>"00000010",
  31774=>"11111111",
  31775=>"00000001",
  31776=>"00000000",
  31777=>"00000000",
  31778=>"00000000",
  31779=>"11111110",
  31780=>"11111110",
  31781=>"11111110",
  31782=>"00000010",
  31783=>"00000010",
  31784=>"00000010",
  31785=>"11111100",
  31786=>"00000001",
  31787=>"00000001",
  31788=>"11111101",
  31789=>"11111110",
  31790=>"00000010",
  31791=>"00000011",
  31792=>"00000001",
  31793=>"11111110",
  31794=>"00000000",
  31795=>"11111111",
  31796=>"00000000",
  31797=>"00000000",
  31798=>"00000000",
  31799=>"00000101",
  31800=>"00000000",
  31801=>"00000010",
  31802=>"00000011",
  31803=>"00000100",
  31804=>"00000000",
  31805=>"11111111",
  31806=>"11111111",
  31807=>"00000100",
  31808=>"00000011",
  31809=>"00000000",
  31810=>"11111111",
  31811=>"11111101",
  31812=>"00000010",
  31813=>"11111111",
  31814=>"00000010",
  31815=>"11111111",
  31816=>"11111110",
  31817=>"00000101",
  31818=>"11111111",
  31819=>"00000000",
  31820=>"00000010",
  31821=>"11111101",
  31822=>"11111111",
  31823=>"11111111",
  31824=>"11111101",
  31825=>"11111011",
  31826=>"11111111",
  31827=>"00000010",
  31828=>"00000000",
  31829=>"11111110",
  31830=>"11111111",
  31831=>"11111101",
  31832=>"00000000",
  31833=>"11111110",
  31834=>"00000010",
  31835=>"11111101",
  31836=>"00000101",
  31837=>"11111110",
  31838=>"11111101",
  31839=>"00000000",
  31840=>"00000010",
  31841=>"00000000",
  31842=>"00000000",
  31843=>"00000000",
  31844=>"00000001",
  31845=>"00000000",
  31846=>"11111101",
  31847=>"11111101",
  31848=>"11111101",
  31849=>"00000010",
  31850=>"11111111",
  31851=>"00000100",
  31852=>"00000000",
  31853=>"00001000",
  31854=>"11111110",
  31855=>"00000010",
  31856=>"00000000",
  31857=>"00000011",
  31858=>"00000010",
  31859=>"00000000",
  31860=>"11111111",
  31861=>"11111101",
  31862=>"11111111",
  31863=>"00000010",
  31864=>"00000000",
  31865=>"00000010",
  31866=>"00000111",
  31867=>"00000000",
  31868=>"00000010",
  31869=>"11111100",
  31870=>"11111101",
  31871=>"00000001",
  31872=>"11111111",
  31873=>"00000100",
  31874=>"11111111",
  31875=>"00000000",
  31876=>"11111101",
  31877=>"00000000",
  31878=>"00000000",
  31879=>"11111111",
  31880=>"11111011",
  31881=>"11111101",
  31882=>"00000000",
  31883=>"00000010",
  31884=>"11111101",
  31885=>"00000010",
  31886=>"00000000",
  31887=>"11111100",
  31888=>"00000000",
  31889=>"11111110",
  31890=>"00000001",
  31891=>"00000010",
  31892=>"11111111",
  31893=>"11111110",
  31894=>"00000000",
  31895=>"00000010",
  31896=>"00000101",
  31897=>"11111111",
  31898=>"11111111",
  31899=>"00000000",
  31900=>"00000010",
  31901=>"00000000",
  31902=>"00000001",
  31903=>"11111111",
  31904=>"11111110",
  31905=>"00000111",
  31906=>"00000011",
  31907=>"11111111",
  31908=>"00000001",
  31909=>"11111111",
  31910=>"00000010",
  31911=>"00000000",
  31912=>"11111111",
  31913=>"11111111",
  31914=>"11111110",
  31915=>"00000001",
  31916=>"00000000",
  31917=>"00000001",
  31918=>"00000000",
  31919=>"00000001",
  31920=>"00000000",
  31921=>"11111111",
  31922=>"00000000",
  31923=>"11111110",
  31924=>"00000010",
  31925=>"00000001",
  31926=>"11111110",
  31927=>"00000001",
  31928=>"11111101",
  31929=>"00000000",
  31930=>"11111110",
  31931=>"00000011",
  31932=>"11111110",
  31933=>"00000010",
  31934=>"11111111",
  31935=>"11111101",
  31936=>"00000011",
  31937=>"11111111",
  31938=>"00000010",
  31939=>"11111111",
  31940=>"00000000",
  31941=>"11111111",
  31942=>"00000100",
  31943=>"11111101",
  31944=>"00000011",
  31945=>"11111100",
  31946=>"00000011",
  31947=>"11111100",
  31948=>"00000001",
  31949=>"00000000",
  31950=>"00000001",
  31951=>"00000000",
  31952=>"00000001",
  31953=>"11111111",
  31954=>"00000001",
  31955=>"00000000",
  31956=>"11111110",
  31957=>"00000100",
  31958=>"00000010",
  31959=>"11111101",
  31960=>"11111111",
  31961=>"11111111",
  31962=>"11111110",
  31963=>"00000000",
  31964=>"11111110",
  31965=>"00000000",
  31966=>"00000010",
  31967=>"11111101",
  31968=>"00000011",
  31969=>"00000000",
  31970=>"00000001",
  31971=>"11111111",
  31972=>"11111101",
  31973=>"00000000",
  31974=>"00000000",
  31975=>"11111101",
  31976=>"00000001",
  31977=>"11111110",
  31978=>"11111110",
  31979=>"11111110",
  31980=>"00000000",
  31981=>"11111100",
  31982=>"00000010",
  31983=>"11111110",
  31984=>"00000000",
  31985=>"11111110",
  31986=>"00000000",
  31987=>"00000011",
  31988=>"11111111",
  31989=>"00000001",
  31990=>"00000010",
  31991=>"00000011",
  31992=>"00000100",
  31993=>"11111101",
  31994=>"11111111",
  31995=>"11111110",
  31996=>"00000001",
  31997=>"11111110",
  31998=>"11111101",
  31999=>"11111111",
  32000=>"00000010",
  32001=>"00000000",
  32002=>"00000011",
  32003=>"11111110",
  32004=>"11111110",
  32005=>"11111110",
  32006=>"11111101",
  32007=>"00000001",
  32008=>"00000000",
  32009=>"11111101",
  32010=>"00000100",
  32011=>"00000011",
  32012=>"11111111",
  32013=>"00000011",
  32014=>"00000011",
  32015=>"00000100",
  32016=>"11111100",
  32017=>"11111110",
  32018=>"11111111",
  32019=>"11111101",
  32020=>"11111101",
  32021=>"11111111",
  32022=>"11111101",
  32023=>"00000001",
  32024=>"11111110",
  32025=>"00000000",
  32026=>"00000010",
  32027=>"00000011",
  32028=>"00000001",
  32029=>"11111110",
  32030=>"11111111",
  32031=>"00000000",
  32032=>"00000100",
  32033=>"11111110",
  32034=>"00000010",
  32035=>"11111100",
  32036=>"11111111",
  32037=>"11111101",
  32038=>"00000010",
  32039=>"11111111",
  32040=>"11111111",
  32041=>"00000100",
  32042=>"11111111",
  32043=>"00000010",
  32044=>"11111111",
  32045=>"11111111",
  32046=>"00000000",
  32047=>"11111111",
  32048=>"00000001",
  32049=>"11111110",
  32050=>"00000011",
  32051=>"11111101",
  32052=>"11111110",
  32053=>"11111011",
  32054=>"00000011",
  32055=>"00000011",
  32056=>"00000100",
  32057=>"00000011",
  32058=>"00000010",
  32059=>"11111111",
  32060=>"00000011",
  32061=>"11111110",
  32062=>"00000001",
  32063=>"00000011",
  32064=>"11111110",
  32065=>"11111111",
  32066=>"11111110",
  32067=>"00000000",
  32068=>"11111111",
  32069=>"00000011",
  32070=>"11111011",
  32071=>"00000100",
  32072=>"00000010",
  32073=>"00000000",
  32074=>"11111110",
  32075=>"11111111",
  32076=>"11111101",
  32077=>"00000011",
  32078=>"00000011",
  32079=>"00000010",
  32080=>"11111101",
  32081=>"00000011",
  32082=>"11111100",
  32083=>"00000000",
  32084=>"11111101",
  32085=>"00000011",
  32086=>"00000000",
  32087=>"00000001",
  32088=>"00000011",
  32089=>"11111111",
  32090=>"00000001",
  32091=>"00000000",
  32092=>"00000000",
  32093=>"11111111",
  32094=>"11111111",
  32095=>"00000000",
  32096=>"11111111",
  32097=>"00000000",
  32098=>"11111111",
  32099=>"11111100",
  32100=>"00000000",
  32101=>"11111111",
  32102=>"00000010",
  32103=>"11111111",
  32104=>"00000101",
  32105=>"11111110",
  32106=>"00000001",
  32107=>"00000011",
  32108=>"11111110",
  32109=>"00000001",
  32110=>"00000100",
  32111=>"11111110",
  32112=>"11111111",
  32113=>"00000011",
  32114=>"00000011",
  32115=>"00000010",
  32116=>"00000010",
  32117=>"11111110",
  32118=>"11111110",
  32119=>"00000000",
  32120=>"00000010",
  32121=>"00000100",
  32122=>"11111110",
  32123=>"00000101",
  32124=>"11111101",
  32125=>"00000001",
  32126=>"00000001",
  32127=>"00000100",
  32128=>"00000000",
  32129=>"00000001",
  32130=>"00000001",
  32131=>"11111101",
  32132=>"11111110",
  32133=>"00000101",
  32134=>"11111111",
  32135=>"11111110",
  32136=>"00000100",
  32137=>"11111101",
  32138=>"11111101",
  32139=>"11111110",
  32140=>"00000001",
  32141=>"11111100",
  32142=>"00000000",
  32143=>"00000010",
  32144=>"00000011",
  32145=>"11111111",
  32146=>"11111101",
  32147=>"00000001",
  32148=>"11111111",
  32149=>"00000001",
  32150=>"00000000",
  32151=>"11111110",
  32152=>"11111101",
  32153=>"11111111",
  32154=>"11111100",
  32155=>"11111111",
  32156=>"00000000",
  32157=>"00000011",
  32158=>"11111101",
  32159=>"00000010",
  32160=>"00000011",
  32161=>"11111101",
  32162=>"11111011",
  32163=>"00000010",
  32164=>"00000010",
  32165=>"11111111",
  32166=>"00000010",
  32167=>"00000010",
  32168=>"00000100",
  32169=>"11111100",
  32170=>"00000011",
  32171=>"11111111",
  32172=>"11111101",
  32173=>"11111111",
  32174=>"11111101",
  32175=>"00000010",
  32176=>"00000011",
  32177=>"11111111",
  32178=>"00000001",
  32179=>"00000010",
  32180=>"00000011",
  32181=>"11111110",
  32182=>"00000001",
  32183=>"11111101",
  32184=>"00000000",
  32185=>"11111101",
  32186=>"00000010",
  32187=>"11111100",
  32188=>"00000010",
  32189=>"00000011",
  32190=>"11111011",
  32191=>"00000000",
  32192=>"00000010",
  32193=>"11111100",
  32194=>"11111110",
  32195=>"11111111",
  32196=>"00000001",
  32197=>"11111101",
  32198=>"11111110",
  32199=>"11111111",
  32200=>"11111111",
  32201=>"11111111",
  32202=>"00000001",
  32203=>"00000010",
  32204=>"00000000",
  32205=>"00000010",
  32206=>"11111110",
  32207=>"00000010",
  32208=>"11111111",
  32209=>"11111101",
  32210=>"11111111",
  32211=>"11111111",
  32212=>"11111110",
  32213=>"11111110",
  32214=>"00000000",
  32215=>"00000001",
  32216=>"11111111",
  32217=>"00000011",
  32218=>"11111101",
  32219=>"11111110",
  32220=>"11111110",
  32221=>"11111110",
  32222=>"00000010",
  32223=>"00000011",
  32224=>"11111111",
  32225=>"00000010",
  32226=>"00000000",
  32227=>"00000001",
  32228=>"11111110",
  32229=>"00000110",
  32230=>"11111100",
  32231=>"11111111",
  32232=>"00000111",
  32233=>"00000000",
  32234=>"11111111",
  32235=>"00000000",
  32236=>"11111111",
  32237=>"00000100",
  32238=>"00000000",
  32239=>"00000010",
  32240=>"00000011",
  32241=>"00000010",
  32242=>"00000000",
  32243=>"11111100",
  32244=>"11111101",
  32245=>"11111100",
  32246=>"00000100",
  32247=>"11111111",
  32248=>"11111111",
  32249=>"00000011",
  32250=>"00000010",
  32251=>"00000000",
  32252=>"11111100",
  32253=>"11111110",
  32254=>"11111110",
  32255=>"11111110",
  32256=>"11111111",
  32257=>"00000010",
  32258=>"00000101",
  32259=>"11111111",
  32260=>"00000001",
  32261=>"00000010",
  32262=>"00001000",
  32263=>"00000000",
  32264=>"00000001",
  32265=>"00000000",
  32266=>"11111111",
  32267=>"11111101",
  32268=>"00000000",
  32269=>"00000010",
  32270=>"11111100",
  32271=>"11111110",
  32272=>"00000001",
  32273=>"00000000",
  32274=>"00000010",
  32275=>"00000010",
  32276=>"11111111",
  32277=>"11111111",
  32278=>"11111111",
  32279=>"00000011",
  32280=>"11111101",
  32281=>"11111100",
  32282=>"11111110",
  32283=>"11111111",
  32284=>"00000000",
  32285=>"00000011",
  32286=>"00000000",
  32287=>"00000010",
  32288=>"00000000",
  32289=>"11111111",
  32290=>"00000000",
  32291=>"11111111",
  32292=>"11111111",
  32293=>"11111111",
  32294=>"00000010",
  32295=>"00000100",
  32296=>"00000001",
  32297=>"00000000",
  32298=>"11111011",
  32299=>"11111100",
  32300=>"11111101",
  32301=>"11111101",
  32302=>"11111110",
  32303=>"00000111",
  32304=>"11111111",
  32305=>"00000001",
  32306=>"00000001",
  32307=>"00000100",
  32308=>"11111100",
  32309=>"11111011",
  32310=>"00000000",
  32311=>"11111111",
  32312=>"11111110",
  32313=>"00000010",
  32314=>"00000001",
  32315=>"00000110",
  32316=>"00000010",
  32317=>"11111101",
  32318=>"00000010",
  32319=>"11111101",
  32320=>"00000000",
  32321=>"11111100",
  32322=>"11111101",
  32323=>"00000010",
  32324=>"11111110",
  32325=>"11111101",
  32326=>"00000000",
  32327=>"11111101",
  32328=>"11111111",
  32329=>"00000010",
  32330=>"11111110",
  32331=>"11111111",
  32332=>"00000010",
  32333=>"00000001",
  32334=>"00000000",
  32335=>"11111110",
  32336=>"11111111",
  32337=>"11111011",
  32338=>"11111101",
  32339=>"11111110",
  32340=>"11111111",
  32341=>"00000101",
  32342=>"00000000",
  32343=>"00000000",
  32344=>"00000000",
  32345=>"11111110",
  32346=>"11111111",
  32347=>"00000010",
  32348=>"11111110",
  32349=>"00000011",
  32350=>"11111101",
  32351=>"00000001",
  32352=>"00000110",
  32353=>"11111110",
  32354=>"00000000",
  32355=>"11111110",
  32356=>"00000000",
  32357=>"11111111",
  32358=>"11111111",
  32359=>"00000010",
  32360=>"11111101",
  32361=>"11111111",
  32362=>"11111111",
  32363=>"00000011",
  32364=>"00000101",
  32365=>"00000001",
  32366=>"11111111",
  32367=>"11111101",
  32368=>"00000011",
  32369=>"11111110",
  32370=>"00000001",
  32371=>"11111100",
  32372=>"00000011",
  32373=>"11111111",
  32374=>"00000001",
  32375=>"11111110",
  32376=>"11111111",
  32377=>"00000010",
  32378=>"11111110",
  32379=>"00000000",
  32380=>"00000010",
  32381=>"11111110",
  32382=>"00000000",
  32383=>"00000010",
  32384=>"00000000",
  32385=>"11111101",
  32386=>"11111110",
  32387=>"11111101",
  32388=>"00000001",
  32389=>"00000000",
  32390=>"00000100",
  32391=>"00000011",
  32392=>"00000010",
  32393=>"11111110",
  32394=>"00000001",
  32395=>"00000100",
  32396=>"00000011",
  32397=>"00000011",
  32398=>"11111110",
  32399=>"00000001",
  32400=>"11111100",
  32401=>"00000001",
  32402=>"00000001",
  32403=>"00000010",
  32404=>"00000101",
  32405=>"00000000",
  32406=>"11111111",
  32407=>"00000000",
  32408=>"11111111",
  32409=>"11111111",
  32410=>"11111110",
  32411=>"11111110",
  32412=>"00000101",
  32413=>"00000000",
  32414=>"11111101",
  32415=>"00000000",
  32416=>"00000001",
  32417=>"11111100",
  32418=>"00000000",
  32419=>"11111110",
  32420=>"00000001",
  32421=>"11111111",
  32422=>"00000101",
  32423=>"00000001",
  32424=>"00000010",
  32425=>"00000000",
  32426=>"00000001",
  32427=>"00000001",
  32428=>"00000000",
  32429=>"00000000",
  32430=>"11111111",
  32431=>"00000000",
  32432=>"00000000",
  32433=>"11111100",
  32434=>"11111111",
  32435=>"11111111",
  32436=>"00000010",
  32437=>"00000001",
  32438=>"00000001",
  32439=>"11111100",
  32440=>"11111111",
  32441=>"00000001",
  32442=>"11111110",
  32443=>"11111111",
  32444=>"11111111",
  32445=>"11111111",
  32446=>"11111101",
  32447=>"11111111",
  32448=>"00000000",
  32449=>"00000000",
  32450=>"11111111",
  32451=>"11111101",
  32452=>"11111110",
  32453=>"00000001",
  32454=>"00000001",
  32455=>"00000000",
  32456=>"11111110",
  32457=>"11111101",
  32458=>"11111100",
  32459=>"00000000",
  32460=>"00000100",
  32461=>"11111110",
  32462=>"11111101",
  32463=>"11111101",
  32464=>"00000001",
  32465=>"00000001",
  32466=>"11111111",
  32467=>"11111111",
  32468=>"11111111",
  32469=>"11111101",
  32470=>"11111111",
  32471=>"00000000",
  32472=>"11111100",
  32473=>"00000001",
  32474=>"11111111",
  32475=>"00000000",
  32476=>"11111111",
  32477=>"11111110",
  32478=>"00000010",
  32479=>"00000000",
  32480=>"00000100",
  32481=>"11111110",
  32482=>"00000001",
  32483=>"00000010",
  32484=>"00000010",
  32485=>"11111111",
  32486=>"00000001",
  32487=>"00000010",
  32488=>"11111110",
  32489=>"00000010",
  32490=>"00000000",
  32491=>"11111101",
  32492=>"11111110",
  32493=>"00000001",
  32494=>"11111101",
  32495=>"00000100",
  32496=>"11111110",
  32497=>"00000000",
  32498=>"11111110",
  32499=>"00000000",
  32500=>"00000000",
  32501=>"00000010",
  32502=>"11111110",
  32503=>"00000001",
  32504=>"11111111",
  32505=>"00000000",
  32506=>"11111111",
  32507=>"00000010",
  32508=>"00000001",
  32509=>"11111110",
  32510=>"11111100",
  32511=>"00000001",
  32512=>"11111110",
  32513=>"00000001",
  32514=>"00000011",
  32515=>"11111101",
  32516=>"00000101",
  32517=>"00000000",
  32518=>"00000010",
  32519=>"11111101",
  32520=>"11111100",
  32521=>"11111111",
  32522=>"11111111",
  32523=>"11111110",
  32524=>"00000011",
  32525=>"11111111",
  32526=>"11111101",
  32527=>"11111110",
  32528=>"11111101",
  32529=>"00000000",
  32530=>"00000000",
  32531=>"00000010",
  32532=>"11111111",
  32533=>"00000011",
  32534=>"00000010",
  32535=>"00000000",
  32536=>"11111111",
  32537=>"11111011",
  32538=>"11111101",
  32539=>"11111110",
  32540=>"11111100",
  32541=>"11111100",
  32542=>"00000011",
  32543=>"00000000",
  32544=>"00000010",
  32545=>"00000001",
  32546=>"11111111",
  32547=>"00000101",
  32548=>"00000011",
  32549=>"00000001",
  32550=>"11111101",
  32551=>"11111100",
  32552=>"00000001",
  32553=>"00000010",
  32554=>"11111111",
  32555=>"00000011",
  32556=>"11111110",
  32557=>"00000010",
  32558=>"00000001",
  32559=>"11111110",
  32560=>"11111110",
  32561=>"11111110",
  32562=>"11111110",
  32563=>"11111111",
  32564=>"11111111",
  32565=>"11111011",
  32566=>"11111110",
  32567=>"00000001",
  32568=>"11111101",
  32569=>"11111111",
  32570=>"00000110",
  32571=>"11111110",
  32572=>"00000001",
  32573=>"00000010",
  32574=>"00000000",
  32575=>"11111111",
  32576=>"11111111",
  32577=>"00000010",
  32578=>"11111111",
  32579=>"11111111",
  32580=>"11111111",
  32581=>"00000001",
  32582=>"00000010",
  32583=>"11111101",
  32584=>"11111111",
  32585=>"00000010",
  32586=>"00000000",
  32587=>"00000000",
  32588=>"00000010",
  32589=>"00000000",
  32590=>"00000100",
  32591=>"00000010",
  32592=>"00000010",
  32593=>"11111110",
  32594=>"11111110",
  32595=>"11111110",
  32596=>"11111110",
  32597=>"11111111",
  32598=>"00000010",
  32599=>"11111111",
  32600=>"00000100",
  32601=>"00000010",
  32602=>"00000000",
  32603=>"11111111",
  32604=>"00000011",
  32605=>"11111101",
  32606=>"00000001",
  32607=>"11111110",
  32608=>"11111100",
  32609=>"11111110",
  32610=>"00000010",
  32611=>"11111111",
  32612=>"11111110",
  32613=>"00000010",
  32614=>"11111110",
  32615=>"00000010",
  32616=>"00000000",
  32617=>"11111100",
  32618=>"11111101",
  32619=>"11111100",
  32620=>"00000000",
  32621=>"00000001",
  32622=>"00000100",
  32623=>"00000000",
  32624=>"11111110",
  32625=>"11111100",
  32626=>"00000010",
  32627=>"00000001",
  32628=>"00000001",
  32629=>"00000000",
  32630=>"00000011",
  32631=>"11111111",
  32632=>"11111110",
  32633=>"00000011",
  32634=>"00000100",
  32635=>"11111101",
  32636=>"11111111",
  32637=>"00000001",
  32638=>"11111111",
  32639=>"00000010",
  32640=>"00000011",
  32641=>"11111110",
  32642=>"11111110",
  32643=>"11111011",
  32644=>"00000000",
  32645=>"11111111",
  32646=>"11111110",
  32647=>"00000101",
  32648=>"11111111",
  32649=>"11111110",
  32650=>"11111101",
  32651=>"11111100",
  32652=>"11111111",
  32653=>"00000010",
  32654=>"11111110",
  32655=>"00000001",
  32656=>"11111110",
  32657=>"11111100",
  32658=>"11111100",
  32659=>"00000010",
  32660=>"00000011",
  32661=>"11111101",
  32662=>"11111110",
  32663=>"11111110",
  32664=>"00000001",
  32665=>"00000100",
  32666=>"11111111",
  32667=>"11111111",
  32668=>"00000000",
  32669=>"00000001",
  32670=>"11111101",
  32671=>"00000011",
  32672=>"11111100",
  32673=>"11111111",
  32674=>"00000000",
  32675=>"00000000",
  32676=>"00000001",
  32677=>"00000101",
  32678=>"00000010",
  32679=>"11111101",
  32680=>"00000000",
  32681=>"00000001",
  32682=>"00000000",
  32683=>"00000011",
  32684=>"00000000",
  32685=>"00000011",
  32686=>"00000010",
  32687=>"00000011",
  32688=>"11111111",
  32689=>"00000110",
  32690=>"00000001",
  32691=>"11111110",
  32692=>"11111111",
  32693=>"00000000",
  32694=>"00000000",
  32695=>"00000110",
  32696=>"00000001",
  32697=>"11111110",
  32698=>"11111111",
  32699=>"11111111",
  32700=>"00000000",
  32701=>"00000000",
  32702=>"00000010",
  32703=>"00000010",
  32704=>"00000001",
  32705=>"11111111",
  32706=>"00000010",
  32707=>"11111111",
  32708=>"11111111",
  32709=>"11111110",
  32710=>"00000001",
  32711=>"00000010",
  32712=>"00000001",
  32713=>"00000100",
  32714=>"00000010",
  32715=>"00000000",
  32716=>"00000011",
  32717=>"11111111",
  32718=>"11111101",
  32719=>"11111110",
  32720=>"00000001",
  32721=>"00000100",
  32722=>"11111101",
  32723=>"00000010",
  32724=>"11111110",
  32725=>"11111100",
  32726=>"00000000",
  32727=>"11111101",
  32728=>"11111110",
  32729=>"11111100",
  32730=>"11111111",
  32731=>"11111100",
  32732=>"00000010",
  32733=>"00000000",
  32734=>"00000011",
  32735=>"00000011",
  32736=>"11111110",
  32737=>"00000000",
  32738=>"11111110",
  32739=>"00000011",
  32740=>"00000001",
  32741=>"00000010",
  32742=>"00000000",
  32743=>"11111110",
  32744=>"00000010",
  32745=>"11111111",
  32746=>"00000100",
  32747=>"00000000",
  32748=>"00000101",
  32749=>"00000010",
  32750=>"00000010",
  32751=>"11111111",
  32752=>"00000010",
  32753=>"11111111",
  32754=>"11111101",
  32755=>"11111101",
  32756=>"11111111",
  32757=>"00000010",
  32758=>"11111101",
  32759=>"00000001",
  32760=>"00000010",
  32761=>"11111111",
  32762=>"00000000",
  32763=>"00000100",
  32764=>"00000000",
  32765=>"11111111",
  32766=>"11111111",
  32767=>"00000100",
  32768=>"00000110",
  32769=>"11111111",
  32770=>"00000011",
  32771=>"00000000",
  32772=>"11111110",
  32773=>"11111101",
  32774=>"00000011",
  32775=>"11111110",
  32776=>"00000010",
  32777=>"00000000",
  32778=>"00000010",
  32779=>"00000000",
  32780=>"00000011",
  32781=>"00000101",
  32782=>"00000001",
  32783=>"11111111",
  32784=>"00000110",
  32785=>"11111100",
  32786=>"11111110",
  32787=>"11111111",
  32788=>"00000011",
  32789=>"11111111",
  32790=>"00000101",
  32791=>"00000100",
  32792=>"00000000",
  32793=>"11111110",
  32794=>"00000001",
  32795=>"11111110",
  32796=>"11111101",
  32797=>"00000010",
  32798=>"11111101",
  32799=>"00000011",
  32800=>"11111110",
  32801=>"00000100",
  32802=>"00000010",
  32803=>"00000000",
  32804=>"11111101",
  32805=>"11111111",
  32806=>"00000001",
  32807=>"00000010",
  32808=>"11111110",
  32809=>"11111110",
  32810=>"11111111",
  32811=>"00000001",
  32812=>"11111110",
  32813=>"11111111",
  32814=>"11111101",
  32815=>"11111110",
  32816=>"11111111",
  32817=>"11111111",
  32818=>"00000000",
  32819=>"11111110",
  32820=>"00000001",
  32821=>"00000001",
  32822=>"11111110",
  32823=>"00000001",
  32824=>"11111100",
  32825=>"00000001",
  32826=>"00000010",
  32827=>"11111110",
  32828=>"00000000",
  32829=>"00000010",
  32830=>"11111100",
  32831=>"11111101",
  32832=>"00000010",
  32833=>"00000001",
  32834=>"00000011",
  32835=>"11111110",
  32836=>"00000100",
  32837=>"00000001",
  32838=>"00000101",
  32839=>"00000100",
  32840=>"11111110",
  32841=>"11111110",
  32842=>"00000001",
  32843=>"00000000",
  32844=>"00000011",
  32845=>"00000001",
  32846=>"00000001",
  32847=>"11111101",
  32848=>"11111100",
  32849=>"00000000",
  32850=>"11111110",
  32851=>"00000010",
  32852=>"00000001",
  32853=>"00000001",
  32854=>"11111111",
  32855=>"00000010",
  32856=>"00000101",
  32857=>"00000100",
  32858=>"00000010",
  32859=>"00000010",
  32860=>"00000011",
  32861=>"00000011",
  32862=>"00000001",
  32863=>"00000011",
  32864=>"11111111",
  32865=>"11111110",
  32866=>"00000000",
  32867=>"11111110",
  32868=>"11111100",
  32869=>"00000000",
  32870=>"11111101",
  32871=>"11111110",
  32872=>"00000101",
  32873=>"11111101",
  32874=>"00000101",
  32875=>"00000000",
  32876=>"00000010",
  32877=>"11111111",
  32878=>"00000001",
  32879=>"00000110",
  32880=>"00000011",
  32881=>"00000010",
  32882=>"00000011",
  32883=>"00000010",
  32884=>"11111110",
  32885=>"00000101",
  32886=>"11111111",
  32887=>"11111101",
  32888=>"00000011",
  32889=>"11111111",
  32890=>"00000000",
  32891=>"00000010",
  32892=>"11111111",
  32893=>"11111111",
  32894=>"11111111",
  32895=>"11111111",
  32896=>"00000011",
  32897=>"00000001",
  32898=>"00000010",
  32899=>"00000001",
  32900=>"11111111",
  32901=>"11111110",
  32902=>"11111110",
  32903=>"11111110",
  32904=>"11111101",
  32905=>"00000011",
  32906=>"00000001",
  32907=>"11111100",
  32908=>"11111110",
  32909=>"11111110",
  32910=>"11111101",
  32911=>"11111110",
  32912=>"00000001",
  32913=>"00000010",
  32914=>"00000011",
  32915=>"11111101",
  32916=>"00000010",
  32917=>"11111111",
  32918=>"11111101",
  32919=>"00000001",
  32920=>"00000100",
  32921=>"00000110",
  32922=>"00000001",
  32923=>"11111101",
  32924=>"11111111",
  32925=>"00000000",
  32926=>"00000001",
  32927=>"00000001",
  32928=>"00000000",
  32929=>"00000011",
  32930=>"00000101",
  32931=>"11111100",
  32932=>"00000010",
  32933=>"00000100",
  32934=>"11111101",
  32935=>"11111110",
  32936=>"00000100",
  32937=>"11111110",
  32938=>"11111101",
  32939=>"11111110",
  32940=>"11111111",
  32941=>"11111111",
  32942=>"11111110",
  32943=>"00000010",
  32944=>"11111110",
  32945=>"11111110",
  32946=>"00000000",
  32947=>"00000001",
  32948=>"11111111",
  32949=>"11111111",
  32950=>"00000001",
  32951=>"11111110",
  32952=>"00000000",
  32953=>"00000001",
  32954=>"11111111",
  32955=>"00000010",
  32956=>"00000101",
  32957=>"11111110",
  32958=>"00000001",
  32959=>"00000001",
  32960=>"00000010",
  32961=>"11111111",
  32962=>"00000001",
  32963=>"11111111",
  32964=>"11111110",
  32965=>"00000101",
  32966=>"11111100",
  32967=>"00000010",
  32968=>"11111101",
  32969=>"11111101",
  32970=>"11111101",
  32971=>"11111110",
  32972=>"00000010",
  32973=>"00000001",
  32974=>"00000000",
  32975=>"00000001",
  32976=>"00000001",
  32977=>"11111100",
  32978=>"00000001",
  32979=>"00000001",
  32980=>"00000001",
  32981=>"11111110",
  32982=>"11111101",
  32983=>"11111110",
  32984=>"11111110",
  32985=>"11111111",
  32986=>"00000010",
  32987=>"11111011",
  32988=>"00000001",
  32989=>"00000000",
  32990=>"00000000",
  32991=>"11111110",
  32992=>"00000011",
  32993=>"00000101",
  32994=>"00000000",
  32995=>"00000101",
  32996=>"00000011",
  32997=>"11111111",
  32998=>"00000011",
  32999=>"00000011",
  33000=>"00000001",
  33001=>"00000110",
  33002=>"11111110",
  33003=>"11111111",
  33004=>"00000000",
  33005=>"00000011",
  33006=>"11111101",
  33007=>"11111111",
  33008=>"11111110",
  33009=>"00000011",
  33010=>"00000010",
  33011=>"00000001",
  33012=>"11111101",
  33013=>"11111100",
  33014=>"11111100",
  33015=>"11111111",
  33016=>"11111111",
  33017=>"00000011",
  33018=>"11111111",
  33019=>"11111110",
  33020=>"11111111",
  33021=>"00000000",
  33022=>"00000000",
  33023=>"11111111",
  33024=>"00000010",
  33025=>"11111101",
  33026=>"00000010",
  33027=>"00000001",
  33028=>"11111111",
  33029=>"11111110",
  33030=>"11111111",
  33031=>"11111110",
  33032=>"11111110",
  33033=>"00000100",
  33034=>"11111101",
  33035=>"00000010",
  33036=>"00000100",
  33037=>"11111111",
  33038=>"11111100",
  33039=>"11111100",
  33040=>"11111111",
  33041=>"11111100",
  33042=>"00000100",
  33043=>"11111111",
  33044=>"11111100",
  33045=>"00000110",
  33046=>"00000110",
  33047=>"00000000",
  33048=>"00000101",
  33049=>"11111110",
  33050=>"00000001",
  33051=>"11111111",
  33052=>"11111101",
  33053=>"00000001",
  33054=>"00000010",
  33055=>"00000111",
  33056=>"00000000",
  33057=>"11111101",
  33058=>"00000000",
  33059=>"00000010",
  33060=>"11111110",
  33061=>"11111101",
  33062=>"00000110",
  33063=>"00000000",
  33064=>"11111110",
  33065=>"11111101",
  33066=>"11111111",
  33067=>"11111110",
  33068=>"11111111",
  33069=>"00000000",
  33070=>"11111110",
  33071=>"00000010",
  33072=>"00000010",
  33073=>"11111111",
  33074=>"11111110",
  33075=>"00000101",
  33076=>"11111101",
  33077=>"11111100",
  33078=>"00000000",
  33079=>"00000011",
  33080=>"11111111",
  33081=>"00000000",
  33082=>"11111111",
  33083=>"00000001",
  33084=>"00000011",
  33085=>"11111110",
  33086=>"00000001",
  33087=>"11111111",
  33088=>"11111110",
  33089=>"11111111",
  33090=>"11111110",
  33091=>"00000001",
  33092=>"00000000",
  33093=>"00000100",
  33094=>"11111100",
  33095=>"00000001",
  33096=>"11111110",
  33097=>"00000001",
  33098=>"11111100",
  33099=>"00000011",
  33100=>"11111110",
  33101=>"11111110",
  33102=>"00000001",
  33103=>"00000100",
  33104=>"11111110",
  33105=>"11111101",
  33106=>"00000000",
  33107=>"00000011",
  33108=>"11111110",
  33109=>"11111111",
  33110=>"00000011",
  33111=>"00000011",
  33112=>"00000000",
  33113=>"11111101",
  33114=>"11111111",
  33115=>"11111111",
  33116=>"11111110",
  33117=>"11111110",
  33118=>"00000010",
  33119=>"00000000",
  33120=>"00000000",
  33121=>"00000001",
  33122=>"11111110",
  33123=>"00000011",
  33124=>"00000001",
  33125=>"00000000",
  33126=>"00000001",
  33127=>"00000100",
  33128=>"11111101",
  33129=>"00000001",
  33130=>"00000001",
  33131=>"11111110",
  33132=>"11111100",
  33133=>"00000000",
  33134=>"11111110",
  33135=>"11111111",
  33136=>"11111111",
  33137=>"11111100",
  33138=>"11111100",
  33139=>"00000010",
  33140=>"00000001",
  33141=>"00000110",
  33142=>"00000001",
  33143=>"11111111",
  33144=>"00000011",
  33145=>"11111101",
  33146=>"00000001",
  33147=>"11111100",
  33148=>"11111111",
  33149=>"00000001",
  33150=>"00000000",
  33151=>"11111111",
  33152=>"00000001",
  33153=>"11111111",
  33154=>"11111111",
  33155=>"11111101",
  33156=>"00000011",
  33157=>"11111101",
  33158=>"11111101",
  33159=>"11111011",
  33160=>"00000010",
  33161=>"00000011",
  33162=>"11111110",
  33163=>"00000001",
  33164=>"11111110",
  33165=>"11111111",
  33166=>"00000000",
  33167=>"00000011",
  33168=>"00000000",
  33169=>"00000010",
  33170=>"00000001",
  33171=>"11111101",
  33172=>"00000001",
  33173=>"11111100",
  33174=>"11111110",
  33175=>"11111110",
  33176=>"11111110",
  33177=>"11111110",
  33178=>"00000001",
  33179=>"11111111",
  33180=>"11111101",
  33181=>"00000010",
  33182=>"00000000",
  33183=>"00000001",
  33184=>"00000000",
  33185=>"00000000",
  33186=>"00000011",
  33187=>"11111110",
  33188=>"00000000",
  33189=>"00000011",
  33190=>"00000001",
  33191=>"00000001",
  33192=>"00000001",
  33193=>"00000110",
  33194=>"00000001",
  33195=>"11111110",
  33196=>"11111110",
  33197=>"11111100",
  33198=>"00000001",
  33199=>"00000010",
  33200=>"00000011",
  33201=>"11111101",
  33202=>"00000001",
  33203=>"11111101",
  33204=>"11111110",
  33205=>"11111111",
  33206=>"00000101",
  33207=>"00000111",
  33208=>"00000100",
  33209=>"11111110",
  33210=>"11111101",
  33211=>"11111100",
  33212=>"11111101",
  33213=>"11111110",
  33214=>"00000001",
  33215=>"00000000",
  33216=>"00000011",
  33217=>"00000000",
  33218=>"00000101",
  33219=>"00000011",
  33220=>"11111110",
  33221=>"11111110",
  33222=>"11111111",
  33223=>"11111101",
  33224=>"00000100",
  33225=>"00000100",
  33226=>"11111111",
  33227=>"11111111",
  33228=>"00000000",
  33229=>"11111101",
  33230=>"11111101",
  33231=>"11111111",
  33232=>"11111110",
  33233=>"00000011",
  33234=>"00000000",
  33235=>"00000001",
  33236=>"11111101",
  33237=>"11111110",
  33238=>"11111101",
  33239=>"00000001",
  33240=>"00000000",
  33241=>"00000000",
  33242=>"00000010",
  33243=>"00000000",
  33244=>"00000000",
  33245=>"00000001",
  33246=>"11111101",
  33247=>"00000001",
  33248=>"11111110",
  33249=>"00000101",
  33250=>"11111110",
  33251=>"00000001",
  33252=>"11111101",
  33253=>"11111111",
  33254=>"00000000",
  33255=>"00000010",
  33256=>"11111100",
  33257=>"00000010",
  33258=>"11111101",
  33259=>"00000101",
  33260=>"00000100",
  33261=>"11111101",
  33262=>"11111110",
  33263=>"11111100",
  33264=>"11111110",
  33265=>"11111011",
  33266=>"00000010",
  33267=>"11111101",
  33268=>"00000001",
  33269=>"11111101",
  33270=>"00000011",
  33271=>"11111101",
  33272=>"00000100",
  33273=>"00000101",
  33274=>"00000001",
  33275=>"11111111",
  33276=>"00000001",
  33277=>"00000000",
  33278=>"00000001",
  33279=>"00000110",
  33280=>"11111111",
  33281=>"00000011",
  33282=>"11111110",
  33283=>"00000000",
  33284=>"11111111",
  33285=>"00000011",
  33286=>"00000000",
  33287=>"00000010",
  33288=>"00000001",
  33289=>"00000000",
  33290=>"11111111",
  33291=>"00000010",
  33292=>"00000011",
  33293=>"00000001",
  33294=>"11111100",
  33295=>"00000100",
  33296=>"00000001",
  33297=>"00000010",
  33298=>"11111101",
  33299=>"11111100",
  33300=>"11111100",
  33301=>"00000011",
  33302=>"11111110",
  33303=>"11111111",
  33304=>"00000011",
  33305=>"00000101",
  33306=>"00000001",
  33307=>"00000010",
  33308=>"11111111",
  33309=>"00000000",
  33310=>"11111110",
  33311=>"00000100",
  33312=>"00000010",
  33313=>"00000001",
  33314=>"11111110",
  33315=>"11111101",
  33316=>"11111101",
  33317=>"00000001",
  33318=>"00000000",
  33319=>"11111110",
  33320=>"11111110",
  33321=>"00000010",
  33322=>"11111010",
  33323=>"11111101",
  33324=>"00000010",
  33325=>"11111110",
  33326=>"11111101",
  33327=>"11111110",
  33328=>"11111101",
  33329=>"11111101",
  33330=>"00000001",
  33331=>"11111100",
  33332=>"11111110",
  33333=>"00000011",
  33334=>"00000011",
  33335=>"11111100",
  33336=>"00000001",
  33337=>"00000000",
  33338=>"00000001",
  33339=>"11111100",
  33340=>"11111101",
  33341=>"00000000",
  33342=>"11111101",
  33343=>"00000010",
  33344=>"11111111",
  33345=>"00000001",
  33346=>"00000111",
  33347=>"11111111",
  33348=>"00000000",
  33349=>"11111111",
  33350=>"00000010",
  33351=>"00000011",
  33352=>"11111111",
  33353=>"00000001",
  33354=>"11111101",
  33355=>"11111101",
  33356=>"11111101",
  33357=>"11111110",
  33358=>"00000000",
  33359=>"11111110",
  33360=>"11111111",
  33361=>"00000000",
  33362=>"11111110",
  33363=>"11111111",
  33364=>"11111101",
  33365=>"11111101",
  33366=>"11111110",
  33367=>"11111100",
  33368=>"00000001",
  33369=>"00000011",
  33370=>"11111111",
  33371=>"00000010",
  33372=>"00000001",
  33373=>"00000000",
  33374=>"00000010",
  33375=>"00000011",
  33376=>"11111101",
  33377=>"00000011",
  33378=>"11111111",
  33379=>"00000010",
  33380=>"11111101",
  33381=>"11111111",
  33382=>"11111111",
  33383=>"00000001",
  33384=>"11111101",
  33385=>"00000010",
  33386=>"00000001",
  33387=>"11111111",
  33388=>"00000011",
  33389=>"00000001",
  33390=>"11111110",
  33391=>"00000001",
  33392=>"00000011",
  33393=>"00000001",
  33394=>"11111111",
  33395=>"00000010",
  33396=>"00000010",
  33397=>"00000000",
  33398=>"00000010",
  33399=>"11111110",
  33400=>"00000001",
  33401=>"11111101",
  33402=>"11111101",
  33403=>"11111110",
  33404=>"00000001",
  33405=>"11111101",
  33406=>"11111101",
  33407=>"00000010",
  33408=>"00000010",
  33409=>"11111111",
  33410=>"11111111",
  33411=>"11111101",
  33412=>"00000011",
  33413=>"00000101",
  33414=>"00000000",
  33415=>"00000011",
  33416=>"11111101",
  33417=>"00000000",
  33418=>"11111100",
  33419=>"00000111",
  33420=>"00000010",
  33421=>"00000000",
  33422=>"00000100",
  33423=>"00000000",
  33424=>"11111101",
  33425=>"11111110",
  33426=>"11111111",
  33427=>"00000001",
  33428=>"00000110",
  33429=>"11111101",
  33430=>"11111111",
  33431=>"00000010",
  33432=>"11111101",
  33433=>"00000010",
  33434=>"00000110",
  33435=>"00000010",
  33436=>"00000001",
  33437=>"11111100",
  33438=>"00000010",
  33439=>"00000000",
  33440=>"00000000",
  33441=>"00000110",
  33442=>"00000001",
  33443=>"11111101",
  33444=>"00000000",
  33445=>"11111110",
  33446=>"11111111",
  33447=>"00000010",
  33448=>"00000001",
  33449=>"11111110",
  33450=>"00000100",
  33451=>"11111110",
  33452=>"00000011",
  33453=>"00000100",
  33454=>"00000001",
  33455=>"00000011",
  33456=>"00000100",
  33457=>"00000001",
  33458=>"00000001",
  33459=>"00000001",
  33460=>"00000010",
  33461=>"00000010",
  33462=>"11111111",
  33463=>"11111101",
  33464=>"00000000",
  33465=>"11111111",
  33466=>"11111110",
  33467=>"11111110",
  33468=>"11111110",
  33469=>"00000001",
  33470=>"00000010",
  33471=>"00000010",
  33472=>"11111110",
  33473=>"11111111",
  33474=>"11111110",
  33475=>"00000000",
  33476=>"00000010",
  33477=>"11111111",
  33478=>"00000000",
  33479=>"00000010",
  33480=>"00000101",
  33481=>"11111110",
  33482=>"00000011",
  33483=>"00000010",
  33484=>"00000100",
  33485=>"00000010",
  33486=>"00000000",
  33487=>"00000001",
  33488=>"00000000",
  33489=>"00000000",
  33490=>"00000001",
  33491=>"11111110",
  33492=>"00000000",
  33493=>"00000011",
  33494=>"00000001",
  33495=>"11111101",
  33496=>"11111110",
  33497=>"00000001",
  33498=>"11111111",
  33499=>"11111111",
  33500=>"11111110",
  33501=>"11111110",
  33502=>"11111111",
  33503=>"11111111",
  33504=>"11111011",
  33505=>"00000000",
  33506=>"00000000",
  33507=>"00000011",
  33508=>"11111110",
  33509=>"00000100",
  33510=>"11111110",
  33511=>"11111101",
  33512=>"11111101",
  33513=>"11111110",
  33514=>"00000011",
  33515=>"00000010",
  33516=>"00000010",
  33517=>"00000000",
  33518=>"00000000",
  33519=>"11111110",
  33520=>"11111101",
  33521=>"11111110",
  33522=>"00000001",
  33523=>"00000000",
  33524=>"11111101",
  33525=>"00000010",
  33526=>"00000010",
  33527=>"00000000",
  33528=>"11111111",
  33529=>"00000100",
  33530=>"00000101",
  33531=>"11111111",
  33532=>"11111111",
  33533=>"11111110",
  33534=>"11111011",
  33535=>"00000000",
  33536=>"00000011",
  33537=>"00000011",
  33538=>"11111101",
  33539=>"11111100",
  33540=>"11111101",
  33541=>"00000000",
  33542=>"11111110",
  33543=>"11111101",
  33544=>"00000100",
  33545=>"11111100",
  33546=>"11111110",
  33547=>"00000001",
  33548=>"00000001",
  33549=>"00000001",
  33550=>"11111101",
  33551=>"00000010",
  33552=>"00000100",
  33553=>"00000110",
  33554=>"00000000",
  33555=>"11111110",
  33556=>"00000000",
  33557=>"00000101",
  33558=>"00000000",
  33559=>"00000011",
  33560=>"00000001",
  33561=>"00000001",
  33562=>"11111111",
  33563=>"11111100",
  33564=>"00000010",
  33565=>"00000001",
  33566=>"00000000",
  33567=>"00000001",
  33568=>"11111100",
  33569=>"00000001",
  33570=>"00000010",
  33571=>"00000000",
  33572=>"11111110",
  33573=>"00000010",
  33574=>"00000001",
  33575=>"11111110",
  33576=>"00000010",
  33577=>"00000000",
  33578=>"00000101",
  33579=>"00000011",
  33580=>"00000000",
  33581=>"00000101",
  33582=>"00000000",
  33583=>"11111111",
  33584=>"00000011",
  33585=>"00000000",
  33586=>"11111111",
  33587=>"00000000",
  33588=>"11111111",
  33589=>"11111111",
  33590=>"00000000",
  33591=>"11111110",
  33592=>"11111110",
  33593=>"11111111",
  33594=>"11111110",
  33595=>"00000110",
  33596=>"00000010",
  33597=>"00000011",
  33598=>"00000010",
  33599=>"11111100",
  33600=>"11111110",
  33601=>"00000001",
  33602=>"00000000",
  33603=>"00000000",
  33604=>"11111110",
  33605=>"11111101",
  33606=>"00000001",
  33607=>"11111110",
  33608=>"00000101",
  33609=>"00000001",
  33610=>"11111111",
  33611=>"00000010",
  33612=>"00000001",
  33613=>"00000001",
  33614=>"11111100",
  33615=>"00000001",
  33616=>"11111110",
  33617=>"00000010",
  33618=>"11111101",
  33619=>"00000001",
  33620=>"11111110",
  33621=>"00000010",
  33622=>"00000000",
  33623=>"11111111",
  33624=>"00000011",
  33625=>"00000010",
  33626=>"11111111",
  33627=>"00000100",
  33628=>"00000000",
  33629=>"11111100",
  33630=>"00000001",
  33631=>"00000100",
  33632=>"11111111",
  33633=>"00000011",
  33634=>"11111110",
  33635=>"00000101",
  33636=>"00000000",
  33637=>"11111110",
  33638=>"11111111",
  33639=>"11111111",
  33640=>"00000011",
  33641=>"00000000",
  33642=>"11111110",
  33643=>"00000100",
  33644=>"00000011",
  33645=>"11111101",
  33646=>"11111101",
  33647=>"11111101",
  33648=>"11111101",
  33649=>"11111110",
  33650=>"00000000",
  33651=>"11111110",
  33652=>"11111101",
  33653=>"11111011",
  33654=>"00000001",
  33655=>"11111101",
  33656=>"00000010",
  33657=>"00000111",
  33658=>"00000010",
  33659=>"11111110",
  33660=>"11111110",
  33661=>"00000001",
  33662=>"00000101",
  33663=>"00000000",
  33664=>"11111110",
  33665=>"11111101",
  33666=>"00000001",
  33667=>"00000010",
  33668=>"00000000",
  33669=>"00000100",
  33670=>"11111111",
  33671=>"11111111",
  33672=>"00000000",
  33673=>"00000001",
  33674=>"11111101",
  33675=>"00000000",
  33676=>"00000011",
  33677=>"11111101",
  33678=>"00000010",
  33679=>"00000001",
  33680=>"00000001",
  33681=>"11111101",
  33682=>"00000110",
  33683=>"00000001",
  33684=>"11111101",
  33685=>"00000000",
  33686=>"00000001",
  33687=>"11111110",
  33688=>"11111111",
  33689=>"00000000",
  33690=>"11111110",
  33691=>"00000100",
  33692=>"00000010",
  33693=>"00000000",
  33694=>"11111110",
  33695=>"00000011",
  33696=>"00000001",
  33697=>"00000001",
  33698=>"00000011",
  33699=>"00000000",
  33700=>"00000001",
  33701=>"11111100",
  33702=>"00000100",
  33703=>"11111101",
  33704=>"00000001",
  33705=>"00000001",
  33706=>"11111111",
  33707=>"11111111",
  33708=>"11111101",
  33709=>"11111110",
  33710=>"11111100",
  33711=>"00000010",
  33712=>"11111111",
  33713=>"00000010",
  33714=>"11111111",
  33715=>"11111111",
  33716=>"00000001",
  33717=>"11111110",
  33718=>"00000010",
  33719=>"11111110",
  33720=>"11111100",
  33721=>"00000011",
  33722=>"00000001",
  33723=>"00000010",
  33724=>"11111111",
  33725=>"00000101",
  33726=>"00000001",
  33727=>"11111101",
  33728=>"00000100",
  33729=>"11111110",
  33730=>"00000001",
  33731=>"11111111",
  33732=>"00000001",
  33733=>"11111111",
  33734=>"00000010",
  33735=>"11111111",
  33736=>"11111110",
  33737=>"11111101",
  33738=>"00000010",
  33739=>"11111111",
  33740=>"11111101",
  33741=>"11111111",
  33742=>"11111111",
  33743=>"11111111",
  33744=>"00000000",
  33745=>"00000001",
  33746=>"00000011",
  33747=>"11111101",
  33748=>"11111111",
  33749=>"00000001",
  33750=>"11111111",
  33751=>"00000000",
  33752=>"11111111",
  33753=>"11111101",
  33754=>"11111110",
  33755=>"00000010",
  33756=>"00000000",
  33757=>"00000001",
  33758=>"00000010",
  33759=>"00000001",
  33760=>"11111110",
  33761=>"11111110",
  33762=>"11111111",
  33763=>"00000010",
  33764=>"00000000",
  33765=>"00000100",
  33766=>"00000000",
  33767=>"00000011",
  33768=>"11111101",
  33769=>"00000001",
  33770=>"11111101",
  33771=>"11111111",
  33772=>"11111111",
  33773=>"00000001",
  33774=>"00000010",
  33775=>"00000011",
  33776=>"11111101",
  33777=>"00000010",
  33778=>"11111100",
  33779=>"11111111",
  33780=>"00000100",
  33781=>"11111111",
  33782=>"00000010",
  33783=>"11111110",
  33784=>"00000011",
  33785=>"00000011",
  33786=>"00000110",
  33787=>"00000010",
  33788=>"00000100",
  33789=>"00000111",
  33790=>"00000010",
  33791=>"11111101",
  33792=>"11111110",
  33793=>"11111101",
  33794=>"00000011",
  33795=>"00000011",
  33796=>"00000111",
  33797=>"11111100",
  33798=>"00000001",
  33799=>"11111110",
  33800=>"00000010",
  33801=>"00000010",
  33802=>"00000000",
  33803=>"11111101",
  33804=>"11111111",
  33805=>"11111101",
  33806=>"00000010",
  33807=>"11111111",
  33808=>"00000001",
  33809=>"11111100",
  33810=>"11111100",
  33811=>"00000000",
  33812=>"00000010",
  33813=>"00000011",
  33814=>"00000010",
  33815=>"11111110",
  33816=>"00000010",
  33817=>"00000010",
  33818=>"00000011",
  33819=>"00000000",
  33820=>"00000000",
  33821=>"00000001",
  33822=>"11111111",
  33823=>"00000011",
  33824=>"00000010",
  33825=>"00000000",
  33826=>"00000000",
  33827=>"00000001",
  33828=>"00000000",
  33829=>"11111111",
  33830=>"00000011",
  33831=>"11111111",
  33832=>"11111110",
  33833=>"11111110",
  33834=>"11111111",
  33835=>"00000000",
  33836=>"11111101",
  33837=>"00000000",
  33838=>"11111111",
  33839=>"00000011",
  33840=>"00000000",
  33841=>"11111110",
  33842=>"00000001",
  33843=>"11111110",
  33844=>"11111110",
  33845=>"00000001",
  33846=>"11111111",
  33847=>"00000100",
  33848=>"11111111",
  33849=>"11111101",
  33850=>"11111111",
  33851=>"00000011",
  33852=>"00000010",
  33853=>"11111111",
  33854=>"00000100",
  33855=>"00000010",
  33856=>"00000101",
  33857=>"00000000",
  33858=>"11111111",
  33859=>"00000000",
  33860=>"00000001",
  33861=>"11111110",
  33862=>"00000001",
  33863=>"11111100",
  33864=>"00000000",
  33865=>"11111110",
  33866=>"00000001",
  33867=>"00000010",
  33868=>"00000000",
  33869=>"00000110",
  33870=>"00000100",
  33871=>"11111110",
  33872=>"11111111",
  33873=>"00000000",
  33874=>"11111110",
  33875=>"11111110",
  33876=>"00000010",
  33877=>"11111110",
  33878=>"11111110",
  33879=>"11111110",
  33880=>"00000010",
  33881=>"00000011",
  33882=>"11111110",
  33883=>"00000000",
  33884=>"11111101",
  33885=>"00000110",
  33886=>"11111111",
  33887=>"11111100",
  33888=>"11111111",
  33889=>"00000001",
  33890=>"11111111",
  33891=>"00000000",
  33892=>"00001001",
  33893=>"11111111",
  33894=>"11111110",
  33895=>"00000000",
  33896=>"00000010",
  33897=>"11111111",
  33898=>"11111101",
  33899=>"11111110",
  33900=>"11111011",
  33901=>"11111101",
  33902=>"00000000",
  33903=>"11111111",
  33904=>"00000011",
  33905=>"00000010",
  33906=>"11111111",
  33907=>"00000000",
  33908=>"00000010",
  33909=>"00000001",
  33910=>"11111111",
  33911=>"11111101",
  33912=>"00000001",
  33913=>"00000000",
  33914=>"00000000",
  33915=>"00000101",
  33916=>"00000011",
  33917=>"00000101",
  33918=>"00000011",
  33919=>"11111101",
  33920=>"00000000",
  33921=>"00000001",
  33922=>"11111110",
  33923=>"00000000",
  33924=>"00000100",
  33925=>"00000001",
  33926=>"11111110",
  33927=>"11111110",
  33928=>"00000011",
  33929=>"00000000",
  33930=>"00000001",
  33931=>"00000100",
  33932=>"00000000",
  33933=>"11111110",
  33934=>"11111101",
  33935=>"11111011",
  33936=>"11111111",
  33937=>"00000001",
  33938=>"11111111",
  33939=>"00000100",
  33940=>"11111111",
  33941=>"00000001",
  33942=>"00000011",
  33943=>"11111110",
  33944=>"11111111",
  33945=>"11111111",
  33946=>"11111101",
  33947=>"11111100",
  33948=>"00000000",
  33949=>"00000110",
  33950=>"11111101",
  33951=>"00000100",
  33952=>"00000000",
  33953=>"11111111",
  33954=>"11111110",
  33955=>"11111101",
  33956=>"11111110",
  33957=>"00000001",
  33958=>"11111111",
  33959=>"00000001",
  33960=>"00000011",
  33961=>"11111110",
  33962=>"00000001",
  33963=>"00000000",
  33964=>"11111110",
  33965=>"00000011",
  33966=>"00000001",
  33967=>"00000000",
  33968=>"11111111",
  33969=>"00000001",
  33970=>"11111110",
  33971=>"00000101",
  33972=>"00000001",
  33973=>"11111101",
  33974=>"00000011",
  33975=>"11111101",
  33976=>"00000000",
  33977=>"11111110",
  33978=>"11111101",
  33979=>"00000000",
  33980=>"11111101",
  33981=>"11111110",
  33982=>"00000000",
  33983=>"11111111",
  33984=>"11111111",
  33985=>"00000010",
  33986=>"00000000",
  33987=>"00000000",
  33988=>"11111111",
  33989=>"00000110",
  33990=>"11111111",
  33991=>"11111111",
  33992=>"11111101",
  33993=>"11111101",
  33994=>"00000010",
  33995=>"00000000",
  33996=>"00000001",
  33997=>"11111101",
  33998=>"00000000",
  33999=>"11111101",
  34000=>"00000001",
  34001=>"00000000",
  34002=>"00000100",
  34003=>"00000000",
  34004=>"00000010",
  34005=>"00000000",
  34006=>"00000000",
  34007=>"11111100",
  34008=>"00000010",
  34009=>"00000001",
  34010=>"00000001",
  34011=>"11111100",
  34012=>"00000011",
  34013=>"11111111",
  34014=>"11111111",
  34015=>"11111111",
  34016=>"11111110",
  34017=>"00000011",
  34018=>"00000010",
  34019=>"00000001",
  34020=>"00000110",
  34021=>"11111110",
  34022=>"11111101",
  34023=>"11111110",
  34024=>"11111110",
  34025=>"00000010",
  34026=>"00000000",
  34027=>"11111110",
  34028=>"00000010",
  34029=>"11111100",
  34030=>"11111101",
  34031=>"00000010",
  34032=>"00000001",
  34033=>"11111110",
  34034=>"11111110",
  34035=>"00000010",
  34036=>"11111101",
  34037=>"00000011",
  34038=>"00000001",
  34039=>"00000011",
  34040=>"11111111",
  34041=>"11111111",
  34042=>"00000101",
  34043=>"11111111",
  34044=>"00000011",
  34045=>"11111110",
  34046=>"00000001",
  34047=>"11111110",
  34048=>"00000001",
  34049=>"00000000",
  34050=>"11111100",
  34051=>"00000010",
  34052=>"00000010",
  34053=>"11111101",
  34054=>"11111111",
  34055=>"11111101",
  34056=>"00000100",
  34057=>"11111110",
  34058=>"11111101",
  34059=>"00000001",
  34060=>"11111111",
  34061=>"00000001",
  34062=>"00000011",
  34063=>"00000010",
  34064=>"00000001",
  34065=>"00000000",
  34066=>"00000001",
  34067=>"00000001",
  34068=>"11111111",
  34069=>"11111100",
  34070=>"00000010",
  34071=>"00000011",
  34072=>"00000010",
  34073=>"00000000",
  34074=>"11111111",
  34075=>"00000001",
  34076=>"11111101",
  34077=>"11111101",
  34078=>"00000010",
  34079=>"00000000",
  34080=>"00000010",
  34081=>"00000101",
  34082=>"00000101",
  34083=>"00000011",
  34084=>"11111100",
  34085=>"11111111",
  34086=>"00000000",
  34087=>"00000001",
  34088=>"00000011",
  34089=>"00000011",
  34090=>"00000001",
  34091=>"00000100",
  34092=>"00000000",
  34093=>"11111101",
  34094=>"00000011",
  34095=>"11111101",
  34096=>"00000000",
  34097=>"11111110",
  34098=>"00000011",
  34099=>"11111101",
  34100=>"00000000",
  34101=>"00000000",
  34102=>"11111110",
  34103=>"11111101",
  34104=>"11111100",
  34105=>"11111111",
  34106=>"00000011",
  34107=>"11111110",
  34108=>"00000000",
  34109=>"00000010",
  34110=>"00000001",
  34111=>"11111111",
  34112=>"00000001",
  34113=>"00000001",
  34114=>"00000001",
  34115=>"00000010",
  34116=>"11111111",
  34117=>"00000000",
  34118=>"00000001",
  34119=>"00000010",
  34120=>"11111111",
  34121=>"11111110",
  34122=>"00000011",
  34123=>"00000011",
  34124=>"11111111",
  34125=>"00000010",
  34126=>"11111110",
  34127=>"11111100",
  34128=>"00000001",
  34129=>"00000011",
  34130=>"11111110",
  34131=>"11111111",
  34132=>"00000001",
  34133=>"11111111",
  34134=>"00000000",
  34135=>"00000000",
  34136=>"00000010",
  34137=>"11111110",
  34138=>"00000001",
  34139=>"11111101",
  34140=>"11111101",
  34141=>"00000001",
  34142=>"11111111",
  34143=>"00000000",
  34144=>"11111111",
  34145=>"11111100",
  34146=>"00000001",
  34147=>"00000010",
  34148=>"00000001",
  34149=>"11111110",
  34150=>"11111111",
  34151=>"11111110",
  34152=>"11111110",
  34153=>"00000000",
  34154=>"11111101",
  34155=>"00000000",
  34156=>"00000001",
  34157=>"00000000",
  34158=>"00000000",
  34159=>"00000001",
  34160=>"11111110",
  34161=>"00000011",
  34162=>"00000100",
  34163=>"00000000",
  34164=>"11111101",
  34165=>"11111111",
  34166=>"11111110",
  34167=>"00000001",
  34168=>"00000001",
  34169=>"00000011",
  34170=>"00000100",
  34171=>"00000000",
  34172=>"00000000",
  34173=>"11111110",
  34174=>"00000000",
  34175=>"00000011",
  34176=>"11111110",
  34177=>"11111100",
  34178=>"00000000",
  34179=>"00000110",
  34180=>"11111101",
  34181=>"11111101",
  34182=>"00000100",
  34183=>"11111110",
  34184=>"11111110",
  34185=>"00000110",
  34186=>"00000101",
  34187=>"00000100",
  34188=>"11111110",
  34189=>"00000011",
  34190=>"00000001",
  34191=>"11111110",
  34192=>"00000001",
  34193=>"00000000",
  34194=>"00000011",
  34195=>"00000010",
  34196=>"00000011",
  34197=>"11111110",
  34198=>"11111111",
  34199=>"00000001",
  34200=>"11111101",
  34201=>"11111101",
  34202=>"11111111",
  34203=>"00000011",
  34204=>"11111110",
  34205=>"11111101",
  34206=>"00000001",
  34207=>"00000001",
  34208=>"11111101",
  34209=>"11111101",
  34210=>"11111111",
  34211=>"11111101",
  34212=>"11111110",
  34213=>"11111110",
  34214=>"11111111",
  34215=>"11111110",
  34216=>"11111110",
  34217=>"00000000",
  34218=>"11111110",
  34219=>"00000000",
  34220=>"00000110",
  34221=>"00000110",
  34222=>"00000010",
  34223=>"00000000",
  34224=>"11111111",
  34225=>"00001000",
  34226=>"11111110",
  34227=>"11111110",
  34228=>"11111101",
  34229=>"00000000",
  34230=>"00000011",
  34231=>"11111101",
  34232=>"00000001",
  34233=>"00000000",
  34234=>"00000010",
  34235=>"11111110",
  34236=>"00000000",
  34237=>"11111111",
  34238=>"00000111",
  34239=>"00000000",
  34240=>"00000101",
  34241=>"00000000",
  34242=>"11111111",
  34243=>"00000101",
  34244=>"11111100",
  34245=>"11111101",
  34246=>"11111110",
  34247=>"11111111",
  34248=>"11111111",
  34249=>"00000001",
  34250=>"11111101",
  34251=>"11111111",
  34252=>"11111111",
  34253=>"11111111",
  34254=>"00000111",
  34255=>"00000100",
  34256=>"11111110",
  34257=>"11111111",
  34258=>"11111111",
  34259=>"11111100",
  34260=>"00000001",
  34261=>"11111111",
  34262=>"00000000",
  34263=>"00000001",
  34264=>"00000001",
  34265=>"11111101",
  34266=>"00000001",
  34267=>"11111101",
  34268=>"00000001",
  34269=>"00000011",
  34270=>"00000001",
  34271=>"00000000",
  34272=>"11111110",
  34273=>"11111111",
  34274=>"11111111",
  34275=>"00000000",
  34276=>"00000001",
  34277=>"11111111",
  34278=>"00000001",
  34279=>"11111110",
  34280=>"11111101",
  34281=>"11111101",
  34282=>"11111111",
  34283=>"00000100",
  34284=>"11111110",
  34285=>"00000010",
  34286=>"00000011",
  34287=>"11111101",
  34288=>"00000001",
  34289=>"00000111",
  34290=>"11111110",
  34291=>"11111111",
  34292=>"11111111",
  34293=>"00000001",
  34294=>"00000010",
  34295=>"00000101",
  34296=>"00000000",
  34297=>"11111111",
  34298=>"00000100",
  34299=>"11111110",
  34300=>"11111111",
  34301=>"00000010",
  34302=>"11111111",
  34303=>"11111111",
  34304=>"11111111",
  34305=>"00000000",
  34306=>"00000001",
  34307=>"00000010",
  34308=>"00000110",
  34309=>"00000011",
  34310=>"11111100",
  34311=>"00000011",
  34312=>"00000011",
  34313=>"00000001",
  34314=>"00000010",
  34315=>"00000011",
  34316=>"11111100",
  34317=>"11111111",
  34318=>"11111101",
  34319=>"00000000",
  34320=>"11111110",
  34321=>"11111110",
  34322=>"11111100",
  34323=>"11111110",
  34324=>"00000010",
  34325=>"00000010",
  34326=>"11111101",
  34327=>"11111110",
  34328=>"00000000",
  34329=>"11111101",
  34330=>"11111111",
  34331=>"11111111",
  34332=>"00000100",
  34333=>"00000010",
  34334=>"11111110",
  34335=>"11111101",
  34336=>"11111101",
  34337=>"00000101",
  34338=>"11111100",
  34339=>"00000001",
  34340=>"00000001",
  34341=>"11111101",
  34342=>"11111110",
  34343=>"11111110",
  34344=>"00000010",
  34345=>"00000011",
  34346=>"11111110",
  34347=>"00000011",
  34348=>"11111101",
  34349=>"00000000",
  34350=>"00000001",
  34351=>"11111111",
  34352=>"00000001",
  34353=>"00000010",
  34354=>"00000010",
  34355=>"00000010",
  34356=>"00000000",
  34357=>"00000001",
  34358=>"11111100",
  34359=>"00000001",
  34360=>"00000011",
  34361=>"00000001",
  34362=>"11111110",
  34363=>"00000010",
  34364=>"11111111",
  34365=>"11111110",
  34366=>"00000011",
  34367=>"00000010",
  34368=>"11111110",
  34369=>"00000011",
  34370=>"00000011",
  34371=>"00000001",
  34372=>"00000011",
  34373=>"11111111",
  34374=>"11111111",
  34375=>"00000010",
  34376=>"00000011",
  34377=>"00000001",
  34378=>"11111110",
  34379=>"11111110",
  34380=>"11111101",
  34381=>"00000010",
  34382=>"00000000",
  34383=>"11111110",
  34384=>"11111111",
  34385=>"11111101",
  34386=>"00000010",
  34387=>"00000000",
  34388=>"11111101",
  34389=>"00000001",
  34390=>"11111110",
  34391=>"00000011",
  34392=>"00000000",
  34393=>"11111111",
  34394=>"00000001",
  34395=>"00000001",
  34396=>"00000001",
  34397=>"00000001",
  34398=>"00000000",
  34399=>"00000010",
  34400=>"00000000",
  34401=>"00000001",
  34402=>"00000010",
  34403=>"11111111",
  34404=>"11111111",
  34405=>"11111101",
  34406=>"11111110",
  34407=>"00000000",
  34408=>"00000010",
  34409=>"00000000",
  34410=>"00000000",
  34411=>"11111111",
  34412=>"00000000",
  34413=>"11111101",
  34414=>"11111101",
  34415=>"00000010",
  34416=>"00000010",
  34417=>"00000100",
  34418=>"11111110",
  34419=>"00000000",
  34420=>"00000001",
  34421=>"11111110",
  34422=>"11111110",
  34423=>"11111100",
  34424=>"00000011",
  34425=>"00000011",
  34426=>"00000101",
  34427=>"00000000",
  34428=>"00000000",
  34429=>"11111111",
  34430=>"11111111",
  34431=>"11111110",
  34432=>"00000010",
  34433=>"11111110",
  34434=>"11111111",
  34435=>"11111110",
  34436=>"11111110",
  34437=>"00000000",
  34438=>"00000011",
  34439=>"11111111",
  34440=>"11111100",
  34441=>"11111111",
  34442=>"11111110",
  34443=>"11111111",
  34444=>"00000000",
  34445=>"00000010",
  34446=>"00000010",
  34447=>"00000001",
  34448=>"00000000",
  34449=>"11111101",
  34450=>"11111101",
  34451=>"00000000",
  34452=>"00000011",
  34453=>"11111110",
  34454=>"00000000",
  34455=>"00000010",
  34456=>"11111111",
  34457=>"11111110",
  34458=>"11111110",
  34459=>"00000100",
  34460=>"00000000",
  34461=>"11111111",
  34462=>"00000010",
  34463=>"11111101",
  34464=>"00000010",
  34465=>"11111110",
  34466=>"00000001",
  34467=>"00000000",
  34468=>"11111101",
  34469=>"00000111",
  34470=>"00000010",
  34471=>"11111111",
  34472=>"11111111",
  34473=>"00000010",
  34474=>"11111111",
  34475=>"00000000",
  34476=>"11111111",
  34477=>"00000001",
  34478=>"11111110",
  34479=>"11111101",
  34480=>"00000001",
  34481=>"00000001",
  34482=>"00000000",
  34483=>"00000001",
  34484=>"00000011",
  34485=>"00000100",
  34486=>"11111110",
  34487=>"11111101",
  34488=>"11111101",
  34489=>"11111111",
  34490=>"00000010",
  34491=>"00000010",
  34492=>"11111100",
  34493=>"00000000",
  34494=>"00000001",
  34495=>"00000010",
  34496=>"11111110",
  34497=>"11111110",
  34498=>"11111110",
  34499=>"11111110",
  34500=>"11111110",
  34501=>"00000000",
  34502=>"00000000",
  34503=>"11111111",
  34504=>"00000000",
  34505=>"00000010",
  34506=>"00000111",
  34507=>"00000011",
  34508=>"11111111",
  34509=>"11111111",
  34510=>"00000011",
  34511=>"11111110",
  34512=>"00000001",
  34513=>"11111110",
  34514=>"00000001",
  34515=>"11111111",
  34516=>"11111111",
  34517=>"11111101",
  34518=>"00000000",
  34519=>"11111110",
  34520=>"11111111",
  34521=>"00000000",
  34522=>"00000010",
  34523=>"00000000",
  34524=>"11111110",
  34525=>"00000011",
  34526=>"11111110",
  34527=>"11111101",
  34528=>"11111100",
  34529=>"00000000",
  34530=>"11111110",
  34531=>"11111101",
  34532=>"11111101",
  34533=>"11111111",
  34534=>"00000001",
  34535=>"00000000",
  34536=>"00000001",
  34537=>"00000010",
  34538=>"00000000",
  34539=>"11111101",
  34540=>"00000100",
  34541=>"11111111",
  34542=>"11111111",
  34543=>"11111111",
  34544=>"00000001",
  34545=>"11111111",
  34546=>"11111111",
  34547=>"00000010",
  34548=>"11111110",
  34549=>"00000001",
  34550=>"11111110",
  34551=>"11111111",
  34552=>"11111101",
  34553=>"11111100",
  34554=>"11111110",
  34555=>"11111100",
  34556=>"00000011",
  34557=>"00000011",
  34558=>"11111110",
  34559=>"00000001",
  34560=>"11111100",
  34561=>"11111111",
  34562=>"11111101",
  34563=>"11111110",
  34564=>"00000101",
  34565=>"00000000",
  34566=>"00000011",
  34567=>"11111111",
  34568=>"00000000",
  34569=>"11111110",
  34570=>"11111111",
  34571=>"11111111",
  34572=>"00000001",
  34573=>"00000100",
  34574=>"00000011",
  34575=>"00000000",
  34576=>"11111101",
  34577=>"11111110",
  34578=>"00000000",
  34579=>"11111111",
  34580=>"00000001",
  34581=>"00000000",
  34582=>"11111100",
  34583=>"00000000",
  34584=>"00000010",
  34585=>"11111101",
  34586=>"00000001",
  34587=>"11111111",
  34588=>"00000001",
  34589=>"00000001",
  34590=>"11111110",
  34591=>"00000001",
  34592=>"11111101",
  34593=>"11111110",
  34594=>"11111110",
  34595=>"11111110",
  34596=>"11111101",
  34597=>"00000011",
  34598=>"11111111",
  34599=>"00000000",
  34600=>"11111101",
  34601=>"00000011",
  34602=>"00000000",
  34603=>"00000011",
  34604=>"00000001",
  34605=>"11111111",
  34606=>"11111111",
  34607=>"00000010",
  34608=>"11111110",
  34609=>"00000011",
  34610=>"11111110",
  34611=>"11111111",
  34612=>"11111111",
  34613=>"11111101",
  34614=>"00000010",
  34615=>"00000011",
  34616=>"11111111",
  34617=>"00000001",
  34618=>"00000000",
  34619=>"11111110",
  34620=>"00000001",
  34621=>"00000001",
  34622=>"00000011",
  34623=>"00000001",
  34624=>"11111110",
  34625=>"00000011",
  34626=>"00000010",
  34627=>"11111100",
  34628=>"00000000",
  34629=>"11111111",
  34630=>"11111111",
  34631=>"00000100",
  34632=>"11111101",
  34633=>"00000100",
  34634=>"00000010",
  34635=>"00000011",
  34636=>"11111110",
  34637=>"11111101",
  34638=>"00000011",
  34639=>"11111111",
  34640=>"00000010",
  34641=>"00000011",
  34642=>"00000000",
  34643=>"11111111",
  34644=>"11111101",
  34645=>"11111110",
  34646=>"11111110",
  34647=>"11111111",
  34648=>"00000010",
  34649=>"00000011",
  34650=>"00000000",
  34651=>"11111101",
  34652=>"11111111",
  34653=>"11111111",
  34654=>"00000100",
  34655=>"11111111",
  34656=>"00000000",
  34657=>"11111111",
  34658=>"00000000",
  34659=>"11111101",
  34660=>"00000010",
  34661=>"00000010",
  34662=>"00000100",
  34663=>"00000010",
  34664=>"00000001",
  34665=>"00000011",
  34666=>"00000010",
  34667=>"00000010",
  34668=>"00000010",
  34669=>"11111111",
  34670=>"11111110",
  34671=>"00000001",
  34672=>"11111110",
  34673=>"00000001",
  34674=>"00000011",
  34675=>"11111110",
  34676=>"11111101",
  34677=>"11111111",
  34678=>"00000001",
  34679=>"00000100",
  34680=>"00000011",
  34681=>"11111110",
  34682=>"11111101",
  34683=>"11111101",
  34684=>"00000100",
  34685=>"00000001",
  34686=>"11111111",
  34687=>"11111101",
  34688=>"00000000",
  34689=>"00000010",
  34690=>"11111110",
  34691=>"11111101",
  34692=>"00000101",
  34693=>"11111110",
  34694=>"11111101",
  34695=>"11111111",
  34696=>"00000100",
  34697=>"00000111",
  34698=>"11111110",
  34699=>"00000001",
  34700=>"11111111",
  34701=>"11111101",
  34702=>"00000000",
  34703=>"00000000",
  34704=>"11111101",
  34705=>"00000001",
  34706=>"00000001",
  34707=>"11111101",
  34708=>"00000001",
  34709=>"00000000",
  34710=>"00000010",
  34711=>"11111110",
  34712=>"00000001",
  34713=>"00000011",
  34714=>"11111110",
  34715=>"11111111",
  34716=>"00000100",
  34717=>"00000010",
  34718=>"00000010",
  34719=>"11111100",
  34720=>"00000001",
  34721=>"00000101",
  34722=>"11111110",
  34723=>"11111111",
  34724=>"11111110",
  34725=>"11111111",
  34726=>"00000000",
  34727=>"11111110",
  34728=>"11111101",
  34729=>"00000010",
  34730=>"00000001",
  34731=>"11111110",
  34732=>"11111100",
  34733=>"11111110",
  34734=>"00000010",
  34735=>"11111101",
  34736=>"00000001",
  34737=>"11111111",
  34738=>"11111100",
  34739=>"11111110",
  34740=>"00000011",
  34741=>"00000010",
  34742=>"00000000",
  34743=>"00000001",
  34744=>"00000100",
  34745=>"00000010",
  34746=>"11111110",
  34747=>"00000001",
  34748=>"00000100",
  34749=>"11111100",
  34750=>"00000000",
  34751=>"11111111",
  34752=>"11111101",
  34753=>"00000001",
  34754=>"00000010",
  34755=>"11111110",
  34756=>"00000011",
  34757=>"00000010",
  34758=>"11111111",
  34759=>"00000011",
  34760=>"11111111",
  34761=>"11111101",
  34762=>"11111100",
  34763=>"00000000",
  34764=>"11111110",
  34765=>"00000010",
  34766=>"00000000",
  34767=>"00000001",
  34768=>"11111110",
  34769=>"00000100",
  34770=>"00000011",
  34771=>"11111110",
  34772=>"00000010",
  34773=>"11111110",
  34774=>"00000001",
  34775=>"00000000",
  34776=>"11111110",
  34777=>"11111101",
  34778=>"00000001",
  34779=>"00000110",
  34780=>"11111101",
  34781=>"11111111",
  34782=>"00000000",
  34783=>"11111101",
  34784=>"00000010",
  34785=>"11111111",
  34786=>"11111111",
  34787=>"00000000",
  34788=>"11111110",
  34789=>"00000001",
  34790=>"00000000",
  34791=>"00000101",
  34792=>"00000100",
  34793=>"00000000",
  34794=>"11111100",
  34795=>"11111110",
  34796=>"00000000",
  34797=>"00000001",
  34798=>"00000101",
  34799=>"11111110",
  34800=>"11111111",
  34801=>"00000010",
  34802=>"00000001",
  34803=>"11111111",
  34804=>"11111111",
  34805=>"11111110",
  34806=>"00000000",
  34807=>"11111110",
  34808=>"11111111",
  34809=>"11111111",
  34810=>"11111111",
  34811=>"11111110",
  34812=>"00000001",
  34813=>"00000010",
  34814=>"00000010",
  34815=>"11111111",
  34816=>"11111111",
  34817=>"00000111",
  34818=>"00000010",
  34819=>"00000000",
  34820=>"00000010",
  34821=>"11111110",
  34822=>"11111110",
  34823=>"00000010",
  34824=>"00000011",
  34825=>"11111111",
  34826=>"00000000",
  34827=>"11111100",
  34828=>"00000000",
  34829=>"00000011",
  34830=>"11111111",
  34831=>"11111100",
  34832=>"00000000",
  34833=>"00000100",
  34834=>"11111101",
  34835=>"00000010",
  34836=>"11111101",
  34837=>"00000010",
  34838=>"11111110",
  34839=>"00000001",
  34840=>"00000000",
  34841=>"00000010",
  34842=>"11111100",
  34843=>"00000100",
  34844=>"00000000",
  34845=>"00000010",
  34846=>"11111111",
  34847=>"00000011",
  34848=>"00000000",
  34849=>"11111110",
  34850=>"11111111",
  34851=>"00000000",
  34852=>"00000000",
  34853=>"00000010",
  34854=>"00000001",
  34855=>"11111110",
  34856=>"11111110",
  34857=>"11111111",
  34858=>"00000000",
  34859=>"00000010",
  34860=>"11111011",
  34861=>"00000000",
  34862=>"00000010",
  34863=>"00000000",
  34864=>"00000000",
  34865=>"11111110",
  34866=>"00000000",
  34867=>"00000011",
  34868=>"00000011",
  34869=>"00000011",
  34870=>"11111101",
  34871=>"11111101",
  34872=>"11111110",
  34873=>"11111110",
  34874=>"11111100",
  34875=>"00000001",
  34876=>"00000001",
  34877=>"11111111",
  34878=>"00000010",
  34879=>"00000000",
  34880=>"11111110",
  34881=>"00000100",
  34882=>"00000001",
  34883=>"00000011",
  34884=>"00000000",
  34885=>"00000001",
  34886=>"00000110",
  34887=>"00000010",
  34888=>"00000011",
  34889=>"11111100",
  34890=>"00000000",
  34891=>"00000010",
  34892=>"00000000",
  34893=>"11111111",
  34894=>"11111111",
  34895=>"11111110",
  34896=>"11111111",
  34897=>"00000100",
  34898=>"00000001",
  34899=>"00000001",
  34900=>"11111110",
  34901=>"00000011",
  34902=>"00000011",
  34903=>"00000000",
  34904=>"11111100",
  34905=>"00000100",
  34906=>"11111110",
  34907=>"00001010",
  34908=>"11111101",
  34909=>"11111111",
  34910=>"11111110",
  34911=>"11111111",
  34912=>"00000011",
  34913=>"11111101",
  34914=>"11111100",
  34915=>"11111110",
  34916=>"00000000",
  34917=>"00000011",
  34918=>"11111110",
  34919=>"11111111",
  34920=>"00000100",
  34921=>"00000001",
  34922=>"11111100",
  34923=>"00000011",
  34924=>"00000010",
  34925=>"00000000",
  34926=>"00000000",
  34927=>"11111101",
  34928=>"11111100",
  34929=>"00000001",
  34930=>"11111111",
  34931=>"11111110",
  34932=>"11111101",
  34933=>"11111110",
  34934=>"00000000",
  34935=>"11111101",
  34936=>"00000011",
  34937=>"00000001",
  34938=>"11111110",
  34939=>"11111101",
  34940=>"00000001",
  34941=>"11111111",
  34942=>"00000000",
  34943=>"11111100",
  34944=>"00000000",
  34945=>"11111110",
  34946=>"11111111",
  34947=>"11111100",
  34948=>"11111110",
  34949=>"00000001",
  34950=>"11111111",
  34951=>"11111111",
  34952=>"00000001",
  34953=>"00000000",
  34954=>"00000011",
  34955=>"11111110",
  34956=>"00000011",
  34957=>"00000001",
  34958=>"00000000",
  34959=>"00000100",
  34960=>"00000010",
  34961=>"11111100",
  34962=>"11111110",
  34963=>"11111101",
  34964=>"00000000",
  34965=>"00000100",
  34966=>"00000010",
  34967=>"11111111",
  34968=>"00000001",
  34969=>"11111111",
  34970=>"11111111",
  34971=>"11111101",
  34972=>"11111101",
  34973=>"00000011",
  34974=>"11111111",
  34975=>"00000010",
  34976=>"11111101",
  34977=>"00000000",
  34978=>"11111111",
  34979=>"00000001",
  34980=>"11111110",
  34981=>"00000010",
  34982=>"00000001",
  34983=>"00000000",
  34984=>"11111101",
  34985=>"00000010",
  34986=>"00000000",
  34987=>"11111100",
  34988=>"11111100",
  34989=>"11111100",
  34990=>"00000011",
  34991=>"00000010",
  34992=>"11111101",
  34993=>"11111110",
  34994=>"00000111",
  34995=>"11111111",
  34996=>"11111101",
  34997=>"11111101",
  34998=>"00000001",
  34999=>"00000001",
  35000=>"00000010",
  35001=>"00000110",
  35002=>"00000011",
  35003=>"00000011",
  35004=>"00000001",
  35005=>"11111110",
  35006=>"00000000",
  35007=>"00000110",
  35008=>"00000010",
  35009=>"00000011",
  35010=>"11111110",
  35011=>"00000100",
  35012=>"00000010",
  35013=>"11111101",
  35014=>"11111111",
  35015=>"11111101",
  35016=>"00000000",
  35017=>"00000011",
  35018=>"11111100",
  35019=>"00000010",
  35020=>"00000101",
  35021=>"11111101",
  35022=>"00000010",
  35023=>"00000010",
  35024=>"11111110",
  35025=>"00000010",
  35026=>"11111110",
  35027=>"11111111",
  35028=>"11111110",
  35029=>"00000100",
  35030=>"11111111",
  35031=>"00000010",
  35032=>"00000010",
  35033=>"00000111",
  35034=>"00000001",
  35035=>"11111111",
  35036=>"11111111",
  35037=>"11111100",
  35038=>"11111101",
  35039=>"00000011",
  35040=>"00000011",
  35041=>"11111111",
  35042=>"00000011",
  35043=>"00000011",
  35044=>"00000001",
  35045=>"11111110",
  35046=>"00000100",
  35047=>"11111110",
  35048=>"00000011",
  35049=>"00000011",
  35050=>"11111101",
  35051=>"00000001",
  35052=>"00000011",
  35053=>"00000011",
  35054=>"00000001",
  35055=>"11111110",
  35056=>"00000001",
  35057=>"00000100",
  35058=>"00000010",
  35059=>"11111111",
  35060=>"00000100",
  35061=>"11111110",
  35062=>"00000010",
  35063=>"00000010",
  35064=>"11111110",
  35065=>"11111110",
  35066=>"11111110",
  35067=>"00000000",
  35068=>"00000000",
  35069=>"00000000",
  35070=>"00000001",
  35071=>"11111110",
  35072=>"00000010",
  35073=>"11111111",
  35074=>"11111111",
  35075=>"11111111",
  35076=>"00000000",
  35077=>"00000100",
  35078=>"00000001",
  35079=>"11111111",
  35080=>"00000010",
  35081=>"00000010",
  35082=>"11111101",
  35083=>"00000010",
  35084=>"00000000",
  35085=>"00000001",
  35086=>"00000010",
  35087=>"11111100",
  35088=>"00000100",
  35089=>"11111110",
  35090=>"00000010",
  35091=>"00000001",
  35092=>"00000011",
  35093=>"11111111",
  35094=>"11111111",
  35095=>"11111100",
  35096=>"11111111",
  35097=>"11111111",
  35098=>"00000000",
  35099=>"00000001",
  35100=>"00000100",
  35101=>"00000100",
  35102=>"00000010",
  35103=>"00000011",
  35104=>"11111111",
  35105=>"11111101",
  35106=>"11111110",
  35107=>"00000010",
  35108=>"00000110",
  35109=>"00000111",
  35110=>"11111110",
  35111=>"00000011",
  35112=>"11111111",
  35113=>"00000001",
  35114=>"00000000",
  35115=>"11111011",
  35116=>"11111110",
  35117=>"11111111",
  35118=>"11111101",
  35119=>"00000011",
  35120=>"00000001",
  35121=>"00000011",
  35122=>"00000010",
  35123=>"11111111",
  35124=>"11111110",
  35125=>"00000100",
  35126=>"11111111",
  35127=>"00000010",
  35128=>"11111110",
  35129=>"00000101",
  35130=>"00000000",
  35131=>"11111110",
  35132=>"00000010",
  35133=>"11111111",
  35134=>"11111110",
  35135=>"11111101",
  35136=>"11111111",
  35137=>"00000000",
  35138=>"00000011",
  35139=>"11111111",
  35140=>"00000000",
  35141=>"00000011",
  35142=>"11111010",
  35143=>"11111101",
  35144=>"11111110",
  35145=>"11111111",
  35146=>"11111101",
  35147=>"11111111",
  35148=>"00000100",
  35149=>"11111110",
  35150=>"11111110",
  35151=>"00000011",
  35152=>"11111101",
  35153=>"00000011",
  35154=>"00000100",
  35155=>"11111110",
  35156=>"00000000",
  35157=>"11111111",
  35158=>"11111100",
  35159=>"11111100",
  35160=>"11111110",
  35161=>"11111110",
  35162=>"00000010",
  35163=>"11111101",
  35164=>"00000101",
  35165=>"00000010",
  35166=>"11111110",
  35167=>"00000000",
  35168=>"11111111",
  35169=>"11111100",
  35170=>"00000001",
  35171=>"00000010",
  35172=>"00000010",
  35173=>"00000001",
  35174=>"11111111",
  35175=>"11111110",
  35176=>"11111101",
  35177=>"11111101",
  35178=>"00000001",
  35179=>"00000010",
  35180=>"00000000",
  35181=>"00000011",
  35182=>"11111111",
  35183=>"00000010",
  35184=>"00000001",
  35185=>"00000000",
  35186=>"00000011",
  35187=>"11111100",
  35188=>"00000100",
  35189=>"00000011",
  35190=>"11111110",
  35191=>"11111110",
  35192=>"11111101",
  35193=>"00000010",
  35194=>"11111101",
  35195=>"11111111",
  35196=>"00000000",
  35197=>"00000001",
  35198=>"00000000",
  35199=>"00000010",
  35200=>"00000001",
  35201=>"00000000",
  35202=>"00000001",
  35203=>"00000001",
  35204=>"00000001",
  35205=>"00000010",
  35206=>"00000010",
  35207=>"00000100",
  35208=>"00000100",
  35209=>"11111111",
  35210=>"00000010",
  35211=>"00000001",
  35212=>"11111101",
  35213=>"11111111",
  35214=>"11111101",
  35215=>"00000001",
  35216=>"00000001",
  35217=>"11111101",
  35218=>"00000011",
  35219=>"00000011",
  35220=>"11111110",
  35221=>"11111100",
  35222=>"00000011",
  35223=>"00000001",
  35224=>"00000011",
  35225=>"11111011",
  35226=>"00000100",
  35227=>"11111101",
  35228=>"11111111",
  35229=>"11111111",
  35230=>"11111101",
  35231=>"11111110",
  35232=>"00000010",
  35233=>"00000010",
  35234=>"00000000",
  35235=>"00000000",
  35236=>"00000000",
  35237=>"11111110",
  35238=>"11111111",
  35239=>"00000000",
  35240=>"00000100",
  35241=>"11111111",
  35242=>"00000101",
  35243=>"00000011",
  35244=>"00000010",
  35245=>"11111101",
  35246=>"00000000",
  35247=>"11111111",
  35248=>"11111101",
  35249=>"11111111",
  35250=>"11111110",
  35251=>"11111101",
  35252=>"11111111",
  35253=>"11111101",
  35254=>"00000010",
  35255=>"11111110",
  35256=>"11111101",
  35257=>"00000010",
  35258=>"11111101",
  35259=>"00000001",
  35260=>"11111101",
  35261=>"11111111",
  35262=>"00000000",
  35263=>"00000001",
  35264=>"11111110",
  35265=>"11111110",
  35266=>"11111110",
  35267=>"00000000",
  35268=>"00000010",
  35269=>"00000001",
  35270=>"11111101",
  35271=>"00000000",
  35272=>"00000110",
  35273=>"00000011",
  35274=>"11111111",
  35275=>"00000000",
  35276=>"11111100",
  35277=>"00000010",
  35278=>"11111110",
  35279=>"11111110",
  35280=>"11111110",
  35281=>"11111111",
  35282=>"00000000",
  35283=>"00000000",
  35284=>"00000001",
  35285=>"11111110",
  35286=>"00000000",
  35287=>"00000000",
  35288=>"00000011",
  35289=>"00000011",
  35290=>"11111110",
  35291=>"11111100",
  35292=>"11111100",
  35293=>"00000001",
  35294=>"00000011",
  35295=>"11111111",
  35296=>"11111101",
  35297=>"11111011",
  35298=>"00000001",
  35299=>"00000010",
  35300=>"00000001",
  35301=>"00000001",
  35302=>"11111111",
  35303=>"00000001",
  35304=>"00000100",
  35305=>"00000100",
  35306=>"11111110",
  35307=>"00000100",
  35308=>"00000010",
  35309=>"00000000",
  35310=>"00000101",
  35311=>"00000011",
  35312=>"00000010",
  35313=>"11111110",
  35314=>"11111111",
  35315=>"11111111",
  35316=>"00000000",
  35317=>"00000101",
  35318=>"00000100",
  35319=>"00000000",
  35320=>"00000011",
  35321=>"00000010",
  35322=>"00000011",
  35323=>"00000001",
  35324=>"00000001",
  35325=>"11111111",
  35326=>"00000001",
  35327=>"00000000",
  35328=>"00000001",
  35329=>"00000000",
  35330=>"00000010",
  35331=>"00000010",
  35332=>"11111100",
  35333=>"00000010",
  35334=>"11111111",
  35335=>"00000010",
  35336=>"00000010",
  35337=>"00000001",
  35338=>"00000001",
  35339=>"00000000",
  35340=>"11111100",
  35341=>"00000000",
  35342=>"00000000",
  35343=>"11111101",
  35344=>"00000010",
  35345=>"00000001",
  35346=>"00000001",
  35347=>"11111110",
  35348=>"00000111",
  35349=>"11111111",
  35350=>"11111100",
  35351=>"11111111",
  35352=>"11111110",
  35353=>"00000001",
  35354=>"11111111",
  35355=>"00000001",
  35356=>"11111111",
  35357=>"11111110",
  35358=>"11111111",
  35359=>"11111110",
  35360=>"00000011",
  35361=>"00000000",
  35362=>"00000011",
  35363=>"11111101",
  35364=>"00000000",
  35365=>"00000011",
  35366=>"00000011",
  35367=>"11111110",
  35368=>"00000000",
  35369=>"00000000",
  35370=>"11111010",
  35371=>"00000011",
  35372=>"11111100",
  35373=>"00000000",
  35374=>"00000011",
  35375=>"00000101",
  35376=>"00000010",
  35377=>"11111111",
  35378=>"11111110",
  35379=>"00000000",
  35380=>"00000001",
  35381=>"11111111",
  35382=>"11111100",
  35383=>"00000001",
  35384=>"11111110",
  35385=>"00000000",
  35386=>"11111110",
  35387=>"00000001",
  35388=>"00000010",
  35389=>"11111111",
  35390=>"00000001",
  35391=>"00000100",
  35392=>"11111110",
  35393=>"11111101",
  35394=>"00000011",
  35395=>"00000111",
  35396=>"11111101",
  35397=>"00000011",
  35398=>"11111110",
  35399=>"00000010",
  35400=>"11111110",
  35401=>"11111100",
  35402=>"00000001",
  35403=>"00000000",
  35404=>"00000010",
  35405=>"11111101",
  35406=>"11111101",
  35407=>"11111101",
  35408=>"11111111",
  35409=>"11111101",
  35410=>"00000001",
  35411=>"00000010",
  35412=>"00000011",
  35413=>"00000011",
  35414=>"11111111",
  35415=>"11111100",
  35416=>"00000001",
  35417=>"00000011",
  35418=>"00000001",
  35419=>"00000000",
  35420=>"11111110",
  35421=>"11111110",
  35422=>"11111101",
  35423=>"11111111",
  35424=>"00000001",
  35425=>"00000010",
  35426=>"00000011",
  35427=>"00000011",
  35428=>"00000011",
  35429=>"00000101",
  35430=>"00000000",
  35431=>"11111110",
  35432=>"11111110",
  35433=>"00000100",
  35434=>"11111111",
  35435=>"00000000",
  35436=>"00000111",
  35437=>"11111110",
  35438=>"00000101",
  35439=>"11111110",
  35440=>"00000010",
  35441=>"00000001",
  35442=>"11111101",
  35443=>"00000101",
  35444=>"11111111",
  35445=>"00000001",
  35446=>"00000000",
  35447=>"11111100",
  35448=>"11111111",
  35449=>"11111101",
  35450=>"00000001",
  35451=>"11111111",
  35452=>"00000001",
  35453=>"00000110",
  35454=>"00000011",
  35455=>"11111110",
  35456=>"00000001",
  35457=>"00000010",
  35458=>"00000011",
  35459=>"11111111",
  35460=>"00000100",
  35461=>"00000000",
  35462=>"11111110",
  35463=>"00000001",
  35464=>"11111111",
  35465=>"00000000",
  35466=>"11111110",
  35467=>"00000001",
  35468=>"11111110",
  35469=>"11111110",
  35470=>"00000001",
  35471=>"00000001",
  35472=>"11111100",
  35473=>"00000011",
  35474=>"00000011",
  35475=>"00000000",
  35476=>"11111111",
  35477=>"11111110",
  35478=>"00000011",
  35479=>"00000101",
  35480=>"00000001",
  35481=>"11111111",
  35482=>"11111110",
  35483=>"00000010",
  35484=>"00000110",
  35485=>"11111110",
  35486=>"11111110",
  35487=>"00000001",
  35488=>"00000010",
  35489=>"11111110",
  35490=>"11111101",
  35491=>"11111111",
  35492=>"00000001",
  35493=>"11111111",
  35494=>"11111110",
  35495=>"11111101",
  35496=>"11111110",
  35497=>"00000011",
  35498=>"00000000",
  35499=>"00000000",
  35500=>"11111101",
  35501=>"11111101",
  35502=>"11111110",
  35503=>"11111101",
  35504=>"00000010",
  35505=>"00000001",
  35506=>"00000011",
  35507=>"11111110",
  35508=>"00000010",
  35509=>"11111111",
  35510=>"00000100",
  35511=>"11111110",
  35512=>"00000010",
  35513=>"11111110",
  35514=>"11111110",
  35515=>"00000000",
  35516=>"00000000",
  35517=>"11111111",
  35518=>"00000001",
  35519=>"11111101",
  35520=>"00000000",
  35521=>"11111111",
  35522=>"00000000",
  35523=>"11111100",
  35524=>"00000010",
  35525=>"00000010",
  35526=>"11111110",
  35527=>"00000100",
  35528=>"00000010",
  35529=>"00000000",
  35530=>"11111100",
  35531=>"00000010",
  35532=>"00000001",
  35533=>"11111100",
  35534=>"00000011",
  35535=>"00000011",
  35536=>"00000000",
  35537=>"00000001",
  35538=>"00000100",
  35539=>"11111111",
  35540=>"11111111",
  35541=>"00000101",
  35542=>"00000001",
  35543=>"11111110",
  35544=>"11111101",
  35545=>"00000011",
  35546=>"00000010",
  35547=>"11111111",
  35548=>"11111111",
  35549=>"11111111",
  35550=>"11111111",
  35551=>"00000100",
  35552=>"00000110",
  35553=>"00000010",
  35554=>"11111110",
  35555=>"00000001",
  35556=>"00000011",
  35557=>"11111111",
  35558=>"00000000",
  35559=>"00000000",
  35560=>"11111110",
  35561=>"11111110",
  35562=>"11111101",
  35563=>"11111101",
  35564=>"00000000",
  35565=>"11111100",
  35566=>"00000011",
  35567=>"11111101",
  35568=>"00000110",
  35569=>"00000000",
  35570=>"00000010",
  35571=>"11111110",
  35572=>"00000000",
  35573=>"00000010",
  35574=>"11111111",
  35575=>"11111111",
  35576=>"00000001",
  35577=>"11111111",
  35578=>"00000011",
  35579=>"00000100",
  35580=>"00000001",
  35581=>"11111101",
  35582=>"00000010",
  35583=>"00000001",
  35584=>"11111110",
  35585=>"11111101",
  35586=>"11111100",
  35587=>"00000011",
  35588=>"11111111",
  35589=>"00000001",
  35590=>"11111110",
  35591=>"00000011",
  35592=>"11111010",
  35593=>"11111110",
  35594=>"00000010",
  35595=>"00000010",
  35596=>"11111111",
  35597=>"00000000",
  35598=>"00000110",
  35599=>"11111110",
  35600=>"11111100",
  35601=>"00000010",
  35602=>"00000001",
  35603=>"00000000",
  35604=>"11111111",
  35605=>"00000000",
  35606=>"11111101",
  35607=>"00000101",
  35608=>"11111101",
  35609=>"11111100",
  35610=>"00000101",
  35611=>"00000100",
  35612=>"11111111",
  35613=>"11111111",
  35614=>"11111100",
  35615=>"00000000",
  35616=>"00000001",
  35617=>"11111110",
  35618=>"00000000",
  35619=>"00000100",
  35620=>"00000010",
  35621=>"00000011",
  35622=>"11111111",
  35623=>"00000000",
  35624=>"11111100",
  35625=>"11111111",
  35626=>"11111111",
  35627=>"11111101",
  35628=>"00000001",
  35629=>"11111111",
  35630=>"00000011",
  35631=>"00000111",
  35632=>"11111101",
  35633=>"11111101",
  35634=>"11111101",
  35635=>"11111111",
  35636=>"00000010",
  35637=>"00000001",
  35638=>"11111101",
  35639=>"00000011",
  35640=>"00000001",
  35641=>"11111111",
  35642=>"11111111",
  35643=>"00000100",
  35644=>"11111110",
  35645=>"00000001",
  35646=>"00000000",
  35647=>"00000000",
  35648=>"00000110",
  35649=>"00000011",
  35650=>"00000010",
  35651=>"00000001",
  35652=>"00000000",
  35653=>"11111111",
  35654=>"11111111",
  35655=>"00000010",
  35656=>"11111111",
  35657=>"00000011",
  35658=>"11111011",
  35659=>"11111111",
  35660=>"11111100",
  35661=>"00000010",
  35662=>"11111101",
  35663=>"11111110",
  35664=>"00000011",
  35665=>"00000000",
  35666=>"11111110",
  35667=>"00000011",
  35668=>"00000101",
  35669=>"11111111",
  35670=>"00000001",
  35671=>"00000001",
  35672=>"11111110",
  35673=>"11111100",
  35674=>"00000100",
  35675=>"11111101",
  35676=>"00000010",
  35677=>"00000010",
  35678=>"00000110",
  35679=>"00000000",
  35680=>"00000001",
  35681=>"00000000",
  35682=>"11111101",
  35683=>"00000000",
  35684=>"00000010",
  35685=>"00000001",
  35686=>"11111101",
  35687=>"11111110",
  35688=>"11111100",
  35689=>"11111101",
  35690=>"00000001",
  35691=>"11111111",
  35692=>"11111101",
  35693=>"11111101",
  35694=>"00000000",
  35695=>"00000100",
  35696=>"00000001",
  35697=>"00000010",
  35698=>"00000001",
  35699=>"00000100",
  35700=>"11111110",
  35701=>"11111110",
  35702=>"11111101",
  35703=>"11111111",
  35704=>"00000000",
  35705=>"00000000",
  35706=>"00000010",
  35707=>"11111100",
  35708=>"00000000",
  35709=>"11111110",
  35710=>"00000001",
  35711=>"00000000",
  35712=>"11111110",
  35713=>"00000100",
  35714=>"00000001",
  35715=>"00000110",
  35716=>"11111110",
  35717=>"00000011",
  35718=>"11111110",
  35719=>"00000010",
  35720=>"00000100",
  35721=>"11111101",
  35722=>"00000010",
  35723=>"00000010",
  35724=>"11111101",
  35725=>"11111110",
  35726=>"00000010",
  35727=>"00000001",
  35728=>"11111110",
  35729=>"00000001",
  35730=>"11111111",
  35731=>"11111111",
  35732=>"00000001",
  35733=>"11111110",
  35734=>"00000000",
  35735=>"11111110",
  35736=>"00000101",
  35737=>"11111101",
  35738=>"11111111",
  35739=>"11111110",
  35740=>"00000001",
  35741=>"00000010",
  35742=>"11111111",
  35743=>"00000011",
  35744=>"00000100",
  35745=>"11111111",
  35746=>"00000101",
  35747=>"11111110",
  35748=>"11111110",
  35749=>"11111110",
  35750=>"00000001",
  35751=>"11111101",
  35752=>"00000000",
  35753=>"00000001",
  35754=>"11111101",
  35755=>"11111101",
  35756=>"00000100",
  35757=>"11111101",
  35758=>"00000010",
  35759=>"11111101",
  35760=>"00000011",
  35761=>"11111110",
  35762=>"11111111",
  35763=>"00000001",
  35764=>"00000000",
  35765=>"11111101",
  35766=>"00000011",
  35767=>"11111111",
  35768=>"11111101",
  35769=>"11111111",
  35770=>"00000011",
  35771=>"11111100",
  35772=>"11111101",
  35773=>"11111101",
  35774=>"00000001",
  35775=>"11111101",
  35776=>"11111111",
  35777=>"00000010",
  35778=>"11111101",
  35779=>"00000100",
  35780=>"11111110",
  35781=>"00000001",
  35782=>"00000011",
  35783=>"00000001",
  35784=>"00000001",
  35785=>"11111101",
  35786=>"00000100",
  35787=>"11111110",
  35788=>"11111111",
  35789=>"00000001",
  35790=>"11111111",
  35791=>"11111101",
  35792=>"00000011",
  35793=>"00000001",
  35794=>"00000100",
  35795=>"11111111",
  35796=>"00000011",
  35797=>"00000100",
  35798=>"00000010",
  35799=>"11111111",
  35800=>"11111101",
  35801=>"11111101",
  35802=>"11111110",
  35803=>"11111110",
  35804=>"11111101",
  35805=>"11111101",
  35806=>"11111111",
  35807=>"00000100",
  35808=>"00000101",
  35809=>"00000001",
  35810=>"00000001",
  35811=>"00000011",
  35812=>"11111110",
  35813=>"00000001",
  35814=>"00000001",
  35815=>"00000011",
  35816=>"00000010",
  35817=>"00000001",
  35818=>"11111100",
  35819=>"00000000",
  35820=>"11111111",
  35821=>"00000001",
  35822=>"11111110",
  35823=>"11111101",
  35824=>"00000001",
  35825=>"11111101",
  35826=>"11111110",
  35827=>"11111110",
  35828=>"00000011",
  35829=>"00000010",
  35830=>"00000100",
  35831=>"00000110",
  35832=>"00000100",
  35833=>"00000011",
  35834=>"11111111",
  35835=>"11111101",
  35836=>"11111111",
  35837=>"00000001",
  35838=>"11111110",
  35839=>"11111101",
  35840=>"11111101",
  35841=>"00000000",
  35842=>"11111101",
  35843=>"11111111",
  35844=>"11111101",
  35845=>"00000100",
  35846=>"11111101",
  35847=>"11111100",
  35848=>"11111110",
  35849=>"11111110",
  35850=>"11111110",
  35851=>"00000000",
  35852=>"00000000",
  35853=>"11111111",
  35854=>"00000000",
  35855=>"11111101",
  35856=>"00000000",
  35857=>"00000101",
  35858=>"00000000",
  35859=>"00000011",
  35860=>"00000000",
  35861=>"11111110",
  35862=>"11111111",
  35863=>"00000001",
  35864=>"11111110",
  35865=>"00000001",
  35866=>"11111101",
  35867=>"11111111",
  35868=>"11111110",
  35869=>"11111101",
  35870=>"11111110",
  35871=>"11111110",
  35872=>"00000100",
  35873=>"11111111",
  35874=>"00000001",
  35875=>"11111101",
  35876=>"11111110",
  35877=>"00000011",
  35878=>"11111101",
  35879=>"00000001",
  35880=>"00000010",
  35881=>"11111110",
  35882=>"11111111",
  35883=>"00000000",
  35884=>"00000010",
  35885=>"00000010",
  35886=>"00000001",
  35887=>"11111111",
  35888=>"00000001",
  35889=>"00000000",
  35890=>"11111100",
  35891=>"00000001",
  35892=>"00000001",
  35893=>"00000000",
  35894=>"00000001",
  35895=>"00000001",
  35896=>"11111110",
  35897=>"00000000",
  35898=>"11111110",
  35899=>"11111110",
  35900=>"00000001",
  35901=>"00000010",
  35902=>"00000001",
  35903=>"00000001",
  35904=>"11111101",
  35905=>"11111110",
  35906=>"00000001",
  35907=>"00000000",
  35908=>"11111100",
  35909=>"00000010",
  35910=>"11111101",
  35911=>"00000101",
  35912=>"11111110",
  35913=>"11111110",
  35914=>"00000000",
  35915=>"11111101",
  35916=>"11111101",
  35917=>"00000000",
  35918=>"00000000",
  35919=>"00000010",
  35920=>"00000101",
  35921=>"00000000",
  35922=>"00000000",
  35923=>"00000000",
  35924=>"00000100",
  35925=>"11111101",
  35926=>"11111101",
  35927=>"11111101",
  35928=>"00000000",
  35929=>"11111110",
  35930=>"11111111",
  35931=>"11111111",
  35932=>"11111100",
  35933=>"11111101",
  35934=>"11111101",
  35935=>"11111110",
  35936=>"11111110",
  35937=>"00000010",
  35938=>"00000010",
  35939=>"00000010",
  35940=>"00000001",
  35941=>"00000011",
  35942=>"00000000",
  35943=>"00000000",
  35944=>"11111110",
  35945=>"00000010",
  35946=>"00000000",
  35947=>"11111110",
  35948=>"11111110",
  35949=>"11111100",
  35950=>"11111110",
  35951=>"11111101",
  35952=>"00000000",
  35953=>"00000010",
  35954=>"00000000",
  35955=>"00000010",
  35956=>"00000000",
  35957=>"00000001",
  35958=>"00000001",
  35959=>"00000001",
  35960=>"11111110",
  35961=>"11111100",
  35962=>"00000010",
  35963=>"11111110",
  35964=>"11111101",
  35965=>"00000010",
  35966=>"00000001",
  35967=>"11111110",
  35968=>"00000000",
  35969=>"00000010",
  35970=>"00000011",
  35971=>"11111101",
  35972=>"00000010",
  35973=>"00000011",
  35974=>"00000001",
  35975=>"00000010",
  35976=>"00000010",
  35977=>"00000000",
  35978=>"11111101",
  35979=>"11111100",
  35980=>"11111111",
  35981=>"11111111",
  35982=>"11111110",
  35983=>"11111101",
  35984=>"11111110",
  35985=>"00000000",
  35986=>"00000001",
  35987=>"11111101",
  35988=>"11111111",
  35989=>"00000000",
  35990=>"11111111",
  35991=>"00000000",
  35992=>"11111110",
  35993=>"11111110",
  35994=>"11111101",
  35995=>"00000011",
  35996=>"11111110",
  35997=>"00000011",
  35998=>"00000001",
  35999=>"00000011",
  36000=>"11111101",
  36001=>"11111110",
  36002=>"00000001",
  36003=>"00000010",
  36004=>"11111110",
  36005=>"11111111",
  36006=>"11111111",
  36007=>"11111101",
  36008=>"00000001",
  36009=>"00000000",
  36010=>"11111101",
  36011=>"11111101",
  36012=>"11111101",
  36013=>"11111110",
  36014=>"00000001",
  36015=>"11111111",
  36016=>"00000101",
  36017=>"11111110",
  36018=>"00000010",
  36019=>"11111111",
  36020=>"00000001",
  36021=>"00000001",
  36022=>"11111111",
  36023=>"00000010",
  36024=>"11111110",
  36025=>"11111101",
  36026=>"11111110",
  36027=>"11111111",
  36028=>"00000000",
  36029=>"00000011",
  36030=>"11111110",
  36031=>"00000100",
  36032=>"11111111",
  36033=>"00000010",
  36034=>"00000000",
  36035=>"00000001",
  36036=>"00000000",
  36037=>"00000000",
  36038=>"00000000",
  36039=>"11111101",
  36040=>"11111101",
  36041=>"11111111",
  36042=>"11111111",
  36043=>"11111111",
  36044=>"00000011",
  36045=>"00000001",
  36046=>"00000010",
  36047=>"00000001",
  36048=>"00000000",
  36049=>"11111110",
  36050=>"11111110",
  36051=>"11111110",
  36052=>"11111110",
  36053=>"11111101",
  36054=>"00000011",
  36055=>"11111110",
  36056=>"11111110",
  36057=>"11111110",
  36058=>"00000010",
  36059=>"00000101",
  36060=>"11111101",
  36061=>"00000001",
  36062=>"00000011",
  36063=>"11111111",
  36064=>"00000001",
  36065=>"00000000",
  36066=>"11111110",
  36067=>"11111110",
  36068=>"00000010",
  36069=>"00000000",
  36070=>"00000000",
  36071=>"00000011",
  36072=>"11111111",
  36073=>"00000001",
  36074=>"11111111",
  36075=>"11111110",
  36076=>"00000000",
  36077=>"00000011",
  36078=>"00000101",
  36079=>"11111111",
  36080=>"11111100",
  36081=>"11111110",
  36082=>"11111111",
  36083=>"11111110",
  36084=>"11111111",
  36085=>"11111111",
  36086=>"00000001",
  36087=>"00000001",
  36088=>"00000001",
  36089=>"00000000",
  36090=>"00000000",
  36091=>"00000001",
  36092=>"00000001",
  36093=>"11111110",
  36094=>"11111110",
  36095=>"11111100",
  36096=>"00000011",
  36097=>"11111111",
  36098=>"11111110",
  36099=>"00000100",
  36100=>"11111101",
  36101=>"00000101",
  36102=>"00000001",
  36103=>"11111111",
  36104=>"11111110",
  36105=>"00000011",
  36106=>"00000011",
  36107=>"00000001",
  36108=>"00000001",
  36109=>"11111111",
  36110=>"11111101",
  36111=>"11111100",
  36112=>"11111111",
  36113=>"11111111",
  36114=>"11111110",
  36115=>"11111101",
  36116=>"00000010",
  36117=>"11111110",
  36118=>"00000000",
  36119=>"00000010",
  36120=>"00000001",
  36121=>"11111101",
  36122=>"00000000",
  36123=>"11111110",
  36124=>"00000001",
  36125=>"00000010",
  36126=>"11111111",
  36127=>"11111111",
  36128=>"11111110",
  36129=>"00000000",
  36130=>"00000000",
  36131=>"11111110",
  36132=>"11111110",
  36133=>"11111100",
  36134=>"00000010",
  36135=>"11111111",
  36136=>"00000100",
  36137=>"11111111",
  36138=>"11111111",
  36139=>"00000011",
  36140=>"00000101",
  36141=>"00000000",
  36142=>"00000001",
  36143=>"00000100",
  36144=>"00000001",
  36145=>"11111110",
  36146=>"00000011",
  36147=>"00000001",
  36148=>"00000000",
  36149=>"11111110",
  36150=>"00000000",
  36151=>"00000011",
  36152=>"00000011",
  36153=>"00000001",
  36154=>"11111110",
  36155=>"11111110",
  36156=>"00000000",
  36157=>"11111110",
  36158=>"00000000",
  36159=>"00000010",
  36160=>"00000011",
  36161=>"00000010",
  36162=>"11111110",
  36163=>"11111110",
  36164=>"11111110",
  36165=>"00000010",
  36166=>"00000000",
  36167=>"00000001",
  36168=>"11111110",
  36169=>"11111101",
  36170=>"11111111",
  36171=>"11111101",
  36172=>"11111110",
  36173=>"11111111",
  36174=>"00000001",
  36175=>"11111101",
  36176=>"11111111",
  36177=>"00000000",
  36178=>"00000101",
  36179=>"00000001",
  36180=>"00000010",
  36181=>"11111111",
  36182=>"00000000",
  36183=>"11111111",
  36184=>"11111101",
  36185=>"00000000",
  36186=>"00000000",
  36187=>"00000010",
  36188=>"11111110",
  36189=>"11111110",
  36190=>"00000001",
  36191=>"11111110",
  36192=>"11111101",
  36193=>"00000010",
  36194=>"11111111",
  36195=>"11111100",
  36196=>"00000011",
  36197=>"11111101",
  36198=>"00000010",
  36199=>"11111101",
  36200=>"11111100",
  36201=>"00000000",
  36202=>"11111110",
  36203=>"11111111",
  36204=>"00000100",
  36205=>"00000101",
  36206=>"00000000",
  36207=>"00000000",
  36208=>"00000001",
  36209=>"00000000",
  36210=>"00000101",
  36211=>"11111110",
  36212=>"00000001",
  36213=>"11111111",
  36214=>"00000001",
  36215=>"11111110",
  36216=>"11111110",
  36217=>"11111100",
  36218=>"11111101",
  36219=>"00000000",
  36220=>"11111110",
  36221=>"00000001",
  36222=>"00000001",
  36223=>"11111111",
  36224=>"00000001",
  36225=>"11111100",
  36226=>"11111111",
  36227=>"00000000",
  36228=>"11111101",
  36229=>"11111110",
  36230=>"00000010",
  36231=>"11111101",
  36232=>"00000001",
  36233=>"00000001",
  36234=>"11111111",
  36235=>"00000010",
  36236=>"00000010",
  36237=>"00000011",
  36238=>"11111100",
  36239=>"11111110",
  36240=>"00000000",
  36241=>"11111101",
  36242=>"11111111",
  36243=>"11111111",
  36244=>"00000000",
  36245=>"11111101",
  36246=>"00000000",
  36247=>"11111101",
  36248=>"11111101",
  36249=>"00000010",
  36250=>"11111111",
  36251=>"00000001",
  36252=>"11111110",
  36253=>"11111110",
  36254=>"00000000",
  36255=>"11111110",
  36256=>"11111110",
  36257=>"00000100",
  36258=>"00000001",
  36259=>"11111110",
  36260=>"11111110",
  36261=>"11111110",
  36262=>"11111111",
  36263=>"11111101",
  36264=>"11111100",
  36265=>"00000001",
  36266=>"00000001",
  36267=>"00000011",
  36268=>"00000101",
  36269=>"00000110",
  36270=>"11111101",
  36271=>"11111110",
  36272=>"00000001",
  36273=>"00000011",
  36274=>"00000010",
  36275=>"00000000",
  36276=>"00000001",
  36277=>"11111110",
  36278=>"11111111",
  36279=>"11111101",
  36280=>"00000010",
  36281=>"11111101",
  36282=>"00000001",
  36283=>"11111110",
  36284=>"00000000",
  36285=>"11111110",
  36286=>"11111100",
  36287=>"00000010",
  36288=>"11111101",
  36289=>"00000000",
  36290=>"11111101",
  36291=>"11111110",
  36292=>"00000100",
  36293=>"00000000",
  36294=>"11111111",
  36295=>"00000011",
  36296=>"11111110",
  36297=>"11111110",
  36298=>"00000111",
  36299=>"11111101",
  36300=>"11111101",
  36301=>"11111101",
  36302=>"11111110",
  36303=>"00000100",
  36304=>"00000011",
  36305=>"11111100",
  36306=>"00000000",
  36307=>"11111111",
  36308=>"11111110",
  36309=>"00000101",
  36310=>"00000001",
  36311=>"00000011",
  36312=>"11111110",
  36313=>"11111110",
  36314=>"11111110",
  36315=>"00000000",
  36316=>"11111110",
  36317=>"11111101",
  36318=>"00000000",
  36319=>"11111111",
  36320=>"00000001",
  36321=>"11111111",
  36322=>"00000001",
  36323=>"00000001",
  36324=>"11111110",
  36325=>"11111111",
  36326=>"00000010",
  36327=>"00000000",
  36328=>"11111111",
  36329=>"00000000",
  36330=>"00000011",
  36331=>"11111111",
  36332=>"00000000",
  36333=>"00000110",
  36334=>"00000001",
  36335=>"00000000",
  36336=>"11111101",
  36337=>"00000011",
  36338=>"11111110",
  36339=>"11111110",
  36340=>"00000010",
  36341=>"00000011",
  36342=>"11111110",
  36343=>"11111101",
  36344=>"11111101",
  36345=>"11111110",
  36346=>"00000001",
  36347=>"11111110",
  36348=>"11111111",
  36349=>"11111111",
  36350=>"00000110",
  36351=>"11111110",
  36352=>"00000010",
  36353=>"00000000",
  36354=>"00000001",
  36355=>"00000010",
  36356=>"00000101",
  36357=>"00000000",
  36358=>"11111110",
  36359=>"00000000",
  36360=>"11111110",
  36361=>"00000001",
  36362=>"11111111",
  36363=>"00000011",
  36364=>"00000101",
  36365=>"00000001",
  36366=>"11111111",
  36367=>"00000001",
  36368=>"00000010",
  36369=>"11111111",
  36370=>"11111101",
  36371=>"11111111",
  36372=>"11111100",
  36373=>"11111111",
  36374=>"00000001",
  36375=>"11111101",
  36376=>"11111111",
  36377=>"11111111",
  36378=>"00000000",
  36379=>"11111101",
  36380=>"00000010",
  36381=>"11111110",
  36382=>"11111111",
  36383=>"11111111",
  36384=>"11111011",
  36385=>"11111110",
  36386=>"11111111",
  36387=>"00000010",
  36388=>"00000000",
  36389=>"00000011",
  36390=>"00000000",
  36391=>"00000010",
  36392=>"00000000",
  36393=>"00000001",
  36394=>"00000000",
  36395=>"11111110",
  36396=>"11111101",
  36397=>"00000010",
  36398=>"00000001",
  36399=>"00000001",
  36400=>"11111101",
  36401=>"00000100",
  36402=>"00000000",
  36403=>"00000000",
  36404=>"11111110",
  36405=>"11111110",
  36406=>"11111111",
  36407=>"00000111",
  36408=>"00000101",
  36409=>"00000010",
  36410=>"00000010",
  36411=>"11111111",
  36412=>"11111110",
  36413=>"11111110",
  36414=>"00000010",
  36415=>"11111110",
  36416=>"11111110",
  36417=>"11111101",
  36418=>"11111110",
  36419=>"00000010",
  36420=>"00000001",
  36421=>"00000011",
  36422=>"00000011",
  36423=>"11111101",
  36424=>"11111111",
  36425=>"11111111",
  36426=>"11111110",
  36427=>"00000010",
  36428=>"11111110",
  36429=>"11111110",
  36430=>"11111111",
  36431=>"11111111",
  36432=>"11111111",
  36433=>"00000001",
  36434=>"00000011",
  36435=>"00000001",
  36436=>"11111110",
  36437=>"11111110",
  36438=>"00000000",
  36439=>"00000011",
  36440=>"11111101",
  36441=>"11111111",
  36442=>"11111111",
  36443=>"00000001",
  36444=>"11111111",
  36445=>"11111111",
  36446=>"00000010",
  36447=>"00000001",
  36448=>"11111110",
  36449=>"11111110",
  36450=>"00000001",
  36451=>"11111111",
  36452=>"00000110",
  36453=>"00000000",
  36454=>"00000000",
  36455=>"11111111",
  36456=>"00000010",
  36457=>"00000010",
  36458=>"00000011",
  36459=>"11111111",
  36460=>"11111101",
  36461=>"11111111",
  36462=>"00000010",
  36463=>"11111110",
  36464=>"00000010",
  36465=>"00000001",
  36466=>"00000011",
  36467=>"00000001",
  36468=>"00000010",
  36469=>"00000000",
  36470=>"11111111",
  36471=>"11111100",
  36472=>"00000010",
  36473=>"00000011",
  36474=>"00000010",
  36475=>"00000000",
  36476=>"11111111",
  36477=>"00000001",
  36478=>"11111100",
  36479=>"00000010",
  36480=>"00000010",
  36481=>"00000011",
  36482=>"11111101",
  36483=>"00000000",
  36484=>"11111110",
  36485=>"11111111",
  36486=>"11111101",
  36487=>"11111110",
  36488=>"11111101",
  36489=>"11111101",
  36490=>"11111111",
  36491=>"11111110",
  36492=>"00000001",
  36493=>"11111110",
  36494=>"00000001",
  36495=>"00000011",
  36496=>"00000010",
  36497=>"00000001",
  36498=>"00000010",
  36499=>"00000010",
  36500=>"11111110",
  36501=>"11111101",
  36502=>"00000010",
  36503=>"11111100",
  36504=>"11111101",
  36505=>"00000001",
  36506=>"11111110",
  36507=>"11111111",
  36508=>"11111110",
  36509=>"11111110",
  36510=>"11111111",
  36511=>"00000011",
  36512=>"11111101",
  36513=>"11111110",
  36514=>"00000001",
  36515=>"11111101",
  36516=>"00000001",
  36517=>"00000001",
  36518=>"11111110",
  36519=>"11111100",
  36520=>"00000011",
  36521=>"00000111",
  36522=>"11111111",
  36523=>"11111111",
  36524=>"11111101",
  36525=>"11111111",
  36526=>"11111110",
  36527=>"00000011",
  36528=>"11111110",
  36529=>"00000100",
  36530=>"00000000",
  36531=>"00000010",
  36532=>"11111110",
  36533=>"00000001",
  36534=>"00000010",
  36535=>"00000010",
  36536=>"11111110",
  36537=>"00000010",
  36538=>"00000010",
  36539=>"00000011",
  36540=>"11111101",
  36541=>"11111110",
  36542=>"11111110",
  36543=>"11111101",
  36544=>"00000010",
  36545=>"00000100",
  36546=>"00000000",
  36547=>"11111111",
  36548=>"00000010",
  36549=>"00000000",
  36550=>"11111110",
  36551=>"00000000",
  36552=>"00000000",
  36553=>"00000110",
  36554=>"00000100",
  36555=>"00000001",
  36556=>"11111110",
  36557=>"11111110",
  36558=>"00000001",
  36559=>"00000000",
  36560=>"11111111",
  36561=>"00000000",
  36562=>"11111101",
  36563=>"11111111",
  36564=>"11111110",
  36565=>"00000000",
  36566=>"00000101",
  36567=>"00000000",
  36568=>"11111111",
  36569=>"00000001",
  36570=>"00000010",
  36571=>"11111111",
  36572=>"11111100",
  36573=>"00000011",
  36574=>"11111111",
  36575=>"00000001",
  36576=>"00000001",
  36577=>"00000111",
  36578=>"00000000",
  36579=>"00000000",
  36580=>"00000000",
  36581=>"11111100",
  36582=>"11111101",
  36583=>"11111110",
  36584=>"11111101",
  36585=>"11111111",
  36586=>"11111110",
  36587=>"00000000",
  36588=>"00000001",
  36589=>"00000110",
  36590=>"11111110",
  36591=>"00000010",
  36592=>"11111110",
  36593=>"11111110",
  36594=>"00000001",
  36595=>"00000000",
  36596=>"00000100",
  36597=>"11111111",
  36598=>"00000001",
  36599=>"11111111",
  36600=>"11111110",
  36601=>"00000000",
  36602=>"00000000",
  36603=>"11111110",
  36604=>"11111111",
  36605=>"11111100",
  36606=>"00000010",
  36607=>"11111110",
  36608=>"00000010",
  36609=>"11111110",
  36610=>"00000101",
  36611=>"00000000",
  36612=>"11111111",
  36613=>"11111111",
  36614=>"11111101",
  36615=>"11111111",
  36616=>"11111111",
  36617=>"11111110",
  36618=>"00000001",
  36619=>"11111101",
  36620=>"11111101",
  36621=>"00000101",
  36622=>"00000100",
  36623=>"11111111",
  36624=>"11111101",
  36625=>"11111111",
  36626=>"00000010",
  36627=>"00000010",
  36628=>"00000010",
  36629=>"11111111",
  36630=>"11111110",
  36631=>"11111101",
  36632=>"00000110",
  36633=>"00000000",
  36634=>"11111111",
  36635=>"11111101",
  36636=>"00000001",
  36637=>"11111101",
  36638=>"00000000",
  36639=>"00000101",
  36640=>"00000001",
  36641=>"00000011",
  36642=>"11111111",
  36643=>"11111100",
  36644=>"00000101",
  36645=>"00000000",
  36646=>"00000001",
  36647=>"11111110",
  36648=>"11111111",
  36649=>"11111110",
  36650=>"00000000",
  36651=>"00000000",
  36652=>"11111111",
  36653=>"11111111",
  36654=>"11111101",
  36655=>"00000000",
  36656=>"00000001",
  36657=>"00000101",
  36658=>"00000000",
  36659=>"00000010",
  36660=>"00000000",
  36661=>"00000010",
  36662=>"00000011",
  36663=>"11111111",
  36664=>"00000000",
  36665=>"11111111",
  36666=>"00000010",
  36667=>"11111101",
  36668=>"11111111",
  36669=>"11111111",
  36670=>"11111101",
  36671=>"11111101",
  36672=>"11111101",
  36673=>"11111111",
  36674=>"11111110",
  36675=>"11111101",
  36676=>"00000100",
  36677=>"00000000",
  36678=>"11111111",
  36679=>"11111110",
  36680=>"11111101",
  36681=>"00000011",
  36682=>"11111101",
  36683=>"00000000",
  36684=>"11111111",
  36685=>"11111101",
  36686=>"11111101",
  36687=>"11111110",
  36688=>"11111101",
  36689=>"00000001",
  36690=>"00000101",
  36691=>"11111111",
  36692=>"11111110",
  36693=>"00000011",
  36694=>"11111101",
  36695=>"00000011",
  36696=>"11111110",
  36697=>"00000011",
  36698=>"11111101",
  36699=>"00000001",
  36700=>"11111110",
  36701=>"11111101",
  36702=>"00000110",
  36703=>"00000000",
  36704=>"00000001",
  36705=>"11111100",
  36706=>"00000000",
  36707=>"11111101",
  36708=>"00000001",
  36709=>"11111100",
  36710=>"00000001",
  36711=>"00000011",
  36712=>"00000011",
  36713=>"00000011",
  36714=>"11111110",
  36715=>"11111111",
  36716=>"00000001",
  36717=>"11111111",
  36718=>"00000000",
  36719=>"00000010",
  36720=>"00000001",
  36721=>"11111111",
  36722=>"00000000",
  36723=>"11111110",
  36724=>"11111111",
  36725=>"00000010",
  36726=>"11111101",
  36727=>"00000001",
  36728=>"11111110",
  36729=>"11111110",
  36730=>"11111111",
  36731=>"00000001",
  36732=>"11111110",
  36733=>"11111110",
  36734=>"11111110",
  36735=>"00000001",
  36736=>"11111111",
  36737=>"00000001",
  36738=>"11111110",
  36739=>"00000011",
  36740=>"00000001",
  36741=>"00000001",
  36742=>"00000010",
  36743=>"00000010",
  36744=>"11111111",
  36745=>"00000101",
  36746=>"11111110",
  36747=>"11111110",
  36748=>"11111110",
  36749=>"00000001",
  36750=>"11111101",
  36751=>"00000010",
  36752=>"11111111",
  36753=>"11111110",
  36754=>"11111101",
  36755=>"00000011",
  36756=>"00000101",
  36757=>"11111101",
  36758=>"00000000",
  36759=>"11111110",
  36760=>"11111101",
  36761=>"00000001",
  36762=>"00000001",
  36763=>"00000000",
  36764=>"11111011",
  36765=>"11111110",
  36766=>"11111111",
  36767=>"11111101",
  36768=>"00000001",
  36769=>"00000000",
  36770=>"11111101",
  36771=>"00000001",
  36772=>"11111110",
  36773=>"00000011",
  36774=>"00000000",
  36775=>"00000100",
  36776=>"00000001",
  36777=>"00000011",
  36778=>"00000100",
  36779=>"00000001",
  36780=>"00000000",
  36781=>"00000011",
  36782=>"11111111",
  36783=>"11111101",
  36784=>"00000001",
  36785=>"11111111",
  36786=>"00000001",
  36787=>"00000100",
  36788=>"00000000",
  36789=>"11111101",
  36790=>"00000010",
  36791=>"00000001",
  36792=>"00000100",
  36793=>"00000010",
  36794=>"11111111",
  36795=>"00000110",
  36796=>"00000110",
  36797=>"00000001",
  36798=>"11111110",
  36799=>"00000011",
  36800=>"11111110",
  36801=>"00000000",
  36802=>"00000001",
  36803=>"11111111",
  36804=>"11111101",
  36805=>"00000000",
  36806=>"11111100",
  36807=>"00000001",
  36808=>"11111111",
  36809=>"00000011",
  36810=>"11111110",
  36811=>"00000010",
  36812=>"00000110",
  36813=>"00000011",
  36814=>"00000011",
  36815=>"11111111",
  36816=>"00000000",
  36817=>"00000001",
  36818=>"00000110",
  36819=>"00000001",
  36820=>"00000011",
  36821=>"00000000",
  36822=>"00000011",
  36823=>"00000010",
  36824=>"00000001",
  36825=>"11111110",
  36826=>"00000000",
  36827=>"11111111",
  36828=>"00000001",
  36829=>"00000000",
  36830=>"11111110",
  36831=>"11111100",
  36832=>"11111110",
  36833=>"00000110",
  36834=>"11111111",
  36835=>"11111110",
  36836=>"11111111",
  36837=>"00000001",
  36838=>"11111101",
  36839=>"00000000",
  36840=>"11111111",
  36841=>"11111111",
  36842=>"11111111",
  36843=>"11111111",
  36844=>"11111110",
  36845=>"11111111",
  36846=>"00000000",
  36847=>"11111111",
  36848=>"11111110",
  36849=>"00000000",
  36850=>"00000000",
  36851=>"11111101",
  36852=>"00000001",
  36853=>"11111101",
  36854=>"00000010",
  36855=>"00000001",
  36856=>"11111101",
  36857=>"00000000",
  36858=>"11111101",
  36859=>"00000010",
  36860=>"11111111",
  36861=>"11111111",
  36862=>"00000010",
  36863=>"00000001",
  36864=>"11111111",
  36865=>"11111110",
  36866=>"11111101",
  36867=>"00000001",
  36868=>"00000011",
  36869=>"11111100",
  36870=>"11111111",
  36871=>"11111100",
  36872=>"00000000",
  36873=>"00000110",
  36874=>"00000000",
  36875=>"00000010",
  36876=>"00000000",
  36877=>"11111100",
  36878=>"11111100",
  36879=>"00000001",
  36880=>"00000000",
  36881=>"11111101",
  36882=>"00000101",
  36883=>"11111110",
  36884=>"11111110",
  36885=>"00000010",
  36886=>"00000100",
  36887=>"00000001",
  36888=>"11111100",
  36889=>"11111100",
  36890=>"11111111",
  36891=>"00000000",
  36892=>"00000000",
  36893=>"11111110",
  36894=>"11111111",
  36895=>"00000100",
  36896=>"00000011",
  36897=>"11111111",
  36898=>"00000001",
  36899=>"00000000",
  36900=>"00000001",
  36901=>"11111100",
  36902=>"00000010",
  36903=>"00000011",
  36904=>"00000011",
  36905=>"11111100",
  36906=>"00000010",
  36907=>"11111110",
  36908=>"11111111",
  36909=>"00000000",
  36910=>"11111110",
  36911=>"00000100",
  36912=>"11111101",
  36913=>"00000011",
  36914=>"11111011",
  36915=>"11111111",
  36916=>"00000000",
  36917=>"00000110",
  36918=>"00000010",
  36919=>"00000001",
  36920=>"00000100",
  36921=>"11111111",
  36922=>"00000010",
  36923=>"11111111",
  36924=>"00000010",
  36925=>"00000001",
  36926=>"11111110",
  36927=>"00000011",
  36928=>"11111011",
  36929=>"00000010",
  36930=>"11111111",
  36931=>"00000001",
  36932=>"00000101",
  36933=>"11111101",
  36934=>"11111110",
  36935=>"00000110",
  36936=>"11111111",
  36937=>"11111110",
  36938=>"11111111",
  36939=>"00000001",
  36940=>"00000001",
  36941=>"11111101",
  36942=>"00000000",
  36943=>"00000001",
  36944=>"11111101",
  36945=>"00000000",
  36946=>"11111110",
  36947=>"00000001",
  36948=>"00000000",
  36949=>"11111100",
  36950=>"11111110",
  36951=>"11111110",
  36952=>"11111101",
  36953=>"00000100",
  36954=>"00000000",
  36955=>"11111101",
  36956=>"00000001",
  36957=>"00000100",
  36958=>"00000010",
  36959=>"11111111",
  36960=>"00000001",
  36961=>"00000100",
  36962=>"11111110",
  36963=>"00000011",
  36964=>"11111110",
  36965=>"00000001",
  36966=>"00000000",
  36967=>"11111101",
  36968=>"00000000",
  36969=>"11111101",
  36970=>"00000000",
  36971=>"11111110",
  36972=>"11111111",
  36973=>"00000000",
  36974=>"11111110",
  36975=>"00000100",
  36976=>"00000010",
  36977=>"00000010",
  36978=>"00000000",
  36979=>"11111101",
  36980=>"00000001",
  36981=>"11111100",
  36982=>"11111110",
  36983=>"00000101",
  36984=>"00000001",
  36985=>"11111100",
  36986=>"11111110",
  36987=>"11111111",
  36988=>"11111101",
  36989=>"00000011",
  36990=>"11111101",
  36991=>"00000011",
  36992=>"00000001",
  36993=>"11111100",
  36994=>"00000011",
  36995=>"00000010",
  36996=>"00000100",
  36997=>"11111111",
  36998=>"11111111",
  36999=>"00000010",
  37000=>"11111111",
  37001=>"00000011",
  37002=>"11111101",
  37003=>"11111101",
  37004=>"00000000",
  37005=>"11111111",
  37006=>"00000011",
  37007=>"11111011",
  37008=>"00000101",
  37009=>"11111111",
  37010=>"11111110",
  37011=>"00000000",
  37012=>"00000000",
  37013=>"00000000",
  37014=>"00000010",
  37015=>"11111111",
  37016=>"00000001",
  37017=>"00000000",
  37018=>"00000001",
  37019=>"00000010",
  37020=>"11111111",
  37021=>"00000010",
  37022=>"00000001",
  37023=>"11111101",
  37024=>"11111101",
  37025=>"00000001",
  37026=>"11111101",
  37027=>"00000101",
  37028=>"11111110",
  37029=>"11111101",
  37030=>"00000001",
  37031=>"00000000",
  37032=>"11111101",
  37033=>"00000011",
  37034=>"00000010",
  37035=>"11111111",
  37036=>"11111100",
  37037=>"00000001",
  37038=>"00000000",
  37039=>"11111101",
  37040=>"11111110",
  37041=>"00000001",
  37042=>"00000000",
  37043=>"00000000",
  37044=>"11111111",
  37045=>"11111100",
  37046=>"00000010",
  37047=>"11111100",
  37048=>"00000001",
  37049=>"00000000",
  37050=>"00000010",
  37051=>"11111101",
  37052=>"11111110",
  37053=>"00000000",
  37054=>"11111111",
  37055=>"00000000",
  37056=>"00000010",
  37057=>"00000001",
  37058=>"11111111",
  37059=>"00000101",
  37060=>"00000101",
  37061=>"00000101",
  37062=>"00000001",
  37063=>"00000010",
  37064=>"00000000",
  37065=>"11111111",
  37066=>"11111110",
  37067=>"00000000",
  37068=>"00000101",
  37069=>"00000011",
  37070=>"00000000",
  37071=>"11111100",
  37072=>"00000001",
  37073=>"11111101",
  37074=>"00000001",
  37075=>"00000010",
  37076=>"00000000",
  37077=>"11111101",
  37078=>"00000011",
  37079=>"11111101",
  37080=>"00000010",
  37081=>"00000000",
  37082=>"00000000",
  37083=>"00000010",
  37084=>"11111110",
  37085=>"11111101",
  37086=>"00000011",
  37087=>"00000010",
  37088=>"00000001",
  37089=>"11111101",
  37090=>"00000001",
  37091=>"11111111",
  37092=>"11111101",
  37093=>"11111110",
  37094=>"00000001",
  37095=>"00000001",
  37096=>"00000010",
  37097=>"00000010",
  37098=>"11111111",
  37099=>"00000001",
  37100=>"00000010",
  37101=>"00000100",
  37102=>"00000010",
  37103=>"11111110",
  37104=>"11111101",
  37105=>"11111110",
  37106=>"11111101",
  37107=>"00000100",
  37108=>"00000000",
  37109=>"11111010",
  37110=>"11111101",
  37111=>"00000011",
  37112=>"00000001",
  37113=>"00000000",
  37114=>"11111110",
  37115=>"00000010",
  37116=>"00000011",
  37117=>"00000100",
  37118=>"00000001",
  37119=>"00000001",
  37120=>"11111110",
  37121=>"11111111",
  37122=>"11111100",
  37123=>"00000000",
  37124=>"00000010",
  37125=>"00000001",
  37126=>"11111100",
  37127=>"00000100",
  37128=>"00000000",
  37129=>"11111110",
  37130=>"00000001",
  37131=>"11111111",
  37132=>"11111111",
  37133=>"11111100",
  37134=>"00000011",
  37135=>"11111110",
  37136=>"00000000",
  37137=>"00000010",
  37138=>"00000000",
  37139=>"11111110",
  37140=>"00000010",
  37141=>"11111111",
  37142=>"00000010",
  37143=>"00000001",
  37144=>"11111101",
  37145=>"11111101",
  37146=>"11111111",
  37147=>"00000010",
  37148=>"00000101",
  37149=>"11111101",
  37150=>"00000000",
  37151=>"11111011",
  37152=>"00000001",
  37153=>"00000001",
  37154=>"00000000",
  37155=>"00000010",
  37156=>"11111101",
  37157=>"00000010",
  37158=>"11111111",
  37159=>"00000010",
  37160=>"00000100",
  37161=>"00000001",
  37162=>"11111101",
  37163=>"00000110",
  37164=>"00000010",
  37165=>"00000001",
  37166=>"00000000",
  37167=>"11111110",
  37168=>"00000000",
  37169=>"00000010",
  37170=>"00000011",
  37171=>"11111111",
  37172=>"11111111",
  37173=>"00000001",
  37174=>"11111110",
  37175=>"11111111",
  37176=>"00000101",
  37177=>"00000000",
  37178=>"00000000",
  37179=>"00000001",
  37180=>"11111111",
  37181=>"00000001",
  37182=>"00000011",
  37183=>"11111111",
  37184=>"11111111",
  37185=>"11111110",
  37186=>"00000011",
  37187=>"00000001",
  37188=>"00000001",
  37189=>"11111111",
  37190=>"00000011",
  37191=>"11111111",
  37192=>"11111101",
  37193=>"00000010",
  37194=>"11111111",
  37195=>"11111110",
  37196=>"11111101",
  37197=>"00000111",
  37198=>"00000000",
  37199=>"11111100",
  37200=>"00000001",
  37201=>"00000000",
  37202=>"00000100",
  37203=>"11111101",
  37204=>"11111111",
  37205=>"00000011",
  37206=>"00000000",
  37207=>"00000011",
  37208=>"11111110",
  37209=>"00000010",
  37210=>"00000001",
  37211=>"00000000",
  37212=>"00000001",
  37213=>"00000001",
  37214=>"00000011",
  37215=>"11111100",
  37216=>"00000011",
  37217=>"00000010",
  37218=>"00000001",
  37219=>"00000000",
  37220=>"11111110",
  37221=>"11111101",
  37222=>"11111101",
  37223=>"11111110",
  37224=>"00000011",
  37225=>"11111111",
  37226=>"11111111",
  37227=>"11111101",
  37228=>"00000001",
  37229=>"11111110",
  37230=>"11111101",
  37231=>"11111110",
  37232=>"00000000",
  37233=>"00000011",
  37234=>"00000001",
  37235=>"00000010",
  37236=>"11111110",
  37237=>"00000010",
  37238=>"00000001",
  37239=>"00000010",
  37240=>"11111111",
  37241=>"00000000",
  37242=>"00000000",
  37243=>"11111101",
  37244=>"11111101",
  37245=>"11111111",
  37246=>"11111101",
  37247=>"00000011",
  37248=>"11111101",
  37249=>"00000000",
  37250=>"11111110",
  37251=>"11111111",
  37252=>"00000011",
  37253=>"00000001",
  37254=>"00000001",
  37255=>"11111111",
  37256=>"00000100",
  37257=>"11111101",
  37258=>"00000010",
  37259=>"00000000",
  37260=>"11111101",
  37261=>"11111111",
  37262=>"00000100",
  37263=>"00000011",
  37264=>"11111101",
  37265=>"00000101",
  37266=>"00000010",
  37267=>"00000001",
  37268=>"00000000",
  37269=>"00000001",
  37270=>"11111111",
  37271=>"11111110",
  37272=>"00000001",
  37273=>"00000100",
  37274=>"11111101",
  37275=>"00000101",
  37276=>"11111111",
  37277=>"11111111",
  37278=>"00000001",
  37279=>"11111110",
  37280=>"00000101",
  37281=>"11111110",
  37282=>"00000000",
  37283=>"00000001",
  37284=>"00000000",
  37285=>"11111111",
  37286=>"11111110",
  37287=>"11111110",
  37288=>"00000000",
  37289=>"11111101",
  37290=>"00000001",
  37291=>"00000010",
  37292=>"11111111",
  37293=>"11111110",
  37294=>"00000011",
  37295=>"11111101",
  37296=>"11111101",
  37297=>"00000001",
  37298=>"11111100",
  37299=>"00000001",
  37300=>"00000000",
  37301=>"00000001",
  37302=>"11111101",
  37303=>"11111111",
  37304=>"11111111",
  37305=>"11111101",
  37306=>"00000010",
  37307=>"00000101",
  37308=>"00000000",
  37309=>"11111111",
  37310=>"11111111",
  37311=>"11111111",
  37312=>"11111111",
  37313=>"11111101",
  37314=>"11111100",
  37315=>"00000111",
  37316=>"00000001",
  37317=>"00000011",
  37318=>"11111110",
  37319=>"11111110",
  37320=>"00000010",
  37321=>"11111110",
  37322=>"11111110",
  37323=>"11111110",
  37324=>"11111110",
  37325=>"00000011",
  37326=>"00000000",
  37327=>"00000010",
  37328=>"11111111",
  37329=>"00000001",
  37330=>"00000011",
  37331=>"11111011",
  37332=>"11111101",
  37333=>"00000001",
  37334=>"00000101",
  37335=>"00000000",
  37336=>"00000011",
  37337=>"11111111",
  37338=>"11111111",
  37339=>"00000000",
  37340=>"00000011",
  37341=>"00000000",
  37342=>"00000010",
  37343=>"11111111",
  37344=>"00000011",
  37345=>"11111011",
  37346=>"11111101",
  37347=>"11111111",
  37348=>"00000010",
  37349=>"00000010",
  37350=>"00000010",
  37351=>"00000001",
  37352=>"00000001",
  37353=>"00000001",
  37354=>"11111110",
  37355=>"11111100",
  37356=>"00000010",
  37357=>"00000011",
  37358=>"00000100",
  37359=>"11111100",
  37360=>"00000000",
  37361=>"11111111",
  37362=>"11111111",
  37363=>"11111111",
  37364=>"11111101",
  37365=>"11111100",
  37366=>"11111101",
  37367=>"00000110",
  37368=>"00000000",
  37369=>"00000000",
  37370=>"11111101",
  37371=>"00000010",
  37372=>"11111101",
  37373=>"11111100",
  37374=>"00000101",
  37375=>"00000010",
  37376=>"11111110",
  37377=>"11111101",
  37378=>"11111110",
  37379=>"11111101",
  37380=>"00000011",
  37381=>"00000101",
  37382=>"11111011",
  37383=>"11111111",
  37384=>"00000000",
  37385=>"11111100",
  37386=>"00000000",
  37387=>"00000000",
  37388=>"11111110",
  37389=>"11111111",
  37390=>"00000001",
  37391=>"11111111",
  37392=>"00000001",
  37393=>"00000011",
  37394=>"11111110",
  37395=>"00000011",
  37396=>"11111011",
  37397=>"11111111",
  37398=>"00000001",
  37399=>"00000010",
  37400=>"00000101",
  37401=>"00000100",
  37402=>"00000001",
  37403=>"11111101",
  37404=>"11111101",
  37405=>"00000011",
  37406=>"11111101",
  37407=>"11111101",
  37408=>"00000001",
  37409=>"11111111",
  37410=>"11111111",
  37411=>"00000000",
  37412=>"11111110",
  37413=>"11111111",
  37414=>"00000001",
  37415=>"00000101",
  37416=>"11111111",
  37417=>"00000000",
  37418=>"11111111",
  37419=>"00000010",
  37420=>"00000000",
  37421=>"00000010",
  37422=>"11111110",
  37423=>"11111111",
  37424=>"00000001",
  37425=>"11111110",
  37426=>"11111101",
  37427=>"00000000",
  37428=>"00000001",
  37429=>"00000001",
  37430=>"00000001",
  37431=>"00000010",
  37432=>"00000010",
  37433=>"00000100",
  37434=>"00000001",
  37435=>"00000001",
  37436=>"11111101",
  37437=>"00000010",
  37438=>"00000101",
  37439=>"00000010",
  37440=>"11111101",
  37441=>"11111100",
  37442=>"11111110",
  37443=>"11111101",
  37444=>"00000000",
  37445=>"11111101",
  37446=>"11111100",
  37447=>"11111101",
  37448=>"11111111",
  37449=>"00000001",
  37450=>"00000010",
  37451=>"00000010",
  37452=>"11111110",
  37453=>"00000010",
  37454=>"00000000",
  37455=>"00000010",
  37456=>"11111110",
  37457=>"11111100",
  37458=>"00000000",
  37459=>"00000010",
  37460=>"00000100",
  37461=>"00000010",
  37462=>"00000000",
  37463=>"00000000",
  37464=>"00000100",
  37465=>"11111101",
  37466=>"11111111",
  37467=>"11111101",
  37468=>"11111100",
  37469=>"11111110",
  37470=>"11111101",
  37471=>"11111110",
  37472=>"00000000",
  37473=>"11111111",
  37474=>"00000001",
  37475=>"11111101",
  37476=>"11111110",
  37477=>"00000010",
  37478=>"00000000",
  37479=>"00000001",
  37480=>"11111110",
  37481=>"11111110",
  37482=>"00000011",
  37483=>"00000000",
  37484=>"11111101",
  37485=>"00000000",
  37486=>"00000000",
  37487=>"00000001",
  37488=>"11111100",
  37489=>"11111110",
  37490=>"11111110",
  37491=>"11111100",
  37492=>"11111110",
  37493=>"00000010",
  37494=>"00000000",
  37495=>"00000001",
  37496=>"00000001",
  37497=>"00000100",
  37498=>"11111101",
  37499=>"00000101",
  37500=>"11111110",
  37501=>"11111110",
  37502=>"11111110",
  37503=>"00000001",
  37504=>"00000000",
  37505=>"00000101",
  37506=>"00000001",
  37507=>"00000011",
  37508=>"00000001",
  37509=>"11111100",
  37510=>"00000001",
  37511=>"11111101",
  37512=>"11111111",
  37513=>"00000000",
  37514=>"00000001",
  37515=>"00000001",
  37516=>"00000000",
  37517=>"11111111",
  37518=>"00000010",
  37519=>"00000001",
  37520=>"11111110",
  37521=>"11111100",
  37522=>"00000010",
  37523=>"11111111",
  37524=>"11111111",
  37525=>"11111101",
  37526=>"11111111",
  37527=>"11111110",
  37528=>"11111110",
  37529=>"00000000",
  37530=>"11111110",
  37531=>"00000001",
  37532=>"00000000",
  37533=>"11111101",
  37534=>"11111101",
  37535=>"00000101",
  37536=>"11111110",
  37537=>"11111011",
  37538=>"00000011",
  37539=>"11111100",
  37540=>"11111110",
  37541=>"00000001",
  37542=>"11111101",
  37543=>"00000001",
  37544=>"11111101",
  37545=>"00000101",
  37546=>"11111101",
  37547=>"00000001",
  37548=>"11111110",
  37549=>"11111110",
  37550=>"11111111",
  37551=>"11111111",
  37552=>"11111110",
  37553=>"11111100",
  37554=>"00000011",
  37555=>"00000011",
  37556=>"11111111",
  37557=>"11111101",
  37558=>"11111110",
  37559=>"00000100",
  37560=>"00000000",
  37561=>"11111111",
  37562=>"11111110",
  37563=>"00000100",
  37564=>"00000010",
  37565=>"11111111",
  37566=>"00000011",
  37567=>"11111111",
  37568=>"00000001",
  37569=>"00000101",
  37570=>"11111101",
  37571=>"00000011",
  37572=>"00000011",
  37573=>"11111101",
  37574=>"11111111",
  37575=>"11111100",
  37576=>"11111110",
  37577=>"00000011",
  37578=>"00000001",
  37579=>"11111111",
  37580=>"11111100",
  37581=>"11111101",
  37582=>"11111110",
  37583=>"11111110",
  37584=>"11111110",
  37585=>"11111101",
  37586=>"11111101",
  37587=>"11111111",
  37588=>"11111101",
  37589=>"11111111",
  37590=>"00000001",
  37591=>"00000010",
  37592=>"00000001",
  37593=>"00000001",
  37594=>"00000001",
  37595=>"00000001",
  37596=>"11111011",
  37597=>"00000010",
  37598=>"00000101",
  37599=>"00000001",
  37600=>"11111111",
  37601=>"00000110",
  37602=>"11111110",
  37603=>"11111111",
  37604=>"11111111",
  37605=>"00000100",
  37606=>"11111111",
  37607=>"00000000",
  37608=>"00000000",
  37609=>"11111101",
  37610=>"00000110",
  37611=>"00000011",
  37612=>"11111111",
  37613=>"11111100",
  37614=>"00000011",
  37615=>"00000100",
  37616=>"11111100",
  37617=>"00000011",
  37618=>"11111111",
  37619=>"00000000",
  37620=>"11111101",
  37621=>"11111011",
  37622=>"11111111",
  37623=>"00000010",
  37624=>"00000000",
  37625=>"00000011",
  37626=>"11111110",
  37627=>"00000100",
  37628=>"00000001",
  37629=>"00000001",
  37630=>"11111110",
  37631=>"11111111",
  37632=>"00000101",
  37633=>"00000100",
  37634=>"00000000",
  37635=>"00000010",
  37636=>"11111111",
  37637=>"00000100",
  37638=>"00000010",
  37639=>"11111100",
  37640=>"11111100",
  37641=>"00000100",
  37642=>"00000001",
  37643=>"11111111",
  37644=>"00000001",
  37645=>"00000011",
  37646=>"11111110",
  37647=>"00000010",
  37648=>"00000000",
  37649=>"00000001",
  37650=>"11111110",
  37651=>"00000001",
  37652=>"00000001",
  37653=>"00000001",
  37654=>"00000000",
  37655=>"00000001",
  37656=>"11111111",
  37657=>"00000100",
  37658=>"11111111",
  37659=>"11111101",
  37660=>"00000011",
  37661=>"00000100",
  37662=>"11111111",
  37663=>"00000110",
  37664=>"00000011",
  37665=>"11111111",
  37666=>"11111101",
  37667=>"00000000",
  37668=>"11111111",
  37669=>"00000101",
  37670=>"00000011",
  37671=>"11111110",
  37672=>"00000000",
  37673=>"00000000",
  37674=>"00000001",
  37675=>"11111111",
  37676=>"11111111",
  37677=>"11111100",
  37678=>"11111110",
  37679=>"00000010",
  37680=>"00000010",
  37681=>"00000011",
  37682=>"00000101",
  37683=>"00000000",
  37684=>"11111110",
  37685=>"11111110",
  37686=>"00000010",
  37687=>"00000000",
  37688=>"11111101",
  37689=>"00000001",
  37690=>"00000010",
  37691=>"11111110",
  37692=>"11111111",
  37693=>"11111111",
  37694=>"11111101",
  37695=>"11111100",
  37696=>"00000010",
  37697=>"11111110",
  37698=>"11111110",
  37699=>"00000001",
  37700=>"00000001",
  37701=>"11111111",
  37702=>"00000011",
  37703=>"11111100",
  37704=>"00000001",
  37705=>"00000001",
  37706=>"11111111",
  37707=>"00000010",
  37708=>"00000100",
  37709=>"00000001",
  37710=>"00000110",
  37711=>"00000000",
  37712=>"11111111",
  37713=>"00000000",
  37714=>"00000110",
  37715=>"00000001",
  37716=>"00000001",
  37717=>"00000100",
  37718=>"11111111",
  37719=>"11111101",
  37720=>"11111110",
  37721=>"11111101",
  37722=>"00000000",
  37723=>"00000001",
  37724=>"11111111",
  37725=>"00000001",
  37726=>"00000001",
  37727=>"00000110",
  37728=>"00000100",
  37729=>"11111101",
  37730=>"11111111",
  37731=>"11111101",
  37732=>"00000000",
  37733=>"00000000",
  37734=>"11111110",
  37735=>"00000110",
  37736=>"11111110",
  37737=>"00000011",
  37738=>"00000010",
  37739=>"11111100",
  37740=>"00000001",
  37741=>"00000010",
  37742=>"11111111",
  37743=>"00000100",
  37744=>"11111101",
  37745=>"00000011",
  37746=>"00000001",
  37747=>"00000101",
  37748=>"11111111",
  37749=>"00000110",
  37750=>"11111011",
  37751=>"00000001",
  37752=>"11111100",
  37753=>"11111110",
  37754=>"00000001",
  37755=>"00000000",
  37756=>"00000010",
  37757=>"00000001",
  37758=>"11111111",
  37759=>"00000100",
  37760=>"00000000",
  37761=>"11111101",
  37762=>"11111110",
  37763=>"00000100",
  37764=>"00000100",
  37765=>"00000000",
  37766=>"00000100",
  37767=>"11111101",
  37768=>"11111111",
  37769=>"00000101",
  37770=>"11111111",
  37771=>"00000011",
  37772=>"00000000",
  37773=>"00000001",
  37774=>"00000001",
  37775=>"00000000",
  37776=>"11111111",
  37777=>"00000000",
  37778=>"11111110",
  37779=>"00000001",
  37780=>"00000000",
  37781=>"11111111",
  37782=>"11111111",
  37783=>"11111111",
  37784=>"00000011",
  37785=>"00000100",
  37786=>"11111101",
  37787=>"00000000",
  37788=>"11111101",
  37789=>"00000001",
  37790=>"00000010",
  37791=>"00000000",
  37792=>"00000010",
  37793=>"00000100",
  37794=>"00000000",
  37795=>"00000001",
  37796=>"11111111",
  37797=>"00000010",
  37798=>"00000000",
  37799=>"00000011",
  37800=>"11111111",
  37801=>"00000010",
  37802=>"00000001",
  37803=>"00000001",
  37804=>"00000001",
  37805=>"00000010",
  37806=>"00000011",
  37807=>"00000011",
  37808=>"00000010",
  37809=>"11111110",
  37810=>"00000000",
  37811=>"11111110",
  37812=>"00000000",
  37813=>"11111100",
  37814=>"00000001",
  37815=>"00000001",
  37816=>"00000111",
  37817=>"00000100",
  37818=>"00000100",
  37819=>"11111100",
  37820=>"00000011",
  37821=>"00000001",
  37822=>"00000010",
  37823=>"00000000",
  37824=>"11111110",
  37825=>"00000011",
  37826=>"11111101",
  37827=>"00000010",
  37828=>"00000011",
  37829=>"11111100",
  37830=>"11111111",
  37831=>"11111110",
  37832=>"11111100",
  37833=>"11111111",
  37834=>"00000011",
  37835=>"00000010",
  37836=>"00000001",
  37837=>"00000011",
  37838=>"00000000",
  37839=>"11111110",
  37840=>"00000100",
  37841=>"11111111",
  37842=>"00000011",
  37843=>"00000001",
  37844=>"11111111",
  37845=>"00000011",
  37846=>"00000001",
  37847=>"11111111",
  37848=>"00000001",
  37849=>"00000101",
  37850=>"11111110",
  37851=>"00000000",
  37852=>"11111111",
  37853=>"11111101",
  37854=>"00000001",
  37855=>"00000010",
  37856=>"11111110",
  37857=>"00000011",
  37858=>"00000001",
  37859=>"11111111",
  37860=>"11111101",
  37861=>"11111110",
  37862=>"00000000",
  37863=>"11111101",
  37864=>"00000000",
  37865=>"00000000",
  37866=>"00000100",
  37867=>"00000100",
  37868=>"11111111",
  37869=>"11111110",
  37870=>"11111110",
  37871=>"11111101",
  37872=>"00000010",
  37873=>"11111110",
  37874=>"00000010",
  37875=>"00000001",
  37876=>"00000100",
  37877=>"11111111",
  37878=>"11111111",
  37879=>"11111111",
  37880=>"11111111",
  37881=>"11111111",
  37882=>"00000001",
  37883=>"00000101",
  37884=>"11111111",
  37885=>"11111110",
  37886=>"00000011",
  37887=>"00000011",
  37888=>"11111111",
  37889=>"11111110",
  37890=>"11111110",
  37891=>"11111111",
  37892=>"00000000",
  37893=>"00000100",
  37894=>"00000000",
  37895=>"11111100",
  37896=>"11111110",
  37897=>"00000000",
  37898=>"00000010",
  37899=>"00000000",
  37900=>"00000001",
  37901=>"00000000",
  37902=>"00000000",
  37903=>"00000001",
  37904=>"00000000",
  37905=>"11111111",
  37906=>"11111100",
  37907=>"00000000",
  37908=>"00000011",
  37909=>"11111111",
  37910=>"00000100",
  37911=>"11111111",
  37912=>"00000001",
  37913=>"00000001",
  37914=>"11111110",
  37915=>"11111100",
  37916=>"11111101",
  37917=>"00000001",
  37918=>"11111101",
  37919=>"11111111",
  37920=>"11111110",
  37921=>"11111111",
  37922=>"00000010",
  37923=>"00000100",
  37924=>"11111101",
  37925=>"00000000",
  37926=>"00000101",
  37927=>"11111111",
  37928=>"00000010",
  37929=>"00000111",
  37930=>"00000000",
  37931=>"11111101",
  37932=>"11111111",
  37933=>"11111111",
  37934=>"00000000",
  37935=>"00000010",
  37936=>"00000000",
  37937=>"00000010",
  37938=>"11111111",
  37939=>"00000000",
  37940=>"00000010",
  37941=>"11111110",
  37942=>"00000001",
  37943=>"00000000",
  37944=>"00000001",
  37945=>"11111100",
  37946=>"00000010",
  37947=>"00000001",
  37948=>"00000100",
  37949=>"00000010",
  37950=>"11111111",
  37951=>"11111110",
  37952=>"11111100",
  37953=>"11111111",
  37954=>"11111111",
  37955=>"11111111",
  37956=>"00000001",
  37957=>"11111100",
  37958=>"11111111",
  37959=>"11111110",
  37960=>"11111101",
  37961=>"11111110",
  37962=>"11111111",
  37963=>"11111111",
  37964=>"11111110",
  37965=>"00000010",
  37966=>"11111101",
  37967=>"11111101",
  37968=>"00000000",
  37969=>"00000000",
  37970=>"11111101",
  37971=>"11111111",
  37972=>"00000001",
  37973=>"00000000",
  37974=>"11111101",
  37975=>"11111111",
  37976=>"11111111",
  37977=>"00000011",
  37978=>"11111110",
  37979=>"11111111",
  37980=>"00000000",
  37981=>"11111110",
  37982=>"00000001",
  37983=>"00000010",
  37984=>"00000000",
  37985=>"00000010",
  37986=>"00000010",
  37987=>"11111110",
  37988=>"00000000",
  37989=>"00000000",
  37990=>"11111111",
  37991=>"00000100",
  37992=>"00000000",
  37993=>"11111100",
  37994=>"00000000",
  37995=>"11111100",
  37996=>"00001000",
  37997=>"11111110",
  37998=>"11111110",
  37999=>"00000001",
  38000=>"00000110",
  38001=>"00000001",
  38002=>"11111101",
  38003=>"11111111",
  38004=>"11111101",
  38005=>"11111111",
  38006=>"00000100",
  38007=>"11111111",
  38008=>"00000111",
  38009=>"00000100",
  38010=>"00000001",
  38011=>"00000001",
  38012=>"00000001",
  38013=>"11111101",
  38014=>"00000000",
  38015=>"00000010",
  38016=>"00000101",
  38017=>"11111111",
  38018=>"11111101",
  38019=>"00000000",
  38020=>"00000010",
  38021=>"00000000",
  38022=>"00000000",
  38023=>"00000010",
  38024=>"00000011",
  38025=>"11111101",
  38026=>"00000001",
  38027=>"00000001",
  38028=>"00000000",
  38029=>"00000011",
  38030=>"11111111",
  38031=>"00000000",
  38032=>"11111111",
  38033=>"11111111",
  38034=>"00000010",
  38035=>"00000001",
  38036=>"11111110",
  38037=>"00000001",
  38038=>"11111101",
  38039=>"00000010",
  38040=>"00000000",
  38041=>"00000111",
  38042=>"11111100",
  38043=>"11111100",
  38044=>"11111101",
  38045=>"00000011",
  38046=>"11111101",
  38047=>"11111100",
  38048=>"11111100",
  38049=>"11111110",
  38050=>"00000101",
  38051=>"00000010",
  38052=>"11111101",
  38053=>"00000011",
  38054=>"00000001",
  38055=>"00000011",
  38056=>"00000010",
  38057=>"11111111",
  38058=>"11111111",
  38059=>"11111100",
  38060=>"11111110",
  38061=>"00000011",
  38062=>"00000001",
  38063=>"00000011",
  38064=>"11111110",
  38065=>"00000001",
  38066=>"00000000",
  38067=>"00000000",
  38068=>"11111101",
  38069=>"00000011",
  38070=>"11111101",
  38071=>"00000110",
  38072=>"00000011",
  38073=>"11111101",
  38074=>"00000101",
  38075=>"00000001",
  38076=>"00000010",
  38077=>"11111101",
  38078=>"00000001",
  38079=>"00000010",
  38080=>"11111111",
  38081=>"11111111",
  38082=>"00000011",
  38083=>"11111110",
  38084=>"11111101",
  38085=>"11111110",
  38086=>"11111100",
  38087=>"00000001",
  38088=>"00000000",
  38089=>"11111111",
  38090=>"00000000",
  38091=>"00000110",
  38092=>"00000000",
  38093=>"11111111",
  38094=>"00000000",
  38095=>"00000001",
  38096=>"00000000",
  38097=>"11111100",
  38098=>"11111111",
  38099=>"11111101",
  38100=>"00000011",
  38101=>"00000000",
  38102=>"00000010",
  38103=>"00000000",
  38104=>"00000010",
  38105=>"00000010",
  38106=>"00000000",
  38107=>"11111110",
  38108=>"00000011",
  38109=>"00000111",
  38110=>"11111101",
  38111=>"11111110",
  38112=>"11111111",
  38113=>"00000101",
  38114=>"00000001",
  38115=>"00000001",
  38116=>"00000011",
  38117=>"00000010",
  38118=>"11111101",
  38119=>"11111111",
  38120=>"00000000",
  38121=>"00000010",
  38122=>"11111110",
  38123=>"11111101",
  38124=>"11111111",
  38125=>"00000100",
  38126=>"00000001",
  38127=>"11111110",
  38128=>"11111100",
  38129=>"11111101",
  38130=>"11111101",
  38131=>"11111100",
  38132=>"00000001",
  38133=>"11111111",
  38134=>"00000001",
  38135=>"11111110",
  38136=>"11111011",
  38137=>"00000011",
  38138=>"00000000",
  38139=>"11111110",
  38140=>"00000010",
  38141=>"00000001",
  38142=>"00000000",
  38143=>"00000000",
  38144=>"11111111",
  38145=>"00000110",
  38146=>"11111011",
  38147=>"11111110",
  38148=>"00000001",
  38149=>"11111100",
  38150=>"00000011",
  38151=>"11111101",
  38152=>"11111110",
  38153=>"11111101",
  38154=>"11111101",
  38155=>"11111110",
  38156=>"11111110",
  38157=>"00000111",
  38158=>"00000000",
  38159=>"11111101",
  38160=>"11111100",
  38161=>"00000001",
  38162=>"00000010",
  38163=>"00000100",
  38164=>"00000110",
  38165=>"11111111",
  38166=>"11111110",
  38167=>"00000001",
  38168=>"11111101",
  38169=>"00000011",
  38170=>"00000100",
  38171=>"11111110",
  38172=>"11111111",
  38173=>"11111111",
  38174=>"00000011",
  38175=>"00000100",
  38176=>"11111110",
  38177=>"00000001",
  38178=>"11111110",
  38179=>"00000010",
  38180=>"00000101",
  38181=>"11111111",
  38182=>"11111101",
  38183=>"11111110",
  38184=>"11111110",
  38185=>"11111101",
  38186=>"11111111",
  38187=>"11111110",
  38188=>"11111110",
  38189=>"11111110",
  38190=>"00000101",
  38191=>"11111111",
  38192=>"00000100",
  38193=>"00000001",
  38194=>"11111101",
  38195=>"00000000",
  38196=>"00000001",
  38197=>"00000000",
  38198=>"00000001",
  38199=>"11111100",
  38200=>"11111110",
  38201=>"00000011",
  38202=>"11111110",
  38203=>"00000001",
  38204=>"00000100",
  38205=>"00000010",
  38206=>"11111110",
  38207=>"00000011",
  38208=>"00000000",
  38209=>"00000001",
  38210=>"00000010",
  38211=>"00000001",
  38212=>"00000000",
  38213=>"00000100",
  38214=>"00000000",
  38215=>"11111101",
  38216=>"11111101",
  38217=>"11111101",
  38218=>"11111111",
  38219=>"11111110",
  38220=>"00000000",
  38221=>"11111111",
  38222=>"11111111",
  38223=>"00000000",
  38224=>"00000100",
  38225=>"11111111",
  38226=>"11111100",
  38227=>"00000011",
  38228=>"00000001",
  38229=>"00000000",
  38230=>"00000100",
  38231=>"00000010",
  38232=>"11111101",
  38233=>"00000100",
  38234=>"11111111",
  38235=>"00000100",
  38236=>"00000011",
  38237=>"11111101",
  38238=>"00000110",
  38239=>"00000000",
  38240=>"11111111",
  38241=>"00000100",
  38242=>"11111101",
  38243=>"00000000",
  38244=>"00000000",
  38245=>"00000001",
  38246=>"00000001",
  38247=>"00000010",
  38248=>"11111101",
  38249=>"11111101",
  38250=>"00000010",
  38251=>"11111111",
  38252=>"00000001",
  38253=>"11111011",
  38254=>"00000100",
  38255=>"00000000",
  38256=>"11111111",
  38257=>"00000010",
  38258=>"11111101",
  38259=>"11111101",
  38260=>"11111110",
  38261=>"00000111",
  38262=>"00000101",
  38263=>"11111111",
  38264=>"00000000",
  38265=>"11111110",
  38266=>"11111111",
  38267=>"00000001",
  38268=>"00000000",
  38269=>"11111110",
  38270=>"11111110",
  38271=>"11111110",
  38272=>"00001000",
  38273=>"00000000",
  38274=>"00000000",
  38275=>"11111111",
  38276=>"11111110",
  38277=>"11111101",
  38278=>"11111101",
  38279=>"11111111",
  38280=>"11111110",
  38281=>"00000100",
  38282=>"00000000",
  38283=>"00000000",
  38284=>"00000010",
  38285=>"11111111",
  38286=>"00000000",
  38287=>"11111110",
  38288=>"11111110",
  38289=>"11111110",
  38290=>"00000001",
  38291=>"00000001",
  38292=>"11111100",
  38293=>"11111111",
  38294=>"11111110",
  38295=>"11111100",
  38296=>"00000100",
  38297=>"11111110",
  38298=>"00000101",
  38299=>"11111111",
  38300=>"00000001",
  38301=>"11111011",
  38302=>"00000000",
  38303=>"11111111",
  38304=>"11111110",
  38305=>"11111110",
  38306=>"11111101",
  38307=>"00000001",
  38308=>"11111110",
  38309=>"11111110",
  38310=>"00000100",
  38311=>"00000001",
  38312=>"11111100",
  38313=>"00000000",
  38314=>"11111110",
  38315=>"00000101",
  38316=>"11111110",
  38317=>"11111110",
  38318=>"11111110",
  38319=>"00000000",
  38320=>"00000001",
  38321=>"11111111",
  38322=>"11111101",
  38323=>"00000100",
  38324=>"00000011",
  38325=>"11111111",
  38326=>"00000111",
  38327=>"00000001",
  38328=>"00000010",
  38329=>"00000001",
  38330=>"11111100",
  38331=>"11111111",
  38332=>"00000000",
  38333=>"00000001",
  38334=>"11111011",
  38335=>"11111110",
  38336=>"00000001",
  38337=>"11111101",
  38338=>"00000000",
  38339=>"11111111",
  38340=>"11111111",
  38341=>"00000110",
  38342=>"00000001",
  38343=>"11111110",
  38344=>"00000101",
  38345=>"00000011",
  38346=>"11111110",
  38347=>"00000010",
  38348=>"00000000",
  38349=>"11111111",
  38350=>"11111111",
  38351=>"11111101",
  38352=>"00000010",
  38353=>"00000010",
  38354=>"00000011",
  38355=>"00000010",
  38356=>"11111101",
  38357=>"00001000",
  38358=>"11111110",
  38359=>"00000100",
  38360=>"00000000",
  38361=>"11111101",
  38362=>"11111111",
  38363=>"11111110",
  38364=>"00000101",
  38365=>"11111111",
  38366=>"00000000",
  38367=>"00000001",
  38368=>"00000000",
  38369=>"11111101",
  38370=>"00000100",
  38371=>"00000010",
  38372=>"11111110",
  38373=>"00000001",
  38374=>"11111110",
  38375=>"00000001",
  38376=>"00000000",
  38377=>"00000001",
  38378=>"00000000",
  38379=>"00000010",
  38380=>"00000010",
  38381=>"11111101",
  38382=>"00000001",
  38383=>"00000010",
  38384=>"00000010",
  38385=>"11111111",
  38386=>"11111111",
  38387=>"00000100",
  38388=>"00000010",
  38389=>"00000000",
  38390=>"00000011",
  38391=>"11111111",
  38392=>"00000111",
  38393=>"11111110",
  38394=>"00000000",
  38395=>"00000010",
  38396=>"00000000",
  38397=>"11111100",
  38398=>"00000001",
  38399=>"11111110",
  38400=>"00000000",
  38401=>"00000000",
  38402=>"11111110",
  38403=>"00000000",
  38404=>"11111111",
  38405=>"11111101",
  38406=>"00000000",
  38407=>"00000010",
  38408=>"00000010",
  38409=>"11111100",
  38410=>"00000000",
  38411=>"00000001",
  38412=>"11111111",
  38413=>"11111111",
  38414=>"11111111",
  38415=>"11111111",
  38416=>"11111101",
  38417=>"00000010",
  38418=>"11111101",
  38419=>"00000010",
  38420=>"11111110",
  38421=>"11111101",
  38422=>"11111110",
  38423=>"11111111",
  38424=>"11111101",
  38425=>"00000010",
  38426=>"11111111",
  38427=>"00000100",
  38428=>"11111110",
  38429=>"11111100",
  38430=>"11111100",
  38431=>"00000010",
  38432=>"00000010",
  38433=>"11111100",
  38434=>"11111111",
  38435=>"00000010",
  38436=>"00000000",
  38437=>"11111101",
  38438=>"00000001",
  38439=>"11111101",
  38440=>"11111110",
  38441=>"11111101",
  38442=>"00000011",
  38443=>"00000010",
  38444=>"11111110",
  38445=>"00000011",
  38446=>"00000010",
  38447=>"11111110",
  38448=>"11111011",
  38449=>"11111110",
  38450=>"11111110",
  38451=>"11111110",
  38452=>"11111101",
  38453=>"00000000",
  38454=>"00000101",
  38455=>"11111110",
  38456=>"00000001",
  38457=>"11111110",
  38458=>"11111110",
  38459=>"00000000",
  38460=>"11111111",
  38461=>"11111101",
  38462=>"11111110",
  38463=>"00000011",
  38464=>"11111111",
  38465=>"00000100",
  38466=>"00000101",
  38467=>"00000010",
  38468=>"00000101",
  38469=>"00000000",
  38470=>"00000001",
  38471=>"11111101",
  38472=>"00000000",
  38473=>"00000001",
  38474=>"00000010",
  38475=>"11111101",
  38476=>"00000111",
  38477=>"00000001",
  38478=>"00000010",
  38479=>"00000011",
  38480=>"11111111",
  38481=>"00000111",
  38482=>"11111110",
  38483=>"00000001",
  38484=>"11111111",
  38485=>"11111101",
  38486=>"00000011",
  38487=>"00000011",
  38488=>"00000001",
  38489=>"11111101",
  38490=>"00000000",
  38491=>"00000001",
  38492=>"11111110",
  38493=>"11111101",
  38494=>"00000011",
  38495=>"00000010",
  38496=>"00000000",
  38497=>"00000001",
  38498=>"11111110",
  38499=>"00000010",
  38500=>"11111110",
  38501=>"00000100",
  38502=>"00000011",
  38503=>"00000010",
  38504=>"00000010",
  38505=>"00000010",
  38506=>"00000011",
  38507=>"11111110",
  38508=>"11111111",
  38509=>"00000010",
  38510=>"11111110",
  38511=>"11111100",
  38512=>"00000000",
  38513=>"00000001",
  38514=>"00000001",
  38515=>"11111101",
  38516=>"00000011",
  38517=>"00000001",
  38518=>"11111101",
  38519=>"00000010",
  38520=>"00000000",
  38521=>"00000000",
  38522=>"11111111",
  38523=>"11111101",
  38524=>"00000001",
  38525=>"11111110",
  38526=>"00000011",
  38527=>"00000001",
  38528=>"00000100",
  38529=>"00000001",
  38530=>"00000010",
  38531=>"11111100",
  38532=>"00000000",
  38533=>"00000001",
  38534=>"00000010",
  38535=>"11111100",
  38536=>"11111110",
  38537=>"00000010",
  38538=>"11111111",
  38539=>"00000001",
  38540=>"11111111",
  38541=>"00000001",
  38542=>"00000000",
  38543=>"11111110",
  38544=>"00000000",
  38545=>"11111110",
  38546=>"11111101",
  38547=>"00000000",
  38548=>"00000001",
  38549=>"11111101",
  38550=>"00000100",
  38551=>"00000001",
  38552=>"00000010",
  38553=>"11111101",
  38554=>"00000011",
  38555=>"00000000",
  38556=>"00000011",
  38557=>"00000000",
  38558=>"00000001",
  38559=>"11111111",
  38560=>"00000001",
  38561=>"00000011",
  38562=>"00000000",
  38563=>"00000000",
  38564=>"11111111",
  38565=>"11111110",
  38566=>"00000000",
  38567=>"00000001",
  38568=>"11111111",
  38569=>"11111101",
  38570=>"11111100",
  38571=>"00000100",
  38572=>"00000010",
  38573=>"00000010",
  38574=>"00000010",
  38575=>"00000001",
  38576=>"00000011",
  38577=>"11111011",
  38578=>"00000001",
  38579=>"00000010",
  38580=>"11111110",
  38581=>"00000010",
  38582=>"11111111",
  38583=>"11111101",
  38584=>"11111110",
  38585=>"11111101",
  38586=>"11111110",
  38587=>"00000010",
  38588=>"00000001",
  38589=>"00000010",
  38590=>"00000000",
  38591=>"11111110",
  38592=>"11111101",
  38593=>"00000100",
  38594=>"00000100",
  38595=>"11111111",
  38596=>"00000000",
  38597=>"00000010",
  38598=>"00000011",
  38599=>"11111011",
  38600=>"11111111",
  38601=>"00000010",
  38602=>"00000001",
  38603=>"11111111",
  38604=>"11111111",
  38605=>"00000101",
  38606=>"00000100",
  38607=>"11111111",
  38608=>"00000011",
  38609=>"00000010",
  38610=>"11111101",
  38611=>"00000010",
  38612=>"00000000",
  38613=>"11111111",
  38614=>"00000000",
  38615=>"00000011",
  38616=>"00000001",
  38617=>"00000011",
  38618=>"00000001",
  38619=>"00000010",
  38620=>"11111110",
  38621=>"11111101",
  38622=>"11111101",
  38623=>"11111111",
  38624=>"11111101",
  38625=>"00000010",
  38626=>"00000001",
  38627=>"00000001",
  38628=>"11111111",
  38629=>"00000000",
  38630=>"00000011",
  38631=>"00000010",
  38632=>"00000010",
  38633=>"11111111",
  38634=>"11111100",
  38635=>"11111111",
  38636=>"11111111",
  38637=>"11111101",
  38638=>"00000001",
  38639=>"00000000",
  38640=>"00000010",
  38641=>"00000011",
  38642=>"00000001",
  38643=>"00000000",
  38644=>"00000000",
  38645=>"00000001",
  38646=>"11111111",
  38647=>"11111100",
  38648=>"11111111",
  38649=>"11111101",
  38650=>"00000010",
  38651=>"11111101",
  38652=>"11111101",
  38653=>"00000001",
  38654=>"00000011",
  38655=>"11111110",
  38656=>"00000000",
  38657=>"00000001",
  38658=>"00000010",
  38659=>"11111100",
  38660=>"11111110",
  38661=>"11111110",
  38662=>"00000001",
  38663=>"11111101",
  38664=>"00000010",
  38665=>"00000010",
  38666=>"00000000",
  38667=>"11111101",
  38668=>"00000011",
  38669=>"11111111",
  38670=>"00000000",
  38671=>"00000010",
  38672=>"00000000",
  38673=>"11111110",
  38674=>"11111110",
  38675=>"00000100",
  38676=>"00000000",
  38677=>"00000000",
  38678=>"00000011",
  38679=>"00000001",
  38680=>"00000010",
  38681=>"00000001",
  38682=>"00000010",
  38683=>"00000011",
  38684=>"00000000",
  38685=>"11111110",
  38686=>"00000100",
  38687=>"11111111",
  38688=>"00000001",
  38689=>"11111111",
  38690=>"11111111",
  38691=>"11111110",
  38692=>"00000001",
  38693=>"11111101",
  38694=>"11111110",
  38695=>"00000010",
  38696=>"00001000",
  38697=>"00000000",
  38698=>"00000101",
  38699=>"00000010",
  38700=>"11111111",
  38701=>"11111111",
  38702=>"00000010",
  38703=>"00000000",
  38704=>"00000010",
  38705=>"11111100",
  38706=>"00000001",
  38707=>"11111111",
  38708=>"00000010",
  38709=>"00000000",
  38710=>"00000010",
  38711=>"00000001",
  38712=>"11111111",
  38713=>"00000001",
  38714=>"11111101",
  38715=>"00000101",
  38716=>"11111101",
  38717=>"11111101",
  38718=>"11111110",
  38719=>"00000100",
  38720=>"00000000",
  38721=>"00000000",
  38722=>"00000001",
  38723=>"11111111",
  38724=>"00000000",
  38725=>"11111100",
  38726=>"11111110",
  38727=>"00000001",
  38728=>"00000011",
  38729=>"00000010",
  38730=>"11111111",
  38731=>"00000000",
  38732=>"11111111",
  38733=>"11111110",
  38734=>"11111100",
  38735=>"11111110",
  38736=>"00000010",
  38737=>"11111101",
  38738=>"11111111",
  38739=>"11111100",
  38740=>"00000001",
  38741=>"00000000",
  38742=>"00000000",
  38743=>"00000101",
  38744=>"11111110",
  38745=>"00000000",
  38746=>"00000010",
  38747=>"11111111",
  38748=>"00000000",
  38749=>"00000101",
  38750=>"11111101",
  38751=>"11111101",
  38752=>"11111111",
  38753=>"11111100",
  38754=>"00000000",
  38755=>"11111100",
  38756=>"11111101",
  38757=>"00000000",
  38758=>"00000000",
  38759=>"00000000",
  38760=>"11111111",
  38761=>"11111101",
  38762=>"11111111",
  38763=>"11111111",
  38764=>"00000000",
  38765=>"00000001",
  38766=>"00000000",
  38767=>"00000010",
  38768=>"00000001",
  38769=>"00000110",
  38770=>"11111101",
  38771=>"11111101",
  38772=>"00000000",
  38773=>"00000000",
  38774=>"00000000",
  38775=>"00000001",
  38776=>"11111101",
  38777=>"11111101",
  38778=>"11111110",
  38779=>"00000101",
  38780=>"11111100",
  38781=>"11111111",
  38782=>"11111100",
  38783=>"11111111",
  38784=>"11111111",
  38785=>"00000011",
  38786=>"00000010",
  38787=>"00000010",
  38788=>"11111111",
  38789=>"00000000",
  38790=>"11111111",
  38791=>"11111101",
  38792=>"00000001",
  38793=>"11111111",
  38794=>"11111111",
  38795=>"11111111",
  38796=>"11111101",
  38797=>"00000010",
  38798=>"11111100",
  38799=>"00000010",
  38800=>"00000001",
  38801=>"11111100",
  38802=>"00000010",
  38803=>"11111101",
  38804=>"00000000",
  38805=>"11111111",
  38806=>"00000001",
  38807=>"00000010",
  38808=>"11111111",
  38809=>"11111101",
  38810=>"00000001",
  38811=>"00000001",
  38812=>"00000000",
  38813=>"00000001",
  38814=>"00000011",
  38815=>"00000001",
  38816=>"11111111",
  38817=>"11111111",
  38818=>"11111111",
  38819=>"00000010",
  38820=>"00000010",
  38821=>"11111110",
  38822=>"00000100",
  38823=>"11111110",
  38824=>"11111110",
  38825=>"11111101",
  38826=>"11111111",
  38827=>"11111110",
  38828=>"00000100",
  38829=>"00000001",
  38830=>"00000011",
  38831=>"11111110",
  38832=>"00000000",
  38833=>"00000010",
  38834=>"11111110",
  38835=>"11111111",
  38836=>"11111110",
  38837=>"00000010",
  38838=>"11111110",
  38839=>"11111111",
  38840=>"00000001",
  38841=>"00000011",
  38842=>"00000010",
  38843=>"11111101",
  38844=>"00000000",
  38845=>"00000001",
  38846=>"00000011",
  38847=>"11111101",
  38848=>"00000000",
  38849=>"11111110",
  38850=>"00000010",
  38851=>"11111101",
  38852=>"00000001",
  38853=>"00000000",
  38854=>"11111111",
  38855=>"00000010",
  38856=>"00000101",
  38857=>"11111101",
  38858=>"11111101",
  38859=>"11111111",
  38860=>"00000001",
  38861=>"11111101",
  38862=>"00000100",
  38863=>"00000001",
  38864=>"00000010",
  38865=>"11111101",
  38866=>"11111101",
  38867=>"11111101",
  38868=>"11111111",
  38869=>"00000000",
  38870=>"00000000",
  38871=>"11111101",
  38872=>"00000000",
  38873=>"11111111",
  38874=>"11111100",
  38875=>"11111101",
  38876=>"11111101",
  38877=>"11111110",
  38878=>"11111110",
  38879=>"11111111",
  38880=>"00000000",
  38881=>"11111101",
  38882=>"00000000",
  38883=>"11111101",
  38884=>"00000001",
  38885=>"11111110",
  38886=>"11111101",
  38887=>"00000001",
  38888=>"11111111",
  38889=>"11111110",
  38890=>"11111011",
  38891=>"00000011",
  38892=>"11111101",
  38893=>"00000011",
  38894=>"11111110",
  38895=>"11111110",
  38896=>"00000001",
  38897=>"11111110",
  38898=>"11111110",
  38899=>"00000010",
  38900=>"00000001",
  38901=>"00000010",
  38902=>"00000000",
  38903=>"11111111",
  38904=>"11111111",
  38905=>"00000000",
  38906=>"11111110",
  38907=>"00000001",
  38908=>"00000011",
  38909=>"00000000",
  38910=>"11111100",
  38911=>"11111101",
  38912=>"00000011",
  38913=>"00000101",
  38914=>"11111110",
  38915=>"00000011",
  38916=>"11111101",
  38917=>"11111110",
  38918=>"11111111",
  38919=>"00000011",
  38920=>"11111110",
  38921=>"11111101",
  38922=>"11111110",
  38923=>"00000010",
  38924=>"11111101",
  38925=>"11111101",
  38926=>"00000011",
  38927=>"11111101",
  38928=>"11111110",
  38929=>"11111100",
  38930=>"11111111",
  38931=>"11111100",
  38932=>"00000010",
  38933=>"11111110",
  38934=>"11111101",
  38935=>"11111110",
  38936=>"00000011",
  38937=>"00000101",
  38938=>"00000101",
  38939=>"00000011",
  38940=>"00000001",
  38941=>"00001000",
  38942=>"00000101",
  38943=>"11111101",
  38944=>"00000010",
  38945=>"11111100",
  38946=>"00000100",
  38947=>"00000100",
  38948=>"00000000",
  38949=>"11111101",
  38950=>"00000000",
  38951=>"00000010",
  38952=>"00000001",
  38953=>"00000010",
  38954=>"11111110",
  38955=>"00000010",
  38956=>"00000100",
  38957=>"11111110",
  38958=>"00000000",
  38959=>"00000000",
  38960=>"11111101",
  38961=>"11111111",
  38962=>"00000010",
  38963=>"00000100",
  38964=>"11111111",
  38965=>"11111100",
  38966=>"11111110",
  38967=>"11111100",
  38968=>"00000010",
  38969=>"11111101",
  38970=>"00000110",
  38971=>"00000011",
  38972=>"11111101",
  38973=>"00000001",
  38974=>"00000011",
  38975=>"00000010",
  38976=>"00000100",
  38977=>"00000001",
  38978=>"00000011",
  38979=>"11111111",
  38980=>"00000011",
  38981=>"00000000",
  38982=>"00000111",
  38983=>"11111100",
  38984=>"11111111",
  38985=>"11111101",
  38986=>"00000100",
  38987=>"11111101",
  38988=>"11111101",
  38989=>"11111111",
  38990=>"11111111",
  38991=>"00000000",
  38992=>"11111111",
  38993=>"11111101",
  38994=>"11111111",
  38995=>"00000011",
  38996=>"00000000",
  38997=>"11111100",
  38998=>"11111110",
  38999=>"11111111",
  39000=>"00000010",
  39001=>"11111001",
  39002=>"00000000",
  39003=>"11111111",
  39004=>"00000010",
  39005=>"11111110",
  39006=>"11111111",
  39007=>"00000011",
  39008=>"00000010",
  39009=>"11111111",
  39010=>"00000101",
  39011=>"00000000",
  39012=>"00000001",
  39013=>"00000010",
  39014=>"00000010",
  39015=>"00000011",
  39016=>"00000110",
  39017=>"00000001",
  39018=>"00000011",
  39019=>"11111101",
  39020=>"00000010",
  39021=>"00000000",
  39022=>"11111111",
  39023=>"11111011",
  39024=>"11111110",
  39025=>"00000000",
  39026=>"00000100",
  39027=>"00000000",
  39028=>"00000100",
  39029=>"00000101",
  39030=>"11111110",
  39031=>"11111111",
  39032=>"00000011",
  39033=>"00000010",
  39034=>"00000011",
  39035=>"00000011",
  39036=>"11111100",
  39037=>"11111101",
  39038=>"00000000",
  39039=>"00000001",
  39040=>"11111110",
  39041=>"11111101",
  39042=>"11111100",
  39043=>"00000011",
  39044=>"11111101",
  39045=>"00000110",
  39046=>"00000000",
  39047=>"00000001",
  39048=>"11111100",
  39049=>"11111101",
  39050=>"11111110",
  39051=>"11111101",
  39052=>"11111110",
  39053=>"00000011",
  39054=>"11111110",
  39055=>"00000011",
  39056=>"11111111",
  39057=>"11111100",
  39058=>"11111110",
  39059=>"00000000",
  39060=>"11111101",
  39061=>"00000011",
  39062=>"00000001",
  39063=>"11111101",
  39064=>"00000010",
  39065=>"11111110",
  39066=>"00000011",
  39067=>"00000011",
  39068=>"00000000",
  39069=>"11111110",
  39070=>"00000000",
  39071=>"00000101",
  39072=>"00000000",
  39073=>"00000010",
  39074=>"00000001",
  39075=>"00000010",
  39076=>"00000001",
  39077=>"11111101",
  39078=>"00000101",
  39079=>"11111110",
  39080=>"00000001",
  39081=>"11111110",
  39082=>"11111111",
  39083=>"00000100",
  39084=>"00000011",
  39085=>"00000000",
  39086=>"11111110",
  39087=>"11111110",
  39088=>"00000011",
  39089=>"00000011",
  39090=>"11111101",
  39091=>"00000011",
  39092=>"00000010",
  39093=>"00000001",
  39094=>"11111100",
  39095=>"00000000",
  39096=>"11111110",
  39097=>"00000100",
  39098=>"11111110",
  39099=>"00000010",
  39100=>"11111011",
  39101=>"00000011",
  39102=>"00000010",
  39103=>"00000001",
  39104=>"00000000",
  39105=>"00000000",
  39106=>"11111111",
  39107=>"11111110",
  39108=>"11111111",
  39109=>"00000000",
  39110=>"00000001",
  39111=>"00000010",
  39112=>"11111110",
  39113=>"00000001",
  39114=>"00000000",
  39115=>"11111101",
  39116=>"00000001",
  39117=>"00000011",
  39118=>"00000000",
  39119=>"11111110",
  39120=>"00000011",
  39121=>"00000001",
  39122=>"11111110",
  39123=>"00000000",
  39124=>"11111110",
  39125=>"11111101",
  39126=>"00000100",
  39127=>"00000001",
  39128=>"11111111",
  39129=>"11111110",
  39130=>"00000000",
  39131=>"11111100",
  39132=>"11111110",
  39133=>"00000100",
  39134=>"11111100",
  39135=>"00000011",
  39136=>"11111111",
  39137=>"00000000",
  39138=>"00000010",
  39139=>"00000001",
  39140=>"11111111",
  39141=>"00000001",
  39142=>"11111100",
  39143=>"00000101",
  39144=>"11111110",
  39145=>"00000001",
  39146=>"11111101",
  39147=>"00000000",
  39148=>"11111111",
  39149=>"11111110",
  39150=>"00000101",
  39151=>"11111101",
  39152=>"00000010",
  39153=>"11111101",
  39154=>"00000001",
  39155=>"00000100",
  39156=>"11111110",
  39157=>"00000000",
  39158=>"00000001",
  39159=>"11111111",
  39160=>"00000000",
  39161=>"00000100",
  39162=>"00000000",
  39163=>"00000001",
  39164=>"00000000",
  39165=>"00000010",
  39166=>"11111111",
  39167=>"00000110",
  39168=>"11111101",
  39169=>"11111101",
  39170=>"00000001",
  39171=>"00000101",
  39172=>"00000001",
  39173=>"00000001",
  39174=>"00000011",
  39175=>"00000011",
  39176=>"11111101",
  39177=>"00000011",
  39178=>"11111100",
  39179=>"00000001",
  39180=>"00000011",
  39181=>"00000000",
  39182=>"00000000",
  39183=>"11111110",
  39184=>"00000000",
  39185=>"00000101",
  39186=>"11111111",
  39187=>"00000000",
  39188=>"00000000",
  39189=>"00000011",
  39190=>"00000110",
  39191=>"00000010",
  39192=>"00000011",
  39193=>"00000000",
  39194=>"11111110",
  39195=>"11111111",
  39196=>"00000011",
  39197=>"00000001",
  39198=>"00000001",
  39199=>"11111011",
  39200=>"00000010",
  39201=>"00000101",
  39202=>"00000001",
  39203=>"11111111",
  39204=>"00000001",
  39205=>"11111101",
  39206=>"11111100",
  39207=>"00000110",
  39208=>"11111100",
  39209=>"11111110",
  39210=>"11111111",
  39211=>"11111100",
  39212=>"00000100",
  39213=>"00000001",
  39214=>"00000011",
  39215=>"00000100",
  39216=>"00000000",
  39217=>"00000000",
  39218=>"00000001",
  39219=>"00000010",
  39220=>"11111101",
  39221=>"11111110",
  39222=>"00000001",
  39223=>"00000001",
  39224=>"00000010",
  39225=>"11111100",
  39226=>"11111101",
  39227=>"00000001",
  39228=>"00000011",
  39229=>"00000001",
  39230=>"00000000",
  39231=>"11111111",
  39232=>"11111111",
  39233=>"11111111",
  39234=>"00000001",
  39235=>"00000100",
  39236=>"00000110",
  39237=>"00000001",
  39238=>"00000001",
  39239=>"11111111",
  39240=>"11111101",
  39241=>"00000011",
  39242=>"00000010",
  39243=>"00000010",
  39244=>"11111101",
  39245=>"11111111",
  39246=>"00000010",
  39247=>"00000010",
  39248=>"11111111",
  39249=>"11111110",
  39250=>"11111111",
  39251=>"00000000",
  39252=>"00000000",
  39253=>"11111101",
  39254=>"11111101",
  39255=>"11111100",
  39256=>"00000010",
  39257=>"11111100",
  39258=>"00000100",
  39259=>"00000100",
  39260=>"00000000",
  39261=>"11111111",
  39262=>"11111101",
  39263=>"00000010",
  39264=>"00000010",
  39265=>"00000011",
  39266=>"00000011",
  39267=>"00000001",
  39268=>"00000001",
  39269=>"00000001",
  39270=>"00000001",
  39271=>"00000010",
  39272=>"00000000",
  39273=>"11111111",
  39274=>"00000000",
  39275=>"00000000",
  39276=>"11111110",
  39277=>"11111011",
  39278=>"11111110",
  39279=>"00000101",
  39280=>"11111111",
  39281=>"00000110",
  39282=>"00000000",
  39283=>"00000100",
  39284=>"11111111",
  39285=>"00000010",
  39286=>"00000001",
  39287=>"00000001",
  39288=>"00000011",
  39289=>"00000000",
  39290=>"00000001",
  39291=>"00000001",
  39292=>"00000011",
  39293=>"11111111",
  39294=>"11111111",
  39295=>"11111111",
  39296=>"11111110",
  39297=>"11111110",
  39298=>"00000010",
  39299=>"00000011",
  39300=>"00000001",
  39301=>"00000000",
  39302=>"00000001",
  39303=>"00000011",
  39304=>"00000100",
  39305=>"00000000",
  39306=>"11111111",
  39307=>"00000000",
  39308=>"00000010",
  39309=>"00000100",
  39310=>"11111111",
  39311=>"11111110",
  39312=>"00000001",
  39313=>"00000011",
  39314=>"00000010",
  39315=>"00000011",
  39316=>"11111110",
  39317=>"00000011",
  39318=>"11111111",
  39319=>"11111101",
  39320=>"00000101",
  39321=>"11111111",
  39322=>"00000001",
  39323=>"11111111",
  39324=>"00000011",
  39325=>"00000011",
  39326=>"00000100",
  39327=>"11111110",
  39328=>"00000010",
  39329=>"00000001",
  39330=>"00000011",
  39331=>"00000000",
  39332=>"11111111",
  39333=>"11111011",
  39334=>"11111101",
  39335=>"00000101",
  39336=>"00000011",
  39337=>"11111110",
  39338=>"11111110",
  39339=>"00000001",
  39340=>"11111011",
  39341=>"11111111",
  39342=>"00000000",
  39343=>"00000011",
  39344=>"11111110",
  39345=>"11111111",
  39346=>"00000010",
  39347=>"11111111",
  39348=>"00000101",
  39349=>"00000010",
  39350=>"00000000",
  39351=>"00000011",
  39352=>"11111101",
  39353=>"11111110",
  39354=>"00000001",
  39355=>"00000001",
  39356=>"00000010",
  39357=>"00000000",
  39358=>"11111110",
  39359=>"00000000",
  39360=>"00000001",
  39361=>"11111101",
  39362=>"00000100",
  39363=>"11111111",
  39364=>"11111110",
  39365=>"00000100",
  39366=>"11111111",
  39367=>"00000100",
  39368=>"11111111",
  39369=>"11111111",
  39370=>"11111111",
  39371=>"11111111",
  39372=>"00000100",
  39373=>"00000100",
  39374=>"11111101",
  39375=>"11111110",
  39376=>"11111111",
  39377=>"00000000",
  39378=>"00000010",
  39379=>"00000001",
  39380=>"11111111",
  39381=>"00000000",
  39382=>"00000000",
  39383=>"11111111",
  39384=>"00000001",
  39385=>"00000011",
  39386=>"00000011",
  39387=>"00000010",
  39388=>"00000010",
  39389=>"00000100",
  39390=>"11111101",
  39391=>"11111111",
  39392=>"00000101",
  39393=>"00000101",
  39394=>"11111100",
  39395=>"11111110",
  39396=>"00000010",
  39397=>"11111110",
  39398=>"00000100",
  39399=>"11111110",
  39400=>"00000010",
  39401=>"00000000",
  39402=>"11111101",
  39403=>"00000011",
  39404=>"00000000",
  39405=>"11111110",
  39406=>"11111011",
  39407=>"00000001",
  39408=>"00000011",
  39409=>"00000110",
  39410=>"00000000",
  39411=>"11111110",
  39412=>"00000001",
  39413=>"00000001",
  39414=>"00000010",
  39415=>"11111101",
  39416=>"11111110",
  39417=>"11111110",
  39418=>"00000001",
  39419=>"11111100",
  39420=>"00000001",
  39421=>"00000001",
  39422=>"11111111",
  39423=>"11111101",
  39424=>"00000000",
  39425=>"00000011",
  39426=>"11111110",
  39427=>"11111110",
  39428=>"11111100",
  39429=>"00000000",
  39430=>"11111101",
  39431=>"11111101",
  39432=>"00000010",
  39433=>"00000110",
  39434=>"11111110",
  39435=>"11111101",
  39436=>"11111111",
  39437=>"11111101",
  39438=>"00000101",
  39439=>"11111111",
  39440=>"11111110",
  39441=>"11111011",
  39442=>"00000000",
  39443=>"00000001",
  39444=>"00000101",
  39445=>"00000001",
  39446=>"00000100",
  39447=>"00000101",
  39448=>"00000001",
  39449=>"11111111",
  39450=>"11111111",
  39451=>"11111111",
  39452=>"00000101",
  39453=>"00000011",
  39454=>"00000000",
  39455=>"00000001",
  39456=>"11111110",
  39457=>"00000100",
  39458=>"00000010",
  39459=>"00000001",
  39460=>"00000001",
  39461=>"11111100",
  39462=>"00000001",
  39463=>"11111101",
  39464=>"00000110",
  39465=>"00000000",
  39466=>"00000001",
  39467=>"11111101",
  39468=>"00000100",
  39469=>"11111111",
  39470=>"00000000",
  39471=>"00000100",
  39472=>"00000010",
  39473=>"11111110",
  39474=>"00000001",
  39475=>"00000000",
  39476=>"00000000",
  39477=>"00000000",
  39478=>"11111110",
  39479=>"11111111",
  39480=>"00000010",
  39481=>"00000010",
  39482=>"11111111",
  39483=>"00000001",
  39484=>"11111111",
  39485=>"00000100",
  39486=>"11111111",
  39487=>"00000100",
  39488=>"00000000",
  39489=>"00000001",
  39490=>"11111101",
  39491=>"11111100",
  39492=>"00000011",
  39493=>"00000001",
  39494=>"00000000",
  39495=>"00000100",
  39496=>"11111110",
  39497=>"11111101",
  39498=>"00000000",
  39499=>"11111110",
  39500=>"00000001",
  39501=>"00000011",
  39502=>"11111101",
  39503=>"11111101",
  39504=>"00000100",
  39505=>"00000011",
  39506=>"00000000",
  39507=>"11111111",
  39508=>"11111011",
  39509=>"00000011",
  39510=>"11111110",
  39511=>"00000011",
  39512=>"11111111",
  39513=>"00000010",
  39514=>"00000001",
  39515=>"00000001",
  39516=>"11111111",
  39517=>"00000010",
  39518=>"11111111",
  39519=>"00000000",
  39520=>"00000001",
  39521=>"00000000",
  39522=>"00000001",
  39523=>"11111110",
  39524=>"00000000",
  39525=>"00000000",
  39526=>"00000001",
  39527=>"00000100",
  39528=>"11111110",
  39529=>"11111111",
  39530=>"00000011",
  39531=>"00000010",
  39532=>"11111110",
  39533=>"11111011",
  39534=>"00000011",
  39535=>"11111101",
  39536=>"00000001",
  39537=>"11111110",
  39538=>"00000000",
  39539=>"00000110",
  39540=>"11111100",
  39541=>"00000011",
  39542=>"00000000",
  39543=>"00000001",
  39544=>"00000000",
  39545=>"11111101",
  39546=>"00000010",
  39547=>"00000011",
  39548=>"00000010",
  39549=>"11111110",
  39550=>"11111101",
  39551=>"11111111",
  39552=>"00000000",
  39553=>"00000100",
  39554=>"00000010",
  39555=>"00000110",
  39556=>"11111101",
  39557=>"11111010",
  39558=>"00000011",
  39559=>"11111101",
  39560=>"00000010",
  39561=>"00000001",
  39562=>"00000100",
  39563=>"00000011",
  39564=>"00000001",
  39565=>"00000001",
  39566=>"00000100",
  39567=>"11111111",
  39568=>"00000011",
  39569=>"00000000",
  39570=>"11111111",
  39571=>"00000001",
  39572=>"00000010",
  39573=>"00000110",
  39574=>"11111101",
  39575=>"11111101",
  39576=>"11111111",
  39577=>"00000101",
  39578=>"11111110",
  39579=>"11111110",
  39580=>"11111100",
  39581=>"00000100",
  39582=>"11111111",
  39583=>"00000011",
  39584=>"00000001",
  39585=>"11111101",
  39586=>"00000001",
  39587=>"00000010",
  39588=>"11111111",
  39589=>"00000001",
  39590=>"00000110",
  39591=>"00000010",
  39592=>"11111100",
  39593=>"00000010",
  39594=>"00000000",
  39595=>"00000010",
  39596=>"11111111",
  39597=>"11111111",
  39598=>"11111111",
  39599=>"11111100",
  39600=>"00000010",
  39601=>"00000000",
  39602=>"00000101",
  39603=>"00000011",
  39604=>"00000000",
  39605=>"11111011",
  39606=>"11111110",
  39607=>"00000010",
  39608=>"11111110",
  39609=>"00000000",
  39610=>"00000010",
  39611=>"11111101",
  39612=>"11111101",
  39613=>"00000000",
  39614=>"00000101",
  39615=>"00000011",
  39616=>"00000000",
  39617=>"00000000",
  39618=>"00000000",
  39619=>"11111110",
  39620=>"00000100",
  39621=>"11111110",
  39622=>"11111110",
  39623=>"00000101",
  39624=>"00000110",
  39625=>"00000011",
  39626=>"00000010",
  39627=>"00000000",
  39628=>"11111111",
  39629=>"11111111",
  39630=>"00000000",
  39631=>"00000010",
  39632=>"00000000",
  39633=>"11111101",
  39634=>"00000011",
  39635=>"00000001",
  39636=>"00000000",
  39637=>"00000001",
  39638=>"00000001",
  39639=>"00000000",
  39640=>"11111110",
  39641=>"11111111",
  39642=>"00000000",
  39643=>"11111101",
  39644=>"00000010",
  39645=>"00000000",
  39646=>"11111100",
  39647=>"00000010",
  39648=>"00000100",
  39649=>"00000000",
  39650=>"00000000",
  39651=>"00000011",
  39652=>"00000011",
  39653=>"11111111",
  39654=>"00000011",
  39655=>"00000101",
  39656=>"00000001",
  39657=>"11111110",
  39658=>"11111101",
  39659=>"00000000",
  39660=>"11111101",
  39661=>"00000001",
  39662=>"00000001",
  39663=>"11111110",
  39664=>"00000101",
  39665=>"00000011",
  39666=>"11111101",
  39667=>"11111101",
  39668=>"00000000",
  39669=>"11111110",
  39670=>"00000010",
  39671=>"00000000",
  39672=>"00000010",
  39673=>"11111101",
  39674=>"00000010",
  39675=>"00000000",
  39676=>"00000001",
  39677=>"11111100",
  39678=>"11111101",
  39679=>"00000000",
  39680=>"00000010",
  39681=>"11111110",
  39682=>"00000100",
  39683=>"00000001",
  39684=>"11111110",
  39685=>"00000001",
  39686=>"00000000",
  39687=>"00000111",
  39688=>"00000000",
  39689=>"00000100",
  39690=>"11111111",
  39691=>"00000100",
  39692=>"11111101",
  39693=>"00000010",
  39694=>"11111110",
  39695=>"00000011",
  39696=>"00000100",
  39697=>"11111101",
  39698=>"11111100",
  39699=>"00000000",
  39700=>"00000010",
  39701=>"00000001",
  39702=>"00000110",
  39703=>"11111111",
  39704=>"00000000",
  39705=>"00000010",
  39706=>"11111110",
  39707=>"00000111",
  39708=>"00000001",
  39709=>"00000000",
  39710=>"11111110",
  39711=>"00000000",
  39712=>"00000100",
  39713=>"11111011",
  39714=>"00000010",
  39715=>"11111110",
  39716=>"00000000",
  39717=>"11111100",
  39718=>"00000011",
  39719=>"11111111",
  39720=>"00000011",
  39721=>"00000110",
  39722=>"00000101",
  39723=>"00000100",
  39724=>"00000010",
  39725=>"00000011",
  39726=>"00000100",
  39727=>"11111111",
  39728=>"11111101",
  39729=>"00000101",
  39730=>"00000011",
  39731=>"00000000",
  39732=>"00000000",
  39733=>"00000010",
  39734=>"00000100",
  39735=>"11111101",
  39736=>"11111111",
  39737=>"11111110",
  39738=>"11111110",
  39739=>"11111100",
  39740=>"00000000",
  39741=>"11111110",
  39742=>"11111111",
  39743=>"00000010",
  39744=>"11111101",
  39745=>"00000000",
  39746=>"11111111",
  39747=>"00000001",
  39748=>"00000100",
  39749=>"00000001",
  39750=>"00000101",
  39751=>"00000001",
  39752=>"11111110",
  39753=>"00000100",
  39754=>"00000000",
  39755=>"11111011",
  39756=>"00000100",
  39757=>"00000000",
  39758=>"11111111",
  39759=>"00000100",
  39760=>"11111111",
  39761=>"11111110",
  39762=>"11111101",
  39763=>"00000011",
  39764=>"00000011",
  39765=>"11111101",
  39766=>"00000010",
  39767=>"11111011",
  39768=>"00000001",
  39769=>"00000001",
  39770=>"00000001",
  39771=>"11111100",
  39772=>"00000100",
  39773=>"00000000",
  39774=>"00000010",
  39775=>"11111111",
  39776=>"11111101",
  39777=>"11111101",
  39778=>"00000011",
  39779=>"00000010",
  39780=>"11111111",
  39781=>"00000011",
  39782=>"00000000",
  39783=>"00000000",
  39784=>"00000000",
  39785=>"00000010",
  39786=>"00000100",
  39787=>"11111110",
  39788=>"11111101",
  39789=>"11111110",
  39790=>"00000010",
  39791=>"00000010",
  39792=>"11111111",
  39793=>"00000010",
  39794=>"00000100",
  39795=>"11111111",
  39796=>"11111110",
  39797=>"00000000",
  39798=>"11111100",
  39799=>"00000001",
  39800=>"00000000",
  39801=>"11111101",
  39802=>"00000011",
  39803=>"11111111",
  39804=>"11111110",
  39805=>"11111111",
  39806=>"00000000",
  39807=>"11111111",
  39808=>"00000001",
  39809=>"00000010",
  39810=>"00000011",
  39811=>"00000100",
  39812=>"11111110",
  39813=>"11111111",
  39814=>"00000001",
  39815=>"00000110",
  39816=>"11111100",
  39817=>"11111101",
  39818=>"11111111",
  39819=>"11111111",
  39820=>"11111101",
  39821=>"00000001",
  39822=>"11111111",
  39823=>"00000011",
  39824=>"00000001",
  39825=>"00000100",
  39826=>"00000011",
  39827=>"00000001",
  39828=>"11111111",
  39829=>"00000011",
  39830=>"11111111",
  39831=>"00000001",
  39832=>"11111101",
  39833=>"11111101",
  39834=>"00000110",
  39835=>"11111100",
  39836=>"11111111",
  39837=>"00000000",
  39838=>"11111011",
  39839=>"00000101",
  39840=>"00000100",
  39841=>"11111101",
  39842=>"11111111",
  39843=>"11111110",
  39844=>"00000000",
  39845=>"11111110",
  39846=>"00000010",
  39847=>"00000001",
  39848=>"11111110",
  39849=>"11111101",
  39850=>"00000011",
  39851=>"00000010",
  39852=>"00000010",
  39853=>"11111101",
  39854=>"11111110",
  39855=>"00000000",
  39856=>"11111111",
  39857=>"00000101",
  39858=>"11111100",
  39859=>"00000001",
  39860=>"00000010",
  39861=>"00000010",
  39862=>"00000000",
  39863=>"11111111",
  39864=>"00000000",
  39865=>"11111110",
  39866=>"00000011",
  39867=>"00000100",
  39868=>"11111111",
  39869=>"11111100",
  39870=>"00000001",
  39871=>"00000000",
  39872=>"11111110",
  39873=>"11111010",
  39874=>"00000000",
  39875=>"00000000",
  39876=>"11111110",
  39877=>"00000000",
  39878=>"11111110",
  39879=>"11111111",
  39880=>"00000000",
  39881=>"00000010",
  39882=>"00000100",
  39883=>"00000000",
  39884=>"00000100",
  39885=>"00000101",
  39886=>"00000011",
  39887=>"00000000",
  39888=>"00000011",
  39889=>"11111101",
  39890=>"11111101",
  39891=>"00000000",
  39892=>"00000000",
  39893=>"00000000",
  39894=>"11111100",
  39895=>"11111101",
  39896=>"00000001",
  39897=>"00000011",
  39898=>"00001000",
  39899=>"11111101",
  39900=>"11111110",
  39901=>"00000001",
  39902=>"00000011",
  39903=>"11111101",
  39904=>"00000000",
  39905=>"11111110",
  39906=>"00000011",
  39907=>"00000011",
  39908=>"00000000",
  39909=>"00000011",
  39910=>"11111101",
  39911=>"11111010",
  39912=>"00000010",
  39913=>"00000100",
  39914=>"00000011",
  39915=>"11111111",
  39916=>"00000100",
  39917=>"11111111",
  39918=>"11111101",
  39919=>"00000011",
  39920=>"00000000",
  39921=>"00000001",
  39922=>"11111100",
  39923=>"00000110",
  39924=>"00000001",
  39925=>"11111100",
  39926=>"11111100",
  39927=>"00000000",
  39928=>"11111011",
  39929=>"11111110",
  39930=>"11111111",
  39931=>"11111101",
  39932=>"00000010",
  39933=>"11111110",
  39934=>"00000000",
  39935=>"11111111",
  39936=>"11111110",
  39937=>"11111110",
  39938=>"11111101",
  39939=>"00000010",
  39940=>"11111101",
  39941=>"11111101",
  39942=>"00000100",
  39943=>"00000011",
  39944=>"11111100",
  39945=>"11111110",
  39946=>"11111111",
  39947=>"00000001",
  39948=>"00000000",
  39949=>"11111110",
  39950=>"00000001",
  39951=>"00000000",
  39952=>"00000101",
  39953=>"00000001",
  39954=>"11111101",
  39955=>"11111110",
  39956=>"00000001",
  39957=>"11111110",
  39958=>"00000101",
  39959=>"11111101",
  39960=>"11111110",
  39961=>"11111111",
  39962=>"11111110",
  39963=>"00000011",
  39964=>"00000011",
  39965=>"00000001",
  39966=>"11111110",
  39967=>"00000010",
  39968=>"11111011",
  39969=>"11111111",
  39970=>"00000011",
  39971=>"11111110",
  39972=>"11111111",
  39973=>"00000000",
  39974=>"11111100",
  39975=>"00000001",
  39976=>"00000010",
  39977=>"11111110",
  39978=>"11111111",
  39979=>"00000000",
  39980=>"00000100",
  39981=>"11111101",
  39982=>"00000010",
  39983=>"00000000",
  39984=>"00000001",
  39985=>"00000001",
  39986=>"11111101",
  39987=>"00000000",
  39988=>"11111101",
  39989=>"00000001",
  39990=>"00000001",
  39991=>"11111110",
  39992=>"11111110",
  39993=>"11111111",
  39994=>"11111110",
  39995=>"00000000",
  39996=>"00000010",
  39997=>"00000000",
  39998=>"00000001",
  39999=>"11111101",
  40000=>"00000010",
  40001=>"00000000",
  40002=>"11111110",
  40003=>"00000000",
  40004=>"11111101",
  40005=>"11111111",
  40006=>"11111100",
  40007=>"00000010",
  40008=>"00000011",
  40009=>"00000001",
  40010=>"00000000",
  40011=>"00000001",
  40012=>"00000000",
  40013=>"11111101",
  40014=>"11111111",
  40015=>"11111110",
  40016=>"00000111",
  40017=>"11111111",
  40018=>"00000110",
  40019=>"00000011",
  40020=>"11111111",
  40021=>"00000010",
  40022=>"11111111",
  40023=>"00000000",
  40024=>"00000001",
  40025=>"11111110",
  40026=>"00000000",
  40027=>"00000000",
  40028=>"11111101",
  40029=>"00000001",
  40030=>"00000011",
  40031=>"11111110",
  40032=>"00000001",
  40033=>"00000011",
  40034=>"00000000",
  40035=>"00000001",
  40036=>"11111101",
  40037=>"00000001",
  40038=>"00000100",
  40039=>"11111110",
  40040=>"00000001",
  40041=>"11111110",
  40042=>"00000100",
  40043=>"00000010",
  40044=>"11111111",
  40045=>"11111101",
  40046=>"11111110",
  40047=>"00000000",
  40048=>"00000111",
  40049=>"11111101",
  40050=>"11111111",
  40051=>"11111111",
  40052=>"00000000",
  40053=>"00000001",
  40054=>"00001000",
  40055=>"11111110",
  40056=>"11111101",
  40057=>"11111111",
  40058=>"11111100",
  40059=>"00000001",
  40060=>"00000011",
  40061=>"00000001",
  40062=>"00000001",
  40063=>"00000011",
  40064=>"00000010",
  40065=>"00000000",
  40066=>"00000000",
  40067=>"00000001",
  40068=>"11111110",
  40069=>"11111111",
  40070=>"11111110",
  40071=>"00000000",
  40072=>"00000000",
  40073=>"11111110",
  40074=>"00000000",
  40075=>"11111100",
  40076=>"11111111",
  40077=>"00000010",
  40078=>"11111111",
  40079=>"00000001",
  40080=>"00000011",
  40081=>"00000001",
  40082=>"00000010",
  40083=>"00000001",
  40084=>"00000010",
  40085=>"00000000",
  40086=>"00000100",
  40087=>"00000010",
  40088=>"11111100",
  40089=>"00000100",
  40090=>"00000001",
  40091=>"11111100",
  40092=>"00000000",
  40093=>"11111101",
  40094=>"00000010",
  40095=>"11111101",
  40096=>"00000000",
  40097=>"11111111",
  40098=>"11111100",
  40099=>"00000001",
  40100=>"00000001",
  40101=>"11111111",
  40102=>"00000000",
  40103=>"11111110",
  40104=>"11111111",
  40105=>"11111110",
  40106=>"00000001",
  40107=>"00000010",
  40108=>"00000100",
  40109=>"11111100",
  40110=>"11111101",
  40111=>"00000100",
  40112=>"00000010",
  40113=>"00000001",
  40114=>"11111111",
  40115=>"00000000",
  40116=>"11111111",
  40117=>"11111111",
  40118=>"00000000",
  40119=>"00000010",
  40120=>"00000000",
  40121=>"11111100",
  40122=>"00000011",
  40123=>"00000000",
  40124=>"11111110",
  40125=>"00000000",
  40126=>"11111110",
  40127=>"11111101",
  40128=>"00000010",
  40129=>"11111111",
  40130=>"00000010",
  40131=>"00000011",
  40132=>"00000001",
  40133=>"11111111",
  40134=>"11111100",
  40135=>"11111110",
  40136=>"00000000",
  40137=>"11111111",
  40138=>"11111100",
  40139=>"00000001",
  40140=>"11111111",
  40141=>"11111111",
  40142=>"00000000",
  40143=>"00000000",
  40144=>"11111101",
  40145=>"00000110",
  40146=>"11111110",
  40147=>"00000010",
  40148=>"11111111",
  40149=>"00000010",
  40150=>"11111110",
  40151=>"00000010",
  40152=>"00000001",
  40153=>"11111101",
  40154=>"00000000",
  40155=>"11111111",
  40156=>"11111111",
  40157=>"00000100",
  40158=>"11111111",
  40159=>"11111101",
  40160=>"11111111",
  40161=>"11111101",
  40162=>"11111100",
  40163=>"11111100",
  40164=>"00000001",
  40165=>"11111101",
  40166=>"11111101",
  40167=>"11111111",
  40168=>"00000000",
  40169=>"11111100",
  40170=>"11111110",
  40171=>"11111110",
  40172=>"00000000",
  40173=>"00000001",
  40174=>"00000000",
  40175=>"00000000",
  40176=>"00000100",
  40177=>"00000101",
  40178=>"11111110",
  40179=>"11111101",
  40180=>"00000001",
  40181=>"00000001",
  40182=>"00000001",
  40183=>"00000001",
  40184=>"00000011",
  40185=>"00000000",
  40186=>"00000011",
  40187=>"11111111",
  40188=>"11111111",
  40189=>"00000010",
  40190=>"00000000",
  40191=>"00000000",
  40192=>"11111110",
  40193=>"00000001",
  40194=>"00000100",
  40195=>"00000001",
  40196=>"00000010",
  40197=>"00000001",
  40198=>"00000001",
  40199=>"11111111",
  40200=>"00000010",
  40201=>"00000001",
  40202=>"00000100",
  40203=>"11111111",
  40204=>"00000001",
  40205=>"00000001",
  40206=>"11111101",
  40207=>"00000011",
  40208=>"00000000",
  40209=>"11111110",
  40210=>"00000000",
  40211=>"00000001",
  40212=>"11111101",
  40213=>"00000000",
  40214=>"00000001",
  40215=>"00000010",
  40216=>"11111101",
  40217=>"00000000",
  40218=>"11111110",
  40219=>"00000000",
  40220=>"11111111",
  40221=>"00000010",
  40222=>"11111110",
  40223=>"00000000",
  40224=>"00000001",
  40225=>"00000001",
  40226=>"00000001",
  40227=>"00000000",
  40228=>"11111111",
  40229=>"11111101",
  40230=>"00000011",
  40231=>"00000000",
  40232=>"00000100",
  40233=>"00000001",
  40234=>"11111110",
  40235=>"00000001",
  40236=>"11111110",
  40237=>"00000000",
  40238=>"00000000",
  40239=>"00000010",
  40240=>"00000011",
  40241=>"11111110",
  40242=>"11111101",
  40243=>"11111011",
  40244=>"00000010",
  40245=>"00000101",
  40246=>"00000001",
  40247=>"11111110",
  40248=>"11111110",
  40249=>"11111110",
  40250=>"00000001",
  40251=>"00000101",
  40252=>"11111100",
  40253=>"11111100",
  40254=>"00000000",
  40255=>"00000000",
  40256=>"00000010",
  40257=>"11111111",
  40258=>"11111101",
  40259=>"00000000",
  40260=>"11111111",
  40261=>"11111100",
  40262=>"00000100",
  40263=>"11111111",
  40264=>"00000011",
  40265=>"00000001",
  40266=>"11111100",
  40267=>"00000011",
  40268=>"11111101",
  40269=>"11111110",
  40270=>"00000000",
  40271=>"00000001",
  40272=>"00000100",
  40273=>"00000001",
  40274=>"00000001",
  40275=>"00000000",
  40276=>"00000011",
  40277=>"00000001",
  40278=>"00000100",
  40279=>"11111110",
  40280=>"00000010",
  40281=>"00000001",
  40282=>"11111110",
  40283=>"11111100",
  40284=>"00000001",
  40285=>"00000001",
  40286=>"00000010",
  40287=>"00000011",
  40288=>"11111101",
  40289=>"00000010",
  40290=>"11111111",
  40291=>"11111110",
  40292=>"00000011",
  40293=>"00000001",
  40294=>"00000001",
  40295=>"00000010",
  40296=>"00000000",
  40297=>"00000001",
  40298=>"00000001",
  40299=>"00000011",
  40300=>"11111110",
  40301=>"00000001",
  40302=>"11111110",
  40303=>"00000011",
  40304=>"11111111",
  40305=>"11111101",
  40306=>"00000000",
  40307=>"11111101",
  40308=>"11111100",
  40309=>"11111110",
  40310=>"11111111",
  40311=>"11111110",
  40312=>"11111100",
  40313=>"00000001",
  40314=>"11111100",
  40315=>"00000010",
  40316=>"11111111",
  40317=>"00000011",
  40318=>"00000000",
  40319=>"11111110",
  40320=>"00000011",
  40321=>"00000010",
  40322=>"00000101",
  40323=>"00000000",
  40324=>"00000001",
  40325=>"00000001",
  40326=>"11111111",
  40327=>"11111110",
  40328=>"11111111",
  40329=>"11111111",
  40330=>"00000101",
  40331=>"00000000",
  40332=>"00000011",
  40333=>"11111111",
  40334=>"11111110",
  40335=>"11111101",
  40336=>"00000001",
  40337=>"11111101",
  40338=>"00000001",
  40339=>"00000001",
  40340=>"00000001",
  40341=>"00000001",
  40342=>"00000001",
  40343=>"00000011",
  40344=>"11111101",
  40345=>"00000111",
  40346=>"11111111",
  40347=>"00000010",
  40348=>"00000110",
  40349=>"00000101",
  40350=>"11111110",
  40351=>"00000110",
  40352=>"00000010",
  40353=>"11111110",
  40354=>"00000011",
  40355=>"11111111",
  40356=>"00000011",
  40357=>"11111110",
  40358=>"00000100",
  40359=>"11111110",
  40360=>"11111110",
  40361=>"00000100",
  40362=>"00000001",
  40363=>"11111101",
  40364=>"11111101",
  40365=>"00000001",
  40366=>"11111111",
  40367=>"00000011",
  40368=>"00000000",
  40369=>"00000000",
  40370=>"11111111",
  40371=>"00000010",
  40372=>"00000001",
  40373=>"11111110",
  40374=>"00000000",
  40375=>"00000011",
  40376=>"11111111",
  40377=>"11111101",
  40378=>"11111111",
  40379=>"11111101",
  40380=>"11111110",
  40381=>"00000011",
  40382=>"00000110",
  40383=>"11111101",
  40384=>"11111100",
  40385=>"00000000",
  40386=>"00000010",
  40387=>"11111101",
  40388=>"00000000",
  40389=>"11111111",
  40390=>"00000000",
  40391=>"00000011",
  40392=>"11111110",
  40393=>"11111110",
  40394=>"11111101",
  40395=>"11111111",
  40396=>"00000010",
  40397=>"11111111",
  40398=>"00000000",
  40399=>"11111100",
  40400=>"11111111",
  40401=>"00000001",
  40402=>"11111101",
  40403=>"00000101",
  40404=>"00000000",
  40405=>"00000001",
  40406=>"00000000",
  40407=>"00000000",
  40408=>"11111101",
  40409=>"11111100",
  40410=>"00000000",
  40411=>"11111111",
  40412=>"00000010",
  40413=>"00000010",
  40414=>"11111110",
  40415=>"11111100",
  40416=>"11111101",
  40417=>"00000100",
  40418=>"11111101",
  40419=>"00000000",
  40420=>"00000000",
  40421=>"11111111",
  40422=>"11111110",
  40423=>"00000010",
  40424=>"11111111",
  40425=>"00000000",
  40426=>"00000000",
  40427=>"11111111",
  40428=>"00000010",
  40429=>"00000000",
  40430=>"11111111",
  40431=>"00000000",
  40432=>"00000001",
  40433=>"11111111",
  40434=>"00000001",
  40435=>"11111101",
  40436=>"00000000",
  40437=>"11111110",
  40438=>"00000000",
  40439=>"11111111",
  40440=>"11111110",
  40441=>"11111111",
  40442=>"00000000",
  40443=>"11111110",
  40444=>"11111101",
  40445=>"00000110",
  40446=>"11111111",
  40447=>"00000001",
  40448=>"00000000",
  40449=>"00000001",
  40450=>"00000001",
  40451=>"11111110",
  40452=>"11111101",
  40453=>"11111101",
  40454=>"11111101",
  40455=>"00000001",
  40456=>"00000001",
  40457=>"11111111",
  40458=>"11111110",
  40459=>"00000000",
  40460=>"11111101",
  40461=>"00000000",
  40462=>"00000010",
  40463=>"00000100",
  40464=>"11111110",
  40465=>"00000010",
  40466=>"11111100",
  40467=>"11111111",
  40468=>"11111100",
  40469=>"00000000",
  40470=>"11111110",
  40471=>"00000010",
  40472=>"11111101",
  40473=>"00000100",
  40474=>"00000110",
  40475=>"11111110",
  40476=>"00000000",
  40477=>"11111111",
  40478=>"11111111",
  40479=>"11111110",
  40480=>"11111101",
  40481=>"11111110",
  40482=>"00000100",
  40483=>"11111111",
  40484=>"11111111",
  40485=>"00000001",
  40486=>"11111101",
  40487=>"00000010",
  40488=>"11111110",
  40489=>"11111111",
  40490=>"00000100",
  40491=>"11111111",
  40492=>"11111100",
  40493=>"11111110",
  40494=>"11111110",
  40495=>"11111101",
  40496=>"00000001",
  40497=>"11111111",
  40498=>"11111110",
  40499=>"00000011",
  40500=>"11111110",
  40501=>"11111111",
  40502=>"00000000",
  40503=>"11111110",
  40504=>"11111100",
  40505=>"11111110",
  40506=>"00000001",
  40507=>"00000000",
  40508=>"00000101",
  40509=>"11111101",
  40510=>"11111100",
  40511=>"11111101",
  40512=>"11111111",
  40513=>"00000110",
  40514=>"11111110",
  40515=>"00000011",
  40516=>"11111111",
  40517=>"11111111",
  40518=>"00000001",
  40519=>"00000000",
  40520=>"00000001",
  40521=>"11111111",
  40522=>"11111101",
  40523=>"11111101",
  40524=>"00000000",
  40525=>"11111110",
  40526=>"11111110",
  40527=>"00000000",
  40528=>"00000010",
  40529=>"00000000",
  40530=>"00000001",
  40531=>"11111110",
  40532=>"00000001",
  40533=>"00000000",
  40534=>"00000000",
  40535=>"00000001",
  40536=>"11111100",
  40537=>"11111101",
  40538=>"11111111",
  40539=>"00000011",
  40540=>"00000001",
  40541=>"00000000",
  40542=>"11111101",
  40543=>"00000010",
  40544=>"11111111",
  40545=>"00000000",
  40546=>"00000000",
  40547=>"00000010",
  40548=>"11111110",
  40549=>"11111111",
  40550=>"00000001",
  40551=>"11111110",
  40552=>"00001001",
  40553=>"00000001",
  40554=>"11111110",
  40555=>"00000000",
  40556=>"11111110",
  40557=>"00000011",
  40558=>"00000001",
  40559=>"11111111",
  40560=>"11111101",
  40561=>"11111111",
  40562=>"11111111",
  40563=>"00000000",
  40564=>"11111110",
  40565=>"00000010",
  40566=>"11111111",
  40567=>"11111100",
  40568=>"00000010",
  40569=>"00000011",
  40570=>"11111101",
  40571=>"11111111",
  40572=>"00000000",
  40573=>"11111101",
  40574=>"11111101",
  40575=>"00000001",
  40576=>"00000000",
  40577=>"00000010",
  40578=>"00000000",
  40579=>"00000001",
  40580=>"00000000",
  40581=>"11111110",
  40582=>"11111011",
  40583=>"00000000",
  40584=>"11111110",
  40585=>"11111110",
  40586=>"00000001",
  40587=>"00000000",
  40588=>"00000010",
  40589=>"00000001",
  40590=>"00000010",
  40591=>"00000100",
  40592=>"11111111",
  40593=>"11111101",
  40594=>"00000000",
  40595=>"11111110",
  40596=>"00000100",
  40597=>"11111100",
  40598=>"00000000",
  40599=>"00000001",
  40600=>"00000011",
  40601=>"11111111",
  40602=>"11111101",
  40603=>"11111111",
  40604=>"11111111",
  40605=>"11111110",
  40606=>"11111101",
  40607=>"11111100",
  40608=>"11111110",
  40609=>"00000011",
  40610=>"11111100",
  40611=>"00000000",
  40612=>"11111101",
  40613=>"11111110",
  40614=>"11111011",
  40615=>"11111100",
  40616=>"11111101",
  40617=>"11111101",
  40618=>"00000100",
  40619=>"11111100",
  40620=>"00000010",
  40621=>"00000000",
  40622=>"00000011",
  40623=>"11111110",
  40624=>"00000000",
  40625=>"00000011",
  40626=>"11111111",
  40627=>"00000000",
  40628=>"00000001",
  40629=>"00000001",
  40630=>"11111111",
  40631=>"00000011",
  40632=>"11111110",
  40633=>"00000001",
  40634=>"11111110",
  40635=>"00000001",
  40636=>"00000100",
  40637=>"11111101",
  40638=>"00000100",
  40639=>"11111110",
  40640=>"00000001",
  40641=>"00000010",
  40642=>"00000100",
  40643=>"00000011",
  40644=>"00000100",
  40645=>"11111011",
  40646=>"11111101",
  40647=>"11111110",
  40648=>"11111101",
  40649=>"00000000",
  40650=>"11111110",
  40651=>"00000001",
  40652=>"11111101",
  40653=>"00000001",
  40654=>"11111101",
  40655=>"00000011",
  40656=>"00000001",
  40657=>"11111110",
  40658=>"11111111",
  40659=>"00000001",
  40660=>"11111110",
  40661=>"00000000",
  40662=>"11111110",
  40663=>"11111111",
  40664=>"11111110",
  40665=>"11111110",
  40666=>"11111101",
  40667=>"11111110",
  40668=>"11111110",
  40669=>"00000010",
  40670=>"00000001",
  40671=>"11111110",
  40672=>"00000011",
  40673=>"11111101",
  40674=>"00000000",
  40675=>"00000001",
  40676=>"11111110",
  40677=>"11111111",
  40678=>"11111100",
  40679=>"11111110",
  40680=>"11111111",
  40681=>"00000000",
  40682=>"11111101",
  40683=>"00000000",
  40684=>"00000000",
  40685=>"11111110",
  40686=>"11111111",
  40687=>"00000000",
  40688=>"00000000",
  40689=>"00000100",
  40690=>"11111101",
  40691=>"00000010",
  40692=>"00000100",
  40693=>"11111110",
  40694=>"11111101",
  40695=>"00000100",
  40696=>"00000000",
  40697=>"11111111",
  40698=>"11111110",
  40699=>"11111011",
  40700=>"11111110",
  40701=>"00000010",
  40702=>"00000011",
  40703=>"11111101",
  40704=>"00000001",
  40705=>"00000001",
  40706=>"00000010",
  40707=>"00000001",
  40708=>"11111110",
  40709=>"00000010",
  40710=>"11111110",
  40711=>"11111111",
  40712=>"11111101",
  40713=>"11111111",
  40714=>"11111100",
  40715=>"00000011",
  40716=>"00000110",
  40717=>"11111111",
  40718=>"11111111",
  40719=>"00000001",
  40720=>"11111100",
  40721=>"00000000",
  40722=>"00000000",
  40723=>"00000001",
  40724=>"00000010",
  40725=>"00000001",
  40726=>"00000100",
  40727=>"11111111",
  40728=>"11111110",
  40729=>"00000110",
  40730=>"11111111",
  40731=>"11111101",
  40732=>"00000000",
  40733=>"00000101",
  40734=>"11111110",
  40735=>"11111111",
  40736=>"00000010",
  40737=>"11111101",
  40738=>"00000000",
  40739=>"11111100",
  40740=>"11111110",
  40741=>"11111100",
  40742=>"00000010",
  40743=>"11111111",
  40744=>"00000000",
  40745=>"11111111",
  40746=>"00000000",
  40747=>"00000000",
  40748=>"00000010",
  40749=>"00000011",
  40750=>"11111111",
  40751=>"11111100",
  40752=>"00000000",
  40753=>"11111011",
  40754=>"00000110",
  40755=>"11111110",
  40756=>"00000010",
  40757=>"00000100",
  40758=>"00000000",
  40759=>"11111110",
  40760=>"00000010",
  40761=>"11111101",
  40762=>"11111111",
  40763=>"11111101",
  40764=>"11111101",
  40765=>"00000010",
  40766=>"00000001",
  40767=>"00000001",
  40768=>"11111100",
  40769=>"11111110",
  40770=>"00000010",
  40771=>"11111101",
  40772=>"11111110",
  40773=>"00000000",
  40774=>"00000000",
  40775=>"11111101",
  40776=>"00000100",
  40777=>"11111101",
  40778=>"00000010",
  40779=>"00000100",
  40780=>"11111101",
  40781=>"11111110",
  40782=>"11111101",
  40783=>"00000000",
  40784=>"11111111",
  40785=>"00000011",
  40786=>"00000001",
  40787=>"11111101",
  40788=>"00000000",
  40789=>"00000000",
  40790=>"11111110",
  40791=>"11111110",
  40792=>"00000000",
  40793=>"00000000",
  40794=>"00000000",
  40795=>"00000100",
  40796=>"00000001",
  40797=>"00000001",
  40798=>"11111111",
  40799=>"00000000",
  40800=>"00000001",
  40801=>"00000001",
  40802=>"11111101",
  40803=>"11111110",
  40804=>"00000010",
  40805=>"00000000",
  40806=>"11111110",
  40807=>"00000000",
  40808=>"11111100",
  40809=>"11111101",
  40810=>"00000000",
  40811=>"11111101",
  40812=>"11111110",
  40813=>"00000010",
  40814=>"00000011",
  40815=>"11111111",
  40816=>"11111111",
  40817=>"00000000",
  40818=>"00000000",
  40819=>"11111101",
  40820=>"11111111",
  40821=>"00000110",
  40822=>"00000001",
  40823=>"00000001",
  40824=>"00000000",
  40825=>"00000000",
  40826=>"00000000",
  40827=>"11111101",
  40828=>"00000101",
  40829=>"11111101",
  40830=>"00000100",
  40831=>"00000001",
  40832=>"00000000",
  40833=>"11111101",
  40834=>"11111101",
  40835=>"11111101",
  40836=>"00000010",
  40837=>"11111110",
  40838=>"11111111",
  40839=>"00000101",
  40840=>"00000000",
  40841=>"00000000",
  40842=>"11111110",
  40843=>"00000001",
  40844=>"00000000",
  40845=>"00000100",
  40846=>"00000001",
  40847=>"11111110",
  40848=>"00000000",
  40849=>"11111101",
  40850=>"00000010",
  40851=>"00000010",
  40852=>"00000001",
  40853=>"11111101",
  40854=>"00000010",
  40855=>"00000011",
  40856=>"00000000",
  40857=>"11111111",
  40858=>"00000000",
  40859=>"00000100",
  40860=>"00000001",
  40861=>"00000001",
  40862=>"00000001",
  40863=>"11111110",
  40864=>"11111111",
  40865=>"11111111",
  40866=>"00000001",
  40867=>"00000000",
  40868=>"00000010",
  40869=>"11111101",
  40870=>"11111101",
  40871=>"00000000",
  40872=>"00000010",
  40873=>"11111111",
  40874=>"11111101",
  40875=>"00000000",
  40876=>"11111110",
  40877=>"00000001",
  40878=>"00000001",
  40879=>"00000001",
  40880=>"11111111",
  40881=>"11111100",
  40882=>"00000110",
  40883=>"00000000",
  40884=>"11111111",
  40885=>"00000100",
  40886=>"11111101",
  40887=>"11111101",
  40888=>"11111110",
  40889=>"00000001",
  40890=>"00000010",
  40891=>"11111111",
  40892=>"00000000",
  40893=>"11111110",
  40894=>"00000001",
  40895=>"11111110",
  40896=>"00000011",
  40897=>"00000001",
  40898=>"00000000",
  40899=>"00000001",
  40900=>"00000010",
  40901=>"00000010",
  40902=>"11111100",
  40903=>"00000010",
  40904=>"11111111",
  40905=>"11111101",
  40906=>"11111111",
  40907=>"00000000",
  40908=>"00000001",
  40909=>"11111100",
  40910=>"00000001",
  40911=>"11111111",
  40912=>"11111101",
  40913=>"00000000",
  40914=>"00000011",
  40915=>"00000001",
  40916=>"00000000",
  40917=>"11111100",
  40918=>"00000000",
  40919=>"11111101",
  40920=>"00000001",
  40921=>"11111110",
  40922=>"11111110",
  40923=>"11111101",
  40924=>"00000010",
  40925=>"11111110",
  40926=>"11111110",
  40927=>"00000001",
  40928=>"11111100",
  40929=>"00000010",
  40930=>"11111111",
  40931=>"00000011",
  40932=>"00000001",
  40933=>"11111110",
  40934=>"00000101",
  40935=>"11111110",
  40936=>"00000000",
  40937=>"11111111",
  40938=>"11111100",
  40939=>"11111111",
  40940=>"11111110",
  40941=>"00000011",
  40942=>"00000010",
  40943=>"00000010",
  40944=>"00000000",
  40945=>"00000100",
  40946=>"11111101",
  40947=>"00000010",
  40948=>"00000001",
  40949=>"00000010",
  40950=>"00000000",
  40951=>"11111111",
  40952=>"11111101",
  40953=>"11111111",
  40954=>"00000010",
  40955=>"00000011",
  40956=>"00000000",
  40957=>"11111110",
  40958=>"11111111",
  40959=>"11111111",
  40960=>"11111110",
  40961=>"00000011",
  40962=>"00000001",
  40963=>"11111101",
  40964=>"00000000",
  40965=>"00000000",
  40966=>"11111111",
  40967=>"00000101",
  40968=>"00000010",
  40969=>"11111111",
  40970=>"11111111",
  40971=>"00000010",
  40972=>"11111110",
  40973=>"11111110",
  40974=>"00000011",
  40975=>"11111111",
  40976=>"11111100",
  40977=>"11111111",
  40978=>"11111111",
  40979=>"00000001",
  40980=>"11111111",
  40981=>"00000000",
  40982=>"11111110",
  40983=>"11111111",
  40984=>"00000010",
  40985=>"11111111",
  40986=>"00000001",
  40987=>"00000000",
  40988=>"11111111",
  40989=>"00000100",
  40990=>"00000101",
  40991=>"11111111",
  40992=>"00000001",
  40993=>"00000000",
  40994=>"00000100",
  40995=>"11111101",
  40996=>"00000011",
  40997=>"11111110",
  40998=>"00000001",
  40999=>"00000001",
  41000=>"00000000",
  41001=>"11111110",
  41002=>"00000000",
  41003=>"00001000",
  41004=>"00000001",
  41005=>"11111110",
  41006=>"00000000",
  41007=>"00000000",
  41008=>"00000000",
  41009=>"00000010",
  41010=>"11111111",
  41011=>"00000010",
  41012=>"11111111",
  41013=>"00000010",
  41014=>"11111110",
  41015=>"11111101",
  41016=>"11111110",
  41017=>"11111111",
  41018=>"00000000",
  41019=>"00000001",
  41020=>"11111111",
  41021=>"00000000",
  41022=>"11111111",
  41023=>"11111101",
  41024=>"11111101",
  41025=>"11111110",
  41026=>"11111101",
  41027=>"00000010",
  41028=>"11111110",
  41029=>"11111110",
  41030=>"11111111",
  41031=>"11111100",
  41032=>"00000000",
  41033=>"11111101",
  41034=>"00000101",
  41035=>"00000011",
  41036=>"11111101",
  41037=>"00000000",
  41038=>"00000000",
  41039=>"00000010",
  41040=>"11111110",
  41041=>"00000010",
  41042=>"11111111",
  41043=>"00000010",
  41044=>"00000010",
  41045=>"00000000",
  41046=>"00000100",
  41047=>"11111111",
  41048=>"11111110",
  41049=>"00000000",
  41050=>"00000011",
  41051=>"00000000",
  41052=>"00000011",
  41053=>"11111101",
  41054=>"11111111",
  41055=>"00000101",
  41056=>"11111110",
  41057=>"00000001",
  41058=>"00000001",
  41059=>"00000000",
  41060=>"00000100",
  41061=>"11111110",
  41062=>"00000010",
  41063=>"11111101",
  41064=>"00000000",
  41065=>"11111110",
  41066=>"11111101",
  41067=>"11111111",
  41068=>"00000001",
  41069=>"11111111",
  41070=>"11111110",
  41071=>"11111101",
  41072=>"11111110",
  41073=>"00000001",
  41074=>"00000011",
  41075=>"11111100",
  41076=>"00000001",
  41077=>"00000000",
  41078=>"11111110",
  41079=>"00000001",
  41080=>"00000010",
  41081=>"00000001",
  41082=>"11111101",
  41083=>"00000000",
  41084=>"11111101",
  41085=>"00000001",
  41086=>"00000001",
  41087=>"11111110",
  41088=>"00000000",
  41089=>"11111110",
  41090=>"00000001",
  41091=>"00000001",
  41092=>"00000000",
  41093=>"00000001",
  41094=>"00000000",
  41095=>"11111100",
  41096=>"00000001",
  41097=>"00000000",
  41098=>"00000000",
  41099=>"00000010",
  41100=>"11111100",
  41101=>"00000010",
  41102=>"00000001",
  41103=>"11111111",
  41104=>"00000000",
  41105=>"00000011",
  41106=>"11111111",
  41107=>"11111111",
  41108=>"11111100",
  41109=>"00000001",
  41110=>"00000110",
  41111=>"00000100",
  41112=>"00000010",
  41113=>"11111101",
  41114=>"00000001",
  41115=>"00000010",
  41116=>"00000011",
  41117=>"11111100",
  41118=>"00000010",
  41119=>"00000001",
  41120=>"00000010",
  41121=>"00000011",
  41122=>"00000100",
  41123=>"11111100",
  41124=>"11111110",
  41125=>"00000001",
  41126=>"11111100",
  41127=>"00000001",
  41128=>"11111101",
  41129=>"00000000",
  41130=>"00000001",
  41131=>"11111101",
  41132=>"00000001",
  41133=>"11111101",
  41134=>"00000000",
  41135=>"11111110",
  41136=>"00000001",
  41137=>"11111110",
  41138=>"11111111",
  41139=>"00000011",
  41140=>"00000000",
  41141=>"11111110",
  41142=>"00000000",
  41143=>"11111111",
  41144=>"00000000",
  41145=>"00000000",
  41146=>"00000010",
  41147=>"11111111",
  41148=>"00000001",
  41149=>"00000010",
  41150=>"00000100",
  41151=>"11111011",
  41152=>"00000001",
  41153=>"00000100",
  41154=>"11111101",
  41155=>"00000000",
  41156=>"00000000",
  41157=>"11111101",
  41158=>"00000001",
  41159=>"00000010",
  41160=>"00000001",
  41161=>"00000010",
  41162=>"00000000",
  41163=>"11111101",
  41164=>"11111110",
  41165=>"11111101",
  41166=>"11111110",
  41167=>"00000100",
  41168=>"11111100",
  41169=>"00000001",
  41170=>"00000000",
  41171=>"00000010",
  41172=>"00000100",
  41173=>"11111110",
  41174=>"11111111",
  41175=>"11111110",
  41176=>"00000010",
  41177=>"11111110",
  41178=>"00000010",
  41179=>"11111101",
  41180=>"11111101",
  41181=>"00000010",
  41182=>"11111111",
  41183=>"00000010",
  41184=>"00000000",
  41185=>"11111110",
  41186=>"11111111",
  41187=>"11111111",
  41188=>"11111111",
  41189=>"00000110",
  41190=>"00000000",
  41191=>"00000111",
  41192=>"00000010",
  41193=>"11111110",
  41194=>"11111110",
  41195=>"00000100",
  41196=>"11111111",
  41197=>"11111110",
  41198=>"00000001",
  41199=>"00000001",
  41200=>"00000110",
  41201=>"11111110",
  41202=>"00000001",
  41203=>"00000011",
  41204=>"11111110",
  41205=>"00000010",
  41206=>"11111111",
  41207=>"11111100",
  41208=>"00000001",
  41209=>"00000000",
  41210=>"11111111",
  41211=>"00000010",
  41212=>"11111100",
  41213=>"00000000",
  41214=>"00000001",
  41215=>"00000011",
  41216=>"11111110",
  41217=>"00000011",
  41218=>"11111100",
  41219=>"00000000",
  41220=>"00000001",
  41221=>"00000010",
  41222=>"11111111",
  41223=>"11111111",
  41224=>"11111101",
  41225=>"00000000",
  41226=>"11111110",
  41227=>"11111111",
  41228=>"00000001",
  41229=>"00000100",
  41230=>"11111110",
  41231=>"00000001",
  41232=>"00000111",
  41233=>"00000001",
  41234=>"00000000",
  41235=>"11111110",
  41236=>"11111111",
  41237=>"00000011",
  41238=>"00000000",
  41239=>"00000100",
  41240=>"00000000",
  41241=>"00000010",
  41242=>"00000001",
  41243=>"11111111",
  41244=>"11111110",
  41245=>"11111111",
  41246=>"11111101",
  41247=>"00000000",
  41248=>"11111110",
  41249=>"11111101",
  41250=>"00000010",
  41251=>"00000010",
  41252=>"00000100",
  41253=>"11111101",
  41254=>"11111110",
  41255=>"00000010",
  41256=>"11111111",
  41257=>"00000000",
  41258=>"11111111",
  41259=>"11111110",
  41260=>"00000001",
  41261=>"00000000",
  41262=>"11111100",
  41263=>"11111111",
  41264=>"11111100",
  41265=>"00000001",
  41266=>"00000001",
  41267=>"11111110",
  41268=>"00000100",
  41269=>"11111100",
  41270=>"11111110",
  41271=>"00000001",
  41272=>"00000010",
  41273=>"11111101",
  41274=>"11111101",
  41275=>"11111110",
  41276=>"11111111",
  41277=>"11111110",
  41278=>"11111111",
  41279=>"00000010",
  41280=>"11111111",
  41281=>"11111111",
  41282=>"00000000",
  41283=>"11111101",
  41284=>"00000001",
  41285=>"00000010",
  41286=>"00000101",
  41287=>"11111110",
  41288=>"00000000",
  41289=>"11111110",
  41290=>"00000100",
  41291=>"00000011",
  41292=>"00000101",
  41293=>"00000011",
  41294=>"11111111",
  41295=>"00000010",
  41296=>"00000001",
  41297=>"11111101",
  41298=>"11111100",
  41299=>"00000000",
  41300=>"11111111",
  41301=>"11111101",
  41302=>"11111110",
  41303=>"00000010",
  41304=>"11111110",
  41305=>"11111111",
  41306=>"11111110",
  41307=>"00000010",
  41308=>"00000001",
  41309=>"00000001",
  41310=>"11111110",
  41311=>"00000011",
  41312=>"00000000",
  41313=>"00000010",
  41314=>"11111101",
  41315=>"00000100",
  41316=>"00000000",
  41317=>"00000100",
  41318=>"11111110",
  41319=>"11111110",
  41320=>"11111111",
  41321=>"00000010",
  41322=>"11111111",
  41323=>"11111101",
  41324=>"00000001",
  41325=>"11111111",
  41326=>"00000100",
  41327=>"11111111",
  41328=>"00000001",
  41329=>"00000101",
  41330=>"00000101",
  41331=>"00000011",
  41332=>"11111101",
  41333=>"00000000",
  41334=>"00000001",
  41335=>"11111111",
  41336=>"00000011",
  41337=>"00000010",
  41338=>"00000101",
  41339=>"00000001",
  41340=>"00000011",
  41341=>"11111101",
  41342=>"11111111",
  41343=>"00000100",
  41344=>"11111101",
  41345=>"00000000",
  41346=>"00000000",
  41347=>"00000011",
  41348=>"00000000",
  41349=>"00000010",
  41350=>"00000110",
  41351=>"00000001",
  41352=>"00000001",
  41353=>"11111110",
  41354=>"00000001",
  41355=>"11111110",
  41356=>"00000001",
  41357=>"00000010",
  41358=>"00000011",
  41359=>"00000010",
  41360=>"00000001",
  41361=>"00000011",
  41362=>"11111110",
  41363=>"00000001",
  41364=>"11111110",
  41365=>"11111110",
  41366=>"11111110",
  41367=>"11111101",
  41368=>"00000101",
  41369=>"11111011",
  41370=>"00000001",
  41371=>"00000000",
  41372=>"11111111",
  41373=>"11111101",
  41374=>"11111110",
  41375=>"11111110",
  41376=>"00000000",
  41377=>"00000001",
  41378=>"11111101",
  41379=>"11111011",
  41380=>"11111110",
  41381=>"11111011",
  41382=>"00000001",
  41383=>"11111011",
  41384=>"11111110",
  41385=>"00000000",
  41386=>"00000000",
  41387=>"11111101",
  41388=>"11111111",
  41389=>"11111111",
  41390=>"00000000",
  41391=>"11111110",
  41392=>"11111110",
  41393=>"00000011",
  41394=>"00000101",
  41395=>"00000000",
  41396=>"11111100",
  41397=>"11111101",
  41398=>"00000000",
  41399=>"11111101",
  41400=>"11111101",
  41401=>"11111101",
  41402=>"00000011",
  41403=>"11111111",
  41404=>"11111110",
  41405=>"00000010",
  41406=>"00000001",
  41407=>"00000001",
  41408=>"00000000",
  41409=>"00000011",
  41410=>"00000010",
  41411=>"00000011",
  41412=>"00000011",
  41413=>"11111111",
  41414=>"00000110",
  41415=>"11111110",
  41416=>"11111110",
  41417=>"11111111",
  41418=>"11111100",
  41419=>"00000001",
  41420=>"00000001",
  41421=>"00000001",
  41422=>"00000010",
  41423=>"11111101",
  41424=>"00000000",
  41425=>"00000000",
  41426=>"00000000",
  41427=>"00000101",
  41428=>"00000001",
  41429=>"11111100",
  41430=>"00000100",
  41431=>"00000010",
  41432=>"11111110",
  41433=>"00000000",
  41434=>"11111101",
  41435=>"11111101",
  41436=>"11111110",
  41437=>"00000011",
  41438=>"11111101",
  41439=>"00000100",
  41440=>"00000011",
  41441=>"00000100",
  41442=>"00000000",
  41443=>"00000000",
  41444=>"11111111",
  41445=>"11111111",
  41446=>"00000001",
  41447=>"00000001",
  41448=>"00000010",
  41449=>"00000000",
  41450=>"11111101",
  41451=>"00000000",
  41452=>"11111111",
  41453=>"11111110",
  41454=>"00000001",
  41455=>"11111100",
  41456=>"00000001",
  41457=>"11111101",
  41458=>"00000011",
  41459=>"00000000",
  41460=>"11111111",
  41461=>"00000010",
  41462=>"11111110",
  41463=>"00000000",
  41464=>"11111110",
  41465=>"11111110",
  41466=>"00000011",
  41467=>"00000001",
  41468=>"11111110",
  41469=>"00000011",
  41470=>"00000010",
  41471=>"00000001",
  41472=>"00000001",
  41473=>"00000001",
  41474=>"00000001",
  41475=>"11111100",
  41476=>"11111101",
  41477=>"00000010",
  41478=>"00000000",
  41479=>"00000010",
  41480=>"00000000",
  41481=>"11111011",
  41482=>"00000001",
  41483=>"00000011",
  41484=>"11111101",
  41485=>"00000000",
  41486=>"00000111",
  41487=>"00000001",
  41488=>"00000000",
  41489=>"00000001",
  41490=>"00000000",
  41491=>"00000101",
  41492=>"00000011",
  41493=>"00000001",
  41494=>"00000001",
  41495=>"00000010",
  41496=>"00000010",
  41497=>"11111110",
  41498=>"11111101",
  41499=>"11111101",
  41500=>"11111111",
  41501=>"11111110",
  41502=>"11111101",
  41503=>"00000011",
  41504=>"00000010",
  41505=>"00000000",
  41506=>"00000011",
  41507=>"00000001",
  41508=>"11111101",
  41509=>"00000001",
  41510=>"00000001",
  41511=>"00000100",
  41512=>"00000000",
  41513=>"11111110",
  41514=>"00000001",
  41515=>"00000000",
  41516=>"00000100",
  41517=>"00000010",
  41518=>"00000001",
  41519=>"11111110",
  41520=>"00000011",
  41521=>"00000010",
  41522=>"11111111",
  41523=>"11111101",
  41524=>"00000000",
  41525=>"00000011",
  41526=>"11111101",
  41527=>"11111111",
  41528=>"11111101",
  41529=>"11111110",
  41530=>"00000001",
  41531=>"11111110",
  41532=>"00000000",
  41533=>"00000011",
  41534=>"11111110",
  41535=>"11111110",
  41536=>"11111111",
  41537=>"11111100",
  41538=>"00000100",
  41539=>"00000000",
  41540=>"00000010",
  41541=>"00000001",
  41542=>"00000000",
  41543=>"00000000",
  41544=>"00000011",
  41545=>"11111110",
  41546=>"00000000",
  41547=>"00000000",
  41548=>"11111101",
  41549=>"11111010",
  41550=>"00000001",
  41551=>"00000101",
  41552=>"00000101",
  41553=>"11111100",
  41554=>"11111111",
  41555=>"00000000",
  41556=>"00000001",
  41557=>"11111111",
  41558=>"00000011",
  41559=>"00000010",
  41560=>"00000101",
  41561=>"11111110",
  41562=>"11111111",
  41563=>"11111111",
  41564=>"11111111",
  41565=>"11111110",
  41566=>"00000000",
  41567=>"11111111",
  41568=>"00000000",
  41569=>"11111111",
  41570=>"00000010",
  41571=>"11111101",
  41572=>"11111100",
  41573=>"00000001",
  41574=>"00000001",
  41575=>"11111101",
  41576=>"00000010",
  41577=>"11111101",
  41578=>"00000001",
  41579=>"11111110",
  41580=>"11111101",
  41581=>"00000000",
  41582=>"11111111",
  41583=>"11111100",
  41584=>"11111111",
  41585=>"00000000",
  41586=>"00000010",
  41587=>"11111110",
  41588=>"00000011",
  41589=>"00000000",
  41590=>"00000011",
  41591=>"00000110",
  41592=>"11111101",
  41593=>"00000011",
  41594=>"11111100",
  41595=>"11111110",
  41596=>"11111110",
  41597=>"00000000",
  41598=>"00000010",
  41599=>"00000000",
  41600=>"11111101",
  41601=>"00000010",
  41602=>"00000010",
  41603=>"11111101",
  41604=>"11111101",
  41605=>"00000000",
  41606=>"11111011",
  41607=>"11111101",
  41608=>"00000010",
  41609=>"00000010",
  41610=>"11111101",
  41611=>"00000011",
  41612=>"11111110",
  41613=>"00000000",
  41614=>"11111101",
  41615=>"11111111",
  41616=>"00000110",
  41617=>"00000001",
  41618=>"00000001",
  41619=>"00000011",
  41620=>"11111101",
  41621=>"00000011",
  41622=>"00000000",
  41623=>"11111100",
  41624=>"00000000",
  41625=>"00000010",
  41626=>"00000000",
  41627=>"00000001",
  41628=>"11111110",
  41629=>"11111101",
  41630=>"11111110",
  41631=>"11111101",
  41632=>"00000011",
  41633=>"11111100",
  41634=>"11111101",
  41635=>"00000011",
  41636=>"00000010",
  41637=>"00000000",
  41638=>"11111100",
  41639=>"11111110",
  41640=>"11111110",
  41641=>"11111111",
  41642=>"11111101",
  41643=>"11111110",
  41644=>"00000010",
  41645=>"11111110",
  41646=>"00000010",
  41647=>"00000001",
  41648=>"00000010",
  41649=>"11111110",
  41650=>"00000001",
  41651=>"11111011",
  41652=>"11111101",
  41653=>"11111101",
  41654=>"11111110",
  41655=>"00000010",
  41656=>"00000100",
  41657=>"00000001",
  41658=>"11111111",
  41659=>"11111101",
  41660=>"00000100",
  41661=>"00000010",
  41662=>"11111111",
  41663=>"00000001",
  41664=>"00000001",
  41665=>"00000000",
  41666=>"00000001",
  41667=>"11111101",
  41668=>"00000010",
  41669=>"00000011",
  41670=>"11111111",
  41671=>"11111101",
  41672=>"11111110",
  41673=>"00000100",
  41674=>"00000000",
  41675=>"00000101",
  41676=>"11111100",
  41677=>"11111110",
  41678=>"00000000",
  41679=>"00000011",
  41680=>"00000010",
  41681=>"11111101",
  41682=>"00000100",
  41683=>"00000010",
  41684=>"00000001",
  41685=>"00000001",
  41686=>"00000000",
  41687=>"11111111",
  41688=>"11111101",
  41689=>"00000010",
  41690=>"00000001",
  41691=>"00000100",
  41692=>"11111110",
  41693=>"00000010",
  41694=>"00000010",
  41695=>"00000010",
  41696=>"00000000",
  41697=>"11111101",
  41698=>"11111101",
  41699=>"11111110",
  41700=>"11111101",
  41701=>"00000000",
  41702=>"00000001",
  41703=>"11111110",
  41704=>"00000001",
  41705=>"00000100",
  41706=>"11111110",
  41707=>"00000000",
  41708=>"11111110",
  41709=>"00000011",
  41710=>"00000000",
  41711=>"11111011",
  41712=>"00000000",
  41713=>"00000000",
  41714=>"00000100",
  41715=>"00000011",
  41716=>"00000010",
  41717=>"11111111",
  41718=>"00000000",
  41719=>"00000010",
  41720=>"00000000",
  41721=>"11111101",
  41722=>"00000011",
  41723=>"00000000",
  41724=>"00000011",
  41725=>"11111111",
  41726=>"00000000",
  41727=>"11111111",
  41728=>"00000001",
  41729=>"11111111",
  41730=>"11111111",
  41731=>"00000010",
  41732=>"11111110",
  41733=>"00000010",
  41734=>"00000010",
  41735=>"00000110",
  41736=>"00000010",
  41737=>"11111101",
  41738=>"00000000",
  41739=>"00000011",
  41740=>"11111101",
  41741=>"11111100",
  41742=>"00000100",
  41743=>"11111111",
  41744=>"00000011",
  41745=>"00000010",
  41746=>"00000000",
  41747=>"00000000",
  41748=>"11111111",
  41749=>"00000011",
  41750=>"11111110",
  41751=>"11111111",
  41752=>"11111110",
  41753=>"11111101",
  41754=>"00000010",
  41755=>"11111110",
  41756=>"00000010",
  41757=>"11111110",
  41758=>"11111101",
  41759=>"11111110",
  41760=>"00000001",
  41761=>"00000000",
  41762=>"11111101",
  41763=>"11111100",
  41764=>"00000001",
  41765=>"11111101",
  41766=>"11111111",
  41767=>"00000101",
  41768=>"11111101",
  41769=>"11111110",
  41770=>"00000000",
  41771=>"11111110",
  41772=>"00000000",
  41773=>"11111111",
  41774=>"00000001",
  41775=>"11111101",
  41776=>"11111111",
  41777=>"00000000",
  41778=>"00000000",
  41779=>"00000010",
  41780=>"11111110",
  41781=>"00000011",
  41782=>"00000011",
  41783=>"00000000",
  41784=>"11111100",
  41785=>"00000001",
  41786=>"00000000",
  41787=>"00000000",
  41788=>"00000110",
  41789=>"00000001",
  41790=>"00000010",
  41791=>"00000101",
  41792=>"11111110",
  41793=>"00000110",
  41794=>"00000011",
  41795=>"11111111",
  41796=>"00000111",
  41797=>"00000001",
  41798=>"00000101",
  41799=>"11111110",
  41800=>"00000011",
  41801=>"11111110",
  41802=>"00000000",
  41803=>"11111111",
  41804=>"00000010",
  41805=>"00000000",
  41806=>"00000000",
  41807=>"11111110",
  41808=>"00000001",
  41809=>"00000001",
  41810=>"00000010",
  41811=>"00000101",
  41812=>"00000011",
  41813=>"00000001",
  41814=>"11111110",
  41815=>"00000001",
  41816=>"11111111",
  41817=>"00000000",
  41818=>"11111110",
  41819=>"11111110",
  41820=>"11111110",
  41821=>"00000001",
  41822=>"11111110",
  41823=>"00000010",
  41824=>"00000100",
  41825=>"00000000",
  41826=>"11111100",
  41827=>"00000101",
  41828=>"11111111",
  41829=>"00000101",
  41830=>"11111110",
  41831=>"11111100",
  41832=>"11111101",
  41833=>"00000010",
  41834=>"11111111",
  41835=>"11111100",
  41836=>"11111101",
  41837=>"00000001",
  41838=>"11111110",
  41839=>"00000100",
  41840=>"00000000",
  41841=>"00000011",
  41842=>"11111111",
  41843=>"00000010",
  41844=>"00000000",
  41845=>"00000000",
  41846=>"00000000",
  41847=>"11111110",
  41848=>"11111101",
  41849=>"00000000",
  41850=>"00000000",
  41851=>"11111110",
  41852=>"00000000",
  41853=>"00000011",
  41854=>"11111101",
  41855=>"00000000",
  41856=>"00000000",
  41857=>"00000001",
  41858=>"00000000",
  41859=>"00000010",
  41860=>"11111101",
  41861=>"00000001",
  41862=>"11111100",
  41863=>"11111110",
  41864=>"11111111",
  41865=>"11111111",
  41866=>"00000000",
  41867=>"11111111",
  41868=>"11111100",
  41869=>"11111111",
  41870=>"11111110",
  41871=>"11111111",
  41872=>"11111111",
  41873=>"00000010",
  41874=>"11111101",
  41875=>"11111101",
  41876=>"11111110",
  41877=>"00000011",
  41878=>"11111111",
  41879=>"11111111",
  41880=>"11111110",
  41881=>"00000000",
  41882=>"00000011",
  41883=>"11111101",
  41884=>"11111111",
  41885=>"00000011",
  41886=>"00000000",
  41887=>"00000100",
  41888=>"11111111",
  41889=>"11111111",
  41890=>"00000001",
  41891=>"11111110",
  41892=>"00000010",
  41893=>"00000001",
  41894=>"00000000",
  41895=>"11111101",
  41896=>"11111110",
  41897=>"00000010",
  41898=>"00000001",
  41899=>"11111110",
  41900=>"11111111",
  41901=>"00000001",
  41902=>"11111111",
  41903=>"00000100",
  41904=>"11111110",
  41905=>"00000101",
  41906=>"11111101",
  41907=>"00000000",
  41908=>"00000001",
  41909=>"11111101",
  41910=>"00000100",
  41911=>"11111101",
  41912=>"11111011",
  41913=>"11111111",
  41914=>"00000000",
  41915=>"11111111",
  41916=>"11111110",
  41917=>"00000011",
  41918=>"00000000",
  41919=>"11111111",
  41920=>"11111110",
  41921=>"11111110",
  41922=>"11111111",
  41923=>"00000101",
  41924=>"11111101",
  41925=>"00000010",
  41926=>"11111011",
  41927=>"00000000",
  41928=>"00000001",
  41929=>"00000010",
  41930=>"00000000",
  41931=>"11111100",
  41932=>"00000001",
  41933=>"11111100",
  41934=>"11111101",
  41935=>"00000010",
  41936=>"00000010",
  41937=>"11111101",
  41938=>"11111100",
  41939=>"00000001",
  41940=>"00000000",
  41941=>"00000010",
  41942=>"00000000",
  41943=>"11111111",
  41944=>"11111110",
  41945=>"00000011",
  41946=>"11111111",
  41947=>"11111111",
  41948=>"00000000",
  41949=>"00001000",
  41950=>"00000011",
  41951=>"00000010",
  41952=>"11111101",
  41953=>"11111101",
  41954=>"00000001",
  41955=>"11111111",
  41956=>"11111110",
  41957=>"00000010",
  41958=>"00000010",
  41959=>"00000110",
  41960=>"00000001",
  41961=>"11111111",
  41962=>"00000000",
  41963=>"11111101",
  41964=>"00000001",
  41965=>"11111110",
  41966=>"00000001",
  41967=>"11111101",
  41968=>"11111110",
  41969=>"00000010",
  41970=>"00000000",
  41971=>"00000001",
  41972=>"11111111",
  41973=>"11111101",
  41974=>"11111110",
  41975=>"00000011",
  41976=>"11111100",
  41977=>"11111111",
  41978=>"11111100",
  41979=>"00000000",
  41980=>"11111111",
  41981=>"00000010",
  41982=>"00000000",
  41983=>"00000001",
  41984=>"11111110",
  41985=>"11111111",
  41986=>"00000010",
  41987=>"11111110",
  41988=>"00000000",
  41989=>"00000001",
  41990=>"11111111",
  41991=>"11111100",
  41992=>"00000011",
  41993=>"11111111",
  41994=>"11111111",
  41995=>"11111110",
  41996=>"00000001",
  41997=>"00000011",
  41998=>"11111111",
  41999=>"00000100",
  42000=>"00000000",
  42001=>"11111101",
  42002=>"11111110",
  42003=>"11111101",
  42004=>"00000000",
  42005=>"00000000",
  42006=>"00000010",
  42007=>"11111111",
  42008=>"11111101",
  42009=>"00000100",
  42010=>"11111101",
  42011=>"11111100",
  42012=>"00000001",
  42013=>"00000001",
  42014=>"00000010",
  42015=>"00000010",
  42016=>"11111110",
  42017=>"11111111",
  42018=>"11111100",
  42019=>"00000001",
  42020=>"11111101",
  42021=>"11111110",
  42022=>"00000011",
  42023=>"00000010",
  42024=>"00000000",
  42025=>"00000101",
  42026=>"11111110",
  42027=>"00000010",
  42028=>"00000100",
  42029=>"00000010",
  42030=>"00000001",
  42031=>"11111111",
  42032=>"00000001",
  42033=>"11111110",
  42034=>"00000000",
  42035=>"11111111",
  42036=>"00000001",
  42037=>"00000000",
  42038=>"00000001",
  42039=>"00000000",
  42040=>"11111110",
  42041=>"00000110",
  42042=>"00000010",
  42043=>"11111100",
  42044=>"00000010",
  42045=>"00000000",
  42046=>"00000001",
  42047=>"00000011",
  42048=>"11111101",
  42049=>"00000101",
  42050=>"00000001",
  42051=>"11111101",
  42052=>"11111101",
  42053=>"11111101",
  42054=>"00000100",
  42055=>"11111111",
  42056=>"11111110",
  42057=>"11111110",
  42058=>"00000000",
  42059=>"11111101",
  42060=>"00000010",
  42061=>"11111110",
  42062=>"11111111",
  42063=>"00000001",
  42064=>"11111110",
  42065=>"11111110",
  42066=>"00000110",
  42067=>"11111101",
  42068=>"00000001",
  42069=>"00000011",
  42070=>"00000010",
  42071=>"00000010",
  42072=>"00000000",
  42073=>"00000011",
  42074=>"11111101",
  42075=>"11111111",
  42076=>"11111111",
  42077=>"11111100",
  42078=>"11111110",
  42079=>"11111111",
  42080=>"00000010",
  42081=>"00000011",
  42082=>"00000000",
  42083=>"11111101",
  42084=>"11111100",
  42085=>"11111111",
  42086=>"00000000",
  42087=>"11111110",
  42088=>"11111111",
  42089=>"11111110",
  42090=>"00000011",
  42091=>"11111110",
  42092=>"00000010",
  42093=>"00000000",
  42094=>"00000011",
  42095=>"00000100",
  42096=>"00000010",
  42097=>"00000001",
  42098=>"11111110",
  42099=>"00000000",
  42100=>"00000000",
  42101=>"00000101",
  42102=>"11111110",
  42103=>"11111101",
  42104=>"00000101",
  42105=>"00000000",
  42106=>"11111111",
  42107=>"11111110",
  42108=>"00000010",
  42109=>"00000010",
  42110=>"00000000",
  42111=>"00000000",
  42112=>"00000010",
  42113=>"00000010",
  42114=>"11111111",
  42115=>"00000001",
  42116=>"11111110",
  42117=>"11111110",
  42118=>"00000010",
  42119=>"00000001",
  42120=>"11111110",
  42121=>"11111111",
  42122=>"11111101",
  42123=>"00000011",
  42124=>"11111111",
  42125=>"11111100",
  42126=>"00000011",
  42127=>"00000101",
  42128=>"00000001",
  42129=>"00000110",
  42130=>"00000001",
  42131=>"11111110",
  42132=>"00000011",
  42133=>"00000011",
  42134=>"11111100",
  42135=>"00000001",
  42136=>"11111110",
  42137=>"00000101",
  42138=>"00000100",
  42139=>"11111101",
  42140=>"00000000",
  42141=>"11111110",
  42142=>"00000000",
  42143=>"11111100",
  42144=>"11111100",
  42145=>"11111100",
  42146=>"00000001",
  42147=>"11111111",
  42148=>"11111101",
  42149=>"00000000",
  42150=>"11111111",
  42151=>"00000001",
  42152=>"00000011",
  42153=>"11111110",
  42154=>"00000010",
  42155=>"00000100",
  42156=>"11111111",
  42157=>"11111111",
  42158=>"00000011",
  42159=>"11111101",
  42160=>"11111100",
  42161=>"00000000",
  42162=>"11111111",
  42163=>"11111111",
  42164=>"11111111",
  42165=>"00000001",
  42166=>"00000010",
  42167=>"00000010",
  42168=>"00000010",
  42169=>"11111111",
  42170=>"00000100",
  42171=>"00000011",
  42172=>"00000010",
  42173=>"00000000",
  42174=>"11111101",
  42175=>"00000010",
  42176=>"00000001",
  42177=>"00000010",
  42178=>"11111100",
  42179=>"00000010",
  42180=>"11111111",
  42181=>"11111110",
  42182=>"11111110",
  42183=>"00000001",
  42184=>"00000011",
  42185=>"00000011",
  42186=>"11111111",
  42187=>"00000110",
  42188=>"11111101",
  42189=>"11111111",
  42190=>"11111101",
  42191=>"00000001",
  42192=>"00000011",
  42193=>"00000010",
  42194=>"00000000",
  42195=>"11111110",
  42196=>"11111101",
  42197=>"00000001",
  42198=>"11111110",
  42199=>"00000010",
  42200=>"00000010",
  42201=>"11111110",
  42202=>"11111111",
  42203=>"00000000",
  42204=>"00000001",
  42205=>"00000000",
  42206=>"00000000",
  42207=>"11111110",
  42208=>"11111110",
  42209=>"00000010",
  42210=>"11111101",
  42211=>"00000001",
  42212=>"00000011",
  42213=>"00000000",
  42214=>"11111110",
  42215=>"11111111",
  42216=>"11111110",
  42217=>"00000010",
  42218=>"11111111",
  42219=>"11111111",
  42220=>"00000001",
  42221=>"11111111",
  42222=>"00000010",
  42223=>"00000000",
  42224=>"00000011",
  42225=>"11111110",
  42226=>"00000000",
  42227=>"11111101",
  42228=>"00000010",
  42229=>"00000111",
  42230=>"00000001",
  42231=>"00000010",
  42232=>"11111110",
  42233=>"11111100",
  42234=>"00000010",
  42235=>"00000001",
  42236=>"11111111",
  42237=>"00000100",
  42238=>"00000000",
  42239=>"00000001",
  42240=>"11111111",
  42241=>"00000001",
  42242=>"00000001",
  42243=>"11111101",
  42244=>"00000000",
  42245=>"11111110",
  42246=>"00000011",
  42247=>"00000010",
  42248=>"00000011",
  42249=>"00000001",
  42250=>"11111100",
  42251=>"00000001",
  42252=>"00000000",
  42253=>"11111101",
  42254=>"11111111",
  42255=>"11111100",
  42256=>"00000001",
  42257=>"11111110",
  42258=>"11111110",
  42259=>"11111111",
  42260=>"11111110",
  42261=>"00000010",
  42262=>"11111111",
  42263=>"11111110",
  42264=>"00000010",
  42265=>"00000010",
  42266=>"11111111",
  42267=>"11111111",
  42268=>"00000001",
  42269=>"00000000",
  42270=>"11111101",
  42271=>"11111101",
  42272=>"00000000",
  42273=>"00000000",
  42274=>"11111110",
  42275=>"11111110",
  42276=>"11111110",
  42277=>"00000001",
  42278=>"11111110",
  42279=>"11111100",
  42280=>"00000000",
  42281=>"00000000",
  42282=>"00000010",
  42283=>"00000011",
  42284=>"00000000",
  42285=>"11111110",
  42286=>"11111101",
  42287=>"11111101",
  42288=>"00000000",
  42289=>"00000001",
  42290=>"00000000",
  42291=>"00000110",
  42292=>"11111110",
  42293=>"00000101",
  42294=>"11111110",
  42295=>"11111100",
  42296=>"00000000",
  42297=>"11111111",
  42298=>"00000001",
  42299=>"11111111",
  42300=>"00000110",
  42301=>"00000000",
  42302=>"11111110",
  42303=>"11111111",
  42304=>"11111110",
  42305=>"00000001",
  42306=>"00000001",
  42307=>"11111110",
  42308=>"11111101",
  42309=>"00000010",
  42310=>"11111110",
  42311=>"00000000",
  42312=>"11111111",
  42313=>"11111100",
  42314=>"00000001",
  42315=>"00000001",
  42316=>"00000000",
  42317=>"00000001",
  42318=>"11111110",
  42319=>"00000111",
  42320=>"11111100",
  42321=>"00000000",
  42322=>"00000001",
  42323=>"00000010",
  42324=>"11111111",
  42325=>"00000011",
  42326=>"00000000",
  42327=>"00000111",
  42328=>"00000000",
  42329=>"11111101",
  42330=>"11111110",
  42331=>"00000001",
  42332=>"00000001",
  42333=>"00000000",
  42334=>"00000100",
  42335=>"00000010",
  42336=>"00000001",
  42337=>"00000010",
  42338=>"11111110",
  42339=>"00000100",
  42340=>"11111110",
  42341=>"11111110",
  42342=>"00000000",
  42343=>"00000000",
  42344=>"11111111",
  42345=>"11111101",
  42346=>"11111111",
  42347=>"00000110",
  42348=>"00000001",
  42349=>"11111111",
  42350=>"00000011",
  42351=>"00000001",
  42352=>"00000001",
  42353=>"11111111",
  42354=>"11111110",
  42355=>"11111101",
  42356=>"11111111",
  42357=>"00000001",
  42358=>"11111111",
  42359=>"00000010",
  42360=>"00000011",
  42361=>"00000000",
  42362=>"11111100",
  42363=>"00000000",
  42364=>"00000100",
  42365=>"00000011",
  42366=>"00000001",
  42367=>"00000001",
  42368=>"11111110",
  42369=>"00000010",
  42370=>"00000010",
  42371=>"00000000",
  42372=>"11111110",
  42373=>"11111101",
  42374=>"11111101",
  42375=>"00000001",
  42376=>"11111110",
  42377=>"11111110",
  42378=>"00000000",
  42379=>"11111101",
  42380=>"00000001",
  42381=>"11111101",
  42382=>"00000001",
  42383=>"00000000",
  42384=>"00000000",
  42385=>"11111101",
  42386=>"00000010",
  42387=>"00000010",
  42388=>"00000111",
  42389=>"11111110",
  42390=>"00000001",
  42391=>"00000110",
  42392=>"00000100",
  42393=>"00000010",
  42394=>"00000010",
  42395=>"00000010",
  42396=>"00000001",
  42397=>"00000000",
  42398=>"00000001",
  42399=>"11111101",
  42400=>"11111010",
  42401=>"11111110",
  42402=>"00000000",
  42403=>"11111100",
  42404=>"00000000",
  42405=>"00000010",
  42406=>"00000001",
  42407=>"00000011",
  42408=>"11111100",
  42409=>"00000000",
  42410=>"00000011",
  42411=>"00000011",
  42412=>"11111110",
  42413=>"00000001",
  42414=>"11111101",
  42415=>"00000000",
  42416=>"00000101",
  42417=>"11111101",
  42418=>"00000000",
  42419=>"00000100",
  42420=>"00000000",
  42421=>"11111111",
  42422=>"00000010",
  42423=>"11111101",
  42424=>"11111101",
  42425=>"11111110",
  42426=>"00000001",
  42427=>"11111100",
  42428=>"00000001",
  42429=>"11111110",
  42430=>"00000001",
  42431=>"00000001",
  42432=>"00000001",
  42433=>"00000100",
  42434=>"00000111",
  42435=>"11111110",
  42436=>"00000000",
  42437=>"00000011",
  42438=>"11111101",
  42439=>"00000010",
  42440=>"00000001",
  42441=>"11111101",
  42442=>"11111111",
  42443=>"11111100",
  42444=>"00000011",
  42445=>"00000001",
  42446=>"00000001",
  42447=>"00000000",
  42448=>"00000010",
  42449=>"11111111",
  42450=>"00000001",
  42451=>"11111110",
  42452=>"00000010",
  42453=>"00000000",
  42454=>"00000001",
  42455=>"11111101",
  42456=>"00000001",
  42457=>"00000001",
  42458=>"11111111",
  42459=>"00000010",
  42460=>"00000010",
  42461=>"11111111",
  42462=>"00000000",
  42463=>"00000000",
  42464=>"11111110",
  42465=>"11111111",
  42466=>"00000011",
  42467=>"00000010",
  42468=>"00000010",
  42469=>"00000011",
  42470=>"11111111",
  42471=>"00000010",
  42472=>"00000111",
  42473=>"00000101",
  42474=>"00000011",
  42475=>"00000001",
  42476=>"00000001",
  42477=>"00000001",
  42478=>"11111111",
  42479=>"00000100",
  42480=>"11111101",
  42481=>"11111100",
  42482=>"11111101",
  42483=>"00000010",
  42484=>"11111111",
  42485=>"00000001",
  42486=>"00000011",
  42487=>"11111110",
  42488=>"11111101",
  42489=>"11111011",
  42490=>"00000010",
  42491=>"00000011",
  42492=>"00000000",
  42493=>"11111100",
  42494=>"11111110",
  42495=>"00000010",
  42496=>"00000000",
  42497=>"11111101",
  42498=>"00000100",
  42499=>"00000000",
  42500=>"11111100",
  42501=>"11111110",
  42502=>"11111111",
  42503=>"11111101",
  42504=>"11111111",
  42505=>"11111100",
  42506=>"00000001",
  42507=>"00000011",
  42508=>"00000001",
  42509=>"11111110",
  42510=>"00000000",
  42511=>"00000100",
  42512=>"11111110",
  42513=>"11111111",
  42514=>"00000001",
  42515=>"00000100",
  42516=>"00000000",
  42517=>"00000001",
  42518=>"11111110",
  42519=>"11111110",
  42520=>"00000010",
  42521=>"00000010",
  42522=>"11111110",
  42523=>"11111110",
  42524=>"11111101",
  42525=>"00000000",
  42526=>"11111100",
  42527=>"00000000",
  42528=>"00000010",
  42529=>"00000011",
  42530=>"11111100",
  42531=>"00000010",
  42532=>"11111111",
  42533=>"11111110",
  42534=>"00000010",
  42535=>"00000000",
  42536=>"11111110",
  42537=>"00000000",
  42538=>"00000011",
  42539=>"11111101",
  42540=>"00000100",
  42541=>"11111110",
  42542=>"00000011",
  42543=>"11111110",
  42544=>"00000010",
  42545=>"00000000",
  42546=>"11111101",
  42547=>"00000011",
  42548=>"11111110",
  42549=>"11111011",
  42550=>"00000001",
  42551=>"11111101",
  42552=>"00000100",
  42553=>"00000001",
  42554=>"11111111",
  42555=>"11111101",
  42556=>"00000001",
  42557=>"11111110",
  42558=>"11111111",
  42559=>"11111100",
  42560=>"11111111",
  42561=>"00000000",
  42562=>"00000001",
  42563=>"00000000",
  42564=>"00000100",
  42565=>"00000010",
  42566=>"11111110",
  42567=>"11111110",
  42568=>"11111111",
  42569=>"00000010",
  42570=>"11111110",
  42571=>"11111110",
  42572=>"00000011",
  42573=>"11111101",
  42574=>"00000010",
  42575=>"00000001",
  42576=>"00000010",
  42577=>"00000100",
  42578=>"00000000",
  42579=>"11111110",
  42580=>"00000001",
  42581=>"00000010",
  42582=>"11111110",
  42583=>"00000000",
  42584=>"00000000",
  42585=>"11111110",
  42586=>"00000000",
  42587=>"00000001",
  42588=>"00000011",
  42589=>"11111110",
  42590=>"00000100",
  42591=>"00000010",
  42592=>"00000010",
  42593=>"00000000",
  42594=>"00000000",
  42595=>"00000010",
  42596=>"11111111",
  42597=>"00000001",
  42598=>"00000000",
  42599=>"00000010",
  42600=>"11111101",
  42601=>"00000010",
  42602=>"11111110",
  42603=>"11111101",
  42604=>"11111101",
  42605=>"00000101",
  42606=>"11111111",
  42607=>"00000100",
  42608=>"00000000",
  42609=>"11111111",
  42610=>"00000010",
  42611=>"11111101",
  42612=>"11111111",
  42613=>"11111100",
  42614=>"00000001",
  42615=>"00000110",
  42616=>"11111111",
  42617=>"11111111",
  42618=>"00000000",
  42619=>"11111101",
  42620=>"00000011",
  42621=>"11111110",
  42622=>"00000001",
  42623=>"11111111",
  42624=>"00000011",
  42625=>"11111111",
  42626=>"11111101",
  42627=>"00000000",
  42628=>"11111100",
  42629=>"00000111",
  42630=>"11111110",
  42631=>"11111111",
  42632=>"00000001",
  42633=>"00000000",
  42634=>"00000000",
  42635=>"00000011",
  42636=>"11111111",
  42637=>"11111110",
  42638=>"00000010",
  42639=>"00000110",
  42640=>"00000000",
  42641=>"00000101",
  42642=>"11111110",
  42643=>"00000010",
  42644=>"00000001",
  42645=>"00000101",
  42646=>"00000001",
  42647=>"11111111",
  42648=>"00000001",
  42649=>"11111111",
  42650=>"11111110",
  42651=>"11111101",
  42652=>"11111111",
  42653=>"11111111",
  42654=>"00000101",
  42655=>"11111110",
  42656=>"00000010",
  42657=>"00000010",
  42658=>"00000001",
  42659=>"11111100",
  42660=>"00000001",
  42661=>"11111110",
  42662=>"11111110",
  42663=>"11111111",
  42664=>"00000010",
  42665=>"00000010",
  42666=>"00000001",
  42667=>"00000000",
  42668=>"11111111",
  42669=>"11111111",
  42670=>"00000011",
  42671=>"00000101",
  42672=>"11111101",
  42673=>"11111110",
  42674=>"00000001",
  42675=>"00000100",
  42676=>"11111101",
  42677=>"11111110",
  42678=>"11111101",
  42679=>"11111111",
  42680=>"11111111",
  42681=>"00000001",
  42682=>"00000001",
  42683=>"11111100",
  42684=>"11111101",
  42685=>"11111110",
  42686=>"11111111",
  42687=>"00000010",
  42688=>"00000011",
  42689=>"00000000",
  42690=>"00000010",
  42691=>"00000000",
  42692=>"11111110",
  42693=>"11111111",
  42694=>"00000001",
  42695=>"00000001",
  42696=>"11111110",
  42697=>"11111101",
  42698=>"00000100",
  42699=>"11111111",
  42700=>"11111111",
  42701=>"00000100",
  42702=>"11111111",
  42703=>"11111111",
  42704=>"00000001",
  42705=>"11111100",
  42706=>"11111110",
  42707=>"00000110",
  42708=>"11111111",
  42709=>"00000010",
  42710=>"11111111",
  42711=>"11111100",
  42712=>"00000001",
  42713=>"11111111",
  42714=>"11111110",
  42715=>"11111110",
  42716=>"11111110",
  42717=>"11111111",
  42718=>"11111101",
  42719=>"11111110",
  42720=>"00000010",
  42721=>"11111101",
  42722=>"00000011",
  42723=>"00000001",
  42724=>"00000000",
  42725=>"00000000",
  42726=>"00000000",
  42727=>"00000000",
  42728=>"00000001",
  42729=>"11111110",
  42730=>"11111101",
  42731=>"11111110",
  42732=>"11111110",
  42733=>"00000000",
  42734=>"00000001",
  42735=>"00000100",
  42736=>"11111111",
  42737=>"11111100",
  42738=>"00000011",
  42739=>"00000011",
  42740=>"00000100",
  42741=>"00000000",
  42742=>"00000100",
  42743=>"00000010",
  42744=>"00000101",
  42745=>"00000010",
  42746=>"11111101",
  42747=>"11111100",
  42748=>"00000000",
  42749=>"11111100",
  42750=>"00000000",
  42751=>"00000011",
  42752=>"11111101",
  42753=>"11111111",
  42754=>"00000010",
  42755=>"00000000",
  42756=>"00000010",
  42757=>"11111110",
  42758=>"11111111",
  42759=>"11111111",
  42760=>"11111111",
  42761=>"11111110",
  42762=>"00000011",
  42763=>"00000010",
  42764=>"00000011",
  42765=>"11111110",
  42766=>"11111110",
  42767=>"11111111",
  42768=>"11111101",
  42769=>"11111111",
  42770=>"11111101",
  42771=>"11111011",
  42772=>"00000001",
  42773=>"11111101",
  42774=>"00000000",
  42775=>"00000001",
  42776=>"11111101",
  42777=>"00000101",
  42778=>"00000001",
  42779=>"00000100",
  42780=>"00000110",
  42781=>"00000100",
  42782=>"00000001",
  42783=>"11111101",
  42784=>"00000011",
  42785=>"11111100",
  42786=>"00000001",
  42787=>"00000010",
  42788=>"11111111",
  42789=>"11111100",
  42790=>"11111111",
  42791=>"00000100",
  42792=>"00000001",
  42793=>"00000011",
  42794=>"11111110",
  42795=>"11111101",
  42796=>"11111111",
  42797=>"00000011",
  42798=>"11111111",
  42799=>"00000010",
  42800=>"11111011",
  42801=>"00000001",
  42802=>"00000000",
  42803=>"00000010",
  42804=>"00000001",
  42805=>"00000000",
  42806=>"11111101",
  42807=>"00000011",
  42808=>"00000001",
  42809=>"11111111",
  42810=>"11111111",
  42811=>"11111111",
  42812=>"11111110",
  42813=>"00000100",
  42814=>"00000000",
  42815=>"11111111",
  42816=>"11111101",
  42817=>"11111110",
  42818=>"00000101",
  42819=>"00000001",
  42820=>"11111110",
  42821=>"11111101",
  42822=>"11111101",
  42823=>"00000001",
  42824=>"00000010",
  42825=>"00000010",
  42826=>"00000110",
  42827=>"11111111",
  42828=>"11111110",
  42829=>"00000000",
  42830=>"11111100",
  42831=>"00000000",
  42832=>"11111101",
  42833=>"00000010",
  42834=>"11111100",
  42835=>"11111100",
  42836=>"11111110",
  42837=>"11111101",
  42838=>"00000011",
  42839=>"00000010",
  42840=>"00000000",
  42841=>"11111110",
  42842=>"11111110",
  42843=>"00000011",
  42844=>"00000000",
  42845=>"00000010",
  42846=>"00000011",
  42847=>"11111111",
  42848=>"00000001",
  42849=>"00000011",
  42850=>"00000011",
  42851=>"11111111",
  42852=>"00000001",
  42853=>"11111101",
  42854=>"11111101",
  42855=>"11111110",
  42856=>"00000000",
  42857=>"11111100",
  42858=>"00000010",
  42859=>"00000101",
  42860=>"00000001",
  42861=>"00000101",
  42862=>"11111100",
  42863=>"00000000",
  42864=>"00000010",
  42865=>"11111100",
  42866=>"00000001",
  42867=>"11111011",
  42868=>"11111111",
  42869=>"00000010",
  42870=>"00000000",
  42871=>"00000010",
  42872=>"11111111",
  42873=>"00000001",
  42874=>"00000000",
  42875=>"00000000",
  42876=>"11111101",
  42877=>"11111111",
  42878=>"11111101",
  42879=>"11111110",
  42880=>"11111101",
  42881=>"11111101",
  42882=>"00000001",
  42883=>"00000001",
  42884=>"11111101",
  42885=>"11111111",
  42886=>"11111111",
  42887=>"00000011",
  42888=>"00000000",
  42889=>"11111110",
  42890=>"00000000",
  42891=>"00001000",
  42892=>"11111110",
  42893=>"00000100",
  42894=>"00000001",
  42895=>"00000011",
  42896=>"11111111",
  42897=>"11111111",
  42898=>"00000110",
  42899=>"11111111",
  42900=>"00000100",
  42901=>"00000001",
  42902=>"11111110",
  42903=>"11111101",
  42904=>"11111111",
  42905=>"00000011",
  42906=>"00000001",
  42907=>"00000010",
  42908=>"11111111",
  42909=>"00000010",
  42910=>"00000011",
  42911=>"11111110",
  42912=>"00000010",
  42913=>"11111111",
  42914=>"00000110",
  42915=>"00000010",
  42916=>"00000010",
  42917=>"11111101",
  42918=>"00000011",
  42919=>"00000000",
  42920=>"00000000",
  42921=>"11111111",
  42922=>"11111110",
  42923=>"00000000",
  42924=>"00000010",
  42925=>"00000011",
  42926=>"00000001",
  42927=>"00000000",
  42928=>"11111101",
  42929=>"00000000",
  42930=>"00000011",
  42931=>"11111110",
  42932=>"11111110",
  42933=>"11111101",
  42934=>"11111110",
  42935=>"11111111",
  42936=>"11111100",
  42937=>"11111101",
  42938=>"11111101",
  42939=>"11111110",
  42940=>"00000001",
  42941=>"11111111",
  42942=>"11111111",
  42943=>"11111111",
  42944=>"00000000",
  42945=>"11111110",
  42946=>"11111110",
  42947=>"11111111",
  42948=>"00000010",
  42949=>"11111101",
  42950=>"00000100",
  42951=>"11111111",
  42952=>"00000001",
  42953=>"11111101",
  42954=>"11111101",
  42955=>"00000010",
  42956=>"11111101",
  42957=>"00000010",
  42958=>"11111111",
  42959=>"00000011",
  42960=>"00000000",
  42961=>"11111111",
  42962=>"00000010",
  42963=>"00000000",
  42964=>"00000001",
  42965=>"11111101",
  42966=>"11111101",
  42967=>"00000100",
  42968=>"11111110",
  42969=>"11111111",
  42970=>"00000010",
  42971=>"00000001",
  42972=>"00000000",
  42973=>"11111110",
  42974=>"11111111",
  42975=>"11111100",
  42976=>"00000001",
  42977=>"00000000",
  42978=>"00000000",
  42979=>"00000001",
  42980=>"00000100",
  42981=>"00000000",
  42982=>"11111100",
  42983=>"11111110",
  42984=>"00000000",
  42985=>"11111110",
  42986=>"11111101",
  42987=>"00000111",
  42988=>"11111100",
  42989=>"00000010",
  42990=>"00000000",
  42991=>"00000000",
  42992=>"11111101",
  42993=>"11111110",
  42994=>"11111101",
  42995=>"00000011",
  42996=>"11111111",
  42997=>"11111111",
  42998=>"11111101",
  42999=>"00000000",
  43000=>"11111111",
  43001=>"11111110",
  43002=>"00000010",
  43003=>"11111110",
  43004=>"11111111",
  43005=>"11111101",
  43006=>"11111110",
  43007=>"11111110",
  43008=>"00000011",
  43009=>"00000001",
  43010=>"00000001",
  43011=>"11111111",
  43012=>"11111110",
  43013=>"00000011",
  43014=>"00000011",
  43015=>"11111101",
  43016=>"11111101",
  43017=>"11111101",
  43018=>"11111110",
  43019=>"11111101",
  43020=>"00000010",
  43021=>"00000010",
  43022=>"00000001",
  43023=>"00000100",
  43024=>"11111101",
  43025=>"00000110",
  43026=>"00000001",
  43027=>"11111111",
  43028=>"11111011",
  43029=>"00000001",
  43030=>"00000000",
  43031=>"00000001",
  43032=>"11111101",
  43033=>"00000001",
  43034=>"00000010",
  43035=>"00000001",
  43036=>"00000101",
  43037=>"11111101",
  43038=>"00000010",
  43039=>"00000011",
  43040=>"00000010",
  43041=>"00000011",
  43042=>"11111101",
  43043=>"11111110",
  43044=>"00000000",
  43045=>"11111111",
  43046=>"11111111",
  43047=>"00000001",
  43048=>"00000001",
  43049=>"00000100",
  43050=>"11111101",
  43051=>"11111110",
  43052=>"00000001",
  43053=>"00000010",
  43054=>"11111111",
  43055=>"11111111",
  43056=>"00000001",
  43057=>"00000010",
  43058=>"11111110",
  43059=>"00000000",
  43060=>"00000001",
  43061=>"11111111",
  43062=>"11111111",
  43063=>"00000001",
  43064=>"11111111",
  43065=>"11111100",
  43066=>"11111101",
  43067=>"11111101",
  43068=>"11111110",
  43069=>"11111101",
  43070=>"11111101",
  43071=>"11111101",
  43072=>"00000101",
  43073=>"00000001",
  43074=>"11111111",
  43075=>"11111111",
  43076=>"11111110",
  43077=>"11111110",
  43078=>"11111111",
  43079=>"00000001",
  43080=>"11111101",
  43081=>"00000000",
  43082=>"11111111",
  43083=>"00000001",
  43084=>"00000011",
  43085=>"00000001",
  43086=>"11111110",
  43087=>"00000001",
  43088=>"00000000",
  43089=>"11111111",
  43090=>"11111111",
  43091=>"11111111",
  43092=>"11111100",
  43093=>"00000110",
  43094=>"11111101",
  43095=>"00000000",
  43096=>"11111100",
  43097=>"00000000",
  43098=>"00000010",
  43099=>"11111101",
  43100=>"11111110",
  43101=>"11111011",
  43102=>"11111111",
  43103=>"11111101",
  43104=>"00000001",
  43105=>"00000001",
  43106=>"11111111",
  43107=>"11111100",
  43108=>"11111101",
  43109=>"00000010",
  43110=>"00000010",
  43111=>"11111101",
  43112=>"00000100",
  43113=>"11111101",
  43114=>"00000101",
  43115=>"00000101",
  43116=>"11111011",
  43117=>"11111110",
  43118=>"00000000",
  43119=>"00000001",
  43120=>"00000011",
  43121=>"11111100",
  43122=>"11111100",
  43123=>"00000010",
  43124=>"00000010",
  43125=>"11111101",
  43126=>"00000001",
  43127=>"00000100",
  43128=>"00000001",
  43129=>"11111101",
  43130=>"11111100",
  43131=>"11111100",
  43132=>"11111111",
  43133=>"11111111",
  43134=>"11111111",
  43135=>"11111111",
  43136=>"11111111",
  43137=>"00000011",
  43138=>"11111110",
  43139=>"00000001",
  43140=>"00000010",
  43141=>"11111111",
  43142=>"00000001",
  43143=>"00000011",
  43144=>"11111111",
  43145=>"00000000",
  43146=>"00000000",
  43147=>"00000001",
  43148=>"00000001",
  43149=>"11111110",
  43150=>"11111101",
  43151=>"00000010",
  43152=>"11111111",
  43153=>"11111101",
  43154=>"11111111",
  43155=>"11111111",
  43156=>"11111111",
  43157=>"00000100",
  43158=>"11111110",
  43159=>"00000001",
  43160=>"11111110",
  43161=>"11111110",
  43162=>"00000011",
  43163=>"00000010",
  43164=>"00000001",
  43165=>"11111110",
  43166=>"11111101",
  43167=>"11111110",
  43168=>"11111110",
  43169=>"11111101",
  43170=>"00000000",
  43171=>"11111011",
  43172=>"00000000",
  43173=>"00000000",
  43174=>"00000001",
  43175=>"11111101",
  43176=>"11111100",
  43177=>"00000000",
  43178=>"00000100",
  43179=>"11111100",
  43180=>"00000011",
  43181=>"00000000",
  43182=>"11111111",
  43183=>"11111110",
  43184=>"00000010",
  43185=>"11111111",
  43186=>"11111111",
  43187=>"11111110",
  43188=>"11111110",
  43189=>"00000000",
  43190=>"11111101",
  43191=>"11111111",
  43192=>"11111100",
  43193=>"11111101",
  43194=>"11111101",
  43195=>"00000100",
  43196=>"00000001",
  43197=>"11111110",
  43198=>"11111101",
  43199=>"00000000",
  43200=>"00000010",
  43201=>"00000001",
  43202=>"00000010",
  43203=>"11111100",
  43204=>"11111111",
  43205=>"11111111",
  43206=>"11111101",
  43207=>"00000000",
  43208=>"00000100",
  43209=>"00000100",
  43210=>"11111110",
  43211=>"00000010",
  43212=>"11111111",
  43213=>"11111101",
  43214=>"00000010",
  43215=>"11111111",
  43216=>"00000000",
  43217=>"00000100",
  43218=>"00000000",
  43219=>"00000000",
  43220=>"11111110",
  43221=>"00001001",
  43222=>"11111100",
  43223=>"11111111",
  43224=>"11111110",
  43225=>"11111110",
  43226=>"00000011",
  43227=>"00000000",
  43228=>"11111111",
  43229=>"11111100",
  43230=>"11111111",
  43231=>"00000001",
  43232=>"00000010",
  43233=>"11111100",
  43234=>"11111101",
  43235=>"11111101",
  43236=>"00000000",
  43237=>"11111101",
  43238=>"00000001",
  43239=>"11111111",
  43240=>"00000010",
  43241=>"11111101",
  43242=>"11111110",
  43243=>"11111111",
  43244=>"00000000",
  43245=>"11111101",
  43246=>"00000001",
  43247=>"00000010",
  43248=>"11111111",
  43249=>"00000010",
  43250=>"11111111",
  43251=>"11111111",
  43252=>"00000000",
  43253=>"00000011",
  43254=>"00000010",
  43255=>"00000001",
  43256=>"00000100",
  43257=>"00000001",
  43258=>"11111100",
  43259=>"11111101",
  43260=>"00000010",
  43261=>"11111111",
  43262=>"11111101",
  43263=>"00000000",
  43264=>"00000000",
  43265=>"11111100",
  43266=>"00000110",
  43267=>"11111101",
  43268=>"11111110",
  43269=>"00000000",
  43270=>"00000010",
  43271=>"11111101",
  43272=>"11111101",
  43273=>"00000011",
  43274=>"00000011",
  43275=>"11111111",
  43276=>"11111110",
  43277=>"00000010",
  43278=>"11111111",
  43279=>"00000101",
  43280=>"11111110",
  43281=>"00000001",
  43282=>"11111110",
  43283=>"00000101",
  43284=>"11111111",
  43285=>"11111100",
  43286=>"11111110",
  43287=>"11111101",
  43288=>"11111100",
  43289=>"00000100",
  43290=>"11111111",
  43291=>"00000001",
  43292=>"11111111",
  43293=>"11111111",
  43294=>"00000000",
  43295=>"11111101",
  43296=>"00000001",
  43297=>"11111110",
  43298=>"11111110",
  43299=>"00000011",
  43300=>"11111101",
  43301=>"11111100",
  43302=>"11111110",
  43303=>"11111101",
  43304=>"11111100",
  43305=>"00000011",
  43306=>"00000001",
  43307=>"11111111",
  43308=>"11111111",
  43309=>"11111111",
  43310=>"00000100",
  43311=>"00000011",
  43312=>"11111111",
  43313=>"11111111",
  43314=>"00000001",
  43315=>"00000100",
  43316=>"00000000",
  43317=>"00000000",
  43318=>"11111110",
  43319=>"00000001",
  43320=>"11111101",
  43321=>"00000000",
  43322=>"00000000",
  43323=>"00000001",
  43324=>"11111110",
  43325=>"00000001",
  43326=>"00000000",
  43327=>"00000001",
  43328=>"11111111",
  43329=>"00000101",
  43330=>"00000000",
  43331=>"00000001",
  43332=>"00000010",
  43333=>"00000010",
  43334=>"00000111",
  43335=>"00000100",
  43336=>"00000000",
  43337=>"00000110",
  43338=>"11111101",
  43339=>"11111110",
  43340=>"11111110",
  43341=>"11111110",
  43342=>"11111101",
  43343=>"00000001",
  43344=>"00000001",
  43345=>"00000101",
  43346=>"11111111",
  43347=>"11111100",
  43348=>"11111111",
  43349=>"00000011",
  43350=>"00000010",
  43351=>"00000011",
  43352=>"11111110",
  43353=>"11111101",
  43354=>"11111101",
  43355=>"11111110",
  43356=>"11111101",
  43357=>"00000001",
  43358=>"11111110",
  43359=>"00000001",
  43360=>"00000000",
  43361=>"00000101",
  43362=>"11111101",
  43363=>"11111111",
  43364=>"00000001",
  43365=>"11111101",
  43366=>"00000001",
  43367=>"11111111",
  43368=>"11111100",
  43369=>"00000001",
  43370=>"00000000",
  43371=>"00000000",
  43372=>"00000011",
  43373=>"00000010",
  43374=>"00000011",
  43375=>"00000000",
  43376=>"00000001",
  43377=>"11111111",
  43378=>"11111111",
  43379=>"11111011",
  43380=>"11111111",
  43381=>"11111101",
  43382=>"00000000",
  43383=>"11111111",
  43384=>"11111110",
  43385=>"00000100",
  43386=>"00000010",
  43387=>"00000001",
  43388=>"11111111",
  43389=>"11111101",
  43390=>"11111100",
  43391=>"11111110",
  43392=>"11111101",
  43393=>"11111110",
  43394=>"00000001",
  43395=>"00000000",
  43396=>"11111110",
  43397=>"00000000",
  43398=>"11111110",
  43399=>"00000000",
  43400=>"11111110",
  43401=>"00000010",
  43402=>"00000001",
  43403=>"11111111",
  43404=>"00000010",
  43405=>"00000000",
  43406=>"00000001",
  43407=>"11111111",
  43408=>"11111110",
  43409=>"11111111",
  43410=>"00000011",
  43411=>"11111111",
  43412=>"00000011",
  43413=>"11111110",
  43414=>"00000000",
  43415=>"11111101",
  43416=>"00000011",
  43417=>"00000101",
  43418=>"00000000",
  43419=>"11111101",
  43420=>"00000011",
  43421=>"00000000",
  43422=>"11111110",
  43423=>"00000010",
  43424=>"00000100",
  43425=>"11111110",
  43426=>"11111111",
  43427=>"11111110",
  43428=>"00000010",
  43429=>"00000110",
  43430=>"00000010",
  43431=>"00000010",
  43432=>"00000010",
  43433=>"00000001",
  43434=>"11111101",
  43435=>"00000000",
  43436=>"11111111",
  43437=>"00000011",
  43438=>"00000001",
  43439=>"00000001",
  43440=>"11111111",
  43441=>"11111100",
  43442=>"11111110",
  43443=>"00000010",
  43444=>"11111101",
  43445=>"00000111",
  43446=>"00000010",
  43447=>"11111100",
  43448=>"00000000",
  43449=>"00000000",
  43450=>"00000000",
  43451=>"11111111",
  43452=>"11111110",
  43453=>"00000011",
  43454=>"00000000",
  43455=>"11111110",
  43456=>"11111110",
  43457=>"00000010",
  43458=>"00000010",
  43459=>"00000001",
  43460=>"00000010",
  43461=>"11111110",
  43462=>"00000101",
  43463=>"00000001",
  43464=>"11111101",
  43465=>"00000011",
  43466=>"11111110",
  43467=>"11111111",
  43468=>"00000100",
  43469=>"00000000",
  43470=>"11111110",
  43471=>"11111100",
  43472=>"00000001",
  43473=>"11111111",
  43474=>"00000001",
  43475=>"00000101",
  43476=>"11111111",
  43477=>"00000010",
  43478=>"11111101",
  43479=>"11111101",
  43480=>"00000000",
  43481=>"11111111",
  43482=>"00000000",
  43483=>"00000011",
  43484=>"11111110",
  43485=>"00000001",
  43486=>"00000010",
  43487=>"00000011",
  43488=>"00000000",
  43489=>"11111111",
  43490=>"11111110",
  43491=>"00000000",
  43492=>"00000001",
  43493=>"00000100",
  43494=>"11111110",
  43495=>"00000001",
  43496=>"00000001",
  43497=>"11111111",
  43498=>"11111111",
  43499=>"11111111",
  43500=>"11111111",
  43501=>"00000000",
  43502=>"11111111",
  43503=>"00000110",
  43504=>"00000010",
  43505=>"11111111",
  43506=>"00000010",
  43507=>"11111101",
  43508=>"11111111",
  43509=>"00000001",
  43510=>"11111111",
  43511=>"00000001",
  43512=>"00000000",
  43513=>"00000101",
  43514=>"00000001",
  43515=>"00000010",
  43516=>"00000010",
  43517=>"00000010",
  43518=>"11111111",
  43519=>"00000001",
  43520=>"00000010",
  43521=>"00000000",
  43522=>"11111100",
  43523=>"00000000",
  43524=>"00000010",
  43525=>"00000000",
  43526=>"00000000",
  43527=>"11111110",
  43528=>"00000010",
  43529=>"00000000",
  43530=>"11111101",
  43531=>"11111110",
  43532=>"11111110",
  43533=>"00000001",
  43534=>"11111011",
  43535=>"11111101",
  43536=>"11111101",
  43537=>"00000010",
  43538=>"11111111",
  43539=>"00000010",
  43540=>"00000011",
  43541=>"00000001",
  43542=>"00000001",
  43543=>"00000000",
  43544=>"00000010",
  43545=>"11111011",
  43546=>"00000000",
  43547=>"00000001",
  43548=>"00000000",
  43549=>"00000010",
  43550=>"11111110",
  43551=>"11111111",
  43552=>"00000000",
  43553=>"11111111",
  43554=>"11111101",
  43555=>"11111110",
  43556=>"00000100",
  43557=>"11111111",
  43558=>"00000010",
  43559=>"00000001",
  43560=>"11111110",
  43561=>"00000010",
  43562=>"00000111",
  43563=>"11111110",
  43564=>"11111111",
  43565=>"00000100",
  43566=>"11111110",
  43567=>"11111111",
  43568=>"00000001",
  43569=>"00000010",
  43570=>"11111111",
  43571=>"00000010",
  43572=>"00000010",
  43573=>"00000100",
  43574=>"11111111",
  43575=>"00000000",
  43576=>"00000001",
  43577=>"00000000",
  43578=>"11111111",
  43579=>"11111111",
  43580=>"00000001",
  43581=>"00000011",
  43582=>"00000010",
  43583=>"11111110",
  43584=>"11111110",
  43585=>"00000101",
  43586=>"11111110",
  43587=>"11111100",
  43588=>"00000000",
  43589=>"11111110",
  43590=>"00000001",
  43591=>"11111111",
  43592=>"11111101",
  43593=>"00000100",
  43594=>"00000001",
  43595=>"00000001",
  43596=>"00000000",
  43597=>"11111111",
  43598=>"11111110",
  43599=>"00000001",
  43600=>"11111110",
  43601=>"00000000",
  43602=>"11111111",
  43603=>"11111101",
  43604=>"11111110",
  43605=>"00000001",
  43606=>"00000010",
  43607=>"11111111",
  43608=>"11111110",
  43609=>"11111101",
  43610=>"00000001",
  43611=>"11111101",
  43612=>"00000001",
  43613=>"00000010",
  43614=>"11111101",
  43615=>"00000010",
  43616=>"00000000",
  43617=>"00000000",
  43618=>"00000010",
  43619=>"11111101",
  43620=>"00000010",
  43621=>"00000010",
  43622=>"00000001",
  43623=>"11111100",
  43624=>"11111110",
  43625=>"00000000",
  43626=>"00000000",
  43627=>"11111111",
  43628=>"11111100",
  43629=>"00000110",
  43630=>"11111100",
  43631=>"11111110",
  43632=>"11111110",
  43633=>"11111111",
  43634=>"00000000",
  43635=>"11111011",
  43636=>"11111111",
  43637=>"11111111",
  43638=>"11111110",
  43639=>"00000010",
  43640=>"11111111",
  43641=>"11111101",
  43642=>"00000010",
  43643=>"11111111",
  43644=>"11111101",
  43645=>"11111101",
  43646=>"11111101",
  43647=>"00000000",
  43648=>"00000010",
  43649=>"11111110",
  43650=>"00000101",
  43651=>"00000010",
  43652=>"11111111",
  43653=>"00000001",
  43654=>"00000011",
  43655=>"00000011",
  43656=>"11111101",
  43657=>"00000000",
  43658=>"11111100",
  43659=>"11111100",
  43660=>"11111110",
  43661=>"11111101",
  43662=>"00000000",
  43663=>"00000011",
  43664=>"00000011",
  43665=>"11111110",
  43666=>"00000010",
  43667=>"11111101",
  43668=>"00000010",
  43669=>"11111101",
  43670=>"11111110",
  43671=>"11111100",
  43672=>"00000000",
  43673=>"11111100",
  43674=>"11111111",
  43675=>"11111111",
  43676=>"11111110",
  43677=>"00000001",
  43678=>"11111111",
  43679=>"11111101",
  43680=>"11111100",
  43681=>"11111101",
  43682=>"00000011",
  43683=>"11111100",
  43684=>"00000001",
  43685=>"00000000",
  43686=>"00000011",
  43687=>"00000110",
  43688=>"00000010",
  43689=>"00000001",
  43690=>"11111101",
  43691=>"11111101",
  43692=>"00000011",
  43693=>"00000011",
  43694=>"00000011",
  43695=>"00000010",
  43696=>"11111110",
  43697=>"00000010",
  43698=>"00000001",
  43699=>"00000100",
  43700=>"00000001",
  43701=>"00000010",
  43702=>"11111101",
  43703=>"11111110",
  43704=>"00000001",
  43705=>"00000001",
  43706=>"00000000",
  43707=>"11111101",
  43708=>"11111110",
  43709=>"00000010",
  43710=>"11111100",
  43711=>"11111111",
  43712=>"11111101",
  43713=>"00000011",
  43714=>"00000000",
  43715=>"00000010",
  43716=>"11111110",
  43717=>"11111110",
  43718=>"00000110",
  43719=>"00000001",
  43720=>"00000010",
  43721=>"11111100",
  43722=>"11111111",
  43723=>"00000001",
  43724=>"11111110",
  43725=>"00000000",
  43726=>"11111111",
  43727=>"11111110",
  43728=>"11111101",
  43729=>"11111110",
  43730=>"11111110",
  43731=>"00000011",
  43732=>"11111111",
  43733=>"11111110",
  43734=>"11111101",
  43735=>"00000000",
  43736=>"11111110",
  43737=>"00000011",
  43738=>"11111111",
  43739=>"00000000",
  43740=>"00000101",
  43741=>"00000000",
  43742=>"00000011",
  43743=>"11111100",
  43744=>"00000001",
  43745=>"11111110",
  43746=>"00000010",
  43747=>"11111110",
  43748=>"11111111",
  43749=>"00000011",
  43750=>"00000000",
  43751=>"00000000",
  43752=>"00000000",
  43753=>"00000011",
  43754=>"11111111",
  43755=>"11111111",
  43756=>"11111111",
  43757=>"00000010",
  43758=>"00000001",
  43759=>"11111101",
  43760=>"11111110",
  43761=>"11111100",
  43762=>"11111101",
  43763=>"11111111",
  43764=>"11111111",
  43765=>"00000000",
  43766=>"00000000",
  43767=>"00000000",
  43768=>"11111101",
  43769=>"11111110",
  43770=>"00000010",
  43771=>"00000000",
  43772=>"00000010",
  43773=>"00000101",
  43774=>"00000000",
  43775=>"11111111",
  43776=>"11111101",
  43777=>"11111110",
  43778=>"00000010",
  43779=>"11111111",
  43780=>"00000001",
  43781=>"11111110",
  43782=>"11111100",
  43783=>"11111101",
  43784=>"11111110",
  43785=>"11111111",
  43786=>"00000000",
  43787=>"00000000",
  43788=>"00000000",
  43789=>"11111111",
  43790=>"00000010",
  43791=>"00000001",
  43792=>"00000001",
  43793=>"11111101",
  43794=>"11111101",
  43795=>"11111101",
  43796=>"00000001",
  43797=>"00000100",
  43798=>"00000001",
  43799=>"11111101",
  43800=>"11111110",
  43801=>"00000010",
  43802=>"11111111",
  43803=>"11111101",
  43804=>"11111100",
  43805=>"00000101",
  43806=>"00000010",
  43807=>"11111110",
  43808=>"11111100",
  43809=>"11111111",
  43810=>"00000001",
  43811=>"00000000",
  43812=>"00000001",
  43813=>"11111110",
  43814=>"00000010",
  43815=>"11111110",
  43816=>"00000010",
  43817=>"00000100",
  43818=>"00000001",
  43819=>"11111101",
  43820=>"11111110",
  43821=>"11111111",
  43822=>"00000001",
  43823=>"00000011",
  43824=>"00000100",
  43825=>"11111101",
  43826=>"00000111",
  43827=>"11111111",
  43828=>"11111110",
  43829=>"00000000",
  43830=>"00000000",
  43831=>"11111110",
  43832=>"00000101",
  43833=>"00000010",
  43834=>"11111110",
  43835=>"11111100",
  43836=>"00000011",
  43837=>"11111100",
  43838=>"11111111",
  43839=>"00000010",
  43840=>"00000001",
  43841=>"11111110",
  43842=>"00000000",
  43843=>"00000010",
  43844=>"11111110",
  43845=>"11111111",
  43846=>"11111110",
  43847=>"11111101",
  43848=>"11111100",
  43849=>"11111101",
  43850=>"11111110",
  43851=>"00000000",
  43852=>"00000010",
  43853=>"11111101",
  43854=>"11111110",
  43855=>"00000000",
  43856=>"11111111",
  43857=>"11111111",
  43858=>"11111110",
  43859=>"11111111",
  43860=>"00000001",
  43861=>"00000001",
  43862=>"00000001",
  43863=>"00000000",
  43864=>"00000000",
  43865=>"11111110",
  43866=>"00000000",
  43867=>"00000010",
  43868=>"11111110",
  43869=>"11111101",
  43870=>"11111101",
  43871=>"00000001",
  43872=>"00000000",
  43873=>"00000010",
  43874=>"11111101",
  43875=>"00000011",
  43876=>"11111101",
  43877=>"00000001",
  43878=>"00000010",
  43879=>"11111111",
  43880=>"00000010",
  43881=>"11111101",
  43882=>"00000000",
  43883=>"00000100",
  43884=>"00000000",
  43885=>"11111101",
  43886=>"00000010",
  43887=>"00000001",
  43888=>"11111111",
  43889=>"00000001",
  43890=>"11111101",
  43891=>"11111100",
  43892=>"11111110",
  43893=>"11111111",
  43894=>"00000011",
  43895=>"11111101",
  43896=>"00000011",
  43897=>"00000001",
  43898=>"11111110",
  43899=>"00000000",
  43900=>"00000001",
  43901=>"11111111",
  43902=>"00000011",
  43903=>"11111101",
  43904=>"11111111",
  43905=>"11111110",
  43906=>"00000010",
  43907=>"11111110",
  43908=>"00000000",
  43909=>"00000001",
  43910=>"00000101",
  43911=>"11111110",
  43912=>"11111101",
  43913=>"00000000",
  43914=>"11111110",
  43915=>"11111111",
  43916=>"00000000",
  43917=>"00000010",
  43918=>"00000101",
  43919=>"00000001",
  43920=>"00000000",
  43921=>"11111100",
  43922=>"00000011",
  43923=>"00000001",
  43924=>"00000001",
  43925=>"11111111",
  43926=>"00000010",
  43927=>"00000001",
  43928=>"00000100",
  43929=>"11111111",
  43930=>"11111100",
  43931=>"00000100",
  43932=>"11111101",
  43933=>"00000010",
  43934=>"00000001",
  43935=>"11111101",
  43936=>"11111100",
  43937=>"00000000",
  43938=>"00000001",
  43939=>"00000010",
  43940=>"00000000",
  43941=>"00000010",
  43942=>"00000000",
  43943=>"00000010",
  43944=>"11111101",
  43945=>"11111111",
  43946=>"00000010",
  43947=>"00000001",
  43948=>"11111111",
  43949=>"00000001",
  43950=>"11111110",
  43951=>"11111101",
  43952=>"00000010",
  43953=>"11111101",
  43954=>"00000111",
  43955=>"00000010",
  43956=>"00000001",
  43957=>"00000101",
  43958=>"00000000",
  43959=>"00000000",
  43960=>"00000000",
  43961=>"00000000",
  43962=>"11111110",
  43963=>"11111111",
  43964=>"00000000",
  43965=>"11111101",
  43966=>"00000001",
  43967=>"00000001",
  43968=>"00000101",
  43969=>"00000000",
  43970=>"11111111",
  43971=>"00000000",
  43972=>"11111101",
  43973=>"00000001",
  43974=>"11111110",
  43975=>"11111110",
  43976=>"00000000",
  43977=>"11111100",
  43978=>"00000011",
  43979=>"00000011",
  43980=>"00000001",
  43981=>"11111110",
  43982=>"11111100",
  43983=>"00000010",
  43984=>"11111111",
  43985=>"11111101",
  43986=>"11111111",
  43987=>"11111100",
  43988=>"00000011",
  43989=>"11111100",
  43990=>"00000001",
  43991=>"11111101",
  43992=>"00000001",
  43993=>"00000100",
  43994=>"00000010",
  43995=>"11111110",
  43996=>"11111101",
  43997=>"00000000",
  43998=>"00000010",
  43999=>"00000110",
  44000=>"11111110",
  44001=>"11111111",
  44002=>"11111110",
  44003=>"11111111",
  44004=>"11111110",
  44005=>"00000000",
  44006=>"11111111",
  44007=>"00000001",
  44008=>"11111111",
  44009=>"00000001",
  44010=>"00000001",
  44011=>"11111101",
  44012=>"00000001",
  44013=>"00000001",
  44014=>"11111100",
  44015=>"11111110",
  44016=>"00000001",
  44017=>"00000001",
  44018=>"11111110",
  44019=>"00000000",
  44020=>"00000001",
  44021=>"00000001",
  44022=>"11111100",
  44023=>"00000000",
  44024=>"00000010",
  44025=>"00000011",
  44026=>"00000011",
  44027=>"00000001",
  44028=>"11111111",
  44029=>"00000010",
  44030=>"00000000",
  44031=>"00000010",
  44032=>"11111101",
  44033=>"11111100",
  44034=>"11111111",
  44035=>"11111110",
  44036=>"11111110",
  44037=>"11111101",
  44038=>"00000010",
  44039=>"00000000",
  44040=>"00000010",
  44041=>"00000001",
  44042=>"11111101",
  44043=>"00000001",
  44044=>"11111101",
  44045=>"11111101",
  44046=>"00000011",
  44047=>"00000001",
  44048=>"00000011",
  44049=>"11111101",
  44050=>"00000011",
  44051=>"00000000",
  44052=>"00000001",
  44053=>"11111111",
  44054=>"11111101",
  44055=>"00000001",
  44056=>"11111101",
  44057=>"11111100",
  44058=>"11111111",
  44059=>"00000010",
  44060=>"00000010",
  44061=>"11111111",
  44062=>"00000001",
  44063=>"11111101",
  44064=>"11111110",
  44065=>"00000010",
  44066=>"11111111",
  44067=>"00000001",
  44068=>"00000010",
  44069=>"11111111",
  44070=>"00000000",
  44071=>"00000000",
  44072=>"00000001",
  44073=>"00000010",
  44074=>"00000000",
  44075=>"11111100",
  44076=>"00000000",
  44077=>"11111110",
  44078=>"00000001",
  44079=>"11111111",
  44080=>"11111110",
  44081=>"11111101",
  44082=>"11111110",
  44083=>"11111101",
  44084=>"00000000",
  44085=>"11111101",
  44086=>"00000001",
  44087=>"00000011",
  44088=>"00000000",
  44089=>"00000011",
  44090=>"11111111",
  44091=>"11111101",
  44092=>"00000001",
  44093=>"00000011",
  44094=>"11111110",
  44095=>"11111110",
  44096=>"00000010",
  44097=>"00000010",
  44098=>"11111101",
  44099=>"00000000",
  44100=>"11111111",
  44101=>"00000001",
  44102=>"11111111",
  44103=>"11111101",
  44104=>"11111101",
  44105=>"00000010",
  44106=>"11111101",
  44107=>"00000010",
  44108=>"00000001",
  44109=>"00000010",
  44110=>"11111111",
  44111=>"00000010",
  44112=>"11111100",
  44113=>"00000001",
  44114=>"11111101",
  44115=>"00000000",
  44116=>"00000010",
  44117=>"00000010",
  44118=>"11111111",
  44119=>"11111111",
  44120=>"11111110",
  44121=>"00000101",
  44122=>"00000001",
  44123=>"11111101",
  44124=>"00000111",
  44125=>"11111100",
  44126=>"11111111",
  44127=>"11111111",
  44128=>"00000011",
  44129=>"11111110",
  44130=>"11111101",
  44131=>"11111101",
  44132=>"00000010",
  44133=>"11111111",
  44134=>"11111110",
  44135=>"11111100",
  44136=>"11111101",
  44137=>"00000001",
  44138=>"11111100",
  44139=>"00000101",
  44140=>"00000001",
  44141=>"00000101",
  44142=>"00000001",
  44143=>"00000000",
  44144=>"11111101",
  44145=>"00000010",
  44146=>"11111100",
  44147=>"11111100",
  44148=>"00000001",
  44149=>"11111111",
  44150=>"11111111",
  44151=>"00000101",
  44152=>"11111110",
  44153=>"11111111",
  44154=>"11111011",
  44155=>"00000011",
  44156=>"11111110",
  44157=>"11111111",
  44158=>"11111111",
  44159=>"11111101",
  44160=>"00000000",
  44161=>"11111111",
  44162=>"00000001",
  44163=>"11111110",
  44164=>"00000001",
  44165=>"00000001",
  44166=>"00000000",
  44167=>"11111011",
  44168=>"11111111",
  44169=>"00000000",
  44170=>"00000010",
  44171=>"00000101",
  44172=>"11111101",
  44173=>"00000001",
  44174=>"11111110",
  44175=>"11111100",
  44176=>"00000000",
  44177=>"00000001",
  44178=>"11111110",
  44179=>"11111110",
  44180=>"00000100",
  44181=>"00000000",
  44182=>"11111101",
  44183=>"11111111",
  44184=>"00000101",
  44185=>"11111101",
  44186=>"11111110",
  44187=>"11111101",
  44188=>"11111111",
  44189=>"11111111",
  44190=>"00000000",
  44191=>"11111110",
  44192=>"00000010",
  44193=>"11111101",
  44194=>"11111111",
  44195=>"00000010",
  44196=>"00000010",
  44197=>"11111101",
  44198=>"00000011",
  44199=>"11111111",
  44200=>"00000001",
  44201=>"00000010",
  44202=>"11111101",
  44203=>"00000011",
  44204=>"00000001",
  44205=>"11111111",
  44206=>"00000000",
  44207=>"11111100",
  44208=>"00000100",
  44209=>"11111100",
  44210=>"11111110",
  44211=>"00000001",
  44212=>"00000100",
  44213=>"00000000",
  44214=>"00000011",
  44215=>"00000001",
  44216=>"00000000",
  44217=>"11111100",
  44218=>"00000011",
  44219=>"11111100",
  44220=>"00000000",
  44221=>"00000000",
  44222=>"11111100",
  44223=>"11111110",
  44224=>"11111111",
  44225=>"00000000",
  44226=>"11111111",
  44227=>"00000000",
  44228=>"00000000",
  44229=>"11111011",
  44230=>"00000011",
  44231=>"11111111",
  44232=>"00000010",
  44233=>"00000110",
  44234=>"00000110",
  44235=>"11111110",
  44236=>"00000001",
  44237=>"00000011",
  44238=>"11111110",
  44239=>"11111110",
  44240=>"00000100",
  44241=>"11111111",
  44242=>"11111110",
  44243=>"00000000",
  44244=>"00000010",
  44245=>"11111101",
  44246=>"00000000",
  44247=>"00000001",
  44248=>"11111101",
  44249=>"11111101",
  44250=>"11111111",
  44251=>"00000000",
  44252=>"00000001",
  44253=>"11111111",
  44254=>"00000010",
  44255=>"11111110",
  44256=>"11111110",
  44257=>"11111101",
  44258=>"00000010",
  44259=>"00000001",
  44260=>"11111101",
  44261=>"11111111",
  44262=>"11111101",
  44263=>"11111101",
  44264=>"00000000",
  44265=>"11111100",
  44266=>"00000001",
  44267=>"00000001",
  44268=>"00000010",
  44269=>"00000011",
  44270=>"11111110",
  44271=>"00000001",
  44272=>"11111110",
  44273=>"11111110",
  44274=>"11111111",
  44275=>"11111011",
  44276=>"11111110",
  44277=>"00000001",
  44278=>"00000001",
  44279=>"11111111",
  44280=>"00000011",
  44281=>"11111100",
  44282=>"00000010",
  44283=>"00000000",
  44284=>"00000001",
  44285=>"00000010",
  44286=>"00000000",
  44287=>"00000010",
  44288=>"00000001",
  44289=>"11111110",
  44290=>"00000000",
  44291=>"11111101",
  44292=>"00000001",
  44293=>"00000000",
  44294=>"11111101",
  44295=>"11111110",
  44296=>"00000011",
  44297=>"00000001",
  44298=>"11111111",
  44299=>"00000001",
  44300=>"11111111",
  44301=>"11111110",
  44302=>"00000000",
  44303=>"11111111",
  44304=>"11111111",
  44305=>"00000010",
  44306=>"00000001",
  44307=>"00000100",
  44308=>"11111101",
  44309=>"11111110",
  44310=>"11111101",
  44311=>"11111101",
  44312=>"11111110",
  44313=>"00000100",
  44314=>"00000000",
  44315=>"11111101",
  44316=>"00000011",
  44317=>"11111101",
  44318=>"00000000",
  44319=>"00000001",
  44320=>"00000000",
  44321=>"11111111",
  44322=>"00000001",
  44323=>"11111110",
  44324=>"00000011",
  44325=>"00000110",
  44326=>"11111110",
  44327=>"11111111",
  44328=>"00000001",
  44329=>"00000001",
  44330=>"11111110",
  44331=>"00000011",
  44332=>"00000010",
  44333=>"11111111",
  44334=>"11111111",
  44335=>"11111111",
  44336=>"11111100",
  44337=>"11111101",
  44338=>"11111110",
  44339=>"11111111",
  44340=>"11111110",
  44341=>"00000001",
  44342=>"11111110",
  44343=>"00000010",
  44344=>"00000000",
  44345=>"00000010",
  44346=>"00000010",
  44347=>"11111101",
  44348=>"11111101",
  44349=>"11111111",
  44350=>"00000010",
  44351=>"11111111",
  44352=>"00000010",
  44353=>"00000000",
  44354=>"00000000",
  44355=>"00000010",
  44356=>"00000000",
  44357=>"11111101",
  44358=>"00000000",
  44359=>"00000011",
  44360=>"00000010",
  44361=>"00000100",
  44362=>"11111111",
  44363=>"00000000",
  44364=>"00000000",
  44365=>"11111100",
  44366=>"11111101",
  44367=>"11111111",
  44368=>"11111110",
  44369=>"11111111",
  44370=>"00000100",
  44371=>"11111111",
  44372=>"00000010",
  44373=>"11111101",
  44374=>"11111110",
  44375=>"11111101",
  44376=>"11111111",
  44377=>"11111111",
  44378=>"11111110",
  44379=>"11111100",
  44380=>"00000010",
  44381=>"11111110",
  44382=>"00000010",
  44383=>"00000001",
  44384=>"11111111",
  44385=>"11111110",
  44386=>"00000001",
  44387=>"11111100",
  44388=>"11111110",
  44389=>"11111110",
  44390=>"00000011",
  44391=>"11111110",
  44392=>"11111101",
  44393=>"00000001",
  44394=>"00000001",
  44395=>"00000000",
  44396=>"00000010",
  44397=>"00000011",
  44398=>"11111100",
  44399=>"00000001",
  44400=>"11111111",
  44401=>"00000010",
  44402=>"00000000",
  44403=>"11111101",
  44404=>"11111101",
  44405=>"00000000",
  44406=>"11111111",
  44407=>"11111110",
  44408=>"00000110",
  44409=>"00000100",
  44410=>"11111110",
  44411=>"00000100",
  44412=>"00000001",
  44413=>"00000110",
  44414=>"11111111",
  44415=>"00000001",
  44416=>"11111101",
  44417=>"11111110",
  44418=>"00000000",
  44419=>"11111110",
  44420=>"11111110",
  44421=>"00000011",
  44422=>"11111110",
  44423=>"11111110",
  44424=>"00000000",
  44425=>"11111101",
  44426=>"00000010",
  44427=>"11111100",
  44428=>"11111101",
  44429=>"00000010",
  44430=>"00000001",
  44431=>"00000000",
  44432=>"00000001",
  44433=>"11111111",
  44434=>"00000000",
  44435=>"00000010",
  44436=>"11111100",
  44437=>"11111110",
  44438=>"11111101",
  44439=>"00000100",
  44440=>"00000010",
  44441=>"00000001",
  44442=>"00000001",
  44443=>"00000010",
  44444=>"11111110",
  44445=>"11111110",
  44446=>"11111110",
  44447=>"11111110",
  44448=>"11111111",
  44449=>"00000010",
  44450=>"11111111",
  44451=>"00000001",
  44452=>"00000000",
  44453=>"00000110",
  44454=>"00000001",
  44455=>"00000001",
  44456=>"00000100",
  44457=>"00000000",
  44458=>"00000010",
  44459=>"11111101",
  44460=>"00000000",
  44461=>"00000010",
  44462=>"00000000",
  44463=>"11111111",
  44464=>"11111110",
  44465=>"11111101",
  44466=>"11111111",
  44467=>"11111110",
  44468=>"11111101",
  44469=>"11111111",
  44470=>"11111101",
  44471=>"11111101",
  44472=>"11111101",
  44473=>"00000001",
  44474=>"00000100",
  44475=>"11111110",
  44476=>"00000010",
  44477=>"11111111",
  44478=>"11111110",
  44479=>"00000010",
  44480=>"11111101",
  44481=>"11111110",
  44482=>"11111101",
  44483=>"00000011",
  44484=>"11111110",
  44485=>"11111101",
  44486=>"00000001",
  44487=>"11111101",
  44488=>"00000001",
  44489=>"00000000",
  44490=>"11111101",
  44491=>"00000011",
  44492=>"11111111",
  44493=>"00000000",
  44494=>"11111110",
  44495=>"00000001",
  44496=>"00000000",
  44497=>"00000000",
  44498=>"00000011",
  44499=>"00000100",
  44500=>"11111110",
  44501=>"11111100",
  44502=>"11111011",
  44503=>"11111110",
  44504=>"00000010",
  44505=>"00000010",
  44506=>"00000000",
  44507=>"00000001",
  44508=>"11111110",
  44509=>"11111110",
  44510=>"00000001",
  44511=>"00000001",
  44512=>"11111111",
  44513=>"11111100",
  44514=>"11111110",
  44515=>"00000000",
  44516=>"11111110",
  44517=>"00000100",
  44518=>"00000010",
  44519=>"11111111",
  44520=>"00000010",
  44521=>"11111111",
  44522=>"00000100",
  44523=>"11111101",
  44524=>"11111101",
  44525=>"11111101",
  44526=>"00000001",
  44527=>"00000100",
  44528=>"00000001",
  44529=>"00000100",
  44530=>"00000000",
  44531=>"00000010",
  44532=>"00000001",
  44533=>"11111111",
  44534=>"11111110",
  44535=>"00000010",
  44536=>"00000000",
  44537=>"00000010",
  44538=>"11111110",
  44539=>"00000110",
  44540=>"11111101",
  44541=>"11111011",
  44542=>"11111110",
  44543=>"11111111",
  44544=>"11111101",
  44545=>"00000001",
  44546=>"00000101",
  44547=>"00000000",
  44548=>"00000000",
  44549=>"11111111",
  44550=>"00000000",
  44551=>"11111111",
  44552=>"11111101",
  44553=>"11111111",
  44554=>"11111111",
  44555=>"11111110",
  44556=>"00000010",
  44557=>"11111110",
  44558=>"00000011",
  44559=>"11111101",
  44560=>"00000011",
  44561=>"00000010",
  44562=>"11111110",
  44563=>"00000010",
  44564=>"11111100",
  44565=>"11111111",
  44566=>"11111110",
  44567=>"00000001",
  44568=>"11111111",
  44569=>"11111111",
  44570=>"00000001",
  44571=>"11111111",
  44572=>"00000000",
  44573=>"00000101",
  44574=>"00000001",
  44575=>"00000010",
  44576=>"00000010",
  44577=>"00000011",
  44578=>"11111111",
  44579=>"11111100",
  44580=>"11111111",
  44581=>"00000001",
  44582=>"00000000",
  44583=>"00000011",
  44584=>"11111110",
  44585=>"00000011",
  44586=>"00000010",
  44587=>"00000100",
  44588=>"11111100",
  44589=>"00000000",
  44590=>"11111101",
  44591=>"00000101",
  44592=>"11111110",
  44593=>"11111101",
  44594=>"11111111",
  44595=>"00000001",
  44596=>"00000001",
  44597=>"11111111",
  44598=>"11111111",
  44599=>"00000011",
  44600=>"11111101",
  44601=>"00000011",
  44602=>"11111110",
  44603=>"00000011",
  44604=>"00000011",
  44605=>"11111101",
  44606=>"00000000",
  44607=>"00000001",
  44608=>"00000100",
  44609=>"00000011",
  44610=>"11111111",
  44611=>"11111111",
  44612=>"00000001",
  44613=>"00000010",
  44614=>"00000001",
  44615=>"11111100",
  44616=>"00000010",
  44617=>"00000000",
  44618=>"00000011",
  44619=>"00000100",
  44620=>"11111111",
  44621=>"00000011",
  44622=>"00000011",
  44623=>"11111111",
  44624=>"11111101",
  44625=>"11111111",
  44626=>"11111100",
  44627=>"00000001",
  44628=>"00000110",
  44629=>"00000001",
  44630=>"00000001",
  44631=>"11111110",
  44632=>"11111101",
  44633=>"00000010",
  44634=>"11111101",
  44635=>"11111110",
  44636=>"00000010",
  44637=>"00000011",
  44638=>"00000000",
  44639=>"00000001",
  44640=>"00000000",
  44641=>"11111101",
  44642=>"11111101",
  44643=>"11111111",
  44644=>"11111110",
  44645=>"00000001",
  44646=>"11111110",
  44647=>"00000001",
  44648=>"11111111",
  44649=>"11111101",
  44650=>"00000000",
  44651=>"00000001",
  44652=>"00000110",
  44653=>"11111111",
  44654=>"11111110",
  44655=>"11111110",
  44656=>"00000000",
  44657=>"11111111",
  44658=>"00000010",
  44659=>"11111110",
  44660=>"00000000",
  44661=>"11111110",
  44662=>"00000010",
  44663=>"00000010",
  44664=>"11111101",
  44665=>"00000001",
  44666=>"00000010",
  44667=>"11111101",
  44668=>"11111111",
  44669=>"11111111",
  44670=>"00000011",
  44671=>"00000010",
  44672=>"00000000",
  44673=>"00000010",
  44674=>"11111110",
  44675=>"00000000",
  44676=>"00000010",
  44677=>"11111111",
  44678=>"11111111",
  44679=>"11111101",
  44680=>"00000001",
  44681=>"11111110",
  44682=>"00000011",
  44683=>"11111111",
  44684=>"00000000",
  44685=>"11111101",
  44686=>"00000000",
  44687=>"11111101",
  44688=>"11111110",
  44689=>"11111111",
  44690=>"00000000",
  44691=>"11111110",
  44692=>"00000100",
  44693=>"11111101",
  44694=>"00000011",
  44695=>"00000100",
  44696=>"11111110",
  44697=>"00000001",
  44698=>"11111100",
  44699=>"11111111",
  44700=>"11111111",
  44701=>"00000001",
  44702=>"11111110",
  44703=>"00000110",
  44704=>"00000001",
  44705=>"00000001",
  44706=>"00000001",
  44707=>"11111111",
  44708=>"00000010",
  44709=>"11111100",
  44710=>"00000010",
  44711=>"11111110",
  44712=>"11111110",
  44713=>"11111111",
  44714=>"00000011",
  44715=>"00000010",
  44716=>"00000001",
  44717=>"11111111",
  44718=>"00000011",
  44719=>"00000010",
  44720=>"00000000",
  44721=>"00000000",
  44722=>"11111101",
  44723=>"00000000",
  44724=>"00000010",
  44725=>"00000011",
  44726=>"11111111",
  44727=>"00000000",
  44728=>"00000001",
  44729=>"00000000",
  44730=>"11111111",
  44731=>"11111110",
  44732=>"11111110",
  44733=>"00000000",
  44734=>"11111110",
  44735=>"00000010",
  44736=>"11111110",
  44737=>"00000000",
  44738=>"11111111",
  44739=>"00000100",
  44740=>"00000001",
  44741=>"00000100",
  44742=>"11111110",
  44743=>"11111110",
  44744=>"11111111",
  44745=>"00000001",
  44746=>"11111100",
  44747=>"00000000",
  44748=>"00000001",
  44749=>"11111100",
  44750=>"00000001",
  44751=>"00000011",
  44752=>"00000000",
  44753=>"00000010",
  44754=>"11111110",
  44755=>"11111111",
  44756=>"00000001",
  44757=>"00000010",
  44758=>"11111111",
  44759=>"00000011",
  44760=>"11111111",
  44761=>"00000000",
  44762=>"11111101",
  44763=>"11111111",
  44764=>"00000001",
  44765=>"11111110",
  44766=>"00000000",
  44767=>"00000000",
  44768=>"11111100",
  44769=>"00000001",
  44770=>"11111111",
  44771=>"11111101",
  44772=>"00000011",
  44773=>"00000101",
  44774=>"11111111",
  44775=>"11111101",
  44776=>"00000000",
  44777=>"11111110",
  44778=>"00000011",
  44779=>"00000010",
  44780=>"00000001",
  44781=>"00000000",
  44782=>"00000000",
  44783=>"00000010",
  44784=>"00000000",
  44785=>"00000010",
  44786=>"00000001",
  44787=>"00000000",
  44788=>"00000000",
  44789=>"11111111",
  44790=>"11111110",
  44791=>"00000010",
  44792=>"11111101",
  44793=>"11111111",
  44794=>"11111111",
  44795=>"00000000",
  44796=>"11111111",
  44797=>"00000011",
  44798=>"11111100",
  44799=>"00000001",
  44800=>"00000001",
  44801=>"00000000",
  44802=>"00000011",
  44803=>"00000000",
  44804=>"11111110",
  44805=>"11111111",
  44806=>"11111111",
  44807=>"00000000",
  44808=>"00000000",
  44809=>"11111111",
  44810=>"00000001",
  44811=>"11111111",
  44812=>"11111110",
  44813=>"11111111",
  44814=>"00000010",
  44815=>"00000001",
  44816=>"11111110",
  44817=>"00000000",
  44818=>"11111110",
  44819=>"11111100",
  44820=>"11111101",
  44821=>"00000001",
  44822=>"00000011",
  44823=>"11111101",
  44824=>"00000000",
  44825=>"11111101",
  44826=>"11111110",
  44827=>"11111111",
  44828=>"11111110",
  44829=>"11111110",
  44830=>"11111100",
  44831=>"00000100",
  44832=>"11111100",
  44833=>"00000010",
  44834=>"11111111",
  44835=>"00000000",
  44836=>"11111111",
  44837=>"00000100",
  44838=>"11111101",
  44839=>"11111100",
  44840=>"11111110",
  44841=>"00000000",
  44842=>"00000001",
  44843=>"00000100",
  44844=>"11111101",
  44845=>"11111111",
  44846=>"11111110",
  44847=>"11111111",
  44848=>"11111101",
  44849=>"11111110",
  44850=>"11111110",
  44851=>"11111101",
  44852=>"11111101",
  44853=>"11111101",
  44854=>"11111101",
  44855=>"00000001",
  44856=>"00000001",
  44857=>"00000010",
  44858=>"11111111",
  44859=>"11111110",
  44860=>"00000000",
  44861=>"11111110",
  44862=>"11111101",
  44863=>"11111110",
  44864=>"11111110",
  44865=>"11111110",
  44866=>"00000010",
  44867=>"00000001",
  44868=>"11111101",
  44869=>"00000011",
  44870=>"00000000",
  44871=>"11111111",
  44872=>"11111111",
  44873=>"11111101",
  44874=>"00000100",
  44875=>"00000000",
  44876=>"00000001",
  44877=>"11111101",
  44878=>"00000010",
  44879=>"00000000",
  44880=>"00000001",
  44881=>"11111110",
  44882=>"00000011",
  44883=>"11111111",
  44884=>"00000001",
  44885=>"00000011",
  44886=>"11111111",
  44887=>"11111110",
  44888=>"11111111",
  44889=>"00000010",
  44890=>"11111111",
  44891=>"00000010",
  44892=>"11111101",
  44893=>"11111111",
  44894=>"11111100",
  44895=>"11111111",
  44896=>"00000000",
  44897=>"00000001",
  44898=>"00000010",
  44899=>"00000110",
  44900=>"11111111",
  44901=>"00000001",
  44902=>"00000000",
  44903=>"00000100",
  44904=>"00000010",
  44905=>"11111110",
  44906=>"11111110",
  44907=>"11111101",
  44908=>"00000000",
  44909=>"00000101",
  44910=>"00000010",
  44911=>"00000001",
  44912=>"11111110",
  44913=>"00000000",
  44914=>"11111111",
  44915=>"00000001",
  44916=>"11111111",
  44917=>"00000010",
  44918=>"00000101",
  44919=>"00000001",
  44920=>"00000010",
  44921=>"00000000",
  44922=>"00000000",
  44923=>"00000011",
  44924=>"00000000",
  44925=>"00000001",
  44926=>"00000010",
  44927=>"00000000",
  44928=>"11111110",
  44929=>"00000011",
  44930=>"00000000",
  44931=>"00000000",
  44932=>"11111110",
  44933=>"00000010",
  44934=>"11111110",
  44935=>"11111100",
  44936=>"11111110",
  44937=>"11111111",
  44938=>"11111110",
  44939=>"11111111",
  44940=>"00000000",
  44941=>"11111101",
  44942=>"11111111",
  44943=>"00000000",
  44944=>"00000000",
  44945=>"11111100",
  44946=>"11111110",
  44947=>"00000010",
  44948=>"00000001",
  44949=>"11111110",
  44950=>"11111111",
  44951=>"00000001",
  44952=>"00000011",
  44953=>"00000011",
  44954=>"11111110",
  44955=>"11111111",
  44956=>"00000000",
  44957=>"11111110",
  44958=>"00000010",
  44959=>"00000010",
  44960=>"11111110",
  44961=>"11111101",
  44962=>"11111101",
  44963=>"00000000",
  44964=>"00000010",
  44965=>"00000001",
  44966=>"00000000",
  44967=>"11111101",
  44968=>"11111110",
  44969=>"00000010",
  44970=>"00000001",
  44971=>"00000001",
  44972=>"11111101",
  44973=>"11111101",
  44974=>"11111110",
  44975=>"00000010",
  44976=>"11111110",
  44977=>"00000011",
  44978=>"11111111",
  44979=>"11111101",
  44980=>"11111101",
  44981=>"00000010",
  44982=>"00000000",
  44983=>"00000010",
  44984=>"00000011",
  44985=>"00000011",
  44986=>"11111101",
  44987=>"11111111",
  44988=>"11111101",
  44989=>"00000100",
  44990=>"11111110",
  44991=>"11111111",
  44992=>"00000001",
  44993=>"00000001",
  44994=>"00000100",
  44995=>"00000010",
  44996=>"11111110",
  44997=>"00000000",
  44998=>"00001000",
  44999=>"11111111",
  45000=>"00000000",
  45001=>"00000000",
  45002=>"00000011",
  45003=>"00000001",
  45004=>"00000101",
  45005=>"11111110",
  45006=>"11111110",
  45007=>"00000011",
  45008=>"00000010",
  45009=>"00000001",
  45010=>"11111011",
  45011=>"00000010",
  45012=>"00000000",
  45013=>"00000100",
  45014=>"00000001",
  45015=>"00000000",
  45016=>"00000001",
  45017=>"00000101",
  45018=>"00000001",
  45019=>"11111101",
  45020=>"00000011",
  45021=>"11111100",
  45022=>"11111110",
  45023=>"11111110",
  45024=>"00000000",
  45025=>"11111110",
  45026=>"11111101",
  45027=>"00000010",
  45028=>"00000001",
  45029=>"11111101",
  45030=>"11111101",
  45031=>"11111110",
  45032=>"00000001",
  45033=>"11111101",
  45034=>"00001000",
  45035=>"11111110",
  45036=>"00000000",
  45037=>"11111101",
  45038=>"11111101",
  45039=>"11111110",
  45040=>"00000100",
  45041=>"11111110",
  45042=>"00000001",
  45043=>"11111111",
  45044=>"11111101",
  45045=>"00000001",
  45046=>"00000101",
  45047=>"00000101",
  45048=>"00000000",
  45049=>"00000011",
  45050=>"00000100",
  45051=>"11111101",
  45052=>"11111101",
  45053=>"11111110",
  45054=>"00000000",
  45055=>"00000000",
  45056=>"00000001",
  45057=>"00000000",
  45058=>"00000000",
  45059=>"11111111",
  45060=>"00000100",
  45061=>"00000011",
  45062=>"00000001",
  45063=>"11111111",
  45064=>"00000100",
  45065=>"00000001",
  45066=>"00000001",
  45067=>"00000001",
  45068=>"00000000",
  45069=>"00000110",
  45070=>"11111010",
  45071=>"11111111",
  45072=>"11111110",
  45073=>"00000001",
  45074=>"00000100",
  45075=>"11111110",
  45076=>"00000000",
  45077=>"00000010",
  45078=>"11111001",
  45079=>"00000011",
  45080=>"00000100",
  45081=>"00000100",
  45082=>"00000111",
  45083=>"00000111",
  45084=>"11111100",
  45085=>"00000010",
  45086=>"11111111",
  45087=>"00000001",
  45088=>"11111101",
  45089=>"00000111",
  45090=>"00000100",
  45091=>"00000110",
  45092=>"00000000",
  45093=>"00000000",
  45094=>"11111101",
  45095=>"11111101",
  45096=>"00000010",
  45097=>"00000101",
  45098=>"11111101",
  45099=>"00000011",
  45100=>"00000101",
  45101=>"11111101",
  45102=>"00000010",
  45103=>"11111101",
  45104=>"00000000",
  45105=>"11111111",
  45106=>"00000000",
  45107=>"00000010",
  45108=>"00000000",
  45109=>"11111111",
  45110=>"00000010",
  45111=>"11111100",
  45112=>"11111110",
  45113=>"00000100",
  45114=>"00000111",
  45115=>"00000001",
  45116=>"11111110",
  45117=>"11111111",
  45118=>"00000101",
  45119=>"11111110",
  45120=>"00000010",
  45121=>"00000010",
  45122=>"11111110",
  45123=>"11111100",
  45124=>"11111111",
  45125=>"00000000",
  45126=>"11111111",
  45127=>"11111100",
  45128=>"11111110",
  45129=>"00000001",
  45130=>"00000010",
  45131=>"11111101",
  45132=>"11111111",
  45133=>"00000000",
  45134=>"11111110",
  45135=>"11111101",
  45136=>"11111111",
  45137=>"11111111",
  45138=>"00000100",
  45139=>"00000001",
  45140=>"00000000",
  45141=>"11111101",
  45142=>"00000010",
  45143=>"11111101",
  45144=>"11111101",
  45145=>"00000010",
  45146=>"00000000",
  45147=>"11111110",
  45148=>"00000000",
  45149=>"11111111",
  45150=>"11111110",
  45151=>"00000010",
  45152=>"11111101",
  45153=>"00000011",
  45154=>"00000011",
  45155=>"11111111",
  45156=>"11111011",
  45157=>"00000011",
  45158=>"00000101",
  45159=>"00000011",
  45160=>"11111100",
  45161=>"00000011",
  45162=>"11111111",
  45163=>"00000110",
  45164=>"11111111",
  45165=>"00000001",
  45166=>"00000100",
  45167=>"11111110",
  45168=>"11111111",
  45169=>"00000001",
  45170=>"00000100",
  45171=>"00000000",
  45172=>"11111101",
  45173=>"00000011",
  45174=>"00000000",
  45175=>"00000001",
  45176=>"00000000",
  45177=>"00000101",
  45178=>"00000111",
  45179=>"00000100",
  45180=>"11111101",
  45181=>"00000011",
  45182=>"00000001",
  45183=>"00000101",
  45184=>"11111110",
  45185=>"00000001",
  45186=>"11111111",
  45187=>"00000000",
  45188=>"11111111",
  45189=>"00000000",
  45190=>"11111111",
  45191=>"00000100",
  45192=>"00000101",
  45193=>"00000001",
  45194=>"00000000",
  45195=>"00000100",
  45196=>"11111101",
  45197=>"11111011",
  45198=>"00000011",
  45199=>"00000100",
  45200=>"00000100",
  45201=>"00000110",
  45202=>"00000000",
  45203=>"11111110",
  45204=>"00000100",
  45205=>"00000101",
  45206=>"00000011",
  45207=>"11111111",
  45208=>"00000100",
  45209=>"00000000",
  45210=>"11111101",
  45211=>"11111111",
  45212=>"11111101",
  45213=>"00000110",
  45214=>"00000010",
  45215=>"11111110",
  45216=>"00000000",
  45217=>"11111101",
  45218=>"11111110",
  45219=>"00000110",
  45220=>"11111100",
  45221=>"00000010",
  45222=>"11111110",
  45223=>"00000010",
  45224=>"11111110",
  45225=>"00000101",
  45226=>"11111011",
  45227=>"00000100",
  45228=>"11111110",
  45229=>"00000000",
  45230=>"00000011",
  45231=>"00000101",
  45232=>"11111111",
  45233=>"00000101",
  45234=>"11111101",
  45235=>"11111010",
  45236=>"00000101",
  45237=>"00000101",
  45238=>"00000000",
  45239=>"00000010",
  45240=>"11111111",
  45241=>"00000110",
  45242=>"00000011",
  45243=>"00000001",
  45244=>"00000110",
  45245=>"00000010",
  45246=>"00000001",
  45247=>"11111101",
  45248=>"00000010",
  45249=>"11111100",
  45250=>"11111110",
  45251=>"00000100",
  45252=>"00000101",
  45253=>"00000000",
  45254=>"00000010",
  45255=>"00000000",
  45256=>"11111111",
  45257=>"00000100",
  45258=>"11111110",
  45259=>"00000000",
  45260=>"11111101",
  45261=>"00000000",
  45262=>"11111111",
  45263=>"00000000",
  45264=>"00000001",
  45265=>"00000001",
  45266=>"00000001",
  45267=>"11111111",
  45268=>"11111111",
  45269=>"00000000",
  45270=>"11111101",
  45271=>"00000011",
  45272=>"11111101",
  45273=>"11111111",
  45274=>"11111110",
  45275=>"00000101",
  45276=>"11111101",
  45277=>"00000100",
  45278=>"11111111",
  45279=>"00000110",
  45280=>"00000011",
  45281=>"11111111",
  45282=>"00000010",
  45283=>"00000010",
  45284=>"00000001",
  45285=>"11111110",
  45286=>"11111111",
  45287=>"11111101",
  45288=>"11111110",
  45289=>"00000010",
  45290=>"00000001",
  45291=>"00000000",
  45292=>"11111110",
  45293=>"00000011",
  45294=>"11111100",
  45295=>"00000010",
  45296=>"00000000",
  45297=>"00000011",
  45298=>"11111110",
  45299=>"00000000",
  45300=>"00000011",
  45301=>"00000011",
  45302=>"00000000",
  45303=>"11111101",
  45304=>"00000001",
  45305=>"11111111",
  45306=>"11111101",
  45307=>"00000001",
  45308=>"11111110",
  45309=>"00000001",
  45310=>"00000010",
  45311=>"11111011",
  45312=>"00000001",
  45313=>"00000010",
  45314=>"11111011",
  45315=>"11111101",
  45316=>"00000011",
  45317=>"00000000",
  45318=>"00000001",
  45319=>"11111111",
  45320=>"11111100",
  45321=>"00000110",
  45322=>"00000101",
  45323=>"11111111",
  45324=>"00000001",
  45325=>"11111100",
  45326=>"11111101",
  45327=>"00000111",
  45328=>"00000011",
  45329=>"00000010",
  45330=>"11111111",
  45331=>"00000000",
  45332=>"00000010",
  45333=>"00000011",
  45334=>"00000100",
  45335=>"00000000",
  45336=>"11111100",
  45337=>"00000011",
  45338=>"11111111",
  45339=>"11111111",
  45340=>"00000000",
  45341=>"11111011",
  45342=>"11111111",
  45343=>"00000100",
  45344=>"00000010",
  45345=>"11111111",
  45346=>"11111101",
  45347=>"00000011",
  45348=>"00000100",
  45349=>"00000011",
  45350=>"00000101",
  45351=>"00000111",
  45352=>"00000100",
  45353=>"00000011",
  45354=>"11111110",
  45355=>"00000011",
  45356=>"11111111",
  45357=>"00000000",
  45358=>"11111111",
  45359=>"00000000",
  45360=>"00000000",
  45361=>"00000011",
  45362=>"11111110",
  45363=>"00000010",
  45364=>"00000011",
  45365=>"00000101",
  45366=>"11111111",
  45367=>"00000010",
  45368=>"00000011",
  45369=>"00000001",
  45370=>"00000100",
  45371=>"00001010",
  45372=>"00000000",
  45373=>"11111100",
  45374=>"00000011",
  45375=>"11111110",
  45376=>"00000010",
  45377=>"00000011",
  45378=>"00000010",
  45379=>"11111111",
  45380=>"00000001",
  45381=>"00000010",
  45382=>"11111110",
  45383=>"11111111",
  45384=>"11111110",
  45385=>"00000001",
  45386=>"00000011",
  45387=>"00000001",
  45388=>"00000100",
  45389=>"11111011",
  45390=>"00000001",
  45391=>"00000000",
  45392=>"11111101",
  45393=>"11111111",
  45394=>"11111101",
  45395=>"00000011",
  45396=>"11111101",
  45397=>"00000010",
  45398=>"11111110",
  45399=>"11111101",
  45400=>"11111110",
  45401=>"00000011",
  45402=>"11111101",
  45403=>"00000101",
  45404=>"11111111",
  45405=>"00000000",
  45406=>"11111101",
  45407=>"11111011",
  45408=>"00000011",
  45409=>"00000100",
  45410=>"11111111",
  45411=>"11111110",
  45412=>"11111110",
  45413=>"00000000",
  45414=>"00000010",
  45415=>"11111111",
  45416=>"00000110",
  45417=>"00000000",
  45418=>"11111111",
  45419=>"00000011",
  45420=>"00000101",
  45421=>"00000000",
  45422=>"11111101",
  45423=>"11111110",
  45424=>"00000001",
  45425=>"11111011",
  45426=>"11111011",
  45427=>"00000100",
  45428=>"00000011",
  45429=>"00000011",
  45430=>"00000010",
  45431=>"00000001",
  45432=>"11111110",
  45433=>"00000100",
  45434=>"00000100",
  45435=>"00000011",
  45436=>"00000000",
  45437=>"00000100",
  45438=>"00000011",
  45439=>"00000011",
  45440=>"00000001",
  45441=>"11111110",
  45442=>"00000010",
  45443=>"11111100",
  45444=>"00000001",
  45445=>"00000100",
  45446=>"11111111",
  45447=>"00000001",
  45448=>"11111110",
  45449=>"11111111",
  45450=>"11111100",
  45451=>"00000000",
  45452=>"00000010",
  45453=>"11111011",
  45454=>"00000001",
  45455=>"11111111",
  45456=>"00000001",
  45457=>"00000100",
  45458=>"11110111",
  45459=>"11111101",
  45460=>"00000100",
  45461=>"00000000",
  45462=>"00000000",
  45463=>"00000010",
  45464=>"00000010",
  45465=>"11111101",
  45466=>"00000001",
  45467=>"00000000",
  45468=>"11111101",
  45469=>"11111101",
  45470=>"00000011",
  45471=>"00000011",
  45472=>"11111111",
  45473=>"00000010",
  45474=>"00000110",
  45475=>"11111110",
  45476=>"00000010",
  45477=>"00000001",
  45478=>"00000001",
  45479=>"00000101",
  45480=>"00000101",
  45481=>"00000000",
  45482=>"11111110",
  45483=>"00000000",
  45484=>"11111100",
  45485=>"11111101",
  45486=>"00000100",
  45487=>"00000100",
  45488=>"00000110",
  45489=>"11111110",
  45490=>"11111101",
  45491=>"00000100",
  45492=>"00000011",
  45493=>"11111111",
  45494=>"11111110",
  45495=>"00000011",
  45496=>"00000010",
  45497=>"00000101",
  45498=>"11111101",
  45499=>"00000100",
  45500=>"11111111",
  45501=>"00000100",
  45502=>"00000001",
  45503=>"00000001",
  45504=>"00000010",
  45505=>"11111111",
  45506=>"00000100",
  45507=>"11111100",
  45508=>"00000100",
  45509=>"00000000",
  45510=>"11111101",
  45511=>"00000101",
  45512=>"11111110",
  45513=>"00000000",
  45514=>"00000000",
  45515=>"00000010",
  45516=>"00000100",
  45517=>"00000000",
  45518=>"11111110",
  45519=>"00000001",
  45520=>"00000000",
  45521=>"11111110",
  45522=>"11111111",
  45523=>"11111111",
  45524=>"00000010",
  45525=>"11111110",
  45526=>"11111101",
  45527=>"11111110",
  45528=>"00000010",
  45529=>"00000001",
  45530=>"00000010",
  45531=>"00000011",
  45532=>"11111101",
  45533=>"11111111",
  45534=>"00000100",
  45535=>"11111101",
  45536=>"11111110",
  45537=>"00000010",
  45538=>"00000000",
  45539=>"00000001",
  45540=>"00000011",
  45541=>"00000000",
  45542=>"00000010",
  45543=>"11111111",
  45544=>"00000101",
  45545=>"00000011",
  45546=>"00000101",
  45547=>"00000010",
  45548=>"00000001",
  45549=>"11111110",
  45550=>"00000000",
  45551=>"11111101",
  45552=>"11111110",
  45553=>"00000010",
  45554=>"00000000",
  45555=>"00000011",
  45556=>"00000000",
  45557=>"00000110",
  45558=>"00000100",
  45559=>"11111101",
  45560=>"11111101",
  45561=>"00000001",
  45562=>"00000011",
  45563=>"00000001",
  45564=>"00000100",
  45565=>"00000100",
  45566=>"00000100",
  45567=>"11111101",
  45568=>"11111101",
  45569=>"11111011",
  45570=>"11111101",
  45571=>"00000101",
  45572=>"00000001",
  45573=>"11111111",
  45574=>"00000001",
  45575=>"11111111",
  45576=>"00000000",
  45577=>"11111110",
  45578=>"11111110",
  45579=>"00000001",
  45580=>"11111011",
  45581=>"11111111",
  45582=>"11111101",
  45583=>"11111111",
  45584=>"11111110",
  45585=>"00000001",
  45586=>"11111110",
  45587=>"11111111",
  45588=>"00000011",
  45589=>"11111110",
  45590=>"00000000",
  45591=>"11111101",
  45592=>"00000100",
  45593=>"00000010",
  45594=>"00000100",
  45595=>"00000010",
  45596=>"11111100",
  45597=>"00000001",
  45598=>"11111111",
  45599=>"00000000",
  45600=>"00000000",
  45601=>"11111100",
  45602=>"11111111",
  45603=>"00000011",
  45604=>"00000100",
  45605=>"00000000",
  45606=>"11111110",
  45607=>"11111110",
  45608=>"11111110",
  45609=>"11111111",
  45610=>"11111110",
  45611=>"00000001",
  45612=>"00000011",
  45613=>"11111101",
  45614=>"00000100",
  45615=>"00000010",
  45616=>"00000100",
  45617=>"11111111",
  45618=>"11111111",
  45619=>"00000001",
  45620=>"00000001",
  45621=>"00000011",
  45622=>"00000011",
  45623=>"11111110",
  45624=>"11111111",
  45625=>"00000001",
  45626=>"11111111",
  45627=>"00000011",
  45628=>"00000100",
  45629=>"00000101",
  45630=>"00000010",
  45631=>"11111111",
  45632=>"00000100",
  45633=>"00000011",
  45634=>"00000000",
  45635=>"00000011",
  45636=>"11111101",
  45637=>"00000001",
  45638=>"00000010",
  45639=>"00000011",
  45640=>"00000010",
  45641=>"00000100",
  45642=>"00000001",
  45643=>"00000010",
  45644=>"00000010",
  45645=>"00000000",
  45646=>"11111110",
  45647=>"00000000",
  45648=>"00000010",
  45649=>"00000010",
  45650=>"11111101",
  45651=>"00000000",
  45652=>"00000010",
  45653=>"00000001",
  45654=>"00000011",
  45655=>"00000100",
  45656=>"11111011",
  45657=>"00000000",
  45658=>"11111110",
  45659=>"00000011",
  45660=>"00000000",
  45661=>"11111011",
  45662=>"11111110",
  45663=>"11111111",
  45664=>"11111101",
  45665=>"00000001",
  45666=>"00000010",
  45667=>"00000000",
  45668=>"11111111",
  45669=>"00000000",
  45670=>"11111110",
  45671=>"11111110",
  45672=>"11111101",
  45673=>"11111011",
  45674=>"11111100",
  45675=>"00000100",
  45676=>"00000011",
  45677=>"11111100",
  45678=>"00000000",
  45679=>"00000010",
  45680=>"11111111",
  45681=>"00000001",
  45682=>"00000100",
  45683=>"00000100",
  45684=>"11111101",
  45685=>"00000100",
  45686=>"00000010",
  45687=>"11111111",
  45688=>"11111100",
  45689=>"00000110",
  45690=>"11111110",
  45691=>"00000000",
  45692=>"11111110",
  45693=>"00000001",
  45694=>"00000101",
  45695=>"11111100",
  45696=>"11111100",
  45697=>"11111111",
  45698=>"00000000",
  45699=>"00000001",
  45700=>"00000011",
  45701=>"00000101",
  45702=>"00000011",
  45703=>"00000100",
  45704=>"00000110",
  45705=>"00000010",
  45706=>"00000011",
  45707=>"00000000",
  45708=>"11111111",
  45709=>"11111101",
  45710=>"11111110",
  45711=>"11111110",
  45712=>"00000011",
  45713=>"11111100",
  45714=>"00000000",
  45715=>"00000010",
  45716=>"11111011",
  45717=>"11111110",
  45718=>"11111110",
  45719=>"00000000",
  45720=>"11111011",
  45721=>"11111111",
  45722=>"00000001",
  45723=>"11111100",
  45724=>"00000010",
  45725=>"00000011",
  45726=>"11111101",
  45727=>"00000011",
  45728=>"11111110",
  45729=>"00000010",
  45730=>"11111111",
  45731=>"00000111",
  45732=>"00000001",
  45733=>"00000000",
  45734=>"00000101",
  45735=>"00000000",
  45736=>"00000100",
  45737=>"00000001",
  45738=>"11111110",
  45739=>"11111111",
  45740=>"00000011",
  45741=>"11111110",
  45742=>"00000001",
  45743=>"11111110",
  45744=>"11111111",
  45745=>"00000010",
  45746=>"11111100",
  45747=>"11111111",
  45748=>"11111111",
  45749=>"00000000",
  45750=>"00000000",
  45751=>"00000001",
  45752=>"00000100",
  45753=>"11111110",
  45754=>"00000000",
  45755=>"11111101",
  45756=>"00000000",
  45757=>"00000001",
  45758=>"11111100",
  45759=>"00000000",
  45760=>"00000000",
  45761=>"11111111",
  45762=>"00000000",
  45763=>"00000110",
  45764=>"00000000",
  45765=>"00000001",
  45766=>"00000001",
  45767=>"00000010",
  45768=>"11111101",
  45769=>"00000001",
  45770=>"00000100",
  45771=>"00000100",
  45772=>"00000100",
  45773=>"00000001",
  45774=>"11111111",
  45775=>"11111111",
  45776=>"11111111",
  45777=>"00000100",
  45778=>"00000011",
  45779=>"00000000",
  45780=>"00000001",
  45781=>"11111101",
  45782=>"11111110",
  45783=>"00000011",
  45784=>"11111110",
  45785=>"00000000",
  45786=>"11111101",
  45787=>"00000010",
  45788=>"00000010",
  45789=>"11111110",
  45790=>"11111011",
  45791=>"00000100",
  45792=>"00000010",
  45793=>"00000100",
  45794=>"11111111",
  45795=>"11111101",
  45796=>"11111101",
  45797=>"00000011",
  45798=>"00000000",
  45799=>"11111111",
  45800=>"00000001",
  45801=>"00000010",
  45802=>"00000010",
  45803=>"00000000",
  45804=>"00000000",
  45805=>"11111111",
  45806=>"11111111",
  45807=>"00000101",
  45808=>"11111101",
  45809=>"11111110",
  45810=>"00000000",
  45811=>"11111110",
  45812=>"11111101",
  45813=>"00000100",
  45814=>"00000011",
  45815=>"11111111",
  45816=>"11111111",
  45817=>"00000110",
  45818=>"11111101",
  45819=>"00000100",
  45820=>"11111111",
  45821=>"00000000",
  45822=>"11111011",
  45823=>"00000000",
  45824=>"11111110",
  45825=>"00000001",
  45826=>"00000100",
  45827=>"00000000",
  45828=>"00000001",
  45829=>"00000000",
  45830=>"00000101",
  45831=>"00000000",
  45832=>"00000010",
  45833=>"00000101",
  45834=>"00000000",
  45835=>"00000010",
  45836=>"00000000",
  45837=>"11111100",
  45838=>"00000010",
  45839=>"11111110",
  45840=>"00000010",
  45841=>"11111110",
  45842=>"00000001",
  45843=>"00000011",
  45844=>"00000010",
  45845=>"11111100",
  45846=>"00000000",
  45847=>"11111101",
  45848=>"11111101",
  45849=>"00000001",
  45850=>"00000100",
  45851=>"11111110",
  45852=>"00000010",
  45853=>"00000111",
  45854=>"00000101",
  45855=>"11111010",
  45856=>"00000011",
  45857=>"00000011",
  45858=>"00000000",
  45859=>"00000000",
  45860=>"11111100",
  45861=>"00000011",
  45862=>"11111111",
  45863=>"00000000",
  45864=>"00000010",
  45865=>"00000101",
  45866=>"11111110",
  45867=>"00000010",
  45868=>"00000010",
  45869=>"00000100",
  45870=>"11111111",
  45871=>"11111100",
  45872=>"11111110",
  45873=>"00000101",
  45874=>"00000011",
  45875=>"11111101",
  45876=>"11111100",
  45877=>"11111110",
  45878=>"11111101",
  45879=>"11111101",
  45880=>"00000001",
  45881=>"11111101",
  45882=>"11111110",
  45883=>"11111101",
  45884=>"11111011",
  45885=>"11111101",
  45886=>"11111111",
  45887=>"00000011",
  45888=>"00000101",
  45889=>"00000101",
  45890=>"11111111",
  45891=>"00000001",
  45892=>"11111011",
  45893=>"11111110",
  45894=>"00000000",
  45895=>"00000001",
  45896=>"11111101",
  45897=>"11111111",
  45898=>"11111111",
  45899=>"11111110",
  45900=>"11111101",
  45901=>"11111111",
  45902=>"11111111",
  45903=>"00000010",
  45904=>"11111100",
  45905=>"11111110",
  45906=>"00000011",
  45907=>"11111110",
  45908=>"00000010",
  45909=>"11111101",
  45910=>"11111110",
  45911=>"00000101",
  45912=>"00000001",
  45913=>"00000001",
  45914=>"11111101",
  45915=>"00000000",
  45916=>"00000001",
  45917=>"11111111",
  45918=>"11111111",
  45919=>"11111101",
  45920=>"00000000",
  45921=>"11111101",
  45922=>"00000010",
  45923=>"11111111",
  45924=>"11111111",
  45925=>"11111011",
  45926=>"11111111",
  45927=>"00000100",
  45928=>"00000000",
  45929=>"00000010",
  45930=>"11111101",
  45931=>"00000011",
  45932=>"00000101",
  45933=>"00000010",
  45934=>"00000001",
  45935=>"00000000",
  45936=>"00000011",
  45937=>"00000010",
  45938=>"00000010",
  45939=>"00000010",
  45940=>"00000010",
  45941=>"11111101",
  45942=>"00000000",
  45943=>"00000010",
  45944=>"00000100",
  45945=>"00000010",
  45946=>"11111100",
  45947=>"00000101",
  45948=>"00000011",
  45949=>"00000001",
  45950=>"00000010",
  45951=>"11111101",
  45952=>"00000000",
  45953=>"11111111",
  45954=>"11111110",
  45955=>"00000110",
  45956=>"00000001",
  45957=>"00000010",
  45958=>"00000010",
  45959=>"11111110",
  45960=>"00000100",
  45961=>"00000100",
  45962=>"11111111",
  45963=>"11111110",
  45964=>"11111101",
  45965=>"00000010",
  45966=>"11111100",
  45967=>"11111101",
  45968=>"11111111",
  45969=>"00000000",
  45970=>"00000010",
  45971=>"11111110",
  45972=>"11111110",
  45973=>"00000001",
  45974=>"11111101",
  45975=>"00000100",
  45976=>"00000011",
  45977=>"00000010",
  45978=>"00000101",
  45979=>"00000011",
  45980=>"00000010",
  45981=>"00000011",
  45982=>"00000110",
  45983=>"11111100",
  45984=>"00000001",
  45985=>"11111011",
  45986=>"11111111",
  45987=>"11111110",
  45988=>"00000001",
  45989=>"00000110",
  45990=>"00000000",
  45991=>"11111101",
  45992=>"00000011",
  45993=>"00000011",
  45994=>"11111110",
  45995=>"11111011",
  45996=>"00000100",
  45997=>"00000001",
  45998=>"11111111",
  45999=>"11111101",
  46000=>"00000111",
  46001=>"11111111",
  46002=>"11111111",
  46003=>"00000000",
  46004=>"11111110",
  46005=>"11111101",
  46006=>"11111110",
  46007=>"00000011",
  46008=>"00000001",
  46009=>"11111100",
  46010=>"11111100",
  46011=>"11111111",
  46012=>"00000011",
  46013=>"00000011",
  46014=>"00000000",
  46015=>"00000000",
  46016=>"00000010",
  46017=>"00000000",
  46018=>"00000101",
  46019=>"00000010",
  46020=>"00000001",
  46021=>"11111111",
  46022=>"00000010",
  46023=>"11111111",
  46024=>"11111111",
  46025=>"11111110",
  46026=>"00000000",
  46027=>"00000101",
  46028=>"00000000",
  46029=>"00000010",
  46030=>"11111111",
  46031=>"00000101",
  46032=>"11111100",
  46033=>"00000001",
  46034=>"00000000",
  46035=>"00000001",
  46036=>"00000010",
  46037=>"11111111",
  46038=>"00000110",
  46039=>"11111111",
  46040=>"11111111",
  46041=>"00000011",
  46042=>"00000010",
  46043=>"00000000",
  46044=>"00000001",
  46045=>"00000001",
  46046=>"00000000",
  46047=>"00000011",
  46048=>"00000111",
  46049=>"11111110",
  46050=>"00000001",
  46051=>"00000000",
  46052=>"00000011",
  46053=>"00000100",
  46054=>"00000100",
  46055=>"11111101",
  46056=>"11111011",
  46057=>"11111110",
  46058=>"11111101",
  46059=>"11111101",
  46060=>"11111110",
  46061=>"11111110",
  46062=>"11111111",
  46063=>"11111111",
  46064=>"00000100",
  46065=>"11111111",
  46066=>"11111111",
  46067=>"11111111",
  46068=>"00000001",
  46069=>"11111101",
  46070=>"00000100",
  46071=>"11111111",
  46072=>"00000110",
  46073=>"00000010",
  46074=>"00000010",
  46075=>"00000100",
  46076=>"00000100",
  46077=>"00000000",
  46078=>"00000000",
  46079=>"00000011",
  46080=>"00000001",
  46081=>"11111111",
  46082=>"00000001",
  46083=>"11111111",
  46084=>"00000001",
  46085=>"11111101",
  46086=>"00000000",
  46087=>"00000011",
  46088=>"00000001",
  46089=>"11111110",
  46090=>"00000011",
  46091=>"00000011",
  46092=>"00000000",
  46093=>"00000100",
  46094=>"11111101",
  46095=>"11111101",
  46096=>"11111101",
  46097=>"00000000",
  46098=>"00000101",
  46099=>"00000101",
  46100=>"00000000",
  46101=>"00000010",
  46102=>"11111100",
  46103=>"11111111",
  46104=>"00000000",
  46105=>"00000000",
  46106=>"11111110",
  46107=>"11111111",
  46108=>"00000000",
  46109=>"00000001",
  46110=>"11111101",
  46111=>"11111111",
  46112=>"11111110",
  46113=>"00000001",
  46114=>"00000000",
  46115=>"00000001",
  46116=>"00000011",
  46117=>"00000100",
  46118=>"00000000",
  46119=>"00000000",
  46120=>"11111111",
  46121=>"00000000",
  46122=>"11111110",
  46123=>"00000110",
  46124=>"11111111",
  46125=>"00000000",
  46126=>"11111110",
  46127=>"00000000",
  46128=>"00000100",
  46129=>"00000011",
  46130=>"00000001",
  46131=>"11111111",
  46132=>"00000001",
  46133=>"00000000",
  46134=>"00000011",
  46135=>"00000010",
  46136=>"11111101",
  46137=>"11111100",
  46138=>"11111101",
  46139=>"00000101",
  46140=>"00000001",
  46141=>"00000000",
  46142=>"00000010",
  46143=>"00000010",
  46144=>"00000101",
  46145=>"11111111",
  46146=>"00000001",
  46147=>"00000010",
  46148=>"11111110",
  46149=>"11111110",
  46150=>"11111101",
  46151=>"00000101",
  46152=>"00000001",
  46153=>"11111110",
  46154=>"00000001",
  46155=>"11111110",
  46156=>"00000101",
  46157=>"00000100",
  46158=>"00000011",
  46159=>"00000011",
  46160=>"00000100",
  46161=>"11111111",
  46162=>"11111101",
  46163=>"00000000",
  46164=>"00000011",
  46165=>"11111101",
  46166=>"00000000",
  46167=>"11111101",
  46168=>"11111110",
  46169=>"00000000",
  46170=>"00000010",
  46171=>"00000010",
  46172=>"11111101",
  46173=>"00000011",
  46174=>"00000011",
  46175=>"11111110",
  46176=>"00000101",
  46177=>"11111101",
  46178=>"00000100",
  46179=>"11111110",
  46180=>"11111110",
  46181=>"11111110",
  46182=>"11111100",
  46183=>"00000100",
  46184=>"00000000",
  46185=>"00000000",
  46186=>"11111010",
  46187=>"00000000",
  46188=>"11111111",
  46189=>"00000010",
  46190=>"11111111",
  46191=>"11111111",
  46192=>"11111110",
  46193=>"00000010",
  46194=>"00000101",
  46195=>"11111111",
  46196=>"00000110",
  46197=>"11111101",
  46198=>"11111101",
  46199=>"11111100",
  46200=>"00000001",
  46201=>"00000110",
  46202=>"00000101",
  46203=>"11111101",
  46204=>"00000000",
  46205=>"00000010",
  46206=>"11111110",
  46207=>"11111111",
  46208=>"00000011",
  46209=>"11111111",
  46210=>"00000100",
  46211=>"11111100",
  46212=>"11111101",
  46213=>"00000010",
  46214=>"00000011",
  46215=>"00000001",
  46216=>"00000010",
  46217=>"11111110",
  46218=>"11111111",
  46219=>"11111101",
  46220=>"00000110",
  46221=>"00000000",
  46222=>"00000011",
  46223=>"11111101",
  46224=>"11111101",
  46225=>"00000001",
  46226=>"11111111",
  46227=>"11111110",
  46228=>"00000100",
  46229=>"11111110",
  46230=>"11111101",
  46231=>"00000010",
  46232=>"11111110",
  46233=>"11111101",
  46234=>"00000100",
  46235=>"00000010",
  46236=>"00000010",
  46237=>"11111100",
  46238=>"00000000",
  46239=>"11111101",
  46240=>"11111110",
  46241=>"00000000",
  46242=>"00000001",
  46243=>"11111110",
  46244=>"00000000",
  46245=>"00000000",
  46246=>"11111100",
  46247=>"00000011",
  46248=>"00000100",
  46249=>"11111111",
  46250=>"11111101",
  46251=>"00000000",
  46252=>"00000010",
  46253=>"00000101",
  46254=>"00000000",
  46255=>"11111100",
  46256=>"00000001",
  46257=>"00000001",
  46258=>"00000000",
  46259=>"11111110",
  46260=>"11111100",
  46261=>"11111110",
  46262=>"11111101",
  46263=>"11111111",
  46264=>"00000001",
  46265=>"11111101",
  46266=>"11111111",
  46267=>"11111111",
  46268=>"11111101",
  46269=>"00000010",
  46270=>"00000010",
  46271=>"11111101",
  46272=>"11111110",
  46273=>"11111111",
  46274=>"00000100",
  46275=>"11111111",
  46276=>"00000011",
  46277=>"00000010",
  46278=>"11111111",
  46279=>"00000000",
  46280=>"11111101",
  46281=>"00000001",
  46282=>"00000110",
  46283=>"00000010",
  46284=>"00000010",
  46285=>"11111111",
  46286=>"11111101",
  46287=>"00000011",
  46288=>"00000011",
  46289=>"11111101",
  46290=>"11111111",
  46291=>"00000011",
  46292=>"00000001",
  46293=>"00000000",
  46294=>"00000000",
  46295=>"11111101",
  46296=>"11111110",
  46297=>"00000001",
  46298=>"11111111",
  46299=>"00000000",
  46300=>"00000001",
  46301=>"11111100",
  46302=>"00000010",
  46303=>"00000001",
  46304=>"00000001",
  46305=>"00000001",
  46306=>"11111111",
  46307=>"00000000",
  46308=>"00000000",
  46309=>"00000011",
  46310=>"00000100",
  46311=>"00000000",
  46312=>"00000001",
  46313=>"00000010",
  46314=>"00000001",
  46315=>"11111110",
  46316=>"11111101",
  46317=>"00000001",
  46318=>"11111101",
  46319=>"00000011",
  46320=>"00000010",
  46321=>"11111111",
  46322=>"00000011",
  46323=>"00000000",
  46324=>"00000011",
  46325=>"11111100",
  46326=>"11111111",
  46327=>"11111110",
  46328=>"00000001",
  46329=>"00000011",
  46330=>"00000000",
  46331=>"11111111",
  46332=>"11111101",
  46333=>"00000000",
  46334=>"11111110",
  46335=>"00000001",
  46336=>"00000000",
  46337=>"00000010",
  46338=>"11111100",
  46339=>"00000010",
  46340=>"11111111",
  46341=>"11111011",
  46342=>"00000000",
  46343=>"00000010",
  46344=>"00000011",
  46345=>"11111100",
  46346=>"11111101",
  46347=>"00000110",
  46348=>"00000000",
  46349=>"11111110",
  46350=>"00000010",
  46351=>"11111111",
  46352=>"00000000",
  46353=>"00000000",
  46354=>"00000010",
  46355=>"11111110",
  46356=>"00000001",
  46357=>"11111100",
  46358=>"00000000",
  46359=>"11111101",
  46360=>"11111101",
  46361=>"00000000",
  46362=>"00000001",
  46363=>"11111111",
  46364=>"11111110",
  46365=>"00000001",
  46366=>"00000001",
  46367=>"00000001",
  46368=>"11111111",
  46369=>"00000100",
  46370=>"00000001",
  46371=>"00000000",
  46372=>"00000010",
  46373=>"11111100",
  46374=>"11111111",
  46375=>"00000001",
  46376=>"11111101",
  46377=>"00000010",
  46378=>"00000000",
  46379=>"00000001",
  46380=>"00000001",
  46381=>"11111110",
  46382=>"00000011",
  46383=>"11111111",
  46384=>"11111111",
  46385=>"00000011",
  46386=>"00000001",
  46387=>"11111110",
  46388=>"00000010",
  46389=>"00000000",
  46390=>"00000000",
  46391=>"00000011",
  46392=>"11111100",
  46393=>"11111110",
  46394=>"11111110",
  46395=>"11111101",
  46396=>"00000010",
  46397=>"00000011",
  46398=>"00000100",
  46399=>"11111111",
  46400=>"00000010",
  46401=>"00000000",
  46402=>"00000001",
  46403=>"00000010",
  46404=>"00000001",
  46405=>"11111111",
  46406=>"11111011",
  46407=>"00000010",
  46408=>"00000101",
  46409=>"11111110",
  46410=>"11111110",
  46411=>"00000001",
  46412=>"00000100",
  46413=>"11111110",
  46414=>"11111110",
  46415=>"11111111",
  46416=>"00000010",
  46417=>"00000010",
  46418=>"00000000",
  46419=>"00000001",
  46420=>"00000000",
  46421=>"11111101",
  46422=>"00000011",
  46423=>"11111111",
  46424=>"11111110",
  46425=>"00000010",
  46426=>"00000010",
  46427=>"11111100",
  46428=>"11111111",
  46429=>"00000001",
  46430=>"11111111",
  46431=>"11111101",
  46432=>"11111111",
  46433=>"11111101",
  46434=>"11111111",
  46435=>"00000100",
  46436=>"00000010",
  46437=>"00000001",
  46438=>"00000001",
  46439=>"00000000",
  46440=>"11111100",
  46441=>"00000101",
  46442=>"11111111",
  46443=>"00000011",
  46444=>"11111110",
  46445=>"11111101",
  46446=>"11111101",
  46447=>"00000010",
  46448=>"11111110",
  46449=>"00000000",
  46450=>"00000000",
  46451=>"00000011",
  46452=>"00000100",
  46453=>"11111111",
  46454=>"11111110",
  46455=>"11111111",
  46456=>"00000110",
  46457=>"00000011",
  46458=>"00000100",
  46459=>"11111111",
  46460=>"00000010",
  46461=>"11111110",
  46462=>"00000000",
  46463=>"11111101",
  46464=>"11111111",
  46465=>"00000001",
  46466=>"11111111",
  46467=>"11111110",
  46468=>"00000000",
  46469=>"11111111",
  46470=>"00000000",
  46471=>"00000001",
  46472=>"11111111",
  46473=>"00000100",
  46474=>"11111111",
  46475=>"00000000",
  46476=>"00000001",
  46477=>"00000000",
  46478=>"11111111",
  46479=>"11111011",
  46480=>"00000001",
  46481=>"00000011",
  46482=>"00000000",
  46483=>"11111111",
  46484=>"11111101",
  46485=>"00000010",
  46486=>"00000010",
  46487=>"11111100",
  46488=>"00000000",
  46489=>"11111101",
  46490=>"00000000",
  46491=>"11111111",
  46492=>"11111110",
  46493=>"00000001",
  46494=>"00000001",
  46495=>"00000010",
  46496=>"00000000",
  46497=>"00000100",
  46498=>"00000010",
  46499=>"00000110",
  46500=>"00000001",
  46501=>"00000001",
  46502=>"00000010",
  46503=>"00000100",
  46504=>"11111110",
  46505=>"00000010",
  46506=>"11111111",
  46507=>"00000001",
  46508=>"00000001",
  46509=>"00000000",
  46510=>"11111101",
  46511=>"11111110",
  46512=>"11111111",
  46513=>"00000100",
  46514=>"00000000",
  46515=>"11111111",
  46516=>"00000000",
  46517=>"11111110",
  46518=>"00000000",
  46519=>"11111101",
  46520=>"00000010",
  46521=>"00000110",
  46522=>"00000001",
  46523=>"11111110",
  46524=>"00000010",
  46525=>"11111111",
  46526=>"11111100",
  46527=>"11111110",
  46528=>"11111110",
  46529=>"00000011",
  46530=>"11111100",
  46531=>"00000010",
  46532=>"00000010",
  46533=>"00000000",
  46534=>"11111111",
  46535=>"00000010",
  46536=>"11111111",
  46537=>"00000001",
  46538=>"00000010",
  46539=>"11111100",
  46540=>"11111101",
  46541=>"00000100",
  46542=>"11111110",
  46543=>"00000100",
  46544=>"00000011",
  46545=>"00000011",
  46546=>"11111111",
  46547=>"11111011",
  46548=>"11111111",
  46549=>"00000110",
  46550=>"11111111",
  46551=>"00000010",
  46552=>"00000010",
  46553=>"11111100",
  46554=>"00000100",
  46555=>"11111111",
  46556=>"00000001",
  46557=>"00000010",
  46558=>"00000001",
  46559=>"11111110",
  46560=>"00000110",
  46561=>"00000011",
  46562=>"00000101",
  46563=>"00000000",
  46564=>"00000000",
  46565=>"00000000",
  46566=>"11111101",
  46567=>"00000011",
  46568=>"11111101",
  46569=>"11111101",
  46570=>"11111101",
  46571=>"00000011",
  46572=>"11111110",
  46573=>"11111111",
  46574=>"11111110",
  46575=>"00000010",
  46576=>"00000011",
  46577=>"00000000",
  46578=>"11111101",
  46579=>"11111100",
  46580=>"00000001",
  46581=>"11111110",
  46582=>"00000010",
  46583=>"11111111",
  46584=>"00000010",
  46585=>"00000001",
  46586=>"11111101",
  46587=>"00000000",
  46588=>"00000001",
  46589=>"11111111",
  46590=>"00000000",
  46591=>"00000000",
  46592=>"00000001",
  46593=>"00000010",
  46594=>"11111101",
  46595=>"00000101",
  46596=>"11111111",
  46597=>"11111111",
  46598=>"00000011",
  46599=>"00000001",
  46600=>"00000000",
  46601=>"00000101",
  46602=>"11111111",
  46603=>"00000001",
  46604=>"00000000",
  46605=>"00000001",
  46606=>"11111110",
  46607=>"11111110",
  46608=>"11111101",
  46609=>"00000001",
  46610=>"11111101",
  46611=>"00000000",
  46612=>"11111011",
  46613=>"11111111",
  46614=>"11111110",
  46615=>"00000100",
  46616=>"00000011",
  46617=>"00000000",
  46618=>"11111111",
  46619=>"00000001",
  46620=>"11111100",
  46621=>"11111101",
  46622=>"00000010",
  46623=>"00000010",
  46624=>"11111110",
  46625=>"00000000",
  46626=>"00000100",
  46627=>"00000000",
  46628=>"00000011",
  46629=>"00000001",
  46630=>"00000010",
  46631=>"11111111",
  46632=>"11111111",
  46633=>"00000000",
  46634=>"00000100",
  46635=>"00000000",
  46636=>"00000011",
  46637=>"00000000",
  46638=>"00000011",
  46639=>"00000011",
  46640=>"00000000",
  46641=>"11111110",
  46642=>"00000001",
  46643=>"00000011",
  46644=>"11111111",
  46645=>"11111100",
  46646=>"11111111",
  46647=>"11111101",
  46648=>"11111111",
  46649=>"11111110",
  46650=>"00000010",
  46651=>"11111111",
  46652=>"11111111",
  46653=>"11111011",
  46654=>"00000110",
  46655=>"00000000",
  46656=>"00000000",
  46657=>"00000000",
  46658=>"00000101",
  46659=>"11111110",
  46660=>"00000001",
  46661=>"00000100",
  46662=>"00000000",
  46663=>"11111111",
  46664=>"11111110",
  46665=>"11111111",
  46666=>"00000000",
  46667=>"00000011",
  46668=>"00000001",
  46669=>"00000000",
  46670=>"00000101",
  46671=>"00000001",
  46672=>"00000000",
  46673=>"00000001",
  46674=>"11111111",
  46675=>"00000001",
  46676=>"00000001",
  46677=>"00000101",
  46678=>"00000011",
  46679=>"00000010",
  46680=>"11111101",
  46681=>"11111111",
  46682=>"00000000",
  46683=>"00000001",
  46684=>"11111111",
  46685=>"00000000",
  46686=>"11111110",
  46687=>"00000011",
  46688=>"00000010",
  46689=>"11111101",
  46690=>"11111101",
  46691=>"00000010",
  46692=>"11111110",
  46693=>"00000001",
  46694=>"00000010",
  46695=>"11111110",
  46696=>"00000100",
  46697=>"00000001",
  46698=>"00000011",
  46699=>"00000001",
  46700=>"11111110",
  46701=>"00000000",
  46702=>"11111110",
  46703=>"00000111",
  46704=>"11111110",
  46705=>"00000001",
  46706=>"11111111",
  46707=>"00000100",
  46708=>"00000000",
  46709=>"11111110",
  46710=>"00000111",
  46711=>"00000001",
  46712=>"00000000",
  46713=>"00000010",
  46714=>"11111101",
  46715=>"11111101",
  46716=>"11111110",
  46717=>"00000000",
  46718=>"11111100",
  46719=>"00000001",
  46720=>"00000000",
  46721=>"11111101",
  46722=>"11111111",
  46723=>"00000000",
  46724=>"00000011",
  46725=>"11111101",
  46726=>"00000001",
  46727=>"00000011",
  46728=>"00000111",
  46729=>"00000001",
  46730=>"00000010",
  46731=>"11111110",
  46732=>"00000000",
  46733=>"00000010",
  46734=>"00000010",
  46735=>"00000000",
  46736=>"11111101",
  46737=>"00000000",
  46738=>"11111101",
  46739=>"00000001",
  46740=>"00000010",
  46741=>"00000000",
  46742=>"11111101",
  46743=>"11111111",
  46744=>"00000010",
  46745=>"11111110",
  46746=>"00000000",
  46747=>"00000001",
  46748=>"00000100",
  46749=>"11111111",
  46750=>"11111110",
  46751=>"11111100",
  46752=>"00000100",
  46753=>"00000010",
  46754=>"00000000",
  46755=>"00000010",
  46756=>"11111110",
  46757=>"11111100",
  46758=>"00000001",
  46759=>"11111110",
  46760=>"00000001",
  46761=>"11111101",
  46762=>"11111110",
  46763=>"00000011",
  46764=>"00000010",
  46765=>"11111111",
  46766=>"00000010",
  46767=>"00000010",
  46768=>"00000001",
  46769=>"00000010",
  46770=>"00000000",
  46771=>"11111110",
  46772=>"11111111",
  46773=>"00000010",
  46774=>"11111111",
  46775=>"11111100",
  46776=>"11111101",
  46777=>"00000100",
  46778=>"00000011",
  46779=>"00000010",
  46780=>"00000010",
  46781=>"11111110",
  46782=>"00000011",
  46783=>"00000000",
  46784=>"11111101",
  46785=>"11111111",
  46786=>"11111110",
  46787=>"11111110",
  46788=>"11111111",
  46789=>"00000100",
  46790=>"00000000",
  46791=>"11111111",
  46792=>"00000010",
  46793=>"00000000",
  46794=>"11111100",
  46795=>"11111111",
  46796=>"00000011",
  46797=>"11111111",
  46798=>"11111111",
  46799=>"00000001",
  46800=>"11111111",
  46801=>"00000010",
  46802=>"00000010",
  46803=>"00000001",
  46804=>"11111110",
  46805=>"11111101",
  46806=>"00000001",
  46807=>"00000001",
  46808=>"11111100",
  46809=>"00000000",
  46810=>"11111110",
  46811=>"00000010",
  46812=>"00000100",
  46813=>"00000101",
  46814=>"11111100",
  46815=>"00000010",
  46816=>"11111100",
  46817=>"11111100",
  46818=>"11111110",
  46819=>"00000010",
  46820=>"00000011",
  46821=>"00000001",
  46822=>"00000010",
  46823=>"00000010",
  46824=>"11111111",
  46825=>"00000010",
  46826=>"00000100",
  46827=>"11111111",
  46828=>"11111111",
  46829=>"11111101",
  46830=>"00000010",
  46831=>"11111110",
  46832=>"00000011",
  46833=>"00000001",
  46834=>"11111100",
  46835=>"00000011",
  46836=>"00000001",
  46837=>"00000001",
  46838=>"11111110",
  46839=>"00000010",
  46840=>"11111111",
  46841=>"11111110",
  46842=>"11111110",
  46843=>"00000011",
  46844=>"11111110",
  46845=>"11111101",
  46846=>"00000001",
  46847=>"00000001",
  46848=>"11111111",
  46849=>"00000100",
  46850=>"11111110",
  46851=>"11111110",
  46852=>"00000000",
  46853=>"00000011",
  46854=>"11111110",
  46855=>"00000010",
  46856=>"00000001",
  46857=>"00000001",
  46858=>"11111111",
  46859=>"00000011",
  46860=>"11111101",
  46861=>"11111110",
  46862=>"11111101",
  46863=>"00000001",
  46864=>"00000001",
  46865=>"11111111",
  46866=>"00000001",
  46867=>"11111111",
  46868=>"11111110",
  46869=>"00000101",
  46870=>"11111110",
  46871=>"11111100",
  46872=>"11111101",
  46873=>"11111101",
  46874=>"11111100",
  46875=>"11111110",
  46876=>"00000001",
  46877=>"00000001",
  46878=>"00000101",
  46879=>"00000000",
  46880=>"11111111",
  46881=>"00000001",
  46882=>"00000000",
  46883=>"00000011",
  46884=>"00000000",
  46885=>"11111111",
  46886=>"00000001",
  46887=>"11111110",
  46888=>"00000001",
  46889=>"00000000",
  46890=>"11111101",
  46891=>"00000011",
  46892=>"00000001",
  46893=>"11111111",
  46894=>"00000000",
  46895=>"11111111",
  46896=>"00000010",
  46897=>"11111100",
  46898=>"00000000",
  46899=>"00000010",
  46900=>"00000100",
  46901=>"00000011",
  46902=>"00000100",
  46903=>"00000011",
  46904=>"00000010",
  46905=>"00000010",
  46906=>"00000010",
  46907=>"00000010",
  46908=>"11111111",
  46909=>"00000001",
  46910=>"00000100",
  46911=>"11111010",
  46912=>"11111110",
  46913=>"11111111",
  46914=>"00000001",
  46915=>"00000011",
  46916=>"00000110",
  46917=>"11111111",
  46918=>"00000010",
  46919=>"00000010",
  46920=>"11111100",
  46921=>"11111101",
  46922=>"00000000",
  46923=>"00000010",
  46924=>"00000000",
  46925=>"00000010",
  46926=>"11111110",
  46927=>"00000100",
  46928=>"00000000",
  46929=>"00000010",
  46930=>"00000000",
  46931=>"00000010",
  46932=>"00000000",
  46933=>"00000001",
  46934=>"11111111",
  46935=>"11111111",
  46936=>"11111111",
  46937=>"00000000",
  46938=>"11111101",
  46939=>"11111100",
  46940=>"00000011",
  46941=>"00000100",
  46942=>"11111100",
  46943=>"11111101",
  46944=>"11111100",
  46945=>"00000001",
  46946=>"00000100",
  46947=>"11111110",
  46948=>"11111111",
  46949=>"00000110",
  46950=>"00000010",
  46951=>"11111110",
  46952=>"00000111",
  46953=>"11111011",
  46954=>"00000101",
  46955=>"00000000",
  46956=>"00000001",
  46957=>"11111101",
  46958=>"11111110",
  46959=>"11111101",
  46960=>"00000011",
  46961=>"11111111",
  46962=>"00000001",
  46963=>"11111100",
  46964=>"00000000",
  46965=>"11111101",
  46966=>"00000001",
  46967=>"00000000",
  46968=>"11111110",
  46969=>"00000010",
  46970=>"00000011",
  46971=>"11111110",
  46972=>"11111111",
  46973=>"00000110",
  46974=>"11111111",
  46975=>"00000011",
  46976=>"00000001",
  46977=>"11111101",
  46978=>"00000010",
  46979=>"00000001",
  46980=>"11111110",
  46981=>"00000010",
  46982=>"11111101",
  46983=>"11111101",
  46984=>"00000001",
  46985=>"11111110",
  46986=>"00000000",
  46987=>"11111110",
  46988=>"11111101",
  46989=>"00000010",
  46990=>"00000011",
  46991=>"00000011",
  46992=>"00000001",
  46993=>"00000100",
  46994=>"11111110",
  46995=>"00000011",
  46996=>"00000001",
  46997=>"00000010",
  46998=>"00000001",
  46999=>"00000011",
  47000=>"00000001",
  47001=>"00000000",
  47002=>"00000011",
  47003=>"11111100",
  47004=>"11111110",
  47005=>"11111110",
  47006=>"00000011",
  47007=>"00000011",
  47008=>"11111111",
  47009=>"00000010",
  47010=>"11111111",
  47011=>"00000001",
  47012=>"11111111",
  47013=>"00000010",
  47014=>"00000010",
  47015=>"11111101",
  47016=>"00000011",
  47017=>"11111111",
  47018=>"00000001",
  47019=>"00000011",
  47020=>"00000101",
  47021=>"11111110",
  47022=>"00000100",
  47023=>"00000001",
  47024=>"11111111",
  47025=>"11111100",
  47026=>"11111111",
  47027=>"11111110",
  47028=>"00000011",
  47029=>"11111101",
  47030=>"00000111",
  47031=>"11111110",
  47032=>"00000000",
  47033=>"00000010",
  47034=>"11111111",
  47035=>"00000010",
  47036=>"11111101",
  47037=>"11111101",
  47038=>"00000010",
  47039=>"00000000",
  47040=>"11111100",
  47041=>"00000000",
  47042=>"11111101",
  47043=>"00000000",
  47044=>"00000000",
  47045=>"00000110",
  47046=>"00000011",
  47047=>"11111101",
  47048=>"11111110",
  47049=>"00000000",
  47050=>"11111101",
  47051=>"11111110",
  47052=>"00000001",
  47053=>"00000100",
  47054=>"00000011",
  47055=>"11111101",
  47056=>"00000011",
  47057=>"11111101",
  47058=>"00000000",
  47059=>"00000001",
  47060=>"00000000",
  47061=>"00000001",
  47062=>"11111110",
  47063=>"00000011",
  47064=>"11111111",
  47065=>"00000000",
  47066=>"00000010",
  47067=>"00000000",
  47068=>"00000101",
  47069=>"00000000",
  47070=>"00000011",
  47071=>"00000010",
  47072=>"00000110",
  47073=>"11111101",
  47074=>"11111111",
  47075=>"11111110",
  47076=>"11111101",
  47077=>"11111111",
  47078=>"11111110",
  47079=>"00000000",
  47080=>"11111110",
  47081=>"11111111",
  47082=>"00000010",
  47083=>"00000010",
  47084=>"11111110",
  47085=>"11111110",
  47086=>"11111111",
  47087=>"11111111",
  47088=>"00000000",
  47089=>"00000001",
  47090=>"00000101",
  47091=>"00000100",
  47092=>"11111110",
  47093=>"11111101",
  47094=>"00000110",
  47095=>"11111101",
  47096=>"00000101",
  47097=>"00000011",
  47098=>"00000010",
  47099=>"00000000",
  47100=>"11111101",
  47101=>"00000000",
  47102=>"00000010",
  47103=>"11111110",
  47104=>"00000010",
  47105=>"00000001",
  47106=>"00000000",
  47107=>"00000011",
  47108=>"00000000",
  47109=>"00000000",
  47110=>"11111101",
  47111=>"11111101",
  47112=>"11111100",
  47113=>"00000101",
  47114=>"11111111",
  47115=>"00000000",
  47116=>"00000010",
  47117=>"00000000",
  47118=>"00000000",
  47119=>"00000001",
  47120=>"00000001",
  47121=>"11111111",
  47122=>"11111110",
  47123=>"11111111",
  47124=>"11111110",
  47125=>"11111110",
  47126=>"00000110",
  47127=>"11111101",
  47128=>"00000001",
  47129=>"00000000",
  47130=>"00000000",
  47131=>"11111101",
  47132=>"00000000",
  47133=>"11111101",
  47134=>"11111110",
  47135=>"11111100",
  47136=>"00000101",
  47137=>"00000010",
  47138=>"00000010",
  47139=>"00000001",
  47140=>"00000000",
  47141=>"11111101",
  47142=>"00000101",
  47143=>"00000000",
  47144=>"00000010",
  47145=>"11111100",
  47146=>"00000000",
  47147=>"11111111",
  47148=>"11111111",
  47149=>"00000100",
  47150=>"11111110",
  47151=>"00000011",
  47152=>"11111111",
  47153=>"11111110",
  47154=>"11111110",
  47155=>"00000000",
  47156=>"00000000",
  47157=>"11111110",
  47158=>"00000001",
  47159=>"00000001",
  47160=>"00000100",
  47161=>"00000000",
  47162=>"11111111",
  47163=>"11111110",
  47164=>"00000000",
  47165=>"00000001",
  47166=>"11111111",
  47167=>"11111111",
  47168=>"11111110",
  47169=>"11111111",
  47170=>"00000100",
  47171=>"00000001",
  47172=>"00000011",
  47173=>"00000010",
  47174=>"11111101",
  47175=>"11111101",
  47176=>"00000010",
  47177=>"00000100",
  47178=>"00000000",
  47179=>"00000000",
  47180=>"00000101",
  47181=>"00000000",
  47182=>"11111111",
  47183=>"00000010",
  47184=>"11111011",
  47185=>"00000000",
  47186=>"00000010",
  47187=>"11111111",
  47188=>"00000011",
  47189=>"00000001",
  47190=>"00000011",
  47191=>"00000010",
  47192=>"00000001",
  47193=>"11111110",
  47194=>"11111110",
  47195=>"11111110",
  47196=>"11111100",
  47197=>"00000010",
  47198=>"00000011",
  47199=>"11111111",
  47200=>"11111101",
  47201=>"00000000",
  47202=>"11111101",
  47203=>"00000000",
  47204=>"11111111",
  47205=>"00000000",
  47206=>"00000001",
  47207=>"11111110",
  47208=>"11111101",
  47209=>"11111111",
  47210=>"00000100",
  47211=>"00000001",
  47212=>"11111100",
  47213=>"11111101",
  47214=>"00000110",
  47215=>"11111110",
  47216=>"00000001",
  47217=>"00000000",
  47218=>"00000010",
  47219=>"00000001",
  47220=>"00000010",
  47221=>"00000011",
  47222=>"00000101",
  47223=>"00000010",
  47224=>"00000010",
  47225=>"00000010",
  47226=>"11111101",
  47227=>"00000010",
  47228=>"00000000",
  47229=>"00000000",
  47230=>"11111110",
  47231=>"00000100",
  47232=>"11111111",
  47233=>"00000000",
  47234=>"11111110",
  47235=>"00000011",
  47236=>"00000001",
  47237=>"11111110",
  47238=>"11111111",
  47239=>"00000011",
  47240=>"11111111",
  47241=>"11111110",
  47242=>"00000100",
  47243=>"00000001",
  47244=>"11111101",
  47245=>"00000100",
  47246=>"00000001",
  47247=>"00000011",
  47248=>"00000000",
  47249=>"11111111",
  47250=>"00000001",
  47251=>"11111111",
  47252=>"00000100",
  47253=>"11111101",
  47254=>"11111101",
  47255=>"00000001",
  47256=>"00000100",
  47257=>"11111111",
  47258=>"00000000",
  47259=>"00000000",
  47260=>"11111110",
  47261=>"00000001",
  47262=>"11111110",
  47263=>"00000000",
  47264=>"11111110",
  47265=>"00000001",
  47266=>"00000000",
  47267=>"11111101",
  47268=>"00000001",
  47269=>"00000001",
  47270=>"11111101",
  47271=>"00000011",
  47272=>"00000000",
  47273=>"11111011",
  47274=>"00000100",
  47275=>"00000010",
  47276=>"00000101",
  47277=>"11111110",
  47278=>"00000000",
  47279=>"11111111",
  47280=>"00000010",
  47281=>"11111110",
  47282=>"00000000",
  47283=>"00000001",
  47284=>"11111111",
  47285=>"00001000",
  47286=>"00000000",
  47287=>"00000000",
  47288=>"00000000",
  47289=>"11111110",
  47290=>"11111110",
  47291=>"11111111",
  47292=>"11111100",
  47293=>"11111111",
  47294=>"11111110",
  47295=>"11111110",
  47296=>"00000001",
  47297=>"00000000",
  47298=>"00000000",
  47299=>"11111110",
  47300=>"11111101",
  47301=>"11111111",
  47302=>"11111100",
  47303=>"00000001",
  47304=>"00000011",
  47305=>"00000010",
  47306=>"11111111",
  47307=>"11111110",
  47308=>"11111101",
  47309=>"11111110",
  47310=>"00000011",
  47311=>"00000010",
  47312=>"11111111",
  47313=>"00000011",
  47314=>"00000001",
  47315=>"11111101",
  47316=>"00000000",
  47317=>"11111100",
  47318=>"00000000",
  47319=>"00000101",
  47320=>"00000000",
  47321=>"11111111",
  47322=>"11111111",
  47323=>"11111110",
  47324=>"00000001",
  47325=>"11111110",
  47326=>"00000100",
  47327=>"11111111",
  47328=>"00000001",
  47329=>"11111100",
  47330=>"00000000",
  47331=>"11111101",
  47332=>"00000000",
  47333=>"00000001",
  47334=>"00000001",
  47335=>"11111101",
  47336=>"00000000",
  47337=>"11111101",
  47338=>"00000000",
  47339=>"00000001",
  47340=>"11111111",
  47341=>"11111111",
  47342=>"11111111",
  47343=>"00000010",
  47344=>"00000001",
  47345=>"11111101",
  47346=>"00000001",
  47347=>"11111110",
  47348=>"11111110",
  47349=>"11111111",
  47350=>"11111110",
  47351=>"11111111",
  47352=>"00000010",
  47353=>"00000000",
  47354=>"00000010",
  47355=>"00000001",
  47356=>"00000011",
  47357=>"11111111",
  47358=>"11111111",
  47359=>"00000001",
  47360=>"00000000",
  47361=>"00000001",
  47362=>"00000011",
  47363=>"11111100",
  47364=>"00000001",
  47365=>"00000000",
  47366=>"11111101",
  47367=>"11111101",
  47368=>"00000001",
  47369=>"00000001",
  47370=>"00000011",
  47371=>"11111101",
  47372=>"11111110",
  47373=>"11111101",
  47374=>"00000101",
  47375=>"00000110",
  47376=>"11111110",
  47377=>"00000001",
  47378=>"11111101",
  47379=>"11111110",
  47380=>"11111101",
  47381=>"11111111",
  47382=>"00000010",
  47383=>"11111101",
  47384=>"00000001",
  47385=>"00000001",
  47386=>"00000100",
  47387=>"00000010",
  47388=>"00000001",
  47389=>"11111101",
  47390=>"00000001",
  47391=>"11111110",
  47392=>"00000100",
  47393=>"00000001",
  47394=>"11111111",
  47395=>"11111111",
  47396=>"11111110",
  47397=>"11111111",
  47398=>"00000010",
  47399=>"11111100",
  47400=>"11111101",
  47401=>"11111101",
  47402=>"11111101",
  47403=>"11111110",
  47404=>"11111111",
  47405=>"11111111",
  47406=>"00000010",
  47407=>"00000010",
  47408=>"00000110",
  47409=>"11111110",
  47410=>"00000001",
  47411=>"11111111",
  47412=>"11111111",
  47413=>"00000000",
  47414=>"11111110",
  47415=>"00000000",
  47416=>"11111101",
  47417=>"11111110",
  47418=>"11111111",
  47419=>"00000010",
  47420=>"11111111",
  47421=>"11111101",
  47422=>"11111111",
  47423=>"11111111",
  47424=>"00000001",
  47425=>"00000010",
  47426=>"00000010",
  47427=>"11111101",
  47428=>"11111101",
  47429=>"00000000",
  47430=>"11111110",
  47431=>"11111110",
  47432=>"00000101",
  47433=>"11111100",
  47434=>"11111110",
  47435=>"00000000",
  47436=>"11111111",
  47437=>"11111111",
  47438=>"00000010",
  47439=>"11111111",
  47440=>"00000100",
  47441=>"00000000",
  47442=>"00000000",
  47443=>"11111110",
  47444=>"11111110",
  47445=>"00000100",
  47446=>"00000000",
  47447=>"00000000",
  47448=>"11111110",
  47449=>"00000011",
  47450=>"11111110",
  47451=>"00000010",
  47452=>"00000010",
  47453=>"00000000",
  47454=>"11111111",
  47455=>"00000010",
  47456=>"11111110",
  47457=>"11111100",
  47458=>"00000001",
  47459=>"11111110",
  47460=>"00000001",
  47461=>"00000010",
  47462=>"00000000",
  47463=>"00000000",
  47464=>"11111110",
  47465=>"00000010",
  47466=>"00000001",
  47467=>"11111101",
  47468=>"11111101",
  47469=>"11111110",
  47470=>"00000101",
  47471=>"00000000",
  47472=>"11111110",
  47473=>"11111110",
  47474=>"00000001",
  47475=>"11111111",
  47476=>"00000011",
  47477=>"11111101",
  47478=>"00000001",
  47479=>"00000001",
  47480=>"11111110",
  47481=>"00000000",
  47482=>"11111111",
  47483=>"11111101",
  47484=>"11111111",
  47485=>"00000001",
  47486=>"00000100",
  47487=>"11111111",
  47488=>"00000001",
  47489=>"00000001",
  47490=>"00000000",
  47491=>"11111110",
  47492=>"00000000",
  47493=>"11111101",
  47494=>"00000000",
  47495=>"00000000",
  47496=>"00000010",
  47497=>"00000001",
  47498=>"00000100",
  47499=>"00000011",
  47500=>"00000101",
  47501=>"00000010",
  47502=>"00000011",
  47503=>"11111101",
  47504=>"00000000",
  47505=>"11111111",
  47506=>"00000100",
  47507=>"00000001",
  47508=>"11111111",
  47509=>"11111101",
  47510=>"00000000",
  47511=>"00000011",
  47512=>"11111100",
  47513=>"00000000",
  47514=>"11111111",
  47515=>"11111110",
  47516=>"00000101",
  47517=>"00000010",
  47518=>"00000011",
  47519=>"00000010",
  47520=>"11111101",
  47521=>"00000000",
  47522=>"00000101",
  47523=>"00000000",
  47524=>"00000010",
  47525=>"00000011",
  47526=>"00000110",
  47527=>"11111111",
  47528=>"00000001",
  47529=>"00000100",
  47530=>"00000001",
  47531=>"00000010",
  47532=>"00000000",
  47533=>"11111101",
  47534=>"11111100",
  47535=>"11111110",
  47536=>"00000000",
  47537=>"11111111",
  47538=>"11111101",
  47539=>"00000011",
  47540=>"00000010",
  47541=>"00000001",
  47542=>"00000010",
  47543=>"00000100",
  47544=>"00000011",
  47545=>"11111110",
  47546=>"11111110",
  47547=>"00000001",
  47548=>"00000010",
  47549=>"11111110",
  47550=>"11111111",
  47551=>"00000011",
  47552=>"00000000",
  47553=>"00000101",
  47554=>"00000000",
  47555=>"11111110",
  47556=>"11111110",
  47557=>"11111111",
  47558=>"11111100",
  47559=>"11111101",
  47560=>"00000000",
  47561=>"00000010",
  47562=>"11111110",
  47563=>"11111110",
  47564=>"00000100",
  47565=>"11111110",
  47566=>"00000001",
  47567=>"11111110",
  47568=>"00000001",
  47569=>"00000001",
  47570=>"11111110",
  47571=>"00000000",
  47572=>"11111110",
  47573=>"00000000",
  47574=>"00000000",
  47575=>"11111111",
  47576=>"11111110",
  47577=>"11111110",
  47578=>"00000010",
  47579=>"00000011",
  47580=>"00000000",
  47581=>"11111100",
  47582=>"00000001",
  47583=>"11111110",
  47584=>"11111101",
  47585=>"11111101",
  47586=>"00000000",
  47587=>"00000000",
  47588=>"00000010",
  47589=>"00000000",
  47590=>"00000001",
  47591=>"11111110",
  47592=>"11111111",
  47593=>"00000011",
  47594=>"11111110",
  47595=>"11111110",
  47596=>"11111110",
  47597=>"00000001",
  47598=>"00000000",
  47599=>"00000010",
  47600=>"11111111",
  47601=>"00000011",
  47602=>"11111111",
  47603=>"00000000",
  47604=>"00000000",
  47605=>"00000000",
  47606=>"00000001",
  47607=>"00000010",
  47608=>"00000100",
  47609=>"00000011",
  47610=>"00000001",
  47611=>"00000000",
  47612=>"00000011",
  47613=>"00000001",
  47614=>"00000000",
  47615=>"00000011",
  47616=>"00000011",
  47617=>"11111111",
  47618=>"11111111",
  47619=>"00000000",
  47620=>"11111101",
  47621=>"11111110",
  47622=>"00000001",
  47623=>"00000011",
  47624=>"11111110",
  47625=>"00000110",
  47626=>"00000011",
  47627=>"11111110",
  47628=>"00000001",
  47629=>"00000001",
  47630=>"00000010",
  47631=>"00000110",
  47632=>"00000011",
  47633=>"11111110",
  47634=>"00000001",
  47635=>"11111101",
  47636=>"00000000",
  47637=>"00000000",
  47638=>"11111111",
  47639=>"11111110",
  47640=>"00000010",
  47641=>"11111110",
  47642=>"11111100",
  47643=>"00000010",
  47644=>"00000001",
  47645=>"00000010",
  47646=>"00000001",
  47647=>"00000001",
  47648=>"11111101",
  47649=>"00000010",
  47650=>"11111101",
  47651=>"11111111",
  47652=>"11111101",
  47653=>"00000011",
  47654=>"11111101",
  47655=>"11111111",
  47656=>"00000010",
  47657=>"11111101",
  47658=>"00000000",
  47659=>"11111111",
  47660=>"00000001",
  47661=>"00000000",
  47662=>"11111111",
  47663=>"11111101",
  47664=>"11111111",
  47665=>"11111101",
  47666=>"00000001",
  47667=>"11111110",
  47668=>"11111111",
  47669=>"00000011",
  47670=>"00000010",
  47671=>"11111111",
  47672=>"00000001",
  47673=>"00000010",
  47674=>"11111110",
  47675=>"00000000",
  47676=>"11111111",
  47677=>"00000001",
  47678=>"11111110",
  47679=>"00000000",
  47680=>"00000001",
  47681=>"00000010",
  47682=>"11111101",
  47683=>"00000011",
  47684=>"00000010",
  47685=>"11111110",
  47686=>"11111101",
  47687=>"11111111",
  47688=>"00000000",
  47689=>"00000000",
  47690=>"11111101",
  47691=>"11111100",
  47692=>"00000011",
  47693=>"00000000",
  47694=>"11111110",
  47695=>"00000000",
  47696=>"00000010",
  47697=>"00000011",
  47698=>"00000011",
  47699=>"11111110",
  47700=>"00000011",
  47701=>"00000000",
  47702=>"00000000",
  47703=>"00000001",
  47704=>"11111110",
  47705=>"00000010",
  47706=>"11111111",
  47707=>"00000100",
  47708=>"00000001",
  47709=>"00000001",
  47710=>"00000010",
  47711=>"11111101",
  47712=>"11111101",
  47713=>"00000100",
  47714=>"11111110",
  47715=>"00000001",
  47716=>"11111101",
  47717=>"11111100",
  47718=>"00000000",
  47719=>"00000000",
  47720=>"00000011",
  47721=>"11111110",
  47722=>"00000000",
  47723=>"00000000",
  47724=>"00000001",
  47725=>"00000111",
  47726=>"11111101",
  47727=>"00000000",
  47728=>"00000010",
  47729=>"00000001",
  47730=>"00000001",
  47731=>"00000000",
  47732=>"11111111",
  47733=>"11111101",
  47734=>"11111111",
  47735=>"00000000",
  47736=>"00000010",
  47737=>"00000000",
  47738=>"11111110",
  47739=>"00000000",
  47740=>"11111110",
  47741=>"00000010",
  47742=>"00000000",
  47743=>"00000000",
  47744=>"00000001",
  47745=>"00000001",
  47746=>"11111101",
  47747=>"11111111",
  47748=>"00000000",
  47749=>"11111111",
  47750=>"11111101",
  47751=>"00000000",
  47752=>"00000010",
  47753=>"00000001",
  47754=>"00000010",
  47755=>"11111111",
  47756=>"00000001",
  47757=>"00000011",
  47758=>"11111110",
  47759=>"11111111",
  47760=>"00000000",
  47761=>"00000110",
  47762=>"11111110",
  47763=>"00000011",
  47764=>"11111100",
  47765=>"00000000",
  47766=>"00000000",
  47767=>"11111101",
  47768=>"11111111",
  47769=>"00000101",
  47770=>"00000101",
  47771=>"00000001",
  47772=>"00000010",
  47773=>"11111101",
  47774=>"00000110",
  47775=>"00000000",
  47776=>"00000010",
  47777=>"11111101",
  47778=>"11111110",
  47779=>"00000000",
  47780=>"00000011",
  47781=>"11111110",
  47782=>"11111011",
  47783=>"11111111",
  47784=>"11111111",
  47785=>"11111101",
  47786=>"00000011",
  47787=>"00000011",
  47788=>"00000011",
  47789=>"11111110",
  47790=>"11111110",
  47791=>"00000000",
  47792=>"00000010",
  47793=>"00000001",
  47794=>"00000010",
  47795=>"11111011",
  47796=>"11111110",
  47797=>"11111101",
  47798=>"11111110",
  47799=>"00000000",
  47800=>"11111100",
  47801=>"00000010",
  47802=>"00000010",
  47803=>"00000100",
  47804=>"00000011",
  47805=>"00000001",
  47806=>"00000000",
  47807=>"00000010",
  47808=>"11111101",
  47809=>"00000001",
  47810=>"00000001",
  47811=>"00000000",
  47812=>"11111111",
  47813=>"00000010",
  47814=>"11111110",
  47815=>"00000010",
  47816=>"00000000",
  47817=>"00000001",
  47818=>"11111111",
  47819=>"11111111",
  47820=>"11111101",
  47821=>"00000111",
  47822=>"11111110",
  47823=>"00000100",
  47824=>"00000000",
  47825=>"00000010",
  47826=>"00000010",
  47827=>"00000011",
  47828=>"00000011",
  47829=>"11111101",
  47830=>"11111101",
  47831=>"11111100",
  47832=>"00000110",
  47833=>"00000001",
  47834=>"11111110",
  47835=>"00000001",
  47836=>"00000000",
  47837=>"00000001",
  47838=>"00000001",
  47839=>"00000000",
  47840=>"11111111",
  47841=>"11111110",
  47842=>"00000001",
  47843=>"00000001",
  47844=>"00000100",
  47845=>"11111111",
  47846=>"11111111",
  47847=>"00000010",
  47848=>"11111111",
  47849=>"11111101",
  47850=>"11111101",
  47851=>"00000000",
  47852=>"11111111",
  47853=>"11111111",
  47854=>"11111101",
  47855=>"00000010",
  47856=>"11111101",
  47857=>"11111111",
  47858=>"11111110",
  47859=>"11111111",
  47860=>"11111101",
  47861=>"11111111",
  47862=>"11111111",
  47863=>"00000000",
  47864=>"11111101",
  47865=>"11111110",
  47866=>"11111111",
  47867=>"00000001",
  47868=>"00000010",
  47869=>"11111100",
  47870=>"11111111",
  47871=>"00000000",
  47872=>"11111111",
  47873=>"00000001",
  47874=>"11111101",
  47875=>"11111111",
  47876=>"11111100",
  47877=>"11111101",
  47878=>"00000010",
  47879=>"11111110",
  47880=>"11111101",
  47881=>"11111110",
  47882=>"00000011",
  47883=>"11111111",
  47884=>"00000011",
  47885=>"11111101",
  47886=>"11111101",
  47887=>"00000010",
  47888=>"00000000",
  47889=>"11111110",
  47890=>"11111101",
  47891=>"00000011",
  47892=>"00000000",
  47893=>"11111110",
  47894=>"11111111",
  47895=>"00000010",
  47896=>"00000001",
  47897=>"00000000",
  47898=>"00000000",
  47899=>"00000000",
  47900=>"00000001",
  47901=>"11111011",
  47902=>"11111011",
  47903=>"11111101",
  47904=>"00000000",
  47905=>"11111111",
  47906=>"00000001",
  47907=>"00000011",
  47908=>"11111111",
  47909=>"11111111",
  47910=>"11111101",
  47911=>"11111111",
  47912=>"00000001",
  47913=>"11111100",
  47914=>"11111011",
  47915=>"11111100",
  47916=>"11111110",
  47917=>"11111101",
  47918=>"00000011",
  47919=>"00000001",
  47920=>"00000000",
  47921=>"11111101",
  47922=>"00000010",
  47923=>"11111101",
  47924=>"00000000",
  47925=>"11111110",
  47926=>"11111101",
  47927=>"11111110",
  47928=>"11111101",
  47929=>"00000010",
  47930=>"00000010",
  47931=>"00000001",
  47932=>"00000010",
  47933=>"00000100",
  47934=>"00000010",
  47935=>"00000000",
  47936=>"11111110",
  47937=>"11111110",
  47938=>"11111111",
  47939=>"00000010",
  47940=>"00000001",
  47941=>"00000001",
  47942=>"11111110",
  47943=>"11111111",
  47944=>"00000101",
  47945=>"11111111",
  47946=>"11111111",
  47947=>"00000011",
  47948=>"00000000",
  47949=>"00000001",
  47950=>"11111111",
  47951=>"11111110",
  47952=>"00000001",
  47953=>"00000011",
  47954=>"11111110",
  47955=>"11111101",
  47956=>"00000000",
  47957=>"11111110",
  47958=>"00000000",
  47959=>"00000001",
  47960=>"11111101",
  47961=>"11111101",
  47962=>"11111110",
  47963=>"00000011",
  47964=>"11111101",
  47965=>"00000101",
  47966=>"11111101",
  47967=>"11111110",
  47968=>"11111110",
  47969=>"00000101",
  47970=>"00000010",
  47971=>"11111101",
  47972=>"00000001",
  47973=>"11111110",
  47974=>"11111111",
  47975=>"11111111",
  47976=>"00000001",
  47977=>"00000011",
  47978=>"00000000",
  47979=>"00000000",
  47980=>"00000000",
  47981=>"00000001",
  47982=>"00000000",
  47983=>"11111100",
  47984=>"00000000",
  47985=>"00000001",
  47986=>"11111110",
  47987=>"11111101",
  47988=>"00000101",
  47989=>"11111111",
  47990=>"11111111",
  47991=>"00000010",
  47992=>"11111111",
  47993=>"00000010",
  47994=>"00000011",
  47995=>"00000000",
  47996=>"00000110",
  47997=>"11111101",
  47998=>"00000111",
  47999=>"11111100",
  48000=>"00000010",
  48001=>"00000110",
  48002=>"11111110",
  48003=>"11111111",
  48004=>"11111101",
  48005=>"00000000",
  48006=>"00000011",
  48007=>"11111100",
  48008=>"11111110",
  48009=>"11111101",
  48010=>"00000000",
  48011=>"00000011",
  48012=>"11111100",
  48013=>"00000101",
  48014=>"00000011",
  48015=>"00000001",
  48016=>"00000000",
  48017=>"00000010",
  48018=>"00000010",
  48019=>"11111111",
  48020=>"11111111",
  48021=>"11111110",
  48022=>"11111111",
  48023=>"00000011",
  48024=>"11111101",
  48025=>"11111100",
  48026=>"00000000",
  48027=>"11111011",
  48028=>"11111100",
  48029=>"11111111",
  48030=>"11111100",
  48031=>"11111101",
  48032=>"11111111",
  48033=>"11111111",
  48034=>"11111111",
  48035=>"00000001",
  48036=>"00000011",
  48037=>"11111111",
  48038=>"00000001",
  48039=>"11111100",
  48040=>"00000000",
  48041=>"11111101",
  48042=>"00000001",
  48043=>"00000001",
  48044=>"00000010",
  48045=>"00000001",
  48046=>"11111110",
  48047=>"11111110",
  48048=>"00000000",
  48049=>"11111011",
  48050=>"00000101",
  48051=>"00000100",
  48052=>"00000000",
  48053=>"00000011",
  48054=>"00000010",
  48055=>"00000000",
  48056=>"00000000",
  48057=>"00000000",
  48058=>"00000000",
  48059=>"11111101",
  48060=>"11111100",
  48061=>"00000010",
  48062=>"11111101",
  48063=>"00000000",
  48064=>"00000101",
  48065=>"00000001",
  48066=>"11111101",
  48067=>"00000000",
  48068=>"11111110",
  48069=>"00000001",
  48070=>"00000000",
  48071=>"00000001",
  48072=>"00000001",
  48073=>"11111111",
  48074=>"11111101",
  48075=>"11111111",
  48076=>"11111101",
  48077=>"11111111",
  48078=>"00000101",
  48079=>"00000001",
  48080=>"00000000",
  48081=>"11111110",
  48082=>"00000000",
  48083=>"00000000",
  48084=>"11111110",
  48085=>"00000001",
  48086=>"00000001",
  48087=>"11111110",
  48088=>"11111110",
  48089=>"11111111",
  48090=>"11111110",
  48091=>"11111101",
  48092=>"11111110",
  48093=>"11111110",
  48094=>"00000001",
  48095=>"00000001",
  48096=>"00000001",
  48097=>"00000001",
  48098=>"00000011",
  48099=>"00000011",
  48100=>"00000001",
  48101=>"11111111",
  48102=>"11111110",
  48103=>"00000000",
  48104=>"11111110",
  48105=>"00000001",
  48106=>"11111101",
  48107=>"11111101",
  48108=>"11111110",
  48109=>"00000101",
  48110=>"11111101",
  48111=>"00000011",
  48112=>"11111110",
  48113=>"00000010",
  48114=>"00000010",
  48115=>"11111111",
  48116=>"11111111",
  48117=>"00000110",
  48118=>"11111111",
  48119=>"00000000",
  48120=>"11111101",
  48121=>"00000001",
  48122=>"00000000",
  48123=>"00000001",
  48124=>"00000001",
  48125=>"11111111",
  48126=>"00000001",
  48127=>"00000001",
  48128=>"11111100",
  48129=>"00000100",
  48130=>"11111111",
  48131=>"00000000",
  48132=>"11111111",
  48133=>"00000011",
  48134=>"11111101",
  48135=>"00000100",
  48136=>"11111111",
  48137=>"11111100",
  48138=>"11111110",
  48139=>"00000001",
  48140=>"00000010",
  48141=>"11111111",
  48142=>"00000000",
  48143=>"11111110",
  48144=>"11111101",
  48145=>"00000000",
  48146=>"00000000",
  48147=>"11111110",
  48148=>"11111110",
  48149=>"11111110",
  48150=>"00000010",
  48151=>"00000001",
  48152=>"00000010",
  48153=>"00000000",
  48154=>"00000001",
  48155=>"00000000",
  48156=>"00000001",
  48157=>"11111101",
  48158=>"11111110",
  48159=>"00000011",
  48160=>"11111101",
  48161=>"00000000",
  48162=>"11111111",
  48163=>"00000001",
  48164=>"00000000",
  48165=>"11111111",
  48166=>"11111110",
  48167=>"11111111",
  48168=>"11111111",
  48169=>"00000000",
  48170=>"11111110",
  48171=>"11111111",
  48172=>"00000010",
  48173=>"00000000",
  48174=>"00000001",
  48175=>"00000001",
  48176=>"11111111",
  48177=>"11111111",
  48178=>"11111110",
  48179=>"00000001",
  48180=>"00000000",
  48181=>"11111101",
  48182=>"11111111",
  48183=>"11111110",
  48184=>"11111111",
  48185=>"11111110",
  48186=>"00000010",
  48187=>"11111110",
  48188=>"00000000",
  48189=>"00000001",
  48190=>"11111111",
  48191=>"00000000",
  48192=>"11111111",
  48193=>"00000000",
  48194=>"11111110",
  48195=>"00000001",
  48196=>"11111100",
  48197=>"00000001",
  48198=>"11111101",
  48199=>"00000001",
  48200=>"00000011",
  48201=>"11111110",
  48202=>"11111100",
  48203=>"00000001",
  48204=>"00000100",
  48205=>"00000001",
  48206=>"11111111",
  48207=>"11111110",
  48208=>"11111111",
  48209=>"00000010",
  48210=>"00000011",
  48211=>"00000000",
  48212=>"00000001",
  48213=>"11111101",
  48214=>"00000010",
  48215=>"00000000",
  48216=>"00000010",
  48217=>"11111111",
  48218=>"00000011",
  48219=>"11111101",
  48220=>"11111111",
  48221=>"11111101",
  48222=>"00000000",
  48223=>"00000101",
  48224=>"00000010",
  48225=>"00000001",
  48226=>"00000110",
  48227=>"00000011",
  48228=>"11111100",
  48229=>"11111101",
  48230=>"00000000",
  48231=>"11111111",
  48232=>"11111110",
  48233=>"11111111",
  48234=>"00000010",
  48235=>"11111110",
  48236=>"00000000",
  48237=>"11111101",
  48238=>"00000000",
  48239=>"11111110",
  48240=>"00000001",
  48241=>"11111111",
  48242=>"11111101",
  48243=>"00000001",
  48244=>"00000000",
  48245=>"11111100",
  48246=>"11111101",
  48247=>"11111110",
  48248=>"00000001",
  48249=>"11111100",
  48250=>"11111110",
  48251=>"11111110",
  48252=>"11111101",
  48253=>"11111101",
  48254=>"11111111",
  48255=>"11111101",
  48256=>"00000001",
  48257=>"11111110",
  48258=>"11111100",
  48259=>"11111101",
  48260=>"11111110",
  48261=>"11111111",
  48262=>"11111111",
  48263=>"00000000",
  48264=>"11111101",
  48265=>"11111110",
  48266=>"00000001",
  48267=>"11111110",
  48268=>"00000000",
  48269=>"11111111",
  48270=>"00000011",
  48271=>"00000000",
  48272=>"00000010",
  48273=>"11111101",
  48274=>"00000011",
  48275=>"11111111",
  48276=>"11111100",
  48277=>"11111100",
  48278=>"00000010",
  48279=>"00000010",
  48280=>"11111100",
  48281=>"11111101",
  48282=>"11111111",
  48283=>"00000000",
  48284=>"11111111",
  48285=>"00000000",
  48286=>"00000000",
  48287=>"11111100",
  48288=>"00000111",
  48289=>"11111110",
  48290=>"11111110",
  48291=>"11111111",
  48292=>"11111110",
  48293=>"11111111",
  48294=>"00000110",
  48295=>"11111110",
  48296=>"00000010",
  48297=>"11111111",
  48298=>"00000010",
  48299=>"11111100",
  48300=>"00000011",
  48301=>"00000001",
  48302=>"11111110",
  48303=>"00000010",
  48304=>"00000001",
  48305=>"11111111",
  48306=>"11111110",
  48307=>"00000101",
  48308=>"11111111",
  48309=>"11111100",
  48310=>"00000101",
  48311=>"11111110",
  48312=>"11111110",
  48313=>"11111101",
  48314=>"00000010",
  48315=>"00000000",
  48316=>"00000011",
  48317=>"00000000",
  48318=>"00000010",
  48319=>"00000010",
  48320=>"00000010",
  48321=>"00000010",
  48322=>"11111101",
  48323=>"11111101",
  48324=>"11111111",
  48325=>"00000011",
  48326=>"00000000",
  48327=>"00000011",
  48328=>"00000000",
  48329=>"11111101",
  48330=>"00000011",
  48331=>"11111110",
  48332=>"00000011",
  48333=>"00000000",
  48334=>"11111111",
  48335=>"00000101",
  48336=>"00000011",
  48337=>"00000001",
  48338=>"00000001",
  48339=>"11111110",
  48340=>"00000001",
  48341=>"11111111",
  48342=>"00000001",
  48343=>"00000010",
  48344=>"00000001",
  48345=>"00000001",
  48346=>"11111111",
  48347=>"11111111",
  48348=>"11111101",
  48349=>"00000100",
  48350=>"00000000",
  48351=>"00001001",
  48352=>"00000001",
  48353=>"00000000",
  48354=>"11111101",
  48355=>"00000011",
  48356=>"11111111",
  48357=>"00000010",
  48358=>"00000001",
  48359=>"00000011",
  48360=>"00000001",
  48361=>"00000011",
  48362=>"00000000",
  48363=>"00000010",
  48364=>"11111110",
  48365=>"00000001",
  48366=>"00000000",
  48367=>"00000010",
  48368=>"11111111",
  48369=>"11111101",
  48370=>"00000010",
  48371=>"00000011",
  48372=>"00000010",
  48373=>"11111111",
  48374=>"00000001",
  48375=>"11111111",
  48376=>"11111110",
  48377=>"00000011",
  48378=>"11111101",
  48379=>"00000000",
  48380=>"00000000",
  48381=>"00000011",
  48382=>"11111111",
  48383=>"11111101",
  48384=>"11111110",
  48385=>"11111111",
  48386=>"11111100",
  48387=>"00000001",
  48388=>"11111110",
  48389=>"00000110",
  48390=>"00000001",
  48391=>"00000011",
  48392=>"00000001",
  48393=>"11111101",
  48394=>"00000000",
  48395=>"00000100",
  48396=>"00000010",
  48397=>"11111111",
  48398=>"00000010",
  48399=>"11111101",
  48400=>"11111111",
  48401=>"00001000",
  48402=>"00000101",
  48403=>"11111100",
  48404=>"00000011",
  48405=>"00000000",
  48406=>"11111111",
  48407=>"00000110",
  48408=>"11111101",
  48409=>"00000000",
  48410=>"11111110",
  48411=>"00000001",
  48412=>"11111110",
  48413=>"00000000",
  48414=>"00000100",
  48415=>"00000000",
  48416=>"11111101",
  48417=>"00000011",
  48418=>"11111101",
  48419=>"11111101",
  48420=>"00000000",
  48421=>"00000010",
  48422=>"11111101",
  48423=>"00000010",
  48424=>"00000000",
  48425=>"00000001",
  48426=>"00000001",
  48427=>"11111111",
  48428=>"00000011",
  48429=>"00000000",
  48430=>"00000001",
  48431=>"11111110",
  48432=>"11111110",
  48433=>"11111111",
  48434=>"11111110",
  48435=>"00000010",
  48436=>"00000100",
  48437=>"00000010",
  48438=>"00000010",
  48439=>"11111110",
  48440=>"00000000",
  48441=>"11111100",
  48442=>"00000001",
  48443=>"00000011",
  48444=>"00000001",
  48445=>"00000000",
  48446=>"11111111",
  48447=>"00000011",
  48448=>"00000000",
  48449=>"00000000",
  48450=>"11111101",
  48451=>"11111110",
  48452=>"00000000",
  48453=>"11111101",
  48454=>"00000100",
  48455=>"11111111",
  48456=>"11111101",
  48457=>"11111110",
  48458=>"00000111",
  48459=>"11111101",
  48460=>"11111100",
  48461=>"00000010",
  48462=>"11111111",
  48463=>"11111110",
  48464=>"11111110",
  48465=>"00000000",
  48466=>"11111111",
  48467=>"11111101",
  48468=>"00000001",
  48469=>"11111100",
  48470=>"11111101",
  48471=>"11111101",
  48472=>"11111110",
  48473=>"00000011",
  48474=>"11111110",
  48475=>"00000111",
  48476=>"11111111",
  48477=>"00000000",
  48478=>"00000010",
  48479=>"00000010",
  48480=>"11111101",
  48481=>"00000001",
  48482=>"11111110",
  48483=>"00000001",
  48484=>"11111110",
  48485=>"11111101",
  48486=>"00000010",
  48487=>"11111110",
  48488=>"00000011",
  48489=>"00000011",
  48490=>"11111101",
  48491=>"00000010",
  48492=>"00000000",
  48493=>"00000000",
  48494=>"11111111",
  48495=>"00000010",
  48496=>"11111111",
  48497=>"00000000",
  48498=>"00000100",
  48499=>"00000011",
  48500=>"00000000",
  48501=>"11111101",
  48502=>"11111101",
  48503=>"00000001",
  48504=>"11111110",
  48505=>"11111100",
  48506=>"11111111",
  48507=>"00000001",
  48508=>"00000001",
  48509=>"00000000",
  48510=>"11111111",
  48511=>"00000001",
  48512=>"11111111",
  48513=>"00000011",
  48514=>"11111111",
  48515=>"00000001",
  48516=>"00000001",
  48517=>"11111110",
  48518=>"00000001",
  48519=>"00000010",
  48520=>"11111110",
  48521=>"11111100",
  48522=>"11111110",
  48523=>"00000001",
  48524=>"00000000",
  48525=>"00000000",
  48526=>"11111111",
  48527=>"00000101",
  48528=>"00000010",
  48529=>"11111111",
  48530=>"00000010",
  48531=>"11111111",
  48532=>"00000010",
  48533=>"00000110",
  48534=>"11111110",
  48535=>"00000001",
  48536=>"11111011",
  48537=>"00000101",
  48538=>"00000000",
  48539=>"00000010",
  48540=>"00000000",
  48541=>"11111100",
  48542=>"11111111",
  48543=>"11111100",
  48544=>"00000011",
  48545=>"11111100",
  48546=>"00000001",
  48547=>"00000100",
  48548=>"11111110",
  48549=>"00000001",
  48550=>"11111111",
  48551=>"11111111",
  48552=>"00000000",
  48553=>"00000000",
  48554=>"11111101",
  48555=>"11111100",
  48556=>"00000010",
  48557=>"00000000",
  48558=>"11111100",
  48559=>"00000110",
  48560=>"11111110",
  48561=>"00000001",
  48562=>"11111101",
  48563=>"00000011",
  48564=>"00000011",
  48565=>"11111110",
  48566=>"00000010",
  48567=>"00000010",
  48568=>"11111110",
  48569=>"11111111",
  48570=>"00000000",
  48571=>"00000011",
  48572=>"00000000",
  48573=>"11111101",
  48574=>"00000001",
  48575=>"11111111",
  48576=>"11111100",
  48577=>"00000010",
  48578=>"11111101",
  48579=>"11111110",
  48580=>"11111100",
  48581=>"00000001",
  48582=>"00000101",
  48583=>"00000000",
  48584=>"11111101",
  48585=>"11111101",
  48586=>"00000100",
  48587=>"00000100",
  48588=>"00000001",
  48589=>"00000010",
  48590=>"00000001",
  48591=>"00000011",
  48592=>"00000001",
  48593=>"00000001",
  48594=>"00000010",
  48595=>"11111111",
  48596=>"11111110",
  48597=>"11111111",
  48598=>"11111101",
  48599=>"00000000",
  48600=>"00000001",
  48601=>"00000001",
  48602=>"11111110",
  48603=>"11111110",
  48604=>"00000101",
  48605=>"11111110",
  48606=>"00000000",
  48607=>"11111011",
  48608=>"00000100",
  48609=>"00000100",
  48610=>"11111111",
  48611=>"11111101",
  48612=>"11111110",
  48613=>"11111101",
  48614=>"00000011",
  48615=>"11111111",
  48616=>"11111110",
  48617=>"00000001",
  48618=>"11111110",
  48619=>"11111100",
  48620=>"11111111",
  48621=>"11111101",
  48622=>"11111101",
  48623=>"11111110",
  48624=>"00000010",
  48625=>"00000011",
  48626=>"00000001",
  48627=>"00000100",
  48628=>"11111111",
  48629=>"00000010",
  48630=>"11111111",
  48631=>"11111110",
  48632=>"11111111",
  48633=>"00000010",
  48634=>"11111110",
  48635=>"11111110",
  48636=>"11111101",
  48637=>"00000100",
  48638=>"11111111",
  48639=>"11111101",
  48640=>"00000001",
  48641=>"00000101",
  48642=>"11111100",
  48643=>"11111101",
  48644=>"11111110",
  48645=>"00000010",
  48646=>"11111110",
  48647=>"00000001",
  48648=>"11111111",
  48649=>"00000100",
  48650=>"00000001",
  48651=>"00000010",
  48652=>"00000011",
  48653=>"00000010",
  48654=>"11111100",
  48655=>"00000000",
  48656=>"00000000",
  48657=>"00000000",
  48658=>"00000001",
  48659=>"00000011",
  48660=>"00000001",
  48661=>"11111110",
  48662=>"11111101",
  48663=>"11111101",
  48664=>"00000010",
  48665=>"00000000",
  48666=>"11111111",
  48667=>"11111100",
  48668=>"11111111",
  48669=>"00000010",
  48670=>"11111110",
  48671=>"11111100",
  48672=>"00000001",
  48673=>"11111101",
  48674=>"11111101",
  48675=>"11111101",
  48676=>"00000100",
  48677=>"00000000",
  48678=>"00000001",
  48679=>"11111101",
  48680=>"11111110",
  48681=>"11111111",
  48682=>"11111100",
  48683=>"00000010",
  48684=>"00000000",
  48685=>"11111110",
  48686=>"11111111",
  48687=>"00000010",
  48688=>"00000100",
  48689=>"11111101",
  48690=>"00000010",
  48691=>"11111110",
  48692=>"11111110",
  48693=>"00000110",
  48694=>"11111111",
  48695=>"11111101",
  48696=>"11111110",
  48697=>"00000010",
  48698=>"11111110",
  48699=>"00000000",
  48700=>"00000000",
  48701=>"11111101",
  48702=>"00000011",
  48703=>"11111111",
  48704=>"11111110",
  48705=>"00000001",
  48706=>"11111111",
  48707=>"11111101",
  48708=>"11111111",
  48709=>"11111111",
  48710=>"11111111",
  48711=>"00000000",
  48712=>"00000001",
  48713=>"00000000",
  48714=>"00000100",
  48715=>"11111110",
  48716=>"00000011",
  48717=>"11111111",
  48718=>"11111110",
  48719=>"00000001",
  48720=>"11111111",
  48721=>"11111110",
  48722=>"00000010",
  48723=>"00000001",
  48724=>"11111101",
  48725=>"11111100",
  48726=>"00000000",
  48727=>"11111111",
  48728=>"11111100",
  48729=>"00000000",
  48730=>"11111110",
  48731=>"00000001",
  48732=>"00000100",
  48733=>"11111101",
  48734=>"11111111",
  48735=>"11111101",
  48736=>"00000010",
  48737=>"00000010",
  48738=>"11111110",
  48739=>"11111110",
  48740=>"11111111",
  48741=>"00000000",
  48742=>"11111101",
  48743=>"11111100",
  48744=>"11111111",
  48745=>"00000001",
  48746=>"11111110",
  48747=>"00000011",
  48748=>"00000000",
  48749=>"11111110",
  48750=>"00000000",
  48751=>"11111101",
  48752=>"11111110",
  48753=>"11111111",
  48754=>"11111111",
  48755=>"00000010",
  48756=>"00000000",
  48757=>"00000100",
  48758=>"00000101",
  48759=>"00000001",
  48760=>"00000010",
  48761=>"11111111",
  48762=>"11111110",
  48763=>"11111111",
  48764=>"11111110",
  48765=>"00000001",
  48766=>"00000000",
  48767=>"11111110",
  48768=>"00000000",
  48769=>"00000001",
  48770=>"00000010",
  48771=>"00000011",
  48772=>"11111111",
  48773=>"00000000",
  48774=>"00000010",
  48775=>"00000000",
  48776=>"11111101",
  48777=>"11111101",
  48778=>"00000010",
  48779=>"11111100",
  48780=>"11111111",
  48781=>"11111110",
  48782=>"11111101",
  48783=>"00000010",
  48784=>"00000000",
  48785=>"00000001",
  48786=>"11111111",
  48787=>"00000010",
  48788=>"00000000",
  48789=>"00000000",
  48790=>"11111111",
  48791=>"11111100",
  48792=>"00000000",
  48793=>"00000010",
  48794=>"11111111",
  48795=>"00000100",
  48796=>"11111111",
  48797=>"00000110",
  48798=>"11111101",
  48799=>"11111101",
  48800=>"00000000",
  48801=>"00000000",
  48802=>"11111100",
  48803=>"11111100",
  48804=>"11111111",
  48805=>"00000011",
  48806=>"00000001",
  48807=>"00000000",
  48808=>"11111101",
  48809=>"11111110",
  48810=>"00000010",
  48811=>"00000000",
  48812=>"11111110",
  48813=>"00000000",
  48814=>"11111111",
  48815=>"00000001",
  48816=>"11111110",
  48817=>"00000010",
  48818=>"00000000",
  48819=>"00000000",
  48820=>"11111110",
  48821=>"00000100",
  48822=>"00000001",
  48823=>"00000101",
  48824=>"00000010",
  48825=>"11111110",
  48826=>"00000010",
  48827=>"11111110",
  48828=>"11111101",
  48829=>"00000010",
  48830=>"11111110",
  48831=>"00000000",
  48832=>"00000000",
  48833=>"11111111",
  48834=>"11111111",
  48835=>"11111100",
  48836=>"11111110",
  48837=>"11111110",
  48838=>"00000001",
  48839=>"11111111",
  48840=>"11111111",
  48841=>"11111110",
  48842=>"00000001",
  48843=>"00000011",
  48844=>"11111101",
  48845=>"11111110",
  48846=>"11111110",
  48847=>"11111101",
  48848=>"11111111",
  48849=>"00000001",
  48850=>"00000100",
  48851=>"00000001",
  48852=>"00000000",
  48853=>"00000010",
  48854=>"11111111",
  48855=>"11111110",
  48856=>"00000010",
  48857=>"11111110",
  48858=>"00000000",
  48859=>"00000011",
  48860=>"11111100",
  48861=>"00000011",
  48862=>"00000001",
  48863=>"00000011",
  48864=>"11111110",
  48865=>"11111101",
  48866=>"00000001",
  48867=>"00000001",
  48868=>"11111111",
  48869=>"11111110",
  48870=>"00000011",
  48871=>"00000001",
  48872=>"00000001",
  48873=>"00000011",
  48874=>"00000010",
  48875=>"00000001",
  48876=>"11111101",
  48877=>"11111101",
  48878=>"00000010",
  48879=>"11111110",
  48880=>"00000100",
  48881=>"00000010",
  48882=>"00000010",
  48883=>"00000000",
  48884=>"00000010",
  48885=>"00000001",
  48886=>"00000001",
  48887=>"00000001",
  48888=>"00000100",
  48889=>"11111110",
  48890=>"00000000",
  48891=>"00000101",
  48892=>"11111111",
  48893=>"11111100",
  48894=>"00000110",
  48895=>"00000001",
  48896=>"11111101",
  48897=>"11111110",
  48898=>"11111101",
  48899=>"00000000",
  48900=>"00000010",
  48901=>"11111101",
  48902=>"11111110",
  48903=>"00000001",
  48904=>"00001011",
  48905=>"00000110",
  48906=>"11111110",
  48907=>"00000010",
  48908=>"11111100",
  48909=>"11111110",
  48910=>"11111101",
  48911=>"00000010",
  48912=>"11111101",
  48913=>"00000000",
  48914=>"00000000",
  48915=>"00000011",
  48916=>"00000000",
  48917=>"11111110",
  48918=>"11111111",
  48919=>"00000010",
  48920=>"00000001",
  48921=>"11111100",
  48922=>"00000010",
  48923=>"11111011",
  48924=>"11111101",
  48925=>"11111110",
  48926=>"00000100",
  48927=>"11111110",
  48928=>"00000001",
  48929=>"00000010",
  48930=>"00000010",
  48931=>"11111110",
  48932=>"00000011",
  48933=>"11111101",
  48934=>"00000010",
  48935=>"00000110",
  48936=>"11111110",
  48937=>"11111101",
  48938=>"00000010",
  48939=>"11111110",
  48940=>"11111110",
  48941=>"11111101",
  48942=>"11111100",
  48943=>"11111111",
  48944=>"00000010",
  48945=>"00000001",
  48946=>"11111101",
  48947=>"00000001",
  48948=>"00000001",
  48949=>"00000000",
  48950=>"11111101",
  48951=>"11111111",
  48952=>"00000000",
  48953=>"00000001",
  48954=>"11111111",
  48955=>"00000001",
  48956=>"11111110",
  48957=>"11111101",
  48958=>"11111110",
  48959=>"00000011",
  48960=>"00000011",
  48961=>"11111101",
  48962=>"11111110",
  48963=>"00000010",
  48964=>"11111110",
  48965=>"11111110",
  48966=>"00000100",
  48967=>"11111110",
  48968=>"00000000",
  48969=>"00000001",
  48970=>"11111111",
  48971=>"11111111",
  48972=>"00000010",
  48973=>"00000000",
  48974=>"00000010",
  48975=>"00000000",
  48976=>"00000011",
  48977=>"11111101",
  48978=>"11111101",
  48979=>"11111111",
  48980=>"00000010",
  48981=>"11111111",
  48982=>"00000011",
  48983=>"11111111",
  48984=>"11111100",
  48985=>"11111110",
  48986=>"11111110",
  48987=>"11111101",
  48988=>"11111111",
  48989=>"00000000",
  48990=>"11111100",
  48991=>"11111111",
  48992=>"00000001",
  48993=>"11111111",
  48994=>"11111110",
  48995=>"00000010",
  48996=>"00000001",
  48997=>"11111110",
  48998=>"11111101",
  48999=>"11111011",
  49000=>"00000010",
  49001=>"11111111",
  49002=>"00000001",
  49003=>"00000001",
  49004=>"11111101",
  49005=>"11111111",
  49006=>"11111110",
  49007=>"00000010",
  49008=>"00000001",
  49009=>"00000001",
  49010=>"00000000",
  49011=>"11111110",
  49012=>"00000010",
  49013=>"11111111",
  49014=>"00000010",
  49015=>"00000010",
  49016=>"00000010",
  49017=>"11111101",
  49018=>"11111100",
  49019=>"11111111",
  49020=>"00000000",
  49021=>"11111101",
  49022=>"00000000",
  49023=>"11111110",
  49024=>"00000000",
  49025=>"00000010",
  49026=>"11111101",
  49027=>"11111100",
  49028=>"11111101",
  49029=>"11111101",
  49030=>"11111100",
  49031=>"11111101",
  49032=>"00000010",
  49033=>"11111111",
  49034=>"00000011",
  49035=>"00000010",
  49036=>"11111101",
  49037=>"11111101",
  49038=>"00000001",
  49039=>"00000010",
  49040=>"00000000",
  49041=>"00000000",
  49042=>"11111011",
  49043=>"11111111",
  49044=>"00000101",
  49045=>"00001000",
  49046=>"11111110",
  49047=>"00000000",
  49048=>"11111100",
  49049=>"11111110",
  49050=>"00000110",
  49051=>"00000000",
  49052=>"11111110",
  49053=>"00000010",
  49054=>"00000000",
  49055=>"00000010",
  49056=>"00000011",
  49057=>"00000011",
  49058=>"00000010",
  49059=>"00000001",
  49060=>"11111110",
  49061=>"00000001",
  49062=>"00000011",
  49063=>"00000101",
  49064=>"11111111",
  49065=>"00000001",
  49066=>"00000010",
  49067=>"00000010",
  49068=>"00000001",
  49069=>"11111111",
  49070=>"11111111",
  49071=>"00000000",
  49072=>"00000001",
  49073=>"00000001",
  49074=>"11111111",
  49075=>"00000001",
  49076=>"00000000",
  49077=>"00000010",
  49078=>"11111101",
  49079=>"00000001",
  49080=>"00000100",
  49081=>"11111101",
  49082=>"11111111",
  49083=>"11111101",
  49084=>"00000001",
  49085=>"11111110",
  49086=>"00000010",
  49087=>"11111110",
  49088=>"11111110",
  49089=>"00000010",
  49090=>"00000010",
  49091=>"11111111",
  49092=>"00000000",
  49093=>"00000001",
  49094=>"11111110",
  49095=>"11111110",
  49096=>"11111110",
  49097=>"00000101",
  49098=>"00000001",
  49099=>"00000011",
  49100=>"11111111",
  49101=>"11111110",
  49102=>"11111110",
  49103=>"11111100",
  49104=>"11111101",
  49105=>"00000001",
  49106=>"11111111",
  49107=>"00000011",
  49108=>"00000000",
  49109=>"00000001",
  49110=>"11111110",
  49111=>"11111111",
  49112=>"00000010",
  49113=>"11111111",
  49114=>"00000010",
  49115=>"11111111",
  49116=>"00000011",
  49117=>"11111111",
  49118=>"00000001",
  49119=>"11111101",
  49120=>"11111110",
  49121=>"00000001",
  49122=>"00000010",
  49123=>"00000010",
  49124=>"11111111",
  49125=>"00000010",
  49126=>"00000001",
  49127=>"00000001",
  49128=>"00000100",
  49129=>"00000000",
  49130=>"00000011",
  49131=>"11111101",
  49132=>"11111101",
  49133=>"00000001",
  49134=>"11111110",
  49135=>"11111100",
  49136=>"00000000",
  49137=>"00000000",
  49138=>"00000001",
  49139=>"11111100",
  49140=>"11111110",
  49141=>"00000100",
  49142=>"00000000",
  49143=>"11111011",
  49144=>"00000000",
  49145=>"11111101",
  49146=>"11111111",
  49147=>"11111110",
  49148=>"00000000",
  49149=>"11111101",
  49150=>"00000000",
  49151=>"00000011",
  49152=>"00000000",
  49153=>"11111101",
  49154=>"00000000",
  49155=>"00000011",
  49156=>"00000001",
  49157=>"00000000",
  49158=>"00000000",
  49159=>"00000000",
  49160=>"11111101",
  49161=>"11111101",
  49162=>"00000001",
  49163=>"11111111",
  49164=>"00000010",
  49165=>"00000000",
  49166=>"00000010",
  49167=>"11111111",
  49168=>"11111111",
  49169=>"11111101",
  49170=>"11111111",
  49171=>"00000100",
  49172=>"00000010",
  49173=>"11111110",
  49174=>"00000010",
  49175=>"11111111",
  49176=>"11111111",
  49177=>"11111110",
  49178=>"00000000",
  49179=>"00000000",
  49180=>"11111111",
  49181=>"11111101",
  49182=>"00000000",
  49183=>"11111100",
  49184=>"00000000",
  49185=>"11111100",
  49186=>"11111101",
  49187=>"11111100",
  49188=>"00000000",
  49189=>"00000000",
  49190=>"00000000",
  49191=>"00000000",
  49192=>"00000001",
  49193=>"11111101",
  49194=>"00000000",
  49195=>"11111111",
  49196=>"00000010",
  49197=>"11111110",
  49198=>"11111110",
  49199=>"11111110",
  49200=>"11111110",
  49201=>"00000001",
  49202=>"00000100",
  49203=>"00000010",
  49204=>"00000011",
  49205=>"00000001",
  49206=>"00000000",
  49207=>"11111110",
  49208=>"00000011",
  49209=>"11111101",
  49210=>"00000010",
  49211=>"11111111",
  49212=>"11111111",
  49213=>"00000000",
  49214=>"00000000",
  49215=>"11111111",
  49216=>"11111111",
  49217=>"00000000",
  49218=>"00000000",
  49219=>"00000001",
  49220=>"11111101",
  49221=>"11111110",
  49222=>"11111111",
  49223=>"00000110",
  49224=>"00000000",
  49225=>"11111110",
  49226=>"00000001",
  49227=>"11111110",
  49228=>"11111101",
  49229=>"00000011",
  49230=>"11111110",
  49231=>"11111110",
  49232=>"00000000",
  49233=>"11111101",
  49234=>"11111100",
  49235=>"11111111",
  49236=>"00000000",
  49237=>"00000000",
  49238=>"11111111",
  49239=>"11111111",
  49240=>"00000000",
  49241=>"11111110",
  49242=>"00000010",
  49243=>"00000010",
  49244=>"11111111",
  49245=>"11111111",
  49246=>"11111111",
  49247=>"11111100",
  49248=>"00000010",
  49249=>"00000001",
  49250=>"00000001",
  49251=>"00000101",
  49252=>"11111110",
  49253=>"11111111",
  49254=>"00000001",
  49255=>"11111110",
  49256=>"00000000",
  49257=>"11111111",
  49258=>"11111110",
  49259=>"11111111",
  49260=>"00000010",
  49261=>"00000100",
  49262=>"00000001",
  49263=>"11111110",
  49264=>"00000010",
  49265=>"00000010",
  49266=>"11111111",
  49267=>"00000001",
  49268=>"11111111",
  49269=>"00000000",
  49270=>"00000011",
  49271=>"11111101",
  49272=>"11111101",
  49273=>"00000000",
  49274=>"00000100",
  49275=>"00000000",
  49276=>"11111110",
  49277=>"11111110",
  49278=>"00000001",
  49279=>"00000011",
  49280=>"11111110",
  49281=>"00000000",
  49282=>"00000101",
  49283=>"11111101",
  49284=>"00000011",
  49285=>"00000000",
  49286=>"00000001",
  49287=>"00000000",
  49288=>"00000001",
  49289=>"11111110",
  49290=>"00000101",
  49291=>"00000001",
  49292=>"00000100",
  49293=>"00000001",
  49294=>"00000001",
  49295=>"00000000",
  49296=>"00000001",
  49297=>"11111101",
  49298=>"00000010",
  49299=>"11111111",
  49300=>"11111101",
  49301=>"00000010",
  49302=>"11111110",
  49303=>"11111110",
  49304=>"00000000",
  49305=>"11111101",
  49306=>"00000001",
  49307=>"00000000",
  49308=>"00000000",
  49309=>"11111111",
  49310=>"11111111",
  49311=>"00000011",
  49312=>"11111101",
  49313=>"11111101",
  49314=>"00000000",
  49315=>"11111100",
  49316=>"00000010",
  49317=>"11111110",
  49318=>"11111111",
  49319=>"00000000",
  49320=>"11111110",
  49321=>"11111110",
  49322=>"11111101",
  49323=>"11111111",
  49324=>"11111101",
  49325=>"00000011",
  49326=>"00000011",
  49327=>"00000010",
  49328=>"00000010",
  49329=>"00000000",
  49330=>"00000000",
  49331=>"11111110",
  49332=>"00000000",
  49333=>"11111111",
  49334=>"11111110",
  49335=>"00000111",
  49336=>"11111111",
  49337=>"11111101",
  49338=>"11111110",
  49339=>"00000001",
  49340=>"11111111",
  49341=>"00000001",
  49342=>"11111111",
  49343=>"00000001",
  49344=>"00000010",
  49345=>"11111101",
  49346=>"00000000",
  49347=>"00000010",
  49348=>"11111111",
  49349=>"00000100",
  49350=>"11111110",
  49351=>"00000001",
  49352=>"11111111",
  49353=>"11111110",
  49354=>"11111101",
  49355=>"00000000",
  49356=>"11111101",
  49357=>"00000001",
  49358=>"11111111",
  49359=>"11111101",
  49360=>"11111111",
  49361=>"11111111",
  49362=>"11111110",
  49363=>"00000001",
  49364=>"00000010",
  49365=>"00000000",
  49366=>"11111111",
  49367=>"11111110",
  49368=>"11111111",
  49369=>"00000001",
  49370=>"11111101",
  49371=>"00001000",
  49372=>"11111111",
  49373=>"11111110",
  49374=>"11111111",
  49375=>"11111111",
  49376=>"00000001",
  49377=>"00000101",
  49378=>"11111111",
  49379=>"11111101",
  49380=>"00000110",
  49381=>"11111111",
  49382=>"00000111",
  49383=>"11111110",
  49384=>"00000010",
  49385=>"11111101",
  49386=>"00000001",
  49387=>"11111101",
  49388=>"00000011",
  49389=>"11111110",
  49390=>"11111111",
  49391=>"00000000",
  49392=>"00000001",
  49393=>"11111110",
  49394=>"11111101",
  49395=>"11111111",
  49396=>"00000000",
  49397=>"11111111",
  49398=>"00000001",
  49399=>"00000011",
  49400=>"11111111",
  49401=>"00000001",
  49402=>"00000011",
  49403=>"00000001",
  49404=>"00000000",
  49405=>"11111100",
  49406=>"11111110",
  49407=>"00000010",
  49408=>"11111101",
  49409=>"11111111",
  49410=>"00000100",
  49411=>"00000100",
  49412=>"11111101",
  49413=>"00000010",
  49414=>"11111101",
  49415=>"00000011",
  49416=>"00000010",
  49417=>"11111101",
  49418=>"00000011",
  49419=>"00000001",
  49420=>"11111110",
  49421=>"11111100",
  49422=>"11111110",
  49423=>"00000011",
  49424=>"11111110",
  49425=>"11111101",
  49426=>"00000001",
  49427=>"00000010",
  49428=>"00000001",
  49429=>"11111101",
  49430=>"00000000",
  49431=>"11111101",
  49432=>"00000100",
  49433=>"11111110",
  49434=>"00000010",
  49435=>"11111111",
  49436=>"00000000",
  49437=>"00000010",
  49438=>"00000010",
  49439=>"11111110",
  49440=>"11111111",
  49441=>"00000001",
  49442=>"00000000",
  49443=>"00000000",
  49444=>"00000000",
  49445=>"00000001",
  49446=>"11111110",
  49447=>"11111110",
  49448=>"00000011",
  49449=>"11111110",
  49450=>"11111101",
  49451=>"00000100",
  49452=>"11111111",
  49453=>"11111111",
  49454=>"00000001",
  49455=>"00000001",
  49456=>"00000000",
  49457=>"11111110",
  49458=>"11111111",
  49459=>"11111111",
  49460=>"11111110",
  49461=>"11111101",
  49462=>"11111111",
  49463=>"11111111",
  49464=>"00000000",
  49465=>"11111101",
  49466=>"00000000",
  49467=>"00000001",
  49468=>"11111101",
  49469=>"00000010",
  49470=>"11111111",
  49471=>"00000000",
  49472=>"11111110",
  49473=>"00000000",
  49474=>"00000010",
  49475=>"00000001",
  49476=>"11111111",
  49477=>"11111101",
  49478=>"11111100",
  49479=>"11111101",
  49480=>"00000000",
  49481=>"11111110",
  49482=>"00000011",
  49483=>"00000001",
  49484=>"00000000",
  49485=>"00000010",
  49486=>"11111111",
  49487=>"11111101",
  49488=>"00000011",
  49489=>"00000011",
  49490=>"00000000",
  49491=>"11111110",
  49492=>"00000001",
  49493=>"00000010",
  49494=>"11111111",
  49495=>"11111110",
  49496=>"11111101",
  49497=>"11111101",
  49498=>"11111110",
  49499=>"11111110",
  49500=>"00000000",
  49501=>"00000000",
  49502=>"00000000",
  49503=>"00000011",
  49504=>"11111101",
  49505=>"11111111",
  49506=>"00000001",
  49507=>"00000001",
  49508=>"00000010",
  49509=>"00000001",
  49510=>"00000000",
  49511=>"11111111",
  49512=>"00000001",
  49513=>"11111111",
  49514=>"11111110",
  49515=>"11111111",
  49516=>"11111110",
  49517=>"00000010",
  49518=>"00000000",
  49519=>"00000011",
  49520=>"11111111",
  49521=>"11111110",
  49522=>"11111110",
  49523=>"11111110",
  49524=>"11111101",
  49525=>"00000000",
  49526=>"00000000",
  49527=>"11111111",
  49528=>"00000001",
  49529=>"00000010",
  49530=>"00000000",
  49531=>"11111111",
  49532=>"11111110",
  49533=>"11111110",
  49534=>"11111110",
  49535=>"11111111",
  49536=>"00000010",
  49537=>"00000001",
  49538=>"00000010",
  49539=>"00000001",
  49540=>"00000001",
  49541=>"00000000",
  49542=>"11111110",
  49543=>"11111110",
  49544=>"11111110",
  49545=>"11111110",
  49546=>"00000001",
  49547=>"11111111",
  49548=>"00000001",
  49549=>"11111111",
  49550=>"11111101",
  49551=>"11111110",
  49552=>"00000000",
  49553=>"11111110",
  49554=>"00000000",
  49555=>"00000001",
  49556=>"00000011",
  49557=>"11111101",
  49558=>"11111110",
  49559=>"00000000",
  49560=>"11111100",
  49561=>"00000011",
  49562=>"11111100",
  49563=>"11111101",
  49564=>"11111110",
  49565=>"11111110",
  49566=>"00000000",
  49567=>"11111110",
  49568=>"00000011",
  49569=>"00000001",
  49570=>"00000001",
  49571=>"11111101",
  49572=>"11111111",
  49573=>"11111101",
  49574=>"11111111",
  49575=>"11111110",
  49576=>"11111111",
  49577=>"11111101",
  49578=>"00000000",
  49579=>"11111101",
  49580=>"00000011",
  49581=>"00000110",
  49582=>"00000000",
  49583=>"11111101",
  49584=>"11111101",
  49585=>"00000011",
  49586=>"00000011",
  49587=>"11111101",
  49588=>"11111110",
  49589=>"11111101",
  49590=>"00000001",
  49591=>"11111101",
  49592=>"00000001",
  49593=>"00000001",
  49594=>"00000001",
  49595=>"11111100",
  49596=>"11111110",
  49597=>"11111101",
  49598=>"11111111",
  49599=>"00000011",
  49600=>"00000001",
  49601=>"11111101",
  49602=>"11111110",
  49603=>"11111100",
  49604=>"11111101",
  49605=>"00000001",
  49606=>"11111111",
  49607=>"11111111",
  49608=>"00000001",
  49609=>"11111101",
  49610=>"00000000",
  49611=>"11111110",
  49612=>"00000000",
  49613=>"11111101",
  49614=>"11111101",
  49615=>"00000101",
  49616=>"00000010",
  49617=>"00000100",
  49618=>"11111101",
  49619=>"11111110",
  49620=>"11111101",
  49621=>"00000100",
  49622=>"11111111",
  49623=>"00000011",
  49624=>"00000001",
  49625=>"00000001",
  49626=>"00000000",
  49627=>"00000011",
  49628=>"00000010",
  49629=>"11111101",
  49630=>"00000001",
  49631=>"00000001",
  49632=>"11111101",
  49633=>"11111100",
  49634=>"00000010",
  49635=>"11111111",
  49636=>"00000001",
  49637=>"11111110",
  49638=>"00000101",
  49639=>"00000000",
  49640=>"11111110",
  49641=>"00000000",
  49642=>"00000001",
  49643=>"11111110",
  49644=>"00000000",
  49645=>"00000001",
  49646=>"11111110",
  49647=>"11111111",
  49648=>"00000001",
  49649=>"11111111",
  49650=>"00000000",
  49651=>"00000101",
  49652=>"11111110",
  49653=>"00000011",
  49654=>"00000000",
  49655=>"11111110",
  49656=>"00000000",
  49657=>"00000010",
  49658=>"00000010",
  49659=>"00000000",
  49660=>"00000000",
  49661=>"00000100",
  49662=>"00000001",
  49663=>"00000010",
  49664=>"00000010",
  49665=>"11111110",
  49666=>"11111101",
  49667=>"11111111",
  49668=>"00000001",
  49669=>"00000010",
  49670=>"00000101",
  49671=>"11111101",
  49672=>"00000000",
  49673=>"11111111",
  49674=>"11111111",
  49675=>"11111101",
  49676=>"11111110",
  49677=>"00000000",
  49678=>"00000001",
  49679=>"11111101",
  49680=>"00000010",
  49681=>"11111111",
  49682=>"00000100",
  49683=>"11111101",
  49684=>"11111100",
  49685=>"00000000",
  49686=>"11111110",
  49687=>"00000001",
  49688=>"00000100",
  49689=>"00000010",
  49690=>"11111111",
  49691=>"11111110",
  49692=>"00000011",
  49693=>"00000001",
  49694=>"11111101",
  49695=>"11111111",
  49696=>"00000110",
  49697=>"11111110",
  49698=>"11111101",
  49699=>"00000000",
  49700=>"11111100",
  49701=>"00000110",
  49702=>"00000001",
  49703=>"00000010",
  49704=>"00000011",
  49705=>"00000011",
  49706=>"00000000",
  49707=>"00000010",
  49708=>"11111111",
  49709=>"11111110",
  49710=>"00000011",
  49711=>"11111101",
  49712=>"11111110",
  49713=>"00000010",
  49714=>"11111110",
  49715=>"11111110",
  49716=>"11111111",
  49717=>"11111101",
  49718=>"11111100",
  49719=>"11111101",
  49720=>"11111100",
  49721=>"11111110",
  49722=>"11111111",
  49723=>"00000010",
  49724=>"11111101",
  49725=>"11111111",
  49726=>"11111111",
  49727=>"11111101",
  49728=>"00000000",
  49729=>"11111101",
  49730=>"11111111",
  49731=>"00000001",
  49732=>"11111110",
  49733=>"11111110",
  49734=>"11111111",
  49735=>"00000100",
  49736=>"11111110",
  49737=>"11111110",
  49738=>"11111111",
  49739=>"00000000",
  49740=>"11111110",
  49741=>"11111111",
  49742=>"00000000",
  49743=>"00000001",
  49744=>"11111101",
  49745=>"00000001",
  49746=>"00000011",
  49747=>"11111110",
  49748=>"11111100",
  49749=>"00000010",
  49750=>"11111110",
  49751=>"11111101",
  49752=>"11111111",
  49753=>"00000101",
  49754=>"00000010",
  49755=>"11111111",
  49756=>"11111101",
  49757=>"11111101",
  49758=>"00000000",
  49759=>"00000010",
  49760=>"00000000",
  49761=>"11111110",
  49762=>"00000000",
  49763=>"11111111",
  49764=>"11111111",
  49765=>"11111101",
  49766=>"11111110",
  49767=>"00000000",
  49768=>"11111110",
  49769=>"00000010",
  49770=>"11111101",
  49771=>"00000000",
  49772=>"11111110",
  49773=>"00000000",
  49774=>"11111111",
  49775=>"11111111",
  49776=>"00000010",
  49777=>"11111110",
  49778=>"00000000",
  49779=>"11111111",
  49780=>"11111110",
  49781=>"00000100",
  49782=>"00000000",
  49783=>"11111111",
  49784=>"00000001",
  49785=>"11111111",
  49786=>"00000100",
  49787=>"00000011",
  49788=>"00000000",
  49789=>"11111111",
  49790=>"00000000",
  49791=>"00000010",
  49792=>"00000000",
  49793=>"11111111",
  49794=>"11111110",
  49795=>"00000011",
  49796=>"00000010",
  49797=>"11111111",
  49798=>"11111111",
  49799=>"00000011",
  49800=>"11111101",
  49801=>"00000000",
  49802=>"00000000",
  49803=>"00000000",
  49804=>"11111110",
  49805=>"00000001",
  49806=>"00000011",
  49807=>"00000001",
  49808=>"00000011",
  49809=>"00000000",
  49810=>"11111111",
  49811=>"11111110",
  49812=>"11111111",
  49813=>"00000010",
  49814=>"00000001",
  49815=>"11111110",
  49816=>"00000000",
  49817=>"00000011",
  49818=>"00000010",
  49819=>"00000011",
  49820=>"11111100",
  49821=>"00000010",
  49822=>"00000000",
  49823=>"00000010",
  49824=>"11111101",
  49825=>"11111100",
  49826=>"00000011",
  49827=>"00000001",
  49828=>"11111111",
  49829=>"11111101",
  49830=>"11111111",
  49831=>"00000011",
  49832=>"00000001",
  49833=>"11111101",
  49834=>"11111110",
  49835=>"00000001",
  49836=>"00000000",
  49837=>"11111101",
  49838=>"11111111",
  49839=>"00000000",
  49840=>"00000000",
  49841=>"00000011",
  49842=>"00000010",
  49843=>"00000011",
  49844=>"00000010",
  49845=>"00000001",
  49846=>"11111110",
  49847=>"11111101",
  49848=>"00000000",
  49849=>"11111101",
  49850=>"11111101",
  49851=>"00000011",
  49852=>"00000010",
  49853=>"00000001",
  49854=>"11111101",
  49855=>"00000010",
  49856=>"00000100",
  49857=>"00000010",
  49858=>"00000000",
  49859=>"00000001",
  49860=>"00000011",
  49861=>"11111100",
  49862=>"11111101",
  49863=>"11111111",
  49864=>"11111101",
  49865=>"00000000",
  49866=>"11111110",
  49867=>"00000010",
  49868=>"11111110",
  49869=>"00000001",
  49870=>"00000000",
  49871=>"00000010",
  49872=>"00000000",
  49873=>"11111111",
  49874=>"00000000",
  49875=>"11111110",
  49876=>"11111110",
  49877=>"00000010",
  49878=>"00000000",
  49879=>"00000001",
  49880=>"11111101",
  49881=>"00000001",
  49882=>"11111110",
  49883=>"00000011",
  49884=>"11111111",
  49885=>"11111110",
  49886=>"00000100",
  49887=>"11111101",
  49888=>"11111110",
  49889=>"11111111",
  49890=>"00000011",
  49891=>"11111101",
  49892=>"11111110",
  49893=>"00000011",
  49894=>"11111111",
  49895=>"11111111",
  49896=>"11111110",
  49897=>"00000010",
  49898=>"11111110",
  49899=>"11111111",
  49900=>"00000000",
  49901=>"00000011",
  49902=>"00000000",
  49903=>"11111110",
  49904=>"11111111",
  49905=>"11111101",
  49906=>"00000010",
  49907=>"00000010",
  49908=>"00000010",
  49909=>"11111101",
  49910=>"11111111",
  49911=>"00000011",
  49912=>"00000001",
  49913=>"00000010",
  49914=>"00000001",
  49915=>"11111101",
  49916=>"11111101",
  49917=>"00000011",
  49918=>"11111111",
  49919=>"11111110",
  49920=>"00000001",
  49921=>"11111100",
  49922=>"11111111",
  49923=>"11111111",
  49924=>"00000100",
  49925=>"00000001",
  49926=>"00000010",
  49927=>"00000001",
  49928=>"11111111",
  49929=>"11111101",
  49930=>"11111111",
  49931=>"11111110",
  49932=>"11111101",
  49933=>"00000010",
  49934=>"00000010",
  49935=>"00000001",
  49936=>"11111111",
  49937=>"00000010",
  49938=>"00000001",
  49939=>"11111111",
  49940=>"11111101",
  49941=>"11111101",
  49942=>"11111111",
  49943=>"00000001",
  49944=>"00000110",
  49945=>"11111111",
  49946=>"00000100",
  49947=>"11111101",
  49948=>"00000001",
  49949=>"11111111",
  49950=>"11111110",
  49951=>"00000001",
  49952=>"11111111",
  49953=>"00000010",
  49954=>"00000011",
  49955=>"11111110",
  49956=>"00000010",
  49957=>"00000010",
  49958=>"00000000",
  49959=>"11111111",
  49960=>"00000000",
  49961=>"00000010",
  49962=>"11111110",
  49963=>"00000001",
  49964=>"11111110",
  49965=>"00000001",
  49966=>"00000000",
  49967=>"00000001",
  49968=>"00000001",
  49969=>"11111100",
  49970=>"11111101",
  49971=>"00000001",
  49972=>"11111110",
  49973=>"00000101",
  49974=>"00000000",
  49975=>"11111101",
  49976=>"11111100",
  49977=>"00000000",
  49978=>"11111110",
  49979=>"00000001",
  49980=>"00000010",
  49981=>"11111111",
  49982=>"00000000",
  49983=>"11111111",
  49984=>"11111100",
  49985=>"00000000",
  49986=>"00000000",
  49987=>"00000000",
  49988=>"00000000",
  49989=>"11111111",
  49990=>"00000001",
  49991=>"11111110",
  49992=>"00000010",
  49993=>"11111110",
  49994=>"00000001",
  49995=>"00000010",
  49996=>"00000100",
  49997=>"11111111",
  49998=>"00000000",
  49999=>"00000001",
  50000=>"00000000",
  50001=>"00000001",
  50002=>"11111111",
  50003=>"00000001",
  50004=>"11111111",
  50005=>"11111110",
  50006=>"00000001",
  50007=>"11111111",
  50008=>"00000010",
  50009=>"00000010",
  50010=>"11111111",
  50011=>"11111111",
  50012=>"11111110",
  50013=>"00000010",
  50014=>"00000101",
  50015=>"11111110",
  50016=>"00000010",
  50017=>"00000001",
  50018=>"00000101",
  50019=>"00000000",
  50020=>"00000001",
  50021=>"11111111",
  50022=>"00000110",
  50023=>"00000010",
  50024=>"00000001",
  50025=>"00000110",
  50026=>"11111110",
  50027=>"11111111",
  50028=>"11111110",
  50029=>"00000000",
  50030=>"11111110",
  50031=>"00000000",
  50032=>"11111111",
  50033=>"00000001",
  50034=>"11111111",
  50035=>"00000101",
  50036=>"11111101",
  50037=>"00000100",
  50038=>"11111111",
  50039=>"00000001",
  50040=>"00000001",
  50041=>"00000001",
  50042=>"11111110",
  50043=>"00000010",
  50044=>"00000010",
  50045=>"11111111",
  50046=>"11111110",
  50047=>"11111111",
  50048=>"00000010",
  50049=>"00000010",
  50050=>"11111110",
  50051=>"11111111",
  50052=>"00000000",
  50053=>"11111110",
  50054=>"00000101",
  50055=>"11111110",
  50056=>"00000001",
  50057=>"11111101",
  50058=>"00000000",
  50059=>"11111110",
  50060=>"00000110",
  50061=>"00000010",
  50062=>"00000001",
  50063=>"11111111",
  50064=>"00000001",
  50065=>"11111100",
  50066=>"11111110",
  50067=>"00000010",
  50068=>"00000100",
  50069=>"00000001",
  50070=>"00000010",
  50071=>"00000001",
  50072=>"00000010",
  50073=>"00000001",
  50074=>"00000001",
  50075=>"11111101",
  50076=>"00000100",
  50077=>"00000001",
  50078=>"00000001",
  50079=>"00000001",
  50080=>"00000001",
  50081=>"00000001",
  50082=>"11111111",
  50083=>"11111110",
  50084=>"00000000",
  50085=>"11111111",
  50086=>"11111110",
  50087=>"00000000",
  50088=>"00000000",
  50089=>"00000010",
  50090=>"00000010",
  50091=>"00000001",
  50092=>"00000001",
  50093=>"11111111",
  50094=>"00000010",
  50095=>"00000000",
  50096=>"00000000",
  50097=>"11111111",
  50098=>"11111110",
  50099=>"11111111",
  50100=>"11111110",
  50101=>"00000001",
  50102=>"11111101",
  50103=>"00000000",
  50104=>"11111110",
  50105=>"00000010",
  50106=>"00000001",
  50107=>"11111110",
  50108=>"00000010",
  50109=>"11111110",
  50110=>"00000010",
  50111=>"00000000",
  50112=>"00000001",
  50113=>"00000010",
  50114=>"00000001",
  50115=>"00000000",
  50116=>"00000000",
  50117=>"11111101",
  50118=>"11111101",
  50119=>"11111110",
  50120=>"00000100",
  50121=>"00000100",
  50122=>"00000001",
  50123=>"00000100",
  50124=>"11111101",
  50125=>"00000100",
  50126=>"11111110",
  50127=>"00000000",
  50128=>"11111101",
  50129=>"11111111",
  50130=>"11111100",
  50131=>"11111110",
  50132=>"11111101",
  50133=>"11111101",
  50134=>"00000011",
  50135=>"00000000",
  50136=>"11111101",
  50137=>"00000010",
  50138=>"00000000",
  50139=>"00000100",
  50140=>"11111101",
  50141=>"11111111",
  50142=>"11111110",
  50143=>"11111100",
  50144=>"00000001",
  50145=>"00000100",
  50146=>"00000000",
  50147=>"00000000",
  50148=>"00000100",
  50149=>"00000001",
  50150=>"00000100",
  50151=>"00000001",
  50152=>"00000000",
  50153=>"11111111",
  50154=>"00000000",
  50155=>"00000001",
  50156=>"11111110",
  50157=>"00000001",
  50158=>"11111110",
  50159=>"11111111",
  50160=>"11111110",
  50161=>"11111111",
  50162=>"00000000",
  50163=>"11111101",
  50164=>"00000001",
  50165=>"00000010",
  50166=>"00000000",
  50167=>"00000000",
  50168=>"11111101",
  50169=>"11111110",
  50170=>"11111110",
  50171=>"11111111",
  50172=>"00000000",
  50173=>"11111111",
  50174=>"11111110",
  50175=>"00000001",
  50176=>"11111111",
  50177=>"00000101",
  50178=>"11111110",
  50179=>"11111111",
  50180=>"11111111",
  50181=>"00000101",
  50182=>"00000100",
  50183=>"00000000",
  50184=>"00000001",
  50185=>"00000001",
  50186=>"00000010",
  50187=>"00000001",
  50188=>"11111110",
  50189=>"11111100",
  50190=>"00000100",
  50191=>"00000000",
  50192=>"11111111",
  50193=>"11111111",
  50194=>"00000011",
  50195=>"00000100",
  50196=>"00000101",
  50197=>"11111110",
  50198=>"00000000",
  50199=>"11111101",
  50200=>"00000011",
  50201=>"00000011",
  50202=>"11111110",
  50203=>"11111111",
  50204=>"00000000",
  50205=>"11111111",
  50206=>"00000110",
  50207=>"00000010",
  50208=>"11111110",
  50209=>"11111100",
  50210=>"00000001",
  50211=>"00000011",
  50212=>"00000100",
  50213=>"00000011",
  50214=>"11111110",
  50215=>"11111111",
  50216=>"11111111",
  50217=>"00000011",
  50218=>"00000101",
  50219=>"11111110",
  50220=>"00000010",
  50221=>"00000010",
  50222=>"00000011",
  50223=>"00000000",
  50224=>"11111111",
  50225=>"00000010",
  50226=>"00000001",
  50227=>"11111111",
  50228=>"11111110",
  50229=>"00000011",
  50230=>"11111111",
  50231=>"00000010",
  50232=>"00000101",
  50233=>"11111111",
  50234=>"11111101",
  50235=>"11111100",
  50236=>"11111110",
  50237=>"11111110",
  50238=>"00000100",
  50239=>"00000000",
  50240=>"11111101",
  50241=>"00000000",
  50242=>"00000001",
  50243=>"00000000",
  50244=>"11111111",
  50245=>"00000010",
  50246=>"11111111",
  50247=>"00000001",
  50248=>"11111111",
  50249=>"11111110",
  50250=>"11111101",
  50251=>"00000000",
  50252=>"11111110",
  50253=>"11111101",
  50254=>"00000011",
  50255=>"00000001",
  50256=>"00000011",
  50257=>"11111110",
  50258=>"00000010",
  50259=>"11111100",
  50260=>"11111110",
  50261=>"11111110",
  50262=>"00000100",
  50263=>"00000100",
  50264=>"00000011",
  50265=>"11111110",
  50266=>"11111111",
  50267=>"00000011",
  50268=>"11111101",
  50269=>"11111111",
  50270=>"11111111",
  50271=>"11111110",
  50272=>"00000010",
  50273=>"00000011",
  50274=>"00000001",
  50275=>"11111111",
  50276=>"00000000",
  50277=>"11111101",
  50278=>"00000101",
  50279=>"00000101",
  50280=>"11111110",
  50281=>"11111101",
  50282=>"11111111",
  50283=>"00000000",
  50284=>"11111110",
  50285=>"11111100",
  50286=>"11111110",
  50287=>"11111101",
  50288=>"11111110",
  50289=>"11111101",
  50290=>"11111110",
  50291=>"00000001",
  50292=>"11111110",
  50293=>"11111101",
  50294=>"11111111",
  50295=>"11111101",
  50296=>"11111110",
  50297=>"00000001",
  50298=>"11111011",
  50299=>"11111111",
  50300=>"00000001",
  50301=>"11111111",
  50302=>"00000011",
  50303=>"11111111",
  50304=>"00000000",
  50305=>"00000001",
  50306=>"00000011",
  50307=>"00001000",
  50308=>"00000010",
  50309=>"00000000",
  50310=>"00000010",
  50311=>"11111100",
  50312=>"00000100",
  50313=>"11111110",
  50314=>"00000001",
  50315=>"11111101",
  50316=>"00000001",
  50317=>"00000101",
  50318=>"00000000",
  50319=>"00000010",
  50320=>"00000011",
  50321=>"00000000",
  50322=>"11111110",
  50323=>"11111110",
  50324=>"00000000",
  50325=>"00000001",
  50326=>"11111110",
  50327=>"00000011",
  50328=>"11111100",
  50329=>"11111111",
  50330=>"11111111",
  50331=>"00000010",
  50332=>"00000011",
  50333=>"11111110",
  50334=>"11111110",
  50335=>"00000001",
  50336=>"00000110",
  50337=>"00000001",
  50338=>"00000000",
  50339=>"00000100",
  50340=>"00000000",
  50341=>"00000000",
  50342=>"00000010",
  50343=>"11111111",
  50344=>"00000001",
  50345=>"00000000",
  50346=>"11111111",
  50347=>"11111100",
  50348=>"11111100",
  50349=>"00000000",
  50350=>"00000001",
  50351=>"11111110",
  50352=>"11111100",
  50353=>"11111110",
  50354=>"11111111",
  50355=>"00000010",
  50356=>"00000001",
  50357=>"00000011",
  50358=>"00000100",
  50359=>"11111111",
  50360=>"11111111",
  50361=>"00000100",
  50362=>"00000000",
  50363=>"11111111",
  50364=>"11111100",
  50365=>"00000000",
  50366=>"00000010",
  50367=>"00000010",
  50368=>"11111111",
  50369=>"11111110",
  50370=>"00000000",
  50371=>"00000000",
  50372=>"11111111",
  50373=>"11111100",
  50374=>"00000010",
  50375=>"11111110",
  50376=>"00000000",
  50377=>"00000100",
  50378=>"11111111",
  50379=>"00000010",
  50380=>"11111111",
  50381=>"11111110",
  50382=>"00000011",
  50383=>"00000000",
  50384=>"11111110",
  50385=>"11111101",
  50386=>"00000000",
  50387=>"00000011",
  50388=>"11111110",
  50389=>"11111100",
  50390=>"00000001",
  50391=>"11111111",
  50392=>"00000100",
  50393=>"00000100",
  50394=>"00000001",
  50395=>"00000010",
  50396=>"11111111",
  50397=>"11111101",
  50398=>"00000010",
  50399=>"00000000",
  50400=>"00000000",
  50401=>"11111111",
  50402=>"11111101",
  50403=>"11111100",
  50404=>"00000001",
  50405=>"00000011",
  50406=>"11111101",
  50407=>"00000011",
  50408=>"00000010",
  50409=>"11111111",
  50410=>"00000011",
  50411=>"11111111",
  50412=>"00000010",
  50413=>"00000000",
  50414=>"00000101",
  50415=>"11111110",
  50416=>"00000010",
  50417=>"00000000",
  50418=>"00000110",
  50419=>"00000011",
  50420=>"00000010",
  50421=>"11111101",
  50422=>"00000000",
  50423=>"00000000",
  50424=>"11111101",
  50425=>"00000011",
  50426=>"00000000",
  50427=>"00000001",
  50428=>"11111110",
  50429=>"11111101",
  50430=>"11111111",
  50431=>"00000011",
  50432=>"00000001",
  50433=>"11111110",
  50434=>"00000000",
  50435=>"11111110",
  50436=>"00000010",
  50437=>"00000010",
  50438=>"00000000",
  50439=>"11111111",
  50440=>"11111111",
  50441=>"00000010",
  50442=>"00000000",
  50443=>"11111101",
  50444=>"11111111",
  50445=>"00000011",
  50446=>"11111100",
  50447=>"11111101",
  50448=>"11111111",
  50449=>"11111101",
  50450=>"11111100",
  50451=>"00000010",
  50452=>"11111110",
  50453=>"11111110",
  50454=>"11111110",
  50455=>"00000011",
  50456=>"11111100",
  50457=>"00000001",
  50458=>"11111110",
  50459=>"11111110",
  50460=>"11111101",
  50461=>"11111111",
  50462=>"00000001",
  50463=>"00000010",
  50464=>"11111110",
  50465=>"11111111",
  50466=>"11111110",
  50467=>"11111100",
  50468=>"11111110",
  50469=>"11111111",
  50470=>"11111111",
  50471=>"00000000",
  50472=>"11111101",
  50473=>"11111101",
  50474=>"00000011",
  50475=>"11111110",
  50476=>"11111110",
  50477=>"00000011",
  50478=>"00000000",
  50479=>"11111111",
  50480=>"00000010",
  50481=>"00000001",
  50482=>"11111100",
  50483=>"11111101",
  50484=>"00000110",
  50485=>"11111101",
  50486=>"00000010",
  50487=>"11111101",
  50488=>"11111100",
  50489=>"00000011",
  50490=>"11111110",
  50491=>"11111101",
  50492=>"11111101",
  50493=>"00001000",
  50494=>"00000101",
  50495=>"00000001",
  50496=>"00000000",
  50497=>"11111101",
  50498=>"00000000",
  50499=>"00000000",
  50500=>"11111111",
  50501=>"00000011",
  50502=>"11111101",
  50503=>"00000000",
  50504=>"11111101",
  50505=>"00000010",
  50506=>"11111101",
  50507=>"11111111",
  50508=>"00000010",
  50509=>"00000010",
  50510=>"00000010",
  50511=>"00000000",
  50512=>"00000001",
  50513=>"00000000",
  50514=>"00000101",
  50515=>"00000001",
  50516=>"00000010",
  50517=>"00000001",
  50518=>"00000000",
  50519=>"00000010",
  50520=>"00000001",
  50521=>"00000101",
  50522=>"00000101",
  50523=>"00000010",
  50524=>"00000011",
  50525=>"00000011",
  50526=>"11111101",
  50527=>"11111110",
  50528=>"00000110",
  50529=>"11111111",
  50530=>"00000001",
  50531=>"11111110",
  50532=>"11111111",
  50533=>"00000011",
  50534=>"00000010",
  50535=>"00000000",
  50536=>"00000010",
  50537=>"00000011",
  50538=>"00000010",
  50539=>"11111110",
  50540=>"00000010",
  50541=>"11111101",
  50542=>"00000001",
  50543=>"11111111",
  50544=>"00000011",
  50545=>"00000011",
  50546=>"00000011",
  50547=>"00000010",
  50548=>"11111111",
  50549=>"11111111",
  50550=>"00000000",
  50551=>"00000011",
  50552=>"11111101",
  50553=>"11111111",
  50554=>"00000000",
  50555=>"11111100",
  50556=>"00000000",
  50557=>"00000001",
  50558=>"11111110",
  50559=>"11111110",
  50560=>"11111110",
  50561=>"00000100",
  50562=>"00000001",
  50563=>"00000000",
  50564=>"00000010",
  50565=>"11111111",
  50566=>"11111101",
  50567=>"00000101",
  50568=>"00000000",
  50569=>"00000011",
  50570=>"11111101",
  50571=>"00000000",
  50572=>"11111101",
  50573=>"00000110",
  50574=>"00000100",
  50575=>"00000100",
  50576=>"00000000",
  50577=>"00000000",
  50578=>"11111111",
  50579=>"00000010",
  50580=>"11111110",
  50581=>"11111110",
  50582=>"00000000",
  50583=>"00000000",
  50584=>"00000011",
  50585=>"11111100",
  50586=>"00000001",
  50587=>"11111100",
  50588=>"00000010",
  50589=>"00000001",
  50590=>"00000010",
  50591=>"00000010",
  50592=>"11111111",
  50593=>"11111111",
  50594=>"11111110",
  50595=>"00000111",
  50596=>"11111101",
  50597=>"00000000",
  50598=>"00000010",
  50599=>"00000000",
  50600=>"11111101",
  50601=>"11111101",
  50602=>"00000011",
  50603=>"11111110",
  50604=>"11111101",
  50605=>"11111111",
  50606=>"00000110",
  50607=>"00000001",
  50608=>"11111111",
  50609=>"00000000",
  50610=>"00000001",
  50611=>"00000001",
  50612=>"00000001",
  50613=>"00000010",
  50614=>"11111101",
  50615=>"11111111",
  50616=>"11111101",
  50617=>"00000100",
  50618=>"00000000",
  50619=>"00000010",
  50620=>"11111111",
  50621=>"11111111",
  50622=>"11111111",
  50623=>"00000010",
  50624=>"00000010",
  50625=>"11111100",
  50626=>"00000001",
  50627=>"11111111",
  50628=>"00000000",
  50629=>"00000001",
  50630=>"11111110",
  50631=>"00000000",
  50632=>"00000000",
  50633=>"11111110",
  50634=>"00000011",
  50635=>"00000011",
  50636=>"00000010",
  50637=>"00000010",
  50638=>"11111111",
  50639=>"11111110",
  50640=>"11111111",
  50641=>"00000010",
  50642=>"00000011",
  50643=>"00000100",
  50644=>"00000011",
  50645=>"00000010",
  50646=>"11111101",
  50647=>"00000010",
  50648=>"00000001",
  50649=>"00000001",
  50650=>"00000010",
  50651=>"11111100",
  50652=>"00000110",
  50653=>"11111111",
  50654=>"00000010",
  50655=>"00000001",
  50656=>"11111101",
  50657=>"11111111",
  50658=>"11111111",
  50659=>"00000001",
  50660=>"11111111",
  50661=>"11111110",
  50662=>"11111101",
  50663=>"00000011",
  50664=>"11111111",
  50665=>"11111101",
  50666=>"00000010",
  50667=>"11111101",
  50668=>"00000001",
  50669=>"11111101",
  50670=>"00000000",
  50671=>"11111100",
  50672=>"11111101",
  50673=>"00000000",
  50674=>"11111110",
  50675=>"00000101",
  50676=>"00000000",
  50677=>"11111110",
  50678=>"00000001",
  50679=>"11111101",
  50680=>"11111100",
  50681=>"11111111",
  50682=>"11111101",
  50683=>"11111101",
  50684=>"00000000",
  50685=>"00000001",
  50686=>"00000001",
  50687=>"00000011",
  50688=>"00000001",
  50689=>"00000010",
  50690=>"00000001",
  50691=>"00000010",
  50692=>"11111100",
  50693=>"00000011",
  50694=>"11111111",
  50695=>"00000000",
  50696=>"00000100",
  50697=>"11111100",
  50698=>"00000011",
  50699=>"00000010",
  50700=>"11111111",
  50701=>"00000001",
  50702=>"00000100",
  50703=>"11111110",
  50704=>"00000110",
  50705=>"00000011",
  50706=>"11111101",
  50707=>"00000001",
  50708=>"11111111",
  50709=>"00000011",
  50710=>"00000001",
  50711=>"11111110",
  50712=>"11111101",
  50713=>"00000000",
  50714=>"11111110",
  50715=>"00000011",
  50716=>"00000000",
  50717=>"00000001",
  50718=>"00000100",
  50719=>"00000010",
  50720=>"00000000",
  50721=>"11111111",
  50722=>"00000000",
  50723=>"00000001",
  50724=>"00000000",
  50725=>"00000001",
  50726=>"11111110",
  50727=>"11111111",
  50728=>"00000101",
  50729=>"11111101",
  50730=>"11111100",
  50731=>"11111110",
  50732=>"11111110",
  50733=>"11111101",
  50734=>"11111101",
  50735=>"11111111",
  50736=>"00000101",
  50737=>"11111111",
  50738=>"00000100",
  50739=>"11111101",
  50740=>"11111101",
  50741=>"00000000",
  50742=>"11111110",
  50743=>"11111111",
  50744=>"11111101",
  50745=>"00000000",
  50746=>"11111110",
  50747=>"00000000",
  50748=>"11111101",
  50749=>"00000110",
  50750=>"11111111",
  50751=>"00000100",
  50752=>"11111111",
  50753=>"00000010",
  50754=>"11111111",
  50755=>"00000000",
  50756=>"00000011",
  50757=>"00000001",
  50758=>"00000110",
  50759=>"00000000",
  50760=>"00000010",
  50761=>"11111110",
  50762=>"00000010",
  50763=>"11111101",
  50764=>"11111101",
  50765=>"00000110",
  50766=>"00000011",
  50767=>"11111101",
  50768=>"11111110",
  50769=>"00000001",
  50770=>"11111110",
  50771=>"11111111",
  50772=>"11111101",
  50773=>"00000000",
  50774=>"00000001",
  50775=>"11111101",
  50776=>"00000110",
  50777=>"00000001",
  50778=>"00000010",
  50779=>"11111111",
  50780=>"00000001",
  50781=>"11111110",
  50782=>"11111101",
  50783=>"11111101",
  50784=>"11111101",
  50785=>"11111111",
  50786=>"00000010",
  50787=>"00000011",
  50788=>"00000110",
  50789=>"00000000",
  50790=>"11111111",
  50791=>"00000000",
  50792=>"00000001",
  50793=>"00000010",
  50794=>"00000010",
  50795=>"00000010",
  50796=>"00000001",
  50797=>"11111111",
  50798=>"00000101",
  50799=>"00000100",
  50800=>"11111100",
  50801=>"00000010",
  50802=>"11111110",
  50803=>"11111101",
  50804=>"00000001",
  50805=>"11111111",
  50806=>"11111110",
  50807=>"00000000",
  50808=>"11111111",
  50809=>"00000011",
  50810=>"00000000",
  50811=>"11111110",
  50812=>"11111110",
  50813=>"00000010",
  50814=>"11111101",
  50815=>"11111110",
  50816=>"11111110",
  50817=>"00000001",
  50818=>"00000010",
  50819=>"00000011",
  50820=>"11111110",
  50821=>"11111100",
  50822=>"00000000",
  50823=>"11111101",
  50824=>"00000011",
  50825=>"11111110",
  50826=>"00000111",
  50827=>"11111111",
  50828=>"00000000",
  50829=>"00000011",
  50830=>"00000000",
  50831=>"00000000",
  50832=>"00000000",
  50833=>"11111110",
  50834=>"00000001",
  50835=>"11111111",
  50836=>"00000001",
  50837=>"00000111",
  50838=>"00000000",
  50839=>"11111101",
  50840=>"00000010",
  50841=>"11111100",
  50842=>"11111111",
  50843=>"00000011",
  50844=>"00000001",
  50845=>"00000010",
  50846=>"11111101",
  50847=>"00000011",
  50848=>"00000000",
  50849=>"00000011",
  50850=>"00000001",
  50851=>"00000101",
  50852=>"11111101",
  50853=>"00000000",
  50854=>"00000000",
  50855=>"00000010",
  50856=>"00000001",
  50857=>"00000000",
  50858=>"11111111",
  50859=>"11111101",
  50860=>"11111111",
  50861=>"00000010",
  50862=>"00000011",
  50863=>"11111110",
  50864=>"11111111",
  50865=>"11111110",
  50866=>"00000000",
  50867=>"11111100",
  50868=>"11111111",
  50869=>"00000010",
  50870=>"00000000",
  50871=>"11111101",
  50872=>"00000011",
  50873=>"00000010",
  50874=>"11111110",
  50875=>"00000000",
  50876=>"11111110",
  50877=>"11111111",
  50878=>"11111111",
  50879=>"00000000",
  50880=>"11111100",
  50881=>"11111110",
  50882=>"11111110",
  50883=>"11111101",
  50884=>"11111110",
  50885=>"11111101",
  50886=>"00000011",
  50887=>"00000001",
  50888=>"00000010",
  50889=>"00000010",
  50890=>"00000001",
  50891=>"11111111",
  50892=>"11111110",
  50893=>"11111111",
  50894=>"00000010",
  50895=>"11111111",
  50896=>"00000001",
  50897=>"00000110",
  50898=>"00000010",
  50899=>"00000001",
  50900=>"00000010",
  50901=>"00000011",
  50902=>"00000010",
  50903=>"00000000",
  50904=>"00000001",
  50905=>"00000010",
  50906=>"11111110",
  50907=>"00000001",
  50908=>"11111100",
  50909=>"00000001",
  50910=>"11111101",
  50911=>"11111110",
  50912=>"00000010",
  50913=>"00000000",
  50914=>"11111110",
  50915=>"00000101",
  50916=>"00000001",
  50917=>"11111100",
  50918=>"00000010",
  50919=>"11111111",
  50920=>"00000000",
  50921=>"00000001",
  50922=>"00000001",
  50923=>"00000100",
  50924=>"00000011",
  50925=>"11111101",
  50926=>"00000010",
  50927=>"11111110",
  50928=>"11111101",
  50929=>"00000011",
  50930=>"11111111",
  50931=>"00000010",
  50932=>"00000010",
  50933=>"11111101",
  50934=>"11111111",
  50935=>"00000000",
  50936=>"11111101",
  50937=>"00000000",
  50938=>"11111111",
  50939=>"11111100",
  50940=>"00000011",
  50941=>"11111101",
  50942=>"11111110",
  50943=>"00000000",
  50944=>"00000100",
  50945=>"11111111",
  50946=>"00000000",
  50947=>"11111111",
  50948=>"00000011",
  50949=>"00000000",
  50950=>"00000000",
  50951=>"00000000",
  50952=>"00000100",
  50953=>"00000101",
  50954=>"11111111",
  50955=>"00000001",
  50956=>"11111101",
  50957=>"00000010",
  50958=>"11111111",
  50959=>"11111111",
  50960=>"00000010",
  50961=>"00000001",
  50962=>"00000101",
  50963=>"00000001",
  50964=>"00000011",
  50965=>"11111110",
  50966=>"11111100",
  50967=>"00000100",
  50968=>"00000010",
  50969=>"11111110",
  50970=>"11111100",
  50971=>"00000010",
  50972=>"00000010",
  50973=>"11111101",
  50974=>"11111111",
  50975=>"00000000",
  50976=>"00000010",
  50977=>"00000100",
  50978=>"00000010",
  50979=>"11111110",
  50980=>"11111111",
  50981=>"11111011",
  50982=>"11111111",
  50983=>"11111100",
  50984=>"11111101",
  50985=>"00000001",
  50986=>"00000001",
  50987=>"11111101",
  50988=>"11111111",
  50989=>"11111110",
  50990=>"00000000",
  50991=>"00000100",
  50992=>"00000010",
  50993=>"11111111",
  50994=>"11111110",
  50995=>"00000011",
  50996=>"00000001",
  50997=>"11111111",
  50998=>"00000001",
  50999=>"00000000",
  51000=>"00000010",
  51001=>"00000001",
  51002=>"00000101",
  51003=>"00000000",
  51004=>"00000010",
  51005=>"11111111",
  51006=>"00000010",
  51007=>"00000001",
  51008=>"11111111",
  51009=>"00000010",
  51010=>"00000000",
  51011=>"00000000",
  51012=>"00000000",
  51013=>"11111110",
  51014=>"11111110",
  51015=>"00000001",
  51016=>"00000001",
  51017=>"11111101",
  51018=>"00000000",
  51019=>"11111110",
  51020=>"11111111",
  51021=>"11111101",
  51022=>"00000000",
  51023=>"11111110",
  51024=>"11111111",
  51025=>"00000000",
  51026=>"00000110",
  51027=>"00000010",
  51028=>"11111101",
  51029=>"00000000",
  51030=>"11111110",
  51031=>"00000101",
  51032=>"00000010",
  51033=>"11111101",
  51034=>"11111111",
  51035=>"00000000",
  51036=>"00000000",
  51037=>"11111101",
  51038=>"11111110",
  51039=>"00000001",
  51040=>"00000000",
  51041=>"00000011",
  51042=>"00000100",
  51043=>"11111110",
  51044=>"11111110",
  51045=>"11111111",
  51046=>"00000001",
  51047=>"00000100",
  51048=>"11111111",
  51049=>"11111110",
  51050=>"11111110",
  51051=>"00000010",
  51052=>"00000001",
  51053=>"11111110",
  51054=>"11111101",
  51055=>"00000011",
  51056=>"00000011",
  51057=>"00000011",
  51058=>"00000001",
  51059=>"00000110",
  51060=>"11111111",
  51061=>"00000000",
  51062=>"00000100",
  51063=>"11111111",
  51064=>"00000001",
  51065=>"11111100",
  51066=>"00000010",
  51067=>"11111111",
  51068=>"11111101",
  51069=>"11111101",
  51070=>"00000001",
  51071=>"00000100",
  51072=>"11111110",
  51073=>"00000000",
  51074=>"11111101",
  51075=>"11111101",
  51076=>"00000011",
  51077=>"00000001",
  51078=>"11111101",
  51079=>"00000000",
  51080=>"11111101",
  51081=>"11111101",
  51082=>"00000000",
  51083=>"11111111",
  51084=>"00000000",
  51085=>"11111111",
  51086=>"11111110",
  51087=>"00000000",
  51088=>"11111111",
  51089=>"00000011",
  51090=>"11111111",
  51091=>"00000000",
  51092=>"00000001",
  51093=>"11111100",
  51094=>"00000001",
  51095=>"00000000",
  51096=>"11111111",
  51097=>"00000000",
  51098=>"11111101",
  51099=>"00000000",
  51100=>"00000011",
  51101=>"11111111",
  51102=>"11111110",
  51103=>"00000010",
  51104=>"00000100",
  51105=>"11111110",
  51106=>"11111100",
  51107=>"00000011",
  51108=>"00000100",
  51109=>"11111101",
  51110=>"11111111",
  51111=>"11111101",
  51112=>"00000000",
  51113=>"00000011",
  51114=>"00000010",
  51115=>"11111110",
  51116=>"11111100",
  51117=>"11111110",
  51118=>"00000000",
  51119=>"00000000",
  51120=>"00000101",
  51121=>"00000010",
  51122=>"00000001",
  51123=>"11111111",
  51124=>"11111110",
  51125=>"11111111",
  51126=>"00000001",
  51127=>"11111110",
  51128=>"00000100",
  51129=>"00000000",
  51130=>"00000010",
  51131=>"00000001",
  51132=>"11111111",
  51133=>"00000100",
  51134=>"00000000",
  51135=>"00000011",
  51136=>"11111101",
  51137=>"11111110",
  51138=>"00000000",
  51139=>"11111110",
  51140=>"00000001",
  51141=>"00000011",
  51142=>"11111111",
  51143=>"11111111",
  51144=>"00000001",
  51145=>"00000101",
  51146=>"11111011",
  51147=>"00000010",
  51148=>"11111100",
  51149=>"00000000",
  51150=>"11111101",
  51151=>"00000011",
  51152=>"00000000",
  51153=>"00000010",
  51154=>"00000000",
  51155=>"00000000",
  51156=>"11111111",
  51157=>"11111111",
  51158=>"00000101",
  51159=>"11111111",
  51160=>"00000010",
  51161=>"00000001",
  51162=>"00000101",
  51163=>"11111101",
  51164=>"00000001",
  51165=>"11111100",
  51166=>"00000011",
  51167=>"00000010",
  51168=>"00000001",
  51169=>"11111111",
  51170=>"00000100",
  51171=>"11111101",
  51172=>"11111111",
  51173=>"11111101",
  51174=>"11111101",
  51175=>"11111110",
  51176=>"11111110",
  51177=>"00000000",
  51178=>"11111011",
  51179=>"11111101",
  51180=>"11111110",
  51181=>"11111110",
  51182=>"11111110",
  51183=>"00000010",
  51184=>"11111100",
  51185=>"00000001",
  51186=>"11111110",
  51187=>"00000001",
  51188=>"00000010",
  51189=>"00000000",
  51190=>"00000010",
  51191=>"00000001",
  51192=>"00000011",
  51193=>"00000001",
  51194=>"00000000",
  51195=>"11111111",
  51196=>"00000010",
  51197=>"00000001",
  51198=>"11111110",
  51199=>"00000000",
  51200=>"11111110",
  51201=>"11111111",
  51202=>"00000000",
  51203=>"00000000",
  51204=>"11111111",
  51205=>"00000001",
  51206=>"00000001",
  51207=>"00000000",
  51208=>"11111111",
  51209=>"00000001",
  51210=>"00000001",
  51211=>"11111111",
  51212=>"00000001",
  51213=>"00000001",
  51214=>"00000001",
  51215=>"00000010",
  51216=>"00000000",
  51217=>"00000000",
  51218=>"00000001",
  51219=>"00000000",
  51220=>"11111111",
  51221=>"11111110",
  51222=>"00000001",
  51223=>"11111110",
  51224=>"00000001",
  51225=>"00000001",
  51226=>"00000000",
  51227=>"00000001",
  51228=>"00000000",
  51229=>"00000001",
  51230=>"00000001",
  51231=>"11111110",
  51232=>"00000000",
  51233=>"11111111",
  51234=>"00000001",
  51235=>"00000010",
  51236=>"11111111",
  51237=>"00000000",
  51238=>"00000000",
  51239=>"11111111",
  51240=>"11111110",
  51241=>"11111111",
  51242=>"11111111",
  51243=>"00000001",
  51244=>"00000001",
  51245=>"11111100",
  51246=>"00000001",
  51247=>"00000000",
  51248=>"11111111",
  51249=>"11111110",
  51250=>"00000001",
  51251=>"00000000",
  51252=>"11111101",
  51253=>"00000000",
  51254=>"00000001",
  51255=>"11111111",
  51256=>"11111111",
  51257=>"11111111",
  51258=>"00000000",
  51259=>"00000000",
  51260=>"00000001",
  51261=>"11111111",
  51262=>"00000001",
  51263=>"00000000",
  51264=>"00000001",
  51265=>"11111111",
  51266=>"00000000",
  51267=>"00000010",
  51268=>"00000010",
  51269=>"00000001",
  51270=>"00000010",
  51271=>"00000010",
  51272=>"00000010",
  51273=>"00000000",
  51274=>"00000010",
  51275=>"00000001",
  51276=>"00000001",
  51277=>"00000001",
  51278=>"11111111",
  51279=>"00000010",
  51280=>"11111111",
  51281=>"00000010",
  51282=>"00000000",
  51283=>"00000000",
  51284=>"00000000",
  51285=>"11111110",
  51286=>"00000001",
  51287=>"00000001",
  51288=>"11111111",
  51289=>"11111111",
  51290=>"11111110",
  51291=>"00000001",
  51292=>"00000001",
  51293=>"00000010",
  51294=>"00000000",
  51295=>"11111111",
  51296=>"00000000",
  51297=>"00000000",
  51298=>"11111110",
  51299=>"11111111",
  51300=>"00000000",
  51301=>"00000010",
  51302=>"11111111",
  51303=>"11111111",
  51304=>"11111111",
  51305=>"11111111",
  51306=>"11111111",
  51307=>"00000001",
  51308=>"00000001",
  51309=>"00000000",
  51310=>"00000000",
  51311=>"11111111",
  51312=>"11111111",
  51313=>"11111111",
  51314=>"00000010",
  51315=>"00000001",
  51316=>"11111110",
  51317=>"00000000",
  51318=>"00000001",
  51319=>"00000000",
  51320=>"00000001",
  51321=>"00000000",
  51322=>"11111111",
  51323=>"00000000",
  51324=>"00000000",
  51325=>"00000001",
  51326=>"00000010",
  51327=>"00000001",
  51328=>"00000000",
  51329=>"00000001",
  51330=>"11111110",
  51331=>"00000011",
  51332=>"00000010",
  51333=>"11111111",
  51334=>"11111111",
  51335=>"11111110",
  51336=>"11111111",
  51337=>"00000000",
  51338=>"00000010",
  51339=>"00000000",
  51340=>"00000010",
  51341=>"00000001",
  51342=>"00000000",
  51343=>"11111110",
  51344=>"00000001",
  51345=>"11111111",
  51346=>"00000001",
  51347=>"00000001",
  51348=>"00000001",
  51349=>"00000001",
  51350=>"11111111",
  51351=>"00000000",
  51352=>"11111111",
  51353=>"00000000",
  51354=>"11111110",
  51355=>"00000001",
  51356=>"00000010",
  51357=>"00000001",
  51358=>"00000001",
  51359=>"00000000",
  51360=>"00000001",
  51361=>"00000001",
  51362=>"11111111",
  51363=>"00000001",
  51364=>"00000010",
  51365=>"00000001",
  51366=>"00000001",
  51367=>"00000000",
  51368=>"11111111",
  51369=>"00000001",
  51370=>"00000000",
  51371=>"00000001",
  51372=>"11111111",
  51373=>"00000001",
  51374=>"00000010",
  51375=>"00000001",
  51376=>"11111111",
  51377=>"00000001",
  51378=>"11111111",
  51379=>"00000001",
  51380=>"11111111",
  51381=>"00000000",
  51382=>"11111111",
  51383=>"11111111",
  51384=>"00000001",
  51385=>"00000000",
  51386=>"11111111",
  51387=>"00000001",
  51388=>"11111110",
  51389=>"00000001",
  51390=>"11111111",
  51391=>"11111111",
  51392=>"11111111",
  51393=>"00000000",
  51394=>"00000001",
  51395=>"00000000",
  51396=>"11111111",
  51397=>"00000000",
  51398=>"00000000",
  51399=>"11111110",
  51400=>"00000000",
  51401=>"11111111",
  51402=>"11111111",
  51403=>"11111111",
  51404=>"00000010",
  51405=>"11111110",
  51406=>"11111110",
  51407=>"11111111",
  51408=>"00000001",
  51409=>"00000001",
  51410=>"11111110",
  51411=>"11111111",
  51412=>"11111110",
  51413=>"00000000",
  51414=>"00000000",
  51415=>"00000001",
  51416=>"00000001",
  51417=>"00000001",
  51418=>"00000001",
  51419=>"11111110",
  51420=>"00000000",
  51421=>"00000010",
  51422=>"11111111",
  51423=>"00000001",
  51424=>"00000000",
  51425=>"00000000",
  51426=>"00000001",
  51427=>"00000001",
  51428=>"11111101",
  51429=>"00000000",
  51430=>"00000010",
  51431=>"11111111",
  51432=>"11111111",
  51433=>"00000001",
  51434=>"00000000",
  51435=>"00000000",
  51436=>"11111111",
  51437=>"00000001",
  51438=>"00000000",
  51439=>"00000010",
  51440=>"00000000",
  51441=>"00000000",
  51442=>"11111111",
  51443=>"00000000",
  51444=>"00000001",
  51445=>"00000000",
  51446=>"00000000",
  51447=>"00000001",
  51448=>"00000000",
  51449=>"11111111",
  51450=>"00000001",
  51451=>"00000001",
  51452=>"11111111",
  51453=>"00000001",
  51454=>"00000000",
  51455=>"00000001",
  51456=>"00000000",
  51457=>"00000000",
  51458=>"11111111",
  51459=>"00000000",
  51460=>"00000010",
  51461=>"11111110",
  51462=>"00000010",
  51463=>"11111111",
  51464=>"11111110",
  51465=>"00000001",
  51466=>"00000001",
  51467=>"11111111",
  51468=>"00000000",
  51469=>"00000000",
  51470=>"11111111",
  51471=>"00000001",
  51472=>"00000001",
  51473=>"11111110",
  51474=>"00000000",
  51475=>"00000010",
  51476=>"00000010",
  51477=>"00000001",
  51478=>"00000000",
  51479=>"00000000",
  51480=>"00000001",
  51481=>"00000001",
  51482=>"00000100",
  51483=>"00000001",
  51484=>"11111111",
  51485=>"00000000",
  51486=>"11111111",
  51487=>"00000000",
  51488=>"00000001",
  51489=>"11111111",
  51490=>"11111111",
  51491=>"00000000",
  51492=>"00000001",
  51493=>"00000000",
  51494=>"00000001",
  51495=>"00000000",
  51496=>"11111111",
  51497=>"00000000",
  51498=>"00000010",
  51499=>"00000001",
  51500=>"11111111",
  51501=>"00000010",
  51502=>"11111111",
  51503=>"11111110",
  51504=>"11111111",
  51505=>"00000000",
  51506=>"00000010",
  51507=>"11111110",
  51508=>"11111111",
  51509=>"00000010",
  51510=>"11111111",
  51511=>"00000010",
  51512=>"11111111",
  51513=>"00000000",
  51514=>"00000010",
  51515=>"00000000",
  51516=>"00000001",
  51517=>"11111111",
  51518=>"11111110",
  51519=>"11111111",
  51520=>"00000001",
  51521=>"00000000",
  51522=>"00000010",
  51523=>"00000000",
  51524=>"11111101",
  51525=>"00000001",
  51526=>"00000001",
  51527=>"11111111",
  51528=>"11111111",
  51529=>"00000010",
  51530=>"00000001",
  51531=>"11111111",
  51532=>"00000001",
  51533=>"00000010",
  51534=>"11111111",
  51535=>"00000001",
  51536=>"00000000",
  51537=>"00000000",
  51538=>"00000010",
  51539=>"00000001",
  51540=>"11111111",
  51541=>"00000000",
  51542=>"00000000",
  51543=>"11111110",
  51544=>"00000000",
  51545=>"11111111",
  51546=>"00000001",
  51547=>"11111111",
  51548=>"11111110",
  51549=>"00000001",
  51550=>"00000001",
  51551=>"00000001",
  51552=>"11111111",
  51553=>"11111111",
  51554=>"11111111",
  51555=>"00000000",
  51556=>"11111110",
  51557=>"11111110",
  51558=>"11111111",
  51559=>"00000000",
  51560=>"00000000",
  51561=>"11111111",
  51562=>"00000001",
  51563=>"00000000",
  51564=>"11111110",
  51565=>"11111111",
  51566=>"11111111",
  51567=>"00000000",
  51568=>"00000000",
  51569=>"11111111",
  51570=>"11111111",
  51571=>"11111111",
  51572=>"00000000",
  51573=>"00000000",
  51574=>"00000001",
  51575=>"11111110",
  51576=>"00000001",
  51577=>"11111110",
  51578=>"00000000",
  51579=>"00000001",
  51580=>"00000001",
  51581=>"11111111",
  51582=>"00000000",
  51583=>"11111111",
  51584=>"00000000",
  51585=>"00000001",
  51586=>"00000000",
  51587=>"00000000",
  51588=>"00000001",
  51589=>"11111111",
  51590=>"00000001",
  51591=>"00000000",
  51592=>"00000000",
  51593=>"00000001",
  51594=>"00000010",
  51595=>"00000000",
  51596=>"00000000",
  51597=>"00000000",
  51598=>"00000001",
  51599=>"00000001",
  51600=>"00000001",
  51601=>"00000010",
  51602=>"11111111",
  51603=>"00000000",
  51604=>"00000000",
  51605=>"00000001",
  51606=>"00000001",
  51607=>"11111111",
  51608=>"00000010",
  51609=>"11111111",
  51610=>"11111111",
  51611=>"00000010",
  51612=>"11111111",
  51613=>"00000001",
  51614=>"00000001",
  51615=>"00000000",
  51616=>"00000000",
  51617=>"00000001",
  51618=>"00000001",
  51619=>"11111111",
  51620=>"11111111",
  51621=>"00000000",
  51622=>"00000000",
  51623=>"00000000",
  51624=>"00000000",
  51625=>"00000000",
  51626=>"00000001",
  51627=>"11111111",
  51628=>"00000001",
  51629=>"00000000",
  51630=>"11111110",
  51631=>"00000001",
  51632=>"11111111",
  51633=>"00000000",
  51634=>"00000010",
  51635=>"00000010",
  51636=>"11111111",
  51637=>"00000000",
  51638=>"11111111",
  51639=>"11111111",
  51640=>"00000000",
  51641=>"11111111",
  51642=>"11111110",
  51643=>"00000001",
  51644=>"00000010",
  51645=>"11111111",
  51646=>"00000000",
  51647=>"11111110",
  51648=>"11111111",
  51649=>"11111111",
  51650=>"00000000",
  51651=>"11111111",
  51652=>"00000000",
  51653=>"00000010",
  51654=>"00000001",
  51655=>"00000000",
  51656=>"00000000",
  51657=>"11111111",
  51658=>"00000000",
  51659=>"00000000",
  51660=>"00000010",
  51661=>"00000000",
  51662=>"11111111",
  51663=>"00000000",
  51664=>"00000001",
  51665=>"11111111",
  51666=>"11111111",
  51667=>"00000001",
  51668=>"00000001",
  51669=>"00000000",
  51670=>"00000001",
  51671=>"00000000",
  51672=>"11111111",
  51673=>"11111110",
  51674=>"00000000",
  51675=>"00000000",
  51676=>"00000000",
  51677=>"00000000",
  51678=>"00000000",
  51679=>"11111111",
  51680=>"00000000",
  51681=>"00000001",
  51682=>"00000000",
  51683=>"11111101",
  51684=>"00000001",
  51685=>"11111110",
  51686=>"11111111",
  51687=>"11111110",
  51688=>"00000000",
  51689=>"00000000",
  51690=>"00000001",
  51691=>"00000000",
  51692=>"00000000",
  51693=>"00000010",
  51694=>"00000001",
  51695=>"00000001",
  51696=>"00000010",
  51697=>"00000010",
  51698=>"00000001",
  51699=>"00000001",
  51700=>"11111111",
  51701=>"00000000",
  51702=>"11111111",
  51703=>"00000000",
  51704=>"00000001",
  51705=>"11111111",
  51706=>"00000001",
  51707=>"00000010",
  51708=>"00000001",
  51709=>"11111111",
  51710=>"11111111",
  51711=>"00000000",
  51712=>"00000010",
  51713=>"00000001",
  51714=>"00000000",
  51715=>"00000000",
  51716=>"11111110",
  51717=>"00000010",
  51718=>"00000000",
  51719=>"11111111",
  51720=>"00000001",
  51721=>"00000001",
  51722=>"00000010",
  51723=>"00000010",
  51724=>"00000000",
  51725=>"00000000",
  51726=>"00000010",
  51727=>"00000000",
  51728=>"11111111",
  51729=>"00000000",
  51730=>"00000001",
  51731=>"11111111",
  51732=>"11111111",
  51733=>"11111111",
  51734=>"00000000",
  51735=>"11111110",
  51736=>"00000000",
  51737=>"11111111",
  51738=>"11111101",
  51739=>"11111110",
  51740=>"00000000",
  51741=>"00000000",
  51742=>"11111110",
  51743=>"11111111",
  51744=>"00000000",
  51745=>"00000001",
  51746=>"00000010",
  51747=>"00000000",
  51748=>"00000001",
  51749=>"00000001",
  51750=>"00000010",
  51751=>"00000000",
  51752=>"11111111",
  51753=>"00000000",
  51754=>"11111111",
  51755=>"00000000",
  51756=>"00000000",
  51757=>"11111111",
  51758=>"00000001",
  51759=>"00000001",
  51760=>"00000001",
  51761=>"00000000",
  51762=>"00000010",
  51763=>"11111101",
  51764=>"00000001",
  51765=>"00000000",
  51766=>"00000000",
  51767=>"11111111",
  51768=>"00000000",
  51769=>"11111110",
  51770=>"00000001",
  51771=>"11111110",
  51772=>"00000001",
  51773=>"00000000",
  51774=>"11111111",
  51775=>"11111110",
  51776=>"00000000",
  51777=>"00000001",
  51778=>"00000000",
  51779=>"11111111",
  51780=>"00000001",
  51781=>"11111110",
  51782=>"00000000",
  51783=>"11111110",
  51784=>"00000000",
  51785=>"00000000",
  51786=>"00000000",
  51787=>"00000000",
  51788=>"00000010",
  51789=>"00000000",
  51790=>"11111111",
  51791=>"00000001",
  51792=>"00000010",
  51793=>"11111111",
  51794=>"00000010",
  51795=>"00000001",
  51796=>"00000001",
  51797=>"11111111",
  51798=>"00000001",
  51799=>"11111110",
  51800=>"00000000",
  51801=>"00000000",
  51802=>"00000000",
  51803=>"11111111",
  51804=>"00000000",
  51805=>"00000001",
  51806=>"11111111",
  51807=>"00000001",
  51808=>"11111111",
  51809=>"00000001",
  51810=>"00000001",
  51811=>"11111111",
  51812=>"00000001",
  51813=>"11111111",
  51814=>"00000000",
  51815=>"00000000",
  51816=>"00000000",
  51817=>"00000001",
  51818=>"00000000",
  51819=>"11111111",
  51820=>"11111111",
  51821=>"00000010",
  51822=>"00000010",
  51823=>"00000001",
  51824=>"00000010",
  51825=>"00000010",
  51826=>"00000001",
  51827=>"11111111",
  51828=>"11111111",
  51829=>"00000001",
  51830=>"00000001",
  51831=>"00000000",
  51832=>"11111111",
  51833=>"00000000",
  51834=>"00000001",
  51835=>"00000000",
  51836=>"11111110",
  51837=>"11111111",
  51838=>"11111111",
  51839=>"11111110",
  51840=>"00000010",
  51841=>"11111111",
  51842=>"00000000",
  51843=>"11111111",
  51844=>"00000000",
  51845=>"00000000",
  51846=>"00000001",
  51847=>"00000000",
  51848=>"11111111",
  51849=>"11111111",
  51850=>"00000001",
  51851=>"11111111",
  51852=>"11111110",
  51853=>"00000001",
  51854=>"11111111",
  51855=>"00000001",
  51856=>"00000000",
  51857=>"00000001",
  51858=>"00000000",
  51859=>"00000001",
  51860=>"00000001",
  51861=>"00000000",
  51862=>"00000000",
  51863=>"00000001",
  51864=>"00000001",
  51865=>"00000000",
  51866=>"00000001",
  51867=>"00000001",
  51868=>"11111110",
  51869=>"11111111",
  51870=>"00000001",
  51871=>"00000001",
  51872=>"11111111",
  51873=>"00000000",
  51874=>"00000010",
  51875=>"00000001",
  51876=>"00000000",
  51877=>"00000000",
  51878=>"11111111",
  51879=>"00000010",
  51880=>"00000001",
  51881=>"11111111",
  51882=>"11111111",
  51883=>"00000011",
  51884=>"00000001",
  51885=>"11111111",
  51886=>"00000001",
  51887=>"00000000",
  51888=>"11111111",
  51889=>"11111111",
  51890=>"11111110",
  51891=>"11111111",
  51892=>"00000001",
  51893=>"11111111",
  51894=>"11111111",
  51895=>"11111111",
  51896=>"11111111",
  51897=>"11111110",
  51898=>"00000010",
  51899=>"00000000",
  51900=>"11111111",
  51901=>"00000000",
  51902=>"11111111",
  51903=>"00000000",
  51904=>"00000000",
  51905=>"11111111",
  51906=>"11111111",
  51907=>"11111111",
  51908=>"00000001",
  51909=>"00000000",
  51910=>"11111111",
  51911=>"00000000",
  51912=>"00000000",
  51913=>"00000000",
  51914=>"11111111",
  51915=>"11111110",
  51916=>"00000000",
  51917=>"11111111",
  51918=>"00000010",
  51919=>"00000001",
  51920=>"11111111",
  51921=>"00000001",
  51922=>"00000000",
  51923=>"11111111",
  51924=>"00000010",
  51925=>"00000001",
  51926=>"11111110",
  51927=>"00000000",
  51928=>"00000000",
  51929=>"11111110",
  51930=>"00000001",
  51931=>"11111111",
  51932=>"00000001",
  51933=>"00000001",
  51934=>"00000000",
  51935=>"00000000",
  51936=>"00000001",
  51937=>"00000001",
  51938=>"00000001",
  51939=>"00000001",
  51940=>"11111111",
  51941=>"00000010",
  51942=>"00000001",
  51943=>"00000001",
  51944=>"11111111",
  51945=>"11111110",
  51946=>"00000000",
  51947=>"00000010",
  51948=>"11111111",
  51949=>"11111111",
  51950=>"00000001",
  51951=>"00000001",
  51952=>"11111110",
  51953=>"11111111",
  51954=>"00000001",
  51955=>"11111101",
  51956=>"00000001",
  51957=>"00000001",
  51958=>"11111111",
  51959=>"00000001",
  51960=>"00000001",
  51961=>"11111110",
  51962=>"00000001",
  51963=>"00000000",
  51964=>"00000010",
  51965=>"00000000",
  51966=>"00000001",
  51967=>"00000000",
  51968=>"11111111",
  51969=>"00000000",
  51970=>"00000010",
  51971=>"00000000",
  51972=>"00000000",
  51973=>"00000001",
  51974=>"11111110",
  51975=>"00000000",
  51976=>"00000010",
  51977=>"00000001",
  51978=>"00000000",
  51979=>"11111111",
  51980=>"11111111",
  51981=>"11111111",
  51982=>"00000000",
  51983=>"11111111",
  51984=>"11111111",
  51985=>"00000000",
  51986=>"11111111",
  51987=>"11111111",
  51988=>"00000000",
  51989=>"00000000",
  51990=>"00000001",
  51991=>"00000000",
  51992=>"00000000",
  51993=>"00000001",
  51994=>"00000001",
  51995=>"11111111",
  51996=>"00000001",
  51997=>"00000000",
  51998=>"00000001",
  51999=>"11111111",
  52000=>"11111111",
  52001=>"00000001",
  52002=>"00000001",
  52003=>"00000001",
  52004=>"00000000",
  52005=>"00000000",
  52006=>"11111111",
  52007=>"11111111",
  52008=>"00000000",
  52009=>"00000000",
  52010=>"00000000",
  52011=>"00000000",
  52012=>"00000001",
  52013=>"11111110",
  52014=>"00000001",
  52015=>"11111110",
  52016=>"00000000",
  52017=>"00000001",
  52018=>"11111111",
  52019=>"00000001",
  52020=>"11111111",
  52021=>"11111111",
  52022=>"11111110",
  52023=>"00000001",
  52024=>"00000001",
  52025=>"00000010",
  52026=>"11111111",
  52027=>"00000001",
  52028=>"00000000",
  52029=>"00000010",
  52030=>"00000000",
  52031=>"00000000",
  52032=>"00000000",
  52033=>"11111111",
  52034=>"11111111",
  52035=>"11111111",
  52036=>"00000001",
  52037=>"00000000",
  52038=>"00000000",
  52039=>"00000000",
  52040=>"11111111",
  52041=>"00000010",
  52042=>"00000001",
  52043=>"00000001",
  52044=>"00000010",
  52045=>"00000000",
  52046=>"00000011",
  52047=>"11111111",
  52048=>"00000000",
  52049=>"11111111",
  52050=>"11111111",
  52051=>"00000000",
  52052=>"11111101",
  52053=>"11111111",
  52054=>"00000000",
  52055=>"00000000",
  52056=>"00000001",
  52057=>"00000000",
  52058=>"11111111",
  52059=>"11111111",
  52060=>"00000000",
  52061=>"00000001",
  52062=>"11111111",
  52063=>"00000000",
  52064=>"11111111",
  52065=>"00000000",
  52066=>"00000000",
  52067=>"00000010",
  52068=>"11111110",
  52069=>"00000001",
  52070=>"11111111",
  52071=>"11111111",
  52072=>"00000001",
  52073=>"11111110",
  52074=>"11111110",
  52075=>"00000001",
  52076=>"00000000",
  52077=>"00000000",
  52078=>"11111111",
  52079=>"00000000",
  52080=>"11111111",
  52081=>"11111111",
  52082=>"11111111",
  52083=>"00000001",
  52084=>"00000000",
  52085=>"00000001",
  52086=>"11111111",
  52087=>"11111111",
  52088=>"11111111",
  52089=>"00000000",
  52090=>"00000001",
  52091=>"11111111",
  52092=>"11111111",
  52093=>"00000001",
  52094=>"11111111",
  52095=>"11111111",
  52096=>"00000000",
  52097=>"00000000",
  52098=>"11111111",
  52099=>"00000000",
  52100=>"00000000",
  52101=>"00000000",
  52102=>"00000000",
  52103=>"00000000",
  52104=>"00000000",
  52105=>"00000010",
  52106=>"11111111",
  52107=>"11111110",
  52108=>"00000001",
  52109=>"11111111",
  52110=>"00000001",
  52111=>"11111110",
  52112=>"00000001",
  52113=>"11111110",
  52114=>"00000000",
  52115=>"00000010",
  52116=>"11111110",
  52117=>"00000000",
  52118=>"11111110",
  52119=>"00000001",
  52120=>"00000010",
  52121=>"00000001",
  52122=>"00000000",
  52123=>"11111111",
  52124=>"00000000",
  52125=>"00000000",
  52126=>"00000000",
  52127=>"11111110",
  52128=>"00000000",
  52129=>"00000001",
  52130=>"00000000",
  52131=>"11111110",
  52132=>"11111111",
  52133=>"11111111",
  52134=>"11111111",
  52135=>"00000010",
  52136=>"11111111",
  52137=>"00000001",
  52138=>"00000001",
  52139=>"00000010",
  52140=>"00000001",
  52141=>"00000000",
  52142=>"00000001",
  52143=>"11111111",
  52144=>"00000001",
  52145=>"11111111",
  52146=>"11111111",
  52147=>"00000000",
  52148=>"11111110",
  52149=>"11111111",
  52150=>"00000000",
  52151=>"00000001",
  52152=>"11111111",
  52153=>"00000001",
  52154=>"11111110",
  52155=>"00000010",
  52156=>"00000000",
  52157=>"00000000",
  52158=>"00000001",
  52159=>"00000010",
  52160=>"00000000",
  52161=>"00000000",
  52162=>"00000001",
  52163=>"00000001",
  52164=>"00000000",
  52165=>"11111111",
  52166=>"00000000",
  52167=>"00000001",
  52168=>"00000001",
  52169=>"11111111",
  52170=>"00000000",
  52171=>"00000010",
  52172=>"00000001",
  52173=>"00000001",
  52174=>"11111111",
  52175=>"00000001",
  52176=>"11111111",
  52177=>"11111111",
  52178=>"00000000",
  52179=>"11111110",
  52180=>"00000000",
  52181=>"00000000",
  52182=>"11111110",
  52183=>"00000000",
  52184=>"11111111",
  52185=>"11111110",
  52186=>"11111111",
  52187=>"00000000",
  52188=>"00000000",
  52189=>"00000010",
  52190=>"00000001",
  52191=>"00000001",
  52192=>"11111111",
  52193=>"00000001",
  52194=>"00000000",
  52195=>"11111110",
  52196=>"00000000",
  52197=>"00000010",
  52198=>"00000001",
  52199=>"11111110",
  52200=>"11111111",
  52201=>"00000000",
  52202=>"00000010",
  52203=>"11111110",
  52204=>"11111110",
  52205=>"00000010",
  52206=>"00000001",
  52207=>"11111111",
  52208=>"11111110",
  52209=>"11111111",
  52210=>"11111111",
  52211=>"00000000",
  52212=>"00000000",
  52213=>"00000000",
  52214=>"11111111",
  52215=>"11111110",
  52216=>"11111111",
  52217=>"11111111",
  52218=>"00000010",
  52219=>"00000010",
  52220=>"00000000",
  52221=>"00000000",
  52222=>"00000010",
  52223=>"00000000",
  52224=>"00000000",
  52225=>"11111111",
  52226=>"00000000",
  52227=>"11111111",
  52228=>"00000000",
  52229=>"00000000",
  52230=>"00000000",
  52231=>"00000001",
  52232=>"00000010",
  52233=>"00000000",
  52234=>"00000001",
  52235=>"00000010",
  52236=>"11111111",
  52237=>"00000000",
  52238=>"11111111",
  52239=>"00000000",
  52240=>"00000000",
  52241=>"00000000",
  52242=>"00000001",
  52243=>"11111111",
  52244=>"00000001",
  52245=>"11111111",
  52246=>"11111111",
  52247=>"11111110",
  52248=>"00000000",
  52249=>"11111111",
  52250=>"11111110",
  52251=>"00000000",
  52252=>"00000000",
  52253=>"00000010",
  52254=>"11111111",
  52255=>"11111110",
  52256=>"00000000",
  52257=>"00000001",
  52258=>"00000000",
  52259=>"00000001",
  52260=>"11111111",
  52261=>"00000001",
  52262=>"11111111",
  52263=>"11111111",
  52264=>"11111110",
  52265=>"11111111",
  52266=>"00000010",
  52267=>"00000000",
  52268=>"00000001",
  52269=>"11111110",
  52270=>"00000010",
  52271=>"11111111",
  52272=>"00000000",
  52273=>"00000010",
  52274=>"00000000",
  52275=>"11111111",
  52276=>"11111110",
  52277=>"00000000",
  52278=>"11111110",
  52279=>"11111111",
  52280=>"00000000",
  52281=>"00000000",
  52282=>"00000000",
  52283=>"00000000",
  52284=>"11111110",
  52285=>"11111111",
  52286=>"00000000",
  52287=>"11111111",
  52288=>"11111110",
  52289=>"00000000",
  52290=>"00000000",
  52291=>"00000000",
  52292=>"00000001",
  52293=>"00000001",
  52294=>"00000000",
  52295=>"11111111",
  52296=>"11111111",
  52297=>"11111111",
  52298=>"00000001",
  52299=>"00000010",
  52300=>"00000000",
  52301=>"00000000",
  52302=>"11111111",
  52303=>"00000001",
  52304=>"00000000",
  52305=>"00000001",
  52306=>"11111110",
  52307=>"00000000",
  52308=>"00000000",
  52309=>"11111111",
  52310=>"11111110",
  52311=>"11111111",
  52312=>"00000000",
  52313=>"11111111",
  52314=>"00000000",
  52315=>"00000000",
  52316=>"11111111",
  52317=>"00000010",
  52318=>"11111111",
  52319=>"11111111",
  52320=>"00000001",
  52321=>"00000000",
  52322=>"00000000",
  52323=>"00000000",
  52324=>"00000000",
  52325=>"00000001",
  52326=>"00000000",
  52327=>"00000000",
  52328=>"11111111",
  52329=>"11111111",
  52330=>"00000000",
  52331=>"00000000",
  52332=>"11111111",
  52333=>"00000001",
  52334=>"00000000",
  52335=>"00000001",
  52336=>"00000001",
  52337=>"00000000",
  52338=>"00000000",
  52339=>"11111111",
  52340=>"00000010",
  52341=>"00000001",
  52342=>"11111111",
  52343=>"11111111",
  52344=>"00000000",
  52345=>"00000001",
  52346=>"00000001",
  52347=>"11111111",
  52348=>"00000001",
  52349=>"11111111",
  52350=>"11111111",
  52351=>"00000000",
  52352=>"00000000",
  52353=>"00000001",
  52354=>"11111111",
  52355=>"00000010",
  52356=>"00000001",
  52357=>"00000001",
  52358=>"00000000",
  52359=>"00000001",
  52360=>"00000000",
  52361=>"11111111",
  52362=>"00000000",
  52363=>"00000000",
  52364=>"11111111",
  52365=>"11111101",
  52366=>"11111111",
  52367=>"00000001",
  52368=>"00000010",
  52369=>"00000001",
  52370=>"11111110",
  52371=>"00000000",
  52372=>"00000000",
  52373=>"00000000",
  52374=>"00000000",
  52375=>"00000000",
  52376=>"11111111",
  52377=>"00000001",
  52378=>"00000000",
  52379=>"11111110",
  52380=>"00000010",
  52381=>"00000000",
  52382=>"11111111",
  52383=>"11111111",
  52384=>"00000001",
  52385=>"00000000",
  52386=>"11111111",
  52387=>"00000000",
  52388=>"00000000",
  52389=>"00000000",
  52390=>"11111111",
  52391=>"00000001",
  52392=>"11111111",
  52393=>"00000010",
  52394=>"11111111",
  52395=>"11111111",
  52396=>"00000000",
  52397=>"00000001",
  52398=>"11111111",
  52399=>"11111110",
  52400=>"00000001",
  52401=>"11111110",
  52402=>"00000001",
  52403=>"00000000",
  52404=>"00000000",
  52405=>"00000000",
  52406=>"00000001",
  52407=>"00000000",
  52408=>"00000000",
  52409=>"11111111",
  52410=>"00000000",
  52411=>"11111111",
  52412=>"11111110",
  52413=>"11111110",
  52414=>"00000001",
  52415=>"00000000",
  52416=>"00000000",
  52417=>"11111110",
  52418=>"00000001",
  52419=>"00000000",
  52420=>"00000001",
  52421=>"11111110",
  52422=>"00000000",
  52423=>"00000001",
  52424=>"00000000",
  52425=>"00000001",
  52426=>"11111111",
  52427=>"00000001",
  52428=>"00000000",
  52429=>"11111111",
  52430=>"00000010",
  52431=>"00000000",
  52432=>"00000000",
  52433=>"00000001",
  52434=>"00000010",
  52435=>"00000001",
  52436=>"11111111",
  52437=>"00000000",
  52438=>"11111111",
  52439=>"00000001",
  52440=>"11111111",
  52441=>"11111111",
  52442=>"11111111",
  52443=>"11111110",
  52444=>"11111111",
  52445=>"00000010",
  52446=>"00000001",
  52447=>"11111111",
  52448=>"00000010",
  52449=>"00000000",
  52450=>"00000000",
  52451=>"00000001",
  52452=>"00000001",
  52453=>"00000010",
  52454=>"00000001",
  52455=>"00000000",
  52456=>"00000001",
  52457=>"11111111",
  52458=>"11111110",
  52459=>"00000000",
  52460=>"11111111",
  52461=>"00000001",
  52462=>"00000010",
  52463=>"00000001",
  52464=>"00000000",
  52465=>"00000001",
  52466=>"11111111",
  52467=>"11111110",
  52468=>"00000000",
  52469=>"00000010",
  52470=>"00000000",
  52471=>"00000000",
  52472=>"11111110",
  52473=>"11111111",
  52474=>"00000001",
  52475=>"11111111",
  52476=>"11111111",
  52477=>"11111111",
  52478=>"00000001",
  52479=>"11111111",
  52480=>"00000010",
  52481=>"11111111",
  52482=>"00000001",
  52483=>"00000001",
  52484=>"11111110",
  52485=>"00000001",
  52486=>"11111111",
  52487=>"00000001",
  52488=>"00000010",
  52489=>"00000000",
  52490=>"11111111",
  52491=>"00000000",
  52492=>"11111111",
  52493=>"11111111",
  52494=>"11111110",
  52495=>"00000001",
  52496=>"00000001",
  52497=>"00000000",
  52498=>"00000001",
  52499=>"00000000",
  52500=>"11111111",
  52501=>"00000001",
  52502=>"11111111",
  52503=>"00000000",
  52504=>"00000001",
  52505=>"00000010",
  52506=>"00000010",
  52507=>"11111110",
  52508=>"11111111",
  52509=>"00000000",
  52510=>"11111111",
  52511=>"11111111",
  52512=>"11111111",
  52513=>"11111111",
  52514=>"11111110",
  52515=>"00000000",
  52516=>"11111111",
  52517=>"00000000",
  52518=>"00000000",
  52519=>"00000001",
  52520=>"00000000",
  52521=>"00000000",
  52522=>"11111111",
  52523=>"00000001",
  52524=>"00000000",
  52525=>"11111111",
  52526=>"11111111",
  52527=>"00000001",
  52528=>"00000001",
  52529=>"00000000",
  52530=>"11111111",
  52531=>"11111111",
  52532=>"11111111",
  52533=>"11111111",
  52534=>"00000001",
  52535=>"11111111",
  52536=>"11111111",
  52537=>"00000001",
  52538=>"11111110",
  52539=>"00000001",
  52540=>"11111101",
  52541=>"00000000",
  52542=>"11111110",
  52543=>"11111111",
  52544=>"00000000",
  52545=>"11111111",
  52546=>"00000001",
  52547=>"00000000",
  52548=>"11111111",
  52549=>"00000000",
  52550=>"00000000",
  52551=>"00000001",
  52552=>"00000001",
  52553=>"00000001",
  52554=>"00000000",
  52555=>"00000000",
  52556=>"11111111",
  52557=>"11111111",
  52558=>"11111111",
  52559=>"11111111",
  52560=>"00000010",
  52561=>"00000000",
  52562=>"00000000",
  52563=>"00000001",
  52564=>"11111110",
  52565=>"00000000",
  52566=>"11111111",
  52567=>"00000000",
  52568=>"00000001",
  52569=>"11111111",
  52570=>"00000000",
  52571=>"00000010",
  52572=>"00000000",
  52573=>"11111111",
  52574=>"11111111",
  52575=>"11111111",
  52576=>"00000000",
  52577=>"00000000",
  52578=>"00000001",
  52579=>"00000001",
  52580=>"00000000",
  52581=>"00000000",
  52582=>"00000000",
  52583=>"11111111",
  52584=>"00000000",
  52585=>"00000000",
  52586=>"00000010",
  52587=>"00000001",
  52588=>"00000001",
  52589=>"11111111",
  52590=>"00000000",
  52591=>"00000001",
  52592=>"00000001",
  52593=>"11111111",
  52594=>"00000000",
  52595=>"00000000",
  52596=>"00000000",
  52597=>"00000001",
  52598=>"11111111",
  52599=>"00000001",
  52600=>"11111111",
  52601=>"11111111",
  52602=>"11111111",
  52603=>"00000001",
  52604=>"00000001",
  52605=>"00000001",
  52606=>"11111111",
  52607=>"00000000",
  52608=>"00000001",
  52609=>"00000001",
  52610=>"00000010",
  52611=>"00000000",
  52612=>"00000000",
  52613=>"00000000",
  52614=>"00000001",
  52615=>"00000001",
  52616=>"11111110",
  52617=>"00000001",
  52618=>"00000000",
  52619=>"00000100",
  52620=>"11111110",
  52621=>"11111111",
  52622=>"00000001",
  52623=>"00000010",
  52624=>"11111110",
  52625=>"11111111",
  52626=>"00000001",
  52627=>"00000000",
  52628=>"00000001",
  52629=>"00000010",
  52630=>"00000001",
  52631=>"00000001",
  52632=>"00000000",
  52633=>"00000001",
  52634=>"00000001",
  52635=>"00000000",
  52636=>"00000001",
  52637=>"00000001",
  52638=>"00000000",
  52639=>"00000000",
  52640=>"00000000",
  52641=>"00000000",
  52642=>"11111110",
  52643=>"11111111",
  52644=>"00000000",
  52645=>"00000001",
  52646=>"00000001",
  52647=>"00000000",
  52648=>"00000001",
  52649=>"00000000",
  52650=>"00000000",
  52651=>"00000001",
  52652=>"00000000",
  52653=>"11111110",
  52654=>"00000000",
  52655=>"00000000",
  52656=>"00000000",
  52657=>"11111111",
  52658=>"11111110",
  52659=>"11111111",
  52660=>"11111111",
  52661=>"00000000",
  52662=>"11111110",
  52663=>"00000001",
  52664=>"00000000",
  52665=>"00000001",
  52666=>"11111111",
  52667=>"11111111",
  52668=>"00000000",
  52669=>"00000001",
  52670=>"00000001",
  52671=>"11111110",
  52672=>"00000000",
  52673=>"00000001",
  52674=>"11111111",
  52675=>"00000000",
  52676=>"00000001",
  52677=>"11111110",
  52678=>"11111111",
  52679=>"00000000",
  52680=>"00000000",
  52681=>"00000001",
  52682=>"00000000",
  52683=>"11111110",
  52684=>"00000000",
  52685=>"11111111",
  52686=>"00000000",
  52687=>"00000010",
  52688=>"11111111",
  52689=>"00000000",
  52690=>"00000001",
  52691=>"00000000",
  52692=>"00000000",
  52693=>"00000000",
  52694=>"00000001",
  52695=>"11111111",
  52696=>"00000001",
  52697=>"00000000",
  52698=>"00000001",
  52699=>"00000010",
  52700=>"00000001",
  52701=>"00000000",
  52702=>"11111111",
  52703=>"11111111",
  52704=>"00000000",
  52705=>"11111111",
  52706=>"00000011",
  52707=>"11111101",
  52708=>"11111110",
  52709=>"11111111",
  52710=>"00000000",
  52711=>"00000001",
  52712=>"00000001",
  52713=>"11111101",
  52714=>"00000001",
  52715=>"00000000",
  52716=>"11111110",
  52717=>"00000000",
  52718=>"11111111",
  52719=>"00000000",
  52720=>"11111111",
  52721=>"11111111",
  52722=>"11111111",
  52723=>"00000001",
  52724=>"00000010",
  52725=>"00000010",
  52726=>"00000001",
  52727=>"00000000",
  52728=>"00000001",
  52729=>"00000000",
  52730=>"00000000",
  52731=>"00000001",
  52732=>"00000001",
  52733=>"00000000",
  52734=>"00000001",
  52735=>"00000000",
  52736=>"00000010",
  52737=>"00000001",
  52738=>"11111111",
  52739=>"11111111",
  52740=>"00000001",
  52741=>"11111110",
  52742=>"11111111",
  52743=>"00000000",
  52744=>"11111110",
  52745=>"00000001",
  52746=>"00000001",
  52747=>"11111111",
  52748=>"00000000",
  52749=>"00000001",
  52750=>"00000000",
  52751=>"00000000",
  52752=>"11111111",
  52753=>"00000001",
  52754=>"11111111",
  52755=>"11111111",
  52756=>"00000000",
  52757=>"11111111",
  52758=>"00000001",
  52759=>"00000000",
  52760=>"00000001",
  52761=>"00000000",
  52762=>"11111111",
  52763=>"00000001",
  52764=>"00000001",
  52765=>"00000001",
  52766=>"11111111",
  52767=>"00000001",
  52768=>"00000001",
  52769=>"00000001",
  52770=>"00000000",
  52771=>"00000000",
  52772=>"00000001",
  52773=>"00000001",
  52774=>"11111110",
  52775=>"00000001",
  52776=>"00000001",
  52777=>"00000001",
  52778=>"00000001",
  52779=>"00000000",
  52780=>"00000001",
  52781=>"00000000",
  52782=>"11111110",
  52783=>"00000010",
  52784=>"00000000",
  52785=>"00000000",
  52786=>"11111110",
  52787=>"11111111",
  52788=>"00000001",
  52789=>"00000000",
  52790=>"00000001",
  52791=>"00000001",
  52792=>"00000001",
  52793=>"00000010",
  52794=>"00000001",
  52795=>"00000000",
  52796=>"00000001",
  52797=>"11111110",
  52798=>"11111111",
  52799=>"00000001",
  52800=>"00000001",
  52801=>"11111110",
  52802=>"00000000",
  52803=>"00000000",
  52804=>"00000001",
  52805=>"00000000",
  52806=>"11111111",
  52807=>"00000001",
  52808=>"11111111",
  52809=>"11111111",
  52810=>"11111110",
  52811=>"11111111",
  52812=>"00000000",
  52813=>"11111111",
  52814=>"11111111",
  52815=>"00000010",
  52816=>"00000001",
  52817=>"11111111",
  52818=>"11111110",
  52819=>"00000000",
  52820=>"00000001",
  52821=>"00000001",
  52822=>"11111111",
  52823=>"00000001",
  52824=>"00000010",
  52825=>"11111110",
  52826=>"00000000",
  52827=>"00000000",
  52828=>"11111110",
  52829=>"11111110",
  52830=>"00000000",
  52831=>"00000001",
  52832=>"00000001",
  52833=>"00000001",
  52834=>"11111111",
  52835=>"00000000",
  52836=>"11111110",
  52837=>"11111111",
  52838=>"00000000",
  52839=>"00000000",
  52840=>"11111111",
  52841=>"00000000",
  52842=>"00000000",
  52843=>"00000001",
  52844=>"00000000",
  52845=>"00000001",
  52846=>"00000001",
  52847=>"11111111",
  52848=>"00000001",
  52849=>"11111111",
  52850=>"00000000",
  52851=>"00000001",
  52852=>"00000001",
  52853=>"00000001",
  52854=>"00000001",
  52855=>"00000000",
  52856=>"00000010",
  52857=>"11111111",
  52858=>"11111111",
  52859=>"11111110",
  52860=>"11111110",
  52861=>"00000010",
  52862=>"00000001",
  52863=>"00000001",
  52864=>"00000010",
  52865=>"00000001",
  52866=>"00000000",
  52867=>"00000000",
  52868=>"11111111",
  52869=>"11111111",
  52870=>"00000001",
  52871=>"11111111",
  52872=>"00000000",
  52873=>"11111111",
  52874=>"11111111",
  52875=>"00000000",
  52876=>"11111101",
  52877=>"00000010",
  52878=>"00000000",
  52879=>"11111110",
  52880=>"11111110",
  52881=>"11111111",
  52882=>"00000001",
  52883=>"00000010",
  52884=>"00000010",
  52885=>"00000001",
  52886=>"00000000",
  52887=>"00000001",
  52888=>"00000010",
  52889=>"11111111",
  52890=>"00000001",
  52891=>"00000010",
  52892=>"11111111",
  52893=>"00000001",
  52894=>"00000001",
  52895=>"00000000",
  52896=>"00000000",
  52897=>"11111111",
  52898=>"11111111",
  52899=>"00000000",
  52900=>"00000000",
  52901=>"11111111",
  52902=>"00000001",
  52903=>"00000000",
  52904=>"00000000",
  52905=>"00000001",
  52906=>"00000000",
  52907=>"00000000",
  52908=>"00000010",
  52909=>"00000001",
  52910=>"00000010",
  52911=>"00000001",
  52912=>"00000001",
  52913=>"00000001",
  52914=>"00000010",
  52915=>"00000001",
  52916=>"00000000",
  52917=>"00000000",
  52918=>"00000001",
  52919=>"00000000",
  52920=>"00000001",
  52921=>"00000001",
  52922=>"11111110",
  52923=>"00000010",
  52924=>"00000000",
  52925=>"00000001",
  52926=>"00000000",
  52927=>"11111110",
  52928=>"11111111",
  52929=>"00000001",
  52930=>"00000000",
  52931=>"00000001",
  52932=>"11111110",
  52933=>"00000000",
  52934=>"11111111",
  52935=>"00000000",
  52936=>"11111111",
  52937=>"00000001",
  52938=>"11111111",
  52939=>"11111111",
  52940=>"11111111",
  52941=>"00000000",
  52942=>"11111111",
  52943=>"11111111",
  52944=>"11111110",
  52945=>"11111111",
  52946=>"11111110",
  52947=>"00000000",
  52948=>"00000001",
  52949=>"00000001",
  52950=>"00000001",
  52951=>"00000001",
  52952=>"00000000",
  52953=>"00000000",
  52954=>"00000000",
  52955=>"00000000",
  52956=>"00000000",
  52957=>"11111110",
  52958=>"11111111",
  52959=>"11111111",
  52960=>"00000001",
  52961=>"00000001",
  52962=>"00000001",
  52963=>"11111111",
  52964=>"11111111",
  52965=>"00000001",
  52966=>"00000001",
  52967=>"00000000",
  52968=>"00000000",
  52969=>"11111111",
  52970=>"11111111",
  52971=>"00000000",
  52972=>"00000000",
  52973=>"11111111",
  52974=>"00000001",
  52975=>"00000000",
  52976=>"00000001",
  52977=>"00000001",
  52978=>"11111110",
  52979=>"00000000",
  52980=>"00000001",
  52981=>"00000000",
  52982=>"00000010",
  52983=>"11111111",
  52984=>"00000000",
  52985=>"00000001",
  52986=>"00000000",
  52987=>"11111111",
  52988=>"00000000",
  52989=>"00000001",
  52990=>"11111111",
  52991=>"00000000",
  52992=>"00000000",
  52993=>"11111110",
  52994=>"11111111",
  52995=>"11111110",
  52996=>"00000001",
  52997=>"00000000",
  52998=>"00000000",
  52999=>"00000000",
  53000=>"00000001",
  53001=>"00000001",
  53002=>"11111111",
  53003=>"11111111",
  53004=>"11111111",
  53005=>"00000001",
  53006=>"11111111",
  53007=>"00000010",
  53008=>"00000000",
  53009=>"11111111",
  53010=>"11111111",
  53011=>"00000000",
  53012=>"00000001",
  53013=>"11111111",
  53014=>"00000001",
  53015=>"00000000",
  53016=>"00000000",
  53017=>"11111111",
  53018=>"11111111",
  53019=>"11111111",
  53020=>"00000000",
  53021=>"00000000",
  53022=>"00000000",
  53023=>"00000010",
  53024=>"11111110",
  53025=>"11111111",
  53026=>"00000001",
  53027=>"11111111",
  53028=>"00000001",
  53029=>"00000000",
  53030=>"00000000",
  53031=>"00000000",
  53032=>"00000000",
  53033=>"00000001",
  53034=>"11111110",
  53035=>"00000001",
  53036=>"00000000",
  53037=>"11111110",
  53038=>"11111111",
  53039=>"00000000",
  53040=>"00000000",
  53041=>"00000001",
  53042=>"11111111",
  53043=>"11111111",
  53044=>"11111110",
  53045=>"00000001",
  53046=>"00000000",
  53047=>"00000001",
  53048=>"00000000",
  53049=>"00000010",
  53050=>"00000010",
  53051=>"00000000",
  53052=>"11111111",
  53053=>"00000001",
  53054=>"11111111",
  53055=>"00000001",
  53056=>"00000001",
  53057=>"11111111",
  53058=>"00000000",
  53059=>"00000000",
  53060=>"00000001",
  53061=>"11111111",
  53062=>"11111111",
  53063=>"00000000",
  53064=>"11111111",
  53065=>"11111110",
  53066=>"11111110",
  53067=>"00000001",
  53068=>"11111111",
  53069=>"00000001",
  53070=>"00000000",
  53071=>"00000000",
  53072=>"00000000",
  53073=>"00000000",
  53074=>"00000010",
  53075=>"00000001",
  53076=>"11111111",
  53077=>"00000000",
  53078=>"11111110",
  53079=>"00000001",
  53080=>"11111111",
  53081=>"00000000",
  53082=>"11111111",
  53083=>"11111111",
  53084=>"00000001",
  53085=>"00000000",
  53086=>"11111111",
  53087=>"00000001",
  53088=>"00000000",
  53089=>"00000001",
  53090=>"00000000",
  53091=>"00000001",
  53092=>"00000010",
  53093=>"11111111",
  53094=>"11111110",
  53095=>"11111110",
  53096=>"00000000",
  53097=>"00000000",
  53098=>"11111110",
  53099=>"00000010",
  53100=>"11111110",
  53101=>"00000000",
  53102=>"00000001",
  53103=>"00000001",
  53104=>"00000001",
  53105=>"00000000",
  53106=>"00000000",
  53107=>"11111111",
  53108=>"00000001",
  53109=>"11111111",
  53110=>"00000001",
  53111=>"00000001",
  53112=>"00000000",
  53113=>"00000001",
  53114=>"00000000",
  53115=>"11111111",
  53116=>"11111111",
  53117=>"00000001",
  53118=>"11111111",
  53119=>"00000010",
  53120=>"00000000",
  53121=>"00000000",
  53122=>"00000001",
  53123=>"11111111",
  53124=>"00000001",
  53125=>"00000001",
  53126=>"11111111",
  53127=>"11111111",
  53128=>"11111110",
  53129=>"11111111",
  53130=>"11111110",
  53131=>"11111111",
  53132=>"00000001",
  53133=>"11111111",
  53134=>"00000010",
  53135=>"00000001",
  53136=>"11111111",
  53137=>"00000001",
  53138=>"11111110",
  53139=>"11111110",
  53140=>"00000000",
  53141=>"00000001",
  53142=>"00000001",
  53143=>"00000001",
  53144=>"00000000",
  53145=>"00000000",
  53146=>"11111111",
  53147=>"00000001",
  53148=>"11111111",
  53149=>"00000000",
  53150=>"00000001",
  53151=>"00000000",
  53152=>"00000001",
  53153=>"00000000",
  53154=>"00000001",
  53155=>"00000000",
  53156=>"11111111",
  53157=>"11111111",
  53158=>"00000001",
  53159=>"11111111",
  53160=>"00000000",
  53161=>"00000001",
  53162=>"11111111",
  53163=>"00000000",
  53164=>"00000001",
  53165=>"11111111",
  53166=>"11111111",
  53167=>"00000001",
  53168=>"00000001",
  53169=>"11111110",
  53170=>"00000001",
  53171=>"11111111",
  53172=>"11111110",
  53173=>"00000001",
  53174=>"11111111",
  53175=>"00000001",
  53176=>"11111110",
  53177=>"00000000",
  53178=>"00000000",
  53179=>"11111111",
  53180=>"11111110",
  53181=>"11111111",
  53182=>"00000000",
  53183=>"00000010",
  53184=>"00000001",
  53185=>"11111111",
  53186=>"00000001",
  53187=>"00000001",
  53188=>"00000000",
  53189=>"00000000",
  53190=>"11111111",
  53191=>"11111110",
  53192=>"00000000",
  53193=>"00000001",
  53194=>"00000000",
  53195=>"11111111",
  53196=>"00000010",
  53197=>"00000010",
  53198=>"11111110",
  53199=>"00000000",
  53200=>"11111101",
  53201=>"00000001",
  53202=>"11111111",
  53203=>"11111111",
  53204=>"00000000",
  53205=>"11111111",
  53206=>"00000001",
  53207=>"00000001",
  53208=>"00000001",
  53209=>"11111111",
  53210=>"11111111",
  53211=>"00000001",
  53212=>"11111111",
  53213=>"00000001",
  53214=>"00000010",
  53215=>"00000000",
  53216=>"11111111",
  53217=>"00000000",
  53218=>"00000000",
  53219=>"00000000",
  53220=>"11111110",
  53221=>"00000001",
  53222=>"00000000",
  53223=>"00000000",
  53224=>"11111111",
  53225=>"11111110",
  53226=>"00000000",
  53227=>"00000000",
  53228=>"00000010",
  53229=>"00000000",
  53230=>"00000001",
  53231=>"00000000",
  53232=>"00000000",
  53233=>"00000001",
  53234=>"11111111",
  53235=>"11111111",
  53236=>"00000000",
  53237=>"11111110",
  53238=>"00000000",
  53239=>"11111110",
  53240=>"00000000",
  53241=>"11111111",
  53242=>"11111111",
  53243=>"11111110",
  53244=>"00000001",
  53245=>"11111111",
  53246=>"00000001",
  53247=>"00000010",
  53248=>"00000000",
  53249=>"00000000",
  53250=>"00000000",
  53251=>"00000000",
  53252=>"00000000",
  53253=>"00000000",
  53254=>"11111111",
  53255=>"00000000",
  53256=>"00000000",
  53257=>"00000000",
  53258=>"00000000",
  53259=>"00000000",
  53260=>"00000000",
  53261=>"00000000",
  53262=>"00000000",
  53263=>"00000000",
  53264=>"00000000",
  53265=>"00000000",
  53266=>"00000000",
  53267=>"00000000",
  53268=>"00000000",
  53269=>"00000000",
  53270=>"00000000",
  53271=>"00000000",
  53272=>"00000000",
  53273=>"00000000",
  53274=>"00000000",
  53275=>"00000000",
  53276=>"00000001",
  53277=>"00000000",
  53278=>"00000000",
  53279=>"00000000",
  53280=>"00000000",
  53281=>"00000000",
  53282=>"00000000",
  53283=>"00000000",
  53284=>"00000000",
  53285=>"00000001",
  53286=>"00000001",
  53287=>"00000000",
  53288=>"00000000",
  53289=>"00000000",
  53290=>"00000000",
  53291=>"00000000",
  53292=>"00000000",
  53293=>"00000000",
  53294=>"00000000",
  53295=>"00000000",
  53296=>"00000000",
  53297=>"00000000",
  53298=>"00000000",
  53299=>"00000000",
  53300=>"00000000",
  53301=>"00000000",
  53302=>"00000000",
  53303=>"00000000",
  53304=>"00000000",
  53305=>"00000000",
  53306=>"00000000",
  53307=>"00000000",
  53308=>"00000000",
  53309=>"00000000",
  53310=>"00000000",
  53311=>"00000001",
  53312=>"00000000",
  53313=>"00000000",
  53314=>"00000000",
  53315=>"00000001",
  53316=>"00000000",
  53317=>"11111111",
  53318=>"00000000",
  53319=>"00000000",
  53320=>"00000000",
  53321=>"00000000",
  53322=>"00000000",
  53323=>"00000000",
  53324=>"00000000",
  53325=>"00000000",
  53326=>"00000000",
  53327=>"00000000",
  53328=>"00000000",
  53329=>"00000000",
  53330=>"00000000",
  53331=>"00000000",
  53332=>"00000000",
  53333=>"00000000",
  53334=>"00000000",
  53335=>"00000000",
  53336=>"00000000",
  53337=>"00000000",
  53338=>"00000000",
  53339=>"00000000",
  53340=>"00000000",
  53341=>"11111111",
  53342=>"00000000",
  53343=>"00000000",
  53344=>"00000000",
  53345=>"00000000",
  53346=>"00000000",
  53347=>"00000000",
  53348=>"00000000",
  53349=>"00000000",
  53350=>"00000000",
  53351=>"11111111",
  53352=>"00000000",
  53353=>"00000001",
  53354=>"00000000",
  53355=>"00000000",
  53356=>"00000000",
  53357=>"00000000",
  53358=>"00000000",
  53359=>"00000000",
  53360=>"00000000",
  53361=>"00000000",
  53362=>"00000000",
  53363=>"00000000",
  53364=>"00000000",
  53365=>"00000000",
  53366=>"00000000",
  53367=>"00000000",
  53368=>"00000000",
  53369=>"00000000",
  53370=>"00000000",
  53371=>"00000000",
  53372=>"00000000",
  53373=>"00000000",
  53374=>"00000001",
  53375=>"00000000",
  53376=>"00000000",
  53377=>"00000000",
  53378=>"00000000",
  53379=>"11111111",
  53380=>"00000000",
  53381=>"00000000",
  53382=>"00000001",
  53383=>"00000000",
  53384=>"00000000",
  53385=>"00000000",
  53386=>"00000001",
  53387=>"00000000",
  53388=>"00000000",
  53389=>"00000000",
  53390=>"00000000",
  53391=>"00000000",
  53392=>"00000000",
  53393=>"00000000",
  53394=>"00000000",
  53395=>"00000000",
  53396=>"00000000",
  53397=>"00000000",
  53398=>"00000000",
  53399=>"00000000",
  53400=>"00000000",
  53401=>"00000000",
  53402=>"00000000",
  53403=>"00000000",
  53404=>"00000001",
  53405=>"00000000",
  53406=>"00000000",
  53407=>"00000000",
  53408=>"00000000",
  53409=>"00000000",
  53410=>"11111111",
  53411=>"00000000",
  53412=>"00000000",
  53413=>"00000000",
  53414=>"00000000",
  53415=>"00000001",
  53416=>"00000000",
  53417=>"00000000",
  53418=>"00000000",
  53419=>"00000000",
  53420=>"00000000",
  53421=>"00000000",
  53422=>"00000000",
  53423=>"00000000",
  53424=>"00000000",
  53425=>"00000000",
  53426=>"11111111",
  53427=>"00000000",
  53428=>"00000000",
  53429=>"00000000",
  53430=>"00000000",
  53431=>"00000000",
  53432=>"00000000",
  53433=>"00000000",
  53434=>"00000000",
  53435=>"00000000",
  53436=>"00000000",
  53437=>"00000000",
  53438=>"00000000",
  53439=>"00000000",
  53440=>"00000000",
  53441=>"11111111",
  53442=>"00000000",
  53443=>"00000000",
  53444=>"11111111",
  53445=>"00000000",
  53446=>"00000000",
  53447=>"00000000",
  53448=>"00000000",
  53449=>"00000000",
  53450=>"11111111",
  53451=>"00000000",
  53452=>"00000000",
  53453=>"00000000",
  53454=>"11111111",
  53455=>"00000000",
  53456=>"00000000",
  53457=>"00000000",
  53458=>"11111100",
  53459=>"00000001",
  53460=>"00000000",
  53461=>"00000000",
  53462=>"00000001",
  53463=>"00000000",
  53464=>"00000000",
  53465=>"00000000",
  53466=>"00000001",
  53467=>"00000000",
  53468=>"00000000",
  53469=>"00000000",
  53470=>"00000000",
  53471=>"11111111",
  53472=>"00000001",
  53473=>"00000000",
  53474=>"00000000",
  53475=>"00000001",
  53476=>"11111111",
  53477=>"00000000",
  53478=>"00000000",
  53479=>"00000000",
  53480=>"00000000",
  53481=>"00000000",
  53482=>"00000001",
  53483=>"11111111",
  53484=>"00000000",
  53485=>"00000000",
  53486=>"00000000",
  53487=>"11111111",
  53488=>"00000000",
  53489=>"00000000",
  53490=>"00000000",
  53491=>"11111111",
  53492=>"00000000",
  53493=>"00000000",
  53494=>"00000000",
  53495=>"00000000",
  53496=>"00000000",
  53497=>"11111111",
  53498=>"00000001",
  53499=>"11111111",
  53500=>"00000001",
  53501=>"00000000",
  53502=>"00000000",
  53503=>"00000000",
  53504=>"00000000",
  53505=>"00000000",
  53506=>"00000000",
  53507=>"11111111",
  53508=>"11111111",
  53509=>"00000000",
  53510=>"00000000",
  53511=>"00000000",
  53512=>"00000000",
  53513=>"00000000",
  53514=>"00000000",
  53515=>"00000000",
  53516=>"00000000",
  53517=>"00000000",
  53518=>"00000000",
  53519=>"00000000",
  53520=>"00000000",
  53521=>"00000000",
  53522=>"00000000",
  53523=>"00000000",
  53524=>"00000000",
  53525=>"00000000",
  53526=>"00000000",
  53527=>"00000000",
  53528=>"00000000",
  53529=>"11111111",
  53530=>"11111111",
  53531=>"11111111",
  53532=>"00000000",
  53533=>"00000000",
  53534=>"00000000",
  53535=>"00000000",
  53536=>"00000000",
  53537=>"00000000",
  53538=>"00000001",
  53539=>"00000000",
  53540=>"00000000",
  53541=>"00000000",
  53542=>"00000000",
  53543=>"00000000",
  53544=>"00000000",
  53545=>"00000000",
  53546=>"00000000",
  53547=>"00000000",
  53548=>"00000000",
  53549=>"11111111",
  53550=>"00000000",
  53551=>"00000000",
  53552=>"11111101",
  53553=>"00000000",
  53554=>"00000000",
  53555=>"00000000",
  53556=>"00000000",
  53557=>"00000000",
  53558=>"00000000",
  53559=>"11111111",
  53560=>"00000000",
  53561=>"00000000",
  53562=>"00000000",
  53563=>"00000000",
  53564=>"00000000",
  53565=>"11111111",
  53566=>"00000000",
  53567=>"00000000",
  53568=>"00000000",
  53569=>"00000000",
  53570=>"00000000",
  53571=>"00000000",
  53572=>"11111111",
  53573=>"00000000",
  53574=>"00000000",
  53575=>"00000000",
  53576=>"00000000",
  53577=>"00000000",
  53578=>"00000000",
  53579=>"00000000",
  53580=>"00000000",
  53581=>"00000000",
  53582=>"00000000",
  53583=>"00000000",
  53584=>"00000000",
  53585=>"00000000",
  53586=>"00000000",
  53587=>"00000000",
  53588=>"00000001",
  53589=>"00000000",
  53590=>"00000000",
  53591=>"00000000",
  53592=>"00000000",
  53593=>"00000000",
  53594=>"00000001",
  53595=>"00000000",
  53596=>"00000000",
  53597=>"00000001",
  53598=>"00000000",
  53599=>"00000000",
  53600=>"00000000",
  53601=>"00000000",
  53602=>"00000000",
  53603=>"00000000",
  53604=>"00000000",
  53605=>"00000000",
  53606=>"00000001",
  53607=>"00000000",
  53608=>"11111111",
  53609=>"00000000",
  53610=>"00000000",
  53611=>"00000000",
  53612=>"00000000",
  53613=>"00000000",
  53614=>"00000000",
  53615=>"00000000",
  53616=>"00000000",
  53617=>"00000000",
  53618=>"00000000",
  53619=>"00000000",
  53620=>"00000000",
  53621=>"00000000",
  53622=>"00000000",
  53623=>"00000000",
  53624=>"00000000",
  53625=>"00000000",
  53626=>"00000000",
  53627=>"00000000",
  53628=>"00000000",
  53629=>"00000000",
  53630=>"00000000",
  53631=>"00000000",
  53632=>"00000000",
  53633=>"00000000",
  53634=>"00000000",
  53635=>"11111111",
  53636=>"00000001",
  53637=>"00000000",
  53638=>"00000000",
  53639=>"00000000",
  53640=>"00000000",
  53641=>"00000000",
  53642=>"00000000",
  53643=>"00000000",
  53644=>"00000000",
  53645=>"00000001",
  53646=>"00000000",
  53647=>"00000000",
  53648=>"11111111",
  53649=>"00000000",
  53650=>"00000000",
  53651=>"00000000",
  53652=>"00000000",
  53653=>"00000000",
  53654=>"00000000",
  53655=>"00000000",
  53656=>"00000000",
  53657=>"00000000",
  53658=>"00000000",
  53659=>"00000000",
  53660=>"00000000",
  53661=>"00000000",
  53662=>"00000000",
  53663=>"00000000",
  53664=>"00000000",
  53665=>"00000000",
  53666=>"00000000",
  53667=>"00000000",
  53668=>"00000000",
  53669=>"00000001",
  53670=>"00000000",
  53671=>"00000000",
  53672=>"00000000",
  53673=>"00000000",
  53674=>"00000000",
  53675=>"00000000",
  53676=>"11111111",
  53677=>"00000000",
  53678=>"00000000",
  53679=>"00000000",
  53680=>"00000000",
  53681=>"00000000",
  53682=>"00000000",
  53683=>"00000000",
  53684=>"00000000",
  53685=>"00000000",
  53686=>"00000000",
  53687=>"00000000",
  53688=>"00000000",
  53689=>"00000000",
  53690=>"11111111",
  53691=>"00000000",
  53692=>"00000000",
  53693=>"00000000",
  53694=>"00000000",
  53695=>"00000000",
  53696=>"00000000",
  53697=>"00000000",
  53698=>"00000000",
  53699=>"00000000",
  53700=>"00000000",
  53701=>"00000000",
  53702=>"00000000",
  53703=>"00000000",
  53704=>"00000000",
  53705=>"00000000",
  53706=>"00000000",
  53707=>"00000000",
  53708=>"00000000",
  53709=>"00000000",
  53710=>"00000000",
  53711=>"00000000",
  53712=>"00000000",
  53713=>"00000000",
  53714=>"00000000",
  53715=>"00000000",
  53716=>"00000000",
  53717=>"00000000",
  53718=>"00000000",
  53719=>"00000000",
  53720=>"00000000",
  53721=>"00000000",
  53722=>"00000000",
  53723=>"00000000",
  53724=>"00000000",
  53725=>"00000000",
  53726=>"00000000",
  53727=>"00000000",
  53728=>"00000000",
  53729=>"11111111",
  53730=>"00000000",
  53731=>"11111111",
  53732=>"00000000",
  53733=>"00000000",
  53734=>"00000000",
  53735=>"00000000",
  53736=>"00000000",
  53737=>"00000000",
  53738=>"00000000",
  53739=>"00000000",
  53740=>"00000001",
  53741=>"00000000",
  53742=>"00000000",
  53743=>"00000000",
  53744=>"00000000",
  53745=>"00000000",
  53746=>"00000000",
  53747=>"00000000",
  53748=>"00000000",
  53749=>"00000000",
  53750=>"00000000",
  53751=>"00000001",
  53752=>"00000000",
  53753=>"00000000",
  53754=>"00000000",
  53755=>"00000000",
  53756=>"11111111",
  53757=>"00000000",
  53758=>"00000000",
  53759=>"00000000",
  53760=>"00000001",
  53761=>"00000001",
  53762=>"00000000",
  53763=>"00000000",
  53764=>"00000000",
  53765=>"00000000",
  53766=>"00000000",
  53767=>"00000000",
  53768=>"00000000",
  53769=>"00000000",
  53770=>"00000000",
  53771=>"00000000",
  53772=>"00000000",
  53773=>"00000000",
  53774=>"00000000",
  53775=>"00000000",
  53776=>"00000000",
  53777=>"00000000",
  53778=>"00000000",
  53779=>"00000000",
  53780=>"00000000",
  53781=>"00000000",
  53782=>"11111111",
  53783=>"00000000",
  53784=>"00000000",
  53785=>"00000000",
  53786=>"00000000",
  53787=>"00000000",
  53788=>"11111111",
  53789=>"00000000",
  53790=>"11111111",
  53791=>"00000000",
  53792=>"00000000",
  53793=>"00000000",
  53794=>"11111111",
  53795=>"00000000",
  53796=>"00000000",
  53797=>"00000000",
  53798=>"00000000",
  53799=>"00000000",
  53800=>"00000000",
  53801=>"00000000",
  53802=>"00000000",
  53803=>"00000000",
  53804=>"00000000",
  53805=>"00000000",
  53806=>"00000000",
  53807=>"11111111",
  53808=>"00000000",
  53809=>"00000000",
  53810=>"00000000",
  53811=>"11111111",
  53812=>"00000000",
  53813=>"00000000",
  53814=>"00000000",
  53815=>"00000000",
  53816=>"00000001",
  53817=>"11111111",
  53818=>"00000000",
  53819=>"11111111",
  53820=>"11111111",
  53821=>"00000000",
  53822=>"00000000",
  53823=>"00000000",
  53824=>"00000000",
  53825=>"00000000",
  53826=>"00000000",
  53827=>"00000000",
  53828=>"00000000",
  53829=>"00000000",
  53830=>"00000000",
  53831=>"00000000",
  53832=>"00000000",
  53833=>"00000000",
  53834=>"00000000",
  53835=>"00000000",
  53836=>"00000000",
  53837=>"00000000",
  53838=>"00000000",
  53839=>"00000000",
  53840=>"00000000",
  53841=>"00000000",
  53842=>"00000000",
  53843=>"00000000",
  53844=>"00000000",
  53845=>"00000000",
  53846=>"00000000",
  53847=>"00000000",
  53848=>"00000000",
  53849=>"00000000",
  53850=>"00000001",
  53851=>"00000000",
  53852=>"00000000",
  53853=>"00000000",
  53854=>"00000000",
  53855=>"00000000",
  53856=>"00000000",
  53857=>"00000000",
  53858=>"00000001",
  53859=>"00000000",
  53860=>"11111111",
  53861=>"00000000",
  53862=>"00000000",
  53863=>"00000000",
  53864=>"00000000",
  53865=>"00000000",
  53866=>"00000000",
  53867=>"00000000",
  53868=>"11111111",
  53869=>"00000000",
  53870=>"00000000",
  53871=>"00000000",
  53872=>"00000001",
  53873=>"00000000",
  53874=>"00000000",
  53875=>"00000000",
  53876=>"00000000",
  53877=>"00000000",
  53878=>"00000000",
  53879=>"00000000",
  53880=>"00000000",
  53881=>"11111111",
  53882=>"00000000",
  53883=>"00000000",
  53884=>"00000000",
  53885=>"00000000",
  53886=>"00000000",
  53887=>"00000000",
  53888=>"00000000",
  53889=>"00000000",
  53890=>"00000000",
  53891=>"00000000",
  53892=>"00000000",
  53893=>"00000000",
  53894=>"00000000",
  53895=>"11111111",
  53896=>"00000000",
  53897=>"00000000",
  53898=>"00000000",
  53899=>"00000000",
  53900=>"00000000",
  53901=>"00000000",
  53902=>"00000001",
  53903=>"00000000",
  53904=>"00000000",
  53905=>"00000000",
  53906=>"00000000",
  53907=>"00000000",
  53908=>"00000000",
  53909=>"00000000",
  53910=>"00000000",
  53911=>"00000000",
  53912=>"00000001",
  53913=>"00000000",
  53914=>"00000000",
  53915=>"00000000",
  53916=>"00000000",
  53917=>"00000000",
  53918=>"11111111",
  53919=>"00000000",
  53920=>"11111111",
  53921=>"00000000",
  53922=>"00000000",
  53923=>"00000000",
  53924=>"00000000",
  53925=>"00000000",
  53926=>"00000000",
  53927=>"00000000",
  53928=>"00000000",
  53929=>"00000000",
  53930=>"00000000",
  53931=>"00000000",
  53932=>"11111111",
  53933=>"00000000",
  53934=>"00000000",
  53935=>"00000000",
  53936=>"00000000",
  53937=>"00000000",
  53938=>"00000000",
  53939=>"11111111",
  53940=>"00000000",
  53941=>"00000000",
  53942=>"11111111",
  53943=>"00000000",
  53944=>"00000000",
  53945=>"00000000",
  53946=>"00000000",
  53947=>"00000000",
  53948=>"00000000",
  53949=>"00000000",
  53950=>"00000000",
  53951=>"00000000",
  53952=>"00000000",
  53953=>"00000000",
  53954=>"00000000",
  53955=>"11111111",
  53956=>"00000000",
  53957=>"00000000",
  53958=>"00000000",
  53959=>"11111111",
  53960=>"00000000",
  53961=>"00000000",
  53962=>"00000000",
  53963=>"00000000",
  53964=>"00000000",
  53965=>"00000000",
  53966=>"00000001",
  53967=>"11111111",
  53968=>"00000000",
  53969=>"00000000",
  53970=>"00000000",
  53971=>"00000000",
  53972=>"00000000",
  53973=>"00000000",
  53974=>"11111111",
  53975=>"00000000",
  53976=>"00000000",
  53977=>"00000000",
  53978=>"00000000",
  53979=>"00000000",
  53980=>"00000000",
  53981=>"11111101",
  53982=>"00000000",
  53983=>"00000000",
  53984=>"00000000",
  53985=>"00000000",
  53986=>"00000001",
  53987=>"00000001",
  53988=>"00000000",
  53989=>"00000000",
  53990=>"00000000",
  53991=>"00000000",
  53992=>"00000000",
  53993=>"00000000",
  53994=>"00000000",
  53995=>"00000000",
  53996=>"00000000",
  53997=>"00000000",
  53998=>"00000000",
  53999=>"00000000",
  54000=>"00000000",
  54001=>"00000000",
  54002=>"00000000",
  54003=>"00000000",
  54004=>"00000000",
  54005=>"00000000",
  54006=>"00000000",
  54007=>"00000000",
  54008=>"00000000",
  54009=>"00000000",
  54010=>"00000000",
  54011=>"00000000",
  54012=>"11111111",
  54013=>"00000000",
  54014=>"00000000",
  54015=>"00000000",
  54016=>"00000000",
  54017=>"00000000",
  54018=>"00000000",
  54019=>"00000000",
  54020=>"00000000",
  54021=>"11111111",
  54022=>"00000000",
  54023=>"00000000",
  54024=>"00000000",
  54025=>"00000000",
  54026=>"00000000",
  54027=>"00000000",
  54028=>"00000000",
  54029=>"00000000",
  54030=>"00000000",
  54031=>"00000000",
  54032=>"00000000",
  54033=>"00000001",
  54034=>"00000000",
  54035=>"00000000",
  54036=>"00000000",
  54037=>"00000000",
  54038=>"00000000",
  54039=>"00000000",
  54040=>"00000000",
  54041=>"00000000",
  54042=>"00000000",
  54043=>"00000001",
  54044=>"11111111",
  54045=>"00000000",
  54046=>"00000000",
  54047=>"00000000",
  54048=>"00000000",
  54049=>"00000000",
  54050=>"11111111",
  54051=>"00000000",
  54052=>"00000000",
  54053=>"00000000",
  54054=>"00000000",
  54055=>"00000000",
  54056=>"00000000",
  54057=>"00000000",
  54058=>"00000000",
  54059=>"00000000",
  54060=>"00000001",
  54061=>"00000000",
  54062=>"00000000",
  54063=>"00000000",
  54064=>"00000000",
  54065=>"00000000",
  54066=>"00000000",
  54067=>"00000001",
  54068=>"00000000",
  54069=>"00000000",
  54070=>"00000000",
  54071=>"00000000",
  54072=>"00000000",
  54073=>"00000001",
  54074=>"00000000",
  54075=>"00000000",
  54076=>"00000000",
  54077=>"00000000",
  54078=>"00000000",
  54079=>"00000000",
  54080=>"00000000",
  54081=>"00000000",
  54082=>"00000000",
  54083=>"00000000",
  54084=>"00000000",
  54085=>"00000000",
  54086=>"11111111",
  54087=>"00000000",
  54088=>"00000000",
  54089=>"11111111",
  54090=>"00000000",
  54091=>"00000000",
  54092=>"00000000",
  54093=>"00000001",
  54094=>"00000000",
  54095=>"00000000",
  54096=>"00000000",
  54097=>"00000000",
  54098=>"00000000",
  54099=>"00000001",
  54100=>"00000000",
  54101=>"00000000",
  54102=>"00000000",
  54103=>"00000000",
  54104=>"00000000",
  54105=>"00000000",
  54106=>"00000000",
  54107=>"00000000",
  54108=>"00000000",
  54109=>"00000000",
  54110=>"00000000",
  54111=>"00000000",
  54112=>"00000000",
  54113=>"00000000",
  54114=>"00000000",
  54115=>"00000001",
  54116=>"00000001",
  54117=>"00000000",
  54118=>"00000000",
  54119=>"11111111",
  54120=>"00000000",
  54121=>"00000000",
  54122=>"00000000",
  54123=>"00000000",
  54124=>"00000000",
  54125=>"00000000",
  54126=>"00000000",
  54127=>"00000000",
  54128=>"00000001",
  54129=>"00000000",
  54130=>"11111111",
  54131=>"00000000",
  54132=>"00000000",
  54133=>"00000000",
  54134=>"00000000",
  54135=>"00000000",
  54136=>"00000000",
  54137=>"11111111",
  54138=>"00000000",
  54139=>"00000000",
  54140=>"00000000",
  54141=>"00000000",
  54142=>"00000000",
  54143=>"00000000",
  54144=>"00000000",
  54145=>"00000000",
  54146=>"00000000",
  54147=>"00000000",
  54148=>"00000000",
  54149=>"00000000",
  54150=>"00000000",
  54151=>"00000000",
  54152=>"00000000",
  54153=>"00000000",
  54154=>"11111111",
  54155=>"11111111",
  54156=>"00000000",
  54157=>"00000001",
  54158=>"00000000",
  54159=>"00000000",
  54160=>"00000000",
  54161=>"00000000",
  54162=>"00000000",
  54163=>"11111111",
  54164=>"00000000",
  54165=>"00000000",
  54166=>"00000000",
  54167=>"00000000",
  54168=>"00000000",
  54169=>"00000000",
  54170=>"11111111",
  54171=>"00000000",
  54172=>"00000000",
  54173=>"00000000",
  54174=>"00000000",
  54175=>"00000000",
  54176=>"00000000",
  54177=>"00000000",
  54178=>"00000001",
  54179=>"00000000",
  54180=>"00000000",
  54181=>"00000000",
  54182=>"00000000",
  54183=>"00000000",
  54184=>"00000000",
  54185=>"00000000",
  54186=>"00000000",
  54187=>"00000000",
  54188=>"00000000",
  54189=>"00000000",
  54190=>"00000000",
  54191=>"00000000",
  54192=>"00000000",
  54193=>"00000000",
  54194=>"00000000",
  54195=>"11111111",
  54196=>"00000000",
  54197=>"00000000",
  54198=>"00000000",
  54199=>"00000000",
  54200=>"00000000",
  54201=>"00000001",
  54202=>"00000000",
  54203=>"00000000",
  54204=>"00000000",
  54205=>"00000000",
  54206=>"00000000",
  54207=>"00000001",
  54208=>"00000000",
  54209=>"00000000",
  54210=>"00000000",
  54211=>"00000000",
  54212=>"00000000",
  54213=>"00000000",
  54214=>"00000000",
  54215=>"00000001",
  54216=>"00000000",
  54217=>"00000000",
  54218=>"00000000",
  54219=>"00000000",
  54220=>"11111111",
  54221=>"00000000",
  54222=>"00000000",
  54223=>"00000000",
  54224=>"00000000",
  54225=>"00000000",
  54226=>"00000000",
  54227=>"00000000",
  54228=>"11111111",
  54229=>"00000000",
  54230=>"00000000",
  54231=>"00000000",
  54232=>"00000001",
  54233=>"00000000",
  54234=>"00000000",
  54235=>"00000000",
  54236=>"00000000",
  54237=>"00000000",
  54238=>"00000000",
  54239=>"00000000",
  54240=>"11111111",
  54241=>"00000000",
  54242=>"00000000",
  54243=>"00000000",
  54244=>"00000000",
  54245=>"00000000",
  54246=>"00000000",
  54247=>"00000000",
  54248=>"00000000",
  54249=>"00000000",
  54250=>"11111111",
  54251=>"00000000",
  54252=>"00000000",
  54253=>"00000000",
  54254=>"00000000",
  54255=>"00000000",
  54256=>"00000000",
  54257=>"00000001",
  54258=>"00000000",
  54259=>"00000001",
  54260=>"00000000",
  54261=>"00000000",
  54262=>"00000000",
  54263=>"00000000",
  54264=>"00000000",
  54265=>"11111111",
  54266=>"00000000",
  54267=>"00000000",
  54268=>"00000001",
  54269=>"00000000",
  54270=>"00000001",
  54271=>"00000000",
  54272=>"00000000",
  54273=>"00000000",
  54274=>"00000000",
  54275=>"00000000",
  54276=>"00000000",
  54277=>"00000000",
  54278=>"00000000",
  54279=>"00000000",
  54280=>"00000000",
  54281=>"00000000",
  54282=>"00000000",
  54283=>"00000000",
  54284=>"00000000",
  54285=>"00000000",
  54286=>"00000000",
  54287=>"00000000",
  54288=>"00000000",
  54289=>"00000000",
  54290=>"00000000",
  54291=>"00000000",
  54292=>"00000000",
  54293=>"00000000",
  54294=>"00000000",
  54295=>"00000000",
  54296=>"00000000",
  54297=>"00000000",
  54298=>"00000000",
  54299=>"00000000",
  54300=>"00000000",
  54301=>"00000000",
  54302=>"00000000",
  54303=>"00000000",
  54304=>"00000000",
  54305=>"00000000",
  54306=>"00000000",
  54307=>"00000000",
  54308=>"00000000",
  54309=>"00000000",
  54310=>"00000000",
  54311=>"00000000",
  54312=>"00000000",
  54313=>"00000000",
  54314=>"00000000",
  54315=>"00000000",
  54316=>"00000000",
  54317=>"00000000",
  54318=>"00000000",
  54319=>"00000000",
  54320=>"00000000",
  54321=>"00000000",
  54322=>"00000000",
  54323=>"00000000",
  54324=>"00000000",
  54325=>"00000000",
  54326=>"00000000",
  54327=>"00000000",
  54328=>"00000000",
  54329=>"00000000",
  54330=>"00000000",
  54331=>"00000000",
  54332=>"00000000",
  54333=>"00000000",
  54334=>"00000000",
  54335=>"00000000",
  54336=>"00000000",
  54337=>"00000000",
  54338=>"00000000",
  54339=>"00000000",
  54340=>"00000000",
  54341=>"00000000",
  54342=>"00000000",
  54343=>"00000000",
  54344=>"00000000",
  54345=>"00000000",
  54346=>"00000000",
  54347=>"00000000",
  54348=>"00000000",
  54349=>"00000000",
  54350=>"00000000",
  54351=>"00000000",
  54352=>"00000000",
  54353=>"00000000",
  54354=>"00000000",
  54355=>"00000000",
  54356=>"00000000",
  54357=>"00000000",
  54358=>"00000000",
  54359=>"00000001",
  54360=>"00000000",
  54361=>"00000000",
  54362=>"00000000",
  54363=>"00000000",
  54364=>"00000000",
  54365=>"00000000",
  54366=>"00000000",
  54367=>"00000000",
  54368=>"00000000",
  54369=>"00000000",
  54370=>"00000000",
  54371=>"00000000",
  54372=>"00000000",
  54373=>"00000000",
  54374=>"00000000",
  54375=>"00000000",
  54376=>"00000000",
  54377=>"00000000",
  54378=>"00000000",
  54379=>"00000000",
  54380=>"00000000",
  54381=>"00000000",
  54382=>"00000000",
  54383=>"00000000",
  54384=>"00000000",
  54385=>"00000000",
  54386=>"00000000",
  54387=>"00000000",
  54388=>"00000000",
  54389=>"00000000",
  54390=>"00000000",
  54391=>"00000000",
  54392=>"00000000",
  54393=>"00000000",
  54394=>"00000000",
  54395=>"00000000",
  54396=>"00000000",
  54397=>"11111111",
  54398=>"00000000",
  54399=>"00000000",
  54400=>"00000000",
  54401=>"00000000",
  54402=>"00000000",
  54403=>"00000000",
  54404=>"00000000",
  54405=>"00000001",
  54406=>"00000000",
  54407=>"00000000",
  54408=>"00000000",
  54409=>"00000000",
  54410=>"00000000",
  54411=>"00000000",
  54412=>"00000000",
  54413=>"00000000",
  54414=>"00000000",
  54415=>"00000000",
  54416=>"00000000",
  54417=>"11111111",
  54418=>"00000000",
  54419=>"00000000",
  54420=>"00000000",
  54421=>"00000000",
  54422=>"00000000",
  54423=>"00000000",
  54424=>"00000000",
  54425=>"00000000",
  54426=>"00000000",
  54427=>"00000000",
  54428=>"11111111",
  54429=>"00000000",
  54430=>"00000000",
  54431=>"00000000",
  54432=>"00000000",
  54433=>"00000000",
  54434=>"00000000",
  54435=>"00000000",
  54436=>"11111111",
  54437=>"00000000",
  54438=>"00000000",
  54439=>"00000000",
  54440=>"00000000",
  54441=>"00000000",
  54442=>"00000000",
  54443=>"00000000",
  54444=>"00000000",
  54445=>"00000000",
  54446=>"00000000",
  54447=>"00000000",
  54448=>"00000000",
  54449=>"00000000",
  54450=>"00000000",
  54451=>"00000000",
  54452=>"00000000",
  54453=>"00000000",
  54454=>"00000000",
  54455=>"00000000",
  54456=>"00000000",
  54457=>"00000000",
  54458=>"00000000",
  54459=>"00000000",
  54460=>"00000000",
  54461=>"11111111",
  54462=>"00000000",
  54463=>"00000000",
  54464=>"00000001",
  54465=>"00000000",
  54466=>"00000000",
  54467=>"00000000",
  54468=>"00000000",
  54469=>"00000000",
  54470=>"00000000",
  54471=>"00000000",
  54472=>"00000000",
  54473=>"00000000",
  54474=>"00000000",
  54475=>"00000000",
  54476=>"00000000",
  54477=>"00000000",
  54478=>"00000000",
  54479=>"00000000",
  54480=>"00000000",
  54481=>"00000000",
  54482=>"00000010",
  54483=>"00000000",
  54484=>"11111111",
  54485=>"00000000",
  54486=>"00000000",
  54487=>"00000000",
  54488=>"00000000",
  54489=>"00000000",
  54490=>"00000001",
  54491=>"00000000",
  54492=>"00000000",
  54493=>"00000000",
  54494=>"00000000",
  54495=>"00000000",
  54496=>"00000000",
  54497=>"00000000",
  54498=>"00000000",
  54499=>"00000000",
  54500=>"00000000",
  54501=>"00000000",
  54502=>"00000000",
  54503=>"00000000",
  54504=>"00000000",
  54505=>"00000000",
  54506=>"00000000",
  54507=>"00000000",
  54508=>"00000000",
  54509=>"00000000",
  54510=>"00000000",
  54511=>"00000001",
  54512=>"00000000",
  54513=>"00000000",
  54514=>"00000000",
  54515=>"00000000",
  54516=>"00000000",
  54517=>"00000000",
  54518=>"00000000",
  54519=>"00000000",
  54520=>"00000000",
  54521=>"00000000",
  54522=>"00000000",
  54523=>"00000001",
  54524=>"00000000",
  54525=>"00000000",
  54526=>"00000000",
  54527=>"11111111",
  54528=>"00000000",
  54529=>"00000000",
  54530=>"00000000",
  54531=>"00000000",
  54532=>"00000001",
  54533=>"00000000",
  54534=>"00000000",
  54535=>"00000000",
  54536=>"00000000",
  54537=>"00000000",
  54538=>"00000000",
  54539=>"00000000",
  54540=>"00000000",
  54541=>"00000000",
  54542=>"00000000",
  54543=>"00000000",
  54544=>"00000000",
  54545=>"11111111",
  54546=>"00000001",
  54547=>"00000000",
  54548=>"00000000",
  54549=>"00000000",
  54550=>"00000000",
  54551=>"00000000",
  54552=>"00000000",
  54553=>"00000000",
  54554=>"00000000",
  54555=>"00000000",
  54556=>"00000000",
  54557=>"00000000",
  54558=>"00000000",
  54559=>"00000000",
  54560=>"00000000",
  54561=>"00000000",
  54562=>"00000001",
  54563=>"00000000",
  54564=>"00000000",
  54565=>"00000000",
  54566=>"00000000",
  54567=>"00000000",
  54568=>"00000000",
  54569=>"00000000",
  54570=>"00000000",
  54571=>"00000000",
  54572=>"00000000",
  54573=>"00000001",
  54574=>"00000000",
  54575=>"00000000",
  54576=>"00000000",
  54577=>"00000001",
  54578=>"11111111",
  54579=>"00000000",
  54580=>"00000000",
  54581=>"00000000",
  54582=>"00000000",
  54583=>"00000001",
  54584=>"00000000",
  54585=>"00000000",
  54586=>"00000000",
  54587=>"00000000",
  54588=>"00000000",
  54589=>"00000000",
  54590=>"00000000",
  54591=>"00000000",
  54592=>"00000000",
  54593=>"00000000",
  54594=>"00000001",
  54595=>"00000000",
  54596=>"00000000",
  54597=>"00000000",
  54598=>"00000000",
  54599=>"00000001",
  54600=>"00000000",
  54601=>"00000000",
  54602=>"00000000",
  54603=>"00000000",
  54604=>"00000000",
  54605=>"00000000",
  54606=>"00000000",
  54607=>"00000000",
  54608=>"00000000",
  54609=>"00000000",
  54610=>"00000000",
  54611=>"00000000",
  54612=>"00000001",
  54613=>"00000000",
  54614=>"00000000",
  54615=>"00000000",
  54616=>"00000000",
  54617=>"00000000",
  54618=>"00000000",
  54619=>"00000000",
  54620=>"00000000",
  54621=>"00000000",
  54622=>"00000000",
  54623=>"00000000",
  54624=>"00000000",
  54625=>"00000000",
  54626=>"00000000",
  54627=>"00000000",
  54628=>"00000000",
  54629=>"00000000",
  54630=>"00000000",
  54631=>"00000000",
  54632=>"00000000",
  54633=>"00000000",
  54634=>"00000000",
  54635=>"00000000",
  54636=>"00000000",
  54637=>"00000000",
  54638=>"00000000",
  54639=>"00000001",
  54640=>"00000000",
  54641=>"00000000",
  54642=>"00000000",
  54643=>"00000000",
  54644=>"00000000",
  54645=>"00000000",
  54646=>"00000000",
  54647=>"00000000",
  54648=>"00000000",
  54649=>"00000000",
  54650=>"00000000",
  54651=>"00000000",
  54652=>"00000000",
  54653=>"00000000",
  54654=>"00000000",
  54655=>"00000000",
  54656=>"00000000",
  54657=>"00000000",
  54658=>"00000000",
  54659=>"00000000",
  54660=>"00000000",
  54661=>"00000000",
  54662=>"00000000",
  54663=>"00000000",
  54664=>"00000000",
  54665=>"00000000",
  54666=>"00000000",
  54667=>"11111111",
  54668=>"00000000",
  54669=>"00000000",
  54670=>"00000000",
  54671=>"00000000",
  54672=>"00000000",
  54673=>"00000000",
  54674=>"00000000",
  54675=>"00000000",
  54676=>"00000000",
  54677=>"00000000",
  54678=>"00000000",
  54679=>"00000000",
  54680=>"00000000",
  54681=>"00000000",
  54682=>"00000000",
  54683=>"00000000",
  54684=>"00000000",
  54685=>"00000000",
  54686=>"00000000",
  54687=>"00000000",
  54688=>"00000000",
  54689=>"00000000",
  54690=>"00000000",
  54691=>"00000000",
  54692=>"00000000",
  54693=>"00000000",
  54694=>"00000000",
  54695=>"00000000",
  54696=>"00000000",
  54697=>"00000000",
  54698=>"00000000",
  54699=>"00000000",
  54700=>"00000000",
  54701=>"00000000",
  54702=>"00000000",
  54703=>"00000000",
  54704=>"00000000",
  54705=>"00000000",
  54706=>"00000000",
  54707=>"11111111",
  54708=>"00000000",
  54709=>"00000000",
  54710=>"00000000",
  54711=>"00000000",
  54712=>"00000000",
  54713=>"00000000",
  54714=>"00000000",
  54715=>"00000000",
  54716=>"00000000",
  54717=>"00000000",
  54718=>"00000000",
  54719=>"00000000",
  54720=>"00000000",
  54721=>"00000000",
  54722=>"00000000",
  54723=>"00000000",
  54724=>"00000000",
  54725=>"00000000",
  54726=>"00000000",
  54727=>"00000000",
  54728=>"00000000",
  54729=>"00000000",
  54730=>"00000000",
  54731=>"00000000",
  54732=>"00000000",
  54733=>"00000000",
  54734=>"00000000",
  54735=>"00000000",
  54736=>"00000000",
  54737=>"00000000",
  54738=>"00000000",
  54739=>"00000000",
  54740=>"00000000",
  54741=>"00000000",
  54742=>"00000000",
  54743=>"00000000",
  54744=>"00000000",
  54745=>"00000000",
  54746=>"00000000",
  54747=>"00000000",
  54748=>"00000000",
  54749=>"00000000",
  54750=>"00000000",
  54751=>"00000000",
  54752=>"00000000",
  54753=>"00000000",
  54754=>"00000000",
  54755=>"11111111",
  54756=>"00000000",
  54757=>"00000000",
  54758=>"00000000",
  54759=>"00000000",
  54760=>"00000000",
  54761=>"00000000",
  54762=>"00000000",
  54763=>"00000000",
  54764=>"00000000",
  54765=>"00000000",
  54766=>"00000000",
  54767=>"00000000",
  54768=>"00000001",
  54769=>"00000000",
  54770=>"00000000",
  54771=>"00000000",
  54772=>"00000000",
  54773=>"00000000",
  54774=>"00000000",
  54775=>"00000000",
  54776=>"00000000",
  54777=>"00000000",
  54778=>"00000000",
  54779=>"00000000",
  54780=>"00000000",
  54781=>"00000000",
  54782=>"00000000",
  54783=>"00000000",
  54784=>"00000000",
  54785=>"00000000",
  54786=>"00000000",
  54787=>"00000000",
  54788=>"00000000",
  54789=>"00000000",
  54790=>"00000000",
  54791=>"00000000",
  54792=>"00000000",
  54793=>"00000000",
  54794=>"00000000",
  54795=>"00000000",
  54796=>"00000000",
  54797=>"00000000",
  54798=>"00000000",
  54799=>"00000000",
  54800=>"00000000",
  54801=>"00000000",
  54802=>"00000000",
  54803=>"00000000",
  54804=>"00000000",
  54805=>"00000000",
  54806=>"00000000",
  54807=>"00000000",
  54808=>"00000000",
  54809=>"00000000",
  54810=>"00000000",
  54811=>"00000000",
  54812=>"11111111",
  54813=>"00000000",
  54814=>"00000000",
  54815=>"00000000",
  54816=>"00000000",
  54817=>"00000000",
  54818=>"00000000",
  54819=>"00000000",
  54820=>"00000000",
  54821=>"00000000",
  54822=>"00000000",
  54823=>"11111111",
  54824=>"00000000",
  54825=>"00000000",
  54826=>"00000000",
  54827=>"00000000",
  54828=>"00000000",
  54829=>"00000000",
  54830=>"00000000",
  54831=>"00000000",
  54832=>"00000000",
  54833=>"00000000",
  54834=>"00000000",
  54835=>"00000000",
  54836=>"00000000",
  54837=>"00000000",
  54838=>"00000000",
  54839=>"00000000",
  54840=>"00000001",
  54841=>"00000000",
  54842=>"00000000",
  54843=>"00000000",
  54844=>"00000000",
  54845=>"00000000",
  54846=>"11111111",
  54847=>"00000000",
  54848=>"00000000",
  54849=>"00000000",
  54850=>"00000000",
  54851=>"00000000",
  54852=>"00000000",
  54853=>"00000000",
  54854=>"00000000",
  54855=>"00000000",
  54856=>"00000001",
  54857=>"00000000",
  54858=>"00000000",
  54859=>"00000000",
  54860=>"00000000",
  54861=>"00000000",
  54862=>"00000000",
  54863=>"00000001",
  54864=>"00000000",
  54865=>"00000000",
  54866=>"00000000",
  54867=>"00000000",
  54868=>"00000000",
  54869=>"00000000",
  54870=>"00000001",
  54871=>"00000000",
  54872=>"00000000",
  54873=>"00000000",
  54874=>"11111111",
  54875=>"00000000",
  54876=>"00000000",
  54877=>"00000000",
  54878=>"00000000",
  54879=>"00000000",
  54880=>"00000000",
  54881=>"00000000",
  54882=>"00000000",
  54883=>"00000000",
  54884=>"00000000",
  54885=>"00000000",
  54886=>"00000001",
  54887=>"00000000",
  54888=>"00000000",
  54889=>"00000000",
  54890=>"00000000",
  54891=>"00000000",
  54892=>"00000000",
  54893=>"00000000",
  54894=>"00000000",
  54895=>"00000000",
  54896=>"00000000",
  54897=>"00000000",
  54898=>"00000000",
  54899=>"00000000",
  54900=>"00000000",
  54901=>"00000000",
  54902=>"00000000",
  54903=>"00000000",
  54904=>"00000000",
  54905=>"00000000",
  54906=>"00000000",
  54907=>"00000000",
  54908=>"00000000",
  54909=>"00000000",
  54910=>"00000000",
  54911=>"00000000",
  54912=>"00000000",
  54913=>"00000000",
  54914=>"00000000",
  54915=>"00000000",
  54916=>"00000000",
  54917=>"00000000",
  54918=>"00000000",
  54919=>"00000000",
  54920=>"00000000",
  54921=>"00000000",
  54922=>"00000000",
  54923=>"00000000",
  54924=>"00000000",
  54925=>"00000000",
  54926=>"00000001",
  54927=>"00000000",
  54928=>"00000000",
  54929=>"00000000",
  54930=>"00000000",
  54931=>"00000000",
  54932=>"00000000",
  54933=>"00000000",
  54934=>"00000000",
  54935=>"00000000",
  54936=>"00000000",
  54937=>"00000000",
  54938=>"00000000",
  54939=>"00000000",
  54940=>"00000000",
  54941=>"00000000",
  54942=>"00000000",
  54943=>"00000000",
  54944=>"00000001",
  54945=>"00000000",
  54946=>"00000000",
  54947=>"00000000",
  54948=>"00000000",
  54949=>"00000000",
  54950=>"00000000",
  54951=>"00000000",
  54952=>"00000000",
  54953=>"00000000",
  54954=>"00000000",
  54955=>"00000000",
  54956=>"00000000",
  54957=>"00000000",
  54958=>"00000000",
  54959=>"00000000",
  54960=>"00000000",
  54961=>"00000000",
  54962=>"00000000",
  54963=>"00000000",
  54964=>"00000001",
  54965=>"00000000",
  54966=>"00000000",
  54967=>"00000000",
  54968=>"00000000",
  54969=>"00000000",
  54970=>"00000001",
  54971=>"00000000",
  54972=>"00000000",
  54973=>"00000000",
  54974=>"00000000",
  54975=>"00000001",
  54976=>"00000000",
  54977=>"00000000",
  54978=>"00000000",
  54979=>"00000000",
  54980=>"00000000",
  54981=>"00000000",
  54982=>"00000000",
  54983=>"00000000",
  54984=>"00000000",
  54985=>"00000000",
  54986=>"00000000",
  54987=>"00000000",
  54988=>"00000000",
  54989=>"00000000",
  54990=>"00000000",
  54991=>"00000000",
  54992=>"00000000",
  54993=>"00000000",
  54994=>"00000000",
  54995=>"00000000",
  54996=>"00000000",
  54997=>"00000000",
  54998=>"00000000",
  54999=>"00000000",
  55000=>"00000000",
  55001=>"00000001",
  55002=>"11111111",
  55003=>"00000000",
  55004=>"00000000",
  55005=>"00000000",
  55006=>"00000000",
  55007=>"00000000",
  55008=>"00000000",
  55009=>"00000000",
  55010=>"00000000",
  55011=>"00000000",
  55012=>"00000000",
  55013=>"00000000",
  55014=>"00000000",
  55015=>"00000000",
  55016=>"00000000",
  55017=>"00000000",
  55018=>"00000000",
  55019=>"00000000",
  55020=>"00000000",
  55021=>"00000000",
  55022=>"00000000",
  55023=>"00000000",
  55024=>"00000000",
  55025=>"00000000",
  55026=>"00000000",
  55027=>"00000001",
  55028=>"00000000",
  55029=>"00000000",
  55030=>"00000000",
  55031=>"00000000",
  55032=>"00000000",
  55033=>"00000000",
  55034=>"00000000",
  55035=>"00000000",
  55036=>"00000000",
  55037=>"00000000",
  55038=>"00000000",
  55039=>"00000000",
  55040=>"00000000",
  55041=>"00000000",
  55042=>"00000000",
  55043=>"00000000",
  55044=>"00000000",
  55045=>"00000000",
  55046=>"00000000",
  55047=>"00000000",
  55048=>"00000000",
  55049=>"00000000",
  55050=>"00000000",
  55051=>"00000000",
  55052=>"00000000",
  55053=>"00000000",
  55054=>"00000000",
  55055=>"00000000",
  55056=>"00000000",
  55057=>"00000000",
  55058=>"00000000",
  55059=>"00000000",
  55060=>"00000000",
  55061=>"00000000",
  55062=>"00000000",
  55063=>"00000000",
  55064=>"00000000",
  55065=>"00000000",
  55066=>"00000000",
  55067=>"00000000",
  55068=>"00000000",
  55069=>"00000000",
  55070=>"00000000",
  55071=>"00000000",
  55072=>"00000000",
  55073=>"00000000",
  55074=>"00000001",
  55075=>"00000000",
  55076=>"00000000",
  55077=>"00000000",
  55078=>"00000000",
  55079=>"00000000",
  55080=>"00000000",
  55081=>"00000000",
  55082=>"00000000",
  55083=>"00000000",
  55084=>"00000000",
  55085=>"00000000",
  55086=>"00000000",
  55087=>"00000000",
  55088=>"00000000",
  55089=>"00000000",
  55090=>"00000000",
  55091=>"00000000",
  55092=>"00000000",
  55093=>"00000000",
  55094=>"00000000",
  55095=>"00000000",
  55096=>"00000000",
  55097=>"00000000",
  55098=>"00000000",
  55099=>"00000000",
  55100=>"00000000",
  55101=>"00000000",
  55102=>"00000000",
  55103=>"00000000",
  55104=>"00000000",
  55105=>"00000000",
  55106=>"00000000",
  55107=>"00000000",
  55108=>"00000000",
  55109=>"00000000",
  55110=>"00000000",
  55111=>"00000000",
  55112=>"00000000",
  55113=>"00000000",
  55114=>"00000000",
  55115=>"00000000",
  55116=>"00000000",
  55117=>"00000001",
  55118=>"00000000",
  55119=>"00000000",
  55120=>"00000000",
  55121=>"00000000",
  55122=>"00000000",
  55123=>"00000000",
  55124=>"00000000",
  55125=>"00000000",
  55126=>"00000000",
  55127=>"00000000",
  55128=>"00000000",
  55129=>"00000000",
  55130=>"00000000",
  55131=>"00000000",
  55132=>"00000000",
  55133=>"00000000",
  55134=>"00000000",
  55135=>"00000000",
  55136=>"00000000",
  55137=>"00000000",
  55138=>"00000000",
  55139=>"00000000",
  55140=>"00000000",
  55141=>"00000000",
  55142=>"00000000",
  55143=>"00000000",
  55144=>"00000000",
  55145=>"00000000",
  55146=>"00000000",
  55147=>"00000000",
  55148=>"00000000",
  55149=>"00000000",
  55150=>"00000000",
  55151=>"00000000",
  55152=>"00000000",
  55153=>"00000000",
  55154=>"00000001",
  55155=>"00000000",
  55156=>"00000000",
  55157=>"00000000",
  55158=>"00000000",
  55159=>"00000000",
  55160=>"00000000",
  55161=>"00000000",
  55162=>"00000000",
  55163=>"00000000",
  55164=>"00000000",
  55165=>"00000000",
  55166=>"00000000",
  55167=>"00000000",
  55168=>"00000001",
  55169=>"00000000",
  55170=>"00000001",
  55171=>"00000000",
  55172=>"00000000",
  55173=>"00000001",
  55174=>"00000000",
  55175=>"00000000",
  55176=>"00000000",
  55177=>"00000000",
  55178=>"00000000",
  55179=>"11111111",
  55180=>"00000000",
  55181=>"00000000",
  55182=>"00000000",
  55183=>"00000000",
  55184=>"00000000",
  55185=>"00000000",
  55186=>"00000000",
  55187=>"00000000",
  55188=>"00000000",
  55189=>"00000000",
  55190=>"00000000",
  55191=>"00000000",
  55192=>"00000000",
  55193=>"00000000",
  55194=>"00000000",
  55195=>"00000000",
  55196=>"00000000",
  55197=>"00000000",
  55198=>"00000000",
  55199=>"00000000",
  55200=>"00000000",
  55201=>"00000000",
  55202=>"00000000",
  55203=>"00000000",
  55204=>"00000000",
  55205=>"00000000",
  55206=>"00000000",
  55207=>"00000000",
  55208=>"00000001",
  55209=>"00000001",
  55210=>"00000000",
  55211=>"00000000",
  55212=>"00000000",
  55213=>"00000000",
  55214=>"00000000",
  55215=>"00000000",
  55216=>"00000000",
  55217=>"00000000",
  55218=>"00000000",
  55219=>"00000000",
  55220=>"00000000",
  55221=>"00000000",
  55222=>"00000000",
  55223=>"00000000",
  55224=>"00000000",
  55225=>"00000000",
  55226=>"00000000",
  55227=>"00000000",
  55228=>"00000000",
  55229=>"00000000",
  55230=>"00000000",
  55231=>"00000000",
  55232=>"00000000",
  55233=>"00000000",
  55234=>"00000000",
  55235=>"00000000",
  55236=>"00000000",
  55237=>"00000000",
  55238=>"00000000",
  55239=>"00000000",
  55240=>"00000000",
  55241=>"00000000",
  55242=>"00000000",
  55243=>"00000000",
  55244=>"00000000",
  55245=>"00000000",
  55246=>"00000000",
  55247=>"00000000",
  55248=>"11111111",
  55249=>"00000000",
  55250=>"00000000",
  55251=>"00000000",
  55252=>"00000000",
  55253=>"00000000",
  55254=>"00000000",
  55255=>"00000000",
  55256=>"00000000",
  55257=>"00000000",
  55258=>"00000000",
  55259=>"00000000",
  55260=>"00000000",
  55261=>"00000000",
  55262=>"00000000",
  55263=>"00000000",
  55264=>"00000000",
  55265=>"00000000",
  55266=>"00000000",
  55267=>"00000000",
  55268=>"00000000",
  55269=>"00000000",
  55270=>"00000000",
  55271=>"00000000",
  55272=>"00000000",
  55273=>"00000000",
  55274=>"00000000",
  55275=>"00000000",
  55276=>"00000000",
  55277=>"00000000",
  55278=>"00000000",
  55279=>"00000000",
  55280=>"00000000",
  55281=>"00000001",
  55282=>"00000000",
  55283=>"00000001",
  55284=>"00000000",
  55285=>"00000000",
  55286=>"00000000",
  55287=>"00000000",
  55288=>"00000000",
  55289=>"00000000",
  55290=>"00000000",
  55291=>"00000000",
  55292=>"00000000",
  55293=>"00000000",
  55294=>"00000000",
  55295=>"00000000",
  55296=>"00000001",
  55297=>"11111110",
  55298=>"11111010",
  55299=>"11111100",
  55300=>"00000011",
  55301=>"00000100",
  55302=>"11111010",
  55303=>"11111101",
  55304=>"00000000",
  55305=>"00000001",
  55306=>"11111110",
  55307=>"00000000",
  55308=>"11111100",
  55309=>"11111111",
  55310=>"00000101",
  55311=>"00000010",
  55312=>"11111110",
  55313=>"00000011",
  55314=>"11111110",
  55315=>"11111101",
  55316=>"00000001",
  55317=>"11111110",
  55318=>"00000000",
  55319=>"00000001",
  55320=>"11111111",
  55321=>"11111111",
  55322=>"00000010",
  55323=>"00000001",
  55324=>"11111011",
  55325=>"11111011",
  55326=>"11111101",
  55327=>"00000000",
  55328=>"00000001",
  55329=>"11111111",
  55330=>"00000000",
  55331=>"11111101",
  55332=>"11111101",
  55333=>"11111101",
  55334=>"11111111",
  55335=>"00000001",
  55336=>"00000100",
  55337=>"00000010",
  55338=>"00000110",
  55339=>"00000010",
  55340=>"00000101",
  55341=>"11110111",
  55342=>"11111101",
  55343=>"00000011",
  55344=>"11111001",
  55345=>"00000000",
  55346=>"11111111",
  55347=>"00000010",
  55348=>"11110101",
  55349=>"00000001",
  55350=>"11111100",
  55351=>"11111111",
  55352=>"11111111",
  55353=>"00000001",
  55354=>"00000000",
  55355=>"00000000",
  55356=>"11111111",
  55357=>"11111100",
  55358=>"11111110",
  55359=>"11111100",
  55360=>"00000110",
  55361=>"00000011",
  55362=>"00000001",
  55363=>"11111001",
  55364=>"11111011",
  55365=>"00000011",
  55366=>"00000001",
  55367=>"00000001",
  55368=>"00000010",
  55369=>"00000001",
  55370=>"00000000",
  55371=>"00000000",
  55372=>"00000010",
  55373=>"00000011",
  55374=>"11111101",
  55375=>"11111001",
  55376=>"00000001",
  55377=>"00000001",
  55378=>"00000010",
  55379=>"00000010",
  55380=>"00000010",
  55381=>"00000010",
  55382=>"00000001",
  55383=>"11111000",
  55384=>"11111100",
  55385=>"11111111",
  55386=>"11111110",
  55387=>"00000010",
  55388=>"00000010",
  55389=>"11111111",
  55390=>"11111100",
  55391=>"00000001",
  55392=>"11111111",
  55393=>"00000001",
  55394=>"00000010",
  55395=>"11111110",
  55396=>"00000000",
  55397=>"00000010",
  55398=>"11111110",
  55399=>"00000001",
  55400=>"11111111",
  55401=>"00000001",
  55402=>"11111111",
  55403=>"11111100",
  55404=>"00000000",
  55405=>"11111111",
  55406=>"11111100",
  55407=>"00000001",
  55408=>"00000000",
  55409=>"11111101",
  55410=>"00000001",
  55411=>"00000000",
  55412=>"11111010",
  55413=>"11111110",
  55414=>"00000001",
  55415=>"00000000",
  55416=>"00000100",
  55417=>"00000010",
  55418=>"11111111",
  55419=>"11111100",
  55420=>"11111100",
  55421=>"11111000",
  55422=>"11111100",
  55423=>"00000000",
  55424=>"00000011",
  55425=>"11111101",
  55426=>"00000011",
  55427=>"00000010",
  55428=>"00000001",
  55429=>"00000101",
  55430=>"11110110",
  55431=>"00000000",
  55432=>"00000001",
  55433=>"11111101",
  55434=>"00000011",
  55435=>"00000001",
  55436=>"00000000",
  55437=>"11111000",
  55438=>"00000010",
  55439=>"11111110",
  55440=>"11111011",
  55441=>"00000000",
  55442=>"11111010",
  55443=>"11111110",
  55444=>"00000000",
  55445=>"00000011",
  55446=>"00000001",
  55447=>"00000000",
  55448=>"00000011",
  55449=>"00000000",
  55450=>"00000001",
  55451=>"00000010",
  55452=>"11111010",
  55453=>"00000001",
  55454=>"11111001",
  55455=>"11111111",
  55456=>"00000000",
  55457=>"11111100",
  55458=>"00000011",
  55459=>"00000000",
  55460=>"11111010",
  55461=>"00000000",
  55462=>"00000000",
  55463=>"00000010",
  55464=>"00000011",
  55465=>"11111110",
  55466=>"00000000",
  55467=>"11111111",
  55468=>"11111101",
  55469=>"11111101",
  55470=>"11111101",
  55471=>"00000000",
  55472=>"00000011",
  55473=>"00000001",
  55474=>"00000010",
  55475=>"00000001",
  55476=>"00000001",
  55477=>"00000000",
  55478=>"00000001",
  55479=>"11111111",
  55480=>"00000000",
  55481=>"11111101",
  55482=>"11111110",
  55483=>"00000001",
  55484=>"11111110",
  55485=>"11111011",
  55486=>"11111100",
  55487=>"00000001",
  55488=>"00000010",
  55489=>"11111001",
  55490=>"11111110",
  55491=>"00000001",
  55492=>"11111110",
  55493=>"00000000",
  55494=>"00000000",
  55495=>"11111110",
  55496=>"11111110",
  55497=>"00000100",
  55498=>"11111011",
  55499=>"00000000",
  55500=>"00000011",
  55501=>"11111010",
  55502=>"11111100",
  55503=>"11111111",
  55504=>"00000011",
  55505=>"11111111",
  55506=>"11111101",
  55507=>"11111101",
  55508=>"11111001",
  55509=>"00000001",
  55510=>"00000000",
  55511=>"11111111",
  55512=>"00000010",
  55513=>"00000000",
  55514=>"00000000",
  55515=>"11111110",
  55516=>"11111101",
  55517=>"11111111",
  55518=>"11111111",
  55519=>"00000101",
  55520=>"11111100",
  55521=>"11111111",
  55522=>"00000001",
  55523=>"11111011",
  55524=>"00000001",
  55525=>"11111111",
  55526=>"00000001",
  55527=>"11111110",
  55528=>"11110111",
  55529=>"00000010",
  55530=>"11111110",
  55531=>"11111010",
  55532=>"11110111",
  55533=>"00000010",
  55534=>"00000000",
  55535=>"11111001",
  55536=>"00000001",
  55537=>"00000000",
  55538=>"00000001",
  55539=>"00000001",
  55540=>"11111110",
  55541=>"00000001",
  55542=>"11111101",
  55543=>"00000001",
  55544=>"00000000",
  55545=>"11111111",
  55546=>"00000100",
  55547=>"11111100",
  55548=>"00000011",
  55549=>"11111001",
  55550=>"00000000",
  55551=>"11111101",
  55552=>"11111110",
  55553=>"00000001",
  55554=>"00000000",
  55555=>"00000010",
  55556=>"11111111",
  55557=>"00000011",
  55558=>"11111110",
  55559=>"11111110",
  55560=>"11111110",
  55561=>"00000010",
  55562=>"11111110",
  55563=>"00000011",
  55564=>"11111100",
  55565=>"11111111",
  55566=>"11111000",
  55567=>"11111111",
  55568=>"00000000",
  55569=>"11111110",
  55570=>"11111001",
  55571=>"00000000",
  55572=>"11111111",
  55573=>"11111000",
  55574=>"11111100",
  55575=>"00000000",
  55576=>"00000110",
  55577=>"11111100",
  55578=>"11111000",
  55579=>"11111101",
  55580=>"00000000",
  55581=>"11111110",
  55582=>"00000000",
  55583=>"00000001",
  55584=>"11111011",
  55585=>"00000011",
  55586=>"11111100",
  55587=>"11111100",
  55588=>"00000000",
  55589=>"00000100",
  55590=>"11111110",
  55591=>"11111111",
  55592=>"00000000",
  55593=>"11111110",
  55594=>"11111011",
  55595=>"00000011",
  55596=>"00000000",
  55597=>"11111010",
  55598=>"11111011",
  55599=>"00000001",
  55600=>"00001001",
  55601=>"11111110",
  55602=>"00000111",
  55603=>"00000010",
  55604=>"00000000",
  55605=>"11111110",
  55606=>"11111110",
  55607=>"00000010",
  55608=>"11111101",
  55609=>"00000000",
  55610=>"11111001",
  55611=>"11111111",
  55612=>"11111101",
  55613=>"11111111",
  55614=>"11111111",
  55615=>"11111101",
  55616=>"11111011",
  55617=>"11111111",
  55618=>"00000001",
  55619=>"11111000",
  55620=>"11110111",
  55621=>"11111011",
  55622=>"00000000",
  55623=>"00000010",
  55624=>"11111111",
  55625=>"11111110",
  55626=>"00000000",
  55627=>"11111100",
  55628=>"00000000",
  55629=>"00000000",
  55630=>"00000001",
  55631=>"11111110",
  55632=>"11111101",
  55633=>"11111111",
  55634=>"11111011",
  55635=>"00000011",
  55636=>"00000000",
  55637=>"11111001",
  55638=>"00000000",
  55639=>"11111110",
  55640=>"11111110",
  55641=>"11110101",
  55642=>"00000001",
  55643=>"00000010",
  55644=>"00000000",
  55645=>"11111101",
  55646=>"11111100",
  55647=>"00000000",
  55648=>"00000001",
  55649=>"00000010",
  55650=>"00000001",
  55651=>"00000001",
  55652=>"11111010",
  55653=>"11111010",
  55654=>"00001001",
  55655=>"11111110",
  55656=>"11111110",
  55657=>"11111001",
  55658=>"11110111",
  55659=>"00000000",
  55660=>"00000010",
  55661=>"11111101",
  55662=>"00000000",
  55663=>"11111011",
  55664=>"11111101",
  55665=>"11111100",
  55666=>"00000110",
  55667=>"00000001",
  55668=>"00000000",
  55669=>"00000001",
  55670=>"11111011",
  55671=>"00000001",
  55672=>"00000001",
  55673=>"11111101",
  55674=>"00000010",
  55675=>"11111101",
  55676=>"11111111",
  55677=>"00000000",
  55678=>"11111011",
  55679=>"00000000",
  55680=>"00000001",
  55681=>"00001001",
  55682=>"11111110",
  55683=>"11111100",
  55684=>"11111011",
  55685=>"00000011",
  55686=>"11111100",
  55687=>"11111100",
  55688=>"11111001",
  55689=>"11111111",
  55690=>"11111111",
  55691=>"11111010",
  55692=>"11111010",
  55693=>"11111100",
  55694=>"00000001",
  55695=>"11111110",
  55696=>"11111000",
  55697=>"00000001",
  55698=>"00000010",
  55699=>"00000001",
  55700=>"00000000",
  55701=>"11111010",
  55702=>"11111101",
  55703=>"11111110",
  55704=>"11111101",
  55705=>"00000101",
  55706=>"11111110",
  55707=>"11111101",
  55708=>"11111100",
  55709=>"00000101",
  55710=>"00000010",
  55711=>"00000001",
  55712=>"00000000",
  55713=>"11111101",
  55714=>"00000010",
  55715=>"00000010",
  55716=>"11110011",
  55717=>"11111110",
  55718=>"11111111",
  55719=>"11111110",
  55720=>"00000001",
  55721=>"00000000",
  55722=>"00000001",
  55723=>"00000000",
  55724=>"00000010",
  55725=>"00000001",
  55726=>"00000101",
  55727=>"11111100",
  55728=>"00000000",
  55729=>"11111111",
  55730=>"11111011",
  55731=>"00000011",
  55732=>"11111111",
  55733=>"00000001",
  55734=>"00000000",
  55735=>"00000001",
  55736=>"00001000",
  55737=>"11111111",
  55738=>"11111010",
  55739=>"11111010",
  55740=>"11111010",
  55741=>"00000000",
  55742=>"00000010",
  55743=>"11111010",
  55744=>"00000011",
  55745=>"00000010",
  55746=>"11111110",
  55747=>"00000010",
  55748=>"11111011",
  55749=>"11111111",
  55750=>"00000001",
  55751=>"00000010",
  55752=>"11111110",
  55753=>"11111110",
  55754=>"00000000",
  55755=>"00000001",
  55756=>"11111100",
  55757=>"11111011",
  55758=>"11111000",
  55759=>"11111111",
  55760=>"00000000",
  55761=>"11111011",
  55762=>"11111011",
  55763=>"11111111",
  55764=>"11111011",
  55765=>"00000001",
  55766=>"11111101",
  55767=>"00000011",
  55768=>"11111000",
  55769=>"11111111",
  55770=>"11110110",
  55771=>"11111101",
  55772=>"00000001",
  55773=>"00000001",
  55774=>"00000000",
  55775=>"11111111",
  55776=>"00000110",
  55777=>"00000001",
  55778=>"11111111",
  55779=>"11111000",
  55780=>"11110110",
  55781=>"00000000",
  55782=>"00000000",
  55783=>"11111000",
  55784=>"00000000",
  55785=>"11111101",
  55786=>"00000110",
  55787=>"11111111",
  55788=>"00001100",
  55789=>"00000110",
  55790=>"00000010",
  55791=>"00000001",
  55792=>"11111011",
  55793=>"00000001",
  55794=>"11111001",
  55795=>"11111100",
  55796=>"11111111",
  55797=>"11111110",
  55798=>"00000010",
  55799=>"00000110",
  55800=>"11111111",
  55801=>"00000100",
  55802=>"11111110",
  55803=>"11111100",
  55804=>"00000010",
  55805=>"00000001",
  55806=>"00000001",
  55807=>"00000010",
  55808=>"11111100",
  55809=>"11111101",
  55810=>"00000001",
  55811=>"11111111",
  55812=>"00000001",
  55813=>"11111110",
  55814=>"00000011",
  55815=>"00000110",
  55816=>"11111100",
  55817=>"00000000",
  55818=>"11111010",
  55819=>"11111000",
  55820=>"11111111",
  55821=>"00000011",
  55822=>"00000010",
  55823=>"00000000",
  55824=>"00000000",
  55825=>"00000010",
  55826=>"00000000",
  55827=>"11111111",
  55828=>"00000000",
  55829=>"11111110",
  55830=>"11111100",
  55831=>"11111011",
  55832=>"11111111",
  55833=>"00000000",
  55834=>"11111000",
  55835=>"11111000",
  55836=>"11111010",
  55837=>"00000010",
  55838=>"11111001",
  55839=>"00000000",
  55840=>"00000011",
  55841=>"11111000",
  55842=>"11111011",
  55843=>"00000001",
  55844=>"11111100",
  55845=>"00000001",
  55846=>"11111100",
  55847=>"11111110",
  55848=>"11111110",
  55849=>"11111111",
  55850=>"11111111",
  55851=>"11111111",
  55852=>"11111111",
  55853=>"00000000",
  55854=>"11111101",
  55855=>"00000011",
  55856=>"00000010",
  55857=>"00000010",
  55858=>"11111011",
  55859=>"00001000",
  55860=>"00000001",
  55861=>"00000000",
  55862=>"11111000",
  55863=>"11111110",
  55864=>"00000001",
  55865=>"11110111",
  55866=>"00000000",
  55867=>"00000011",
  55868=>"11111011",
  55869=>"11111111",
  55870=>"11111001",
  55871=>"11111100",
  55872=>"00000010",
  55873=>"00000000",
  55874=>"00000010",
  55875=>"00000001",
  55876=>"00000001",
  55877=>"00000011",
  55878=>"00000100",
  55879=>"00000010",
  55880=>"11111110",
  55881=>"11110111",
  55882=>"11111111",
  55883=>"00000010",
  55884=>"11111111",
  55885=>"11111111",
  55886=>"00000001",
  55887=>"11111111",
  55888=>"11111100",
  55889=>"00000000",
  55890=>"11111100",
  55891=>"11111000",
  55892=>"11111010",
  55893=>"11111100",
  55894=>"11111101",
  55895=>"11111110",
  55896=>"00000000",
  55897=>"11111100",
  55898=>"11111101",
  55899=>"00000000",
  55900=>"00000000",
  55901=>"11111010",
  55902=>"00000001",
  55903=>"00000100",
  55904=>"11111100",
  55905=>"11111101",
  55906=>"11111111",
  55907=>"00000000",
  55908=>"11111101",
  55909=>"00000011",
  55910=>"11111001",
  55911=>"00000010",
  55912=>"00000001",
  55913=>"11111111",
  55914=>"11111001",
  55915=>"11111111",
  55916=>"11111100",
  55917=>"11111111",
  55918=>"00000001",
  55919=>"00000010",
  55920=>"11111111",
  55921=>"00000001",
  55922=>"11111111",
  55923=>"00000000",
  55924=>"11111000",
  55925=>"11111001",
  55926=>"11111101",
  55927=>"00000000",
  55928=>"11111110",
  55929=>"00000001",
  55930=>"11111111",
  55931=>"00000010",
  55932=>"11111001",
  55933=>"11111101",
  55934=>"00000001",
  55935=>"11111010",
  55936=>"11111100",
  55937=>"11111101",
  55938=>"00000010",
  55939=>"00000000",
  55940=>"00000011",
  55941=>"00000010",
  55942=>"11111110",
  55943=>"11111111",
  55944=>"11111111",
  55945=>"00000100",
  55946=>"00000001",
  55947=>"00000000",
  55948=>"11111001",
  55949=>"11111011",
  55950=>"00000111",
  55951=>"00000010",
  55952=>"11111101",
  55953=>"00000001",
  55954=>"11111111",
  55955=>"11111011",
  55956=>"00000001",
  55957=>"11111111",
  55958=>"11111001",
  55959=>"11111111",
  55960=>"11111110",
  55961=>"00000001",
  55962=>"00000001",
  55963=>"11111011",
  55964=>"00000010",
  55965=>"00000001",
  55966=>"00000000",
  55967=>"11111101",
  55968=>"11111001",
  55969=>"11111111",
  55970=>"00000000",
  55971=>"11111111",
  55972=>"11111110",
  55973=>"11111110",
  55974=>"00000000",
  55975=>"00000000",
  55976=>"11111111",
  55977=>"00000001",
  55978=>"11111110",
  55979=>"11111101",
  55980=>"11111001",
  55981=>"11111010",
  55982=>"11110110",
  55983=>"11111110",
  55984=>"00000001",
  55985=>"11111111",
  55986=>"11111111",
  55987=>"11111010",
  55988=>"11111101",
  55989=>"00000010",
  55990=>"11111101",
  55991=>"00000101",
  55992=>"11111111",
  55993=>"11111100",
  55994=>"11111000",
  55995=>"00000000",
  55996=>"11111110",
  55997=>"00000010",
  55998=>"00000101",
  55999=>"11111010",
  56000=>"11111000",
  56001=>"00000010",
  56002=>"00000000",
  56003=>"11111101",
  56004=>"11111011",
  56005=>"11111110",
  56006=>"11111101",
  56007=>"11111111",
  56008=>"00000000",
  56009=>"11111111",
  56010=>"00000010",
  56011=>"11111100",
  56012=>"00000010",
  56013=>"00000011",
  56014=>"11111001",
  56015=>"11111111",
  56016=>"11111001",
  56017=>"11111011",
  56018=>"00000011",
  56019=>"00000001",
  56020=>"00000011",
  56021=>"11111110",
  56022=>"11111010",
  56023=>"00000101",
  56024=>"00000001",
  56025=>"11111111",
  56026=>"11111101",
  56027=>"00000000",
  56028=>"00000000",
  56029=>"11111101",
  56030=>"11111010",
  56031=>"11111111",
  56032=>"00000000",
  56033=>"11111101",
  56034=>"00000010",
  56035=>"00000100",
  56036=>"11111110",
  56037=>"11111110",
  56038=>"11111111",
  56039=>"00000001",
  56040=>"11111111",
  56041=>"11111100",
  56042=>"00000001",
  56043=>"11111101",
  56044=>"11111010",
  56045=>"00000000",
  56046=>"00000000",
  56047=>"11111111",
  56048=>"11111101",
  56049=>"11111101",
  56050=>"11111011",
  56051=>"11111001",
  56052=>"00000000",
  56053=>"00000000",
  56054=>"11111100",
  56055=>"00000000",
  56056=>"00000010",
  56057=>"00000011",
  56058=>"11111001",
  56059=>"11111111",
  56060=>"11111011",
  56061=>"11111111",
  56062=>"11111110",
  56063=>"11111100",
  56064=>"00000001",
  56065=>"11111111",
  56066=>"11111100",
  56067=>"11111111",
  56068=>"00000000",
  56069=>"11111111",
  56070=>"11111010",
  56071=>"11111100",
  56072=>"00000011",
  56073=>"00000001",
  56074=>"11111101",
  56075=>"00000100",
  56076=>"00000001",
  56077=>"00000010",
  56078=>"11111111",
  56079=>"11111010",
  56080=>"11111110",
  56081=>"11111111",
  56082=>"11111110",
  56083=>"00000000",
  56084=>"11111111",
  56085=>"00000000",
  56086=>"11111111",
  56087=>"00000001",
  56088=>"00000011",
  56089=>"11111111",
  56090=>"00000001",
  56091=>"11111111",
  56092=>"00000000",
  56093=>"00000000",
  56094=>"00000000",
  56095=>"11111100",
  56096=>"00000001",
  56097=>"00000001",
  56098=>"11111101",
  56099=>"11110111",
  56100=>"11111011",
  56101=>"00000001",
  56102=>"11111110",
  56103=>"00000010",
  56104=>"00000000",
  56105=>"00000000",
  56106=>"00000001",
  56107=>"11111010",
  56108=>"00000001",
  56109=>"11111110",
  56110=>"11111110",
  56111=>"00000110",
  56112=>"00000000",
  56113=>"00000011",
  56114=>"00000000",
  56115=>"00000011",
  56116=>"11110111",
  56117=>"00000001",
  56118=>"11111011",
  56119=>"00000010",
  56120=>"00000001",
  56121=>"11111000",
  56122=>"11111111",
  56123=>"00000010",
  56124=>"11111110",
  56125=>"11111111",
  56126=>"00000010",
  56127=>"11111101",
  56128=>"00000001",
  56129=>"00000000",
  56130=>"11111110",
  56131=>"00000000",
  56132=>"00000001",
  56133=>"11111100",
  56134=>"00000001",
  56135=>"00000110",
  56136=>"00000000",
  56137=>"11110101",
  56138=>"11111111",
  56139=>"00000001",
  56140=>"11111000",
  56141=>"00000010",
  56142=>"11111111",
  56143=>"00000000",
  56144=>"11111110",
  56145=>"11111001",
  56146=>"11111101",
  56147=>"00000011",
  56148=>"00000000",
  56149=>"11111110",
  56150=>"11111100",
  56151=>"00000001",
  56152=>"11111111",
  56153=>"11111010",
  56154=>"11111111",
  56155=>"00000000",
  56156=>"11111001",
  56157=>"00000000",
  56158=>"11111110",
  56159=>"00000000",
  56160=>"00000001",
  56161=>"00000000",
  56162=>"11111110",
  56163=>"11111011",
  56164=>"11111100",
  56165=>"11111010",
  56166=>"00000010",
  56167=>"11111110",
  56168=>"11111111",
  56169=>"11111111",
  56170=>"11111100",
  56171=>"00000000",
  56172=>"11111101",
  56173=>"00000000",
  56174=>"00000000",
  56175=>"00000000",
  56176=>"00000010",
  56177=>"11111110",
  56178=>"11111011",
  56179=>"00000000",
  56180=>"11111011",
  56181=>"00000001",
  56182=>"11111101",
  56183=>"11111110",
  56184=>"11111110",
  56185=>"11111101",
  56186=>"00000000",
  56187=>"11111110",
  56188=>"11111111",
  56189=>"00000000",
  56190=>"00000001",
  56191=>"11111111",
  56192=>"11111000",
  56193=>"00000100",
  56194=>"11111111",
  56195=>"00000001",
  56196=>"11111011",
  56197=>"00000001",
  56198=>"11111111",
  56199=>"00000001",
  56200=>"00000001",
  56201=>"00000010",
  56202=>"11111001",
  56203=>"00000001",
  56204=>"00000001",
  56205=>"11111100",
  56206=>"00000011",
  56207=>"11111001",
  56208=>"11110100",
  56209=>"00000000",
  56210=>"11111111",
  56211=>"11111000",
  56212=>"11111101",
  56213=>"11111111",
  56214=>"00000001",
  56215=>"00000001",
  56216=>"11111111",
  56217=>"11111110",
  56218=>"11111111",
  56219=>"11111111",
  56220=>"00000010",
  56221=>"11111010",
  56222=>"00000011",
  56223=>"11111000",
  56224=>"00000001",
  56225=>"11110111",
  56226=>"00000000",
  56227=>"11111000",
  56228=>"11111010",
  56229=>"00000001",
  56230=>"00000001",
  56231=>"11111010",
  56232=>"11111100",
  56233=>"00000010",
  56234=>"00000100",
  56235=>"00000000",
  56236=>"11111111",
  56237=>"00000001",
  56238=>"11111001",
  56239=>"11111001",
  56240=>"00000110",
  56241=>"11111111",
  56242=>"11111111",
  56243=>"11111110",
  56244=>"11111000",
  56245=>"00000010",
  56246=>"11111110",
  56247=>"00000110",
  56248=>"11111010",
  56249=>"11111101",
  56250=>"11111101",
  56251=>"11111010",
  56252=>"11111110",
  56253=>"00000001",
  56254=>"11111001",
  56255=>"11111101",
  56256=>"00000010",
  56257=>"11111101",
  56258=>"00000001",
  56259=>"11111100",
  56260=>"11111010",
  56261=>"11111010",
  56262=>"11111101",
  56263=>"11111100",
  56264=>"00001010",
  56265=>"11111110",
  56266=>"00000010",
  56267=>"11111010",
  56268=>"11111010",
  56269=>"11111111",
  56270=>"00000000",
  56271=>"00000010",
  56272=>"11110101",
  56273=>"11111110",
  56274=>"00000000",
  56275=>"11111001",
  56276=>"11111010",
  56277=>"00000011",
  56278=>"00000010",
  56279=>"00000101",
  56280=>"11111011",
  56281=>"11111111",
  56282=>"00000011",
  56283=>"11111011",
  56284=>"11111110",
  56285=>"00000010",
  56286=>"00000010",
  56287=>"00000000",
  56288=>"00000000",
  56289=>"11111100",
  56290=>"11111010",
  56291=>"11111010",
  56292=>"11111101",
  56293=>"11111111",
  56294=>"00000011",
  56295=>"11111111",
  56296=>"00000000",
  56297=>"11111011",
  56298=>"00000100",
  56299=>"00000000",
  56300=>"11111100",
  56301=>"00000010",
  56302=>"00000101",
  56303=>"11111101",
  56304=>"00000001",
  56305=>"11111100",
  56306=>"11111111",
  56307=>"11111101",
  56308=>"11111001",
  56309=>"00000101",
  56310=>"11111110",
  56311=>"11111101",
  56312=>"00000001",
  56313=>"11110001",
  56314=>"11111111",
  56315=>"11111101",
  56316=>"00000110",
  56317=>"00000011",
  56318=>"00000011",
  56319=>"11111001",
  56320=>"11111101",
  56321=>"00000010",
  56322=>"11111111",
  56323=>"00000000",
  56324=>"11111110",
  56325=>"11111110",
  56326=>"00000010",
  56327=>"11111110",
  56328=>"00000001",
  56329=>"00000000",
  56330=>"11111101",
  56331=>"00000001",
  56332=>"00000000",
  56333=>"00000001",
  56334=>"11111111",
  56335=>"11111101",
  56336=>"11111110",
  56337=>"00000010",
  56338=>"00000000",
  56339=>"11111101",
  56340=>"00000000",
  56341=>"00000001",
  56342=>"11111111",
  56343=>"11111101",
  56344=>"00000001",
  56345=>"00000010",
  56346=>"11111111",
  56347=>"11111111",
  56348=>"00000000",
  56349=>"11111110",
  56350=>"00000010",
  56351=>"00000100",
  56352=>"11111101",
  56353=>"11111110",
  56354=>"11111110",
  56355=>"11111111",
  56356=>"00000000",
  56357=>"00000000",
  56358=>"00000000",
  56359=>"11111110",
  56360=>"00000010",
  56361=>"11111111",
  56362=>"11111110",
  56363=>"11111111",
  56364=>"11111110",
  56365=>"11111110",
  56366=>"00000001",
  56367=>"00000010",
  56368=>"00000010",
  56369=>"11111110",
  56370=>"00000000",
  56371=>"11111111",
  56372=>"00000011",
  56373=>"00000010",
  56374=>"00000001",
  56375=>"00000001",
  56376=>"00000000",
  56377=>"11111100",
  56378=>"11111110",
  56379=>"00000000",
  56380=>"11111110",
  56381=>"11111110",
  56382=>"11111110",
  56383=>"11111110",
  56384=>"11111110",
  56385=>"11111111",
  56386=>"00000001",
  56387=>"00000010",
  56388=>"00000001",
  56389=>"11111110",
  56390=>"11111110",
  56391=>"00000000",
  56392=>"11111101",
  56393=>"11111110",
  56394=>"11111110",
  56395=>"11111111",
  56396=>"11111111",
  56397=>"00000011",
  56398=>"00000010",
  56399=>"11111110",
  56400=>"11111101",
  56401=>"11111111",
  56402=>"00000001",
  56403=>"11111101",
  56404=>"11111110",
  56405=>"00000000",
  56406=>"00000001",
  56407=>"00000011",
  56408=>"00000001",
  56409=>"11111101",
  56410=>"11111110",
  56411=>"00000000",
  56412=>"11111111",
  56413=>"11111111",
  56414=>"11111101",
  56415=>"00000011",
  56416=>"00000010",
  56417=>"00000001",
  56418=>"00000000",
  56419=>"00000001",
  56420=>"00000000",
  56421=>"00000001",
  56422=>"11111101",
  56423=>"11111110",
  56424=>"11111101",
  56425=>"00000001",
  56426=>"00000010",
  56427=>"00000000",
  56428=>"00000000",
  56429=>"00000010",
  56430=>"00000001",
  56431=>"11111111",
  56432=>"11111110",
  56433=>"00000001",
  56434=>"11111110",
  56435=>"00000010",
  56436=>"11111110",
  56437=>"11111110",
  56438=>"11111110",
  56439=>"00000011",
  56440=>"11111111",
  56441=>"11111111",
  56442=>"00000001",
  56443=>"00000010",
  56444=>"00000001",
  56445=>"11111111",
  56446=>"00000000",
  56447=>"11111110",
  56448=>"11111101",
  56449=>"11111110",
  56450=>"00000010",
  56451=>"11111111",
  56452=>"00000010",
  56453=>"00000001",
  56454=>"00000001",
  56455=>"00000100",
  56456=>"11111110",
  56457=>"00000000",
  56458=>"00000010",
  56459=>"11111110",
  56460=>"11111111",
  56461=>"11111111",
  56462=>"11111111",
  56463=>"00000000",
  56464=>"00000011",
  56465=>"00000011",
  56466=>"11111110",
  56467=>"11111101",
  56468=>"11111101",
  56469=>"00000000",
  56470=>"00000000",
  56471=>"11111110",
  56472=>"11111100",
  56473=>"11111111",
  56474=>"11111100",
  56475=>"00000001",
  56476=>"00000001",
  56477=>"11111111",
  56478=>"11111101",
  56479=>"00000011",
  56480=>"00000000",
  56481=>"00000011",
  56482=>"00000000",
  56483=>"11111111",
  56484=>"00000000",
  56485=>"11111111",
  56486=>"11111111",
  56487=>"00000010",
  56488=>"00000010",
  56489=>"00000001",
  56490=>"11111101",
  56491=>"11111111",
  56492=>"11111110",
  56493=>"00000000",
  56494=>"11111110",
  56495=>"11111110",
  56496=>"00000001",
  56497=>"11111110",
  56498=>"11111111",
  56499=>"00000000",
  56500=>"00000010",
  56501=>"11111110",
  56502=>"00000011",
  56503=>"00000001",
  56504=>"00000000",
  56505=>"00000011",
  56506=>"11111111",
  56507=>"11111110",
  56508=>"11111111",
  56509=>"11111111",
  56510=>"11111110",
  56511=>"00000011",
  56512=>"11111101",
  56513=>"00000000",
  56514=>"11111111",
  56515=>"00000001",
  56516=>"00000000",
  56517=>"00000010",
  56518=>"00000101",
  56519=>"00000000",
  56520=>"00000000",
  56521=>"11111111",
  56522=>"00000010",
  56523=>"00000010",
  56524=>"11111110",
  56525=>"11111101",
  56526=>"00000011",
  56527=>"00000100",
  56528=>"11111110",
  56529=>"11111110",
  56530=>"11111111",
  56531=>"00000010",
  56532=>"11111111",
  56533=>"11111110",
  56534=>"00000000",
  56535=>"00000001",
  56536=>"11111110",
  56537=>"11111101",
  56538=>"00000010",
  56539=>"00000001",
  56540=>"00000001",
  56541=>"11111101",
  56542=>"00000000",
  56543=>"00000001",
  56544=>"11111111",
  56545=>"00000001",
  56546=>"00000001",
  56547=>"11111110",
  56548=>"00000000",
  56549=>"11111111",
  56550=>"00000001",
  56551=>"11111110",
  56552=>"11111101",
  56553=>"00000000",
  56554=>"00000100",
  56555=>"11111111",
  56556=>"00000001",
  56557=>"00000001",
  56558=>"11111110",
  56559=>"11111101",
  56560=>"11111101",
  56561=>"00000010",
  56562=>"11111100",
  56563=>"00000010",
  56564=>"11111101",
  56565=>"00000001",
  56566=>"11111111",
  56567=>"11111110",
  56568=>"00000101",
  56569=>"11111111",
  56570=>"00000001",
  56571=>"11111111",
  56572=>"00000000",
  56573=>"00000010",
  56574=>"11111101",
  56575=>"00000110",
  56576=>"00000000",
  56577=>"00000001",
  56578=>"11111101",
  56579=>"11111100",
  56580=>"11111111",
  56581=>"00000010",
  56582=>"11111110",
  56583=>"00000001",
  56584=>"00000001",
  56585=>"11111110",
  56586=>"00000010",
  56587=>"00000000",
  56588=>"11111110",
  56589=>"11111100",
  56590=>"00000001",
  56591=>"11111110",
  56592=>"00000000",
  56593=>"00000001",
  56594=>"00000011",
  56595=>"00000000",
  56596=>"11111111",
  56597=>"00000001",
  56598=>"11111110",
  56599=>"00000000",
  56600=>"00000101",
  56601=>"00000010",
  56602=>"00000000",
  56603=>"11111111",
  56604=>"00000011",
  56605=>"00000100",
  56606=>"11111111",
  56607=>"00000101",
  56608=>"00000010",
  56609=>"11111111",
  56610=>"11111101",
  56611=>"11111111",
  56612=>"11111110",
  56613=>"11111101",
  56614=>"00000000",
  56615=>"11111101",
  56616=>"00000001",
  56617=>"11111110",
  56618=>"00000100",
  56619=>"00000000",
  56620=>"11111111",
  56621=>"11111111",
  56622=>"11111110",
  56623=>"11111101",
  56624=>"11111110",
  56625=>"11111101",
  56626=>"00000101",
  56627=>"11111111",
  56628=>"00000000",
  56629=>"00000010",
  56630=>"00000011",
  56631=>"00000000",
  56632=>"00000010",
  56633=>"11111111",
  56634=>"00000010",
  56635=>"11111111",
  56636=>"11111111",
  56637=>"11111110",
  56638=>"11111111",
  56639=>"11111111",
  56640=>"00000001",
  56641=>"11111111",
  56642=>"00000010",
  56643=>"11111111",
  56644=>"00000001",
  56645=>"11111111",
  56646=>"00000000",
  56647=>"11111110",
  56648=>"00000000",
  56649=>"11111111",
  56650=>"00000010",
  56651=>"11111110",
  56652=>"11111111",
  56653=>"11111110",
  56654=>"11111111",
  56655=>"11111111",
  56656=>"11111110",
  56657=>"11111110",
  56658=>"11111101",
  56659=>"00000000",
  56660=>"11111101",
  56661=>"00000001",
  56662=>"11111110",
  56663=>"00000001",
  56664=>"00000001",
  56665=>"11111110",
  56666=>"11111111",
  56667=>"00000000",
  56668=>"11111111",
  56669=>"00000001",
  56670=>"00000010",
  56671=>"11111111",
  56672=>"11111110",
  56673=>"00000000",
  56674=>"00000001",
  56675=>"00000000",
  56676=>"00000010",
  56677=>"00000010",
  56678=>"11111110",
  56679=>"00000000",
  56680=>"00000001",
  56681=>"11111110",
  56682=>"00000001",
  56683=>"11111110",
  56684=>"11111101",
  56685=>"00000011",
  56686=>"00000010",
  56687=>"11111111",
  56688=>"11111101",
  56689=>"00000010",
  56690=>"11111101",
  56691=>"11111101",
  56692=>"00000000",
  56693=>"00000000",
  56694=>"00000010",
  56695=>"00000001",
  56696=>"00000001",
  56697=>"11111110",
  56698=>"11111111",
  56699=>"11111111",
  56700=>"11111101",
  56701=>"11111111",
  56702=>"00000010",
  56703=>"11111110",
  56704=>"00000010",
  56705=>"00000011",
  56706=>"11111101",
  56707=>"00000010",
  56708=>"00000010",
  56709=>"11111101",
  56710=>"11111111",
  56711=>"00000000",
  56712=>"11111101",
  56713=>"11111101",
  56714=>"00000011",
  56715=>"11111111",
  56716=>"00000010",
  56717=>"00000010",
  56718=>"00000001",
  56719=>"00000010",
  56720=>"00000010",
  56721=>"00000001",
  56722=>"11111100",
  56723=>"00000010",
  56724=>"11111101",
  56725=>"11111101",
  56726=>"00000000",
  56727=>"11111101",
  56728=>"11111111",
  56729=>"00000011",
  56730=>"11111110",
  56731=>"00000010",
  56732=>"11111110",
  56733=>"00000010",
  56734=>"00000001",
  56735=>"11111110",
  56736=>"00000000",
  56737=>"00000001",
  56738=>"11111100",
  56739=>"11111111",
  56740=>"00000001",
  56741=>"11111111",
  56742=>"11111100",
  56743=>"00000010",
  56744=>"00000011",
  56745=>"11111110",
  56746=>"11111110",
  56747=>"11111111",
  56748=>"00000010",
  56749=>"00000010",
  56750=>"11111110",
  56751=>"00000001",
  56752=>"00000001",
  56753=>"11111110",
  56754=>"00000001",
  56755=>"00000010",
  56756=>"00000000",
  56757=>"00000100",
  56758=>"11111101",
  56759=>"00000010",
  56760=>"00000101",
  56761=>"11111110",
  56762=>"11111111",
  56763=>"00000001",
  56764=>"11111101",
  56765=>"11111101",
  56766=>"11111101",
  56767=>"00000001",
  56768=>"00000010",
  56769=>"11111110",
  56770=>"11111110",
  56771=>"00000010",
  56772=>"00000000",
  56773=>"11111110",
  56774=>"00000001",
  56775=>"00000010",
  56776=>"11111101",
  56777=>"00000011",
  56778=>"11111111",
  56779=>"11111101",
  56780=>"00000001",
  56781=>"00000001",
  56782=>"00000100",
  56783=>"00000001",
  56784=>"11111111",
  56785=>"11111111",
  56786=>"00000001",
  56787=>"00000001",
  56788=>"11111101",
  56789=>"00000000",
  56790=>"00000100",
  56791=>"00000010",
  56792=>"00000010",
  56793=>"00000100",
  56794=>"00000000",
  56795=>"00000101",
  56796=>"00000000",
  56797=>"00000000",
  56798=>"00000000",
  56799=>"00000001",
  56800=>"00000001",
  56801=>"00000001",
  56802=>"00000001",
  56803=>"11111110",
  56804=>"00000011",
  56805=>"11111111",
  56806=>"11111111",
  56807=>"11111101",
  56808=>"11111110",
  56809=>"11111110",
  56810=>"00000001",
  56811=>"00000000",
  56812=>"11111110",
  56813=>"11111110",
  56814=>"00000011",
  56815=>"11111110",
  56816=>"00000000",
  56817=>"00000000",
  56818=>"00000010",
  56819=>"00000001",
  56820=>"11111101",
  56821=>"00000000",
  56822=>"11111110",
  56823=>"00000101",
  56824=>"11111111",
  56825=>"00000001",
  56826=>"00000001",
  56827=>"00000010",
  56828=>"11111111",
  56829=>"11111111",
  56830=>"00000000",
  56831=>"11111110",
  56832=>"11111110",
  56833=>"11111110",
  56834=>"11111110",
  56835=>"11111101",
  56836=>"00000011",
  56837=>"00000000",
  56838=>"11111111",
  56839=>"11111101",
  56840=>"00000000",
  56841=>"00000000",
  56842=>"11111111",
  56843=>"00000001",
  56844=>"00000010",
  56845=>"11111110",
  56846=>"11111110",
  56847=>"11111110",
  56848=>"00000001",
  56849=>"00000111",
  56850=>"00000001",
  56851=>"00000001",
  56852=>"00000000",
  56853=>"00000010",
  56854=>"00000001",
  56855=>"00000110",
  56856=>"00000001",
  56857=>"11111111",
  56858=>"00000001",
  56859=>"11111111",
  56860=>"00000010",
  56861=>"11111100",
  56862=>"11111111",
  56863=>"00000010",
  56864=>"11111110",
  56865=>"00000000",
  56866=>"11111101",
  56867=>"00000110",
  56868=>"00000010",
  56869=>"11111110",
  56870=>"00000010",
  56871=>"11111111",
  56872=>"00000001",
  56873=>"11111111",
  56874=>"11111110",
  56875=>"00000000",
  56876=>"00000001",
  56877=>"11111110",
  56878=>"00000110",
  56879=>"11111110",
  56880=>"11111101",
  56881=>"00000000",
  56882=>"00000010",
  56883=>"00000000",
  56884=>"00000000",
  56885=>"00000000",
  56886=>"00000001",
  56887=>"11111110",
  56888=>"11111110",
  56889=>"11111101",
  56890=>"00000000",
  56891=>"00000010",
  56892=>"11111101",
  56893=>"00000000",
  56894=>"00000000",
  56895=>"11111111",
  56896=>"11111111",
  56897=>"00000001",
  56898=>"11111110",
  56899=>"11111101",
  56900=>"11111101",
  56901=>"11111101",
  56902=>"00000001",
  56903=>"00000101",
  56904=>"00000000",
  56905=>"00000010",
  56906=>"11111111",
  56907=>"00000010",
  56908=>"11111111",
  56909=>"11111110",
  56910=>"11111100",
  56911=>"11111111",
  56912=>"00000000",
  56913=>"00000010",
  56914=>"00000011",
  56915=>"00000010",
  56916=>"00000000",
  56917=>"00000001",
  56918=>"11111101",
  56919=>"00000011",
  56920=>"00000010",
  56921=>"00000010",
  56922=>"11111111",
  56923=>"00000001",
  56924=>"11111101",
  56925=>"11111110",
  56926=>"11111110",
  56927=>"11111111",
  56928=>"00000100",
  56929=>"11111111",
  56930=>"00000001",
  56931=>"00000110",
  56932=>"11111111",
  56933=>"11111111",
  56934=>"00000001",
  56935=>"00000101",
  56936=>"11111110",
  56937=>"00000000",
  56938=>"00000000",
  56939=>"11111111",
  56940=>"11111101",
  56941=>"00000000",
  56942=>"00000001",
  56943=>"00000001",
  56944=>"00000000",
  56945=>"00000000",
  56946=>"00000000",
  56947=>"11111110",
  56948=>"11111111",
  56949=>"00000000",
  56950=>"00000010",
  56951=>"00000010",
  56952=>"00000011",
  56953=>"11111110",
  56954=>"00000101",
  56955=>"00000010",
  56956=>"11111111",
  56957=>"00000001",
  56958=>"00000000",
  56959=>"11111111",
  56960=>"11111110",
  56961=>"11111111",
  56962=>"11111101",
  56963=>"00000000",
  56964=>"00000000",
  56965=>"00000011",
  56966=>"00000001",
  56967=>"00000010",
  56968=>"11111110",
  56969=>"11111110",
  56970=>"11111111",
  56971=>"11111111",
  56972=>"00000010",
  56973=>"00000010",
  56974=>"11111101",
  56975=>"00000000",
  56976=>"00000000",
  56977=>"11111111",
  56978=>"00000001",
  56979=>"00000001",
  56980=>"11111101",
  56981=>"00000001",
  56982=>"00000010",
  56983=>"00000110",
  56984=>"11111111",
  56985=>"11111111",
  56986=>"11111101",
  56987=>"00000000",
  56988=>"11111111",
  56989=>"11111111",
  56990=>"00000001",
  56991=>"00000001",
  56992=>"00000010",
  56993=>"00000100",
  56994=>"11111111",
  56995=>"00000001",
  56996=>"00000001",
  56997=>"00000100",
  56998=>"11111110",
  56999=>"00000100",
  57000=>"11111101",
  57001=>"00000000",
  57002=>"11111110",
  57003=>"11111101",
  57004=>"11111111",
  57005=>"11111111",
  57006=>"00000001",
  57007=>"11111110",
  57008=>"00000100",
  57009=>"00000000",
  57010=>"00000010",
  57011=>"00000001",
  57012=>"00000000",
  57013=>"00000101",
  57014=>"00000011",
  57015=>"11111111",
  57016=>"11111101",
  57017=>"00000001",
  57018=>"11111101",
  57019=>"00000000",
  57020=>"11111111",
  57021=>"00000001",
  57022=>"00000001",
  57023=>"11111111",
  57024=>"00000001",
  57025=>"11111110",
  57026=>"00000001",
  57027=>"00000000",
  57028=>"11111101",
  57029=>"00000010",
  57030=>"11111111",
  57031=>"11111101",
  57032=>"11111111",
  57033=>"00000000",
  57034=>"11111110",
  57035=>"00000001",
  57036=>"11111110",
  57037=>"11111101",
  57038=>"00000010",
  57039=>"00000010",
  57040=>"00000001",
  57041=>"00000011",
  57042=>"00000000",
  57043=>"11111110",
  57044=>"11111111",
  57045=>"11111111",
  57046=>"00000010",
  57047=>"00000001",
  57048=>"11111110",
  57049=>"00000010",
  57050=>"00000001",
  57051=>"00000010",
  57052=>"00000010",
  57053=>"00000000",
  57054=>"00000011",
  57055=>"11111111",
  57056=>"00000001",
  57057=>"00000001",
  57058=>"00000011",
  57059=>"00000101",
  57060=>"00000001",
  57061=>"11111111",
  57062=>"11111110",
  57063=>"11111101",
  57064=>"11111101",
  57065=>"11111111",
  57066=>"00000011",
  57067=>"11111101",
  57068=>"00000000",
  57069=>"00000101",
  57070=>"00000010",
  57071=>"00000000",
  57072=>"00000011",
  57073=>"00000000",
  57074=>"00000000",
  57075=>"11111110",
  57076=>"11111101",
  57077=>"00000000",
  57078=>"00000000",
  57079=>"11111111",
  57080=>"11111110",
  57081=>"00000000",
  57082=>"11111110",
  57083=>"11111101",
  57084=>"11111110",
  57085=>"11111111",
  57086=>"00000000",
  57087=>"00000010",
  57088=>"00000110",
  57089=>"11111111",
  57090=>"00000001",
  57091=>"11111111",
  57092=>"00000010",
  57093=>"00000010",
  57094=>"00000000",
  57095=>"00000001",
  57096=>"11111111",
  57097=>"11111111",
  57098=>"00000010",
  57099=>"00000001",
  57100=>"11111111",
  57101=>"00000100",
  57102=>"11111110",
  57103=>"11111110",
  57104=>"11111111",
  57105=>"00000010",
  57106=>"11111111",
  57107=>"11111111",
  57108=>"11111111",
  57109=>"11111101",
  57110=>"00000001",
  57111=>"00000010",
  57112=>"00000000",
  57113=>"11111101",
  57114=>"00000100",
  57115=>"11111111",
  57116=>"11111110",
  57117=>"00000000",
  57118=>"11111111",
  57119=>"00000001",
  57120=>"00000010",
  57121=>"11111111",
  57122=>"11111111",
  57123=>"00000000",
  57124=>"11111111",
  57125=>"00000010",
  57126=>"00000010",
  57127=>"00000000",
  57128=>"11111110",
  57129=>"11111110",
  57130=>"00000000",
  57131=>"00000001",
  57132=>"11111101",
  57133=>"00000001",
  57134=>"00000100",
  57135=>"11111111",
  57136=>"00000100",
  57137=>"11111101",
  57138=>"11111101",
  57139=>"11111101",
  57140=>"11111111",
  57141=>"00000010",
  57142=>"00000010",
  57143=>"00000000",
  57144=>"00000010",
  57145=>"00000010",
  57146=>"11111110",
  57147=>"11111111",
  57148=>"11111111",
  57149=>"00000000",
  57150=>"11111101",
  57151=>"11111110",
  57152=>"00000101",
  57153=>"11111111",
  57154=>"00000001",
  57155=>"11111101",
  57156=>"11111111",
  57157=>"11111111",
  57158=>"00000001",
  57159=>"00000010",
  57160=>"00000001",
  57161=>"11111111",
  57162=>"11111110",
  57163=>"00000000",
  57164=>"11111110",
  57165=>"00000001",
  57166=>"11111111",
  57167=>"00000010",
  57168=>"11111101",
  57169=>"11111111",
  57170=>"00000011",
  57171=>"11111110",
  57172=>"11111101",
  57173=>"00000011",
  57174=>"00000001",
  57175=>"11111110",
  57176=>"00000010",
  57177=>"11111101",
  57178=>"11111111",
  57179=>"00000001",
  57180=>"00000010",
  57181=>"11111111",
  57182=>"11111111",
  57183=>"11111111",
  57184=>"00000011",
  57185=>"11111101",
  57186=>"00000000",
  57187=>"11111101",
  57188=>"00000010",
  57189=>"11111111",
  57190=>"00000000",
  57191=>"11111110",
  57192=>"00000011",
  57193=>"00000010",
  57194=>"00000010",
  57195=>"11111101",
  57196=>"11111111",
  57197=>"11111101",
  57198=>"00000010",
  57199=>"11111111",
  57200=>"11111110",
  57201=>"00000010",
  57202=>"00000001",
  57203=>"00000000",
  57204=>"00000000",
  57205=>"00000000",
  57206=>"00000100",
  57207=>"00000001",
  57208=>"00000000",
  57209=>"11111101",
  57210=>"11111110",
  57211=>"11111110",
  57212=>"00000000",
  57213=>"00000000",
  57214=>"00000000",
  57215=>"11111110",
  57216=>"00000010",
  57217=>"11111110",
  57218=>"11111111",
  57219=>"11111110",
  57220=>"00000010",
  57221=>"00000001",
  57222=>"00000000",
  57223=>"00000001",
  57224=>"11111111",
  57225=>"00000000",
  57226=>"00000001",
  57227=>"00000010",
  57228=>"00000101",
  57229=>"00000000",
  57230=>"11111111",
  57231=>"11111111",
  57232=>"00000001",
  57233=>"11111101",
  57234=>"00000011",
  57235=>"11111111",
  57236=>"00000000",
  57237=>"00000001",
  57238=>"00000001",
  57239=>"11111101",
  57240=>"00000000",
  57241=>"00000100",
  57242=>"11111110",
  57243=>"11111110",
  57244=>"00000000",
  57245=>"00000011",
  57246=>"00000010",
  57247=>"11111111",
  57248=>"11111111",
  57249=>"11111110",
  57250=>"00000010",
  57251=>"11111110",
  57252=>"11111101",
  57253=>"00000000",
  57254=>"00000001",
  57255=>"00000000",
  57256=>"00000010",
  57257=>"00000011",
  57258=>"11111111",
  57259=>"00000001",
  57260=>"11111111",
  57261=>"00000001",
  57262=>"00000000",
  57263=>"11111101",
  57264=>"00000010",
  57265=>"11111111",
  57266=>"11111111",
  57267=>"11111110",
  57268=>"11111101",
  57269=>"11111101",
  57270=>"11111111",
  57271=>"00000100",
  57272=>"11111101",
  57273=>"00000001",
  57274=>"11111101",
  57275=>"00000000",
  57276=>"00000001",
  57277=>"00000101",
  57278=>"00000010",
  57279=>"00000010",
  57280=>"00000011",
  57281=>"00000001",
  57282=>"11111101",
  57283=>"00000001",
  57284=>"00000010",
  57285=>"11111110",
  57286=>"11111111",
  57287=>"00000010",
  57288=>"00000001",
  57289=>"00000010",
  57290=>"00000000",
  57291=>"11111111",
  57292=>"00000000",
  57293=>"00000011",
  57294=>"11111111",
  57295=>"11111110",
  57296=>"11111111",
  57297=>"00000011",
  57298=>"00000100",
  57299=>"11111111",
  57300=>"00000001",
  57301=>"11111101",
  57302=>"11111101",
  57303=>"00000001",
  57304=>"00000010",
  57305=>"11111110",
  57306=>"11111111",
  57307=>"11111111",
  57308=>"00000010",
  57309=>"00000000",
  57310=>"11111110",
  57311=>"00000000",
  57312=>"11111100",
  57313=>"00000000",
  57314=>"00000000",
  57315=>"11111101",
  57316=>"11111111",
  57317=>"00000001",
  57318=>"00000011",
  57319=>"11111110",
  57320=>"00000010",
  57321=>"11111110",
  57322=>"11111111",
  57323=>"11111111",
  57324=>"11111110",
  57325=>"00000000",
  57326=>"00000110",
  57327=>"00000000",
  57328=>"00000010",
  57329=>"11111110",
  57330=>"00000100",
  57331=>"00000001",
  57332=>"00000000",
  57333=>"11111110",
  57334=>"11111111",
  57335=>"11111101",
  57336=>"11111110",
  57337=>"00000001",
  57338=>"11111111",
  57339=>"11111111",
  57340=>"00000000",
  57341=>"00000010",
  57342=>"00000011",
  57343=>"11111110",
  57344=>"11111101",
  57345=>"00000000",
  57346=>"11111110",
  57347=>"00000001",
  57348=>"00000001",
  57349=>"11111100",
  57350=>"00000001",
  57351=>"11111101",
  57352=>"11111110",
  57353=>"11111111",
  57354=>"11111111",
  57355=>"11111111",
  57356=>"00000010",
  57357=>"00000000",
  57358=>"00000011",
  57359=>"11111111",
  57360=>"11111110",
  57361=>"00000011",
  57362=>"11111101",
  57363=>"00000000",
  57364=>"00000101",
  57365=>"11111111",
  57366=>"00000001",
  57367=>"11111101",
  57368=>"11111110",
  57369=>"00000100",
  57370=>"11111110",
  57371=>"11111111",
  57372=>"00000000",
  57373=>"11111111",
  57374=>"00000001",
  57375=>"00000000",
  57376=>"00000001",
  57377=>"00000101",
  57378=>"11111101",
  57379=>"11111110",
  57380=>"00000010",
  57381=>"00000001",
  57382=>"11111110",
  57383=>"11111110",
  57384=>"11111110",
  57385=>"11111110",
  57386=>"00000000",
  57387=>"00000010",
  57388=>"11111110",
  57389=>"11111111",
  57390=>"00000000",
  57391=>"00000010",
  57392=>"11111101",
  57393=>"11111111",
  57394=>"11111101",
  57395=>"00000001",
  57396=>"00000011",
  57397=>"00000001",
  57398=>"00000010",
  57399=>"11111110",
  57400=>"00000010",
  57401=>"00000000",
  57402=>"00000001",
  57403=>"00000010",
  57404=>"00000000",
  57405=>"11111101",
  57406=>"11111101",
  57407=>"11111111",
  57408=>"00000100",
  57409=>"11111101",
  57410=>"11111111",
  57411=>"00000010",
  57412=>"00000011",
  57413=>"00000001",
  57414=>"11111101",
  57415=>"00000001",
  57416=>"11111101",
  57417=>"00000011",
  57418=>"00000010",
  57419=>"00000000",
  57420=>"11111110",
  57421=>"11111111",
  57422=>"11111111",
  57423=>"11111110",
  57424=>"11111101",
  57425=>"11111111",
  57426=>"11111101",
  57427=>"00000011",
  57428=>"11111110",
  57429=>"00000011",
  57430=>"11111100",
  57431=>"11111110",
  57432=>"11111110",
  57433=>"00000000",
  57434=>"11111111",
  57435=>"00000011",
  57436=>"00000100",
  57437=>"00000000",
  57438=>"11111101",
  57439=>"11111111",
  57440=>"00000001",
  57441=>"00000000",
  57442=>"11111111",
  57443=>"00000000",
  57444=>"00000000",
  57445=>"00000000",
  57446=>"11111110",
  57447=>"00000000",
  57448=>"11111110",
  57449=>"00000000",
  57450=>"11111110",
  57451=>"00000001",
  57452=>"00000010",
  57453=>"00000011",
  57454=>"11111111",
  57455=>"00000001",
  57456=>"11111101",
  57457=>"00000000",
  57458=>"00000010",
  57459=>"11111110",
  57460=>"00000000",
  57461=>"00000000",
  57462=>"11111110",
  57463=>"00000001",
  57464=>"11111110",
  57465=>"00000011",
  57466=>"00000010",
  57467=>"00000001",
  57468=>"11111110",
  57469=>"00000000",
  57470=>"11111110",
  57471=>"00000001",
  57472=>"11111111",
  57473=>"00000000",
  57474=>"11111110",
  57475=>"00000010",
  57476=>"11111101",
  57477=>"00000000",
  57478=>"11111111",
  57479=>"11111110",
  57480=>"00000010",
  57481=>"00000001",
  57482=>"00000000",
  57483=>"00000010",
  57484=>"11111111",
  57485=>"11111111",
  57486=>"11111111",
  57487=>"11111110",
  57488=>"00000000",
  57489=>"11111110",
  57490=>"00000001",
  57491=>"11111101",
  57492=>"00000100",
  57493=>"11111100",
  57494=>"00000000",
  57495=>"11111101",
  57496=>"00000101",
  57497=>"11111110",
  57498=>"00000010",
  57499=>"11111100",
  57500=>"00000010",
  57501=>"00000010",
  57502=>"00000011",
  57503=>"11111111",
  57504=>"11111111",
  57505=>"00000000",
  57506=>"00000011",
  57507=>"00000000",
  57508=>"00000010",
  57509=>"00000000",
  57510=>"00000001",
  57511=>"00000100",
  57512=>"11111110",
  57513=>"00000000",
  57514=>"00000000",
  57515=>"00000000",
  57516=>"00000001",
  57517=>"11111101",
  57518=>"00000010",
  57519=>"00000000",
  57520=>"11111110",
  57521=>"00000000",
  57522=>"11111110",
  57523=>"11111110",
  57524=>"00000010",
  57525=>"11111110",
  57526=>"11111101",
  57527=>"00000000",
  57528=>"00000000",
  57529=>"11111101",
  57530=>"00000000",
  57531=>"00000000",
  57532=>"11111101",
  57533=>"00000000",
  57534=>"00000001",
  57535=>"00000000",
  57536=>"00000001",
  57537=>"00000001",
  57538=>"11111111",
  57539=>"11111111",
  57540=>"11111101",
  57541=>"11111101",
  57542=>"00000000",
  57543=>"11111110",
  57544=>"00000010",
  57545=>"00000010",
  57546=>"00000010",
  57547=>"11111110",
  57548=>"00000010",
  57549=>"00000001",
  57550=>"00000001",
  57551=>"11111101",
  57552=>"00000000",
  57553=>"11111101",
  57554=>"11111111",
  57555=>"00000010",
  57556=>"11111111",
  57557=>"00000011",
  57558=>"00000000",
  57559=>"00000001",
  57560=>"00000000",
  57561=>"00000001",
  57562=>"11111110",
  57563=>"00000010",
  57564=>"11111111",
  57565=>"00000010",
  57566=>"11111111",
  57567=>"00000010",
  57568=>"11111111",
  57569=>"00000000",
  57570=>"00000000",
  57571=>"00000000",
  57572=>"11111111",
  57573=>"00000001",
  57574=>"00000001",
  57575=>"11111110",
  57576=>"00000000",
  57577=>"00000000",
  57578=>"11111111",
  57579=>"00000000",
  57580=>"11111110",
  57581=>"11111110",
  57582=>"00000001",
  57583=>"11111111",
  57584=>"11111110",
  57585=>"11111101",
  57586=>"11111111",
  57587=>"00000001",
  57588=>"00000001",
  57589=>"11111111",
  57590=>"00000000",
  57591=>"00000001",
  57592=>"00000001",
  57593=>"00000000",
  57594=>"11111110",
  57595=>"00000001",
  57596=>"00000001",
  57597=>"00000000",
  57598=>"11111111",
  57599=>"00000010",
  57600=>"11111110",
  57601=>"11111100",
  57602=>"00000011",
  57603=>"00000000",
  57604=>"00000010",
  57605=>"11111111",
  57606=>"00000001",
  57607=>"11111111",
  57608=>"00000001",
  57609=>"11111111",
  57610=>"11111101",
  57611=>"00000011",
  57612=>"00000000",
  57613=>"00000010",
  57614=>"11111110",
  57615=>"11111110",
  57616=>"00000001",
  57617=>"11111110",
  57618=>"00000011",
  57619=>"11111111",
  57620=>"00000000",
  57621=>"11111110",
  57622=>"11111111",
  57623=>"11111110",
  57624=>"00000010",
  57625=>"11111111",
  57626=>"00000001",
  57627=>"11111111",
  57628=>"11111100",
  57629=>"11111111",
  57630=>"11111101",
  57631=>"11111101",
  57632=>"00000000",
  57633=>"00000001",
  57634=>"00000001",
  57635=>"11111110",
  57636=>"00000001",
  57637=>"00000001",
  57638=>"00000010",
  57639=>"11111111",
  57640=>"11111101",
  57641=>"00000100",
  57642=>"00000000",
  57643=>"00000011",
  57644=>"11111111",
  57645=>"00000001",
  57646=>"00000010",
  57647=>"11111110",
  57648=>"11111100",
  57649=>"00000000",
  57650=>"00000101",
  57651=>"00000001",
  57652=>"00000000",
  57653=>"11111011",
  57654=>"00000011",
  57655=>"00000010",
  57656=>"00000000",
  57657=>"00000001",
  57658=>"00000001",
  57659=>"11111111",
  57660=>"11111101",
  57661=>"00000010",
  57662=>"00000010",
  57663=>"11111111",
  57664=>"00000000",
  57665=>"00000000",
  57666=>"00000001",
  57667=>"11111111",
  57668=>"11111110",
  57669=>"11111111",
  57670=>"11111100",
  57671=>"00000000",
  57672=>"11111110",
  57673=>"00000000",
  57674=>"11111100",
  57675=>"00000001",
  57676=>"00000000",
  57677=>"00000010",
  57678=>"00000100",
  57679=>"11111111",
  57680=>"11111111",
  57681=>"00000011",
  57682=>"11111110",
  57683=>"11111110",
  57684=>"00000010",
  57685=>"11111110",
  57686=>"00000010",
  57687=>"11111111",
  57688=>"00000011",
  57689=>"00000001",
  57690=>"11111110",
  57691=>"00000001",
  57692=>"00000000",
  57693=>"00000010",
  57694=>"11111110",
  57695=>"11111101",
  57696=>"11111110",
  57697=>"00000010",
  57698=>"00000000",
  57699=>"11111111",
  57700=>"11111111",
  57701=>"00000001",
  57702=>"00000010",
  57703=>"00000000",
  57704=>"00000000",
  57705=>"00000001",
  57706=>"11111110",
  57707=>"00000010",
  57708=>"00000000",
  57709=>"11111101",
  57710=>"11111111",
  57711=>"11111101",
  57712=>"00000010",
  57713=>"11111111",
  57714=>"11111111",
  57715=>"00000101",
  57716=>"00000000",
  57717=>"11111101",
  57718=>"11111111",
  57719=>"11111110",
  57720=>"00000001",
  57721=>"00000010",
  57722=>"11111100",
  57723=>"00000001",
  57724=>"11111110",
  57725=>"11111101",
  57726=>"00000000",
  57727=>"00000001",
  57728=>"11111111",
  57729=>"11111100",
  57730=>"11111110",
  57731=>"11111111",
  57732=>"00000001",
  57733=>"00000111",
  57734=>"00000001",
  57735=>"11111110",
  57736=>"00000010",
  57737=>"11111101",
  57738=>"00000001",
  57739=>"11111111",
  57740=>"11111110",
  57741=>"11111110",
  57742=>"11111111",
  57743=>"11111110",
  57744=>"00000000",
  57745=>"00000010",
  57746=>"11111110",
  57747=>"11111110",
  57748=>"11111100",
  57749=>"00000001",
  57750=>"00000000",
  57751=>"00000010",
  57752=>"11111101",
  57753=>"11111110",
  57754=>"11111101",
  57755=>"00000000",
  57756=>"00000010",
  57757=>"00000000",
  57758=>"11111101",
  57759=>"00000001",
  57760=>"00000001",
  57761=>"11111111",
  57762=>"11111111",
  57763=>"11111110",
  57764=>"11111110",
  57765=>"11111110",
  57766=>"11111111",
  57767=>"00000010",
  57768=>"00000001",
  57769=>"11111110",
  57770=>"11111111",
  57771=>"00000000",
  57772=>"11111111",
  57773=>"00000001",
  57774=>"11111111",
  57775=>"11111101",
  57776=>"00000000",
  57777=>"00000001",
  57778=>"11111101",
  57779=>"00000001",
  57780=>"00000010",
  57781=>"00000000",
  57782=>"11111110",
  57783=>"11111110",
  57784=>"00000010",
  57785=>"11111111",
  57786=>"00000010",
  57787=>"00000000",
  57788=>"00000010",
  57789=>"00000100",
  57790=>"11111110",
  57791=>"11111111",
  57792=>"11111101",
  57793=>"00000010",
  57794=>"00000000",
  57795=>"11111111",
  57796=>"11111101",
  57797=>"11111101",
  57798=>"11111101",
  57799=>"11111110",
  57800=>"11111111",
  57801=>"11111111",
  57802=>"00000011",
  57803=>"00000010",
  57804=>"11111110",
  57805=>"00000001",
  57806=>"00000010",
  57807=>"00000001",
  57808=>"11111110",
  57809=>"00000010",
  57810=>"11111111",
  57811=>"00000010",
  57812=>"11111111",
  57813=>"00000010",
  57814=>"11111101",
  57815=>"11111110",
  57816=>"11111110",
  57817=>"00000101",
  57818=>"00000001",
  57819=>"11111101",
  57820=>"00000010",
  57821=>"11111111",
  57822=>"00000000",
  57823=>"00000100",
  57824=>"00000011",
  57825=>"11111110",
  57826=>"11111110",
  57827=>"00000011",
  57828=>"11111110",
  57829=>"00000001",
  57830=>"11111111",
  57831=>"00000000",
  57832=>"00000110",
  57833=>"11111110",
  57834=>"11111110",
  57835=>"11111100",
  57836=>"00000010",
  57837=>"11111110",
  57838=>"00000001",
  57839=>"11111100",
  57840=>"11111110",
  57841=>"11111110",
  57842=>"00000001",
  57843=>"00000000",
  57844=>"11111100",
  57845=>"00000000",
  57846=>"00000010",
  57847=>"11111111",
  57848=>"11111111",
  57849=>"00000001",
  57850=>"00000000",
  57851=>"11111110",
  57852=>"00000000",
  57853=>"00000011",
  57854=>"11111101",
  57855=>"00000000",
  57856=>"11111110",
  57857=>"11111111",
  57858=>"00000110",
  57859=>"11111111",
  57860=>"00000010",
  57861=>"11111101",
  57862=>"00000110",
  57863=>"11111111",
  57864=>"11111111",
  57865=>"11111111",
  57866=>"00000000",
  57867=>"11111110",
  57868=>"11111111",
  57869=>"11111111",
  57870=>"11111101",
  57871=>"00000000",
  57872=>"00000001",
  57873=>"00000010",
  57874=>"00000100",
  57875=>"00000010",
  57876=>"11111111",
  57877=>"00000001",
  57878=>"00000011",
  57879=>"00000011",
  57880=>"11111101",
  57881=>"11111110",
  57882=>"11111110",
  57883=>"00000010",
  57884=>"11111110",
  57885=>"00000001",
  57886=>"00000000",
  57887=>"11111111",
  57888=>"00000010",
  57889=>"11111110",
  57890=>"00000010",
  57891=>"11111111",
  57892=>"11111110",
  57893=>"00000001",
  57894=>"11111101",
  57895=>"00000001",
  57896=>"11111101",
  57897=>"00000011",
  57898=>"11111111",
  57899=>"00000000",
  57900=>"11111110",
  57901=>"00000001",
  57902=>"11111101",
  57903=>"00000100",
  57904=>"11111111",
  57905=>"11111110",
  57906=>"11111111",
  57907=>"00000100",
  57908=>"00000001",
  57909=>"11111101",
  57910=>"00000010",
  57911=>"00000010",
  57912=>"11111111",
  57913=>"00000011",
  57914=>"00000000",
  57915=>"00000100",
  57916=>"11111111",
  57917=>"11111101",
  57918=>"11111110",
  57919=>"00000001",
  57920=>"11111110",
  57921=>"11111101",
  57922=>"11111111",
  57923=>"00000000",
  57924=>"00000010",
  57925=>"11111110",
  57926=>"11111100",
  57927=>"11111101",
  57928=>"11111101",
  57929=>"00000001",
  57930=>"00000010",
  57931=>"11111101",
  57932=>"11111111",
  57933=>"00000011",
  57934=>"00000011",
  57935=>"11111101",
  57936=>"11111110",
  57937=>"11111100",
  57938=>"00000010",
  57939=>"00000001",
  57940=>"00000000",
  57941=>"00000011",
  57942=>"00000010",
  57943=>"00000010",
  57944=>"00000010",
  57945=>"11111111",
  57946=>"00000000",
  57947=>"00000001",
  57948=>"11111111",
  57949=>"00000010",
  57950=>"00000001",
  57951=>"00000001",
  57952=>"00000100",
  57953=>"11111101",
  57954=>"11111110",
  57955=>"00000010",
  57956=>"00000001",
  57957=>"11111110",
  57958=>"11111101",
  57959=>"11111111",
  57960=>"11111110",
  57961=>"00000010",
  57962=>"00000010",
  57963=>"00000001",
  57964=>"00000100",
  57965=>"00000001",
  57966=>"00000010",
  57967=>"00000000",
  57968=>"00000010",
  57969=>"00000000",
  57970=>"00000000",
  57971=>"11111101",
  57972=>"00000000",
  57973=>"11111110",
  57974=>"11111100",
  57975=>"11111101",
  57976=>"00000000",
  57977=>"00000000",
  57978=>"00000010",
  57979=>"11111101",
  57980=>"11111111",
  57981=>"00000001",
  57982=>"00000010",
  57983=>"00000000",
  57984=>"00000001",
  57985=>"11111110",
  57986=>"11111111",
  57987=>"11111110",
  57988=>"00000010",
  57989=>"00000000",
  57990=>"00000101",
  57991=>"00000010",
  57992=>"11111110",
  57993=>"00000000",
  57994=>"11111111",
  57995=>"00000111",
  57996=>"11111111",
  57997=>"00000010",
  57998=>"00000001",
  57999=>"11111101",
  58000=>"11111111",
  58001=>"11111110",
  58002=>"11111111",
  58003=>"00000010",
  58004=>"00000010",
  58005=>"11111111",
  58006=>"11111110",
  58007=>"00000101",
  58008=>"00000111",
  58009=>"11111101",
  58010=>"11111101",
  58011=>"11111111",
  58012=>"00000100",
  58013=>"00000010",
  58014=>"00000010",
  58015=>"00000010",
  58016=>"11111110",
  58017=>"11111101",
  58018=>"00000100",
  58019=>"00000010",
  58020=>"00000000",
  58021=>"00000010",
  58022=>"00000001",
  58023=>"00000010",
  58024=>"00000010",
  58025=>"00000011",
  58026=>"00000101",
  58027=>"00000010",
  58028=>"00000010",
  58029=>"00000000",
  58030=>"11111110",
  58031=>"11111111",
  58032=>"00000001",
  58033=>"11111111",
  58034=>"11111110",
  58035=>"11111101",
  58036=>"00000001",
  58037=>"11111111",
  58038=>"11111110",
  58039=>"00000000",
  58040=>"11111111",
  58041=>"11111110",
  58042=>"11111101",
  58043=>"11111101",
  58044=>"11111101",
  58045=>"00000010",
  58046=>"00000000",
  58047=>"11111111",
  58048=>"11111110",
  58049=>"00000001",
  58050=>"11111100",
  58051=>"00000001",
  58052=>"00000001",
  58053=>"00000000",
  58054=>"00000010",
  58055=>"11111110",
  58056=>"11111111",
  58057=>"00000000",
  58058=>"11111101",
  58059=>"11111110",
  58060=>"00000110",
  58061=>"11111110",
  58062=>"00000000",
  58063=>"00000001",
  58064=>"00000000",
  58065=>"00000011",
  58066=>"00000001",
  58067=>"11111101",
  58068=>"11111110",
  58069=>"00000001",
  58070=>"00000010",
  58071=>"00000000",
  58072=>"11111100",
  58073=>"00000010",
  58074=>"00000001",
  58075=>"11111101",
  58076=>"00000101",
  58077=>"11111111",
  58078=>"11111111",
  58079=>"11111100",
  58080=>"00000000",
  58081=>"11111110",
  58082=>"00000011",
  58083=>"00000011",
  58084=>"00000011",
  58085=>"00000001",
  58086=>"00000010",
  58087=>"00000001",
  58088=>"11111101",
  58089=>"00000001",
  58090=>"11111111",
  58091=>"11111110",
  58092=>"11111110",
  58093=>"11111101",
  58094=>"00000001",
  58095=>"00000001",
  58096=>"00000001",
  58097=>"00000000",
  58098=>"00000010",
  58099=>"11111110",
  58100=>"11111111",
  58101=>"00000011",
  58102=>"00000001",
  58103=>"11111111",
  58104=>"11111111",
  58105=>"11111111",
  58106=>"00000000",
  58107=>"00000001",
  58108=>"00000010",
  58109=>"00000011",
  58110=>"00000000",
  58111=>"00000010",
  58112=>"00000000",
  58113=>"11111111",
  58114=>"00000001",
  58115=>"11111110",
  58116=>"11111101",
  58117=>"00000000",
  58118=>"00000000",
  58119=>"11111110",
  58120=>"11111110",
  58121=>"00000001",
  58122=>"00000000",
  58123=>"00000000",
  58124=>"00000101",
  58125=>"11111111",
  58126=>"11111110",
  58127=>"00000010",
  58128=>"00000010",
  58129=>"00000011",
  58130=>"11111101",
  58131=>"11111110",
  58132=>"00000001",
  58133=>"00000001",
  58134=>"00000011",
  58135=>"11111110",
  58136=>"11111101",
  58137=>"11111110",
  58138=>"00000001",
  58139=>"11111100",
  58140=>"11111101",
  58141=>"11111101",
  58142=>"00000001",
  58143=>"11111111",
  58144=>"00000000",
  58145=>"00000000",
  58146=>"00000000",
  58147=>"00000010",
  58148=>"00000010",
  58149=>"00001000",
  58150=>"00000100",
  58151=>"11111100",
  58152=>"00000010",
  58153=>"11111110",
  58154=>"11111110",
  58155=>"00000010",
  58156=>"00000001",
  58157=>"00000000",
  58158=>"00000001",
  58159=>"11111111",
  58160=>"11111110",
  58161=>"00000001",
  58162=>"00000010",
  58163=>"00000010",
  58164=>"00000000",
  58165=>"11111111",
  58166=>"11111110",
  58167=>"00000010",
  58168=>"00000001",
  58169=>"00000010",
  58170=>"00000011",
  58171=>"11111110",
  58172=>"11111110",
  58173=>"00000000",
  58174=>"00000001",
  58175=>"00000001",
  58176=>"11111101",
  58177=>"11111110",
  58178=>"11111111",
  58179=>"00000000",
  58180=>"11111101",
  58181=>"00000000",
  58182=>"00000010",
  58183=>"00000100",
  58184=>"00000010",
  58185=>"11111111",
  58186=>"00000001",
  58187=>"00000000",
  58188=>"00000000",
  58189=>"00000000",
  58190=>"11111101",
  58191=>"00000001",
  58192=>"11111111",
  58193=>"11111110",
  58194=>"00000010",
  58195=>"00000010",
  58196=>"00000000",
  58197=>"11111101",
  58198=>"00000000",
  58199=>"00000000",
  58200=>"00001000",
  58201=>"11111110",
  58202=>"00000100",
  58203=>"11111100",
  58204=>"00000100",
  58205=>"11111111",
  58206=>"00000010",
  58207=>"00000011",
  58208=>"11111111",
  58209=>"11111110",
  58210=>"00000001",
  58211=>"00000010",
  58212=>"00000001",
  58213=>"00000000",
  58214=>"00000010",
  58215=>"00000001",
  58216=>"00000000",
  58217=>"11111111",
  58218=>"11111111",
  58219=>"11111101",
  58220=>"11111110",
  58221=>"00000000",
  58222=>"11111111",
  58223=>"11111111",
  58224=>"00000001",
  58225=>"00000001",
  58226=>"00000000",
  58227=>"11111111",
  58228=>"00000011",
  58229=>"00000010",
  58230=>"00000011",
  58231=>"00000010",
  58232=>"11111101",
  58233=>"00000011",
  58234=>"00000101",
  58235=>"11111101",
  58236=>"11111110",
  58237=>"00000011",
  58238=>"11111101",
  58239=>"00000001",
  58240=>"11111110",
  58241=>"00000010",
  58242=>"11111111",
  58243=>"11111101",
  58244=>"11111110",
  58245=>"11111101",
  58246=>"00000001",
  58247=>"00000100",
  58248=>"11111111",
  58249=>"11111110",
  58250=>"11111101",
  58251=>"00000001",
  58252=>"00000010",
  58253=>"11111110",
  58254=>"11111101",
  58255=>"11111110",
  58256=>"11111101",
  58257=>"11111111",
  58258=>"11111111",
  58259=>"00000011",
  58260=>"11111110",
  58261=>"11111110",
  58262=>"00000001",
  58263=>"00000000",
  58264=>"11111101",
  58265=>"00000011",
  58266=>"00000001",
  58267=>"11111111",
  58268=>"00000001",
  58269=>"00000010",
  58270=>"11111101",
  58271=>"00000101",
  58272=>"00000000",
  58273=>"00000001",
  58274=>"00000001",
  58275=>"00000010",
  58276=>"00000001",
  58277=>"00000010",
  58278=>"00000001",
  58279=>"11111111",
  58280=>"00000010",
  58281=>"00000010",
  58282=>"00000011",
  58283=>"00000000",
  58284=>"00000001",
  58285=>"11111101",
  58286=>"00000001",
  58287=>"00000001",
  58288=>"00000010",
  58289=>"11111110",
  58290=>"00000010",
  58291=>"00000001",
  58292=>"00000010",
  58293=>"00000000",
  58294=>"00000000",
  58295=>"00000101",
  58296=>"00000000",
  58297=>"11111111",
  58298=>"11111110",
  58299=>"11111111",
  58300=>"11111110",
  58301=>"11111111",
  58302=>"11111110",
  58303=>"00000001",
  58304=>"11111100",
  58305=>"11111110",
  58306=>"00000001",
  58307=>"00000001",
  58308=>"00000011",
  58309=>"11111110",
  58310=>"11111101",
  58311=>"00000000",
  58312=>"00000010",
  58313=>"11111110",
  58314=>"11111101",
  58315=>"00000001",
  58316=>"11111110",
  58317=>"00000001",
  58318=>"11111111",
  58319=>"00000000",
  58320=>"00000011",
  58321=>"11111111",
  58322=>"11111111",
  58323=>"11111111",
  58324=>"00000001",
  58325=>"11111101",
  58326=>"11111101",
  58327=>"11111111",
  58328=>"11111111",
  58329=>"11111110",
  58330=>"00000001",
  58331=>"11111111",
  58332=>"00000010",
  58333=>"00000101",
  58334=>"11111110",
  58335=>"00000101",
  58336=>"11111101",
  58337=>"00000001",
  58338=>"00000000",
  58339=>"00000011",
  58340=>"00000010",
  58341=>"00000001",
  58342=>"00000001",
  58343=>"00000001",
  58344=>"00000001",
  58345=>"00000001",
  58346=>"00000000",
  58347=>"00000001",
  58348=>"00000000",
  58349=>"00000001",
  58350=>"11111110",
  58351=>"11111110",
  58352=>"00000001",
  58353=>"00000010",
  58354=>"00000001",
  58355=>"11111111",
  58356=>"00000010",
  58357=>"00000010",
  58358=>"00000000",
  58359=>"00000000",
  58360=>"11111101",
  58361=>"00000000",
  58362=>"00000001",
  58363=>"00000101",
  58364=>"00000011",
  58365=>"00000011",
  58366=>"00000000",
  58367=>"00000001",
  58368=>"00000100",
  58369=>"11111101",
  58370=>"00000010",
  58371=>"11111111",
  58372=>"00000001",
  58373=>"11111101",
  58374=>"00000000",
  58375=>"00000000",
  58376=>"00000010",
  58377=>"00000000",
  58378=>"00000000",
  58379=>"11111110",
  58380=>"00000001",
  58381=>"00000100",
  58382=>"11111101",
  58383=>"11111101",
  58384=>"00000101",
  58385=>"00000010",
  58386=>"00000001",
  58387=>"00000001",
  58388=>"00000000",
  58389=>"00000001",
  58390=>"00000101",
  58391=>"00000011",
  58392=>"11111110",
  58393=>"00000000",
  58394=>"00000000",
  58395=>"00000010",
  58396=>"00000001",
  58397=>"11111101",
  58398=>"11111111",
  58399=>"11111111",
  58400=>"11111110",
  58401=>"00000000",
  58402=>"00000010",
  58403=>"11111100",
  58404=>"00000000",
  58405=>"11111110",
  58406=>"00000001",
  58407=>"11111110",
  58408=>"00000010",
  58409=>"11111011",
  58410=>"11111111",
  58411=>"11111111",
  58412=>"00000011",
  58413=>"00000011",
  58414=>"00000000",
  58415=>"00000010",
  58416=>"00000010",
  58417=>"11111110",
  58418=>"00000000",
  58419=>"00000000",
  58420=>"00000010",
  58421=>"00000001",
  58422=>"11111110",
  58423=>"11111101",
  58424=>"00000001",
  58425=>"00000000",
  58426=>"00000011",
  58427=>"00000001",
  58428=>"11111111",
  58429=>"00000000",
  58430=>"00000010",
  58431=>"00000000",
  58432=>"00000000",
  58433=>"00000011",
  58434=>"00000010",
  58435=>"11111110",
  58436=>"00000011",
  58437=>"00000000",
  58438=>"00000010",
  58439=>"00000010",
  58440=>"00000000",
  58441=>"11111110",
  58442=>"11111101",
  58443=>"11111111",
  58444=>"11111111",
  58445=>"11111111",
  58446=>"11111110",
  58447=>"11111101",
  58448=>"00000000",
  58449=>"11111111",
  58450=>"11111101",
  58451=>"00000000",
  58452=>"00000000",
  58453=>"00000001",
  58454=>"00000001",
  58455=>"00000010",
  58456=>"00000100",
  58457=>"00000010",
  58458=>"11111111",
  58459=>"00000001",
  58460=>"00000101",
  58461=>"11111110",
  58462=>"11111111",
  58463=>"00000001",
  58464=>"00000001",
  58465=>"00000010",
  58466=>"00000001",
  58467=>"11111111",
  58468=>"11111111",
  58469=>"00000000",
  58470=>"11111110",
  58471=>"00000001",
  58472=>"00000010",
  58473=>"11111110",
  58474=>"00000000",
  58475=>"00000001",
  58476=>"00000010",
  58477=>"11111111",
  58478=>"00000001",
  58479=>"00000010",
  58480=>"11111110",
  58481=>"11111110",
  58482=>"00000011",
  58483=>"00000010",
  58484=>"00000001",
  58485=>"11111111",
  58486=>"11111111",
  58487=>"00000010",
  58488=>"00000011",
  58489=>"11111110",
  58490=>"11111110",
  58491=>"00000011",
  58492=>"11111111",
  58493=>"11111111",
  58494=>"00000001",
  58495=>"11111100",
  58496=>"00000000",
  58497=>"11111111",
  58498=>"11111111",
  58499=>"00000000",
  58500=>"00000001",
  58501=>"00000001",
  58502=>"11111111",
  58503=>"11111111",
  58504=>"11111101",
  58505=>"00000101",
  58506=>"11111111",
  58507=>"11111100",
  58508=>"11111110",
  58509=>"00000010",
  58510=>"11111110",
  58511=>"11111101",
  58512=>"11111110",
  58513=>"11111110",
  58514=>"11111111",
  58515=>"00000010",
  58516=>"00000010",
  58517=>"00000100",
  58518=>"00000000",
  58519=>"00000001",
  58520=>"00000110",
  58521=>"00000101",
  58522=>"00000011",
  58523=>"11111101",
  58524=>"11111111",
  58525=>"00000000",
  58526=>"11111111",
  58527=>"11111110",
  58528=>"00000010",
  58529=>"00000100",
  58530=>"00000110",
  58531=>"00000001",
  58532=>"00000010",
  58533=>"00000001",
  58534=>"11111110",
  58535=>"11111101",
  58536=>"11111111",
  58537=>"11111111",
  58538=>"11111100",
  58539=>"00000001",
  58540=>"11111111",
  58541=>"00000000",
  58542=>"11111101",
  58543=>"00000010",
  58544=>"00000001",
  58545=>"11111110",
  58546=>"00000001",
  58547=>"00000001",
  58548=>"11111100",
  58549=>"11111111",
  58550=>"11111111",
  58551=>"11111101",
  58552=>"11111111",
  58553=>"11111110",
  58554=>"11111101",
  58555=>"00000000",
  58556=>"00000100",
  58557=>"00000001",
  58558=>"00000011",
  58559=>"00000010",
  58560=>"00000010",
  58561=>"00000011",
  58562=>"00000010",
  58563=>"11111101",
  58564=>"00000001",
  58565=>"11111110",
  58566=>"11111101",
  58567=>"00000001",
  58568=>"00000000",
  58569=>"11111101",
  58570=>"11111111",
  58571=>"11111100",
  58572=>"00000001",
  58573=>"11111111",
  58574=>"00000001",
  58575=>"11111111",
  58576=>"00000000",
  58577=>"11111110",
  58578=>"11111111",
  58579=>"00000100",
  58580=>"00000010",
  58581=>"00000000",
  58582=>"11111100",
  58583=>"11111011",
  58584=>"11111101",
  58585=>"11111111",
  58586=>"00000001",
  58587=>"11111110",
  58588=>"11111101",
  58589=>"11111111",
  58590=>"11111100",
  58591=>"00000000",
  58592=>"00000001",
  58593=>"00000011",
  58594=>"00000100",
  58595=>"00000100",
  58596=>"00000001",
  58597=>"11111101",
  58598=>"00000011",
  58599=>"00000000",
  58600=>"00000000",
  58601=>"11111111",
  58602=>"11111111",
  58603=>"11111110",
  58604=>"00000000",
  58605=>"11111100",
  58606=>"00000001",
  58607=>"11111110",
  58608=>"11111110",
  58609=>"11111110",
  58610=>"11111101",
  58611=>"11111110",
  58612=>"00000001",
  58613=>"11111100",
  58614=>"11111110",
  58615=>"11111100",
  58616=>"11111111",
  58617=>"00000010",
  58618=>"11111110",
  58619=>"00000001",
  58620=>"11111111",
  58621=>"11111111",
  58622=>"11111101",
  58623=>"00000011",
  58624=>"11111110",
  58625=>"11111011",
  58626=>"00000101",
  58627=>"11111101",
  58628=>"11111110",
  58629=>"00000000",
  58630=>"00000000",
  58631=>"00000000",
  58632=>"00000001",
  58633=>"00000011",
  58634=>"00000001",
  58635=>"11111110",
  58636=>"11111101",
  58637=>"11111111",
  58638=>"11111111",
  58639=>"11111111",
  58640=>"00000011",
  58641=>"11111111",
  58642=>"00000010",
  58643=>"00000001",
  58644=>"11111110",
  58645=>"00000100",
  58646=>"00000100",
  58647=>"11111101",
  58648=>"00000101",
  58649=>"11111101",
  58650=>"00000011",
  58651=>"00000011",
  58652=>"00000000",
  58653=>"11111110",
  58654=>"00000101",
  58655=>"00000100",
  58656=>"11111111",
  58657=>"00000010",
  58658=>"00000001",
  58659=>"11111111",
  58660=>"11111101",
  58661=>"11111100",
  58662=>"00000111",
  58663=>"11111100",
  58664=>"00000010",
  58665=>"00000001",
  58666=>"11111110",
  58667=>"00000011",
  58668=>"11111111",
  58669=>"00000001",
  58670=>"11111111",
  58671=>"00000000",
  58672=>"11111111",
  58673=>"11111101",
  58674=>"11111111",
  58675=>"00000011",
  58676=>"00000010",
  58677=>"11111101",
  58678=>"00000010",
  58679=>"00000001",
  58680=>"11111111",
  58681=>"11111110",
  58682=>"00000001",
  58683=>"00000011",
  58684=>"00000000",
  58685=>"00000000",
  58686=>"00000000",
  58687=>"00000001",
  58688=>"11111111",
  58689=>"11111110",
  58690=>"11111100",
  58691=>"00000000",
  58692=>"00000000",
  58693=>"00000011",
  58694=>"00000000",
  58695=>"00000001",
  58696=>"00000001",
  58697=>"00000100",
  58698=>"11111111",
  58699=>"00000100",
  58700=>"00000000",
  58701=>"00000001",
  58702=>"00000011",
  58703=>"00000000",
  58704=>"11111110",
  58705=>"00000000",
  58706=>"11111111",
  58707=>"00000101",
  58708=>"00000001",
  58709=>"11111110",
  58710=>"00000011",
  58711=>"11111110",
  58712=>"00000001",
  58713=>"11111110",
  58714=>"11111101",
  58715=>"11111111",
  58716=>"00000000",
  58717=>"00000000",
  58718=>"11111110",
  58719=>"00000001",
  58720=>"00000101",
  58721=>"11111110",
  58722=>"00000000",
  58723=>"11111111",
  58724=>"11111101",
  58725=>"11111111",
  58726=>"00000001",
  58727=>"00000010",
  58728=>"11111110",
  58729=>"11111110",
  58730=>"00000001",
  58731=>"00000010",
  58732=>"11111100",
  58733=>"11111111",
  58734=>"00000001",
  58735=>"11111101",
  58736=>"00000011",
  58737=>"00000010",
  58738=>"11111101",
  58739=>"00000001",
  58740=>"11111101",
  58741=>"00000100",
  58742=>"00000001",
  58743=>"00000011",
  58744=>"00000010",
  58745=>"00000001",
  58746=>"11111111",
  58747=>"00000000",
  58748=>"00000000",
  58749=>"11111111",
  58750=>"00000000",
  58751=>"11111110",
  58752=>"00000001",
  58753=>"11111011",
  58754=>"00000001",
  58755=>"11111111",
  58756=>"00000000",
  58757=>"11111110",
  58758=>"11111101",
  58759=>"11111111",
  58760=>"00000001",
  58761=>"00000100",
  58762=>"11111111",
  58763=>"00000000",
  58764=>"11111110",
  58765=>"00000010",
  58766=>"00000001",
  58767=>"11111101",
  58768=>"00000010",
  58769=>"00000011",
  58770=>"00000011",
  58771=>"11111100",
  58772=>"11111111",
  58773=>"00000000",
  58774=>"00000010",
  58775=>"11111111",
  58776=>"11111111",
  58777=>"11111100",
  58778=>"00000011",
  58779=>"00000001",
  58780=>"11111111",
  58781=>"11111111",
  58782=>"00000100",
  58783=>"00000100",
  58784=>"00000000",
  58785=>"00000001",
  58786=>"00000000",
  58787=>"00000001",
  58788=>"11111101",
  58789=>"00000000",
  58790=>"00000001",
  58791=>"11111111",
  58792=>"11111101",
  58793=>"00000111",
  58794=>"11111101",
  58795=>"11111110",
  58796=>"00000010",
  58797=>"00000010",
  58798=>"00000010",
  58799=>"00000010",
  58800=>"00000011",
  58801=>"00000000",
  58802=>"00000001",
  58803=>"11111101",
  58804=>"11111110",
  58805=>"00000011",
  58806=>"00000000",
  58807=>"00000011",
  58808=>"00000100",
  58809=>"00000000",
  58810=>"11111110",
  58811=>"11111110",
  58812=>"11111110",
  58813=>"11111100",
  58814=>"11111110",
  58815=>"00000000",
  58816=>"00000011",
  58817=>"00000000",
  58818=>"00000010",
  58819=>"00000011",
  58820=>"11111100",
  58821=>"11111101",
  58822=>"00000001",
  58823=>"11111110",
  58824=>"00000101",
  58825=>"00000010",
  58826=>"00000100",
  58827=>"00000011",
  58828=>"00000000",
  58829=>"00000000",
  58830=>"00000000",
  58831=>"11111110",
  58832=>"11111110",
  58833=>"11111111",
  58834=>"11111111",
  58835=>"11111111",
  58836=>"00000010",
  58837=>"11111100",
  58838=>"11111110",
  58839=>"00000010",
  58840=>"00000001",
  58841=>"11111111",
  58842=>"11111101",
  58843=>"00000010",
  58844=>"11111111",
  58845=>"11111111",
  58846=>"11111111",
  58847=>"11111111",
  58848=>"00000010",
  58849=>"00000101",
  58850=>"00000000",
  58851=>"00000011",
  58852=>"11111110",
  58853=>"00000001",
  58854=>"11111110",
  58855=>"11111101",
  58856=>"11111100",
  58857=>"11111111",
  58858=>"00000000",
  58859=>"00000101",
  58860=>"00000010",
  58861=>"11111111",
  58862=>"11111110",
  58863=>"11111010",
  58864=>"00000001",
  58865=>"00000000",
  58866=>"00000000",
  58867=>"00000000",
  58868=>"00000010",
  58869=>"00000000",
  58870=>"11111110",
  58871=>"11111111",
  58872=>"00000101",
  58873=>"00000011",
  58874=>"11111110",
  58875=>"00000000",
  58876=>"00000101",
  58877=>"00000001",
  58878=>"00000010",
  58879=>"00000100",
  58880=>"11111111",
  58881=>"11111111",
  58882=>"11111111",
  58883=>"11111111",
  58884=>"00000011",
  58885=>"00000010",
  58886=>"11111111",
  58887=>"11111111",
  58888=>"11111110",
  58889=>"11111111",
  58890=>"11111111",
  58891=>"00000010",
  58892=>"00000001",
  58893=>"00000000",
  58894=>"11111011",
  58895=>"00000001",
  58896=>"11111111",
  58897=>"00000000",
  58898=>"11111100",
  58899=>"11111101",
  58900=>"11111101",
  58901=>"00000000",
  58902=>"00000001",
  58903=>"11111101",
  58904=>"11111111",
  58905=>"00000101",
  58906=>"00000001",
  58907=>"00000011",
  58908=>"11111110",
  58909=>"11111111",
  58910=>"00000001",
  58911=>"00000001",
  58912=>"00000000",
  58913=>"00000000",
  58914=>"11111101",
  58915=>"00000000",
  58916=>"11111110",
  58917=>"11111111",
  58918=>"00000011",
  58919=>"11111111",
  58920=>"00000000",
  58921=>"11111110",
  58922=>"11111110",
  58923=>"11111110",
  58924=>"00000010",
  58925=>"11111111",
  58926=>"00000001",
  58927=>"11111100",
  58928=>"11111011",
  58929=>"00000011",
  58930=>"11111111",
  58931=>"11111101",
  58932=>"00000000",
  58933=>"00000100",
  58934=>"11111111",
  58935=>"00000001",
  58936=>"00000001",
  58937=>"00000010",
  58938=>"00000011",
  58939=>"00000000",
  58940=>"11111111",
  58941=>"11111111",
  58942=>"11111111",
  58943=>"11111101",
  58944=>"00000011",
  58945=>"11111111",
  58946=>"00000100",
  58947=>"11111100",
  58948=>"00000001",
  58949=>"00000000",
  58950=>"11111110",
  58951=>"00000011",
  58952=>"00000000",
  58953=>"00000010",
  58954=>"00000010",
  58955=>"11111111",
  58956=>"11111101",
  58957=>"00000001",
  58958=>"00000000",
  58959=>"11111111",
  58960=>"00000010",
  58961=>"00000010",
  58962=>"00000000",
  58963=>"11111111",
  58964=>"00000000",
  58965=>"00000001",
  58966=>"11111110",
  58967=>"11111101",
  58968=>"00000000",
  58969=>"00000010",
  58970=>"00000010",
  58971=>"11111101",
  58972=>"11111110",
  58973=>"11111111",
  58974=>"11111101",
  58975=>"11111110",
  58976=>"00000000",
  58977=>"00000010",
  58978=>"11111110",
  58979=>"11111110",
  58980=>"11111101",
  58981=>"00000010",
  58982=>"00000010",
  58983=>"00000100",
  58984=>"11111111",
  58985=>"00000101",
  58986=>"11111110",
  58987=>"00000011",
  58988=>"00000001",
  58989=>"00000001",
  58990=>"11111101",
  58991=>"11111111",
  58992=>"00000001",
  58993=>"00000100",
  58994=>"11111101",
  58995=>"11111101",
  58996=>"00000001",
  58997=>"11111111",
  58998=>"11111110",
  58999=>"11111110",
  59000=>"00000000",
  59001=>"11111101",
  59002=>"00000000",
  59003=>"00000000",
  59004=>"00000000",
  59005=>"00000001",
  59006=>"00000001",
  59007=>"00000011",
  59008=>"00000000",
  59009=>"11111101",
  59010=>"11111101",
  59011=>"11111111",
  59012=>"00000010",
  59013=>"00000001",
  59014=>"00000000",
  59015=>"00000000",
  59016=>"11111101",
  59017=>"00000011",
  59018=>"11111111",
  59019=>"00000010",
  59020=>"00000000",
  59021=>"00000001",
  59022=>"00000011",
  59023=>"00000110",
  59024=>"11111111",
  59025=>"11111110",
  59026=>"00000101",
  59027=>"11111110",
  59028=>"00000100",
  59029=>"11111101",
  59030=>"00000000",
  59031=>"00000010",
  59032=>"11111101",
  59033=>"00000000",
  59034=>"00000100",
  59035=>"00000000",
  59036=>"11111100",
  59037=>"11111111",
  59038=>"00000010",
  59039=>"00000000",
  59040=>"00000000",
  59041=>"00000011",
  59042=>"11111111",
  59043=>"11111110",
  59044=>"11111101",
  59045=>"11111101",
  59046=>"00000010",
  59047=>"11111100",
  59048=>"00000010",
  59049=>"11111101",
  59050=>"00000100",
  59051=>"11111110",
  59052=>"11111110",
  59053=>"00000001",
  59054=>"11111110",
  59055=>"00000001",
  59056=>"00000010",
  59057=>"11111101",
  59058=>"00000010",
  59059=>"11111111",
  59060=>"11111110",
  59061=>"11111110",
  59062=>"11111111",
  59063=>"11111110",
  59064=>"00000000",
  59065=>"00000101",
  59066=>"00000100",
  59067=>"00000001",
  59068=>"11111111",
  59069=>"11111111",
  59070=>"00000000",
  59071=>"00000010",
  59072=>"11111111",
  59073=>"11111101",
  59074=>"11111110",
  59075=>"11111110",
  59076=>"11111111",
  59077=>"11111101",
  59078=>"11111111",
  59079=>"11111111",
  59080=>"00000011",
  59081=>"11111111",
  59082=>"00000010",
  59083=>"00000000",
  59084=>"00000010",
  59085=>"00000110",
  59086=>"11111111",
  59087=>"11111111",
  59088=>"11111110",
  59089=>"00000010",
  59090=>"00000001",
  59091=>"11111101",
  59092=>"11111110",
  59093=>"11111110",
  59094=>"00000001",
  59095=>"00000001",
  59096=>"00000001",
  59097=>"00000011",
  59098=>"00000010",
  59099=>"11111111",
  59100=>"11111110",
  59101=>"11111111",
  59102=>"00000000",
  59103=>"00000000",
  59104=>"11111110",
  59105=>"00000001",
  59106=>"00000101",
  59107=>"00000010",
  59108=>"11111101",
  59109=>"11111111",
  59110=>"00000001",
  59111=>"00000010",
  59112=>"00000001",
  59113=>"00000000",
  59114=>"00000010",
  59115=>"11111111",
  59116=>"00000000",
  59117=>"00000001",
  59118=>"00000001",
  59119=>"11111111",
  59120=>"00000001",
  59121=>"11111111",
  59122=>"00000010",
  59123=>"11111110",
  59124=>"11111101",
  59125=>"00000010",
  59126=>"00000100",
  59127=>"11111111",
  59128=>"00000000",
  59129=>"00000011",
  59130=>"00000001",
  59131=>"00000000",
  59132=>"11111101",
  59133=>"11111110",
  59134=>"11111101",
  59135=>"11111111",
  59136=>"00000010",
  59137=>"11111110",
  59138=>"11111110",
  59139=>"00000011",
  59140=>"11111111",
  59141=>"11111101",
  59142=>"00000001",
  59143=>"11111110",
  59144=>"00000010",
  59145=>"11111110",
  59146=>"00000000",
  59147=>"11111101",
  59148=>"00000000",
  59149=>"11111110",
  59150=>"11111111",
  59151=>"00000100",
  59152=>"11111111",
  59153=>"00000001",
  59154=>"00000011",
  59155=>"00000001",
  59156=>"11111100",
  59157=>"00000100",
  59158=>"11111110",
  59159=>"11111110",
  59160=>"00000001",
  59161=>"11111100",
  59162=>"11111100",
  59163=>"11111111",
  59164=>"11111110",
  59165=>"11111110",
  59166=>"11111101",
  59167=>"00000011",
  59168=>"11111110",
  59169=>"11111110",
  59170=>"00000010",
  59171=>"00000010",
  59172=>"11111111",
  59173=>"00000010",
  59174=>"11111110",
  59175=>"00000001",
  59176=>"11111101",
  59177=>"00000001",
  59178=>"00000111",
  59179=>"11111111",
  59180=>"00000011",
  59181=>"00000010",
  59182=>"11111111",
  59183=>"11111110",
  59184=>"00000011",
  59185=>"11111110",
  59186=>"11111111",
  59187=>"00000000",
  59188=>"11111110",
  59189=>"00000000",
  59190=>"11111111",
  59191=>"00000011",
  59192=>"00000010",
  59193=>"00000000",
  59194=>"11111111",
  59195=>"00000110",
  59196=>"00000001",
  59197=>"00000010",
  59198=>"00000011",
  59199=>"11111100",
  59200=>"11111100",
  59201=>"00000010",
  59202=>"00000010",
  59203=>"11111111",
  59204=>"11111111",
  59205=>"11111110",
  59206=>"11111101",
  59207=>"11111111",
  59208=>"00000010",
  59209=>"11111111",
  59210=>"00000010",
  59211=>"00000001",
  59212=>"00000001",
  59213=>"11111111",
  59214=>"11111101",
  59215=>"00000000",
  59216=>"00000000",
  59217=>"00000000",
  59218=>"00000000",
  59219=>"00000001",
  59220=>"11111100",
  59221=>"00000011",
  59222=>"00000000",
  59223=>"00000000",
  59224=>"00000000",
  59225=>"11111101",
  59226=>"00000001",
  59227=>"00000101",
  59228=>"00000001",
  59229=>"11111110",
  59230=>"11111100",
  59231=>"00000001",
  59232=>"11111101",
  59233=>"00000101",
  59234=>"11111101",
  59235=>"00000000",
  59236=>"11111110",
  59237=>"11111111",
  59238=>"11111101",
  59239=>"00000010",
  59240=>"00000010",
  59241=>"00000011",
  59242=>"00000000",
  59243=>"00000001",
  59244=>"11111111",
  59245=>"11111110",
  59246=>"11111110",
  59247=>"00000000",
  59248=>"11111011",
  59249=>"00000001",
  59250=>"00000000",
  59251=>"11111100",
  59252=>"00000001",
  59253=>"11111100",
  59254=>"00000011",
  59255=>"11111101",
  59256=>"11111101",
  59257=>"00000100",
  59258=>"11111110",
  59259=>"00000010",
  59260=>"00000110",
  59261=>"11111110",
  59262=>"00000011",
  59263=>"00000001",
  59264=>"11111110",
  59265=>"11111101",
  59266=>"00000001",
  59267=>"11111111",
  59268=>"11111110",
  59269=>"00000001",
  59270=>"11111101",
  59271=>"00000001",
  59272=>"11111111",
  59273=>"00000001",
  59274=>"11111111",
  59275=>"00000010",
  59276=>"00000010",
  59277=>"11111111",
  59278=>"00000010",
  59279=>"11111111",
  59280=>"00000001",
  59281=>"11111101",
  59282=>"00000000",
  59283=>"11111111",
  59284=>"11111101",
  59285=>"00000000",
  59286=>"11111111",
  59287=>"11111110",
  59288=>"11111100",
  59289=>"00000000",
  59290=>"11111101",
  59291=>"00000111",
  59292=>"00000011",
  59293=>"00000001",
  59294=>"00000010",
  59295=>"00000001",
  59296=>"11111110",
  59297=>"11111111",
  59298=>"00000100",
  59299=>"00000001",
  59300=>"00000010",
  59301=>"11111101",
  59302=>"00000100",
  59303=>"11111110",
  59304=>"00000001",
  59305=>"00000001",
  59306=>"11111100",
  59307=>"11111101",
  59308=>"11111111",
  59309=>"00000000",
  59310=>"00000000",
  59311=>"11111101",
  59312=>"00000001",
  59313=>"11111101",
  59314=>"00000000",
  59315=>"00000001",
  59316=>"00000001",
  59317=>"11111111",
  59318=>"00000011",
  59319=>"00000001",
  59320=>"11111110",
  59321=>"11111110",
  59322=>"00000000",
  59323=>"00000010",
  59324=>"00000001",
  59325=>"11111111",
  59326=>"00000000",
  59327=>"11111110",
  59328=>"00000100",
  59329=>"00000000",
  59330=>"00000010",
  59331=>"00000001",
  59332=>"00000001",
  59333=>"11111110",
  59334=>"11111101",
  59335=>"11111111",
  59336=>"11111101",
  59337=>"11111101",
  59338=>"00000000",
  59339=>"00000001",
  59340=>"00000000",
  59341=>"11111101",
  59342=>"00000010",
  59343=>"11111110",
  59344=>"11111101",
  59345=>"11111101",
  59346=>"00000001",
  59347=>"00000001",
  59348=>"00000010",
  59349=>"00000011",
  59350=>"11111110",
  59351=>"11111101",
  59352=>"11111110",
  59353=>"00000011",
  59354=>"00000011",
  59355=>"00000001",
  59356=>"11111110",
  59357=>"11111111",
  59358=>"11111101",
  59359=>"11111101",
  59360=>"00000010",
  59361=>"00000001",
  59362=>"00000011",
  59363=>"00000001",
  59364=>"11111101",
  59365=>"00000010",
  59366=>"00000110",
  59367=>"00000000",
  59368=>"00000011",
  59369=>"11111111",
  59370=>"11111101",
  59371=>"11111111",
  59372=>"11111111",
  59373=>"00000011",
  59374=>"00000110",
  59375=>"00000001",
  59376=>"11111101",
  59377=>"00000011",
  59378=>"11111101",
  59379=>"00000010",
  59380=>"00000010",
  59381=>"11111111",
  59382=>"11111100",
  59383=>"00000010",
  59384=>"11111110",
  59385=>"00000010",
  59386=>"00000101",
  59387=>"00000001",
  59388=>"00000001",
  59389=>"00000110",
  59390=>"00000000",
  59391=>"11111110",
  59392=>"11111111",
  59393=>"00000001",
  59394=>"00000001",
  59395=>"00000010",
  59396=>"00000100",
  59397=>"00000000",
  59398=>"00000010",
  59399=>"00000000",
  59400=>"11111111",
  59401=>"11111110",
  59402=>"11111110",
  59403=>"00000000",
  59404=>"00000010",
  59405=>"11111101",
  59406=>"11111101",
  59407=>"11111100",
  59408=>"00000010",
  59409=>"11111110",
  59410=>"11111101",
  59411=>"00000000",
  59412=>"00000011",
  59413=>"11111111",
  59414=>"11111111",
  59415=>"00000010",
  59416=>"00000011",
  59417=>"11111110",
  59418=>"00000001",
  59419=>"11111110",
  59420=>"00000001",
  59421=>"11111110",
  59422=>"11111111",
  59423=>"00000000",
  59424=>"00000011",
  59425=>"11111111",
  59426=>"11111101",
  59427=>"11111111",
  59428=>"11111110",
  59429=>"11111101",
  59430=>"00000011",
  59431=>"00000000",
  59432=>"11111110",
  59433=>"11111100",
  59434=>"11111100",
  59435=>"11111101",
  59436=>"11111100",
  59437=>"11111101",
  59438=>"11111110",
  59439=>"00000010",
  59440=>"11111111",
  59441=>"11111110",
  59442=>"00000010",
  59443=>"00000011",
  59444=>"11111110",
  59445=>"00000100",
  59446=>"00000001",
  59447=>"11111110",
  59448=>"11111110",
  59449=>"11111101",
  59450=>"00000000",
  59451=>"11111101",
  59452=>"11111111",
  59453=>"11111110",
  59454=>"00000011",
  59455=>"11111111",
  59456=>"00000011",
  59457=>"11111111",
  59458=>"00000000",
  59459=>"00000001",
  59460=>"00000000",
  59461=>"11111111",
  59462=>"11111110",
  59463=>"11111111",
  59464=>"11111111",
  59465=>"11111111",
  59466=>"00000000",
  59467=>"00000000",
  59468=>"11111111",
  59469=>"00000101",
  59470=>"00000010",
  59471=>"00000001",
  59472=>"00000100",
  59473=>"00000010",
  59474=>"00000000",
  59475=>"11111100",
  59476=>"00000010",
  59477=>"11111110",
  59478=>"11111110",
  59479=>"11111101",
  59480=>"00000000",
  59481=>"00000010",
  59482=>"11111101",
  59483=>"11111101",
  59484=>"00000010",
  59485=>"00000010",
  59486=>"11111110",
  59487=>"00000000",
  59488=>"11111101",
  59489=>"00000010",
  59490=>"00000000",
  59491=>"00000010",
  59492=>"00000010",
  59493=>"00000010",
  59494=>"11111101",
  59495=>"00000010",
  59496=>"11111101",
  59497=>"00000101",
  59498=>"11111111",
  59499=>"11111111",
  59500=>"11111111",
  59501=>"00000001",
  59502=>"11111101",
  59503=>"00000000",
  59504=>"00000011",
  59505=>"00000011",
  59506=>"00000000",
  59507=>"00000011",
  59508=>"00000011",
  59509=>"11111101",
  59510=>"00000001",
  59511=>"00000000",
  59512=>"00000010",
  59513=>"11111100",
  59514=>"00000001",
  59515=>"00000100",
  59516=>"00000010",
  59517=>"00000100",
  59518=>"00000000",
  59519=>"00000000",
  59520=>"00000000",
  59521=>"00000101",
  59522=>"11111110",
  59523=>"11111101",
  59524=>"00000010",
  59525=>"11111111",
  59526=>"00000001",
  59527=>"00000010",
  59528=>"11111111",
  59529=>"11111110",
  59530=>"11111110",
  59531=>"00000110",
  59532=>"11111110",
  59533=>"11111110",
  59534=>"00000001",
  59535=>"00000001",
  59536=>"00000001",
  59537=>"00000000",
  59538=>"00000010",
  59539=>"00000011",
  59540=>"11111110",
  59541=>"00000000",
  59542=>"00000000",
  59543=>"11111110",
  59544=>"11111111",
  59545=>"00000001",
  59546=>"11111110",
  59547=>"11111101",
  59548=>"00000001",
  59549=>"00000010",
  59550=>"00000001",
  59551=>"11111110",
  59552=>"00000010",
  59553=>"11111111",
  59554=>"11111101",
  59555=>"11111111",
  59556=>"00000001",
  59557=>"11111110",
  59558=>"11111101",
  59559=>"11111101",
  59560=>"00000000",
  59561=>"11111110",
  59562=>"11111101",
  59563=>"00000001",
  59564=>"11111111",
  59565=>"00000010",
  59566=>"00000001",
  59567=>"11111101",
  59568=>"00000010",
  59569=>"11111111",
  59570=>"00000010",
  59571=>"00000001",
  59572=>"11111110",
  59573=>"11111101",
  59574=>"00000001",
  59575=>"00000001",
  59576=>"00000010",
  59577=>"00000011",
  59578=>"11111101",
  59579=>"11111111",
  59580=>"11111111",
  59581=>"00000010",
  59582=>"00000010",
  59583=>"11111111",
  59584=>"11111101",
  59585=>"11111110",
  59586=>"00000000",
  59587=>"00000011",
  59588=>"11111111",
  59589=>"00000001",
  59590=>"00000000",
  59591=>"00000011",
  59592=>"00000001",
  59593=>"00000001",
  59594=>"00000001",
  59595=>"11111101",
  59596=>"11111111",
  59597=>"11111110",
  59598=>"11111110",
  59599=>"11111101",
  59600=>"00000000",
  59601=>"11111101",
  59602=>"00000000",
  59603=>"00000001",
  59604=>"11111110",
  59605=>"11111101",
  59606=>"11111110",
  59607=>"11111101",
  59608=>"11111110",
  59609=>"00000001",
  59610=>"00000000",
  59611=>"00000001",
  59612=>"11111111",
  59613=>"00000000",
  59614=>"00000001",
  59615=>"00000000",
  59616=>"00000000",
  59617=>"00000001",
  59618=>"00000001",
  59619=>"11111110",
  59620=>"11111111",
  59621=>"11111110",
  59622=>"11111100",
  59623=>"11111101",
  59624=>"11111110",
  59625=>"00000001",
  59626=>"11111110",
  59627=>"00000000",
  59628=>"00000011",
  59629=>"11111110",
  59630=>"00000001",
  59631=>"00000000",
  59632=>"11111111",
  59633=>"11111111",
  59634=>"11111110",
  59635=>"00000001",
  59636=>"00000000",
  59637=>"00000001",
  59638=>"11111111",
  59639=>"11111111",
  59640=>"11111101",
  59641=>"11111101",
  59642=>"00000000",
  59643=>"00000000",
  59644=>"00000010",
  59645=>"11111110",
  59646=>"11111111",
  59647=>"00000001",
  59648=>"00000001",
  59649=>"00000001",
  59650=>"00000000",
  59651=>"00000011",
  59652=>"00000011",
  59653=>"11111101",
  59654=>"00000010",
  59655=>"11111101",
  59656=>"00000011",
  59657=>"11111101",
  59658=>"00000000",
  59659=>"00000001",
  59660=>"11111111",
  59661=>"11111111",
  59662=>"11111111",
  59663=>"00000000",
  59664=>"00000000",
  59665=>"00000000",
  59666=>"11111110",
  59667=>"11111110",
  59668=>"11111110",
  59669=>"00000000",
  59670=>"00000001",
  59671=>"00000010",
  59672=>"00000101",
  59673=>"00000010",
  59674=>"11111101",
  59675=>"00000001",
  59676=>"00000011",
  59677=>"11111111",
  59678=>"11111111",
  59679=>"00000000",
  59680=>"11111101",
  59681=>"11111110",
  59682=>"00000010",
  59683=>"00000101",
  59684=>"11111110",
  59685=>"00000000",
  59686=>"11111101",
  59687=>"11111110",
  59688=>"00000010",
  59689=>"00000010",
  59690=>"00000010",
  59691=>"11111111",
  59692=>"00000010",
  59693=>"11111101",
  59694=>"00000010",
  59695=>"11111111",
  59696=>"00000000",
  59697=>"00000010",
  59698=>"00000011",
  59699=>"00000010",
  59700=>"00000001",
  59701=>"11111111",
  59702=>"11111110",
  59703=>"11111111",
  59704=>"11111101",
  59705=>"11111110",
  59706=>"11111111",
  59707=>"11111100",
  59708=>"00000000",
  59709=>"00000001",
  59710=>"00000010",
  59711=>"00000000",
  59712=>"00000010",
  59713=>"11111111",
  59714=>"11111111",
  59715=>"11111111",
  59716=>"00000010",
  59717=>"00000001",
  59718=>"00000000",
  59719=>"00000000",
  59720=>"11111101",
  59721=>"11111111",
  59722=>"00000011",
  59723=>"11111110",
  59724=>"00000001",
  59725=>"00000000",
  59726=>"00000000",
  59727=>"11111101",
  59728=>"11111110",
  59729=>"11111111",
  59730=>"11111110",
  59731=>"00000001",
  59732=>"11111111",
  59733=>"11111110",
  59734=>"11111111",
  59735=>"00000000",
  59736=>"00000001",
  59737=>"00000001",
  59738=>"00000000",
  59739=>"11111101",
  59740=>"11111110",
  59741=>"00000001",
  59742=>"00000000",
  59743=>"11111110",
  59744=>"00000001",
  59745=>"11111101",
  59746=>"00000001",
  59747=>"00000100",
  59748=>"00000010",
  59749=>"00000010",
  59750=>"11111110",
  59751=>"00000010",
  59752=>"00000000",
  59753=>"00000011",
  59754=>"11111101",
  59755=>"00000010",
  59756=>"11111110",
  59757=>"00000100",
  59758=>"11111110",
  59759=>"00000000",
  59760=>"00000011",
  59761=>"11111110",
  59762=>"00000000",
  59763=>"11111110",
  59764=>"00000000",
  59765=>"00000000",
  59766=>"11111101",
  59767=>"11111110",
  59768=>"00000000",
  59769=>"00000010",
  59770=>"11111110",
  59771=>"00000000",
  59772=>"11111101",
  59773=>"00000000",
  59774=>"00000010",
  59775=>"00000101",
  59776=>"11111101",
  59777=>"11111110",
  59778=>"11111111",
  59779=>"00000011",
  59780=>"00000000",
  59781=>"00000001",
  59782=>"00000100",
  59783=>"00000010",
  59784=>"00000001",
  59785=>"00000101",
  59786=>"00000011",
  59787=>"00000101",
  59788=>"00000000",
  59789=>"00000011",
  59790=>"00000001",
  59791=>"11111111",
  59792=>"11111111",
  59793=>"00000011",
  59794=>"00000100",
  59795=>"00000100",
  59796=>"00000001",
  59797=>"00000011",
  59798=>"11111101",
  59799=>"11111110",
  59800=>"11111111",
  59801=>"11111110",
  59802=>"00000001",
  59803=>"00000010",
  59804=>"11111101",
  59805=>"00000000",
  59806=>"11111111",
  59807=>"11111110",
  59808=>"11111101",
  59809=>"11111100",
  59810=>"11111101",
  59811=>"00000000",
  59812=>"00000001",
  59813=>"00000010",
  59814=>"11111111",
  59815=>"11111111",
  59816=>"00000001",
  59817=>"11111101",
  59818=>"11111111",
  59819=>"00000000",
  59820=>"00000000",
  59821=>"00000110",
  59822=>"11111101",
  59823=>"11111111",
  59824=>"00000010",
  59825=>"00000111",
  59826=>"11111111",
  59827=>"00000000",
  59828=>"00000010",
  59829=>"00000010",
  59830=>"00000001",
  59831=>"00000000",
  59832=>"00000010",
  59833=>"00000000",
  59834=>"11111110",
  59835=>"00000001",
  59836=>"11111111",
  59837=>"00000000",
  59838=>"00000101",
  59839=>"00000000",
  59840=>"00000011",
  59841=>"11111101",
  59842=>"11111110",
  59843=>"00000001",
  59844=>"00000010",
  59845=>"00000000",
  59846=>"00000100",
  59847=>"00000011",
  59848=>"11111111",
  59849=>"00000000",
  59850=>"11111111",
  59851=>"00000011",
  59852=>"11111111",
  59853=>"11111111",
  59854=>"00000010",
  59855=>"00000000",
  59856=>"11111111",
  59857=>"00000011",
  59858=>"00000010",
  59859=>"11111110",
  59860=>"11111110",
  59861=>"00000000",
  59862=>"00000011",
  59863=>"00000100",
  59864=>"11111111",
  59865=>"00000011",
  59866=>"00000001",
  59867=>"11111111",
  59868=>"00000000",
  59869=>"00000010",
  59870=>"11111110",
  59871=>"11111110",
  59872=>"00000000",
  59873=>"11111110",
  59874=>"00000010",
  59875=>"00000001",
  59876=>"00000010",
  59877=>"00000001",
  59878=>"00000000",
  59879=>"00000000",
  59880=>"11111110",
  59881=>"00000010",
  59882=>"11111110",
  59883=>"00000100",
  59884=>"11111111",
  59885=>"00000100",
  59886=>"00000011",
  59887=>"00000001",
  59888=>"00000000",
  59889=>"00000101",
  59890=>"11111101",
  59891=>"00000010",
  59892=>"00000001",
  59893=>"00000010",
  59894=>"11111111",
  59895=>"00000101",
  59896=>"00000010",
  59897=>"11111110",
  59898=>"00000000",
  59899=>"00000000",
  59900=>"00000011",
  59901=>"00000001",
  59902=>"00000010",
  59903=>"00000000",
  59904=>"00000010",
  59905=>"00000000",
  59906=>"11111110",
  59907=>"00000011",
  59908=>"00000010",
  59909=>"00000101",
  59910=>"11111101",
  59911=>"00000000",
  59912=>"00000011",
  59913=>"00000010",
  59914=>"00000011",
  59915=>"11111111",
  59916=>"11111111",
  59917=>"00000010",
  59918=>"00000011",
  59919=>"11111101",
  59920=>"00000010",
  59921=>"11111110",
  59922=>"00000000",
  59923=>"11111110",
  59924=>"00000011",
  59925=>"00000000",
  59926=>"11111101",
  59927=>"00000001",
  59928=>"00000000",
  59929=>"00000010",
  59930=>"11111110",
  59931=>"00000000",
  59932=>"00000000",
  59933=>"11111101",
  59934=>"11111111",
  59935=>"11111110",
  59936=>"11111111",
  59937=>"00000001",
  59938=>"11111110",
  59939=>"00000110",
  59940=>"00000000",
  59941=>"00000000",
  59942=>"11111101",
  59943=>"11111110",
  59944=>"11111111",
  59945=>"11111110",
  59946=>"00000000",
  59947=>"00000001",
  59948=>"00000001",
  59949=>"00000000",
  59950=>"00000011",
  59951=>"00000000",
  59952=>"00000000",
  59953=>"00000010",
  59954=>"00000011",
  59955=>"00000000",
  59956=>"00000100",
  59957=>"11111110",
  59958=>"11111111",
  59959=>"00000000",
  59960=>"00000011",
  59961=>"00000000",
  59962=>"11111110",
  59963=>"00000000",
  59964=>"11111111",
  59965=>"11111111",
  59966=>"00000100",
  59967=>"11111101",
  59968=>"11111110",
  59969=>"11111111",
  59970=>"00000011",
  59971=>"00000000",
  59972=>"00000000",
  59973=>"00000100",
  59974=>"11111100",
  59975=>"00000011",
  59976=>"00000011",
  59977=>"00000001",
  59978=>"00000000",
  59979=>"00000011",
  59980=>"11111110",
  59981=>"00000000",
  59982=>"11111111",
  59983=>"00000001",
  59984=>"11111110",
  59985=>"11111111",
  59986=>"11111110",
  59987=>"00000010",
  59988=>"00000000",
  59989=>"00000000",
  59990=>"00000000",
  59991=>"00000010",
  59992=>"00000011",
  59993=>"00000001",
  59994=>"00000010",
  59995=>"00000000",
  59996=>"00000000",
  59997=>"00000010",
  59998=>"11111111",
  59999=>"00000000",
  60000=>"00000010",
  60001=>"11111110",
  60002=>"11111111",
  60003=>"11111111",
  60004=>"11111101",
  60005=>"11111110",
  60006=>"11111111",
  60007=>"11111100",
  60008=>"11111110",
  60009=>"00000010",
  60010=>"00000010",
  60011=>"11111111",
  60012=>"00000000",
  60013=>"11111111",
  60014=>"11111100",
  60015=>"00000001",
  60016=>"00000100",
  60017=>"11111110",
  60018=>"00000000",
  60019=>"11111111",
  60020=>"00000001",
  60021=>"11111110",
  60022=>"11111101",
  60023=>"00000001",
  60024=>"00000011",
  60025=>"11111110",
  60026=>"00000000",
  60027=>"11111111",
  60028=>"00000010",
  60029=>"00000000",
  60030=>"00000001",
  60031=>"00000010",
  60032=>"00000001",
  60033=>"11111110",
  60034=>"11111100",
  60035=>"00000010",
  60036=>"00000001",
  60037=>"11111111",
  60038=>"00000100",
  60039=>"00000010",
  60040=>"11111111",
  60041=>"00000001",
  60042=>"00000011",
  60043=>"00000001",
  60044=>"11111111",
  60045=>"00000011",
  60046=>"11111110",
  60047=>"11111110",
  60048=>"11111111",
  60049=>"00000001",
  60050=>"00000001",
  60051=>"11111101",
  60052=>"00000011",
  60053=>"00000010",
  60054=>"00000000",
  60055=>"00000011",
  60056=>"11111101",
  60057=>"00000001",
  60058=>"11111110",
  60059=>"00000011",
  60060=>"11111111",
  60061=>"11111101",
  60062=>"00000001",
  60063=>"11111101",
  60064=>"11111111",
  60065=>"00000000",
  60066=>"00000100",
  60067=>"00000010",
  60068=>"11111101",
  60069=>"00000101",
  60070=>"00000011",
  60071=>"11111111",
  60072=>"00000011",
  60073=>"00000001",
  60074=>"11111101",
  60075=>"00000000",
  60076=>"00000001",
  60077=>"00000000",
  60078=>"11111110",
  60079=>"00000010",
  60080=>"11111110",
  60081=>"00000001",
  60082=>"00000001",
  60083=>"11111111",
  60084=>"00000011",
  60085=>"00000100",
  60086=>"11111110",
  60087=>"00000001",
  60088=>"11111111",
  60089=>"00000000",
  60090=>"00000001",
  60091=>"00000100",
  60092=>"00000000",
  60093=>"11111110",
  60094=>"00000001",
  60095=>"00000010",
  60096=>"00000011",
  60097=>"00000000",
  60098=>"00000001",
  60099=>"00000010",
  60100=>"00000000",
  60101=>"00000000",
  60102=>"11111111",
  60103=>"11111101",
  60104=>"11111110",
  60105=>"11111111",
  60106=>"00000101",
  60107=>"00000010",
  60108=>"11111111",
  60109=>"00000011",
  60110=>"00000000",
  60111=>"00000000",
  60112=>"00000010",
  60113=>"11111111",
  60114=>"11111101",
  60115=>"00000000",
  60116=>"11111110",
  60117=>"11111110",
  60118=>"00000000",
  60119=>"11111110",
  60120=>"00000001",
  60121=>"11111110",
  60122=>"11111111",
  60123=>"11111110",
  60124=>"00000000",
  60125=>"11111110",
  60126=>"11111110",
  60127=>"00000000",
  60128=>"00000010",
  60129=>"11111101",
  60130=>"00000000",
  60131=>"11111111",
  60132=>"00000000",
  60133=>"00000001",
  60134=>"00000000",
  60135=>"00000000",
  60136=>"00000000",
  60137=>"00000000",
  60138=>"11111111",
  60139=>"00000001",
  60140=>"00000000",
  60141=>"11111101",
  60142=>"11111101",
  60143=>"11111111",
  60144=>"00000010",
  60145=>"11111111",
  60146=>"00000010",
  60147=>"00000000",
  60148=>"11111111",
  60149=>"11111110",
  60150=>"11111110",
  60151=>"11111110",
  60152=>"00000000",
  60153=>"11111111",
  60154=>"11111111",
  60155=>"11111101",
  60156=>"00000001",
  60157=>"00000010",
  60158=>"00000001",
  60159=>"11111111",
  60160=>"00000000",
  60161=>"11111101",
  60162=>"00000100",
  60163=>"00000000",
  60164=>"00000101",
  60165=>"11111111",
  60166=>"11111111",
  60167=>"11111110",
  60168=>"00000100",
  60169=>"00000000",
  60170=>"00000001",
  60171=>"11111111",
  60172=>"00000011",
  60173=>"00000110",
  60174=>"00000000",
  60175=>"11111110",
  60176=>"11111110",
  60177=>"00000010",
  60178=>"00000001",
  60179=>"00000000",
  60180=>"11111111",
  60181=>"00000001",
  60182=>"00000001",
  60183=>"00000001",
  60184=>"11111110",
  60185=>"11111111",
  60186=>"11111110",
  60187=>"00000001",
  60188=>"11111111",
  60189=>"00000011",
  60190=>"11111101",
  60191=>"00000011",
  60192=>"00000010",
  60193=>"11111110",
  60194=>"11111110",
  60195=>"00000000",
  60196=>"00000000",
  60197=>"00000001",
  60198=>"00000010",
  60199=>"00000000",
  60200=>"11111100",
  60201=>"00000010",
  60202=>"11111101",
  60203=>"00000001",
  60204=>"00000001",
  60205=>"00000011",
  60206=>"00000001",
  60207=>"00000010",
  60208=>"00000000",
  60209=>"00000010",
  60210=>"00000001",
  60211=>"00000010",
  60212=>"11111111",
  60213=>"00000000",
  60214=>"00000010",
  60215=>"00000010",
  60216=>"11111101",
  60217=>"00000011",
  60218=>"00000000",
  60219=>"11111101",
  60220=>"00000011",
  60221=>"00000000",
  60222=>"11111110",
  60223=>"11111111",
  60224=>"00000101",
  60225=>"11111111",
  60226=>"11111101",
  60227=>"11111101",
  60228=>"00000010",
  60229=>"00000011",
  60230=>"00000001",
  60231=>"00000011",
  60232=>"00000000",
  60233=>"00000011",
  60234=>"00000000",
  60235=>"11111111",
  60236=>"00000001",
  60237=>"11111111",
  60238=>"11111111",
  60239=>"11111111",
  60240=>"11111101",
  60241=>"00000001",
  60242=>"11111111",
  60243=>"00000000",
  60244=>"11111110",
  60245=>"11111110",
  60246=>"11111110",
  60247=>"11111110",
  60248=>"11111111",
  60249=>"00000001",
  60250=>"00000000",
  60251=>"00000010",
  60252=>"11111111",
  60253=>"00000000",
  60254=>"00000000",
  60255=>"00000011",
  60256=>"11111110",
  60257=>"11111111",
  60258=>"11111111",
  60259=>"11111101",
  60260=>"00000000",
  60261=>"11111101",
  60262=>"00000100",
  60263=>"11111101",
  60264=>"00000010",
  60265=>"11111111",
  60266=>"11111111",
  60267=>"00000000",
  60268=>"00000010",
  60269=>"00000000",
  60270=>"11111100",
  60271=>"00000001",
  60272=>"11111101",
  60273=>"00000000",
  60274=>"00000000",
  60275=>"11111110",
  60276=>"00000001",
  60277=>"00000010",
  60278=>"00000011",
  60279=>"00000011",
  60280=>"00000000",
  60281=>"11111110",
  60282=>"00000001",
  60283=>"00000001",
  60284=>"00000101",
  60285=>"11111110",
  60286=>"00000001",
  60287=>"11111110",
  60288=>"00000000",
  60289=>"00000010",
  60290=>"11111101",
  60291=>"11111101",
  60292=>"00000100",
  60293=>"11111110",
  60294=>"11111101",
  60295=>"00000010",
  60296=>"00000001",
  60297=>"00000100",
  60298=>"00000000",
  60299=>"00000000",
  60300=>"00000010",
  60301=>"00000000",
  60302=>"11111111",
  60303=>"00000010",
  60304=>"11111110",
  60305=>"00000101",
  60306=>"00000000",
  60307=>"00000010",
  60308=>"00000001",
  60309=>"11111110",
  60310=>"00000010",
  60311=>"11111110",
  60312=>"11111110",
  60313=>"00000100",
  60314=>"00000001",
  60315=>"11111110",
  60316=>"00000100",
  60317=>"00000010",
  60318=>"00000000",
  60319=>"11111110",
  60320=>"11111111",
  60321=>"00000001",
  60322=>"11111111",
  60323=>"00000000",
  60324=>"00000001",
  60325=>"00000010",
  60326=>"11111110",
  60327=>"11111111",
  60328=>"11111101",
  60329=>"00000100",
  60330=>"00000000",
  60331=>"00000001",
  60332=>"11111111",
  60333=>"11111110",
  60334=>"00000011",
  60335=>"00000001",
  60336=>"11111110",
  60337=>"11111111",
  60338=>"00000000",
  60339=>"00000011",
  60340=>"00000000",
  60341=>"11111111",
  60342=>"11111101",
  60343=>"00000001",
  60344=>"00000101",
  60345=>"00000010",
  60346=>"00000001",
  60347=>"00000011",
  60348=>"00000010",
  60349=>"11111110",
  60350=>"11111110",
  60351=>"11111110",
  60352=>"11111101",
  60353=>"00000001",
  60354=>"00000001",
  60355=>"00000001",
  60356=>"00000000",
  60357=>"00000011",
  60358=>"11111101",
  60359=>"11111111",
  60360=>"00000010",
  60361=>"00000001",
  60362=>"11111101",
  60363=>"11111111",
  60364=>"11111110",
  60365=>"11111101",
  60366=>"00000010",
  60367=>"11111101",
  60368=>"11111110",
  60369=>"00000010",
  60370=>"11111101",
  60371=>"00000000",
  60372=>"00000010",
  60373=>"11111100",
  60374=>"11111110",
  60375=>"00000001",
  60376=>"00000010",
  60377=>"11111110",
  60378=>"11111111",
  60379=>"00000001",
  60380=>"00000000",
  60381=>"00000010",
  60382=>"11111111",
  60383=>"11111111",
  60384=>"11111111",
  60385=>"11111110",
  60386=>"11111111",
  60387=>"00000001",
  60388=>"11111110",
  60389=>"11111111",
  60390=>"11111110",
  60391=>"00000110",
  60392=>"11111111",
  60393=>"11111111",
  60394=>"11111101",
  60395=>"00000000",
  60396=>"11111111",
  60397=>"11111101",
  60398=>"00000100",
  60399=>"00000001",
  60400=>"00000000",
  60401=>"00000000",
  60402=>"00000010",
  60403=>"00000000",
  60404=>"00000001",
  60405=>"00000000",
  60406=>"11111110",
  60407=>"11111111",
  60408=>"00000011",
  60409=>"00000010",
  60410=>"11111100",
  60411=>"11111111",
  60412=>"00000001",
  60413=>"00000001",
  60414=>"00000110",
  60415=>"11111110",
  60416=>"00000011",
  60417=>"11111111",
  60418=>"00000011",
  60419=>"11111100",
  60420=>"00000010",
  60421=>"11111101",
  60422=>"11111101",
  60423=>"11111110",
  60424=>"00000001",
  60425=>"11111110",
  60426=>"00000001",
  60427=>"00000001",
  60428=>"00000000",
  60429=>"11111101",
  60430=>"00000000",
  60431=>"11111110",
  60432=>"00000001",
  60433=>"00000011",
  60434=>"00000010",
  60435=>"00000000",
  60436=>"11111110",
  60437=>"00000011",
  60438=>"00000001",
  60439=>"11111110",
  60440=>"00000001",
  60441=>"11111100",
  60442=>"00000000",
  60443=>"00000011",
  60444=>"00000001",
  60445=>"00000000",
  60446=>"00000000",
  60447=>"00000010",
  60448=>"00000001",
  60449=>"11111111",
  60450=>"00000000",
  60451=>"11111111",
  60452=>"00000001",
  60453=>"00000011",
  60454=>"00000000",
  60455=>"11111100",
  60456=>"00000010",
  60457=>"11111101",
  60458=>"00000100",
  60459=>"00000001",
  60460=>"11111101",
  60461=>"00000000",
  60462=>"00000001",
  60463=>"11111101",
  60464=>"11111111",
  60465=>"11111111",
  60466=>"00000000",
  60467=>"00000100",
  60468=>"11111111",
  60469=>"00000001",
  60470=>"11111110",
  60471=>"11111101",
  60472=>"11111111",
  60473=>"00000000",
  60474=>"00000000",
  60475=>"11111110",
  60476=>"00000011",
  60477=>"11111110",
  60478=>"00000001",
  60479=>"00000000",
  60480=>"00000010",
  60481=>"11111111",
  60482=>"11111110",
  60483=>"11111111",
  60484=>"11111110",
  60485=>"00000011",
  60486=>"00000010",
  60487=>"11111110",
  60488=>"00000011",
  60489=>"11111111",
  60490=>"11111111",
  60491=>"11111110",
  60492=>"00000010",
  60493=>"11111111",
  60494=>"11111111",
  60495=>"11111111",
  60496=>"00000001",
  60497=>"00000011",
  60498=>"11111100",
  60499=>"00000011",
  60500=>"11111110",
  60501=>"11111110",
  60502=>"00000110",
  60503=>"00000000",
  60504=>"00000001",
  60505=>"00000010",
  60506=>"00000001",
  60507=>"00000101",
  60508=>"00000010",
  60509=>"00000000",
  60510=>"00000000",
  60511=>"00000000",
  60512=>"00000110",
  60513=>"00000001",
  60514=>"11111100",
  60515=>"11111101",
  60516=>"11111111",
  60517=>"00000001",
  60518=>"11111110",
  60519=>"00000000",
  60520=>"00000011",
  60521=>"00000001",
  60522=>"00000000",
  60523=>"00000010",
  60524=>"11111011",
  60525=>"11111101",
  60526=>"11111101",
  60527=>"00000001",
  60528=>"00000010",
  60529=>"11111111",
  60530=>"11111111",
  60531=>"11111100",
  60532=>"00000000",
  60533=>"11111110",
  60534=>"00000000",
  60535=>"11111101",
  60536=>"00000101",
  60537=>"00000001",
  60538=>"00000001",
  60539=>"00000010",
  60540=>"11111101",
  60541=>"11111110",
  60542=>"00000001",
  60543=>"11111100",
  60544=>"00000010",
  60545=>"00000000",
  60546=>"11111110",
  60547=>"11111110",
  60548=>"11111110",
  60549=>"00000000",
  60550=>"00000010",
  60551=>"11111101",
  60552=>"11111111",
  60553=>"00000001",
  60554=>"11111101",
  60555=>"11111111",
  60556=>"00000100",
  60557=>"11111110",
  60558=>"00000010",
  60559=>"00000001",
  60560=>"11111111",
  60561=>"11111110",
  60562=>"00000010",
  60563=>"00000001",
  60564=>"00000000",
  60565=>"00000001",
  60566=>"00000110",
  60567=>"00000011",
  60568=>"11111100",
  60569=>"00000000",
  60570=>"00000000",
  60571=>"11111101",
  60572=>"00000010",
  60573=>"11111101",
  60574=>"11111110",
  60575=>"00000010",
  60576=>"00000001",
  60577=>"11111110",
  60578=>"11111100",
  60579=>"00000101",
  60580=>"00000001",
  60581=>"00000001",
  60582=>"11111110",
  60583=>"00000011",
  60584=>"00000000",
  60585=>"11111110",
  60586=>"11111111",
  60587=>"11111101",
  60588=>"11111111",
  60589=>"11111110",
  60590=>"00000001",
  60591=>"00000010",
  60592=>"11111111",
  60593=>"00000000",
  60594=>"00000100",
  60595=>"11111110",
  60596=>"11111011",
  60597=>"11111111",
  60598=>"00000010",
  60599=>"11111101",
  60600=>"11111101",
  60601=>"00000001",
  60602=>"11111101",
  60603=>"00000101",
  60604=>"00000000",
  60605=>"11111111",
  60606=>"00000001",
  60607=>"11111110",
  60608=>"00000000",
  60609=>"00000001",
  60610=>"11111101",
  60611=>"11111111",
  60612=>"00000010",
  60613=>"11111111",
  60614=>"11111110",
  60615=>"00000010",
  60616=>"00000001",
  60617=>"00000001",
  60618=>"11111101",
  60619=>"11111101",
  60620=>"00000100",
  60621=>"00000001",
  60622=>"00000011",
  60623=>"11111111",
  60624=>"11111101",
  60625=>"00000000",
  60626=>"00000000",
  60627=>"00000000",
  60628=>"00000011",
  60629=>"00000000",
  60630=>"11111110",
  60631=>"11111101",
  60632=>"11111100",
  60633=>"00000001",
  60634=>"00000010",
  60635=>"00000001",
  60636=>"00000100",
  60637=>"00000000",
  60638=>"00000001",
  60639=>"00000011",
  60640=>"11111111",
  60641=>"11111110",
  60642=>"00000100",
  60643=>"00000011",
  60644=>"00000010",
  60645=>"11111101",
  60646=>"00000110",
  60647=>"00000001",
  60648=>"00000010",
  60649=>"00000011",
  60650=>"00000001",
  60651=>"00000000",
  60652=>"00000010",
  60653=>"00000011",
  60654=>"00000011",
  60655=>"11111110",
  60656=>"11111110",
  60657=>"11111111",
  60658=>"00000010",
  60659=>"11111101",
  60660=>"00000011",
  60661=>"11111101",
  60662=>"11111111",
  60663=>"00000011",
  60664=>"00000000",
  60665=>"11111101",
  60666=>"11111111",
  60667=>"00000001",
  60668=>"00000000",
  60669=>"11111111",
  60670=>"11111100",
  60671=>"11111110",
  60672=>"00000010",
  60673=>"00000001",
  60674=>"00000011",
  60675=>"00000000",
  60676=>"00000010",
  60677=>"00000101",
  60678=>"11111110",
  60679=>"00000000",
  60680=>"00000011",
  60681=>"00000100",
  60682=>"00000010",
  60683=>"00000010",
  60684=>"00000001",
  60685=>"00000011",
  60686=>"00000011",
  60687=>"00000000",
  60688=>"11111101",
  60689=>"11111111",
  60690=>"00000010",
  60691=>"00000010",
  60692=>"00000000",
  60693=>"00000011",
  60694=>"00000001",
  60695=>"11111101",
  60696=>"11111110",
  60697=>"11111101",
  60698=>"00000010",
  60699=>"00000010",
  60700=>"00000000",
  60701=>"00000011",
  60702=>"00000011",
  60703=>"11111111",
  60704=>"00000001",
  60705=>"00000011",
  60706=>"00000001",
  60707=>"00000010",
  60708=>"00000110",
  60709=>"00000110",
  60710=>"11111111",
  60711=>"00000010",
  60712=>"00000010",
  60713=>"11111110",
  60714=>"00000000",
  60715=>"11111110",
  60716=>"00000101",
  60717=>"11111111",
  60718=>"11111101",
  60719=>"00000011",
  60720=>"00000100",
  60721=>"00000011",
  60722=>"00000010",
  60723=>"11111110",
  60724=>"00000010",
  60725=>"11111111",
  60726=>"00000000",
  60727=>"00000110",
  60728=>"00000000",
  60729=>"00000100",
  60730=>"00000010",
  60731=>"11111100",
  60732=>"00000000",
  60733=>"00000010",
  60734=>"11111111",
  60735=>"00000000",
  60736=>"00000010",
  60737=>"11111110",
  60738=>"11111100",
  60739=>"00000001",
  60740=>"11111111",
  60741=>"11111111",
  60742=>"11111101",
  60743=>"11111101",
  60744=>"11111111",
  60745=>"00000001",
  60746=>"11111111",
  60747=>"00000000",
  60748=>"11111110",
  60749=>"00000000",
  60750=>"11111110",
  60751=>"00000100",
  60752=>"11111111",
  60753=>"11111110",
  60754=>"11111110",
  60755=>"11111110",
  60756=>"00000001",
  60757=>"00000010",
  60758=>"11111111",
  60759=>"11111101",
  60760=>"11111110",
  60761=>"11111110",
  60762=>"11111111",
  60763=>"00000001",
  60764=>"00000110",
  60765=>"00000001",
  60766=>"11111101",
  60767=>"00000010",
  60768=>"00000101",
  60769=>"11111100",
  60770=>"11111111",
  60771=>"00000000",
  60772=>"11111111",
  60773=>"00000010",
  60774=>"11111110",
  60775=>"00000010",
  60776=>"11111111",
  60777=>"00000010",
  60778=>"11111111",
  60779=>"11111111",
  60780=>"11111111",
  60781=>"00000001",
  60782=>"11111110",
  60783=>"00000010",
  60784=>"00000001",
  60785=>"00000001",
  60786=>"11111110",
  60787=>"11111110",
  60788=>"00000001",
  60789=>"11111111",
  60790=>"11111111",
  60791=>"00000001",
  60792=>"00000000",
  60793=>"00000001",
  60794=>"00000000",
  60795=>"00000000",
  60796=>"00000000",
  60797=>"00000000",
  60798=>"11111110",
  60799=>"00000001",
  60800=>"00000001",
  60801=>"11111111",
  60802=>"00000001",
  60803=>"00000100",
  60804=>"11111110",
  60805=>"11111101",
  60806=>"00000010",
  60807=>"00000010",
  60808=>"00000100",
  60809=>"11111101",
  60810=>"11111111",
  60811=>"11111110",
  60812=>"00000010",
  60813=>"00000010",
  60814=>"11111110",
  60815=>"00000000",
  60816=>"00000001",
  60817=>"11111110",
  60818=>"00000011",
  60819=>"11111101",
  60820=>"00000000",
  60821=>"11111110",
  60822=>"00000011",
  60823=>"11111111",
  60824=>"11111100",
  60825=>"11111110",
  60826=>"00000010",
  60827=>"11111111",
  60828=>"11111101",
  60829=>"00000010",
  60830=>"00000001",
  60831=>"00000000",
  60832=>"00000010",
  60833=>"00000000",
  60834=>"00000000",
  60835=>"00000011",
  60836=>"11111111",
  60837=>"00000000",
  60838=>"00000001",
  60839=>"11111110",
  60840=>"00000000",
  60841=>"11111101",
  60842=>"00000010",
  60843=>"00000000",
  60844=>"00000100",
  60845=>"00000001",
  60846=>"00000100",
  60847=>"11111111",
  60848=>"11111101",
  60849=>"00000010",
  60850=>"00000000",
  60851=>"00000001",
  60852=>"11111101",
  60853=>"11111111",
  60854=>"00000010",
  60855=>"11111101",
  60856=>"11111100",
  60857=>"00000011",
  60858=>"00000010",
  60859=>"11111110",
  60860=>"00000001",
  60861=>"11111111",
  60862=>"00000001",
  60863=>"11111110",
  60864=>"00000010",
  60865=>"11111111",
  60866=>"11111101",
  60867=>"11111110",
  60868=>"00000010",
  60869=>"00000001",
  60870=>"11111111",
  60871=>"11111101",
  60872=>"00000100",
  60873=>"11111101",
  60874=>"00000000",
  60875=>"00000000",
  60876=>"00000010",
  60877=>"00000000",
  60878=>"11111110",
  60879=>"11111100",
  60880=>"00000000",
  60881=>"00000011",
  60882=>"00000001",
  60883=>"00000000",
  60884=>"00000001",
  60885=>"00000010",
  60886=>"00000010",
  60887=>"00000000",
  60888=>"00000000",
  60889=>"00000000",
  60890=>"00000000",
  60891=>"11111100",
  60892=>"11111100",
  60893=>"11111110",
  60894=>"00000001",
  60895=>"00000011",
  60896=>"11111110",
  60897=>"11111110",
  60898=>"11111110",
  60899=>"11111110",
  60900=>"11111110",
  60901=>"00000001",
  60902=>"11111110",
  60903=>"00000010",
  60904=>"00000010",
  60905=>"00000010",
  60906=>"11111111",
  60907=>"00000010",
  60908=>"11111101",
  60909=>"00000100",
  60910=>"00000011",
  60911=>"00000001",
  60912=>"00000010",
  60913=>"11111111",
  60914=>"11111111",
  60915=>"11111101",
  60916=>"11111111",
  60917=>"11111111",
  60918=>"00000100",
  60919=>"00000010",
  60920=>"00000011",
  60921=>"11111110",
  60922=>"00000100",
  60923=>"00000011",
  60924=>"00000001",
  60925=>"11111110",
  60926=>"00000010",
  60927=>"11111110",
  60928=>"00000001",
  60929=>"00000010",
  60930=>"11111101",
  60931=>"11111111",
  60932=>"11111110",
  60933=>"11111110",
  60934=>"11111111",
  60935=>"11111101",
  60936=>"11111101",
  60937=>"00000011",
  60938=>"00000010",
  60939=>"00000000",
  60940=>"00000010",
  60941=>"00000001",
  60942=>"00000011",
  60943=>"11111111",
  60944=>"11111110",
  60945=>"11111101",
  60946=>"00000011",
  60947=>"11111111",
  60948=>"00000000",
  60949=>"00000000",
  60950=>"11111110",
  60951=>"11111110",
  60952=>"00000011",
  60953=>"11111101",
  60954=>"11111110",
  60955=>"11111111",
  60956=>"00000000",
  60957=>"11111100",
  60958=>"00000001",
  60959=>"00000011",
  60960=>"00000100",
  60961=>"00000001",
  60962=>"00000001",
  60963=>"11111101",
  60964=>"00000100",
  60965=>"00000011",
  60966=>"00000001",
  60967=>"11111101",
  60968=>"00000010",
  60969=>"11111111",
  60970=>"11111111",
  60971=>"00000001",
  60972=>"00000011",
  60973=>"00000001",
  60974=>"00000011",
  60975=>"11111111",
  60976=>"00000001",
  60977=>"00000010",
  60978=>"00000001",
  60979=>"11111111",
  60980=>"11111110",
  60981=>"00000001",
  60982=>"11111111",
  60983=>"11111111",
  60984=>"11111110",
  60985=>"00000010",
  60986=>"00000001",
  60987=>"00000000",
  60988=>"00000001",
  60989=>"11111110",
  60990=>"00000001",
  60991=>"00000100",
  60992=>"00000001",
  60993=>"11111101",
  60994=>"00000100",
  60995=>"00000100",
  60996=>"00000001",
  60997=>"00000010",
  60998=>"00000100",
  60999=>"00000001",
  61000=>"00000011",
  61001=>"11111111",
  61002=>"11111110",
  61003=>"00000100",
  61004=>"00000011",
  61005=>"11111110",
  61006=>"11111110",
  61007=>"00000001",
  61008=>"00000010",
  61009=>"00000000",
  61010=>"00000010",
  61011=>"11111110",
  61012=>"00000001",
  61013=>"11111111",
  61014=>"11111111",
  61015=>"11111111",
  61016=>"00000010",
  61017=>"00000100",
  61018=>"11111111",
  61019=>"00000001",
  61020=>"11111110",
  61021=>"00000010",
  61022=>"11111110",
  61023=>"11111101",
  61024=>"00000011",
  61025=>"11111110",
  61026=>"00000010",
  61027=>"00000001",
  61028=>"00000011",
  61029=>"00000100",
  61030=>"00000000",
  61031=>"00000000",
  61032=>"11111110",
  61033=>"11111111",
  61034=>"00000000",
  61035=>"11111110",
  61036=>"00000001",
  61037=>"00000000",
  61038=>"00000100",
  61039=>"11111111",
  61040=>"11111101",
  61041=>"00000001",
  61042=>"11111111",
  61043=>"00000101",
  61044=>"00000010",
  61045=>"00000010",
  61046=>"00000000",
  61047=>"00000001",
  61048=>"00000010",
  61049=>"00000001",
  61050=>"11111111",
  61051=>"11111100",
  61052=>"00000001",
  61053=>"00000100",
  61054=>"11111101",
  61055=>"00000000",
  61056=>"00000011",
  61057=>"00000101",
  61058=>"11111111",
  61059=>"00000010",
  61060=>"00000101",
  61061=>"00000010",
  61062=>"11111111",
  61063=>"11111110",
  61064=>"11111111",
  61065=>"11111101",
  61066=>"11111110",
  61067=>"00000001",
  61068=>"00000001",
  61069=>"11111101",
  61070=>"11111110",
  61071=>"11111101",
  61072=>"00000000",
  61073=>"00000011",
  61074=>"00000110",
  61075=>"00000001",
  61076=>"00000001",
  61077=>"11111110",
  61078=>"00000000",
  61079=>"00000000",
  61080=>"11111100",
  61081=>"00000010",
  61082=>"11111111",
  61083=>"00000001",
  61084=>"00000011",
  61085=>"00000010",
  61086=>"11111101",
  61087=>"00000010",
  61088=>"00000001",
  61089=>"11111110",
  61090=>"11111110",
  61091=>"00000000",
  61092=>"11111110",
  61093=>"00000010",
  61094=>"00000001",
  61095=>"11111101",
  61096=>"00000010",
  61097=>"00000101",
  61098=>"11111110",
  61099=>"00000010",
  61100=>"00000011",
  61101=>"00000000",
  61102=>"00000010",
  61103=>"00000000",
  61104=>"11111110",
  61105=>"00000000",
  61106=>"11111110",
  61107=>"00000010",
  61108=>"00000010",
  61109=>"11111111",
  61110=>"00000001",
  61111=>"00000010",
  61112=>"00000001",
  61113=>"11111101",
  61114=>"00000000",
  61115=>"11111110",
  61116=>"00000011",
  61117=>"00000001",
  61118=>"00000101",
  61119=>"00000000",
  61120=>"00000011",
  61121=>"11111111",
  61122=>"11111101",
  61123=>"11111101",
  61124=>"11111111",
  61125=>"00000001",
  61126=>"11111111",
  61127=>"11111111",
  61128=>"00000001",
  61129=>"00000001",
  61130=>"00000001",
  61131=>"00000001",
  61132=>"11111100",
  61133=>"00000000",
  61134=>"11111110",
  61135=>"00000000",
  61136=>"00000000",
  61137=>"11111111",
  61138=>"00000000",
  61139=>"11111110",
  61140=>"00000011",
  61141=>"00000101",
  61142=>"11111110",
  61143=>"11111101",
  61144=>"00000010",
  61145=>"00000001",
  61146=>"00000001",
  61147=>"00000011",
  61148=>"11111110",
  61149=>"00000000",
  61150=>"00000000",
  61151=>"11111110",
  61152=>"00000001",
  61153=>"00000000",
  61154=>"11111101",
  61155=>"00000011",
  61156=>"11111110",
  61157=>"00000001",
  61158=>"11111110",
  61159=>"00000000",
  61160=>"00000000",
  61161=>"11111110",
  61162=>"11111110",
  61163=>"11111111",
  61164=>"00000011",
  61165=>"11111111",
  61166=>"00000100",
  61167=>"11111110",
  61168=>"00000011",
  61169=>"11111110",
  61170=>"00000001",
  61171=>"00000001",
  61172=>"11111101",
  61173=>"00000001",
  61174=>"00000001",
  61175=>"11111101",
  61176=>"11111101",
  61177=>"11111111",
  61178=>"00000010",
  61179=>"00000000",
  61180=>"00000001",
  61181=>"11111101",
  61182=>"00000010",
  61183=>"00000000",
  61184=>"00000001",
  61185=>"00000100",
  61186=>"11111110",
  61187=>"00000011",
  61188=>"00000000",
  61189=>"00000001",
  61190=>"11111111",
  61191=>"11111110",
  61192=>"00000000",
  61193=>"00000001",
  61194=>"00000000",
  61195=>"00000001",
  61196=>"11111101",
  61197=>"11111110",
  61198=>"11111111",
  61199=>"11111110",
  61200=>"11111111",
  61201=>"00000001",
  61202=>"00000010",
  61203=>"00000000",
  61204=>"11111110",
  61205=>"00000001",
  61206=>"00000000",
  61207=>"00000001",
  61208=>"11111101",
  61209=>"11111111",
  61210=>"00000110",
  61211=>"00000010",
  61212=>"00000000",
  61213=>"11111111",
  61214=>"11111101",
  61215=>"11111110",
  61216=>"11111111",
  61217=>"00000001",
  61218=>"11111110",
  61219=>"11111101",
  61220=>"11111110",
  61221=>"00000010",
  61222=>"11111100",
  61223=>"11111100",
  61224=>"11111110",
  61225=>"11111111",
  61226=>"00000011",
  61227=>"00000001",
  61228=>"00000011",
  61229=>"11111101",
  61230=>"00000010",
  61231=>"00000101",
  61232=>"11111111",
  61233=>"00000000",
  61234=>"11111100",
  61235=>"00000100",
  61236=>"00000000",
  61237=>"00000100",
  61238=>"00000000",
  61239=>"00000000",
  61240=>"11111111",
  61241=>"00000000",
  61242=>"11111110",
  61243=>"11111101",
  61244=>"00000010",
  61245=>"11111110",
  61246=>"00000000",
  61247=>"00000000",
  61248=>"00000011",
  61249=>"00000010",
  61250=>"00000001",
  61251=>"11111101",
  61252=>"11111110",
  61253=>"00000000",
  61254=>"11111101",
  61255=>"00000000",
  61256=>"11111101",
  61257=>"00000011",
  61258=>"11111110",
  61259=>"11111100",
  61260=>"00000011",
  61261=>"11111111",
  61262=>"00000000",
  61263=>"00000000",
  61264=>"11111101",
  61265=>"00000011",
  61266=>"00000000",
  61267=>"11111111",
  61268=>"00000010",
  61269=>"11111100",
  61270=>"00000010",
  61271=>"11111101",
  61272=>"11111110",
  61273=>"11111110",
  61274=>"11111110",
  61275=>"11111110",
  61276=>"11111111",
  61277=>"00000001",
  61278=>"00000100",
  61279=>"11111110",
  61280=>"11111101",
  61281=>"11111110",
  61282=>"11111101",
  61283=>"11111101",
  61284=>"00000010",
  61285=>"00000000",
  61286=>"00000000",
  61287=>"11111101",
  61288=>"11111101",
  61289=>"00000010",
  61290=>"11111110",
  61291=>"11111110",
  61292=>"11111110",
  61293=>"00000000",
  61294=>"00000011",
  61295=>"00000010",
  61296=>"00000001",
  61297=>"11111111",
  61298=>"00000010",
  61299=>"00000010",
  61300=>"11111111",
  61301=>"00000001",
  61302=>"11111110",
  61303=>"00000001",
  61304=>"00000001",
  61305=>"00000000",
  61306=>"11111110",
  61307=>"11111101",
  61308=>"11111101",
  61309=>"11111101",
  61310=>"11111110",
  61311=>"11111101",
  61312=>"00000000",
  61313=>"11111111",
  61314=>"11111110",
  61315=>"11111111",
  61316=>"00000001",
  61317=>"00000010",
  61318=>"11111110",
  61319=>"00000010",
  61320=>"00000001",
  61321=>"11111110",
  61322=>"11111111",
  61323=>"11111110",
  61324=>"11111101",
  61325=>"11111101",
  61326=>"00000000",
  61327=>"00000001",
  61328=>"00000000",
  61329=>"11111110",
  61330=>"11111100",
  61331=>"00000010",
  61332=>"11111101",
  61333=>"00000000",
  61334=>"00000001",
  61335=>"00000001",
  61336=>"11111100",
  61337=>"11111100",
  61338=>"00000011",
  61339=>"11111101",
  61340=>"11111101",
  61341=>"11111101",
  61342=>"11111100",
  61343=>"00000000",
  61344=>"00000010",
  61345=>"00000000",
  61346=>"00000010",
  61347=>"11111111",
  61348=>"11111111",
  61349=>"11111101",
  61350=>"11111101",
  61351=>"11111110",
  61352=>"11111111",
  61353=>"11111110",
  61354=>"11111101",
  61355=>"00000000",
  61356=>"00000000",
  61357=>"00000001",
  61358=>"11111111",
  61359=>"00000001",
  61360=>"00000100",
  61361=>"11111110",
  61362=>"00000000",
  61363=>"00000011",
  61364=>"00000001",
  61365=>"11111110",
  61366=>"00000010",
  61367=>"00000010",
  61368=>"11111111",
  61369=>"00000000",
  61370=>"00000100",
  61371=>"00000000",
  61372=>"00000001",
  61373=>"11111101",
  61374=>"11111101",
  61375=>"11111110",
  61376=>"00000000",
  61377=>"00000010",
  61378=>"11111111",
  61379=>"00000100",
  61380=>"00000010",
  61381=>"00000001",
  61382=>"11111110",
  61383=>"11111111",
  61384=>"00000001",
  61385=>"11111110",
  61386=>"00000011",
  61387=>"11111111",
  61388=>"00000010",
  61389=>"00000100",
  61390=>"11111101",
  61391=>"00000000",
  61392=>"11111111",
  61393=>"00000001",
  61394=>"00000011",
  61395=>"11111110",
  61396=>"11111111",
  61397=>"00000000",
  61398=>"00000100",
  61399=>"00000001",
  61400=>"11111110",
  61401=>"00000011",
  61402=>"11111101",
  61403=>"00000010",
  61404=>"11111100",
  61405=>"11111101",
  61406=>"11111110",
  61407=>"00000100",
  61408=>"00000110",
  61409=>"00000001",
  61410=>"00000001",
  61411=>"00000010",
  61412=>"11111110",
  61413=>"00000011",
  61414=>"00000010",
  61415=>"11111101",
  61416=>"11111101",
  61417=>"00000001",
  61418=>"00000000",
  61419=>"00000011",
  61420=>"00000000",
  61421=>"00000000",
  61422=>"00000000",
  61423=>"00000001",
  61424=>"11111110",
  61425=>"11111111",
  61426=>"11111101",
  61427=>"11111111",
  61428=>"00000010",
  61429=>"11111100",
  61430=>"00000101",
  61431=>"11111101",
  61432=>"11111101",
  61433=>"11111110",
  61434=>"00000100",
  61435=>"11111101",
  61436=>"11111101",
  61437=>"11111101",
  61438=>"00000100",
  61439=>"11111111",
  61440=>"00000001",
  61441=>"00000000",
  61442=>"11111101",
  61443=>"11111101",
  61444=>"00000000",
  61445=>"00000110",
  61446=>"11111110",
  61447=>"11111111",
  61448=>"00000001",
  61449=>"00000000",
  61450=>"11111111",
  61451=>"11111110",
  61452=>"11111101",
  61453=>"11111101",
  61454=>"11111101",
  61455=>"11111101",
  61456=>"00000001",
  61457=>"11111110",
  61458=>"00000000",
  61459=>"00000001",
  61460=>"11111110",
  61461=>"00000000",
  61462=>"00000000",
  61463=>"11111110",
  61464=>"00000001",
  61465=>"00000001",
  61466=>"00000000",
  61467=>"00000001",
  61468=>"00000001",
  61469=>"11111110",
  61470=>"11111101",
  61471=>"11111111",
  61472=>"00000100",
  61473=>"11111110",
  61474=>"00000000",
  61475=>"00000000",
  61476=>"11111110",
  61477=>"00000000",
  61478=>"11111101",
  61479=>"00000001",
  61480=>"11111110",
  61481=>"11111111",
  61482=>"00000111",
  61483=>"11111110",
  61484=>"00000001",
  61485=>"11111110",
  61486=>"11111111",
  61487=>"11111110",
  61488=>"11111110",
  61489=>"00000011",
  61490=>"00000001",
  61491=>"11111111",
  61492=>"11111111",
  61493=>"11111111",
  61494=>"00000010",
  61495=>"00000010",
  61496=>"00000101",
  61497=>"11111100",
  61498=>"00000010",
  61499=>"00000000",
  61500=>"11111111",
  61501=>"11111110",
  61502=>"11111101",
  61503=>"00000001",
  61504=>"11111101",
  61505=>"00000000",
  61506=>"00000000",
  61507=>"11111111",
  61508=>"11111110",
  61509=>"00000010",
  61510=>"11111101",
  61511=>"00000000",
  61512=>"11111111",
  61513=>"11111101",
  61514=>"00000001",
  61515=>"00000010",
  61516=>"11111101",
  61517=>"00000011",
  61518=>"11111110",
  61519=>"11111110",
  61520=>"00000011",
  61521=>"00000010",
  61522=>"00000001",
  61523=>"00000000",
  61524=>"11111111",
  61525=>"11111110",
  61526=>"11111101",
  61527=>"11111111",
  61528=>"11111111",
  61529=>"11111101",
  61530=>"00000010",
  61531=>"00000000",
  61532=>"11111101",
  61533=>"00000011",
  61534=>"11111101",
  61535=>"11111110",
  61536=>"00000000",
  61537=>"00000001",
  61538=>"00000010",
  61539=>"00000010",
  61540=>"00000001",
  61541=>"00000010",
  61542=>"00000100",
  61543=>"00000010",
  61544=>"00000001",
  61545=>"00000010",
  61546=>"00000010",
  61547=>"00000010",
  61548=>"11111111",
  61549=>"11111110",
  61550=>"11111110",
  61551=>"11111111",
  61552=>"11111101",
  61553=>"00000101",
  61554=>"00000000",
  61555=>"00000011",
  61556=>"11111110",
  61557=>"00000010",
  61558=>"00000001",
  61559=>"00000000",
  61560=>"00000000",
  61561=>"00000000",
  61562=>"00000000",
  61563=>"00000000",
  61564=>"00000000",
  61565=>"11111111",
  61566=>"11111101",
  61567=>"11111110",
  61568=>"11111101",
  61569=>"00000101",
  61570=>"00000110",
  61571=>"00000000",
  61572=>"00000011",
  61573=>"00000001",
  61574=>"00000001",
  61575=>"00000010",
  61576=>"11111111",
  61577=>"11111111",
  61578=>"11111111",
  61579=>"00000010",
  61580=>"11111111",
  61581=>"00000001",
  61582=>"11111100",
  61583=>"00000000",
  61584=>"00000000",
  61585=>"00000000",
  61586=>"00000010",
  61587=>"00000010",
  61588=>"11111101",
  61589=>"00000000",
  61590=>"11111111",
  61591=>"00000001",
  61592=>"11111110",
  61593=>"00000000",
  61594=>"11111111",
  61595=>"00000111",
  61596=>"00000010",
  61597=>"00000011",
  61598=>"11111101",
  61599=>"00000011",
  61600=>"11111111",
  61601=>"00000001",
  61602=>"00000000",
  61603=>"00000011",
  61604=>"00000000",
  61605=>"11111101",
  61606=>"00000000",
  61607=>"00000100",
  61608=>"00000001",
  61609=>"11111100",
  61610=>"00000001",
  61611=>"11111110",
  61612=>"00000001",
  61613=>"00000000",
  61614=>"00000010",
  61615=>"11111110",
  61616=>"00000000",
  61617=>"00000001",
  61618=>"00000000",
  61619=>"11111111",
  61620=>"00000001",
  61621=>"00000000",
  61622=>"00000001",
  61623=>"11111111",
  61624=>"11111101",
  61625=>"00000000",
  61626=>"11111111",
  61627=>"00000101",
  61628=>"11111101",
  61629=>"11111111",
  61630=>"00000001",
  61631=>"00000000",
  61632=>"11111101",
  61633=>"11111111",
  61634=>"11111111",
  61635=>"00000011",
  61636=>"00000000",
  61637=>"00000100",
  61638=>"00000001",
  61639=>"11111110",
  61640=>"00000001",
  61641=>"11111101",
  61642=>"11111111",
  61643=>"00000000",
  61644=>"11111101",
  61645=>"11111110",
  61646=>"11111101",
  61647=>"11111111",
  61648=>"00000001",
  61649=>"11111110",
  61650=>"00000001",
  61651=>"00000010",
  61652=>"00000000",
  61653=>"11111111",
  61654=>"00000000",
  61655=>"00000001",
  61656=>"11111110",
  61657=>"00000010",
  61658=>"00000000",
  61659=>"00000000",
  61660=>"11111101",
  61661=>"11111111",
  61662=>"00000000",
  61663=>"11111110",
  61664=>"00000001",
  61665=>"00000010",
  61666=>"11111101",
  61667=>"11111110",
  61668=>"00000011",
  61669=>"00000001",
  61670=>"00000001",
  61671=>"00000010",
  61672=>"11111110",
  61673=>"00000001",
  61674=>"00000001",
  61675=>"11111111",
  61676=>"00000011",
  61677=>"00000001",
  61678=>"00000000",
  61679=>"00000001",
  61680=>"11111111",
  61681=>"11111110",
  61682=>"00000001",
  61683=>"11111110",
  61684=>"00000010",
  61685=>"11111101",
  61686=>"00000010",
  61687=>"00000011",
  61688=>"00000010",
  61689=>"00000000",
  61690=>"11111101",
  61691=>"11111101",
  61692=>"00000100",
  61693=>"00000000",
  61694=>"11111110",
  61695=>"11111111",
  61696=>"00000000",
  61697=>"00000000",
  61698=>"11111101",
  61699=>"00000010",
  61700=>"11111111",
  61701=>"00000000",
  61702=>"00000001",
  61703=>"00000001",
  61704=>"11111110",
  61705=>"00000011",
  61706=>"00000011",
  61707=>"11111111",
  61708=>"11111110",
  61709=>"11111110",
  61710=>"00000010",
  61711=>"00000001",
  61712=>"11111110",
  61713=>"00000000",
  61714=>"11111101",
  61715=>"11111101",
  61716=>"00000001",
  61717=>"11111110",
  61718=>"11111101",
  61719=>"00000010",
  61720=>"00000000",
  61721=>"11111101",
  61722=>"00000001",
  61723=>"00000001",
  61724=>"00000100",
  61725=>"11111101",
  61726=>"11111111",
  61727=>"11111110",
  61728=>"00000000",
  61729=>"00000000",
  61730=>"00000010",
  61731=>"00000010",
  61732=>"00000100",
  61733=>"11111100",
  61734=>"11111111",
  61735=>"11111111",
  61736=>"00000010",
  61737=>"11111110",
  61738=>"00000001",
  61739=>"00000100",
  61740=>"11111111",
  61741=>"00000000",
  61742=>"00000001",
  61743=>"00000011",
  61744=>"11111101",
  61745=>"00000001",
  61746=>"00000011",
  61747=>"00000001",
  61748=>"00000101",
  61749=>"00000010",
  61750=>"00000000",
  61751=>"00000001",
  61752=>"00000101",
  61753=>"11111110",
  61754=>"00000000",
  61755=>"00000000",
  61756=>"11111111",
  61757=>"00000001",
  61758=>"00000011",
  61759=>"00000011",
  61760=>"11111111",
  61761=>"00000001",
  61762=>"00000010",
  61763=>"11111110",
  61764=>"00000001",
  61765=>"00000001",
  61766=>"11111110",
  61767=>"00000000",
  61768=>"11111111",
  61769=>"00000001",
  61770=>"11111111",
  61771=>"00000001",
  61772=>"11111110",
  61773=>"11111110",
  61774=>"00000001",
  61775=>"11111111",
  61776=>"00000011",
  61777=>"11111111",
  61778=>"00000001",
  61779=>"00000010",
  61780=>"11111110",
  61781=>"00000001",
  61782=>"00000001",
  61783=>"11111101",
  61784=>"00000010",
  61785=>"00000010",
  61786=>"00000001",
  61787=>"11111110",
  61788=>"00000010",
  61789=>"00000001",
  61790=>"11111101",
  61791=>"00000010",
  61792=>"11111111",
  61793=>"11111101",
  61794=>"11111101",
  61795=>"11111101",
  61796=>"00000000",
  61797=>"00000000",
  61798=>"00000000",
  61799=>"11111101",
  61800=>"00000000",
  61801=>"00000010",
  61802=>"00000001",
  61803=>"00000000",
  61804=>"11111111",
  61805=>"11111111",
  61806=>"11111101",
  61807=>"11111110",
  61808=>"00000010",
  61809=>"11111111",
  61810=>"11111111",
  61811=>"00000010",
  61812=>"00000001",
  61813=>"00000000",
  61814=>"00000001",
  61815=>"00000001",
  61816=>"00000000",
  61817=>"11111111",
  61818=>"00000001",
  61819=>"11111111",
  61820=>"11111101",
  61821=>"11111100",
  61822=>"11111111",
  61823=>"00000000",
  61824=>"11111110",
  61825=>"11111111",
  61826=>"00000000",
  61827=>"00000001",
  61828=>"00000010",
  61829=>"11111110",
  61830=>"00000000",
  61831=>"11111110",
  61832=>"11111111",
  61833=>"00000000",
  61834=>"00000010",
  61835=>"11111111",
  61836=>"00000001",
  61837=>"00000011",
  61838=>"00000001",
  61839=>"11111111",
  61840=>"11111110",
  61841=>"11111111",
  61842=>"11111111",
  61843=>"11111110",
  61844=>"11111101",
  61845=>"11111101",
  61846=>"00000011",
  61847=>"00000000",
  61848=>"11111111",
  61849=>"00000010",
  61850=>"00000010",
  61851=>"00000001",
  61852=>"00000010",
  61853=>"11111110",
  61854=>"11111101",
  61855=>"00000010",
  61856=>"00000000",
  61857=>"00000001",
  61858=>"00000001",
  61859=>"11111111",
  61860=>"00000001",
  61861=>"11111110",
  61862=>"00000000",
  61863=>"11111110",
  61864=>"00000010",
  61865=>"11111111",
  61866=>"11111111",
  61867=>"00000001",
  61868=>"00000001",
  61869=>"00000100",
  61870=>"11111101",
  61871=>"00000001",
  61872=>"11111110",
  61873=>"00000001",
  61874=>"00000010",
  61875=>"11111111",
  61876=>"11111110",
  61877=>"11111111",
  61878=>"11111110",
  61879=>"00000001",
  61880=>"00000000",
  61881=>"11111101",
  61882=>"00000000",
  61883=>"11111111",
  61884=>"11111111",
  61885=>"11111111",
  61886=>"11111110",
  61887=>"00000010",
  61888=>"11111110",
  61889=>"00000100",
  61890=>"11111110",
  61891=>"11111100",
  61892=>"11111110",
  61893=>"11111110",
  61894=>"11111101",
  61895=>"00000011",
  61896=>"00000000",
  61897=>"00000000",
  61898=>"00000010",
  61899=>"11111100",
  61900=>"00000000",
  61901=>"00000000",
  61902=>"00000001",
  61903=>"00000101",
  61904=>"00000011",
  61905=>"11111111",
  61906=>"11111111",
  61907=>"11111101",
  61908=>"11111101",
  61909=>"00000001",
  61910=>"11111101",
  61911=>"00000001",
  61912=>"00000001",
  61913=>"00000000",
  61914=>"00000010",
  61915=>"00000010",
  61916=>"11111101",
  61917=>"11111101",
  61918=>"00000010",
  61919=>"11111110",
  61920=>"00000011",
  61921=>"11111110",
  61922=>"11111111",
  61923=>"11111110",
  61924=>"11111111",
  61925=>"11111111",
  61926=>"11111111",
  61927=>"00000010",
  61928=>"11111111",
  61929=>"11111111",
  61930=>"00000100",
  61931=>"00000001",
  61932=>"00000010",
  61933=>"00000100",
  61934=>"00000011",
  61935=>"00000101",
  61936=>"00000010",
  61937=>"11111110",
  61938=>"00000010",
  61939=>"00000011",
  61940=>"00000000",
  61941=>"00000101",
  61942=>"11111110",
  61943=>"11111110",
  61944=>"11111111",
  61945=>"11111101",
  61946=>"11111101",
  61947=>"00000000",
  61948=>"11111101",
  61949=>"00000010",
  61950=>"00000101",
  61951=>"11111110",
  61952=>"11111110",
  61953=>"11111110",
  61954=>"11111111",
  61955=>"00000011",
  61956=>"00000010",
  61957=>"11111111",
  61958=>"11111110",
  61959=>"00000011",
  61960=>"00000010",
  61961=>"11111110",
  61962=>"00000001",
  61963=>"00000011",
  61964=>"00000011",
  61965=>"11111111",
  61966=>"00000001",
  61967=>"00000000",
  61968=>"00000001",
  61969=>"00000000",
  61970=>"00000001",
  61971=>"11111101",
  61972=>"11111110",
  61973=>"11111101",
  61974=>"11111110",
  61975=>"00000011",
  61976=>"11111110",
  61977=>"11111111",
  61978=>"00000000",
  61979=>"11111111",
  61980=>"11111111",
  61981=>"00000000",
  61982=>"00000001",
  61983=>"11111111",
  61984=>"11111110",
  61985=>"11111101",
  61986=>"00000011",
  61987=>"11111110",
  61988=>"00000001",
  61989=>"00000001",
  61990=>"11111110",
  61991=>"11111111",
  61992=>"00000000",
  61993=>"00000010",
  61994=>"11111110",
  61995=>"11111111",
  61996=>"11111110",
  61997=>"00000010",
  61998=>"11111110",
  61999=>"00000010",
  62000=>"11111101",
  62001=>"00000001",
  62002=>"00000001",
  62003=>"00000010",
  62004=>"00000000",
  62005=>"00000010",
  62006=>"00000010",
  62007=>"00000011",
  62008=>"00000000",
  62009=>"11111111",
  62010=>"11111111",
  62011=>"00000001",
  62012=>"00000000",
  62013=>"00000010",
  62014=>"11111110",
  62015=>"11111110",
  62016=>"00000001",
  62017=>"11111110",
  62018=>"11111110",
  62019=>"00000000",
  62020=>"00000000",
  62021=>"00000000",
  62022=>"00000110",
  62023=>"11111101",
  62024=>"11111110",
  62025=>"00000010",
  62026=>"11111111",
  62027=>"11111111",
  62028=>"00000001",
  62029=>"11111111",
  62030=>"00000011",
  62031=>"11111101",
  62032=>"00000010",
  62033=>"00000000",
  62034=>"00000001",
  62035=>"00000001",
  62036=>"00000000",
  62037=>"00000000",
  62038=>"00000001",
  62039=>"00000101",
  62040=>"00000000",
  62041=>"00000001",
  62042=>"00000001",
  62043=>"11111111",
  62044=>"00000000",
  62045=>"00000001",
  62046=>"11111111",
  62047=>"00000000",
  62048=>"11111101",
  62049=>"00000000",
  62050=>"11111101",
  62051=>"00000000",
  62052=>"00000101",
  62053=>"00000001",
  62054=>"00000001",
  62055=>"00000010",
  62056=>"00000001",
  62057=>"00000011",
  62058=>"11111110",
  62059=>"11111111",
  62060=>"11111111",
  62061=>"11111101",
  62062=>"00000000",
  62063=>"11111110",
  62064=>"00000010",
  62065=>"11111110",
  62066=>"00000010",
  62067=>"11111110",
  62068=>"00000001",
  62069=>"00000000",
  62070=>"11111110",
  62071=>"11111111",
  62072=>"11111110",
  62073=>"00000010",
  62074=>"00000001",
  62075=>"00000010",
  62076=>"00000001",
  62077=>"00000100",
  62078=>"11111110",
  62079=>"00000000",
  62080=>"00000000",
  62081=>"00000001",
  62082=>"11111101",
  62083=>"11111111",
  62084=>"11111101",
  62085=>"00000001",
  62086=>"11111110",
  62087=>"00000010",
  62088=>"00000001",
  62089=>"11111110",
  62090=>"11111111",
  62091=>"11111101",
  62092=>"11111111",
  62093=>"00000010",
  62094=>"11111111",
  62095=>"11111101",
  62096=>"11111110",
  62097=>"11111111",
  62098=>"11111111",
  62099=>"00000010",
  62100=>"00000001",
  62101=>"11111111",
  62102=>"11111110",
  62103=>"00000011",
  62104=>"11111101",
  62105=>"00000001",
  62106=>"00000000",
  62107=>"00000001",
  62108=>"00000101",
  62109=>"11111101",
  62110=>"11111111",
  62111=>"11111111",
  62112=>"00000000",
  62113=>"00000001",
  62114=>"00000000",
  62115=>"11111111",
  62116=>"11111111",
  62117=>"00000000",
  62118=>"11111111",
  62119=>"11111101",
  62120=>"00000100",
  62121=>"00000100",
  62122=>"11111110",
  62123=>"11111110",
  62124=>"00000001",
  62125=>"00000000",
  62126=>"11111110",
  62127=>"00000011",
  62128=>"11111101",
  62129=>"11111111",
  62130=>"00000001",
  62131=>"00000010",
  62132=>"00000011",
  62133=>"11111110",
  62134=>"00000100",
  62135=>"00000100",
  62136=>"00000100",
  62137=>"00000001",
  62138=>"00000001",
  62139=>"00000011",
  62140=>"00000001",
  62141=>"11111101",
  62142=>"11111101",
  62143=>"11111110",
  62144=>"00000001",
  62145=>"00000001",
  62146=>"00000010",
  62147=>"00000101",
  62148=>"00000010",
  62149=>"11111110",
  62150=>"00000011",
  62151=>"00000000",
  62152=>"11111101",
  62153=>"11111110",
  62154=>"00000011",
  62155=>"00000100",
  62156=>"00000001",
  62157=>"11111110",
  62158=>"00000010",
  62159=>"00000001",
  62160=>"00000001",
  62161=>"00000011",
  62162=>"00000001",
  62163=>"11111110",
  62164=>"00000101",
  62165=>"00000001",
  62166=>"11111111",
  62167=>"00000010",
  62168=>"11111110",
  62169=>"11111101",
  62170=>"00000000",
  62171=>"11111100",
  62172=>"11111101",
  62173=>"00000001",
  62174=>"11111110",
  62175=>"00000011",
  62176=>"11111101",
  62177=>"00000100",
  62178=>"00000001",
  62179=>"00000010",
  62180=>"11111101",
  62181=>"00000000",
  62182=>"00000001",
  62183=>"11111100",
  62184=>"00000001",
  62185=>"00000001",
  62186=>"11111101",
  62187=>"00000010",
  62188=>"00000010",
  62189=>"00000111",
  62190=>"00000000",
  62191=>"11111111",
  62192=>"00000000",
  62193=>"11111101",
  62194=>"00000011",
  62195=>"00000000",
  62196=>"00000010",
  62197=>"11111101",
  62198=>"11111111",
  62199=>"11111101",
  62200=>"11111101",
  62201=>"00000100",
  62202=>"11111110",
  62203=>"11111110",
  62204=>"00000000",
  62205=>"11111110",
  62206=>"00000010",
  62207=>"00000000",
  62208=>"00000010",
  62209=>"00000000",
  62210=>"00000011",
  62211=>"11111101",
  62212=>"11111110",
  62213=>"11111111",
  62214=>"11111111",
  62215=>"11111101",
  62216=>"11111101",
  62217=>"11111101",
  62218=>"00000001",
  62219=>"00000001",
  62220=>"11111101",
  62221=>"11111110",
  62222=>"11111111",
  62223=>"00000010",
  62224=>"11111110",
  62225=>"00000010",
  62226=>"11111111",
  62227=>"00000010",
  62228=>"11111110",
  62229=>"00000000",
  62230=>"11111100",
  62231=>"11111101",
  62232=>"00000010",
  62233=>"11111100",
  62234=>"11111111",
  62235=>"11111110",
  62236=>"11111111",
  62237=>"11111110",
  62238=>"00000011",
  62239=>"00000000",
  62240=>"00000100",
  62241=>"00000100",
  62242=>"11111110",
  62243=>"11111110",
  62244=>"11111111",
  62245=>"00000000",
  62246=>"00000000",
  62247=>"11111101",
  62248=>"00000000",
  62249=>"11111101",
  62250=>"00000101",
  62251=>"00000010",
  62252=>"11111111",
  62253=>"11111110",
  62254=>"00000000",
  62255=>"00000000",
  62256=>"11111101",
  62257=>"00000111",
  62258=>"00000001",
  62259=>"00000000",
  62260=>"00000001",
  62261=>"00000000",
  62262=>"11111111",
  62263=>"11111111",
  62264=>"00000000",
  62265=>"00000000",
  62266=>"00000011",
  62267=>"00000010",
  62268=>"00000001",
  62269=>"00000001",
  62270=>"11111101",
  62271=>"00000000",
  62272=>"11111111",
  62273=>"11111111",
  62274=>"00000010",
  62275=>"11111111",
  62276=>"00000011",
  62277=>"11111110",
  62278=>"11111111",
  62279=>"11111111",
  62280=>"11111111",
  62281=>"00000000",
  62282=>"11111110",
  62283=>"00000000",
  62284=>"00000000",
  62285=>"00000001",
  62286=>"11111111",
  62287=>"00000000",
  62288=>"00000000",
  62289=>"00000001",
  62290=>"00000010",
  62291=>"00000000",
  62292=>"11111101",
  62293=>"00000011",
  62294=>"00000010",
  62295=>"00000100",
  62296=>"11111111",
  62297=>"00000001",
  62298=>"11111111",
  62299=>"11111101",
  62300=>"11111111",
  62301=>"00000011",
  62302=>"00000100",
  62303=>"00000010",
  62304=>"11111110",
  62305=>"00000000",
  62306=>"11111101",
  62307=>"11111110",
  62308=>"00000010",
  62309=>"00000001",
  62310=>"00000000",
  62311=>"00000001",
  62312=>"11111110",
  62313=>"00000000",
  62314=>"11111101",
  62315=>"00000000",
  62316=>"11111111",
  62317=>"11111110",
  62318=>"11111110",
  62319=>"11111110",
  62320=>"00000010",
  62321=>"11111100",
  62322=>"00000000",
  62323=>"11111101",
  62324=>"11111101",
  62325=>"00000010",
  62326=>"00000010",
  62327=>"11111111",
  62328=>"11111110",
  62329=>"00000000",
  62330=>"00000000",
  62331=>"00000000",
  62332=>"11111110",
  62333=>"00000000",
  62334=>"11111111",
  62335=>"00000001",
  62336=>"11111110",
  62337=>"11111111",
  62338=>"00000000",
  62339=>"11111111",
  62340=>"11111110",
  62341=>"11111101",
  62342=>"00000000",
  62343=>"11111111",
  62344=>"00000001",
  62345=>"00000100",
  62346=>"11111110",
  62347=>"11111111",
  62348=>"00000010",
  62349=>"11111110",
  62350=>"00000000",
  62351=>"00000001",
  62352=>"11111111",
  62353=>"11111101",
  62354=>"00000000",
  62355=>"00000001",
  62356=>"00000011",
  62357=>"11111111",
  62358=>"00000100",
  62359=>"00000001",
  62360=>"00000010",
  62361=>"00000001",
  62362=>"11111110",
  62363=>"11111110",
  62364=>"11111100",
  62365=>"00000001",
  62366=>"00000011",
  62367=>"11111110",
  62368=>"11111101",
  62369=>"00000000",
  62370=>"11111110",
  62371=>"11111111",
  62372=>"00000000",
  62373=>"00000101",
  62374=>"00000000",
  62375=>"00000001",
  62376=>"00000000",
  62377=>"00000010",
  62378=>"00000010",
  62379=>"00000000",
  62380=>"11111110",
  62381=>"11111110",
  62382=>"11111101",
  62383=>"00000000",
  62384=>"11111111",
  62385=>"00000010",
  62386=>"11111101",
  62387=>"00000110",
  62388=>"11111101",
  62389=>"00000010",
  62390=>"00000010",
  62391=>"11111100",
  62392=>"00000000",
  62393=>"00000100",
  62394=>"11111110",
  62395=>"00000001",
  62396=>"00000001",
  62397=>"11111110",
  62398=>"00000001",
  62399=>"00000010",
  62400=>"00000001",
  62401=>"11111110",
  62402=>"11111101",
  62403=>"11111110",
  62404=>"11111110",
  62405=>"00000010",
  62406=>"00000001",
  62407=>"00000001",
  62408=>"00000011",
  62409=>"00000001",
  62410=>"00000010",
  62411=>"00000010",
  62412=>"00000011",
  62413=>"11111110",
  62414=>"00000000",
  62415=>"11111101",
  62416=>"00000010",
  62417=>"00000000",
  62418=>"00000101",
  62419=>"00000001",
  62420=>"00000000",
  62421=>"00000000",
  62422=>"00000110",
  62423=>"00000010",
  62424=>"00000001",
  62425=>"11111110",
  62426=>"11111111",
  62427=>"11111110",
  62428=>"00000000",
  62429=>"11111101",
  62430=>"00000011",
  62431=>"00000001",
  62432=>"11111110",
  62433=>"00000100",
  62434=>"11111110",
  62435=>"11111110",
  62436=>"00000001",
  62437=>"00000110",
  62438=>"00000001",
  62439=>"11111111",
  62440=>"11111111",
  62441=>"00000010",
  62442=>"11111101",
  62443=>"11111110",
  62444=>"00000010",
  62445=>"11111110",
  62446=>"11111101",
  62447=>"00000000",
  62448=>"00000010",
  62449=>"11111101",
  62450=>"00000000",
  62451=>"11111110",
  62452=>"00000010",
  62453=>"11111110",
  62454=>"00000011",
  62455=>"11111101",
  62456=>"00000000",
  62457=>"00000000",
  62458=>"11111101",
  62459=>"00000010",
  62460=>"11111110",
  62461=>"00000000",
  62462=>"00000000",
  62463=>"00000000",
  62464=>"00000000",
  62465=>"00000001",
  62466=>"00000001",
  62467=>"11111111",
  62468=>"00000100",
  62469=>"00000001",
  62470=>"00000001",
  62471=>"11111100",
  62472=>"00000000",
  62473=>"00000010",
  62474=>"11111101",
  62475=>"00000000",
  62476=>"11111101",
  62477=>"11111110",
  62478=>"00000001",
  62479=>"00000011",
  62480=>"11111101",
  62481=>"11111101",
  62482=>"11111101",
  62483=>"00000001",
  62484=>"00000000",
  62485=>"11111101",
  62486=>"00000011",
  62487=>"11111101",
  62488=>"11111111",
  62489=>"00000011",
  62490=>"00000011",
  62491=>"00000000",
  62492=>"00000001",
  62493=>"11111111",
  62494=>"00000001",
  62495=>"00000010",
  62496=>"11111111",
  62497=>"11111100",
  62498=>"00000001",
  62499=>"00000010",
  62500=>"00000010",
  62501=>"00000000",
  62502=>"00000010",
  62503=>"11111110",
  62504=>"11111101",
  62505=>"11111101",
  62506=>"00000011",
  62507=>"11111110",
  62508=>"00000000",
  62509=>"00000000",
  62510=>"11111110",
  62511=>"00000001",
  62512=>"00000010",
  62513=>"11111111",
  62514=>"11111100",
  62515=>"11111111",
  62516=>"11111111",
  62517=>"00000101",
  62518=>"11111111",
  62519=>"00000000",
  62520=>"00000011",
  62521=>"11111101",
  62522=>"11111111",
  62523=>"00000000",
  62524=>"00000000",
  62525=>"00000000",
  62526=>"11111101",
  62527=>"00000110",
  62528=>"11111111",
  62529=>"00000001",
  62530=>"00000001",
  62531=>"11111111",
  62532=>"00000000",
  62533=>"00000000",
  62534=>"11111101",
  62535=>"00000001",
  62536=>"00000000",
  62537=>"00000001",
  62538=>"00000011",
  62539=>"00000011",
  62540=>"11111111",
  62541=>"11111101",
  62542=>"11111111",
  62543=>"11111101",
  62544=>"11111110",
  62545=>"00000000",
  62546=>"00000000",
  62547=>"00000000",
  62548=>"00000000",
  62549=>"00000000",
  62550=>"11111101",
  62551=>"00000000",
  62552=>"00000001",
  62553=>"00000001",
  62554=>"11111111",
  62555=>"11111110",
  62556=>"11111110",
  62557=>"11111111",
  62558=>"11111111",
  62559=>"00000001",
  62560=>"11111101",
  62561=>"00000101",
  62562=>"00000100",
  62563=>"00000011",
  62564=>"00000000",
  62565=>"00000001",
  62566=>"11111111",
  62567=>"11111110",
  62568=>"11111111",
  62569=>"11111100",
  62570=>"11111111",
  62571=>"00000000",
  62572=>"00000000",
  62573=>"00000001",
  62574=>"00000001",
  62575=>"00000001",
  62576=>"11111110",
  62577=>"11111110",
  62578=>"11111110",
  62579=>"00000010",
  62580=>"00000010",
  62581=>"00000010",
  62582=>"11111100",
  62583=>"00000000",
  62584=>"11111101",
  62585=>"11111101",
  62586=>"00000011",
  62587=>"11111111",
  62588=>"11111111",
  62589=>"11111110",
  62590=>"11111101",
  62591=>"00000010",
  62592=>"11111100",
  62593=>"11111101",
  62594=>"11111111",
  62595=>"00000000",
  62596=>"00000010",
  62597=>"11111111",
  62598=>"00000010",
  62599=>"00000100",
  62600=>"00000000",
  62601=>"11111101",
  62602=>"11111111",
  62603=>"00000110",
  62604=>"00000010",
  62605=>"11111101",
  62606=>"00000011",
  62607=>"00000001",
  62608=>"00000011",
  62609=>"00000100",
  62610=>"00000000",
  62611=>"11111110",
  62612=>"11111111",
  62613=>"00000001",
  62614=>"00000100",
  62615=>"00000010",
  62616=>"00000001",
  62617=>"00000001",
  62618=>"11111101",
  62619=>"11111110",
  62620=>"00000010",
  62621=>"11111110",
  62622=>"00000010",
  62623=>"00000010",
  62624=>"00000000",
  62625=>"11111101",
  62626=>"11111111",
  62627=>"00000010",
  62628=>"00000000",
  62629=>"00000000",
  62630=>"11111111",
  62631=>"11111110",
  62632=>"11111111",
  62633=>"00000010",
  62634=>"11111101",
  62635=>"11111110",
  62636=>"00000001",
  62637=>"00000010",
  62638=>"11111101",
  62639=>"11111101",
  62640=>"00000001",
  62641=>"00000000",
  62642=>"11111111",
  62643=>"11111111",
  62644=>"00000000",
  62645=>"11111101",
  62646=>"11111111",
  62647=>"11111101",
  62648=>"11111100",
  62649=>"11111111",
  62650=>"11111111",
  62651=>"00000011",
  62652=>"00000000",
  62653=>"11111110",
  62654=>"00000010",
  62655=>"00000010",
  62656=>"11111101",
  62657=>"00000000",
  62658=>"00000000",
  62659=>"00000100",
  62660=>"00000011",
  62661=>"00000110",
  62662=>"00000010",
  62663=>"00000000",
  62664=>"00000000",
  62665=>"00000101",
  62666=>"00000001",
  62667=>"11111111",
  62668=>"00000010",
  62669=>"00000010",
  62670=>"11111111",
  62671=>"11111110",
  62672=>"11111111",
  62673=>"00000001",
  62674=>"00000010",
  62675=>"00000001",
  62676=>"00000010",
  62677=>"00000001",
  62678=>"00000100",
  62679=>"00000010",
  62680=>"11111110",
  62681=>"11111111",
  62682=>"00000010",
  62683=>"00000011",
  62684=>"00000000",
  62685=>"00000001",
  62686=>"00000001",
  62687=>"00000000",
  62688=>"00000000",
  62689=>"11111110",
  62690=>"11111111",
  62691=>"11111111",
  62692=>"00000010",
  62693=>"11111110",
  62694=>"00000011",
  62695=>"00000000",
  62696=>"00000000",
  62697=>"00000001",
  62698=>"00000011",
  62699=>"00000010",
  62700=>"00000000",
  62701=>"00000010",
  62702=>"11111110",
  62703=>"00000010",
  62704=>"11111100",
  62705=>"11111100",
  62706=>"00000001",
  62707=>"00000100",
  62708=>"11111101",
  62709=>"00000000",
  62710=>"00000010",
  62711=>"11111111",
  62712=>"11111110",
  62713=>"00000010",
  62714=>"11111101",
  62715=>"00000000",
  62716=>"00000100",
  62717=>"00000011",
  62718=>"11111110",
  62719=>"11111111",
  62720=>"00000011",
  62721=>"00000000",
  62722=>"00000000",
  62723=>"00000010",
  62724=>"00000010",
  62725=>"00000001",
  62726=>"00000000",
  62727=>"00000110",
  62728=>"11111111",
  62729=>"11111100",
  62730=>"00000011",
  62731=>"00000011",
  62732=>"00000000",
  62733=>"11111101",
  62734=>"00000010",
  62735=>"11111111",
  62736=>"11111111",
  62737=>"00000001",
  62738=>"11111111",
  62739=>"11111111",
  62740=>"11111111",
  62741=>"11111111",
  62742=>"00000000",
  62743=>"00000000",
  62744=>"11111110",
  62745=>"00000001",
  62746=>"00000011",
  62747=>"11111110",
  62748=>"00000011",
  62749=>"11111110",
  62750=>"00000001",
  62751=>"11111111",
  62752=>"00000000",
  62753=>"11111110",
  62754=>"11111111",
  62755=>"00000000",
  62756=>"11111101",
  62757=>"00000100",
  62758=>"00000000",
  62759=>"00000000",
  62760=>"00000100",
  62761=>"11111111",
  62762=>"11111111",
  62763=>"00000000",
  62764=>"11111110",
  62765=>"11111110",
  62766=>"00000010",
  62767=>"00000000",
  62768=>"00000010",
  62769=>"11111110",
  62770=>"00000001",
  62771=>"11111101",
  62772=>"00000010",
  62773=>"00000000",
  62774=>"00000000",
  62775=>"11111101",
  62776=>"11111101",
  62777=>"11111110",
  62778=>"11111110",
  62779=>"00000000",
  62780=>"11111111",
  62781=>"00000000",
  62782=>"00000111",
  62783=>"11111110",
  62784=>"11111110",
  62785=>"00000000",
  62786=>"00000100",
  62787=>"11111110",
  62788=>"11111110",
  62789=>"00000010",
  62790=>"00000000",
  62791=>"11111101",
  62792=>"11111101",
  62793=>"00000101",
  62794=>"00000001",
  62795=>"11111111",
  62796=>"11111110",
  62797=>"00000000",
  62798=>"00000010",
  62799=>"00000010",
  62800=>"00000001",
  62801=>"00000001",
  62802=>"00000100",
  62803=>"11111111",
  62804=>"00000100",
  62805=>"00000000",
  62806=>"00000000",
  62807=>"00000011",
  62808=>"00000011",
  62809=>"00000010",
  62810=>"11111111",
  62811=>"11111110",
  62812=>"00000001",
  62813=>"00000000",
  62814=>"11111111",
  62815=>"00000000",
  62816=>"00000100",
  62817=>"00000000",
  62818=>"00000001",
  62819=>"11111101",
  62820=>"00000001",
  62821=>"11111111",
  62822=>"11111110",
  62823=>"00000001",
  62824=>"00000000",
  62825=>"00000010",
  62826=>"11111110",
  62827=>"11111110",
  62828=>"00000010",
  62829=>"11111110",
  62830=>"11111101",
  62831=>"11111110",
  62832=>"00000001",
  62833=>"00000011",
  62834=>"00000100",
  62835=>"00000010",
  62836=>"11111110",
  62837=>"11111110",
  62838=>"00000001",
  62839=>"11111111",
  62840=>"11111101",
  62841=>"11111111",
  62842=>"11111110",
  62843=>"00000000",
  62844=>"11111111",
  62845=>"00000001",
  62846=>"11111101",
  62847=>"00000001",
  62848=>"11111111",
  62849=>"00000010",
  62850=>"00000000",
  62851=>"00000010",
  62852=>"11111110",
  62853=>"00000001",
  62854=>"00000001",
  62855=>"00000000",
  62856=>"00000010",
  62857=>"00000010",
  62858=>"00000010",
  62859=>"11111111",
  62860=>"00000010",
  62861=>"00000011",
  62862=>"00000001",
  62863=>"00000010",
  62864=>"00000010",
  62865=>"00000000",
  62866=>"00000000",
  62867=>"11111101",
  62868=>"00000010",
  62869=>"00000101",
  62870=>"11111111",
  62871=>"00000011",
  62872=>"11111111",
  62873=>"00000010",
  62874=>"11111111",
  62875=>"00000001",
  62876=>"11111110",
  62877=>"11111111",
  62878=>"11111111",
  62879=>"00000000",
  62880=>"11111111",
  62881=>"00000001",
  62882=>"00000000",
  62883=>"00000000",
  62884=>"00000001",
  62885=>"11111110",
  62886=>"11111100",
  62887=>"11111111",
  62888=>"11111110",
  62889=>"00000001",
  62890=>"00000001",
  62891=>"11111110",
  62892=>"00000001",
  62893=>"00000010",
  62894=>"00000011",
  62895=>"11111111",
  62896=>"11111110",
  62897=>"11111101",
  62898=>"00000010",
  62899=>"11111101",
  62900=>"11111110",
  62901=>"11111110",
  62902=>"00000001",
  62903=>"11111110",
  62904=>"00000100",
  62905=>"11111110",
  62906=>"00000011",
  62907=>"11111111",
  62908=>"00000001",
  62909=>"11111101",
  62910=>"00000000",
  62911=>"11111101",
  62912=>"00000001",
  62913=>"00000010",
  62914=>"00000000",
  62915=>"00000001",
  62916=>"11111111",
  62917=>"00000010",
  62918=>"00000010",
  62919=>"00000000",
  62920=>"11111111",
  62921=>"00000010",
  62922=>"11111111",
  62923=>"11111110",
  62924=>"00000001",
  62925=>"11111110",
  62926=>"00000010",
  62927=>"00000010",
  62928=>"11111111",
  62929=>"00000000",
  62930=>"00000011",
  62931=>"11111111",
  62932=>"00000011",
  62933=>"00000000",
  62934=>"00000010",
  62935=>"00000010",
  62936=>"11111101",
  62937=>"00000000",
  62938=>"00000011",
  62939=>"00000011",
  62940=>"00000011",
  62941=>"11111111",
  62942=>"00000010",
  62943=>"00000010",
  62944=>"00000000",
  62945=>"11111110",
  62946=>"11111110",
  62947=>"00000001",
  62948=>"11111110",
  62949=>"11111101",
  62950=>"00000011",
  62951=>"00000000",
  62952=>"00000101",
  62953=>"11111111",
  62954=>"00000010",
  62955=>"11111111",
  62956=>"00000001",
  62957=>"00000010",
  62958=>"11111111",
  62959=>"11111100",
  62960=>"11111111",
  62961=>"11111100",
  62962=>"00000000",
  62963=>"11111110",
  62964=>"00000010",
  62965=>"11111111",
  62966=>"11111100",
  62967=>"00000101",
  62968=>"11111110",
  62969=>"11111101",
  62970=>"00000000",
  62971=>"11111110",
  62972=>"11111111",
  62973=>"11111110",
  62974=>"00000010",
  62975=>"00000010",
  62976=>"00000010",
  62977=>"00000010",
  62978=>"00000001",
  62979=>"00000011",
  62980=>"11111101",
  62981=>"00000010",
  62982=>"11111111",
  62983=>"00000100",
  62984=>"11111101",
  62985=>"11111101",
  62986=>"00000000",
  62987=>"00000000",
  62988=>"00000011",
  62989=>"00000001",
  62990=>"00000011",
  62991=>"11111100",
  62992=>"00000100",
  62993=>"11111111",
  62994=>"00000001",
  62995=>"00000011",
  62996=>"00000001",
  62997=>"11111111",
  62998=>"00000000",
  62999=>"11111101",
  63000=>"00000001",
  63001=>"11111111",
  63002=>"11111110",
  63003=>"00000011",
  63004=>"00000000",
  63005=>"00000101",
  63006=>"00000010",
  63007=>"11111110",
  63008=>"00000010",
  63009=>"00000000",
  63010=>"11111111",
  63011=>"00000100",
  63012=>"11111101",
  63013=>"00000100",
  63014=>"00000011",
  63015=>"00000010",
  63016=>"11111101",
  63017=>"00000001",
  63018=>"00000010",
  63019=>"00000010",
  63020=>"11111110",
  63021=>"00000000",
  63022=>"00000010",
  63023=>"11111111",
  63024=>"00000110",
  63025=>"11111101",
  63026=>"11111110",
  63027=>"00000000",
  63028=>"11111111",
  63029=>"00000001",
  63030=>"00000001",
  63031=>"00000011",
  63032=>"00000011",
  63033=>"00000001",
  63034=>"00000001",
  63035=>"00000010",
  63036=>"00000001",
  63037=>"11111111",
  63038=>"11111111",
  63039=>"00000001",
  63040=>"11111100",
  63041=>"11111111",
  63042=>"11111111",
  63043=>"11111110",
  63044=>"11111110",
  63045=>"00000000",
  63046=>"11111101",
  63047=>"11111110",
  63048=>"11111110",
  63049=>"11111110",
  63050=>"11111110",
  63051=>"11111110",
  63052=>"00000001",
  63053=>"11111101",
  63054=>"00000011",
  63055=>"00000000",
  63056=>"11111110",
  63057=>"00000000",
  63058=>"11111110",
  63059=>"00000010",
  63060=>"00000001",
  63061=>"00000001",
  63062=>"00000001",
  63063=>"00000000",
  63064=>"00000011",
  63065=>"11111101",
  63066=>"11111101",
  63067=>"11111111",
  63068=>"00000000",
  63069=>"11111110",
  63070=>"11111101",
  63071=>"00000001",
  63072=>"00000001",
  63073=>"00000001",
  63074=>"00000010",
  63075=>"00000101",
  63076=>"11111111",
  63077=>"11111110",
  63078=>"11111110",
  63079=>"00000001",
  63080=>"00000000",
  63081=>"00000000",
  63082=>"00000010",
  63083=>"11111110",
  63084=>"00000000",
  63085=>"00000000",
  63086=>"00000001",
  63087=>"00000110",
  63088=>"11111110",
  63089=>"00000010",
  63090=>"00000010",
  63091=>"00000001",
  63092=>"00000010",
  63093=>"00000010",
  63094=>"11111111",
  63095=>"00000001",
  63096=>"11111110",
  63097=>"11111111",
  63098=>"00000001",
  63099=>"00000010",
  63100=>"00000000",
  63101=>"11111110",
  63102=>"00000010",
  63103=>"11111110",
  63104=>"00000010",
  63105=>"00000001",
  63106=>"11111100",
  63107=>"00000000",
  63108=>"11111111",
  63109=>"11111110",
  63110=>"00000001",
  63111=>"11111110",
  63112=>"00000010",
  63113=>"00000000",
  63114=>"11111111",
  63115=>"00000000",
  63116=>"11111110",
  63117=>"11111110",
  63118=>"11111110",
  63119=>"11111110",
  63120=>"00000010",
  63121=>"00000001",
  63122=>"11111111",
  63123=>"00000001",
  63124=>"00000010",
  63125=>"00000000",
  63126=>"11111101",
  63127=>"00000100",
  63128=>"11111101",
  63129=>"00000111",
  63130=>"00000000",
  63131=>"00000001",
  63132=>"00000101",
  63133=>"11111101",
  63134=>"00000001",
  63135=>"00000011",
  63136=>"00000001",
  63137=>"00000010",
  63138=>"11111110",
  63139=>"11111111",
  63140=>"11111110",
  63141=>"00000001",
  63142=>"00000001",
  63143=>"00000000",
  63144=>"11111101",
  63145=>"00000000",
  63146=>"00000010",
  63147=>"00000000",
  63148=>"11111110",
  63149=>"11111101",
  63150=>"00000010",
  63151=>"11111111",
  63152=>"00000001",
  63153=>"11111110",
  63154=>"00000011",
  63155=>"00000001",
  63156=>"00000010",
  63157=>"11111101",
  63158=>"00000000",
  63159=>"00000101",
  63160=>"00000010",
  63161=>"11111101",
  63162=>"00000001",
  63163=>"00000010",
  63164=>"11111111",
  63165=>"11111111",
  63166=>"00000000",
  63167=>"11111101",
  63168=>"00000000",
  63169=>"00000001",
  63170=>"00000011",
  63171=>"00000001",
  63172=>"11111111",
  63173=>"11111111",
  63174=>"00000010",
  63175=>"00000000",
  63176=>"00000010",
  63177=>"00000001",
  63178=>"11111110",
  63179=>"11111110",
  63180=>"00000001",
  63181=>"11111101",
  63182=>"00000000",
  63183=>"00000000",
  63184=>"11111111",
  63185=>"00000000",
  63186=>"11111110",
  63187=>"11111110",
  63188=>"00000001",
  63189=>"00000011",
  63190=>"11111110",
  63191=>"00000000",
  63192=>"00000010",
  63193=>"00000010",
  63194=>"11111110",
  63195=>"00000101",
  63196=>"11111101",
  63197=>"00000001",
  63198=>"11111110",
  63199=>"00000100",
  63200=>"11111110",
  63201=>"00000100",
  63202=>"11111111",
  63203=>"11111111",
  63204=>"11111111",
  63205=>"00000000",
  63206=>"11111110",
  63207=>"11111110",
  63208=>"11111111",
  63209=>"11111111",
  63210=>"00000010",
  63211=>"11111110",
  63212=>"00000000",
  63213=>"11111100",
  63214=>"00000100",
  63215=>"00000010",
  63216=>"00000000",
  63217=>"11111101",
  63218=>"11111101",
  63219=>"11111111",
  63220=>"00000001",
  63221=>"11111101",
  63222=>"00000010",
  63223=>"00000000",
  63224=>"11111101",
  63225=>"00000010",
  63226=>"11111111",
  63227=>"00000001",
  63228=>"00000000",
  63229=>"11111111",
  63230=>"11111111",
  63231=>"00000001",
  63232=>"11111111",
  63233=>"00000011",
  63234=>"11111110",
  63235=>"00000100",
  63236=>"11111110",
  63237=>"00000010",
  63238=>"00000011",
  63239=>"11111111",
  63240=>"00000000",
  63241=>"00000001",
  63242=>"00000010",
  63243=>"11111100",
  63244=>"11111111",
  63245=>"00000000",
  63246=>"00000010",
  63247=>"00000010",
  63248=>"11111111",
  63249=>"00000011",
  63250=>"11111110",
  63251=>"11111110",
  63252=>"11111110",
  63253=>"00000001",
  63254=>"00000000",
  63255=>"00000001",
  63256=>"11111111",
  63257=>"00000100",
  63258=>"00000100",
  63259=>"11111111",
  63260=>"11111111",
  63261=>"11111111",
  63262=>"11111101",
  63263=>"00000010",
  63264=>"00000101",
  63265=>"11111111",
  63266=>"11111110",
  63267=>"11111110",
  63268=>"00000100",
  63269=>"11111100",
  63270=>"00000000",
  63271=>"00000000",
  63272=>"11111111",
  63273=>"11111110",
  63274=>"00000001",
  63275=>"00000000",
  63276=>"00000001",
  63277=>"00000000",
  63278=>"00000000",
  63279=>"11111110",
  63280=>"00000000",
  63281=>"00000011",
  63282=>"11111111",
  63283=>"00000010",
  63284=>"11111111",
  63285=>"11111100",
  63286=>"11111111",
  63287=>"11111101",
  63288=>"11111100",
  63289=>"11111111",
  63290=>"11111110",
  63291=>"11111111",
  63292=>"00000000",
  63293=>"11111111",
  63294=>"11111101",
  63295=>"11111111",
  63296=>"00000100",
  63297=>"11111110",
  63298=>"00000000",
  63299=>"00000011",
  63300=>"11111111",
  63301=>"00000001",
  63302=>"11111110",
  63303=>"00000000",
  63304=>"00000001",
  63305=>"11111101",
  63306=>"11111110",
  63307=>"00000000",
  63308=>"00000001",
  63309=>"00000010",
  63310=>"00000111",
  63311=>"11111111",
  63312=>"11111111",
  63313=>"11111101",
  63314=>"11111111",
  63315=>"00000010",
  63316=>"11111101",
  63317=>"00000001",
  63318=>"00000010",
  63319=>"11111101",
  63320=>"00000000",
  63321=>"11111110",
  63322=>"00000010",
  63323=>"11111100",
  63324=>"00000001",
  63325=>"00000011",
  63326=>"00000000",
  63327=>"00000011",
  63328=>"11111111",
  63329=>"00000010",
  63330=>"11111110",
  63331=>"11111111",
  63332=>"11111110",
  63333=>"11111110",
  63334=>"11111100",
  63335=>"00000110",
  63336=>"11111111",
  63337=>"11111111",
  63338=>"00000000",
  63339=>"11111110",
  63340=>"11111101",
  63341=>"11111110",
  63342=>"11111111",
  63343=>"11111111",
  63344=>"11111110",
  63345=>"00000011",
  63346=>"11111110",
  63347=>"11111111",
  63348=>"11111101",
  63349=>"00000111",
  63350=>"00000000",
  63351=>"00000000",
  63352=>"11111111",
  63353=>"00000010",
  63354=>"00000100",
  63355=>"00000010",
  63356=>"00000000",
  63357=>"11111110",
  63358=>"11111110",
  63359=>"00000100",
  63360=>"11111110",
  63361=>"11111110",
  63362=>"11111101",
  63363=>"11111111",
  63364=>"00000010",
  63365=>"11111111",
  63366=>"11111111",
  63367=>"11111101",
  63368=>"00000001",
  63369=>"00000011",
  63370=>"11111111",
  63371=>"00000000",
  63372=>"00000010",
  63373=>"00000010",
  63374=>"11111100",
  63375=>"11111110",
  63376=>"11111111",
  63377=>"11111110",
  63378=>"00000000",
  63379=>"11111111",
  63380=>"11111111",
  63381=>"00000001",
  63382=>"11111101",
  63383=>"11111110",
  63384=>"00000110",
  63385=>"00000100",
  63386=>"11111110",
  63387=>"00000000",
  63388=>"11111100",
  63389=>"00000001",
  63390=>"00000001",
  63391=>"11111101",
  63392=>"11111101",
  63393=>"00000000",
  63394=>"11111111",
  63395=>"00000010",
  63396=>"00000000",
  63397=>"00000001",
  63398=>"11111101",
  63399=>"11111111",
  63400=>"00000001",
  63401=>"11111111",
  63402=>"00000100",
  63403=>"00000000",
  63404=>"11111110",
  63405=>"00000100",
  63406=>"00000010",
  63407=>"00000000",
  63408=>"11111101",
  63409=>"11111111",
  63410=>"00000011",
  63411=>"00000000",
  63412=>"11111101",
  63413=>"11111101",
  63414=>"00000000",
  63415=>"00000111",
  63416=>"11111110",
  63417=>"00000011",
  63418=>"00000001",
  63419=>"11111100",
  63420=>"11111111",
  63421=>"00000011",
  63422=>"11111110",
  63423=>"11111111",
  63424=>"11111101",
  63425=>"00000010",
  63426=>"11111111",
  63427=>"00000011",
  63428=>"00000000",
  63429=>"11111111",
  63430=>"11111110",
  63431=>"11111110",
  63432=>"00000001",
  63433=>"11111101",
  63434=>"00000010",
  63435=>"00000010",
  63436=>"00000011",
  63437=>"00000001",
  63438=>"11111111",
  63439=>"11111101",
  63440=>"00000011",
  63441=>"11111111",
  63442=>"11111110",
  63443=>"00000010",
  63444=>"00000000",
  63445=>"00000011",
  63446=>"00000101",
  63447=>"00000010",
  63448=>"00000001",
  63449=>"00000000",
  63450=>"11111111",
  63451=>"00000100",
  63452=>"11111110",
  63453=>"00000001",
  63454=>"11111110",
  63455=>"00000000",
  63456=>"11111111",
  63457=>"00000000",
  63458=>"00000000",
  63459=>"00000010",
  63460=>"00000010",
  63461=>"00000000",
  63462=>"11111101",
  63463=>"00000010",
  63464=>"00000001",
  63465=>"00000010",
  63466=>"00000011",
  63467=>"00000011",
  63468=>"11111111",
  63469=>"11111101",
  63470=>"11111111",
  63471=>"11111110",
  63472=>"00000010",
  63473=>"00000001",
  63474=>"11111111",
  63475=>"11111111",
  63476=>"11111111",
  63477=>"11111110",
  63478=>"00000010",
  63479=>"11111100",
  63480=>"00000001",
  63481=>"00000000",
  63482=>"00000011",
  63483=>"00000100",
  63484=>"00000010",
  63485=>"11111100",
  63486=>"11111111",
  63487=>"11111110",
  63488=>"00000010",
  63489=>"00000001",
  63490=>"11111110",
  63491=>"00000000",
  63492=>"11111110",
  63493=>"11111111",
  63494=>"00000001",
  63495=>"11111110",
  63496=>"11111101",
  63497=>"00000110",
  63498=>"00000001",
  63499=>"00000010",
  63500=>"00000001",
  63501=>"00000000",
  63502=>"00000010",
  63503=>"00000101",
  63504=>"11111110",
  63505=>"11111101",
  63506=>"11111101",
  63507=>"00000011",
  63508=>"11111110",
  63509=>"00000000",
  63510=>"00000000",
  63511=>"00000110",
  63512=>"11111101",
  63513=>"00000000",
  63514=>"00000000",
  63515=>"11111011",
  63516=>"00000001",
  63517=>"11111110",
  63518=>"11111110",
  63519=>"11111101",
  63520=>"11111101",
  63521=>"00000000",
  63522=>"00000010",
  63523=>"00000001",
  63524=>"00000001",
  63525=>"00000011",
  63526=>"00000101",
  63527=>"00000100",
  63528=>"00000100",
  63529=>"00000010",
  63530=>"11111110",
  63531=>"11111100",
  63532=>"00000010",
  63533=>"00000000",
  63534=>"00000100",
  63535=>"11111110",
  63536=>"11111111",
  63537=>"00000111",
  63538=>"00000001",
  63539=>"00000011",
  63540=>"00000010",
  63541=>"00000000",
  63542=>"00000001",
  63543=>"00000000",
  63544=>"11111110",
  63545=>"11111111",
  63546=>"00000011",
  63547=>"00000010",
  63548=>"00000110",
  63549=>"11111101",
  63550=>"00000010",
  63551=>"00000001",
  63552=>"00000000",
  63553=>"00000010",
  63554=>"00000000",
  63555=>"00000001",
  63556=>"00000000",
  63557=>"11111110",
  63558=>"11111110",
  63559=>"11111110",
  63560=>"00000011",
  63561=>"00000100",
  63562=>"00000000",
  63563=>"00000101",
  63564=>"11111101",
  63565=>"11111111",
  63566=>"11111101",
  63567=>"00000000",
  63568=>"11111110",
  63569=>"00000110",
  63570=>"11111100",
  63571=>"11111100",
  63572=>"00000011",
  63573=>"00000001",
  63574=>"00000001",
  63575=>"00000001",
  63576=>"11111110",
  63577=>"00000000",
  63578=>"00000000",
  63579=>"11111101",
  63580=>"00000001",
  63581=>"11111111",
  63582=>"00000010",
  63583=>"11111101",
  63584=>"11111101",
  63585=>"00000010",
  63586=>"11111111",
  63587=>"00000000",
  63588=>"11111101",
  63589=>"00000011",
  63590=>"11111101",
  63591=>"00000110",
  63592=>"00000000",
  63593=>"11111111",
  63594=>"00000001",
  63595=>"00000010",
  63596=>"00000000",
  63597=>"11111100",
  63598=>"11111111",
  63599=>"11111111",
  63600=>"00000110",
  63601=>"11111111",
  63602=>"11111110",
  63603=>"11111111",
  63604=>"11111111",
  63605=>"11111111",
  63606=>"00000000",
  63607=>"00000010",
  63608=>"00000111",
  63609=>"00000101",
  63610=>"00000000",
  63611=>"11111111",
  63612=>"00000011",
  63613=>"00000000",
  63614=>"00000000",
  63615=>"11111111",
  63616=>"00000000",
  63617=>"11111110",
  63618=>"11111101",
  63619=>"11111110",
  63620=>"11111110",
  63621=>"11111101",
  63622=>"11111111",
  63623=>"00000011",
  63624=>"00000010",
  63625=>"11111111",
  63626=>"11111111",
  63627=>"11111111",
  63628=>"11111110",
  63629=>"00000010",
  63630=>"00000010",
  63631=>"11111101",
  63632=>"11111110",
  63633=>"11111100",
  63634=>"00000000",
  63635=>"11111111",
  63636=>"11111110",
  63637=>"00000101",
  63638=>"11111100",
  63639=>"00000110",
  63640=>"00000000",
  63641=>"00000011",
  63642=>"11111101",
  63643=>"11111101",
  63644=>"11111111",
  63645=>"00000011",
  63646=>"00000001",
  63647=>"00000000",
  63648=>"11111101",
  63649=>"00000001",
  63650=>"00000100",
  63651=>"11111110",
  63652=>"00000010",
  63653=>"00000101",
  63654=>"11111111",
  63655=>"00000010",
  63656=>"00000011",
  63657=>"00000010",
  63658=>"11111110",
  63659=>"11111101",
  63660=>"11111110",
  63661=>"00000011",
  63662=>"11111111",
  63663=>"00000001",
  63664=>"00000010",
  63665=>"00000110",
  63666=>"11111101",
  63667=>"11111110",
  63668=>"00000001",
  63669=>"11111111",
  63670=>"11111101",
  63671=>"00000010",
  63672=>"00000101",
  63673=>"11111111",
  63674=>"00000100",
  63675=>"11111101",
  63676=>"11111111",
  63677=>"00000001",
  63678=>"00000001",
  63679=>"11111111",
  63680=>"00000000",
  63681=>"00000000",
  63682=>"00000100",
  63683=>"11111110",
  63684=>"00000000",
  63685=>"00000001",
  63686=>"11111100",
  63687=>"11111111",
  63688=>"00000000",
  63689=>"11111011",
  63690=>"00000000",
  63691=>"00000101",
  63692=>"11111100",
  63693=>"00000001",
  63694=>"11111111",
  63695=>"11111100",
  63696=>"00000000",
  63697=>"11111110",
  63698=>"11111111",
  63699=>"11111111",
  63700=>"00000010",
  63701=>"00000001",
  63702=>"11111100",
  63703=>"00000000",
  63704=>"00000111",
  63705=>"11111110",
  63706=>"00000110",
  63707=>"11111110",
  63708=>"00000001",
  63709=>"00000010",
  63710=>"00000010",
  63711=>"11111101",
  63712=>"00000000",
  63713=>"00000010",
  63714=>"11111111",
  63715=>"00000010",
  63716=>"00000001",
  63717=>"00000000",
  63718=>"00000010",
  63719=>"00000010",
  63720=>"00000001",
  63721=>"00000010",
  63722=>"00000001",
  63723=>"00000001",
  63724=>"11111101",
  63725=>"11111110",
  63726=>"00000010",
  63727=>"00000001",
  63728=>"00000001",
  63729=>"11111100",
  63730=>"11111100",
  63731=>"11111111",
  63732=>"11111111",
  63733=>"11111111",
  63734=>"11111100",
  63735=>"00000000",
  63736=>"11111101",
  63737=>"00000100",
  63738=>"00000010",
  63739=>"00000010",
  63740=>"00000001",
  63741=>"11111111",
  63742=>"00000100",
  63743=>"00000010",
  63744=>"11111110",
  63745=>"00000000",
  63746=>"11111110",
  63747=>"11111111",
  63748=>"00000010",
  63749=>"11111110",
  63750=>"11111111",
  63751=>"00000000",
  63752=>"00000010",
  63753=>"11111101",
  63754=>"11111111",
  63755=>"11111100",
  63756=>"11111110",
  63757=>"11111111",
  63758=>"00000001",
  63759=>"11111100",
  63760=>"11111100",
  63761=>"00000000",
  63762=>"00000000",
  63763=>"00000011",
  63764=>"00000100",
  63765=>"00000000",
  63766=>"11111100",
  63767=>"00000011",
  63768=>"11111111",
  63769=>"00000001",
  63770=>"00000010",
  63771=>"11111110",
  63772=>"11111101",
  63773=>"00000011",
  63774=>"11111101",
  63775=>"11111101",
  63776=>"11111110",
  63777=>"11111111",
  63778=>"00000000",
  63779=>"11111101",
  63780=>"00000100",
  63781=>"00001000",
  63782=>"00000001",
  63783=>"00000010",
  63784=>"11111110",
  63785=>"11111101",
  63786=>"00000001",
  63787=>"11111111",
  63788=>"11111111",
  63789=>"00000000",
  63790=>"00000011",
  63791=>"00000000",
  63792=>"11111111",
  63793=>"11111101",
  63794=>"11111110",
  63795=>"11111100",
  63796=>"00000001",
  63797=>"11111101",
  63798=>"11111101",
  63799=>"11111101",
  63800=>"00000010",
  63801=>"00000101",
  63802=>"11111110",
  63803=>"00000011",
  63804=>"00000000",
  63805=>"11111110",
  63806=>"00000010",
  63807=>"00000001",
  63808=>"00000001",
  63809=>"00000000",
  63810=>"00000001",
  63811=>"00000010",
  63812=>"11111111",
  63813=>"11111111",
  63814=>"11111111",
  63815=>"00000001",
  63816=>"11111111",
  63817=>"11111110",
  63818=>"11111110",
  63819=>"00000001",
  63820=>"00000001",
  63821=>"00000011",
  63822=>"11111101",
  63823=>"00000010",
  63824=>"11111110",
  63825=>"11111111",
  63826=>"00000010",
  63827=>"00000011",
  63828=>"11111111",
  63829=>"11111101",
  63830=>"00000001",
  63831=>"00000000",
  63832=>"00000001",
  63833=>"00000000",
  63834=>"11111100",
  63835=>"11111111",
  63836=>"00000010",
  63837=>"11111101",
  63838=>"00000100",
  63839=>"00000001",
  63840=>"00000001",
  63841=>"00000011",
  63842=>"11111101",
  63843=>"00000011",
  63844=>"00000010",
  63845=>"00000000",
  63846=>"00000000",
  63847=>"11111111",
  63848=>"00000001",
  63849=>"00000001",
  63850=>"00000011",
  63851=>"00000000",
  63852=>"00000011",
  63853=>"11111101",
  63854=>"00000010",
  63855=>"00000010",
  63856=>"00000000",
  63857=>"00000000",
  63858=>"11111110",
  63859=>"00000001",
  63860=>"00000001",
  63861=>"00000101",
  63862=>"00000010",
  63863=>"11111111",
  63864=>"11111111",
  63865=>"11111110",
  63866=>"00000010",
  63867=>"00000000",
  63868=>"11111111",
  63869=>"00000001",
  63870=>"11111110",
  63871=>"00000001",
  63872=>"00000001",
  63873=>"11111110",
  63874=>"00000010",
  63875=>"11111110",
  63876=>"11111101",
  63877=>"11111101",
  63878=>"11111111",
  63879=>"00000010",
  63880=>"11111110",
  63881=>"00000000",
  63882=>"11111111",
  63883=>"00000001",
  63884=>"00000001",
  63885=>"00000010",
  63886=>"00000001",
  63887=>"11111100",
  63888=>"00000000",
  63889=>"00000011",
  63890=>"00000100",
  63891=>"00000010",
  63892=>"00000001",
  63893=>"11111101",
  63894=>"00000000",
  63895=>"11111110",
  63896=>"00000010",
  63897=>"11111110",
  63898=>"00000100",
  63899=>"00000010",
  63900=>"11111111",
  63901=>"11111100",
  63902=>"00000000",
  63903=>"11111110",
  63904=>"11111111",
  63905=>"00000000",
  63906=>"00000010",
  63907=>"00000010",
  63908=>"00000001",
  63909=>"11111111",
  63910=>"11111111",
  63911=>"00000011",
  63912=>"00000010",
  63913=>"11111100",
  63914=>"00000001",
  63915=>"11111111",
  63916=>"11111101",
  63917=>"11111110",
  63918=>"11111110",
  63919=>"11111111",
  63920=>"11111100",
  63921=>"11111111",
  63922=>"00000000",
  63923=>"00000101",
  63924=>"00000001",
  63925=>"00000010",
  63926=>"00000000",
  63927=>"11111101",
  63928=>"11111101",
  63929=>"11111101",
  63930=>"11111101",
  63931=>"11111111",
  63932=>"11111110",
  63933=>"00000011",
  63934=>"00000010",
  63935=>"00000010",
  63936=>"11111110",
  63937=>"00000001",
  63938=>"11111101",
  63939=>"00000100",
  63940=>"11111111",
  63941=>"00000100",
  63942=>"00000011",
  63943=>"11111100",
  63944=>"00000111",
  63945=>"00000001",
  63946=>"00000000",
  63947=>"00000011",
  63948=>"00000000",
  63949=>"11111101",
  63950=>"11111111",
  63951=>"00000010",
  63952=>"00000000",
  63953=>"00000011",
  63954=>"00000001",
  63955=>"11111110",
  63956=>"00000001",
  63957=>"00000110",
  63958=>"11111111",
  63959=>"11111101",
  63960=>"11111101",
  63961=>"00000000",
  63962=>"11111111",
  63963=>"11111111",
  63964=>"00000000",
  63965=>"11111111",
  63966=>"11111101",
  63967=>"00000000",
  63968=>"11111101",
  63969=>"11111111",
  63970=>"00000000",
  63971=>"00000000",
  63972=>"11111111",
  63973=>"00000000",
  63974=>"11111111",
  63975=>"11111110",
  63976=>"00000001",
  63977=>"00000101",
  63978=>"11111110",
  63979=>"00000001",
  63980=>"11111110",
  63981=>"00000000",
  63982=>"00000000",
  63983=>"00000000",
  63984=>"11111111",
  63985=>"11111101",
  63986=>"00000011",
  63987=>"11111111",
  63988=>"00000100",
  63989=>"11111110",
  63990=>"00000000",
  63991=>"00000001",
  63992=>"00000101",
  63993=>"00000001",
  63994=>"11111110",
  63995=>"11111111",
  63996=>"11111110",
  63997=>"11111101",
  63998=>"00000010",
  63999=>"00000001",
  64000=>"00000000",
  64001=>"00000001",
  64002=>"00000000",
  64003=>"00000010",
  64004=>"11111110",
  64005=>"11111110",
  64006=>"11111011",
  64007=>"00000100",
  64008=>"11111110",
  64009=>"11111101",
  64010=>"00000001",
  64011=>"11111101",
  64012=>"00000001",
  64013=>"00000100",
  64014=>"11111111",
  64015=>"11111101",
  64016=>"11111101",
  64017=>"00000000",
  64018=>"11111111",
  64019=>"00000100",
  64020=>"00000001",
  64021=>"00000001",
  64022=>"00000011",
  64023=>"00000001",
  64024=>"11111111",
  64025=>"11111101",
  64026=>"11111110",
  64027=>"00000010",
  64028=>"11111111",
  64029=>"11111101",
  64030=>"11111110",
  64031=>"00000001",
  64032=>"00000001",
  64033=>"00000001",
  64034=>"00000001",
  64035=>"00000010",
  64036=>"00000100",
  64037=>"00000001",
  64038=>"00000100",
  64039=>"11111110",
  64040=>"00000010",
  64041=>"11111110",
  64042=>"11111111",
  64043=>"00000010",
  64044=>"11111110",
  64045=>"00001000",
  64046=>"00000010",
  64047=>"11111110",
  64048=>"11111110",
  64049=>"00000001",
  64050=>"11111110",
  64051=>"11111111",
  64052=>"11111101",
  64053=>"11111110",
  64054=>"11111111",
  64055=>"00000001",
  64056=>"11111111",
  64057=>"11111111",
  64058=>"11111111",
  64059=>"11111111",
  64060=>"00000000",
  64061=>"11111111",
  64062=>"11111111",
  64063=>"11111101",
  64064=>"00000000",
  64065=>"11111111",
  64066=>"00000100",
  64067=>"00000001",
  64068=>"00000101",
  64069=>"00000011",
  64070=>"00000010",
  64071=>"00000000",
  64072=>"11111101",
  64073=>"00000001",
  64074=>"11111110",
  64075=>"11111111",
  64076=>"00000010",
  64077=>"11111110",
  64078=>"00000001",
  64079=>"11111110",
  64080=>"11111111",
  64081=>"11111111",
  64082=>"00000010",
  64083=>"00000000",
  64084=>"11111110",
  64085=>"00000001",
  64086=>"00000000",
  64087=>"11111111",
  64088=>"11111111",
  64089=>"00000001",
  64090=>"00000010",
  64091=>"00000000",
  64092=>"11111111",
  64093=>"11111110",
  64094=>"00000100",
  64095=>"00000011",
  64096=>"11111111",
  64097=>"00000010",
  64098=>"00000000",
  64099=>"11111101",
  64100=>"11111111",
  64101=>"00000101",
  64102=>"00000010",
  64103=>"11111110",
  64104=>"00000000",
  64105=>"00000101",
  64106=>"00000010",
  64107=>"11111110",
  64108=>"00000011",
  64109=>"00000000",
  64110=>"00000000",
  64111=>"11111101",
  64112=>"00000011",
  64113=>"11111110",
  64114=>"00000001",
  64115=>"00000000",
  64116=>"11111111",
  64117=>"11111111",
  64118=>"11111101",
  64119=>"00000000",
  64120=>"11111101",
  64121=>"11111110",
  64122=>"11111111",
  64123=>"11111111",
  64124=>"00000001",
  64125=>"11111101",
  64126=>"11111111",
  64127=>"00000010",
  64128=>"00000010",
  64129=>"00000000",
  64130=>"00000111",
  64131=>"11111100",
  64132=>"11111110",
  64133=>"00000000",
  64134=>"11111111",
  64135=>"00000010",
  64136=>"00000000",
  64137=>"00000000",
  64138=>"11111110",
  64139=>"11111111",
  64140=>"00000001",
  64141=>"00000011",
  64142=>"00000010",
  64143=>"00000001",
  64144=>"11111111",
  64145=>"00000000",
  64146=>"11111011",
  64147=>"00000001",
  64148=>"11111011",
  64149=>"11111101",
  64150=>"11111111",
  64151=>"11111100",
  64152=>"11111110",
  64153=>"11111111",
  64154=>"00000100",
  64155=>"00000001",
  64156=>"00000010",
  64157=>"00000101",
  64158=>"00000000",
  64159=>"11111111",
  64160=>"00000000",
  64161=>"00000011",
  64162=>"00000001",
  64163=>"00000010",
  64164=>"11111111",
  64165=>"11111110",
  64166=>"00000001",
  64167=>"00000011",
  64168=>"11111111",
  64169=>"11111101",
  64170=>"11111111",
  64171=>"11111110",
  64172=>"11111101",
  64173=>"11111110",
  64174=>"11111111",
  64175=>"00000000",
  64176=>"00000010",
  64177=>"11111101",
  64178=>"11111111",
  64179=>"00000010",
  64180=>"00000000",
  64181=>"00000000",
  64182=>"11111101",
  64183=>"00000001",
  64184=>"11111100",
  64185=>"00000000",
  64186=>"00000000",
  64187=>"00000001",
  64188=>"00000000",
  64189=>"00000101",
  64190=>"00000000",
  64191=>"11111101",
  64192=>"11111111",
  64193=>"00000100",
  64194=>"00000111",
  64195=>"00000001",
  64196=>"00000010",
  64197=>"00000100",
  64198=>"00000011",
  64199=>"00000001",
  64200=>"11111100",
  64201=>"00000010",
  64202=>"11111101",
  64203=>"00000000",
  64204=>"11111100",
  64205=>"00000001",
  64206=>"00000100",
  64207=>"11111101",
  64208=>"00000010",
  64209=>"11111101",
  64210=>"00000001",
  64211=>"11111111",
  64212=>"00000000",
  64213=>"11111101",
  64214=>"11111101",
  64215=>"00000001",
  64216=>"00000001",
  64217=>"00000011",
  64218=>"00000000",
  64219=>"11111101",
  64220=>"00000000",
  64221=>"00000000",
  64222=>"11111110",
  64223=>"00000001",
  64224=>"11111110",
  64225=>"11111110",
  64226=>"11111111",
  64227=>"00000010",
  64228=>"11111110",
  64229=>"11111101",
  64230=>"00000100",
  64231=>"11111110",
  64232=>"11111101",
  64233=>"00000011",
  64234=>"00000000",
  64235=>"11111100",
  64236=>"11111111",
  64237=>"11111111",
  64238=>"11111101",
  64239=>"11111100",
  64240=>"00000000",
  64241=>"11111110",
  64242=>"00000000",
  64243=>"11111111",
  64244=>"11111110",
  64245=>"00000001",
  64246=>"00000000",
  64247=>"00000010",
  64248=>"00000100",
  64249=>"11111110",
  64250=>"00000011",
  64251=>"00000000",
  64252=>"00000001",
  64253=>"11111101",
  64254=>"00000000",
  64255=>"00000100",
  64256=>"11111110",
  64257=>"11111110",
  64258=>"00000001",
  64259=>"00000000",
  64260=>"11111110",
  64261=>"00000001",
  64262=>"00000010",
  64263=>"11111111",
  64264=>"00000010",
  64265=>"00000000",
  64266=>"11111111",
  64267=>"11111100",
  64268=>"11111101",
  64269=>"00000000",
  64270=>"11111110",
  64271=>"00000010",
  64272=>"00000011",
  64273=>"00000000",
  64274=>"00000100",
  64275=>"00000100",
  64276=>"11111101",
  64277=>"00000010",
  64278=>"11111111",
  64279=>"11111101",
  64280=>"00000111",
  64281=>"00000010",
  64282=>"00000000",
  64283=>"00000001",
  64284=>"00000000",
  64285=>"11111011",
  64286=>"11111111",
  64287=>"00000011",
  64288=>"11111110",
  64289=>"11111111",
  64290=>"00000000",
  64291=>"11111111",
  64292=>"11111110",
  64293=>"11111111",
  64294=>"00000010",
  64295=>"00000001",
  64296=>"00000111",
  64297=>"11111101",
  64298=>"00000100",
  64299=>"11111110",
  64300=>"00000110",
  64301=>"00000010",
  64302=>"00000010",
  64303=>"00000001",
  64304=>"00000001",
  64305=>"00000001",
  64306=>"11111011",
  64307=>"00000000",
  64308=>"00000001",
  64309=>"11111111",
  64310=>"00000001",
  64311=>"00000001",
  64312=>"00000011",
  64313=>"11111111",
  64314=>"11111110",
  64315=>"11111111",
  64316=>"11111111",
  64317=>"00000010",
  64318=>"11111110",
  64319=>"00000010",
  64320=>"11111100",
  64321=>"00000000",
  64322=>"11111111",
  64323=>"11111100",
  64324=>"00000010",
  64325=>"11111110",
  64326=>"00000001",
  64327=>"00000010",
  64328=>"00000010",
  64329=>"00000010",
  64330=>"11111110",
  64331=>"00000000",
  64332=>"00000000",
  64333=>"11111101",
  64334=>"11111101",
  64335=>"11111110",
  64336=>"00000111",
  64337=>"11111101",
  64338=>"00000010",
  64339=>"00000001",
  64340=>"00000000",
  64341=>"00000001",
  64342=>"00000000",
  64343=>"00000001",
  64344=>"11111100",
  64345=>"00000001",
  64346=>"00000000",
  64347=>"00000000",
  64348=>"11111111",
  64349=>"00000011",
  64350=>"11111101",
  64351=>"11111111",
  64352=>"11111110",
  64353=>"00000000",
  64354=>"00000000",
  64355=>"11111110",
  64356=>"11111111",
  64357=>"11111111",
  64358=>"11111101",
  64359=>"11111110",
  64360=>"11111101",
  64361=>"11111111",
  64362=>"00000000",
  64363=>"00000010",
  64364=>"00000000",
  64365=>"00000010",
  64366=>"00000101",
  64367=>"11111110",
  64368=>"11111111",
  64369=>"00000101",
  64370=>"11111110",
  64371=>"11111111",
  64372=>"00000000",
  64373=>"00000000",
  64374=>"00000010",
  64375=>"00000000",
  64376=>"11111111",
  64377=>"11111110",
  64378=>"11111100",
  64379=>"00000011",
  64380=>"11111101",
  64381=>"11111101",
  64382=>"11111101",
  64383=>"11111111",
  64384=>"00000000",
  64385=>"00000011",
  64386=>"00000011",
  64387=>"00000011",
  64388=>"11111110",
  64389=>"11111111",
  64390=>"00000011",
  64391=>"11111101",
  64392=>"00000000",
  64393=>"00000000",
  64394=>"00000010",
  64395=>"00000011",
  64396=>"11111110",
  64397=>"00000011",
  64398=>"11111110",
  64399=>"00000011",
  64400=>"00000001",
  64401=>"11111110",
  64402=>"11111111",
  64403=>"11111111",
  64404=>"11111101",
  64405=>"00000011",
  64406=>"00000010",
  64407=>"11111111",
  64408=>"11111111",
  64409=>"11111101",
  64410=>"00000101",
  64411=>"00000011",
  64412=>"11111111",
  64413=>"11111110",
  64414=>"00000100",
  64415=>"11111111",
  64416=>"00000000",
  64417=>"00000001",
  64418=>"00000001",
  64419=>"00000001",
  64420=>"00000001",
  64421=>"11111111",
  64422=>"00000100",
  64423=>"11111111",
  64424=>"11111100",
  64425=>"00000001",
  64426=>"11111110",
  64427=>"11111110",
  64428=>"00000100",
  64429=>"11111111",
  64430=>"11111110",
  64431=>"11111111",
  64432=>"11111101",
  64433=>"11111111",
  64434=>"11111111",
  64435=>"11111110",
  64436=>"11111111",
  64437=>"00000011",
  64438=>"11111110",
  64439=>"00000001",
  64440=>"00000010",
  64441=>"11111110",
  64442=>"11111110",
  64443=>"00000001",
  64444=>"11111111",
  64445=>"11111101",
  64446=>"00000000",
  64447=>"11111100",
  64448=>"00000011",
  64449=>"00000011",
  64450=>"00000010",
  64451=>"00000010",
  64452=>"11111111",
  64453=>"00000000",
  64454=>"11111111",
  64455=>"00000000",
  64456=>"00000010",
  64457=>"11111111",
  64458=>"11111111",
  64459=>"11111110",
  64460=>"11111101",
  64461=>"00000000",
  64462=>"00000100",
  64463=>"11111110",
  64464=>"00000011",
  64465=>"11111110",
  64466=>"11111101",
  64467=>"11111111",
  64468=>"00000010",
  64469=>"00000000",
  64470=>"11111100",
  64471=>"00000010",
  64472=>"00000010",
  64473=>"11111111",
  64474=>"11111111",
  64475=>"11111110",
  64476=>"11111111",
  64477=>"00000001",
  64478=>"11111110",
  64479=>"11111111",
  64480=>"00000001",
  64481=>"00000010",
  64482=>"00000000",
  64483=>"11111101",
  64484=>"00000001",
  64485=>"00000010",
  64486=>"11111111",
  64487=>"11111110",
  64488=>"11111101",
  64489=>"11111101",
  64490=>"11111101",
  64491=>"11111101",
  64492=>"00000000",
  64493=>"00000100",
  64494=>"11111111",
  64495=>"00000010",
  64496=>"11111100",
  64497=>"00000000",
  64498=>"11111101",
  64499=>"00000010",
  64500=>"11111101",
  64501=>"11111101",
  64502=>"00000001",
  64503=>"00000100",
  64504=>"00000000",
  64505=>"11111101",
  64506=>"11111100",
  64507=>"00000010",
  64508=>"00000100",
  64509=>"11111100",
  64510=>"11111110",
  64511=>"00000001");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;