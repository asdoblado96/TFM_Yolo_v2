LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_12_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_12_BNROM;

ARCHITECTURE RTL OF L8_12_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0001100111010000"&"0001111100001111",
  1=>"0001110011001011"&"0010011011010000",
  2=>"0010000101110111"&"0010010011000111",
  3=>"0000001001010001"&"0001100111111011",
  4=>"0000101111010100"&"0010000100000100",
  5=>"0001010010101000"&"0010001111000111",
  6=>"0001011001010100"&"0010001001001101",
  7=>"0010000111101100"&"0010010100101010",
  8=>"0000011000010011"&"0010010011100100",
  9=>"0000101110010011"&"0010011111110000",
  10=>"0001010010010100"&"0010011011110011",
  11=>"0000001110110100"&"0010001011001001",
  12=>"0001100010000111"&"0010001101100100",
  13=>"0010011110001111"&"0010010110000100",
  14=>"0010010010001001"&"0001110010111101",
  15=>"0001101010100010"&"0010000011011010",
  16=>"0001011110000010"&"0001101101111110",
  17=>"0001100000110101"&"0010001000100101",
  18=>"0010011101101010"&"0010001110111101",
  19=>"0000110100111100"&"0010100110010000",
  20=>"0001001101000101"&"0010001101101010",
  21=>"0000111010000111"&"0010001101101010",
  22=>"0000100111001001"&"0001101011110010",
  23=>"1111110001100000"&"0001111011000111",
  24=>"0001101111100011"&"0010010101100001",
  25=>"0000110111110101"&"0010001100001110",
  26=>"0001000000000110"&"0010000011011011",
  27=>"0000100110000111"&"0010010001101000",
  28=>"0001001101001101"&"0010001000001010",
  29=>"0001100111101000"&"0001110111001100",
  30=>"0001011100111001"&"0010001011010000",
  31=>"0000001100000010"&"0010000110111111",
  32=>"0010000110111001"&"0010011000100111",
  33=>"0001100101100110"&"0010000101111100",
  34=>"0000100110111000"&"0010011111000010",
  35=>"0000100000010110"&"0010001100001010",
  36=>"1111101111100111"&"0001111110000100",
  37=>"0001001001110000"&"0010001000111010",
  38=>"0000110101011010"&"0010011010111000",
  39=>"0001011110001000"&"0010011010010110",
  40=>"0010011100011100"&"0001111001110101",
  41=>"0000110001110110"&"0010000111011110",
  42=>"0001100010000111"&"0010011000101001",
  43=>"0010001010100111"&"0010011011011101",
  44=>"0010001100100000"&"0001110100111001",
  45=>"0000011101101000"&"0010011100101101",
  46=>"0000010100000110"&"0010001011101001",
  47=>"0000110000011111"&"0010010011101010",
  48=>"0000101010101001"&"0010001110101101",
  49=>"0010000011011011"&"0010001011000010",
  50=>"0000110111111111"&"0010000011000111",
  51=>"0001011010010101"&"0001110011001011",
  52=>"0001000001100110"&"0010011100011001",
  53=>"1111110010111011"&"0010010010110001",
  54=>"0001011100100110"&"0001110010110001",
  55=>"0001100101111001"&"0010010011101000",
  56=>"0000110111111101"&"0010001100100100",
  57=>"0000110110100001"&"0010000000101001",
  58=>"0001101000100000"&"0001111001000111",
  59=>"0001100011000100"&"0010010011011010",
  60=>"1111111100001111"&"0001110000011010",
  61=>"0010011011111101"&"0010011010110111",
  62=>"0001100100001111"&"0010011101110011",
  63=>"0010010110000101"&"0001111011010111");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;