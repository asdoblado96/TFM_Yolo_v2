LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_15_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_15_BNROM;

ARCHITECTURE RTL OF L8_15_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0010000110101111"&"0001110010000001",
  1=>"0000100110101011"&"0010010001100011",
  2=>"0001100010100101"&"0001110110001011",
  3=>"0001111110100010"&"0010010001011101",
  4=>"0010010000011001"&"0010001111101011",
  5=>"0010100010110110"&"0010010001111000",
  6=>"1111101111001111"&"0010000111101110",
  7=>"0001110010010110"&"0010011100111111",
  8=>"1111100100110110"&"0010000110000011",
  9=>"0001111111110100"&"0010011000010100",
  10=>"0001100000100111"&"0001110101001001",
  11=>"0001000111110000"&"0010000101000010",
  12=>"0000111111101001"&"0010010011110001",
  13=>"1110110110111101"&"0001100100101000",
  14=>"0000001110011110"&"0010011001111000",
  15=>"0001101000011110"&"0001101010111101",
  16=>"0001001100010101"&"0001100010100110",
  17=>"0000010110000010"&"0010100011100111",
  18=>"0000000101000111"&"0010011010101111",
  19=>"0001101011110000"&"0001110110001010",
  20=>"0000101000110101"&"0010000111000010",
  21=>"0000000110100101"&"0010010001010101",
  22=>"0001011011000010"&"0001110101110110",
  23=>"0001111001111100"&"0010010100100110",
  24=>"0000110110101101"&"0010000010110010",
  25=>"0000010000101011"&"0010000001100011",
  26=>"0001011100010101"&"0010010111100100",
  27=>"0001101001110111"&"0010010110111001",
  28=>"0001001100000011"&"0010010000010111",
  29=>"0000011010110100"&"0010000011101111",
  30=>"0000111011001111"&"0010010001000010",
  31=>"0001110010011010"&"0001110001111001",
  32=>"0001100011000100"&"0010100111100010",
  33=>"0001011100000101"&"0001110001010110",
  34=>"0000110101111100"&"0010010111001000",
  35=>"0010010101111000"&"0001110110100110",
  36=>"0001001000010011"&"0001110100010010",
  37=>"0000000111001101"&"0001110011110111",
  38=>"0000111110110100"&"0010010101110000",
  39=>"0000001011100111"&"0010010000100001",
  40=>"0001110100011100"&"0001110111111000",
  41=>"0001110101001110"&"0010001111100110",
  42=>"0000011100011100"&"0010010010110111",
  43=>"0010000110010101"&"0001111101110110",
  44=>"0001100110000101"&"0010001110011000",
  45=>"0001010110010000"&"0010001101001011",
  46=>"0010001000011011"&"0010000110111010",
  47=>"0001010100100100"&"0010000001001000",
  48=>"0011010011000011"&"0010001010001110",
  49=>"1111100101010011"&"0001101100010001",
  50=>"0001011000100011"&"0010011101100100",
  51=>"0001000111010011"&"0010011001010000",
  52=>"0001110111010001"&"0001111010101100",
  53=>"0000010111100011"&"0010011000111000",
  54=>"0000111010100100"&"0010010011001100",
  55=>"0010011110011100"&"0010001010000000",
  56=>"0001000001111000"&"0010000111110101",
  57=>"0001111100100000"&"0001110001101101",
  58=>"0001100110001110"&"0001111010000101",
  59=>"0000110010111110"&"0001110000000110",
  60=>"0001100101011101"&"0010010101100101",
  61=>"0000101010100001"&"0010100001001010",
  62=>"0001111100110110"&"0001111100011101",
  63=>"0001111001111111"&"0010001000001111");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;