LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_16_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_16_WROM;

ARCHITECTURE RTL OF L8_16_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"000110000",
  1=>"001101011",
  2=>"010101001",
  3=>"110101101",
  4=>"101001101",
  5=>"111001110",
  6=>"110010111",
  7=>"110000111",
  8=>"001000100",
  9=>"100110111",
  10=>"110101100",
  11=>"001100100",
  12=>"101011010",
  13=>"000101000",
  14=>"011011010",
  15=>"001101000",
  16=>"100001001",
  17=>"001000011",
  18=>"110001111",
  19=>"101010110",
  20=>"001101001",
  21=>"011010011",
  22=>"010110110",
  23=>"100011101",
  24=>"001110111",
  25=>"101011110",
  26=>"011000101",
  27=>"010001100",
  28=>"010001010",
  29=>"101100110",
  30=>"001111001",
  31=>"101000011",
  32=>"110011100",
  33=>"100001001",
  34=>"011010011",
  35=>"100101000",
  36=>"011010001",
  37=>"001110101",
  38=>"111011001",
  39=>"000111011",
  40=>"000100000",
  41=>"001001100",
  42=>"110101110",
  43=>"110101100",
  44=>"011111000",
  45=>"110100010",
  46=>"111111101",
  47=>"011011001",
  48=>"011001011",
  49=>"001100010",
  50=>"101100110",
  51=>"111000101",
  52=>"011001011",
  53=>"000100011",
  54=>"010100000",
  55=>"000100010",
  56=>"110000000",
  57=>"000110110",
  58=>"011000101",
  59=>"101110100",
  60=>"001010110",
  61=>"101001010",
  62=>"000100010",
  63=>"111101001",
  64=>"111110111",
  65=>"100001111",
  66=>"011001111",
  67=>"100000011",
  68=>"011001000",
  69=>"001001111",
  70=>"011000110",
  71=>"100111011",
  72=>"000101001",
  73=>"101110101",
  74=>"111010010",
  75=>"011000010",
  76=>"001111011",
  77=>"001111111",
  78=>"101001101",
  79=>"111011110",
  80=>"110000000",
  81=>"110000000",
  82=>"110110011",
  83=>"110011101",
  84=>"110001100",
  85=>"101000001",
  86=>"101100001",
  87=>"110001111",
  88=>"100111100",
  89=>"100110001",
  90=>"111011000",
  91=>"000010000",
  92=>"001101111",
  93=>"001100100",
  94=>"000010010",
  95=>"100000100",
  96=>"110001101",
  97=>"000001110",
  98=>"011010111",
  99=>"001011110",
  100=>"011001010",
  101=>"001101111",
  102=>"101101111",
  103=>"101011111",
  104=>"100111110",
  105=>"101100001",
  106=>"010010011",
  107=>"111001111",
  108=>"000101101",
  109=>"010110001",
  110=>"001000111",
  111=>"100011101",
  112=>"011100010",
  113=>"000100100",
  114=>"000100000",
  115=>"110010111",
  116=>"000000101",
  117=>"010010100",
  118=>"001000100",
  119=>"111011011",
  120=>"111010101",
  121=>"111011000",
  122=>"111010101",
  123=>"001000000",
  124=>"110110011",
  125=>"000011011",
  126=>"011000000",
  127=>"111111110",
  128=>"100100110",
  129=>"100111011",
  130=>"111001110",
  131=>"110000101",
  132=>"111101100",
  133=>"000000100",
  134=>"100111000",
  135=>"001001100",
  136=>"100101010",
  137=>"000110110",
  138=>"111000101",
  139=>"011100001",
  140=>"001011101",
  141=>"010110100",
  142=>"000110111",
  143=>"001000010",
  144=>"000110001",
  145=>"100100011",
  146=>"001101100",
  147=>"001000000",
  148=>"110101111",
  149=>"110011010",
  150=>"101101100",
  151=>"111101110",
  152=>"101011101",
  153=>"110100001",
  154=>"100010100",
  155=>"011011001",
  156=>"110001100",
  157=>"111111011",
  158=>"001000001",
  159=>"101101110",
  160=>"000100011",
  161=>"010111000",
  162=>"100001001",
  163=>"110000110",
  164=>"100100100",
  165=>"110101110",
  166=>"100000000",
  167=>"010100011",
  168=>"011011101",
  169=>"000000100",
  170=>"111000001",
  171=>"000001100",
  172=>"010110001",
  173=>"000111111",
  174=>"011110010",
  175=>"110110011",
  176=>"000010001",
  177=>"111111100",
  178=>"111000000",
  179=>"001010110",
  180=>"111110111",
  181=>"010011010",
  182=>"001000011",
  183=>"011101001",
  184=>"011100100",
  185=>"111111100",
  186=>"100111101",
  187=>"000001101",
  188=>"000011100",
  189=>"000001001",
  190=>"111101100",
  191=>"100100100",
  192=>"101010101",
  193=>"101000100",
  194=>"101111000",
  195=>"000101101",
  196=>"111110111",
  197=>"111001101",
  198=>"110101011",
  199=>"111011101",
  200=>"100010110",
  201=>"111010000",
  202=>"100011001",
  203=>"001110000",
  204=>"000011110",
  205=>"011111111",
  206=>"111011111",
  207=>"010000000",
  208=>"010010001",
  209=>"110110010",
  210=>"011110000",
  211=>"101101011",
  212=>"011101000",
  213=>"100111101",
  214=>"111000010",
  215=>"010001001",
  216=>"001001000",
  217=>"011110101",
  218=>"100000111",
  219=>"111110100",
  220=>"111010010",
  221=>"010111010",
  222=>"101011010",
  223=>"001100000",
  224=>"100111011",
  225=>"101110100",
  226=>"100111101",
  227=>"011000101",
  228=>"111011010",
  229=>"010001010",
  230=>"101101110",
  231=>"111101010",
  232=>"010111001",
  233=>"100001100",
  234=>"101101111",
  235=>"001000000",
  236=>"001010111",
  237=>"110100100",
  238=>"010001100",
  239=>"110010110",
  240=>"010000111",
  241=>"111110010",
  242=>"111100111",
  243=>"100011111",
  244=>"101010110",
  245=>"110001000",
  246=>"101100001",
  247=>"110110111",
  248=>"111011010",
  249=>"000011011",
  250=>"000110011",
  251=>"001010111",
  252=>"101100000",
  253=>"110110101",
  254=>"000010100",
  255=>"011000000",
  256=>"010100110",
  257=>"110111000",
  258=>"110000111",
  259=>"000101100",
  260=>"010001101",
  261=>"001011100",
  262=>"111111110",
  263=>"000110101",
  264=>"111100110",
  265=>"100001111",
  266=>"100010110",
  267=>"110100100",
  268=>"111111110",
  269=>"111000011",
  270=>"011100100",
  271=>"111000100",
  272=>"101111010",
  273=>"110001011",
  274=>"011010110",
  275=>"010001010",
  276=>"100011000",
  277=>"100110111",
  278=>"011010101",
  279=>"011101101",
  280=>"111011000",
  281=>"001001111",
  282=>"011100111",
  283=>"101011000",
  284=>"101111100",
  285=>"010100110",
  286=>"100001011",
  287=>"001010010",
  288=>"100011000",
  289=>"101100011",
  290=>"000000010",
  291=>"001000001",
  292=>"010101001",
  293=>"000011010",
  294=>"100000010",
  295=>"001010001",
  296=>"011100010",
  297=>"000000001",
  298=>"101100010",
  299=>"101100101",
  300=>"000000111",
  301=>"110010001",
  302=>"011011001",
  303=>"100101111",
  304=>"010000011",
  305=>"000000111",
  306=>"010100110",
  307=>"101011110",
  308=>"110100111",
  309=>"100110000",
  310=>"010101110",
  311=>"110001000",
  312=>"011110011",
  313=>"011100111",
  314=>"001100001",
  315=>"010110010",
  316=>"111101011",
  317=>"110101111",
  318=>"101100101",
  319=>"011001101",
  320=>"111000110",
  321=>"000100001",
  322=>"000001101",
  323=>"100011001",
  324=>"011100011",
  325=>"000110011",
  326=>"110000110",
  327=>"010000000",
  328=>"000010010",
  329=>"111101110",
  330=>"011101111",
  331=>"010101110",
  332=>"111001011",
  333=>"111010100",
  334=>"101000001",
  335=>"011000100",
  336=>"010101010",
  337=>"000100001",
  338=>"101101011",
  339=>"010111111",
  340=>"000011001",
  341=>"000000011",
  342=>"111100111",
  343=>"000011010",
  344=>"111111110",
  345=>"000000011",
  346=>"111100000",
  347=>"011001000",
  348=>"011000100",
  349=>"010001111",
  350=>"110011100",
  351=>"000100011",
  352=>"101111110",
  353=>"101001101",
  354=>"100111110",
  355=>"001001000",
  356=>"001111100",
  357=>"010001010",
  358=>"001010001",
  359=>"111000110",
  360=>"110110000",
  361=>"010111100",
  362=>"101101100",
  363=>"101111111",
  364=>"001110110",
  365=>"000100000",
  366=>"000000011",
  367=>"100111101",
  368=>"110101100",
  369=>"110110110",
  370=>"100110011",
  371=>"000110111",
  372=>"101000010",
  373=>"110010011",
  374=>"110110100",
  375=>"110001101",
  376=>"010000001",
  377=>"111010000",
  378=>"110111100",
  379=>"001000110",
  380=>"101111011",
  381=>"100101001",
  382=>"101111010",
  383=>"010100110",
  384=>"101111101",
  385=>"101000000",
  386=>"111010011",
  387=>"100110010",
  388=>"101011001",
  389=>"001000000",
  390=>"101010110",
  391=>"101010100",
  392=>"000011101",
  393=>"110001001",
  394=>"010010010",
  395=>"010010101",
  396=>"000001001",
  397=>"100000011",
  398=>"011101110",
  399=>"001011110",
  400=>"000011010",
  401=>"101110001",
  402=>"001000110",
  403=>"101100001",
  404=>"011001100",
  405=>"111011000",
  406=>"000000001",
  407=>"011011101",
  408=>"011100010",
  409=>"011001101",
  410=>"001101110",
  411=>"010100101",
  412=>"010010100",
  413=>"001001000",
  414=>"100111011",
  415=>"101011111",
  416=>"111101001",
  417=>"001001101",
  418=>"010111100",
  419=>"010100010",
  420=>"101100011",
  421=>"011110010",
  422=>"111010000",
  423=>"110110100",
  424=>"111011011",
  425=>"110000011",
  426=>"101010011",
  427=>"011100010",
  428=>"010011010",
  429=>"000000111",
  430=>"110101110",
  431=>"101011000",
  432=>"101010100",
  433=>"101001111",
  434=>"010110010",
  435=>"101001001",
  436=>"011101101",
  437=>"011000010",
  438=>"010010000",
  439=>"111101000",
  440=>"010001100",
  441=>"011011101",
  442=>"100100010",
  443=>"110010010",
  444=>"010011011",
  445=>"111000110",
  446=>"001011101",
  447=>"101010001",
  448=>"000001010",
  449=>"000000010",
  450=>"110111001",
  451=>"011110001",
  452=>"000111101",
  453=>"001000111",
  454=>"101100010",
  455=>"110000110",
  456=>"110011101",
  457=>"101001001",
  458=>"111101111",
  459=>"100111110",
  460=>"001000010",
  461=>"111100111",
  462=>"010000000",
  463=>"001100110",
  464=>"111111111",
  465=>"101111111",
  466=>"101111100",
  467=>"110110111",
  468=>"011011000",
  469=>"010010011",
  470=>"000110111",
  471=>"010010101",
  472=>"110001000",
  473=>"000000100",
  474=>"101011111",
  475=>"101010011",
  476=>"001110101",
  477=>"111100101",
  478=>"011100001",
  479=>"101001010",
  480=>"010001100",
  481=>"010110010",
  482=>"001010100",
  483=>"000111111",
  484=>"111111001",
  485=>"000000000",
  486=>"110011001",
  487=>"100100111",
  488=>"110101010",
  489=>"111100000",
  490=>"101001111",
  491=>"000011111",
  492=>"001110000",
  493=>"110010101",
  494=>"110001001",
  495=>"001011111",
  496=>"100000001",
  497=>"101011100",
  498=>"110110010",
  499=>"001000000",
  500=>"111011111",
  501=>"111000100",
  502=>"001110010",
  503=>"101010010",
  504=>"010101010",
  505=>"011110101",
  506=>"100010110",
  507=>"011111111",
  508=>"110101011",
  509=>"110100101",
  510=>"001011001",
  511=>"100000111",
  512=>"110001101",
  513=>"110100111",
  514=>"000100010",
  515=>"000101000",
  516=>"010010001",
  517=>"100010110",
  518=>"111000110",
  519=>"011111101",
  520=>"000101110",
  521=>"011111001",
  522=>"110111111",
  523=>"011110000",
  524=>"101101111",
  525=>"011001011",
  526=>"000100100",
  527=>"011111111",
  528=>"100101000",
  529=>"011110111",
  530=>"000110010",
  531=>"011001100",
  532=>"010001011",
  533=>"110110001",
  534=>"111111100",
  535=>"000011100",
  536=>"111001010",
  537=>"111111000",
  538=>"101000011",
  539=>"000010001",
  540=>"010000000",
  541=>"111000101",
  542=>"111111101",
  543=>"100001110",
  544=>"010001110",
  545=>"010011111",
  546=>"001001000",
  547=>"011010111",
  548=>"101011011",
  549=>"000111011",
  550=>"001001111",
  551=>"111010011",
  552=>"101001000",
  553=>"110110100",
  554=>"000011110",
  555=>"100110010",
  556=>"000100111",
  557=>"010101100",
  558=>"111111000",
  559=>"110110101",
  560=>"101100000",
  561=>"100110011",
  562=>"011100101",
  563=>"010111110",
  564=>"110111011",
  565=>"110100111",
  566=>"111111001",
  567=>"100100000",
  568=>"001111101",
  569=>"011110010",
  570=>"010111001",
  571=>"010010001",
  572=>"100110110",
  573=>"001001000",
  574=>"000011001",
  575=>"000001101",
  576=>"101100000",
  577=>"000101110",
  578=>"111100000",
  579=>"101010001",
  580=>"000100001",
  581=>"100010110",
  582=>"111010101",
  583=>"011001010",
  584=>"000011111",
  585=>"010110111",
  586=>"110101011",
  587=>"001001110",
  588=>"101000011",
  589=>"011011111",
  590=>"001001010",
  591=>"010101011",
  592=>"101111101",
  593=>"110110101",
  594=>"001100101",
  595=>"110000000",
  596=>"000101111",
  597=>"001011101",
  598=>"010001000",
  599=>"100000001",
  600=>"010101100",
  601=>"001101100",
  602=>"110111110",
  603=>"000110100",
  604=>"101011110",
  605=>"111010110",
  606=>"101100001",
  607=>"011111011",
  608=>"100001011",
  609=>"110110111",
  610=>"110100011",
  611=>"110111011",
  612=>"101000010",
  613=>"000001100",
  614=>"101001110",
  615=>"010111011",
  616=>"011010001",
  617=>"111110010",
  618=>"100001100",
  619=>"100000101",
  620=>"011000010",
  621=>"001010001",
  622=>"110100110",
  623=>"111111101",
  624=>"001001111",
  625=>"001100001",
  626=>"101110101",
  627=>"010010101",
  628=>"001001100",
  629=>"000000000",
  630=>"011011101",
  631=>"111101010",
  632=>"110001111",
  633=>"101011001",
  634=>"111011000",
  635=>"011011010",
  636=>"001100111",
  637=>"011111010",
  638=>"001000010",
  639=>"101101100",
  640=>"111100011",
  641=>"101000111",
  642=>"110010011",
  643=>"001001111",
  644=>"001011100",
  645=>"100011110",
  646=>"100000011",
  647=>"000010110",
  648=>"110110011",
  649=>"001101100",
  650=>"111101101",
  651=>"100100010",
  652=>"010001011",
  653=>"000001111",
  654=>"110001100",
  655=>"111001001",
  656=>"111110010",
  657=>"110111000",
  658=>"010011110",
  659=>"101000011",
  660=>"011010110",
  661=>"010010101",
  662=>"101111000",
  663=>"001001001",
  664=>"010000010",
  665=>"101110110",
  666=>"000011000",
  667=>"000100010",
  668=>"101111001",
  669=>"010101111",
  670=>"001110100",
  671=>"110100111",
  672=>"000010100",
  673=>"110000111",
  674=>"100000110",
  675=>"110100101",
  676=>"101010011",
  677=>"010000110",
  678=>"101101011",
  679=>"000101110",
  680=>"010101011",
  681=>"001101001",
  682=>"001100101",
  683=>"100000010",
  684=>"101100110",
  685=>"000100001",
  686=>"010011111",
  687=>"000110111",
  688=>"001000000",
  689=>"011110011",
  690=>"101011011",
  691=>"011111111",
  692=>"110111110",
  693=>"110111010",
  694=>"100101000",
  695=>"010100000",
  696=>"111010101",
  697=>"000001011",
  698=>"000001010",
  699=>"111011100",
  700=>"111110000",
  701=>"110110100",
  702=>"110000011",
  703=>"011011011",
  704=>"101111111",
  705=>"011100111",
  706=>"100101001",
  707=>"011101010",
  708=>"110001011",
  709=>"010010011",
  710=>"110001110",
  711=>"000000100",
  712=>"111001010",
  713=>"101000011",
  714=>"010000100",
  715=>"111100101",
  716=>"110110111",
  717=>"100111001",
  718=>"011011111",
  719=>"100011011",
  720=>"101000011",
  721=>"111111110",
  722=>"001000000",
  723=>"011000100",
  724=>"101101010",
  725=>"100111111",
  726=>"100110101",
  727=>"110010000",
  728=>"111111101",
  729=>"110101100",
  730=>"110000111",
  731=>"011100110",
  732=>"100101111",
  733=>"111111000",
  734=>"101001000",
  735=>"000111101",
  736=>"100010110",
  737=>"011001010",
  738=>"110000001",
  739=>"100010110",
  740=>"001111000",
  741=>"111001101",
  742=>"100100100",
  743=>"000000001",
  744=>"100100100",
  745=>"111110000",
  746=>"101100011",
  747=>"011001101",
  748=>"110001110",
  749=>"011101110",
  750=>"011001000",
  751=>"100001100",
  752=>"100000101",
  753=>"111100100",
  754=>"111100110",
  755=>"100011111",
  756=>"111001001",
  757=>"001111001",
  758=>"110111010",
  759=>"011000001",
  760=>"000110000",
  761=>"110000111",
  762=>"110010101",
  763=>"011010000",
  764=>"011001010",
  765=>"100001101",
  766=>"101110000",
  767=>"010110010",
  768=>"111011000",
  769=>"010101010",
  770=>"100110010",
  771=>"100100110",
  772=>"110111110",
  773=>"110110000",
  774=>"111100010",
  775=>"011110110",
  776=>"111101101",
  777=>"011001000",
  778=>"000011001",
  779=>"000111011",
  780=>"000010001",
  781=>"000010010",
  782=>"010101110",
  783=>"101101111",
  784=>"011100111",
  785=>"101000110",
  786=>"000000000",
  787=>"111001010",
  788=>"011101001",
  789=>"100011011",
  790=>"100100110",
  791=>"110100110",
  792=>"101011101",
  793=>"110000100",
  794=>"110011001",
  795=>"001100110",
  796=>"110001110",
  797=>"011110111",
  798=>"100011100",
  799=>"100010001",
  800=>"010011010",
  801=>"100010011",
  802=>"010110010",
  803=>"110101001",
  804=>"010110100",
  805=>"101110010",
  806=>"010000110",
  807=>"101001110",
  808=>"000000100",
  809=>"101100110",
  810=>"110000101",
  811=>"000000101",
  812=>"001010010",
  813=>"110110110",
  814=>"101001010",
  815=>"100001110",
  816=>"100111011",
  817=>"000100101",
  818=>"010000100",
  819=>"000000010",
  820=>"001001010",
  821=>"101011101",
  822=>"000011010",
  823=>"100100001",
  824=>"011111001",
  825=>"110101000",
  826=>"011010100",
  827=>"011101010",
  828=>"000000010",
  829=>"000000110",
  830=>"101111001",
  831=>"110101101",
  832=>"011001111",
  833=>"010101000",
  834=>"101101001",
  835=>"100001000",
  836=>"110111010",
  837=>"101110111",
  838=>"111111111",
  839=>"101101100",
  840=>"010010110",
  841=>"001111000",
  842=>"110101000",
  843=>"010100111",
  844=>"011010001",
  845=>"100101100",
  846=>"110101000",
  847=>"010011111",
  848=>"101100101",
  849=>"111111100",
  850=>"111010001",
  851=>"001101111",
  852=>"011101100",
  853=>"101101111",
  854=>"111111110",
  855=>"001001010",
  856=>"111111010",
  857=>"001100010",
  858=>"111011010",
  859=>"110111001",
  860=>"010110010",
  861=>"000101010",
  862=>"000000000",
  863=>"011110000",
  864=>"011101110",
  865=>"100011100",
  866=>"011001011",
  867=>"110001111",
  868=>"101010101",
  869=>"011011101",
  870=>"111101001",
  871=>"000101101",
  872=>"101001011",
  873=>"111101011",
  874=>"100100101",
  875=>"000010101",
  876=>"001100111",
  877=>"001001010",
  878=>"111101101",
  879=>"101100000",
  880=>"100001101",
  881=>"111000010",
  882=>"001111111",
  883=>"100000001",
  884=>"001111111",
  885=>"110010000",
  886=>"001011000",
  887=>"101011011",
  888=>"100100000",
  889=>"111110000",
  890=>"100001000",
  891=>"111010100",
  892=>"100100110",
  893=>"110111011",
  894=>"110010110",
  895=>"011000100",
  896=>"111111110",
  897=>"010010111",
  898=>"111010000",
  899=>"011100010",
  900=>"111110000",
  901=>"001001110",
  902=>"110011101",
  903=>"001000010",
  904=>"100100000",
  905=>"001001100",
  906=>"001000100",
  907=>"110000111",
  908=>"111011011",
  909=>"100110011",
  910=>"010111111",
  911=>"101110001",
  912=>"111111000",
  913=>"111001010",
  914=>"100110010",
  915=>"000101010",
  916=>"110101101",
  917=>"011100111",
  918=>"111101001",
  919=>"001100011",
  920=>"010011101",
  921=>"001111110",
  922=>"000001101",
  923=>"001000010",
  924=>"001001101",
  925=>"000111000",
  926=>"111101000",
  927=>"111100000",
  928=>"101010110",
  929=>"111000100",
  930=>"111100110",
  931=>"111011100",
  932=>"000010001",
  933=>"110111001",
  934=>"100010100",
  935=>"010010000",
  936=>"010001000",
  937=>"011101111",
  938=>"001001001",
  939=>"011001101",
  940=>"011110111",
  941=>"110101011",
  942=>"011101000",
  943=>"011101111",
  944=>"010101010",
  945=>"001100110",
  946=>"001100101",
  947=>"101010111",
  948=>"000010100",
  949=>"001100011",
  950=>"101010011",
  951=>"001101010",
  952=>"110101110",
  953=>"001001111",
  954=>"011000011",
  955=>"100100001",
  956=>"110001101",
  957=>"110001000",
  958=>"001010010",
  959=>"111001111",
  960=>"111000010",
  961=>"000010010",
  962=>"000101111",
  963=>"100010010",
  964=>"100110001",
  965=>"111101001",
  966=>"100100000",
  967=>"010101100",
  968=>"011001101",
  969=>"001100110",
  970=>"010100110",
  971=>"001111111",
  972=>"011111111",
  973=>"111110000",
  974=>"011101100",
  975=>"010110010",
  976=>"101100001",
  977=>"011101100",
  978=>"010101111",
  979=>"000011010",
  980=>"000100101",
  981=>"101111100",
  982=>"111011001",
  983=>"101000000",
  984=>"011100101",
  985=>"100111111",
  986=>"110011110",
  987=>"011110011",
  988=>"010010001",
  989=>"010010011",
  990=>"111000010",
  991=>"011001000",
  992=>"111011110",
  993=>"101100001",
  994=>"100100111",
  995=>"000111001",
  996=>"000011101",
  997=>"111011111",
  998=>"100010000",
  999=>"001101001",
  1000=>"000000011",
  1001=>"000111111",
  1002=>"010110000",
  1003=>"001111110",
  1004=>"100110101",
  1005=>"100100001",
  1006=>"011001010",
  1007=>"110011001",
  1008=>"100110111",
  1009=>"111110000",
  1010=>"000000101",
  1011=>"000011001",
  1012=>"101000110",
  1013=>"001010101",
  1014=>"111100011",
  1015=>"110110010",
  1016=>"010101000",
  1017=>"100010011",
  1018=>"010010001",
  1019=>"000110100",
  1020=>"011111111",
  1021=>"011101101",
  1022=>"111110101",
  1023=>"101011000",
  1024=>"101001011",
  1025=>"110101110",
  1026=>"111011010",
  1027=>"101111001",
  1028=>"011010001",
  1029=>"000110001",
  1030=>"001001001",
  1031=>"110101000",
  1032=>"011111001",
  1033=>"011011010",
  1034=>"110111101",
  1035=>"100000110",
  1036=>"100000010",
  1037=>"011100101",
  1038=>"101001100",
  1039=>"100100011",
  1040=>"110101011",
  1041=>"111100110",
  1042=>"010110110",
  1043=>"000110010",
  1044=>"000111110",
  1045=>"000011100",
  1046=>"000101101",
  1047=>"110100100",
  1048=>"110100111",
  1049=>"100000111",
  1050=>"110001100",
  1051=>"001110010",
  1052=>"001000010",
  1053=>"111100110",
  1054=>"001110011",
  1055=>"011100110",
  1056=>"000001111",
  1057=>"011101010",
  1058=>"110001000",
  1059=>"001001100",
  1060=>"110011101",
  1061=>"010110100",
  1062=>"101111101",
  1063=>"110101111",
  1064=>"001110011",
  1065=>"010001000",
  1066=>"111000011",
  1067=>"100011100",
  1068=>"110111001",
  1069=>"101010101",
  1070=>"001101010",
  1071=>"101110011",
  1072=>"110000110",
  1073=>"010011101",
  1074=>"110001101",
  1075=>"000100100",
  1076=>"000001011",
  1077=>"000101010",
  1078=>"110000101",
  1079=>"101001100",
  1080=>"110001110",
  1081=>"001000111",
  1082=>"010110100",
  1083=>"101001001",
  1084=>"011000000",
  1085=>"000001001",
  1086=>"001110110",
  1087=>"001100111",
  1088=>"110000001",
  1089=>"000110000",
  1090=>"010110011",
  1091=>"100000000",
  1092=>"111110111",
  1093=>"000011111",
  1094=>"111100000",
  1095=>"011111101",
  1096=>"100100011",
  1097=>"110101001",
  1098=>"000101111",
  1099=>"011110001",
  1100=>"111001000",
  1101=>"010111110",
  1102=>"100001111",
  1103=>"000101011",
  1104=>"001001110",
  1105=>"110100100",
  1106=>"100000110",
  1107=>"110010000",
  1108=>"100011001",
  1109=>"000100100",
  1110=>"011111101",
  1111=>"101011011",
  1112=>"110000111",
  1113=>"101111100",
  1114=>"110011100",
  1115=>"110000110",
  1116=>"100101000",
  1117=>"110000100",
  1118=>"000110001",
  1119=>"010110100",
  1120=>"111100111",
  1121=>"001011011",
  1122=>"001001100",
  1123=>"001010101",
  1124=>"000001001",
  1125=>"010100110",
  1126=>"010111101",
  1127=>"001100000",
  1128=>"100100001",
  1129=>"100100001",
  1130=>"000000010",
  1131=>"101101010",
  1132=>"111001000",
  1133=>"000000010",
  1134=>"100000110",
  1135=>"100011110",
  1136=>"100010011",
  1137=>"001111010",
  1138=>"011110101",
  1139=>"101100111",
  1140=>"000100000",
  1141=>"101101110",
  1142=>"011000010",
  1143=>"011111111",
  1144=>"101111101",
  1145=>"111101101",
  1146=>"110011110",
  1147=>"011100001",
  1148=>"011100100",
  1149=>"011110001",
  1150=>"111000001",
  1151=>"001001110",
  1152=>"001111111",
  1153=>"011111011",
  1154=>"001000001",
  1155=>"010010100",
  1156=>"001000111",
  1157=>"011101110",
  1158=>"111111101",
  1159=>"110100001",
  1160=>"100101100",
  1161=>"011000010",
  1162=>"000110111",
  1163=>"000110000",
  1164=>"101110101",
  1165=>"100111011",
  1166=>"000111000",
  1167=>"011100101",
  1168=>"110010111",
  1169=>"010100001",
  1170=>"101100100",
  1171=>"111001110",
  1172=>"000110110",
  1173=>"010000001",
  1174=>"010101111",
  1175=>"111110001",
  1176=>"000100111",
  1177=>"111100101",
  1178=>"000000110",
  1179=>"011001100",
  1180=>"110000100",
  1181=>"010001100",
  1182=>"111011110",
  1183=>"100100111",
  1184=>"001011110",
  1185=>"001100000",
  1186=>"001010110",
  1187=>"101011000",
  1188=>"110101010",
  1189=>"100101100",
  1190=>"110101110",
  1191=>"000100110",
  1192=>"100110111",
  1193=>"101110111",
  1194=>"001011100",
  1195=>"100111110",
  1196=>"011101101",
  1197=>"011010101",
  1198=>"110010001",
  1199=>"011101111",
  1200=>"001101100",
  1201=>"001110010",
  1202=>"001110101",
  1203=>"110000011",
  1204=>"110010110",
  1205=>"011001001",
  1206=>"011011000",
  1207=>"111111111",
  1208=>"100111100",
  1209=>"100001000",
  1210=>"101100111",
  1211=>"111110010",
  1212=>"101101001",
  1213=>"100001101",
  1214=>"001010011",
  1215=>"010010111",
  1216=>"111110110",
  1217=>"011000101",
  1218=>"001110100",
  1219=>"000101101",
  1220=>"101111011",
  1221=>"011010101",
  1222=>"000010010",
  1223=>"011010100",
  1224=>"001100110",
  1225=>"000111001",
  1226=>"011000101",
  1227=>"011000001",
  1228=>"101000100",
  1229=>"100001011",
  1230=>"000110101",
  1231=>"101101001",
  1232=>"011110110",
  1233=>"111100110",
  1234=>"010000011",
  1235=>"100111100",
  1236=>"111111100",
  1237=>"001000011",
  1238=>"111001100",
  1239=>"011101100",
  1240=>"000000100",
  1241=>"010001100",
  1242=>"011100011",
  1243=>"100010010",
  1244=>"111000101",
  1245=>"101010100",
  1246=>"010011010",
  1247=>"010100010",
  1248=>"000001010",
  1249=>"111011111",
  1250=>"001000100",
  1251=>"110010011",
  1252=>"100011000",
  1253=>"110010101",
  1254=>"101010101",
  1255=>"100001111",
  1256=>"111100101",
  1257=>"000100010",
  1258=>"110001010",
  1259=>"001110011",
  1260=>"000001000",
  1261=>"010001110",
  1262=>"110111000",
  1263=>"101010001",
  1264=>"000011101",
  1265=>"111011000",
  1266=>"011100111",
  1267=>"001110101",
  1268=>"100010011",
  1269=>"101001100",
  1270=>"110110111",
  1271=>"000000010",
  1272=>"011110111",
  1273=>"001101101",
  1274=>"010000000",
  1275=>"100111111",
  1276=>"001000001",
  1277=>"011111011",
  1278=>"100101110",
  1279=>"111111100",
  1280=>"010010110",
  1281=>"110111101",
  1282=>"000010011",
  1283=>"110111011",
  1284=>"110100101",
  1285=>"001111101",
  1286=>"100111111",
  1287=>"100010101",
  1288=>"001111100",
  1289=>"101001011",
  1290=>"010101111",
  1291=>"011010010",
  1292=>"001110110",
  1293=>"000101110",
  1294=>"011101110",
  1295=>"101011011",
  1296=>"100011010",
  1297=>"011001000",
  1298=>"011100100",
  1299=>"011010101",
  1300=>"010010011",
  1301=>"001010101",
  1302=>"010000101",
  1303=>"011000000",
  1304=>"100000001",
  1305=>"000010010",
  1306=>"011011011",
  1307=>"101100111",
  1308=>"110101111",
  1309=>"110001010",
  1310=>"011111100",
  1311=>"101101111",
  1312=>"100000000",
  1313=>"100010110",
  1314=>"111111100",
  1315=>"101011100",
  1316=>"011101010",
  1317=>"110101000",
  1318=>"001011010",
  1319=>"101101000",
  1320=>"000101010",
  1321=>"101011010",
  1322=>"101011111",
  1323=>"100101001",
  1324=>"101000001",
  1325=>"111011010",
  1326=>"000000001",
  1327=>"011110110",
  1328=>"010000111",
  1329=>"111001011",
  1330=>"100001000",
  1331=>"101011110",
  1332=>"111101101",
  1333=>"010110010",
  1334=>"110000000",
  1335=>"101111111",
  1336=>"000001101",
  1337=>"000100111",
  1338=>"010000000",
  1339=>"101111011",
  1340=>"111010100",
  1341=>"001100111",
  1342=>"011010111",
  1343=>"011010110",
  1344=>"111111000",
  1345=>"100001001",
  1346=>"000000101",
  1347=>"101100101",
  1348=>"011110110",
  1349=>"101111000",
  1350=>"010010001",
  1351=>"100011000",
  1352=>"000100110",
  1353=>"010010111",
  1354=>"101001011",
  1355=>"001000010",
  1356=>"101000100",
  1357=>"100111011",
  1358=>"001101000",
  1359=>"011001010",
  1360=>"001101101",
  1361=>"000010110",
  1362=>"101001110",
  1363=>"111000110",
  1364=>"100101010",
  1365=>"111010000",
  1366=>"100110110",
  1367=>"001111010",
  1368=>"100111100",
  1369=>"100001000",
  1370=>"110100101",
  1371=>"001101101",
  1372=>"101110001",
  1373=>"011100000",
  1374=>"011001010",
  1375=>"000100100",
  1376=>"001000000",
  1377=>"000110010",
  1378=>"011111111",
  1379=>"001000001",
  1380=>"001000100",
  1381=>"100000111",
  1382=>"101000111",
  1383=>"011101110",
  1384=>"010010111",
  1385=>"011001010",
  1386=>"110111110",
  1387=>"000110111",
  1388=>"001011100",
  1389=>"110011011",
  1390=>"000011110",
  1391=>"110110100",
  1392=>"010110110",
  1393=>"101010011",
  1394=>"111101111",
  1395=>"001011110",
  1396=>"010000001",
  1397=>"011010100",
  1398=>"000011111",
  1399=>"011100000",
  1400=>"010000101",
  1401=>"011001100",
  1402=>"000110110",
  1403=>"111101011",
  1404=>"000000000",
  1405=>"011110110",
  1406=>"001001001",
  1407=>"000011101",
  1408=>"101000010",
  1409=>"010010000",
  1410=>"101110001",
  1411=>"010110111",
  1412=>"011111101",
  1413=>"111101101",
  1414=>"111111110",
  1415=>"101101101",
  1416=>"001000001",
  1417=>"110001110",
  1418=>"101101100",
  1419=>"110001001",
  1420=>"111101111",
  1421=>"000011110",
  1422=>"010001010",
  1423=>"010011100",
  1424=>"111111011",
  1425=>"011000011",
  1426=>"011001000",
  1427=>"001110011",
  1428=>"101100000",
  1429=>"010000000",
  1430=>"111010110",
  1431=>"001011111",
  1432=>"010100110",
  1433=>"001000001",
  1434=>"101101001",
  1435=>"100100010",
  1436=>"110110000",
  1437=>"010111110",
  1438=>"100100101",
  1439=>"100011011",
  1440=>"000100001",
  1441=>"011011101",
  1442=>"100000100",
  1443=>"110000110",
  1444=>"101001010",
  1445=>"100101110",
  1446=>"011000000",
  1447=>"101011100",
  1448=>"100101010",
  1449=>"011111001",
  1450=>"110010111",
  1451=>"010000000",
  1452=>"100101111",
  1453=>"001001000",
  1454=>"010001000",
  1455=>"110111011",
  1456=>"101000000",
  1457=>"000000110",
  1458=>"100101100",
  1459=>"000001001",
  1460=>"101000111",
  1461=>"011101100",
  1462=>"101110000",
  1463=>"111010010",
  1464=>"000001100",
  1465=>"000001000",
  1466=>"001001010",
  1467=>"010000001",
  1468=>"000000010",
  1469=>"110011000",
  1470=>"111100111",
  1471=>"111011000",
  1472=>"011001111",
  1473=>"001010000",
  1474=>"100011011",
  1475=>"010110111",
  1476=>"011101110",
  1477=>"100010000",
  1478=>"011111111",
  1479=>"100000000",
  1480=>"011010011",
  1481=>"100001111",
  1482=>"110001001",
  1483=>"010010011",
  1484=>"000110010",
  1485=>"110010100",
  1486=>"000000011",
  1487=>"011011011",
  1488=>"100010100",
  1489=>"101101000",
  1490=>"011001100",
  1491=>"111011110",
  1492=>"000000111",
  1493=>"010000111",
  1494=>"110111001",
  1495=>"110111011",
  1496=>"101100011",
  1497=>"100011011",
  1498=>"110101001",
  1499=>"101000000",
  1500=>"110101011",
  1501=>"111110111",
  1502=>"111011000",
  1503=>"001101010",
  1504=>"010111011",
  1505=>"000010101",
  1506=>"110111011",
  1507=>"001101101",
  1508=>"000000000",
  1509=>"111110101",
  1510=>"001001010",
  1511=>"110001101",
  1512=>"011101010",
  1513=>"001011000",
  1514=>"110101010",
  1515=>"100111101",
  1516=>"001110001",
  1517=>"000001101",
  1518=>"100111101",
  1519=>"111100000",
  1520=>"011000110",
  1521=>"001100110",
  1522=>"111000111",
  1523=>"001010110",
  1524=>"100011011",
  1525=>"101101011",
  1526=>"101001010",
  1527=>"101001001",
  1528=>"100110110",
  1529=>"110101011",
  1530=>"001110000",
  1531=>"011100100",
  1532=>"111000010",
  1533=>"000000110",
  1534=>"110100111",
  1535=>"101101011",
  1536=>"111001001",
  1537=>"111101101",
  1538=>"011101100",
  1539=>"001011110",
  1540=>"100010000",
  1541=>"001111010",
  1542=>"000010110",
  1543=>"010100010",
  1544=>"111010101",
  1545=>"110101111",
  1546=>"000010001",
  1547=>"101000011",
  1548=>"010010101",
  1549=>"000100010",
  1550=>"110110011",
  1551=>"110000000",
  1552=>"001110101",
  1553=>"011000111",
  1554=>"100100010",
  1555=>"010101010",
  1556=>"101011001",
  1557=>"011011001",
  1558=>"100000000",
  1559=>"000011000",
  1560=>"101101111",
  1561=>"001010011",
  1562=>"000000111",
  1563=>"111100101",
  1564=>"010110000",
  1565=>"110100110",
  1566=>"010000001",
  1567=>"001111100",
  1568=>"011111111",
  1569=>"110010010",
  1570=>"101000001",
  1571=>"000001111",
  1572=>"000101010",
  1573=>"111110011",
  1574=>"011011000",
  1575=>"001110100",
  1576=>"111101000",
  1577=>"001111101",
  1578=>"001000000",
  1579=>"101101101",
  1580=>"001000010",
  1581=>"001111101",
  1582=>"011101010",
  1583=>"111111100",
  1584=>"111010111",
  1585=>"111011001",
  1586=>"011000101",
  1587=>"010011000",
  1588=>"010010010",
  1589=>"100001100",
  1590=>"101110100",
  1591=>"010101100",
  1592=>"101111011",
  1593=>"110001110",
  1594=>"000010010",
  1595=>"010100000",
  1596=>"100011101",
  1597=>"111111011",
  1598=>"000000110",
  1599=>"010011110",
  1600=>"010101001",
  1601=>"001111001",
  1602=>"011011100",
  1603=>"010011100",
  1604=>"110010110",
  1605=>"110101011",
  1606=>"001001010",
  1607=>"001010001",
  1608=>"101100000",
  1609=>"011110101",
  1610=>"101110000",
  1611=>"010000100",
  1612=>"100000001",
  1613=>"010000011",
  1614=>"110001101",
  1615=>"010010100",
  1616=>"111110000",
  1617=>"000111101",
  1618=>"100111111",
  1619=>"101001111",
  1620=>"110110000",
  1621=>"100111110",
  1622=>"001010100",
  1623=>"110101101",
  1624=>"000000110",
  1625=>"111101101",
  1626=>"101010011",
  1627=>"001000010",
  1628=>"110111011",
  1629=>"001000000",
  1630=>"010011001",
  1631=>"000110101",
  1632=>"010100101",
  1633=>"101111010",
  1634=>"000101111",
  1635=>"010011010",
  1636=>"110111010",
  1637=>"000001001",
  1638=>"001110110",
  1639=>"111011000",
  1640=>"000000000",
  1641=>"000101100",
  1642=>"001001001",
  1643=>"111000011",
  1644=>"111011110",
  1645=>"000100011",
  1646=>"111011000",
  1647=>"000001100",
  1648=>"110101011",
  1649=>"010010100",
  1650=>"100011101",
  1651=>"000111010",
  1652=>"001010000",
  1653=>"101111001",
  1654=>"111101111",
  1655=>"100110101",
  1656=>"001011101",
  1657=>"111011001",
  1658=>"111111011",
  1659=>"110011001",
  1660=>"000011001",
  1661=>"100100111",
  1662=>"001101011",
  1663=>"010100100",
  1664=>"100110111",
  1665=>"111100010",
  1666=>"000001000",
  1667=>"000010010",
  1668=>"111011111",
  1669=>"011101000",
  1670=>"100000110",
  1671=>"110001110",
  1672=>"001001111",
  1673=>"001110101",
  1674=>"001000100",
  1675=>"110110111",
  1676=>"010001001",
  1677=>"010010100",
  1678=>"011101111",
  1679=>"001100000",
  1680=>"101111111",
  1681=>"111001011",
  1682=>"011110111",
  1683=>"101100011",
  1684=>"001100111",
  1685=>"100100001",
  1686=>"111101110",
  1687=>"100100100",
  1688=>"011111000",
  1689=>"000011000",
  1690=>"101101110",
  1691=>"000000001",
  1692=>"001001111",
  1693=>"000010011",
  1694=>"001010111",
  1695=>"101010111",
  1696=>"110110100",
  1697=>"011111001",
  1698=>"010001110",
  1699=>"100001011",
  1700=>"110101011",
  1701=>"111010111",
  1702=>"010111010",
  1703=>"001010111",
  1704=>"101011111",
  1705=>"011100100",
  1706=>"101100100",
  1707=>"001110111",
  1708=>"001000101",
  1709=>"001011000",
  1710=>"001110000",
  1711=>"011011110",
  1712=>"010001111",
  1713=>"110000111",
  1714=>"001000000",
  1715=>"100011111",
  1716=>"010110101",
  1717=>"110111010",
  1718=>"101110011",
  1719=>"111111000",
  1720=>"110010101",
  1721=>"111101001",
  1722=>"101100001",
  1723=>"100011101",
  1724=>"101111000",
  1725=>"011000011",
  1726=>"011001011",
  1727=>"011011000",
  1728=>"111000100",
  1729=>"110000101",
  1730=>"101001010",
  1731=>"010010010",
  1732=>"001100010",
  1733=>"011001010",
  1734=>"100100011",
  1735=>"011100101",
  1736=>"100010000",
  1737=>"001101011",
  1738=>"111010101",
  1739=>"010111001",
  1740=>"011100000",
  1741=>"100000101",
  1742=>"010000011",
  1743=>"000101100",
  1744=>"100000101",
  1745=>"001011001",
  1746=>"001000001",
  1747=>"111110100",
  1748=>"011110110",
  1749=>"000011111",
  1750=>"001111100",
  1751=>"100001101",
  1752=>"111101001",
  1753=>"011001111",
  1754=>"010000010",
  1755=>"000100000",
  1756=>"001111111",
  1757=>"110000101",
  1758=>"000100001",
  1759=>"011011011",
  1760=>"100010100",
  1761=>"011100101",
  1762=>"101000010",
  1763=>"011110011",
  1764=>"110111000",
  1765=>"100000010",
  1766=>"111001010",
  1767=>"001001111",
  1768=>"001100010",
  1769=>"001110101",
  1770=>"010001010",
  1771=>"001110111",
  1772=>"110110010",
  1773=>"001110001",
  1774=>"010011011",
  1775=>"000000100",
  1776=>"011110011",
  1777=>"110001101",
  1778=>"000001000",
  1779=>"000001011",
  1780=>"000010000",
  1781=>"111100000",
  1782=>"110101011",
  1783=>"001111010",
  1784=>"110000100",
  1785=>"101001100",
  1786=>"000000001",
  1787=>"110010111",
  1788=>"100000001",
  1789=>"001100111",
  1790=>"010001111",
  1791=>"100111101",
  1792=>"001111100",
  1793=>"111000001",
  1794=>"100011010",
  1795=>"101000101",
  1796=>"110111100",
  1797=>"000001000",
  1798=>"010100101",
  1799=>"100110110",
  1800=>"110110010",
  1801=>"011111101",
  1802=>"001000011",
  1803=>"001000100",
  1804=>"111011000",
  1805=>"101101101",
  1806=>"001000010",
  1807=>"000000011",
  1808=>"111010111",
  1809=>"111110001",
  1810=>"100101011",
  1811=>"110010011",
  1812=>"111000011",
  1813=>"100010111",
  1814=>"000010111",
  1815=>"011100111",
  1816=>"000010000",
  1817=>"001101000",
  1818=>"010011101",
  1819=>"100000000",
  1820=>"011111011",
  1821=>"110000001",
  1822=>"010111001",
  1823=>"110011001",
  1824=>"000001000",
  1825=>"110010110",
  1826=>"010010011",
  1827=>"011110000",
  1828=>"110010101",
  1829=>"001110111",
  1830=>"001100110",
  1831=>"100110011",
  1832=>"010010111",
  1833=>"100101101",
  1834=>"101110011",
  1835=>"111111100",
  1836=>"111111111",
  1837=>"110110110",
  1838=>"010000000",
  1839=>"110011110",
  1840=>"011010011",
  1841=>"100100100",
  1842=>"110010010",
  1843=>"011011001",
  1844=>"111111110",
  1845=>"111110010",
  1846=>"111010100",
  1847=>"101101011",
  1848=>"110011100",
  1849=>"010010000",
  1850=>"100100010",
  1851=>"111010011",
  1852=>"010100111",
  1853=>"100011001",
  1854=>"111100110",
  1855=>"001000001",
  1856=>"100100000",
  1857=>"111100101",
  1858=>"101001110",
  1859=>"010111000",
  1860=>"101001000",
  1861=>"111011110",
  1862=>"111101011",
  1863=>"000111101",
  1864=>"000010100",
  1865=>"110110100",
  1866=>"111010000",
  1867=>"100110001",
  1868=>"000011110",
  1869=>"101101101",
  1870=>"100101110",
  1871=>"010000010",
  1872=>"001110110",
  1873=>"000101011",
  1874=>"111001001",
  1875=>"110111000",
  1876=>"111000100",
  1877=>"000001001",
  1878=>"100001000",
  1879=>"101101101",
  1880=>"111010000",
  1881=>"001000010",
  1882=>"010101101",
  1883=>"001001001",
  1884=>"010110011",
  1885=>"000011010",
  1886=>"100100010",
  1887=>"011000010",
  1888=>"000000010",
  1889=>"011011110",
  1890=>"010110101",
  1891=>"100110011",
  1892=>"101101000",
  1893=>"100001000",
  1894=>"011101100",
  1895=>"000111001",
  1896=>"101001100",
  1897=>"010111000",
  1898=>"100001010",
  1899=>"101111110",
  1900=>"000001000",
  1901=>"001000010",
  1902=>"000000000",
  1903=>"010011110",
  1904=>"000100111",
  1905=>"100100000",
  1906=>"111110101",
  1907=>"010011110",
  1908=>"001011110",
  1909=>"000110100",
  1910=>"000001101",
  1911=>"010111101",
  1912=>"101111110",
  1913=>"110111111",
  1914=>"100011111",
  1915=>"011010101",
  1916=>"000000010",
  1917=>"010000010",
  1918=>"011110011",
  1919=>"111110101",
  1920=>"011100000",
  1921=>"000101101",
  1922=>"010011001",
  1923=>"000110010",
  1924=>"000101110",
  1925=>"110110000",
  1926=>"001010001",
  1927=>"010111110",
  1928=>"000111111",
  1929=>"000001110",
  1930=>"011000110",
  1931=>"111100001",
  1932=>"101100100",
  1933=>"010100011",
  1934=>"010101001",
  1935=>"000001010",
  1936=>"010010111",
  1937=>"011101110",
  1938=>"111111011",
  1939=>"011111100",
  1940=>"001001010",
  1941=>"110110010",
  1942=>"110101100",
  1943=>"101001011",
  1944=>"011000111",
  1945=>"100000000",
  1946=>"011111100",
  1947=>"001010100",
  1948=>"010000010",
  1949=>"100100100",
  1950=>"100001010",
  1951=>"010010111",
  1952=>"000001000",
  1953=>"110100010",
  1954=>"111010000",
  1955=>"100000001",
  1956=>"001011111",
  1957=>"011010010",
  1958=>"111101010",
  1959=>"101001011",
  1960=>"101011000",
  1961=>"100111110",
  1962=>"111101110",
  1963=>"110011100",
  1964=>"111100010",
  1965=>"101100001",
  1966=>"010000011",
  1967=>"111000100",
  1968=>"000101011",
  1969=>"000111010",
  1970=>"000101100",
  1971=>"000100011",
  1972=>"011001000",
  1973=>"100000000",
  1974=>"001011101",
  1975=>"011110000",
  1976=>"010110110",
  1977=>"100001110",
  1978=>"001000011",
  1979=>"101100011",
  1980=>"100110011",
  1981=>"110010110",
  1982=>"000000110",
  1983=>"110001100",
  1984=>"000001011",
  1985=>"000101111",
  1986=>"101010000",
  1987=>"000111111",
  1988=>"001110011",
  1989=>"100101101",
  1990=>"111111100",
  1991=>"011100010",
  1992=>"011010110",
  1993=>"011100100",
  1994=>"101001111",
  1995=>"000010010",
  1996=>"000111001",
  1997=>"100000101",
  1998=>"001101000",
  1999=>"100010000",
  2000=>"111111110",
  2001=>"100010110",
  2002=>"101001000",
  2003=>"001000111",
  2004=>"111101001",
  2005=>"000101001",
  2006=>"011100000",
  2007=>"101101111",
  2008=>"000100001",
  2009=>"100000000",
  2010=>"010001001",
  2011=>"000010011",
  2012=>"101110101",
  2013=>"111111001",
  2014=>"101010100",
  2015=>"001001101",
  2016=>"010111111",
  2017=>"011111101",
  2018=>"111100100",
  2019=>"100110001",
  2020=>"000000000",
  2021=>"010100000",
  2022=>"101000111",
  2023=>"110110000",
  2024=>"100100001",
  2025=>"110000101",
  2026=>"010110001",
  2027=>"111001101",
  2028=>"111101101",
  2029=>"000001111",
  2030=>"111101011",
  2031=>"100100010",
  2032=>"000100101",
  2033=>"111110101",
  2034=>"100000111",
  2035=>"000101100",
  2036=>"001100011",
  2037=>"000111111",
  2038=>"111011110",
  2039=>"100010100",
  2040=>"010010100",
  2041=>"001110110",
  2042=>"001100100",
  2043=>"001101010",
  2044=>"001101101",
  2045=>"110101111",
  2046=>"110000100",
  2047=>"100100000",
  2048=>"111011111",
  2049=>"101001001",
  2050=>"001111110",
  2051=>"011110001",
  2052=>"110101111",
  2053=>"010100110",
  2054=>"011100010",
  2055=>"010010011",
  2056=>"111110110",
  2057=>"110100010",
  2058=>"001011111",
  2059=>"011010111",
  2060=>"000000100",
  2061=>"110001101",
  2062=>"000011101",
  2063=>"100101101",
  2064=>"100000100",
  2065=>"111110111",
  2066=>"111010110",
  2067=>"000101011",
  2068=>"000100101",
  2069=>"111011011",
  2070=>"000011011",
  2071=>"111001101",
  2072=>"110001110",
  2073=>"110101011",
  2074=>"011011000",
  2075=>"100110101",
  2076=>"000010110",
  2077=>"010000011",
  2078=>"010010000",
  2079=>"110000011",
  2080=>"000110100",
  2081=>"000100101",
  2082=>"010010010",
  2083=>"110100010",
  2084=>"110010101",
  2085=>"000110011",
  2086=>"001110100",
  2087=>"110111110",
  2088=>"011110011",
  2089=>"010001110",
  2090=>"111001000",
  2091=>"110011011",
  2092=>"010000100",
  2093=>"010110111",
  2094=>"001110100",
  2095=>"100010110",
  2096=>"111111010",
  2097=>"010100110",
  2098=>"110011010",
  2099=>"000101011",
  2100=>"101100000",
  2101=>"000000000",
  2102=>"000110000",
  2103=>"000000111",
  2104=>"101001010",
  2105=>"000011100",
  2106=>"001110110",
  2107=>"100000111",
  2108=>"100101010",
  2109=>"011110100",
  2110=>"101000001",
  2111=>"000100001",
  2112=>"110010111",
  2113=>"001001010",
  2114=>"011001100",
  2115=>"111100100",
  2116=>"100111101",
  2117=>"101111001",
  2118=>"010010001",
  2119=>"000101110",
  2120=>"101011011",
  2121=>"100111101",
  2122=>"000010000",
  2123=>"100001000",
  2124=>"101101110",
  2125=>"111000001",
  2126=>"110101101",
  2127=>"110001011",
  2128=>"101001101",
  2129=>"001010110",
  2130=>"011000001",
  2131=>"100111111",
  2132=>"010111100",
  2133=>"010001101",
  2134=>"011110001",
  2135=>"011111010",
  2136=>"110011000",
  2137=>"100101010",
  2138=>"101100100",
  2139=>"000001000",
  2140=>"111000111",
  2141=>"000011001",
  2142=>"110010001",
  2143=>"111010100",
  2144=>"001110111",
  2145=>"010000100",
  2146=>"010110100",
  2147=>"110011011",
  2148=>"000010001",
  2149=>"110111011",
  2150=>"001001101",
  2151=>"001010010",
  2152=>"110100110",
  2153=>"101111011",
  2154=>"000110000",
  2155=>"110010101",
  2156=>"101101110",
  2157=>"101100110",
  2158=>"010000001",
  2159=>"010110011",
  2160=>"100010111",
  2161=>"001000100",
  2162=>"101101101",
  2163=>"000111001",
  2164=>"110110010",
  2165=>"010111110",
  2166=>"100000100",
  2167=>"000100111",
  2168=>"011011010",
  2169=>"101000000",
  2170=>"011100000",
  2171=>"111001010",
  2172=>"100001101",
  2173=>"111111010",
  2174=>"010100010",
  2175=>"010000000",
  2176=>"001110101",
  2177=>"101110101",
  2178=>"110001010",
  2179=>"100001001",
  2180=>"001000000",
  2181=>"110101110",
  2182=>"011111100",
  2183=>"111000100",
  2184=>"111110101",
  2185=>"110100011",
  2186=>"010100000",
  2187=>"000000011",
  2188=>"011100111",
  2189=>"100110000",
  2190=>"011111111",
  2191=>"111101101",
  2192=>"101100001",
  2193=>"000111000",
  2194=>"000000111",
  2195=>"101000111",
  2196=>"100101101",
  2197=>"111110010",
  2198=>"010100101",
  2199=>"101101010",
  2200=>"110001100",
  2201=>"100010001",
  2202=>"011001100",
  2203=>"001011010",
  2204=>"010110011",
  2205=>"011111010",
  2206=>"100101110",
  2207=>"000010111",
  2208=>"110100101",
  2209=>"010100111",
  2210=>"010111000",
  2211=>"011101000",
  2212=>"110101110",
  2213=>"010001101",
  2214=>"001101100",
  2215=>"010010000",
  2216=>"000010110",
  2217=>"111011010",
  2218=>"010010101",
  2219=>"101010100",
  2220=>"100011010",
  2221=>"001000101",
  2222=>"001000001",
  2223=>"110010000",
  2224=>"100000111",
  2225=>"001001111",
  2226=>"100100101",
  2227=>"000000001",
  2228=>"101010011",
  2229=>"100101011",
  2230=>"010010000",
  2231=>"111001101",
  2232=>"100101101",
  2233=>"111010010",
  2234=>"000011110",
  2235=>"111011100",
  2236=>"001010110",
  2237=>"000010111",
  2238=>"111101011",
  2239=>"001110001",
  2240=>"001101110",
  2241=>"010001000",
  2242=>"111100010",
  2243=>"101011110",
  2244=>"111110111",
  2245=>"111110101",
  2246=>"010101010",
  2247=>"100101101",
  2248=>"111111110",
  2249=>"001110010",
  2250=>"111011000",
  2251=>"010110101",
  2252=>"001001101",
  2253=>"010100000",
  2254=>"011011111",
  2255=>"101100010",
  2256=>"000110011",
  2257=>"111010100",
  2258=>"111010000",
  2259=>"001100000",
  2260=>"011000000",
  2261=>"000110101",
  2262=>"100011001",
  2263=>"100111011",
  2264=>"111100111",
  2265=>"111100111",
  2266=>"000011010",
  2267=>"100110001",
  2268=>"100101010",
  2269=>"010101000",
  2270=>"000100101",
  2271=>"010100000",
  2272=>"100110010",
  2273=>"110001110",
  2274=>"110110100",
  2275=>"011100100",
  2276=>"101001011",
  2277=>"000100010",
  2278=>"011010111",
  2279=>"001101011",
  2280=>"100101011",
  2281=>"111110000",
  2282=>"101000010",
  2283=>"111010110",
  2284=>"000111011",
  2285=>"100010100",
  2286=>"000010000",
  2287=>"111001001",
  2288=>"010000001",
  2289=>"000101111",
  2290=>"100010111",
  2291=>"100110011",
  2292=>"011000011",
  2293=>"111011110",
  2294=>"000011110",
  2295=>"111001001",
  2296=>"100000101",
  2297=>"010111101",
  2298=>"101101011",
  2299=>"101010000",
  2300=>"011100010",
  2301=>"011101111",
  2302=>"110000000",
  2303=>"000100001",
  2304=>"111110000",
  2305=>"011010000",
  2306=>"100010010",
  2307=>"111010101",
  2308=>"110011011",
  2309=>"101100110",
  2310=>"001111000",
  2311=>"001000000",
  2312=>"000101000",
  2313=>"101101011",
  2314=>"100100000",
  2315=>"111110010",
  2316=>"111111101",
  2317=>"001001100",
  2318=>"101010110",
  2319=>"011011000",
  2320=>"110001000",
  2321=>"010011011",
  2322=>"000110101",
  2323=>"001101011",
  2324=>"110100001",
  2325=>"111011000",
  2326=>"001010000",
  2327=>"001100111",
  2328=>"010010111",
  2329=>"100110111",
  2330=>"010110000",
  2331=>"100100001",
  2332=>"000111010",
  2333=>"101010110",
  2334=>"010010101",
  2335=>"000010000",
  2336=>"011001011",
  2337=>"110110101",
  2338=>"000001000",
  2339=>"110101100",
  2340=>"110001011",
  2341=>"011000100",
  2342=>"010100000",
  2343=>"000010110",
  2344=>"100011001",
  2345=>"010101100",
  2346=>"000001110",
  2347=>"100001000",
  2348=>"110100100",
  2349=>"111111010",
  2350=>"000000100",
  2351=>"001100001",
  2352=>"000011111",
  2353=>"110011001",
  2354=>"110000101",
  2355=>"001001000",
  2356=>"001101000",
  2357=>"100100101",
  2358=>"101010010",
  2359=>"101101111",
  2360=>"010000101",
  2361=>"001001010",
  2362=>"010110001",
  2363=>"111110101",
  2364=>"000011010",
  2365=>"110011001",
  2366=>"000111101",
  2367=>"000001110",
  2368=>"000011111",
  2369=>"111001101",
  2370=>"000100110",
  2371=>"000100010",
  2372=>"101011011",
  2373=>"010110010",
  2374=>"011100110",
  2375=>"110010100",
  2376=>"001011110",
  2377=>"110011011",
  2378=>"001101101",
  2379=>"001110100",
  2380=>"010110110",
  2381=>"011100011",
  2382=>"011100001",
  2383=>"111101000",
  2384=>"101111100",
  2385=>"111011001",
  2386=>"110011011",
  2387=>"000010010",
  2388=>"001001011",
  2389=>"111111111",
  2390=>"100001101",
  2391=>"010010001",
  2392=>"100000001",
  2393=>"110100011",
  2394=>"110010010",
  2395=>"000001001",
  2396=>"100101010",
  2397=>"010101000",
  2398=>"010011110",
  2399=>"011011000",
  2400=>"011011111",
  2401=>"011110101",
  2402=>"010111000",
  2403=>"001000011",
  2404=>"100110000",
  2405=>"010100010",
  2406=>"000110000",
  2407=>"000000100",
  2408=>"000010111",
  2409=>"111001010",
  2410=>"101011000",
  2411=>"000101001",
  2412=>"011011000",
  2413=>"010010111",
  2414=>"101001001",
  2415=>"010000100",
  2416=>"101100100",
  2417=>"000010001",
  2418=>"000011011",
  2419=>"000111010",
  2420=>"110010000",
  2421=>"000001010",
  2422=>"010011010",
  2423=>"000001101",
  2424=>"001010100",
  2425=>"011110100",
  2426=>"111110110",
  2427=>"110010110",
  2428=>"110001010",
  2429=>"011100101",
  2430=>"100010101",
  2431=>"111110100",
  2432=>"100011110",
  2433=>"100011110",
  2434=>"100100010",
  2435=>"111011011",
  2436=>"000000100",
  2437=>"001100010",
  2438=>"000100001",
  2439=>"001110100",
  2440=>"111000101",
  2441=>"000111001",
  2442=>"111100011",
  2443=>"111111111",
  2444=>"010111011",
  2445=>"000100110",
  2446=>"000011110",
  2447=>"100101001",
  2448=>"000111101",
  2449=>"000001010",
  2450=>"010111100",
  2451=>"010111100",
  2452=>"000111000",
  2453=>"010011010",
  2454=>"101100111",
  2455=>"010011010",
  2456=>"000011011",
  2457=>"000010110",
  2458=>"101100111",
  2459=>"000011101",
  2460=>"001011101",
  2461=>"011011110",
  2462=>"100001010",
  2463=>"000111110",
  2464=>"000000100",
  2465=>"101111101",
  2466=>"011000101",
  2467=>"011000100",
  2468=>"111001001",
  2469=>"010101111",
  2470=>"100101000",
  2471=>"101001001",
  2472=>"011011011",
  2473=>"011011001",
  2474=>"000000010",
  2475=>"110101101",
  2476=>"001111111",
  2477=>"100110001",
  2478=>"011101111",
  2479=>"100110000",
  2480=>"100100011",
  2481=>"010001000",
  2482=>"100101011",
  2483=>"000010010",
  2484=>"010000011",
  2485=>"001000110",
  2486=>"001101101",
  2487=>"011100001",
  2488=>"010100111",
  2489=>"101101100",
  2490=>"101110010",
  2491=>"011010011",
  2492=>"100001100",
  2493=>"100111010",
  2494=>"111101000",
  2495=>"100111101",
  2496=>"000010100",
  2497=>"101010011",
  2498=>"110010000",
  2499=>"101011010",
  2500=>"010001001",
  2501=>"110100100",
  2502=>"001001110",
  2503=>"010001100",
  2504=>"001001111",
  2505=>"000001111",
  2506=>"000001010",
  2507=>"011001111",
  2508=>"011111010",
  2509=>"111011001",
  2510=>"011110001",
  2511=>"111110011",
  2512=>"011010011",
  2513=>"100001110",
  2514=>"010110010",
  2515=>"100111010",
  2516=>"010010000",
  2517=>"000100010",
  2518=>"001110000",
  2519=>"110000000",
  2520=>"000101011",
  2521=>"011010000",
  2522=>"000110010",
  2523=>"101001100",
  2524=>"111010001",
  2525=>"001110000",
  2526=>"011100111",
  2527=>"101100111",
  2528=>"000000001",
  2529=>"100110100",
  2530=>"101010010",
  2531=>"101001000",
  2532=>"111001101",
  2533=>"000010101",
  2534=>"100110000",
  2535=>"010110011",
  2536=>"000000000",
  2537=>"000011101",
  2538=>"000000000",
  2539=>"111001100",
  2540=>"110100010",
  2541=>"011100011",
  2542=>"000100011",
  2543=>"000001001",
  2544=>"111111111",
  2545=>"010110011",
  2546=>"010011000",
  2547=>"011011101",
  2548=>"110010011",
  2549=>"101010110",
  2550=>"101100010",
  2551=>"000110000",
  2552=>"011000111",
  2553=>"110001011",
  2554=>"000000010",
  2555=>"111100100",
  2556=>"110111000",
  2557=>"000000100",
  2558=>"010110010",
  2559=>"000100010",
  2560=>"110110100",
  2561=>"011001000",
  2562=>"100110011",
  2563=>"111111110",
  2564=>"010010001",
  2565=>"111011111",
  2566=>"110111000",
  2567=>"100001111",
  2568=>"110110011",
  2569=>"000010001",
  2570=>"011011010",
  2571=>"110010101",
  2572=>"101011111",
  2573=>"110010001",
  2574=>"111100111",
  2575=>"110011000",
  2576=>"110100111",
  2577=>"111110110",
  2578=>"101111100",
  2579=>"100100011",
  2580=>"010000101",
  2581=>"010010010",
  2582=>"101011111",
  2583=>"000110011",
  2584=>"010111101",
  2585=>"000001111",
  2586=>"000011101",
  2587=>"100001001",
  2588=>"001000111",
  2589=>"000101110",
  2590=>"000110001",
  2591=>"111101100",
  2592=>"111000101",
  2593=>"000010110",
  2594=>"010110100",
  2595=>"011111001",
  2596=>"111001010",
  2597=>"101001100",
  2598=>"001110100",
  2599=>"110100000",
  2600=>"110000011",
  2601=>"000100000",
  2602=>"011000111",
  2603=>"100000001",
  2604=>"000001110",
  2605=>"110100001",
  2606=>"101110000",
  2607=>"001010100",
  2608=>"010011100",
  2609=>"101111011",
  2610=>"001110100",
  2611=>"000100011",
  2612=>"100000010",
  2613=>"000001000",
  2614=>"001111010",
  2615=>"111110010",
  2616=>"100010001",
  2617=>"000111110",
  2618=>"010001011",
  2619=>"111111011",
  2620=>"011011011",
  2621=>"111100111",
  2622=>"010010111",
  2623=>"111000000",
  2624=>"011111111",
  2625=>"101011110",
  2626=>"000010000",
  2627=>"100100111",
  2628=>"111001111",
  2629=>"010110010",
  2630=>"000000001",
  2631=>"011100011",
  2632=>"010110110",
  2633=>"010000111",
  2634=>"011111100",
  2635=>"111110111",
  2636=>"101111111",
  2637=>"010111111",
  2638=>"110101111",
  2639=>"100110111",
  2640=>"001110110",
  2641=>"100000011",
  2642=>"110001101",
  2643=>"111110010",
  2644=>"001000100",
  2645=>"000101010",
  2646=>"100111101",
  2647=>"011110000",
  2648=>"011100111",
  2649=>"100100100",
  2650=>"100100111",
  2651=>"000110100",
  2652=>"110110010",
  2653=>"111001000",
  2654=>"001001001",
  2655=>"001110010",
  2656=>"011010101",
  2657=>"100010010",
  2658=>"101001010",
  2659=>"000000000",
  2660=>"001001110",
  2661=>"110010111",
  2662=>"001100011",
  2663=>"010101110",
  2664=>"000001111",
  2665=>"111111111",
  2666=>"001000001",
  2667=>"010110100",
  2668=>"111000100",
  2669=>"110100000",
  2670=>"010100111",
  2671=>"001011000",
  2672=>"100101000",
  2673=>"100010100",
  2674=>"111100000",
  2675=>"100110111",
  2676=>"101101000",
  2677=>"011000011",
  2678=>"001010010",
  2679=>"010000101",
  2680=>"110010111",
  2681=>"010001001",
  2682=>"100111010",
  2683=>"110011100",
  2684=>"110000110",
  2685=>"010101001",
  2686=>"001011100",
  2687=>"110000001",
  2688=>"000001100",
  2689=>"101011111",
  2690=>"011010111",
  2691=>"111011010",
  2692=>"010101000",
  2693=>"000100111",
  2694=>"110110011",
  2695=>"001100011",
  2696=>"100000100",
  2697=>"110101000",
  2698=>"000011000",
  2699=>"001001000",
  2700=>"000010011",
  2701=>"111100011",
  2702=>"110001111",
  2703=>"010000000",
  2704=>"010101010",
  2705=>"100011010",
  2706=>"010100011",
  2707=>"111010011",
  2708=>"001001011",
  2709=>"001000100",
  2710=>"001111101",
  2711=>"100100001",
  2712=>"010011101",
  2713=>"100000010",
  2714=>"100101110",
  2715=>"000111011",
  2716=>"000000010",
  2717=>"111110000",
  2718=>"011010110",
  2719=>"001000110",
  2720=>"111011000",
  2721=>"010010000",
  2722=>"011000001",
  2723=>"110110111",
  2724=>"000001101",
  2725=>"111110101",
  2726=>"101011010",
  2727=>"000000010",
  2728=>"100001010",
  2729=>"111011001",
  2730=>"101111010",
  2731=>"011010001",
  2732=>"100011101",
  2733=>"101110011",
  2734=>"011001001",
  2735=>"001100001",
  2736=>"100010001",
  2737=>"010010101",
  2738=>"111100100",
  2739=>"101101101",
  2740=>"000110010",
  2741=>"011100101",
  2742=>"111111101",
  2743=>"100001101",
  2744=>"000110010",
  2745=>"110101000",
  2746=>"001001000",
  2747=>"000111011",
  2748=>"001011110",
  2749=>"110001101",
  2750=>"100110011",
  2751=>"101011101",
  2752=>"111101111",
  2753=>"110011000",
  2754=>"100001000",
  2755=>"000110111",
  2756=>"110101110",
  2757=>"011010100",
  2758=>"111110010",
  2759=>"011001011",
  2760=>"000111110",
  2761=>"110011011",
  2762=>"000010011",
  2763=>"100101010",
  2764=>"001101100",
  2765=>"100110000",
  2766=>"111001000",
  2767=>"000011011",
  2768=>"111000001",
  2769=>"010011011",
  2770=>"000000010",
  2771=>"011111111",
  2772=>"100111111",
  2773=>"010011000",
  2774=>"111011111",
  2775=>"000101111",
  2776=>"010110010",
  2777=>"100010111",
  2778=>"110010110",
  2779=>"110110011",
  2780=>"010010110",
  2781=>"110100101",
  2782=>"011100010",
  2783=>"000100011",
  2784=>"000111111",
  2785=>"001001100",
  2786=>"100110000",
  2787=>"111000110",
  2788=>"100100111",
  2789=>"000000101",
  2790=>"110101001",
  2791=>"101111110",
  2792=>"011101000",
  2793=>"010011101",
  2794=>"110000001",
  2795=>"010110110",
  2796=>"110100111",
  2797=>"010001010",
  2798=>"000111001",
  2799=>"010001110",
  2800=>"111110110",
  2801=>"110101011",
  2802=>"110011001",
  2803=>"011000011",
  2804=>"110000000",
  2805=>"100100000",
  2806=>"110101010",
  2807=>"100010111",
  2808=>"001001001",
  2809=>"000100100",
  2810=>"110000001",
  2811=>"001100010",
  2812=>"000011001",
  2813=>"000001001",
  2814=>"110100001",
  2815=>"000111010",
  2816=>"101110110",
  2817=>"101010111",
  2818=>"001110000",
  2819=>"101000100",
  2820=>"001011100",
  2821=>"010110110",
  2822=>"110111111",
  2823=>"010010101",
  2824=>"101011110",
  2825=>"100100001",
  2826=>"101101101",
  2827=>"100100110",
  2828=>"011100100",
  2829=>"101110100",
  2830=>"101011110",
  2831=>"101001101",
  2832=>"010010010",
  2833=>"010101010",
  2834=>"001000001",
  2835=>"101101111",
  2836=>"010001110",
  2837=>"001101011",
  2838=>"111010100",
  2839=>"111111011",
  2840=>"011011100",
  2841=>"111001000",
  2842=>"000011000",
  2843=>"100011111",
  2844=>"111110000",
  2845=>"101011100",
  2846=>"001110000",
  2847=>"101110000",
  2848=>"110111001",
  2849=>"011110001",
  2850=>"110110000",
  2851=>"001100011",
  2852=>"001001110",
  2853=>"001010000",
  2854=>"010011010",
  2855=>"110001100",
  2856=>"001110111",
  2857=>"010010000",
  2858=>"000100000",
  2859=>"111100111",
  2860=>"001101001",
  2861=>"011110110",
  2862=>"100000100",
  2863=>"111011001",
  2864=>"110011000",
  2865=>"001111110",
  2866=>"111100100",
  2867=>"111010001",
  2868=>"100010000",
  2869=>"110011010",
  2870=>"101111001",
  2871=>"111001110",
  2872=>"011010000",
  2873=>"101011111",
  2874=>"001010110",
  2875=>"111011110",
  2876=>"001011101",
  2877=>"111111010",
  2878=>"010101110",
  2879=>"010110011",
  2880=>"011011110",
  2881=>"100101111",
  2882=>"110010111",
  2883=>"001110101",
  2884=>"011001000",
  2885=>"010111101",
  2886=>"110011011",
  2887=>"001001010",
  2888=>"010010011",
  2889=>"001111001",
  2890=>"000110101",
  2891=>"101110101",
  2892=>"111111000",
  2893=>"001111010",
  2894=>"101111001",
  2895=>"001011110",
  2896=>"100001100",
  2897=>"100111010",
  2898=>"011001011",
  2899=>"110100110",
  2900=>"111111010",
  2901=>"100010010",
  2902=>"101010101",
  2903=>"100111011",
  2904=>"110011001",
  2905=>"001101110",
  2906=>"011010001",
  2907=>"001110010",
  2908=>"001110010",
  2909=>"010110001",
  2910=>"001011101",
  2911=>"000001010",
  2912=>"000101011",
  2913=>"011100001",
  2914=>"000000110",
  2915=>"001111010",
  2916=>"010110100",
  2917=>"010100111",
  2918=>"000101010",
  2919=>"000001000",
  2920=>"011100111",
  2921=>"011010110",
  2922=>"111011101",
  2923=>"010011001",
  2924=>"111011001",
  2925=>"110101001",
  2926=>"111100111",
  2927=>"100110000",
  2928=>"001110010",
  2929=>"101111000",
  2930=>"100111100",
  2931=>"101000100",
  2932=>"100100110",
  2933=>"001011011",
  2934=>"100101001",
  2935=>"100110111",
  2936=>"001011111",
  2937=>"110111000",
  2938=>"101111111",
  2939=>"011010111",
  2940=>"001000010",
  2941=>"111001101",
  2942=>"101000111",
  2943=>"110111000",
  2944=>"000101001",
  2945=>"001011100",
  2946=>"110010110",
  2947=>"110101111",
  2948=>"100111011",
  2949=>"001101011",
  2950=>"110010010",
  2951=>"010011100",
  2952=>"111000011",
  2953=>"101000000",
  2954=>"110011000",
  2955=>"111100100",
  2956=>"100100010",
  2957=>"011100100",
  2958=>"100000110",
  2959=>"000000111",
  2960=>"001110000",
  2961=>"110001000",
  2962=>"111100011",
  2963=>"111100011",
  2964=>"001110001",
  2965=>"000001000",
  2966=>"110000100",
  2967=>"111110111",
  2968=>"000011111",
  2969=>"111010011",
  2970=>"000100111",
  2971=>"110101100",
  2972=>"001001000",
  2973=>"111000000",
  2974=>"010011001",
  2975=>"100110010",
  2976=>"011001110",
  2977=>"111000000",
  2978=>"000111110",
  2979=>"000100001",
  2980=>"001000100",
  2981=>"000001110",
  2982=>"100110100",
  2983=>"001101010",
  2984=>"011111000",
  2985=>"101110111",
  2986=>"110010111",
  2987=>"111110110",
  2988=>"100101111",
  2989=>"101101001",
  2990=>"010001111",
  2991=>"110101011",
  2992=>"100000011",
  2993=>"111000000",
  2994=>"111100000",
  2995=>"100010001",
  2996=>"111011101",
  2997=>"000001100",
  2998=>"100010000",
  2999=>"111111011",
  3000=>"010010111",
  3001=>"110110110",
  3002=>"111100110",
  3003=>"011011000",
  3004=>"110100101",
  3005=>"000010010",
  3006=>"100110111",
  3007=>"010001101",
  3008=>"101100010",
  3009=>"011110001",
  3010=>"010010001",
  3011=>"000100110",
  3012=>"011001010",
  3013=>"000110011",
  3014=>"000000000",
  3015=>"000111110",
  3016=>"110100111",
  3017=>"010001000",
  3018=>"110000010",
  3019=>"011011011",
  3020=>"001010101",
  3021=>"110110010",
  3022=>"110011101",
  3023=>"100010110",
  3024=>"011001111",
  3025=>"110111011",
  3026=>"111010111",
  3027=>"011101011",
  3028=>"110010110",
  3029=>"010101100",
  3030=>"010001000",
  3031=>"110010010",
  3032=>"101000001",
  3033=>"110001011",
  3034=>"001011110",
  3035=>"000000101",
  3036=>"001101100",
  3037=>"111111101",
  3038=>"111011011",
  3039=>"111111110",
  3040=>"011010010",
  3041=>"000101001",
  3042=>"010011101",
  3043=>"111101111",
  3044=>"110000010",
  3045=>"111100011",
  3046=>"000101100",
  3047=>"011110111",
  3048=>"001110001",
  3049=>"110011011",
  3050=>"001010110",
  3051=>"111010101",
  3052=>"101000110",
  3053=>"111011001",
  3054=>"010101000",
  3055=>"011011000",
  3056=>"000000010",
  3057=>"010100011",
  3058=>"101011110",
  3059=>"111101010",
  3060=>"111111010",
  3061=>"011110111",
  3062=>"010100000",
  3063=>"011001011",
  3064=>"110000111",
  3065=>"111100101",
  3066=>"111010000",
  3067=>"100000000",
  3068=>"000001110",
  3069=>"010010010",
  3070=>"010101000",
  3071=>"000111110",
  3072=>"111101000",
  3073=>"000110111",
  3074=>"110110000",
  3075=>"111111111",
  3076=>"101000000",
  3077=>"011001000",
  3078=>"101101101",
  3079=>"001111110",
  3080=>"000111010",
  3081=>"100011111",
  3082=>"111101000",
  3083=>"110000011",
  3084=>"011111111",
  3085=>"001001111",
  3086=>"101001001",
  3087=>"100110011",
  3088=>"010100110",
  3089=>"010100100",
  3090=>"011011100",
  3091=>"110110010",
  3092=>"010111111",
  3093=>"000110000",
  3094=>"011010110",
  3095=>"111001000",
  3096=>"100111001",
  3097=>"111111011",
  3098=>"100000100",
  3099=>"011100001",
  3100=>"110111010",
  3101=>"000110001",
  3102=>"011100001",
  3103=>"101000111",
  3104=>"001101101",
  3105=>"011111011",
  3106=>"101110101",
  3107=>"111101110",
  3108=>"001101101",
  3109=>"010000000",
  3110=>"110000100",
  3111=>"111111111",
  3112=>"101110001",
  3113=>"101001110",
  3114=>"010001010",
  3115=>"011000100",
  3116=>"010111110",
  3117=>"001011111",
  3118=>"100101100",
  3119=>"100100001",
  3120=>"010001111",
  3121=>"100011001",
  3122=>"000101101",
  3123=>"010111001",
  3124=>"000101010",
  3125=>"101110001",
  3126=>"101000001",
  3127=>"000010111",
  3128=>"111110111",
  3129=>"110000100",
  3130=>"011100100",
  3131=>"001011000",
  3132=>"010001001",
  3133=>"101001101",
  3134=>"000010001",
  3135=>"100011010",
  3136=>"101001000",
  3137=>"000011010",
  3138=>"110111110",
  3139=>"100000100",
  3140=>"111111010",
  3141=>"100100011",
  3142=>"100001001",
  3143=>"101010000",
  3144=>"100001101",
  3145=>"100001100",
  3146=>"011101011",
  3147=>"010111001",
  3148=>"110000110",
  3149=>"111010100",
  3150=>"111011011",
  3151=>"101101010",
  3152=>"000100001",
  3153=>"110100101",
  3154=>"110010111",
  3155=>"110001101",
  3156=>"110101100",
  3157=>"000111001",
  3158=>"000010010",
  3159=>"001101101",
  3160=>"110001011",
  3161=>"011011010",
  3162=>"000001110",
  3163=>"111111001",
  3164=>"101011010",
  3165=>"100100110",
  3166=>"100001011",
  3167=>"101110001",
  3168=>"011111101",
  3169=>"100100100",
  3170=>"111101011",
  3171=>"000101001",
  3172=>"011000100",
  3173=>"101000110",
  3174=>"000011001",
  3175=>"001110101",
  3176=>"010011011",
  3177=>"011101101",
  3178=>"001010000",
  3179=>"100100101",
  3180=>"011010111",
  3181=>"001110111",
  3182=>"010010111",
  3183=>"110001011",
  3184=>"100010100",
  3185=>"001101010",
  3186=>"100000000",
  3187=>"011101100",
  3188=>"011001000",
  3189=>"100010001",
  3190=>"000010001",
  3191=>"101101001",
  3192=>"001100100",
  3193=>"010101110",
  3194=>"111000100",
  3195=>"111101010",
  3196=>"111110110",
  3197=>"110001010",
  3198=>"111100110",
  3199=>"001100110",
  3200=>"110111010",
  3201=>"011101001",
  3202=>"101110000",
  3203=>"100100101",
  3204=>"110011001",
  3205=>"100000011",
  3206=>"001011000",
  3207=>"101000101",
  3208=>"001110101",
  3209=>"011111110",
  3210=>"100010101",
  3211=>"010110100",
  3212=>"000011110",
  3213=>"000000000",
  3214=>"101000000",
  3215=>"000011110",
  3216=>"101110010",
  3217=>"111010111",
  3218=>"011000100",
  3219=>"101011110",
  3220=>"001001011",
  3221=>"010110100",
  3222=>"011011111",
  3223=>"110011000",
  3224=>"101000100",
  3225=>"100000100",
  3226=>"101000011",
  3227=>"111110101",
  3228=>"000010111",
  3229=>"000001000",
  3230=>"101000001",
  3231=>"010010000",
  3232=>"101111111",
  3233=>"110010111",
  3234=>"100011001",
  3235=>"110100110",
  3236=>"011110011",
  3237=>"011001010",
  3238=>"001111000",
  3239=>"100101001",
  3240=>"100110010",
  3241=>"000100110",
  3242=>"100111011",
  3243=>"101101010",
  3244=>"000110110",
  3245=>"101100001",
  3246=>"100100010",
  3247=>"111011011",
  3248=>"001000110",
  3249=>"101101111",
  3250=>"010100010",
  3251=>"111101001",
  3252=>"001110000",
  3253=>"111111001",
  3254=>"011010111",
  3255=>"011000011",
  3256=>"000001011",
  3257=>"110110011",
  3258=>"110001001",
  3259=>"001011101",
  3260=>"111110110",
  3261=>"110101111",
  3262=>"110101100",
  3263=>"101111000",
  3264=>"101101110",
  3265=>"110010000",
  3266=>"101001001",
  3267=>"100110111",
  3268=>"001111010",
  3269=>"011101010",
  3270=>"111000100",
  3271=>"010100001",
  3272=>"101010100",
  3273=>"010101110",
  3274=>"101101100",
  3275=>"110111110",
  3276=>"100010011",
  3277=>"000101110",
  3278=>"011010110",
  3279=>"101000100",
  3280=>"011010100",
  3281=>"010111011",
  3282=>"100100100",
  3283=>"101111110",
  3284=>"000001001",
  3285=>"001011001",
  3286=>"110100100",
  3287=>"011111110",
  3288=>"100010110",
  3289=>"000010011",
  3290=>"110111100",
  3291=>"000111110",
  3292=>"100111001",
  3293=>"010011111",
  3294=>"100101111",
  3295=>"001110010",
  3296=>"100000001",
  3297=>"000000101",
  3298=>"110100010",
  3299=>"101011100",
  3300=>"111011000",
  3301=>"000000011",
  3302=>"101001100",
  3303=>"110100001",
  3304=>"011000101",
  3305=>"011010111",
  3306=>"111101001",
  3307=>"000011011",
  3308=>"100110010",
  3309=>"101011011",
  3310=>"100001111",
  3311=>"010011101",
  3312=>"100101101",
  3313=>"111001011",
  3314=>"111011100",
  3315=>"111011011",
  3316=>"010111001",
  3317=>"111100110",
  3318=>"000110010",
  3319=>"101101101",
  3320=>"111001001",
  3321=>"100111100",
  3322=>"111100100",
  3323=>"011000110",
  3324=>"000011111",
  3325=>"000111110",
  3326=>"110010111",
  3327=>"100010110",
  3328=>"101011101",
  3329=>"011011111",
  3330=>"100000101",
  3331=>"010101010",
  3332=>"001011110",
  3333=>"001100000",
  3334=>"111110111",
  3335=>"011100101",
  3336=>"010011010",
  3337=>"011100101",
  3338=>"010110100",
  3339=>"110000110",
  3340=>"011111001",
  3341=>"001000001",
  3342=>"110110000",
  3343=>"011000000",
  3344=>"011011001",
  3345=>"000001100",
  3346=>"100010101",
  3347=>"010101000",
  3348=>"100110100",
  3349=>"110011110",
  3350=>"011010001",
  3351=>"111001111",
  3352=>"111001001",
  3353=>"101000100",
  3354=>"100000110",
  3355=>"100001000",
  3356=>"010101110",
  3357=>"000000011",
  3358=>"000011101",
  3359=>"000010111",
  3360=>"101101010",
  3361=>"011110100",
  3362=>"010001100",
  3363=>"101110000",
  3364=>"000010001",
  3365=>"000101111",
  3366=>"110111100",
  3367=>"101000111",
  3368=>"100110101",
  3369=>"101100010",
  3370=>"110011111",
  3371=>"011011011",
  3372=>"000000111",
  3373=>"011010011",
  3374=>"011011111",
  3375=>"100001101",
  3376=>"001101000",
  3377=>"100001001",
  3378=>"001011000",
  3379=>"000001111",
  3380=>"000110100",
  3381=>"101011011",
  3382=>"100100011",
  3383=>"101111011",
  3384=>"000001110",
  3385=>"110110101",
  3386=>"010101000",
  3387=>"100111101",
  3388=>"101111110",
  3389=>"001110011",
  3390=>"111010000",
  3391=>"010000110",
  3392=>"011010011",
  3393=>"010010001",
  3394=>"110110110",
  3395=>"010011111",
  3396=>"000000100",
  3397=>"100111101",
  3398=>"101000000",
  3399=>"001000111",
  3400=>"101110001",
  3401=>"000110111",
  3402=>"101010110",
  3403=>"000000001",
  3404=>"000010100",
  3405=>"010110111",
  3406=>"111001011",
  3407=>"011000011",
  3408=>"100011001",
  3409=>"101110000",
  3410=>"110100100",
  3411=>"110111110",
  3412=>"011001011",
  3413=>"101000010",
  3414=>"011111100",
  3415=>"100010101",
  3416=>"111001001",
  3417=>"111100010",
  3418=>"010000110",
  3419=>"111101110",
  3420=>"111110010",
  3421=>"100100011",
  3422=>"100101001",
  3423=>"000001111",
  3424=>"001111101",
  3425=>"101111110",
  3426=>"011010100",
  3427=>"101101011",
  3428=>"001100011",
  3429=>"011000010",
  3430=>"010000001",
  3431=>"010111110",
  3432=>"101101011",
  3433=>"000110101",
  3434=>"011010010",
  3435=>"001000000",
  3436=>"110000000",
  3437=>"011110011",
  3438=>"100011010",
  3439=>"001100110",
  3440=>"111010000",
  3441=>"010010010",
  3442=>"100101111",
  3443=>"100101111",
  3444=>"010110111",
  3445=>"001100100",
  3446=>"111000101",
  3447=>"000000001",
  3448=>"011000111",
  3449=>"010100110",
  3450=>"100010111",
  3451=>"100110110",
  3452=>"000010001",
  3453=>"010011100",
  3454=>"000000001",
  3455=>"011100001",
  3456=>"110110000",
  3457=>"110001110",
  3458=>"011011001",
  3459=>"010001000",
  3460=>"100100010",
  3461=>"001001100",
  3462=>"111110111",
  3463=>"111001000",
  3464=>"000101100",
  3465=>"111100100",
  3466=>"100011111",
  3467=>"101110011",
  3468=>"111111100",
  3469=>"010011001",
  3470=>"111110010",
  3471=>"101011110",
  3472=>"111111010",
  3473=>"110110011",
  3474=>"000011011",
  3475=>"011000110",
  3476=>"001011000",
  3477=>"100101000",
  3478=>"010110010",
  3479=>"100110110",
  3480=>"001100110",
  3481=>"001101011",
  3482=>"000001111",
  3483=>"011000010",
  3484=>"010100101",
  3485=>"000101011",
  3486=>"011110000",
  3487=>"000110010",
  3488=>"000111001",
  3489=>"101000000",
  3490=>"011101111",
  3491=>"011001101",
  3492=>"101101011",
  3493=>"010101011",
  3494=>"000011101",
  3495=>"010000001",
  3496=>"000010110",
  3497=>"011010000",
  3498=>"000101000",
  3499=>"000000100",
  3500=>"110111111",
  3501=>"001001001",
  3502=>"000011100",
  3503=>"110011011",
  3504=>"000010011",
  3505=>"000001101",
  3506=>"011011010",
  3507=>"000011100",
  3508=>"000101000",
  3509=>"000100111",
  3510=>"101010010",
  3511=>"100010100",
  3512=>"010000111",
  3513=>"110111110",
  3514=>"011010010",
  3515=>"111110101",
  3516=>"010110010",
  3517=>"101101110",
  3518=>"010001100",
  3519=>"011110010",
  3520=>"010011000",
  3521=>"111011100",
  3522=>"110001111",
  3523=>"010010101",
  3524=>"000000000",
  3525=>"100000100",
  3526=>"001001000",
  3527=>"111100110",
  3528=>"000001000",
  3529=>"011101100",
  3530=>"000100110",
  3531=>"111011101",
  3532=>"001100000",
  3533=>"011000100",
  3534=>"111011111",
  3535=>"001101111",
  3536=>"001110001",
  3537=>"011000000",
  3538=>"011110010",
  3539=>"000100101",
  3540=>"010001110",
  3541=>"000100111",
  3542=>"111111110",
  3543=>"001010011",
  3544=>"010010101",
  3545=>"011110111",
  3546=>"000111010",
  3547=>"100000111",
  3548=>"010110110",
  3549=>"101000011",
  3550=>"111011110",
  3551=>"001010011",
  3552=>"010101101",
  3553=>"011011110",
  3554=>"110111110",
  3555=>"111101100",
  3556=>"011100001",
  3557=>"001000111",
  3558=>"000100101",
  3559=>"011111011",
  3560=>"001000010",
  3561=>"000011001",
  3562=>"101000000",
  3563=>"101011010",
  3564=>"001110111",
  3565=>"110011011",
  3566=>"111100110",
  3567=>"110100101",
  3568=>"001000111",
  3569=>"110111010",
  3570=>"101111010",
  3571=>"001011000",
  3572=>"011011000",
  3573=>"010111000",
  3574=>"010100010",
  3575=>"100110011",
  3576=>"001011000",
  3577=>"111010000",
  3578=>"111101010",
  3579=>"000111111",
  3580=>"101100011",
  3581=>"100001000",
  3582=>"000000100",
  3583=>"100011101",
  3584=>"111110000",
  3585=>"101001010",
  3586=>"111100100",
  3587=>"001010100",
  3588=>"001001001",
  3589=>"011000001",
  3590=>"100100111",
  3591=>"100011101",
  3592=>"100110001",
  3593=>"100110010",
  3594=>"001000000",
  3595=>"100111001",
  3596=>"101011111",
  3597=>"011110100",
  3598=>"001001100",
  3599=>"111100010",
  3600=>"111101101",
  3601=>"111110000",
  3602=>"100011100",
  3603=>"000000000",
  3604=>"110000000",
  3605=>"011101111",
  3606=>"101100010",
  3607=>"111010101",
  3608=>"101010101",
  3609=>"010111110",
  3610=>"011001000",
  3611=>"111111111",
  3612=>"101111011",
  3613=>"111101110",
  3614=>"001001110",
  3615=>"100001110",
  3616=>"111011010",
  3617=>"110001111",
  3618=>"000110100",
  3619=>"001011110",
  3620=>"111110011",
  3621=>"100010000",
  3622=>"111001000",
  3623=>"111001100",
  3624=>"111010001",
  3625=>"100010010",
  3626=>"001011001",
  3627=>"000001001",
  3628=>"111100101",
  3629=>"010001111",
  3630=>"010011101",
  3631=>"110001110",
  3632=>"111010100",
  3633=>"001101011",
  3634=>"001110000",
  3635=>"110110100",
  3636=>"100010011",
  3637=>"101000000",
  3638=>"100000111",
  3639=>"000000100",
  3640=>"001000010",
  3641=>"010001111",
  3642=>"101010100",
  3643=>"010101101",
  3644=>"100011110",
  3645=>"010100010",
  3646=>"100110010",
  3647=>"101111111",
  3648=>"100100100",
  3649=>"011100000",
  3650=>"000011000",
  3651=>"010101000",
  3652=>"001111010",
  3653=>"010110101",
  3654=>"000110011",
  3655=>"000001010",
  3656=>"110101111",
  3657=>"010000001",
  3658=>"001101010",
  3659=>"101001010",
  3660=>"011101101",
  3661=>"001010100",
  3662=>"111100100",
  3663=>"111110101",
  3664=>"000101100",
  3665=>"101010110",
  3666=>"001100001",
  3667=>"110000100",
  3668=>"011011101",
  3669=>"110001100",
  3670=>"001100001",
  3671=>"001000010",
  3672=>"000100110",
  3673=>"110111011",
  3674=>"110110001",
  3675=>"110111011",
  3676=>"001000100",
  3677=>"001111101",
  3678=>"000110110",
  3679=>"011010000",
  3680=>"110101100",
  3681=>"000000010",
  3682=>"110101111",
  3683=>"111111001",
  3684=>"110100110",
  3685=>"000110110",
  3686=>"110110000",
  3687=>"001101000",
  3688=>"011100011",
  3689=>"011101110",
  3690=>"100001100",
  3691=>"100110110",
  3692=>"110111110",
  3693=>"000010101",
  3694=>"100110010",
  3695=>"101101011",
  3696=>"000110111",
  3697=>"101001010",
  3698=>"000011001",
  3699=>"111111100",
  3700=>"000110000",
  3701=>"010110001",
  3702=>"000100000",
  3703=>"010100100",
  3704=>"001111111",
  3705=>"011010111",
  3706=>"001011110",
  3707=>"100011001",
  3708=>"000110100",
  3709=>"001100101",
  3710=>"100111000",
  3711=>"101000100",
  3712=>"110110111",
  3713=>"111100110",
  3714=>"110111100",
  3715=>"000000010",
  3716=>"100000110",
  3717=>"000010110",
  3718=>"010110000",
  3719=>"000000100",
  3720=>"000101001",
  3721=>"001011011",
  3722=>"001101110",
  3723=>"100001100",
  3724=>"111110101",
  3725=>"000110001",
  3726=>"110101100",
  3727=>"101100001",
  3728=>"010000000",
  3729=>"011100010",
  3730=>"111100011",
  3731=>"101010111",
  3732=>"111010101",
  3733=>"100011010",
  3734=>"010111100",
  3735=>"000101000",
  3736=>"100001111",
  3737=>"010000100",
  3738=>"010111110",
  3739=>"001101010",
  3740=>"001011101",
  3741=>"001011000",
  3742=>"010000001",
  3743=>"010011010",
  3744=>"111010011",
  3745=>"101001010",
  3746=>"100101110",
  3747=>"010101110",
  3748=>"100011000",
  3749=>"000000000",
  3750=>"100000011",
  3751=>"111001111",
  3752=>"001100100",
  3753=>"111101000",
  3754=>"110011011",
  3755=>"111111001",
  3756=>"010001000",
  3757=>"111110000",
  3758=>"001001111",
  3759=>"010011000",
  3760=>"000110011",
  3761=>"111100110",
  3762=>"100011010",
  3763=>"001101001",
  3764=>"111000000",
  3765=>"111011000",
  3766=>"100110001",
  3767=>"101110001",
  3768=>"110101001",
  3769=>"011110111",
  3770=>"101010001",
  3771=>"010000000",
  3772=>"011101100",
  3773=>"010110100",
  3774=>"101000111",
  3775=>"111001001",
  3776=>"011001111",
  3777=>"101101110",
  3778=>"110000010",
  3779=>"100110010",
  3780=>"000101001",
  3781=>"011100111",
  3782=>"100011110",
  3783=>"111000010",
  3784=>"011000101",
  3785=>"110010110",
  3786=>"111111011",
  3787=>"110110011",
  3788=>"000000000",
  3789=>"110000111",
  3790=>"101010111",
  3791=>"111110010",
  3792=>"001100101",
  3793=>"000011100",
  3794=>"111111000",
  3795=>"001110000",
  3796=>"100101110",
  3797=>"110111001",
  3798=>"001011011",
  3799=>"001011000",
  3800=>"000110000",
  3801=>"011110100",
  3802=>"111001111",
  3803=>"010110010",
  3804=>"111001111",
  3805=>"101100000",
  3806=>"110010001",
  3807=>"010101001",
  3808=>"111010011",
  3809=>"100010010",
  3810=>"000010000",
  3811=>"110110011",
  3812=>"110001100",
  3813=>"010000110",
  3814=>"001010101",
  3815=>"100101000",
  3816=>"111100011",
  3817=>"111011100",
  3818=>"111111100",
  3819=>"101000101",
  3820=>"001000100",
  3821=>"100000010",
  3822=>"111000110",
  3823=>"000011110",
  3824=>"010111101",
  3825=>"001000101",
  3826=>"110101000",
  3827=>"110101010",
  3828=>"101111111",
  3829=>"100110110",
  3830=>"010110110",
  3831=>"111011111",
  3832=>"000010000",
  3833=>"001111110",
  3834=>"101010011",
  3835=>"110010110",
  3836=>"001101111",
  3837=>"010001111",
  3838=>"011100011",
  3839=>"111010111",
  3840=>"100101010",
  3841=>"111011111",
  3842=>"110111011",
  3843=>"110011000",
  3844=>"001100001",
  3845=>"001100010",
  3846=>"000110111",
  3847=>"000010101",
  3848=>"011010110",
  3849=>"011010111",
  3850=>"101001000",
  3851=>"001101110",
  3852=>"111111100",
  3853=>"110110100",
  3854=>"110010101",
  3855=>"010101000",
  3856=>"000010111",
  3857=>"100111010",
  3858=>"011101011",
  3859=>"100100010",
  3860=>"101110110",
  3861=>"000111011",
  3862=>"111110010",
  3863=>"110100111",
  3864=>"111011001",
  3865=>"100100101",
  3866=>"000010011",
  3867=>"000000101",
  3868=>"100001101",
  3869=>"011011011",
  3870=>"111001100",
  3871=>"001010111",
  3872=>"011111110",
  3873=>"001000111",
  3874=>"111001010",
  3875=>"100000010",
  3876=>"101010010",
  3877=>"111000111",
  3878=>"110000001",
  3879=>"110110101",
  3880=>"001011010",
  3881=>"101101100",
  3882=>"001001110",
  3883=>"110111000",
  3884=>"111001011",
  3885=>"101000100",
  3886=>"000111001",
  3887=>"111010010",
  3888=>"010011111",
  3889=>"010000001",
  3890=>"000101100",
  3891=>"100010110",
  3892=>"011011000",
  3893=>"000001111",
  3894=>"000101110",
  3895=>"110101111",
  3896=>"011110101",
  3897=>"111011000",
  3898=>"011101101",
  3899=>"110101111",
  3900=>"111001110",
  3901=>"100000101",
  3902=>"011010101",
  3903=>"111101011",
  3904=>"101001100",
  3905=>"011000010",
  3906=>"100001000",
  3907=>"111111001",
  3908=>"010101010",
  3909=>"111110000",
  3910=>"101100010",
  3911=>"000000010",
  3912=>"101011111",
  3913=>"111110110",
  3914=>"110000001",
  3915=>"101101100",
  3916=>"110111010",
  3917=>"000001000",
  3918=>"110000100",
  3919=>"100100011",
  3920=>"101011010",
  3921=>"000010000",
  3922=>"111100000",
  3923=>"011000111",
  3924=>"101111001",
  3925=>"011101100",
  3926=>"101110111",
  3927=>"111100011",
  3928=>"001100101",
  3929=>"110010000",
  3930=>"101011001",
  3931=>"011011110",
  3932=>"111100110",
  3933=>"110001110",
  3934=>"111010001",
  3935=>"001110011",
  3936=>"110101000",
  3937=>"101000100",
  3938=>"010010101",
  3939=>"011100101",
  3940=>"100011111",
  3941=>"010100111",
  3942=>"010011010",
  3943=>"110111111",
  3944=>"100101010",
  3945=>"011101001",
  3946=>"000001101",
  3947=>"100000111",
  3948=>"110010010",
  3949=>"101000000",
  3950=>"111111100",
  3951=>"001101001",
  3952=>"000111111",
  3953=>"100110000",
  3954=>"001001011",
  3955=>"111100001",
  3956=>"111110101",
  3957=>"100110000",
  3958=>"000100110",
  3959=>"101111111",
  3960=>"000001100",
  3961=>"010111111",
  3962=>"100011001",
  3963=>"111101011",
  3964=>"001001010",
  3965=>"001100010",
  3966=>"010100100",
  3967=>"011110100",
  3968=>"110011011",
  3969=>"011000101",
  3970=>"100001001",
  3971=>"101000000",
  3972=>"101110101",
  3973=>"011011000",
  3974=>"101011011",
  3975=>"100001010",
  3976=>"010110111",
  3977=>"111110110",
  3978=>"110111111",
  3979=>"000100001",
  3980=>"010110101",
  3981=>"010111101",
  3982=>"000100000",
  3983=>"100001100",
  3984=>"101111000",
  3985=>"000111011",
  3986=>"100111000",
  3987=>"011111010",
  3988=>"011011100",
  3989=>"011010011",
  3990=>"011111101",
  3991=>"111011100",
  3992=>"110000001",
  3993=>"011110111",
  3994=>"000110100",
  3995=>"010110011",
  3996=>"001100001",
  3997=>"001001101",
  3998=>"001001100",
  3999=>"000000001",
  4000=>"011001111",
  4001=>"001000111",
  4002=>"111100000",
  4003=>"101100110",
  4004=>"000110111",
  4005=>"110100000",
  4006=>"011101111",
  4007=>"010111110",
  4008=>"010100001",
  4009=>"000011010",
  4010=>"000101111",
  4011=>"011110001",
  4012=>"011010000",
  4013=>"011010110",
  4014=>"000011000",
  4015=>"111100100",
  4016=>"011000010",
  4017=>"001110111",
  4018=>"111000101",
  4019=>"011011100",
  4020=>"011000010",
  4021=>"010010111",
  4022=>"101000010",
  4023=>"101110111",
  4024=>"010000100",
  4025=>"011110111",
  4026=>"000101010",
  4027=>"110110000",
  4028=>"110111011",
  4029=>"111011001",
  4030=>"101101111",
  4031=>"111000000",
  4032=>"010101000",
  4033=>"011011100",
  4034=>"000100100",
  4035=>"000111110",
  4036=>"000100100",
  4037=>"101111011",
  4038=>"101100010",
  4039=>"000010110",
  4040=>"001011100",
  4041=>"010010010",
  4042=>"010111101",
  4043=>"110010100",
  4044=>"111111110",
  4045=>"011100110",
  4046=>"111000110",
  4047=>"100010100",
  4048=>"110111100",
  4049=>"011110001",
  4050=>"010011010",
  4051=>"111000001",
  4052=>"011001110",
  4053=>"000000111",
  4054=>"001010010",
  4055=>"010010111",
  4056=>"110000001",
  4057=>"100001011",
  4058=>"010100000",
  4059=>"100011100",
  4060=>"101101011",
  4061=>"110000101",
  4062=>"110100100",
  4063=>"111110011",
  4064=>"110100011",
  4065=>"001001001",
  4066=>"100000110",
  4067=>"001100001",
  4068=>"101011000",
  4069=>"110001111",
  4070=>"100010100",
  4071=>"100010100",
  4072=>"100111000",
  4073=>"111011110",
  4074=>"111000010",
  4075=>"010001100",
  4076=>"101111100",
  4077=>"011110111",
  4078=>"011110011",
  4079=>"111011101",
  4080=>"000110010",
  4081=>"011110011",
  4082=>"001100100",
  4083=>"001111001",
  4084=>"111100100",
  4085=>"010011111",
  4086=>"000101000",
  4087=>"010101100",
  4088=>"000100100",
  4089=>"001010101",
  4090=>"001110001",
  4091=>"110110111",
  4092=>"001001011",
  4093=>"101010011",
  4094=>"110001001",
  4095=>"000110001",
  4096=>"010101000",
  4097=>"110111101",
  4098=>"111100000",
  4099=>"110010011",
  4100=>"100000111",
  4101=>"110011000",
  4102=>"000110001",
  4103=>"101001111",
  4104=>"111101000",
  4105=>"000111001",
  4106=>"011011111",
  4107=>"000010010",
  4108=>"100110100",
  4109=>"111011001",
  4110=>"111001111",
  4111=>"110000000",
  4112=>"110010111",
  4113=>"011001000",
  4114=>"001101101",
  4115=>"010000110",
  4116=>"110111110",
  4117=>"011010001",
  4118=>"100101101",
  4119=>"110000010",
  4120=>"101100110",
  4121=>"110111101",
  4122=>"101001011",
  4123=>"101111100",
  4124=>"010010101",
  4125=>"010101111",
  4126=>"100100010",
  4127=>"000000010",
  4128=>"000000001",
  4129=>"000111001",
  4130=>"110111110",
  4131=>"001111110",
  4132=>"010111110",
  4133=>"101010101",
  4134=>"100101111",
  4135=>"000111000",
  4136=>"101010100",
  4137=>"100000101",
  4138=>"100010111",
  4139=>"110000000",
  4140=>"000110101",
  4141=>"001101011",
  4142=>"001000011",
  4143=>"110101110",
  4144=>"111101110",
  4145=>"000011110",
  4146=>"011100001",
  4147=>"111011111",
  4148=>"101111000",
  4149=>"010000101",
  4150=>"001000000",
  4151=>"100101010",
  4152=>"010100100",
  4153=>"100001000",
  4154=>"111101001",
  4155=>"001101101",
  4156=>"111010000",
  4157=>"101111011",
  4158=>"000100111",
  4159=>"011001000",
  4160=>"010001011",
  4161=>"101101100",
  4162=>"010101100",
  4163=>"101101010",
  4164=>"010110100",
  4165=>"110100110",
  4166=>"110100101",
  4167=>"000111111",
  4168=>"111001011",
  4169=>"001000001",
  4170=>"110001111",
  4171=>"111100100",
  4172=>"011001111",
  4173=>"001100001",
  4174=>"111101000",
  4175=>"011001001",
  4176=>"111011011",
  4177=>"000101000",
  4178=>"100101110",
  4179=>"000001101",
  4180=>"111000110",
  4181=>"010010111",
  4182=>"011110100",
  4183=>"111100010",
  4184=>"100110001",
  4185=>"011010100",
  4186=>"100100111",
  4187=>"100001000",
  4188=>"000000001",
  4189=>"100101001",
  4190=>"011111111",
  4191=>"001110011",
  4192=>"000111001",
  4193=>"000100001",
  4194=>"010100111",
  4195=>"111001111",
  4196=>"001110001",
  4197=>"011010011",
  4198=>"100100110",
  4199=>"000001010",
  4200=>"101111110",
  4201=>"001100001",
  4202=>"010100111",
  4203=>"111000111",
  4204=>"111110101",
  4205=>"111110111",
  4206=>"110001100",
  4207=>"001000101",
  4208=>"010111001",
  4209=>"100001111",
  4210=>"110110011",
  4211=>"011011010",
  4212=>"001001110",
  4213=>"001010111",
  4214=>"110010000",
  4215=>"101010010",
  4216=>"101110111",
  4217=>"100101001",
  4218=>"111111110",
  4219=>"010000000",
  4220=>"000110000",
  4221=>"010011010",
  4222=>"100100101",
  4223=>"111111100",
  4224=>"110011010",
  4225=>"010110101",
  4226=>"100101100",
  4227=>"101111101",
  4228=>"111111100",
  4229=>"110000011",
  4230=>"111001001",
  4231=>"101110001",
  4232=>"111110111",
  4233=>"001101001",
  4234=>"110110100",
  4235=>"111101010",
  4236=>"111110000",
  4237=>"111100101",
  4238=>"111010100",
  4239=>"010011001",
  4240=>"000000110",
  4241=>"011111111",
  4242=>"000101100",
  4243=>"001001010",
  4244=>"010111111",
  4245=>"111111101",
  4246=>"100000001",
  4247=>"001110100",
  4248=>"111010110",
  4249=>"100101100",
  4250=>"010101110",
  4251=>"111111110",
  4252=>"000001011",
  4253=>"001011100",
  4254=>"000010111",
  4255=>"000001111",
  4256=>"101110111",
  4257=>"010111010",
  4258=>"010011100",
  4259=>"101000000",
  4260=>"000111101",
  4261=>"100111111",
  4262=>"010100110",
  4263=>"010010001",
  4264=>"111011010",
  4265=>"010001010",
  4266=>"101101101",
  4267=>"010101101",
  4268=>"010101101",
  4269=>"101010000",
  4270=>"101001111",
  4271=>"101010000",
  4272=>"001001001",
  4273=>"100100011",
  4274=>"100101011",
  4275=>"101110110",
  4276=>"101001001",
  4277=>"000001111",
  4278=>"001011111",
  4279=>"101011110",
  4280=>"000010101",
  4281=>"110100000",
  4282=>"101110101",
  4283=>"011100100",
  4284=>"010110010",
  4285=>"111011001",
  4286=>"011000010",
  4287=>"111111110",
  4288=>"100001101",
  4289=>"101011011",
  4290=>"101100101",
  4291=>"001111101",
  4292=>"100011001",
  4293=>"001011110",
  4294=>"110110110",
  4295=>"110111110",
  4296=>"001001001",
  4297=>"001000101",
  4298=>"110101000",
  4299=>"000011011",
  4300=>"000101111",
  4301=>"001011110",
  4302=>"001100111",
  4303=>"010011110",
  4304=>"001011111",
  4305=>"001110101",
  4306=>"101110110",
  4307=>"010001000",
  4308=>"000111100",
  4309=>"001100011",
  4310=>"101111101",
  4311=>"011111110",
  4312=>"011111101",
  4313=>"011100111",
  4314=>"110001111",
  4315=>"000101000",
  4316=>"101000101",
  4317=>"010110010",
  4318=>"011110011",
  4319=>"100010000",
  4320=>"100000101",
  4321=>"000011010",
  4322=>"011011001",
  4323=>"000100101",
  4324=>"011010010",
  4325=>"111001000",
  4326=>"100101001",
  4327=>"100010011",
  4328=>"100101110",
  4329=>"010010100",
  4330=>"110111001",
  4331=>"000100110",
  4332=>"111111010",
  4333=>"111110010",
  4334=>"110010100",
  4335=>"100001100",
  4336=>"000111001",
  4337=>"000101001",
  4338=>"100110010",
  4339=>"011111101",
  4340=>"001011010",
  4341=>"001111011",
  4342=>"001101110",
  4343=>"000100010",
  4344=>"100111011",
  4345=>"010001111",
  4346=>"010001110",
  4347=>"000101000",
  4348=>"101000101",
  4349=>"001000100",
  4350=>"010111111",
  4351=>"101101111",
  4352=>"000100101",
  4353=>"111000111",
  4354=>"000011111",
  4355=>"000000001",
  4356=>"000101100",
  4357=>"011100010",
  4358=>"100100111",
  4359=>"010101101",
  4360=>"111111110",
  4361=>"011011000",
  4362=>"001111011",
  4363=>"100000000",
  4364=>"011000010",
  4365=>"001000101",
  4366=>"010011001",
  4367=>"101001010",
  4368=>"100000011",
  4369=>"010001000",
  4370=>"010101010",
  4371=>"100010000",
  4372=>"101011111",
  4373=>"000101100",
  4374=>"101101101",
  4375=>"101000011",
  4376=>"101111101",
  4377=>"111100101",
  4378=>"010010101",
  4379=>"100100111",
  4380=>"011001000",
  4381=>"011110000",
  4382=>"110111111",
  4383=>"101110110",
  4384=>"110100001",
  4385=>"010001111",
  4386=>"100000000",
  4387=>"011101001",
  4388=>"000011001",
  4389=>"011111000",
  4390=>"100100110",
  4391=>"011011111",
  4392=>"010010110",
  4393=>"100010010",
  4394=>"110000110",
  4395=>"110010111",
  4396=>"011011111",
  4397=>"100010000",
  4398=>"001010001",
  4399=>"111101010",
  4400=>"100100010",
  4401=>"001011001",
  4402=>"111001001",
  4403=>"010011100",
  4404=>"111010111",
  4405=>"101010100",
  4406=>"010111000",
  4407=>"011010010",
  4408=>"010001000",
  4409=>"101010000",
  4410=>"000011011",
  4411=>"000110010",
  4412=>"101111101",
  4413=>"111010000",
  4414=>"100000110",
  4415=>"111011100",
  4416=>"101100100",
  4417=>"100101111",
  4418=>"001110011",
  4419=>"110100110",
  4420=>"000001101",
  4421=>"000100010",
  4422=>"110001100",
  4423=>"000001110",
  4424=>"110010111",
  4425=>"010000000",
  4426=>"011011100",
  4427=>"001000111",
  4428=>"100000101",
  4429=>"101001011",
  4430=>"000010010",
  4431=>"011010010",
  4432=>"011111100",
  4433=>"001111111",
  4434=>"000001000",
  4435=>"110110111",
  4436=>"100100001",
  4437=>"001101000",
  4438=>"011000100",
  4439=>"011110100",
  4440=>"000000010",
  4441=>"100001111",
  4442=>"110011011",
  4443=>"010111000",
  4444=>"100100100",
  4445=>"100101101",
  4446=>"000011001",
  4447=>"010000001",
  4448=>"100011101",
  4449=>"010100100",
  4450=>"100001010",
  4451=>"000110000",
  4452=>"100011011",
  4453=>"110001110",
  4454=>"000010110",
  4455=>"010001010",
  4456=>"111110101",
  4457=>"100111110",
  4458=>"011010010",
  4459=>"101101010",
  4460=>"111110001",
  4461=>"001111011",
  4462=>"000100111",
  4463=>"001111110",
  4464=>"110110101",
  4465=>"011111111",
  4466=>"000001100",
  4467=>"110110101",
  4468=>"100000000",
  4469=>"101111010",
  4470=>"100010001",
  4471=>"100100111",
  4472=>"111111101",
  4473=>"000101100",
  4474=>"011100110",
  4475=>"111111111",
  4476=>"001110110",
  4477=>"001001100",
  4478=>"010110111",
  4479=>"001100101",
  4480=>"100011011",
  4481=>"011011100",
  4482=>"110000001",
  4483=>"011011011",
  4484=>"101100111",
  4485=>"011100110",
  4486=>"111010011",
  4487=>"001111010",
  4488=>"100101101",
  4489=>"110011100",
  4490=>"100000101",
  4491=>"000000001",
  4492=>"001101000",
  4493=>"010101111",
  4494=>"000101000",
  4495=>"010111111",
  4496=>"111111000",
  4497=>"110100010",
  4498=>"011011100",
  4499=>"001010010",
  4500=>"111111111",
  4501=>"100011010",
  4502=>"101011011",
  4503=>"111110010",
  4504=>"101001101",
  4505=>"100001101",
  4506=>"110000000",
  4507=>"010110100",
  4508=>"001010011",
  4509=>"010010101",
  4510=>"110100111",
  4511=>"010100100",
  4512=>"010101100",
  4513=>"101111100",
  4514=>"110111101",
  4515=>"001001000",
  4516=>"011101100",
  4517=>"011110011",
  4518=>"100100111",
  4519=>"011110110",
  4520=>"010110101",
  4521=>"110111000",
  4522=>"101000100",
  4523=>"000001001",
  4524=>"100101100",
  4525=>"101111111",
  4526=>"001110111",
  4527=>"100000011",
  4528=>"011001000",
  4529=>"111110101",
  4530=>"101010101",
  4531=>"000010100",
  4532=>"101000010",
  4533=>"000011000",
  4534=>"110000001",
  4535=>"101110101",
  4536=>"110111010",
  4537=>"000100000",
  4538=>"000000000",
  4539=>"011101101",
  4540=>"000010101",
  4541=>"011101101",
  4542=>"000111100",
  4543=>"100100011",
  4544=>"010010100",
  4545=>"000000000",
  4546=>"010100011",
  4547=>"011001111",
  4548=>"111000001",
  4549=>"110110000",
  4550=>"110000011",
  4551=>"111100100",
  4552=>"010000001",
  4553=>"000100101",
  4554=>"100011100",
  4555=>"011000101",
  4556=>"110100101",
  4557=>"010011101",
  4558=>"101101111",
  4559=>"000100010",
  4560=>"110000010",
  4561=>"000111100",
  4562=>"001001111",
  4563=>"010010010",
  4564=>"111101101",
  4565=>"011101011",
  4566=>"111111100",
  4567=>"110011100",
  4568=>"000110111",
  4569=>"000000010",
  4570=>"101001001",
  4571=>"001001001",
  4572=>"011100001",
  4573=>"101101110",
  4574=>"011011011",
  4575=>"001111111",
  4576=>"010111110",
  4577=>"011101000",
  4578=>"000100000",
  4579=>"011011010",
  4580=>"001101111",
  4581=>"000001011",
  4582=>"101101101",
  4583=>"110100110",
  4584=>"010110110",
  4585=>"100010110",
  4586=>"111100110",
  4587=>"100001001",
  4588=>"100110110",
  4589=>"010100000",
  4590=>"110011110",
  4591=>"101011100",
  4592=>"100011000",
  4593=>"110000111",
  4594=>"110101011",
  4595=>"110011010",
  4596=>"010000111",
  4597=>"111000110",
  4598=>"001001101",
  4599=>"010110001",
  4600=>"111100011",
  4601=>"111111111",
  4602=>"101100000",
  4603=>"000000110",
  4604=>"101011100",
  4605=>"000110110",
  4606=>"100011010",
  4607=>"110100111",
  4608=>"011101011",
  4609=>"101101000",
  4610=>"011011000",
  4611=>"100101001",
  4612=>"111100001",
  4613=>"000110101",
  4614=>"000100111",
  4615=>"110110000",
  4616=>"111000100",
  4617=>"010001010",
  4618=>"111101011",
  4619=>"010111100",
  4620=>"110101000",
  4621=>"001000010",
  4622=>"000001011",
  4623=>"001011111",
  4624=>"000011000",
  4625=>"110110011",
  4626=>"100000010",
  4627=>"100111001",
  4628=>"101010000",
  4629=>"110000111",
  4630=>"001000111",
  4631=>"111111110",
  4632=>"001000101",
  4633=>"111111001",
  4634=>"111010110",
  4635=>"110011111",
  4636=>"001011101",
  4637=>"011001101",
  4638=>"010011111",
  4639=>"010101101",
  4640=>"010000000",
  4641=>"100000101",
  4642=>"110000110",
  4643=>"100000101",
  4644=>"101001011",
  4645=>"110010100",
  4646=>"100101111",
  4647=>"000100110",
  4648=>"100000011",
  4649=>"100000101",
  4650=>"000001100",
  4651=>"011001000",
  4652=>"010011001",
  4653=>"111001001",
  4654=>"000000000",
  4655=>"011011101",
  4656=>"111001001",
  4657=>"110010101",
  4658=>"010111111",
  4659=>"001110111",
  4660=>"001111101",
  4661=>"010101111",
  4662=>"100000010",
  4663=>"101000101",
  4664=>"101001101",
  4665=>"001111101",
  4666=>"001010011",
  4667=>"011111110",
  4668=>"001011110",
  4669=>"100001010",
  4670=>"010110001",
  4671=>"000111001",
  4672=>"000000001",
  4673=>"111010111",
  4674=>"111011110",
  4675=>"110000001",
  4676=>"011111111",
  4677=>"111100101",
  4678=>"000101110",
  4679=>"001010111",
  4680=>"011110101",
  4681=>"101101101",
  4682=>"101001100",
  4683=>"011011110",
  4684=>"010101110",
  4685=>"110000111",
  4686=>"110010110",
  4687=>"111110010",
  4688=>"000001011",
  4689=>"100101101",
  4690=>"110111111",
  4691=>"010101001",
  4692=>"010000100",
  4693=>"101001000",
  4694=>"001101101",
  4695=>"011010010",
  4696=>"100001101",
  4697=>"110111001",
  4698=>"100110100",
  4699=>"111000110",
  4700=>"010001000",
  4701=>"001001001",
  4702=>"111110111",
  4703=>"101101000",
  4704=>"000011010",
  4705=>"000111000",
  4706=>"001010010",
  4707=>"111111101",
  4708=>"110110110",
  4709=>"111111101",
  4710=>"100000110",
  4711=>"010101100",
  4712=>"010000000",
  4713=>"000111010",
  4714=>"001010011",
  4715=>"111110101",
  4716=>"010000111",
  4717=>"111001100",
  4718=>"111101010",
  4719=>"110101110",
  4720=>"101101101",
  4721=>"010011001",
  4722=>"111000011",
  4723=>"010001001",
  4724=>"010010001",
  4725=>"110101010",
  4726=>"100011110",
  4727=>"000011011",
  4728=>"110111100",
  4729=>"111010000",
  4730=>"010001000",
  4731=>"011001010",
  4732=>"111111111",
  4733=>"101001101",
  4734=>"111101101",
  4735=>"101001010",
  4736=>"010111111",
  4737=>"011110111",
  4738=>"011101110",
  4739=>"010111011",
  4740=>"100101110",
  4741=>"011100000",
  4742=>"001011111",
  4743=>"010101111",
  4744=>"011100111",
  4745=>"000011000",
  4746=>"011111011",
  4747=>"101010011",
  4748=>"011111000",
  4749=>"110010111",
  4750=>"101011100",
  4751=>"001010000",
  4752=>"011111010",
  4753=>"000010100",
  4754=>"010101101",
  4755=>"111001110",
  4756=>"111000000",
  4757=>"010000110",
  4758=>"111101110",
  4759=>"111111111",
  4760=>"111001011",
  4761=>"111010011",
  4762=>"011001001",
  4763=>"110110100",
  4764=>"000100000",
  4765=>"100011010",
  4766=>"110010100",
  4767=>"110011011",
  4768=>"110101100",
  4769=>"101100000",
  4770=>"011010110",
  4771=>"010100110",
  4772=>"111111000",
  4773=>"100010001",
  4774=>"100110110",
  4775=>"010000011",
  4776=>"000001110",
  4777=>"010001001",
  4778=>"101100001",
  4779=>"000110001",
  4780=>"010000000",
  4781=>"110000101",
  4782=>"001111011",
  4783=>"110100110",
  4784=>"000011100",
  4785=>"100000110",
  4786=>"101110101",
  4787=>"100100010",
  4788=>"001001011",
  4789=>"111011101",
  4790=>"000110111",
  4791=>"000001100",
  4792=>"010011110",
  4793=>"111011011",
  4794=>"000111001",
  4795=>"000101111",
  4796=>"000101101",
  4797=>"000010111",
  4798=>"111101110",
  4799=>"100011010",
  4800=>"000011111",
  4801=>"110000010",
  4802=>"000001101",
  4803=>"000111010",
  4804=>"000111000",
  4805=>"101100000",
  4806=>"110001100",
  4807=>"000101101",
  4808=>"111100001",
  4809=>"100001110",
  4810=>"100010001",
  4811=>"100011001",
  4812=>"101000100",
  4813=>"001010111",
  4814=>"000100000",
  4815=>"101101111",
  4816=>"101111001",
  4817=>"110001111",
  4818=>"010011111",
  4819=>"001001010",
  4820=>"011111001",
  4821=>"011111010",
  4822=>"001110100",
  4823=>"000111111",
  4824=>"111010010",
  4825=>"000101101",
  4826=>"111000010",
  4827=>"001101011",
  4828=>"111101101",
  4829=>"011101111",
  4830=>"110111010",
  4831=>"001111000",
  4832=>"110110101",
  4833=>"000010110",
  4834=>"111111111",
  4835=>"111011100",
  4836=>"100010111",
  4837=>"100110110",
  4838=>"101011000",
  4839=>"111111111",
  4840=>"100100000",
  4841=>"001010001",
  4842=>"111011100",
  4843=>"110011001",
  4844=>"000111100",
  4845=>"000010011",
  4846=>"110011000",
  4847=>"111100101",
  4848=>"010100010",
  4849=>"010011001",
  4850=>"001111111",
  4851=>"111111101",
  4852=>"100011000",
  4853=>"111111111",
  4854=>"000111101",
  4855=>"001000100",
  4856=>"000101001",
  4857=>"110010101",
  4858=>"010000000",
  4859=>"111100110",
  4860=>"100001110",
  4861=>"101011101",
  4862=>"001110000",
  4863=>"000010100",
  4864=>"100000110",
  4865=>"000010100",
  4866=>"010110010",
  4867=>"110101111",
  4868=>"001100000",
  4869=>"010000000",
  4870=>"100110010",
  4871=>"111111111",
  4872=>"101001111",
  4873=>"100110011",
  4874=>"010111111",
  4875=>"001101100",
  4876=>"011001001",
  4877=>"100010000",
  4878=>"001101100",
  4879=>"110101010",
  4880=>"010111110",
  4881=>"101101100",
  4882=>"011001101",
  4883=>"110010111",
  4884=>"010000000",
  4885=>"000010001",
  4886=>"101100001",
  4887=>"011010001",
  4888=>"000100010",
  4889=>"111111001",
  4890=>"011100011",
  4891=>"011000010",
  4892=>"110111111",
  4893=>"100110110",
  4894=>"100110110",
  4895=>"000101101",
  4896=>"101100011",
  4897=>"000011111",
  4898=>"111011011",
  4899=>"111010001",
  4900=>"000001011",
  4901=>"010110110",
  4902=>"111000011",
  4903=>"110011100",
  4904=>"100001101",
  4905=>"111010111",
  4906=>"000000000",
  4907=>"000011010",
  4908=>"000110011",
  4909=>"001010100",
  4910=>"101001010",
  4911=>"000101100",
  4912=>"001110100",
  4913=>"110011110",
  4914=>"100000111",
  4915=>"011010000",
  4916=>"000100100",
  4917=>"101010111",
  4918=>"000101010",
  4919=>"111111101",
  4920=>"000010000",
  4921=>"010010011",
  4922=>"000110011",
  4923=>"111111111",
  4924=>"000110000",
  4925=>"111000011",
  4926=>"011010101",
  4927=>"001111100",
  4928=>"111101111",
  4929=>"110110001",
  4930=>"100111001",
  4931=>"010111110",
  4932=>"001101010",
  4933=>"010100010",
  4934=>"000100110",
  4935=>"111100100",
  4936=>"001001100",
  4937=>"110110001",
  4938=>"011000000",
  4939=>"011100010",
  4940=>"111001010",
  4941=>"001011100",
  4942=>"101001011",
  4943=>"001010011",
  4944=>"001101000",
  4945=>"100110000",
  4946=>"100100010",
  4947=>"100100011",
  4948=>"011000100",
  4949=>"010010001",
  4950=>"111111110",
  4951=>"111010001",
  4952=>"010000101",
  4953=>"010000000",
  4954=>"011000010",
  4955=>"000000110",
  4956=>"101111011",
  4957=>"000101010",
  4958=>"110000111",
  4959=>"110011100",
  4960=>"100010011",
  4961=>"010111000",
  4962=>"110010001",
  4963=>"111000011",
  4964=>"101100010",
  4965=>"111100100",
  4966=>"110111110",
  4967=>"111010101",
  4968=>"010111011",
  4969=>"000010000",
  4970=>"011100110",
  4971=>"110001111",
  4972=>"101101111",
  4973=>"100100101",
  4974=>"000010101",
  4975=>"001011100",
  4976=>"001000001",
  4977=>"001110000",
  4978=>"110001101",
  4979=>"010000010",
  4980=>"011100100",
  4981=>"000010101",
  4982=>"000110100",
  4983=>"001011011",
  4984=>"110111010",
  4985=>"101011100",
  4986=>"000001011",
  4987=>"100110111",
  4988=>"001010001",
  4989=>"110000111",
  4990=>"110000101",
  4991=>"100111010",
  4992=>"010010111",
  4993=>"101011110",
  4994=>"101011101",
  4995=>"011100100",
  4996=>"011101011",
  4997=>"101101001",
  4998=>"111000110",
  4999=>"111010011",
  5000=>"000111011",
  5001=>"001011111",
  5002=>"010101011",
  5003=>"000000100",
  5004=>"010010010",
  5005=>"001011000",
  5006=>"011100100",
  5007=>"000110101",
  5008=>"101100101",
  5009=>"101100100",
  5010=>"100101010",
  5011=>"011011011",
  5012=>"001001001",
  5013=>"100100010",
  5014=>"001001111",
  5015=>"100101000",
  5016=>"100111101",
  5017=>"101100101",
  5018=>"100001111",
  5019=>"111111100",
  5020=>"010110111",
  5021=>"100011111",
  5022=>"010000101",
  5023=>"001011110",
  5024=>"001110100",
  5025=>"000010101",
  5026=>"010010000",
  5027=>"111101111",
  5028=>"111101000",
  5029=>"011010010",
  5030=>"010110010",
  5031=>"100100010",
  5032=>"111000101",
  5033=>"111011000",
  5034=>"110110011",
  5035=>"000010101",
  5036=>"001000000",
  5037=>"111000111",
  5038=>"001101001",
  5039=>"000110100",
  5040=>"100001111",
  5041=>"101101110",
  5042=>"001101111",
  5043=>"001001000",
  5044=>"001000010",
  5045=>"000000101",
  5046=>"101001010",
  5047=>"011011101",
  5048=>"101001100",
  5049=>"010111010",
  5050=>"011011100",
  5051=>"000100000",
  5052=>"011001010",
  5053=>"010011001",
  5054=>"010100000",
  5055=>"111101101",
  5056=>"000010000",
  5057=>"000010000",
  5058=>"100111011",
  5059=>"100100010",
  5060=>"100110011",
  5061=>"100111000",
  5062=>"010010101",
  5063=>"110101000",
  5064=>"100001100",
  5065=>"110111101",
  5066=>"011111111",
  5067=>"010101011",
  5068=>"110101100",
  5069=>"100011111",
  5070=>"111000011",
  5071=>"010000010",
  5072=>"101011000",
  5073=>"001010000",
  5074=>"011000000",
  5075=>"111000000",
  5076=>"011011001",
  5077=>"100010010",
  5078=>"110001101",
  5079=>"110101101",
  5080=>"011010001",
  5081=>"001000100",
  5082=>"101111111",
  5083=>"111001001",
  5084=>"111111000",
  5085=>"100010100",
  5086=>"100011001",
  5087=>"010101010",
  5088=>"101110110",
  5089=>"100100100",
  5090=>"100100100",
  5091=>"010100101",
  5092=>"111010100",
  5093=>"100101010",
  5094=>"000010111",
  5095=>"111111110",
  5096=>"111100000",
  5097=>"001000110",
  5098=>"100001010",
  5099=>"101011110",
  5100=>"000001011",
  5101=>"101100010",
  5102=>"110101001",
  5103=>"100001010",
  5104=>"111101110",
  5105=>"111000001",
  5106=>"001110011",
  5107=>"110110111",
  5108=>"000010010",
  5109=>"000001100",
  5110=>"001110110",
  5111=>"101001101",
  5112=>"100011110",
  5113=>"000000100",
  5114=>"011001011",
  5115=>"111111110",
  5116=>"001100111",
  5117=>"011011000",
  5118=>"000101011",
  5119=>"000011000",
  5120=>"110111000",
  5121=>"000010011",
  5122=>"000001110",
  5123=>"111100011",
  5124=>"111010000",
  5125=>"111111101",
  5126=>"011100001",
  5127=>"101100011",
  5128=>"000000010",
  5129=>"000000111",
  5130=>"100100011",
  5131=>"000011011",
  5132=>"101100000",
  5133=>"100001001",
  5134=>"111101101",
  5135=>"010010101",
  5136=>"100010000",
  5137=>"011101111",
  5138=>"010101001",
  5139=>"101000100",
  5140=>"011110111",
  5141=>"000011000",
  5142=>"011101111",
  5143=>"101100010",
  5144=>"001001100",
  5145=>"111110011",
  5146=>"100011010",
  5147=>"111010001",
  5148=>"001101001",
  5149=>"110000110",
  5150=>"101100110",
  5151=>"111010001",
  5152=>"111000011",
  5153=>"111010101",
  5154=>"100111101",
  5155=>"000111011",
  5156=>"101011010",
  5157=>"011101111",
  5158=>"110011100",
  5159=>"010000111",
  5160=>"101100000",
  5161=>"110001101",
  5162=>"110001000",
  5163=>"000010110",
  5164=>"001001010",
  5165=>"011100100",
  5166=>"111100011",
  5167=>"001001011",
  5168=>"100101000",
  5169=>"101000001",
  5170=>"001000111",
  5171=>"100110101",
  5172=>"010100001",
  5173=>"101001100",
  5174=>"110000011",
  5175=>"110101101",
  5176=>"011011110",
  5177=>"101100011",
  5178=>"000000000",
  5179=>"011001000",
  5180=>"101010110",
  5181=>"101000101",
  5182=>"110011000",
  5183=>"111000000",
  5184=>"000010111",
  5185=>"110111011",
  5186=>"001010000",
  5187=>"001000001",
  5188=>"111010010",
  5189=>"111010001",
  5190=>"001010101",
  5191=>"111100110",
  5192=>"000001000",
  5193=>"011000001",
  5194=>"100001110",
  5195=>"000110000",
  5196=>"111111101",
  5197=>"101111111",
  5198=>"111000110",
  5199=>"100011011",
  5200=>"111001000",
  5201=>"110010010",
  5202=>"101100010",
  5203=>"010111100",
  5204=>"000110101",
  5205=>"111100101",
  5206=>"000000101",
  5207=>"101110010",
  5208=>"001100110",
  5209=>"110001110",
  5210=>"101101111",
  5211=>"011100000",
  5212=>"010010100",
  5213=>"111111011",
  5214=>"001011111",
  5215=>"110000011",
  5216=>"111101110",
  5217=>"000100001",
  5218=>"101011000",
  5219=>"011010000",
  5220=>"001101100",
  5221=>"010100010",
  5222=>"111100111",
  5223=>"010011010",
  5224=>"000001100",
  5225=>"100111000",
  5226=>"001110010",
  5227=>"111100010",
  5228=>"000000000",
  5229=>"010101001",
  5230=>"100000001",
  5231=>"010010100",
  5232=>"000001101",
  5233=>"111110011",
  5234=>"011000111",
  5235=>"111111001",
  5236=>"010011111",
  5237=>"110000111",
  5238=>"000110110",
  5239=>"010110101",
  5240=>"111101011",
  5241=>"001011011",
  5242=>"101110110",
  5243=>"000101100",
  5244=>"101100111",
  5245=>"010001010",
  5246=>"111110001",
  5247=>"101001000",
  5248=>"111100001",
  5249=>"110000001",
  5250=>"000001001",
  5251=>"001101011",
  5252=>"111011100",
  5253=>"100111001",
  5254=>"111110101",
  5255=>"010010000",
  5256=>"100101011",
  5257=>"101110010",
  5258=>"111011100",
  5259=>"001111111",
  5260=>"010100010",
  5261=>"100101011",
  5262=>"011110000",
  5263=>"101111011",
  5264=>"101001011",
  5265=>"010011001",
  5266=>"011000010",
  5267=>"100010111",
  5268=>"101001001",
  5269=>"000011111",
  5270=>"111000000",
  5271=>"100001101",
  5272=>"001000001",
  5273=>"100100111",
  5274=>"100011110",
  5275=>"000111110",
  5276=>"100111100",
  5277=>"100110100",
  5278=>"000000010",
  5279=>"010010001",
  5280=>"111001011",
  5281=>"101101111",
  5282=>"011110111",
  5283=>"111111011",
  5284=>"101001010",
  5285=>"110101110",
  5286=>"000101101",
  5287=>"000101011",
  5288=>"001111010",
  5289=>"000001000",
  5290=>"000100000",
  5291=>"010000000",
  5292=>"000011010",
  5293=>"001011100",
  5294=>"110010101",
  5295=>"111000010",
  5296=>"101000011",
  5297=>"000001101",
  5298=>"010111110",
  5299=>"011010011",
  5300=>"100011111",
  5301=>"110011111",
  5302=>"000000010",
  5303=>"001010011",
  5304=>"101100100",
  5305=>"101000011",
  5306=>"011000010",
  5307=>"011011001",
  5308=>"011100000",
  5309=>"110101010",
  5310=>"101110111",
  5311=>"000100100",
  5312=>"101001000",
  5313=>"011001001",
  5314=>"010000111",
  5315=>"001010001",
  5316=>"100101110",
  5317=>"100010000",
  5318=>"011000110",
  5319=>"010110110",
  5320=>"101110011",
  5321=>"001101100",
  5322=>"101001111",
  5323=>"011000000",
  5324=>"001110101",
  5325=>"110111110",
  5326=>"101100101",
  5327=>"000001000",
  5328=>"001110001",
  5329=>"001111010",
  5330=>"010011110",
  5331=>"001101000",
  5332=>"001010000",
  5333=>"001001111",
  5334=>"100111001",
  5335=>"100111110",
  5336=>"101101100",
  5337=>"101010100",
  5338=>"011000011",
  5339=>"101011011",
  5340=>"000010001",
  5341=>"010110000",
  5342=>"001000100",
  5343=>"110110101",
  5344=>"001110100",
  5345=>"100100111",
  5346=>"111011000",
  5347=>"000101000",
  5348=>"000111111",
  5349=>"110010111",
  5350=>"100000111",
  5351=>"100110100",
  5352=>"011001110",
  5353=>"100111100",
  5354=>"000010001",
  5355=>"001111110",
  5356=>"000100010",
  5357=>"110001100",
  5358=>"100011010",
  5359=>"101110100",
  5360=>"100101011",
  5361=>"100000110",
  5362=>"101010111",
  5363=>"000001000",
  5364=>"000100000",
  5365=>"100110101",
  5366=>"100101101",
  5367=>"000100111",
  5368=>"001111111",
  5369=>"101011111",
  5370=>"000011001",
  5371=>"000101001",
  5372=>"000000101",
  5373=>"101100111",
  5374=>"010000000",
  5375=>"010001101",
  5376=>"101000011",
  5377=>"110011010",
  5378=>"000111110",
  5379=>"000101111",
  5380=>"111000011",
  5381=>"011010000",
  5382=>"010010110",
  5383=>"101011000",
  5384=>"000000111",
  5385=>"010111100",
  5386=>"110001011",
  5387=>"101110010",
  5388=>"000010100",
  5389=>"000101100",
  5390=>"000011111",
  5391=>"110000100",
  5392=>"010011111",
  5393=>"110100000",
  5394=>"011101011",
  5395=>"000111101",
  5396=>"001000010",
  5397=>"000001001",
  5398=>"000111011",
  5399=>"100101001",
  5400=>"011011000",
  5401=>"010110110",
  5402=>"011011000",
  5403=>"100001101",
  5404=>"010011101",
  5405=>"101111110",
  5406=>"010110110",
  5407=>"110100101",
  5408=>"000100101",
  5409=>"010000001",
  5410=>"111000100",
  5411=>"111101111",
  5412=>"001110010",
  5413=>"001100011",
  5414=>"101100001",
  5415=>"001000111",
  5416=>"001100100",
  5417=>"011000100",
  5418=>"110111010",
  5419=>"011011010",
  5420=>"000110010",
  5421=>"111011101",
  5422=>"100101001",
  5423=>"101110001",
  5424=>"111110011",
  5425=>"001100010",
  5426=>"010000100",
  5427=>"011101010",
  5428=>"000100100",
  5429=>"110111101",
  5430=>"110001000",
  5431=>"000110101",
  5432=>"100000110",
  5433=>"110001010",
  5434=>"000000100",
  5435=>"110111001",
  5436=>"000011000",
  5437=>"001010101",
  5438=>"101101100",
  5439=>"000011101",
  5440=>"111110111",
  5441=>"101110001",
  5442=>"100111000",
  5443=>"111110100",
  5444=>"111110101",
  5445=>"010100111",
  5446=>"011111010",
  5447=>"100100100",
  5448=>"110110110",
  5449=>"010100111",
  5450=>"101011110",
  5451=>"000010111",
  5452=>"001100100",
  5453=>"100111001",
  5454=>"110000001",
  5455=>"000011100",
  5456=>"011111011",
  5457=>"110011110",
  5458=>"011001000",
  5459=>"001000000",
  5460=>"001010001",
  5461=>"000000110",
  5462=>"111001000",
  5463=>"010110000",
  5464=>"001110010",
  5465=>"010011100",
  5466=>"001110100",
  5467=>"110111110",
  5468=>"111011101",
  5469=>"111000011",
  5470=>"110101001",
  5471=>"111110100",
  5472=>"110100111",
  5473=>"100100010",
  5474=>"011011100",
  5475=>"101111011",
  5476=>"001101000",
  5477=>"001000010",
  5478=>"111011011",
  5479=>"111011100",
  5480=>"010001000",
  5481=>"100110110",
  5482=>"001100100",
  5483=>"011010000",
  5484=>"000000111",
  5485=>"100101011",
  5486=>"100001101",
  5487=>"010101011",
  5488=>"010001110",
  5489=>"000000000",
  5490=>"011111010",
  5491=>"111010110",
  5492=>"000101101",
  5493=>"010101101",
  5494=>"001011100",
  5495=>"001111001",
  5496=>"000000000",
  5497=>"000111000",
  5498=>"011001001",
  5499=>"000010001",
  5500=>"101000000",
  5501=>"101100111",
  5502=>"001101000",
  5503=>"111111010",
  5504=>"101101010",
  5505=>"010001001",
  5506=>"100110001",
  5507=>"001111111",
  5508=>"010110100",
  5509=>"110100010",
  5510=>"000001110",
  5511=>"101110100",
  5512=>"000000010",
  5513=>"110001000",
  5514=>"100100110",
  5515=>"000001001",
  5516=>"100000100",
  5517=>"011001001",
  5518=>"101001000",
  5519=>"000110110",
  5520=>"001000011",
  5521=>"000000001",
  5522=>"001100100",
  5523=>"001100011",
  5524=>"011011011",
  5525=>"101110011",
  5526=>"111111101",
  5527=>"101010010",
  5528=>"111110000",
  5529=>"001000110",
  5530=>"110100111",
  5531=>"111111100",
  5532=>"100111111",
  5533=>"011000010",
  5534=>"110011000",
  5535=>"110011011",
  5536=>"000100110",
  5537=>"110000011",
  5538=>"001101100",
  5539=>"010011010",
  5540=>"001100101",
  5541=>"001101110",
  5542=>"000001000",
  5543=>"010001101",
  5544=>"001000100",
  5545=>"110101100",
  5546=>"110100111",
  5547=>"101011010",
  5548=>"010100111",
  5549=>"111111001",
  5550=>"000011110",
  5551=>"000001100",
  5552=>"000000011",
  5553=>"101011111",
  5554=>"010101110",
  5555=>"110110001",
  5556=>"001111101",
  5557=>"101000100",
  5558=>"011011111",
  5559=>"011011110",
  5560=>"100001000",
  5561=>"010000001",
  5562=>"000010011",
  5563=>"001001111",
  5564=>"110110000",
  5565=>"101110011",
  5566=>"000011100",
  5567=>"111001101",
  5568=>"111000111",
  5569=>"011100001",
  5570=>"010011000",
  5571=>"001000101",
  5572=>"000000110",
  5573=>"001111110",
  5574=>"111001101",
  5575=>"000100000",
  5576=>"100001111",
  5577=>"110110011",
  5578=>"011111110",
  5579=>"010110110",
  5580=>"010000101",
  5581=>"011111000",
  5582=>"110110101",
  5583=>"001100111",
  5584=>"011010000",
  5585=>"101000001",
  5586=>"000100011",
  5587=>"010001100",
  5588=>"101110001",
  5589=>"101101100",
  5590=>"111001111",
  5591=>"010110100",
  5592=>"110001010",
  5593=>"101101111",
  5594=>"110100110",
  5595=>"011000010",
  5596=>"000001001",
  5597=>"110010000",
  5598=>"100011100",
  5599=>"010110101",
  5600=>"001010010",
  5601=>"001111101",
  5602=>"100101011",
  5603=>"001111010",
  5604=>"100010100",
  5605=>"100010010",
  5606=>"011100100",
  5607=>"010110110",
  5608=>"011001011",
  5609=>"101101101",
  5610=>"010000001",
  5611=>"101101001",
  5612=>"000001110",
  5613=>"010010000",
  5614=>"001001010",
  5615=>"100101001",
  5616=>"001000110",
  5617=>"010001101",
  5618=>"101101010",
  5619=>"101101010",
  5620=>"111101000",
  5621=>"000001111",
  5622=>"101110110",
  5623=>"110001101",
  5624=>"010110010",
  5625=>"100110010",
  5626=>"111101001",
  5627=>"000011010",
  5628=>"011111001",
  5629=>"101110111",
  5630=>"010010010",
  5631=>"000001101",
  5632=>"100110001",
  5633=>"000000010",
  5634=>"101001110",
  5635=>"000000011",
  5636=>"000001110",
  5637=>"001000010",
  5638=>"111011000",
  5639=>"001011100",
  5640=>"000000001",
  5641=>"000001011",
  5642=>"111010111",
  5643=>"010110010",
  5644=>"111001101",
  5645=>"000000000",
  5646=>"000011111",
  5647=>"000100010",
  5648=>"001011100",
  5649=>"100101010",
  5650=>"101011011",
  5651=>"001101001",
  5652=>"010010010",
  5653=>"110010010",
  5654=>"100111001",
  5655=>"000100011",
  5656=>"111101010",
  5657=>"010110011",
  5658=>"001001000",
  5659=>"001011111",
  5660=>"011101000",
  5661=>"000000110",
  5662=>"110001110",
  5663=>"100111011",
  5664=>"010100101",
  5665=>"100000100",
  5666=>"000111110",
  5667=>"111001001",
  5668=>"100011101",
  5669=>"011111110",
  5670=>"000110001",
  5671=>"001101011",
  5672=>"001101001",
  5673=>"010111100",
  5674=>"010110110",
  5675=>"110000001",
  5676=>"011101011",
  5677=>"110001110",
  5678=>"111100100",
  5679=>"010010010",
  5680=>"100000000",
  5681=>"010111001",
  5682=>"000001001",
  5683=>"111001111",
  5684=>"000101000",
  5685=>"001101100",
  5686=>"110111010",
  5687=>"001011000",
  5688=>"000101001",
  5689=>"101111110",
  5690=>"010001100",
  5691=>"111010000",
  5692=>"011011101",
  5693=>"111010000",
  5694=>"101010010",
  5695=>"001100100",
  5696=>"111100011",
  5697=>"100110001",
  5698=>"101000000",
  5699=>"111111110",
  5700=>"000100010",
  5701=>"000000100",
  5702=>"010100010",
  5703=>"011010010",
  5704=>"011100101",
  5705=>"001011100",
  5706=>"101001111",
  5707=>"100110101",
  5708=>"101001100",
  5709=>"101000100",
  5710=>"110000110",
  5711=>"000000010",
  5712=>"011111011",
  5713=>"011100010",
  5714=>"101110100",
  5715=>"011011000",
  5716=>"011100111",
  5717=>"010101111",
  5718=>"000110100",
  5719=>"011010000",
  5720=>"100000101",
  5721=>"111101100",
  5722=>"100011101",
  5723=>"100010101",
  5724=>"110011010",
  5725=>"010101111",
  5726=>"101001001",
  5727=>"111111101",
  5728=>"100001011",
  5729=>"000100010",
  5730=>"011000110",
  5731=>"110110000",
  5732=>"110000111",
  5733=>"110000100",
  5734=>"000011011",
  5735=>"010101011",
  5736=>"001001001",
  5737=>"010110001",
  5738=>"100111100",
  5739=>"111100001",
  5740=>"111101101",
  5741=>"001100011",
  5742=>"001010000",
  5743=>"101000010",
  5744=>"111111010",
  5745=>"011001101",
  5746=>"011100100",
  5747=>"100000111",
  5748=>"100110010",
  5749=>"011000000",
  5750=>"011110010",
  5751=>"010011100",
  5752=>"010110111",
  5753=>"111000011",
  5754=>"001000111",
  5755=>"000111100",
  5756=>"110111000",
  5757=>"100000011",
  5758=>"100100000",
  5759=>"011011100",
  5760=>"110100111",
  5761=>"011111111",
  5762=>"010110000",
  5763=>"000010110",
  5764=>"101110000",
  5765=>"110001111",
  5766=>"010010101",
  5767=>"110011100",
  5768=>"000000101",
  5769=>"000010011",
  5770=>"111101010",
  5771=>"110011001",
  5772=>"010101110",
  5773=>"011000010",
  5774=>"110111001",
  5775=>"111111111",
  5776=>"011100101",
  5777=>"000010010",
  5778=>"100110111",
  5779=>"111100111",
  5780=>"001100001",
  5781=>"011110101",
  5782=>"111101001",
  5783=>"100000000",
  5784=>"011010111",
  5785=>"001000101",
  5786=>"000001000",
  5787=>"101010110",
  5788=>"101000010",
  5789=>"100111101",
  5790=>"010101100",
  5791=>"001110011",
  5792=>"100111011",
  5793=>"101111011",
  5794=>"110011100",
  5795=>"001110000",
  5796=>"001100101",
  5797=>"111110101",
  5798=>"111011010",
  5799=>"011111010",
  5800=>"011000111",
  5801=>"110010100",
  5802=>"101011000",
  5803=>"100000110",
  5804=>"001101110",
  5805=>"011001011",
  5806=>"000111000",
  5807=>"100101001",
  5808=>"000011110",
  5809=>"010000110",
  5810=>"110000001",
  5811=>"100100101",
  5812=>"111001011",
  5813=>"001001100",
  5814=>"110100101",
  5815=>"001010001",
  5816=>"000111111",
  5817=>"100101100",
  5818=>"001101011",
  5819=>"101100111",
  5820=>"011010001",
  5821=>"110010100",
  5822=>"100000100",
  5823=>"000111011",
  5824=>"001101001",
  5825=>"000011011",
  5826=>"010110000",
  5827=>"100000000",
  5828=>"011010001",
  5829=>"101111011",
  5830=>"110010100",
  5831=>"011111010",
  5832=>"000000100",
  5833=>"110110001",
  5834=>"011100100",
  5835=>"010010010",
  5836=>"011101011",
  5837=>"011001111",
  5838=>"010000011",
  5839=>"001011011",
  5840=>"001101100",
  5841=>"001011110",
  5842=>"111110000",
  5843=>"010000011",
  5844=>"110110100",
  5845=>"010110100",
  5846=>"111000010",
  5847=>"110011011",
  5848=>"101111100",
  5849=>"011011100",
  5850=>"101010000",
  5851=>"001110100",
  5852=>"101101111",
  5853=>"111111100",
  5854=>"010011010",
  5855=>"001011011",
  5856=>"110110010",
  5857=>"100001010",
  5858=>"111001111",
  5859=>"010010101",
  5860=>"111101000",
  5861=>"110110110",
  5862=>"000100000",
  5863=>"001001000",
  5864=>"101001111",
  5865=>"111110110",
  5866=>"011000111",
  5867=>"011110000",
  5868=>"000000101",
  5869=>"110100111",
  5870=>"001111101",
  5871=>"110000101",
  5872=>"110010110",
  5873=>"000100100",
  5874=>"010010011",
  5875=>"110011100",
  5876=>"111010010",
  5877=>"110100001",
  5878=>"011000010",
  5879=>"011100100",
  5880=>"111001001",
  5881=>"001011011",
  5882=>"101101001",
  5883=>"110111100",
  5884=>"100001010",
  5885=>"010000100",
  5886=>"110100111",
  5887=>"100000111",
  5888=>"010010000",
  5889=>"011100011",
  5890=>"010001000",
  5891=>"000011010",
  5892=>"001110111",
  5893=>"011100010",
  5894=>"010101111",
  5895=>"011101101",
  5896=>"100100011",
  5897=>"000000111",
  5898=>"110011110",
  5899=>"101101111",
  5900=>"001101010",
  5901=>"011000010",
  5902=>"011100010",
  5903=>"110000110",
  5904=>"100111111",
  5905=>"100101100",
  5906=>"100110000",
  5907=>"011110001",
  5908=>"011011010",
  5909=>"000011110",
  5910=>"110100011",
  5911=>"101111011",
  5912=>"100010010",
  5913=>"001001011",
  5914=>"101001011",
  5915=>"010111110",
  5916=>"010011001",
  5917=>"111100010",
  5918=>"010110101",
  5919=>"001100100",
  5920=>"110101000",
  5921=>"111010010",
  5922=>"001001110",
  5923=>"010001000",
  5924=>"010000000",
  5925=>"010000000",
  5926=>"001000110",
  5927=>"111001110",
  5928=>"101100011",
  5929=>"001000000",
  5930=>"111101100",
  5931=>"100010001",
  5932=>"111001011",
  5933=>"000110011",
  5934=>"001011011",
  5935=>"110100110",
  5936=>"010000111",
  5937=>"000001110",
  5938=>"100011110",
  5939=>"001111100",
  5940=>"111100101",
  5941=>"100000010",
  5942=>"111010000",
  5943=>"100101110",
  5944=>"010111110",
  5945=>"111011111",
  5946=>"010011011",
  5947=>"001101000",
  5948=>"111111110",
  5949=>"001001101",
  5950=>"011000011",
  5951=>"011111110",
  5952=>"000000010",
  5953=>"011101111",
  5954=>"011001111",
  5955=>"110111000",
  5956=>"011000010",
  5957=>"000011010",
  5958=>"011100100",
  5959=>"100110100",
  5960=>"000011100",
  5961=>"101101001",
  5962=>"001010011",
  5963=>"111111100",
  5964=>"000101110",
  5965=>"010110110",
  5966=>"101010111",
  5967=>"111101011",
  5968=>"011010011",
  5969=>"000101111",
  5970=>"101100100",
  5971=>"000001111",
  5972=>"100111000",
  5973=>"011111010",
  5974=>"110111111",
  5975=>"000001110",
  5976=>"000100000",
  5977=>"011000010",
  5978=>"111100001",
  5979=>"110001110",
  5980=>"101000100",
  5981=>"001000110",
  5982=>"001101101",
  5983=>"101110010",
  5984=>"110111110",
  5985=>"110010111",
  5986=>"011000001",
  5987=>"011000101",
  5988=>"101111100",
  5989=>"010100101",
  5990=>"101111010",
  5991=>"111001000",
  5992=>"101000000",
  5993=>"010110110",
  5994=>"100110000",
  5995=>"110010101",
  5996=>"010110111",
  5997=>"001101011",
  5998=>"000111110",
  5999=>"001010011",
  6000=>"000000100",
  6001=>"000100011",
  6002=>"111000000",
  6003=>"011000100",
  6004=>"110000001",
  6005=>"001010000",
  6006=>"010001011",
  6007=>"011111010",
  6008=>"101101111",
  6009=>"011100101",
  6010=>"110000011",
  6011=>"001011110",
  6012=>"000100100",
  6013=>"000001001",
  6014=>"011010100",
  6015=>"111100101",
  6016=>"011111111",
  6017=>"011110111",
  6018=>"001001111",
  6019=>"001001100",
  6020=>"110001100",
  6021=>"110110000",
  6022=>"100001000",
  6023=>"001110111",
  6024=>"010101111",
  6025=>"001101011",
  6026=>"000111000",
  6027=>"100101100",
  6028=>"100001001",
  6029=>"100101111",
  6030=>"110110101",
  6031=>"101011100",
  6032=>"010100011",
  6033=>"111100011",
  6034=>"000100111",
  6035=>"111110110",
  6036=>"010011010",
  6037=>"111110010",
  6038=>"101000110",
  6039=>"011000100",
  6040=>"111101010",
  6041=>"110100111",
  6042=>"010010111",
  6043=>"001110111",
  6044=>"101001000",
  6045=>"111000100",
  6046=>"000100110",
  6047=>"011100000",
  6048=>"000000010",
  6049=>"111010010",
  6050=>"110011010",
  6051=>"001011010",
  6052=>"011010000",
  6053=>"110111011",
  6054=>"011010110",
  6055=>"011101100",
  6056=>"010000100",
  6057=>"000001010",
  6058=>"001101101",
  6059=>"111110111",
  6060=>"110111001",
  6061=>"111100101",
  6062=>"111000110",
  6063=>"111111101",
  6064=>"000001110",
  6065=>"110000011",
  6066=>"100010111",
  6067=>"100000001",
  6068=>"101110000",
  6069=>"001011011",
  6070=>"010000001",
  6071=>"110010110",
  6072=>"110001101",
  6073=>"001110001",
  6074=>"000011100",
  6075=>"101100000",
  6076=>"101101001",
  6077=>"111010100",
  6078=>"010001000",
  6079=>"100100111",
  6080=>"000010101",
  6081=>"011010101",
  6082=>"001010111",
  6083=>"100101100",
  6084=>"111111101",
  6085=>"100111011",
  6086=>"000101010",
  6087=>"101010010",
  6088=>"110110100",
  6089=>"001100110",
  6090=>"100110001",
  6091=>"111101111",
  6092=>"011111110",
  6093=>"100000010",
  6094=>"100011000",
  6095=>"001111011",
  6096=>"100011101",
  6097=>"101011100",
  6098=>"001001011",
  6099=>"100100111",
  6100=>"000000000",
  6101=>"011001010",
  6102=>"010111101",
  6103=>"000000100",
  6104=>"011001111",
  6105=>"110110010",
  6106=>"100010001",
  6107=>"110000000",
  6108=>"101110010",
  6109=>"011000111",
  6110=>"001001010",
  6111=>"100100110",
  6112=>"100110011",
  6113=>"111001000",
  6114=>"110100000",
  6115=>"110010001",
  6116=>"000110000",
  6117=>"001101111",
  6118=>"101001000",
  6119=>"011010011",
  6120=>"100010010",
  6121=>"000001101",
  6122=>"000011001",
  6123=>"011001011",
  6124=>"010110100",
  6125=>"110111101",
  6126=>"001111101",
  6127=>"111010001",
  6128=>"001111000",
  6129=>"010101110",
  6130=>"001000101",
  6131=>"010101000",
  6132=>"001001111",
  6133=>"001110010",
  6134=>"011010101",
  6135=>"100011010",
  6136=>"101111001",
  6137=>"100011110",
  6138=>"111100100",
  6139=>"010010100",
  6140=>"110011110",
  6141=>"011010100",
  6142=>"011010000",
  6143=>"100100000",
  6144=>"000110011",
  6145=>"011100100",
  6146=>"111111000",
  6147=>"111101011",
  6148=>"011101001",
  6149=>"100000101",
  6150=>"110010000",
  6151=>"010010010",
  6152=>"100100011",
  6153=>"011100011",
  6154=>"100010001",
  6155=>"011010001",
  6156=>"101100001",
  6157=>"000111010",
  6158=>"001000000",
  6159=>"111110101",
  6160=>"001100001",
  6161=>"111011110",
  6162=>"111000010",
  6163=>"111011111",
  6164=>"010111010",
  6165=>"111100011",
  6166=>"000111000",
  6167=>"001001010",
  6168=>"000111010",
  6169=>"110000100",
  6170=>"010110110",
  6171=>"000101110",
  6172=>"101100111",
  6173=>"001001000",
  6174=>"110101101",
  6175=>"001111010",
  6176=>"010100111",
  6177=>"100100011",
  6178=>"101111101",
  6179=>"111011011",
  6180=>"111100101",
  6181=>"011111101",
  6182=>"111111010",
  6183=>"000111110",
  6184=>"100001100",
  6185=>"010100101",
  6186=>"111101011",
  6187=>"100100011",
  6188=>"101011101",
  6189=>"000010100",
  6190=>"111011001",
  6191=>"101000110",
  6192=>"000101001",
  6193=>"000111110",
  6194=>"001010000",
  6195=>"111100001",
  6196=>"101111110",
  6197=>"100110010",
  6198=>"011101111",
  6199=>"101010010",
  6200=>"101010001",
  6201=>"010000001",
  6202=>"111011011",
  6203=>"100100110",
  6204=>"000110000",
  6205=>"110000100",
  6206=>"010101111",
  6207=>"111111011",
  6208=>"100110011",
  6209=>"010010110",
  6210=>"010011101",
  6211=>"100001110",
  6212=>"110001101",
  6213=>"100111111",
  6214=>"100011101",
  6215=>"111111001",
  6216=>"110000101",
  6217=>"011010110",
  6218=>"110001001",
  6219=>"101100101",
  6220=>"111010011",
  6221=>"011000110",
  6222=>"011100100",
  6223=>"101110111",
  6224=>"111101011",
  6225=>"101001100",
  6226=>"110111000",
  6227=>"010001100",
  6228=>"000000001",
  6229=>"111101011",
  6230=>"100010011",
  6231=>"010010010",
  6232=>"111100110",
  6233=>"110010010",
  6234=>"100000000",
  6235=>"111011001",
  6236=>"011000000",
  6237=>"110000000",
  6238=>"010011100",
  6239=>"101001111",
  6240=>"101001011",
  6241=>"001110110",
  6242=>"110110100",
  6243=>"111110001",
  6244=>"000110101",
  6245=>"011010110",
  6246=>"010110110",
  6247=>"000111110",
  6248=>"011000101",
  6249=>"111001101",
  6250=>"010010000",
  6251=>"100010110",
  6252=>"101000111",
  6253=>"001100000",
  6254=>"110001010",
  6255=>"001101110",
  6256=>"101110001",
  6257=>"010111110",
  6258=>"111101000",
  6259=>"011001110",
  6260=>"011100001",
  6261=>"100110001",
  6262=>"011100011",
  6263=>"001001100",
  6264=>"100111111",
  6265=>"001101101",
  6266=>"100000111",
  6267=>"000100000",
  6268=>"101000011",
  6269=>"111110111",
  6270=>"010000010",
  6271=>"111111111",
  6272=>"111111000",
  6273=>"101010011",
  6274=>"110001100",
  6275=>"100111110",
  6276=>"011100101",
  6277=>"011101001",
  6278=>"100110101",
  6279=>"110010001",
  6280=>"001101001",
  6281=>"011101100",
  6282=>"101100000",
  6283=>"000001000",
  6284=>"101000001",
  6285=>"111001100",
  6286=>"111100000",
  6287=>"111010101",
  6288=>"010001100",
  6289=>"100100010",
  6290=>"010101100",
  6291=>"101101011",
  6292=>"000101111",
  6293=>"101100000",
  6294=>"111111010",
  6295=>"111010100",
  6296=>"111001101",
  6297=>"000001000",
  6298=>"110000011",
  6299=>"101011101",
  6300=>"010010000",
  6301=>"011100011",
  6302=>"010001011",
  6303=>"111001111",
  6304=>"100000001",
  6305=>"101000001",
  6306=>"011100101",
  6307=>"000010001",
  6308=>"101010000",
  6309=>"010011010",
  6310=>"111001101",
  6311=>"011100110",
  6312=>"101110100",
  6313=>"100101110",
  6314=>"101010001",
  6315=>"001001010",
  6316=>"100001001",
  6317=>"010101001",
  6318=>"110111111",
  6319=>"001001100",
  6320=>"000111101",
  6321=>"001000000",
  6322=>"100001101",
  6323=>"000000001",
  6324=>"000110111",
  6325=>"010010110",
  6326=>"100010000",
  6327=>"110111110",
  6328=>"001110000",
  6329=>"111001010",
  6330=>"101100110",
  6331=>"010011111",
  6332=>"011010011",
  6333=>"100001001",
  6334=>"110000001",
  6335=>"000000110",
  6336=>"000100001",
  6337=>"110100000",
  6338=>"010111010",
  6339=>"011111010",
  6340=>"000001011",
  6341=>"110001111",
  6342=>"000100101",
  6343=>"001001110",
  6344=>"111101101",
  6345=>"011101000",
  6346=>"011000011",
  6347=>"111000101",
  6348=>"111101000",
  6349=>"010101111",
  6350=>"101101100",
  6351=>"100000010",
  6352=>"101101011",
  6353=>"101010100",
  6354=>"110011101",
  6355=>"100101011",
  6356=>"011110001",
  6357=>"100101101",
  6358=>"011011101",
  6359=>"001001011",
  6360=>"001001011",
  6361=>"000111001",
  6362=>"000010111",
  6363=>"101001101",
  6364=>"101110110",
  6365=>"101101100",
  6366=>"010100101",
  6367=>"101111000",
  6368=>"110000111",
  6369=>"110100000",
  6370=>"011110001",
  6371=>"000001000",
  6372=>"101110111",
  6373=>"011111100",
  6374=>"111101110",
  6375=>"001100010",
  6376=>"101110110",
  6377=>"100000110",
  6378=>"110101111",
  6379=>"000000011",
  6380=>"000000101",
  6381=>"001111111",
  6382=>"001001111",
  6383=>"111000010",
  6384=>"011011111",
  6385=>"100011010",
  6386=>"001010001",
  6387=>"011100100",
  6388=>"100010111",
  6389=>"000000110",
  6390=>"011001101",
  6391=>"111101100",
  6392=>"001100101",
  6393=>"100110110",
  6394=>"010000011",
  6395=>"110000011",
  6396=>"010101001",
  6397=>"010100000",
  6398=>"000100010",
  6399=>"111101111",
  6400=>"101101001",
  6401=>"000111001",
  6402=>"000100011",
  6403=>"011110101",
  6404=>"100100111",
  6405=>"000001111",
  6406=>"100111000",
  6407=>"100010001",
  6408=>"111100101",
  6409=>"110010001",
  6410=>"011011101",
  6411=>"011011101",
  6412=>"001110110",
  6413=>"001011110",
  6414=>"110010010",
  6415=>"111101111",
  6416=>"110011010",
  6417=>"110110001",
  6418=>"101101101",
  6419=>"100001111",
  6420=>"110110111",
  6421=>"111001011",
  6422=>"111111111",
  6423=>"100010111",
  6424=>"100001010",
  6425=>"111010000",
  6426=>"011010011",
  6427=>"111101000",
  6428=>"010011010",
  6429=>"110110011",
  6430=>"001000000",
  6431=>"011111110",
  6432=>"000111000",
  6433=>"110100111",
  6434=>"110010000",
  6435=>"110010001",
  6436=>"010010001",
  6437=>"111110100",
  6438=>"101101100",
  6439=>"101100010",
  6440=>"100100010",
  6441=>"111001001",
  6442=>"011111010",
  6443=>"101111010",
  6444=>"011111010",
  6445=>"101101011",
  6446=>"110000111",
  6447=>"101111100",
  6448=>"110100001",
  6449=>"100001000",
  6450=>"100100111",
  6451=>"001000100",
  6452=>"001100111",
  6453=>"110100100",
  6454=>"110111001",
  6455=>"101000011",
  6456=>"010010001",
  6457=>"001101111",
  6458=>"111010011",
  6459=>"111001100",
  6460=>"000111100",
  6461=>"100010001",
  6462=>"000100000",
  6463=>"011011101",
  6464=>"110010000",
  6465=>"100001101",
  6466=>"110101011",
  6467=>"011101101",
  6468=>"011001000",
  6469=>"100000010",
  6470=>"111010000",
  6471=>"001101101",
  6472=>"110010000",
  6473=>"111111110",
  6474=>"101000101",
  6475=>"111010011",
  6476=>"101011110",
  6477=>"000100101",
  6478=>"101111111",
  6479=>"010010010",
  6480=>"011000111",
  6481=>"101001100",
  6482=>"001101010",
  6483=>"000000010",
  6484=>"100011110",
  6485=>"111111100",
  6486=>"101000100",
  6487=>"111000001",
  6488=>"011111010",
  6489=>"100000001",
  6490=>"000101001",
  6491=>"111001010",
  6492=>"101111001",
  6493=>"100111110",
  6494=>"000011010",
  6495=>"110000000",
  6496=>"110111110",
  6497=>"100010110",
  6498=>"010100011",
  6499=>"101110011",
  6500=>"100010011",
  6501=>"110110011",
  6502=>"111101011",
  6503=>"001000001",
  6504=>"111000111",
  6505=>"111111111",
  6506=>"000111110",
  6507=>"111111100",
  6508=>"000111000",
  6509=>"010100011",
  6510=>"001000000",
  6511=>"000000100",
  6512=>"001001011",
  6513=>"110110110",
  6514=>"101110001",
  6515=>"100100110",
  6516=>"000001111",
  6517=>"001000000",
  6518=>"101011100",
  6519=>"001001011",
  6520=>"001010000",
  6521=>"011101011",
  6522=>"010111111",
  6523=>"100111110",
  6524=>"101000000",
  6525=>"001010001",
  6526=>"101101011",
  6527=>"111001100",
  6528=>"000001001",
  6529=>"011000100",
  6530=>"100000100",
  6531=>"111100100",
  6532=>"101010011",
  6533=>"010010001",
  6534=>"100001111",
  6535=>"010111100",
  6536=>"100100111",
  6537=>"100010100",
  6538=>"000001011",
  6539=>"101110110",
  6540=>"111101101",
  6541=>"111011001",
  6542=>"001111011",
  6543=>"110010100",
  6544=>"001101101",
  6545=>"001001101",
  6546=>"110000111",
  6547=>"010000001",
  6548=>"110010101",
  6549=>"101111100",
  6550=>"110101100",
  6551=>"000100011",
  6552=>"001001011",
  6553=>"111011001",
  6554=>"010001010",
  6555=>"001110110",
  6556=>"111000101",
  6557=>"111011001",
  6558=>"001011100",
  6559=>"000011010",
  6560=>"111100111",
  6561=>"110111000",
  6562=>"010010100",
  6563=>"101101101",
  6564=>"001111101",
  6565=>"111110000",
  6566=>"101001010",
  6567=>"111011010",
  6568=>"111101000",
  6569=>"111011111",
  6570=>"001001101",
  6571=>"001010011",
  6572=>"101101001",
  6573=>"010010000",
  6574=>"001111001",
  6575=>"111100110",
  6576=>"010101011",
  6577=>"100100110",
  6578=>"000001111",
  6579=>"010010011",
  6580=>"001001000",
  6581=>"111110110",
  6582=>"110011111",
  6583=>"000100111",
  6584=>"110100101",
  6585=>"000010111",
  6586=>"101011010",
  6587=>"001001110",
  6588=>"111011100",
  6589=>"111010110",
  6590=>"100111110",
  6591=>"111101000",
  6592=>"111111000",
  6593=>"111110011",
  6594=>"001000001",
  6595=>"111011100",
  6596=>"010101110",
  6597=>"111111100",
  6598=>"100100001",
  6599=>"000110011",
  6600=>"011101001",
  6601=>"101010110",
  6602=>"110111010",
  6603=>"011001010",
  6604=>"000111101",
  6605=>"110111011",
  6606=>"000011000",
  6607=>"111011011",
  6608=>"110110111",
  6609=>"011000010",
  6610=>"111110100",
  6611=>"000111100",
  6612=>"101110001",
  6613=>"010000110",
  6614=>"000010001",
  6615=>"111111011",
  6616=>"111000111",
  6617=>"100111101",
  6618=>"011011011",
  6619=>"001111110",
  6620=>"011100000",
  6621=>"001100011",
  6622=>"011001110",
  6623=>"100010101",
  6624=>"011100001",
  6625=>"010011010",
  6626=>"110000111",
  6627=>"100010000",
  6628=>"010001011",
  6629=>"010001010",
  6630=>"100101000",
  6631=>"011111010",
  6632=>"101101100",
  6633=>"111110000",
  6634=>"101010101",
  6635=>"111010110",
  6636=>"010000011",
  6637=>"001110011",
  6638=>"010011011",
  6639=>"011001111",
  6640=>"111001011",
  6641=>"101101001",
  6642=>"100111111",
  6643=>"111111111",
  6644=>"110100101",
  6645=>"000111110",
  6646=>"100000100",
  6647=>"011100101",
  6648=>"011101011",
  6649=>"010111101",
  6650=>"111110110",
  6651=>"100011010",
  6652=>"010101101",
  6653=>"001110000",
  6654=>"000001010",
  6655=>"000011101",
  6656=>"011111000",
  6657=>"110011000",
  6658=>"110010011",
  6659=>"101000100",
  6660=>"000100010",
  6661=>"010001000",
  6662=>"110010011",
  6663=>"110001101",
  6664=>"000010000",
  6665=>"101000001",
  6666=>"111110101",
  6667=>"000011001",
  6668=>"000100110",
  6669=>"011000100",
  6670=>"111000001",
  6671=>"101110111",
  6672=>"101011110",
  6673=>"011000011",
  6674=>"111110111",
  6675=>"100000011",
  6676=>"001101000",
  6677=>"111000110",
  6678=>"111110010",
  6679=>"010111100",
  6680=>"000001000",
  6681=>"100101111",
  6682=>"101101100",
  6683=>"010001110",
  6684=>"111001101",
  6685=>"011011110",
  6686=>"110000111",
  6687=>"000001011",
  6688=>"101101001",
  6689=>"011011011",
  6690=>"101010001",
  6691=>"010000010",
  6692=>"100001111",
  6693=>"110110000",
  6694=>"001000110",
  6695=>"000001001",
  6696=>"100100001",
  6697=>"011110100",
  6698=>"100000110",
  6699=>"001100000",
  6700=>"011110111",
  6701=>"100110001",
  6702=>"010110011",
  6703=>"100101101",
  6704=>"110111111",
  6705=>"111010000",
  6706=>"110011101",
  6707=>"011000000",
  6708=>"010110000",
  6709=>"111001010",
  6710=>"110100001",
  6711=>"011111101",
  6712=>"111100111",
  6713=>"011011001",
  6714=>"110011011",
  6715=>"110011100",
  6716=>"100100100",
  6717=>"010000010",
  6718=>"011100111",
  6719=>"100100011",
  6720=>"101110001",
  6721=>"100111111",
  6722=>"000100001",
  6723=>"010100010",
  6724=>"000111110",
  6725=>"101000101",
  6726=>"111100110",
  6727=>"010110100",
  6728=>"001100111",
  6729=>"001001010",
  6730=>"011101110",
  6731=>"001001000",
  6732=>"111001111",
  6733=>"110100110",
  6734=>"000110010",
  6735=>"001011000",
  6736=>"010010100",
  6737=>"000111100",
  6738=>"000110010",
  6739=>"010000101",
  6740=>"010010100",
  6741=>"110001010",
  6742=>"100100100",
  6743=>"010011001",
  6744=>"000010110",
  6745=>"000110111",
  6746=>"100100100",
  6747=>"111111100",
  6748=>"010000011",
  6749=>"110110000",
  6750=>"001111000",
  6751=>"101001001",
  6752=>"111001111",
  6753=>"010100100",
  6754=>"011101011",
  6755=>"100001001",
  6756=>"011011010",
  6757=>"100001110",
  6758=>"011011000",
  6759=>"001011010",
  6760=>"101100100",
  6761=>"010110111",
  6762=>"000000110",
  6763=>"110100101",
  6764=>"111011000",
  6765=>"011101110",
  6766=>"011111010",
  6767=>"110100101",
  6768=>"001001100",
  6769=>"100011111",
  6770=>"101111100",
  6771=>"100101010",
  6772=>"011100111",
  6773=>"100100010",
  6774=>"010000111",
  6775=>"000001010",
  6776=>"111100100",
  6777=>"011110101",
  6778=>"011100000",
  6779=>"010101001",
  6780=>"111010100",
  6781=>"000010000",
  6782=>"011001111",
  6783=>"101000100",
  6784=>"001000110",
  6785=>"111110001",
  6786=>"101101101",
  6787=>"111110000",
  6788=>"100111101",
  6789=>"010111011",
  6790=>"011110101",
  6791=>"101011101",
  6792=>"101001111",
  6793=>"010001011",
  6794=>"010111101",
  6795=>"011101110",
  6796=>"111001101",
  6797=>"111011100",
  6798=>"111101101",
  6799=>"111110010",
  6800=>"000011110",
  6801=>"011101001",
  6802=>"111111000",
  6803=>"100101001",
  6804=>"000001000",
  6805=>"110100011",
  6806=>"100010001",
  6807=>"010110101",
  6808=>"111110001",
  6809=>"111001101",
  6810=>"011111010",
  6811=>"111011111",
  6812=>"011110100",
  6813=>"001101001",
  6814=>"001110111",
  6815=>"110111011",
  6816=>"000000110",
  6817=>"100100000",
  6818=>"101100111",
  6819=>"100111111",
  6820=>"111000101",
  6821=>"001000110",
  6822=>"010100010",
  6823=>"100011010",
  6824=>"011110100",
  6825=>"000101100",
  6826=>"000001100",
  6827=>"111110010",
  6828=>"111111000",
  6829=>"100111011",
  6830=>"011101010",
  6831=>"100111011",
  6832=>"111011010",
  6833=>"110011101",
  6834=>"111101001",
  6835=>"100001100",
  6836=>"011001000",
  6837=>"001111010",
  6838=>"010101000",
  6839=>"001100110",
  6840=>"011110011",
  6841=>"100011110",
  6842=>"111011111",
  6843=>"011111001",
  6844=>"011011111",
  6845=>"010110001",
  6846=>"110010010",
  6847=>"011000101",
  6848=>"111001100",
  6849=>"110100100",
  6850=>"111001100",
  6851=>"101101001",
  6852=>"100011000",
  6853=>"001001100",
  6854=>"011011100",
  6855=>"001001001",
  6856=>"010111111",
  6857=>"111101011",
  6858=>"001010111",
  6859=>"101001101",
  6860=>"000110100",
  6861=>"111011001",
  6862=>"101010011",
  6863=>"000010000",
  6864=>"111100010",
  6865=>"010000110",
  6866=>"111010111",
  6867=>"000110010",
  6868=>"000000010",
  6869=>"111001001",
  6870=>"110001111",
  6871=>"010101100",
  6872=>"011111100",
  6873=>"000110101",
  6874=>"000100010",
  6875=>"001010000",
  6876=>"000011101",
  6877=>"011100010",
  6878=>"110101110",
  6879=>"001101110",
  6880=>"100000000",
  6881=>"100010000",
  6882=>"000101001",
  6883=>"001011100",
  6884=>"000001110",
  6885=>"001011100",
  6886=>"000000110",
  6887=>"101000001",
  6888=>"010011110",
  6889=>"101111110",
  6890=>"110101101",
  6891=>"110100100",
  6892=>"001001110",
  6893=>"111000000",
  6894=>"011011101",
  6895=>"110101011",
  6896=>"111001100",
  6897=>"000001010",
  6898=>"000010010",
  6899=>"100111100",
  6900=>"110110100",
  6901=>"111000110",
  6902=>"111011111",
  6903=>"011101101",
  6904=>"000010110",
  6905=>"111111110",
  6906=>"101010001",
  6907=>"101101101",
  6908=>"101001100",
  6909=>"010100110",
  6910=>"010110000",
  6911=>"111111111",
  6912=>"111001000",
  6913=>"111110000",
  6914=>"001000110",
  6915=>"111011011",
  6916=>"001001011",
  6917=>"111000111",
  6918=>"000000001",
  6919=>"111111111",
  6920=>"011011011",
  6921=>"010111011",
  6922=>"010110000",
  6923=>"010010101",
  6924=>"101011110",
  6925=>"011011010",
  6926=>"001000100",
  6927=>"001111100",
  6928=>"010011011",
  6929=>"001101110",
  6930=>"011011101",
  6931=>"001100110",
  6932=>"111001110",
  6933=>"001100011",
  6934=>"001111100",
  6935=>"001001111",
  6936=>"111111100",
  6937=>"101101000",
  6938=>"111001100",
  6939=>"010100000",
  6940=>"000001100",
  6941=>"100000000",
  6942=>"101010001",
  6943=>"111100001",
  6944=>"001000001",
  6945=>"010111011",
  6946=>"010000000",
  6947=>"111010010",
  6948=>"111111100",
  6949=>"000010101",
  6950=>"011001010",
  6951=>"000011000",
  6952=>"001001011",
  6953=>"000011001",
  6954=>"100100010",
  6955=>"100000110",
  6956=>"100100100",
  6957=>"100001000",
  6958=>"100111000",
  6959=>"111101110",
  6960=>"111110001",
  6961=>"011000100",
  6962=>"000000010",
  6963=>"110010011",
  6964=>"110011011",
  6965=>"011000011",
  6966=>"011011011",
  6967=>"000000011",
  6968=>"101111111",
  6969=>"101000101",
  6970=>"110110000",
  6971=>"101110111",
  6972=>"011010111",
  6973=>"000001101",
  6974=>"101011111",
  6975=>"000010111",
  6976=>"001100100",
  6977=>"000001111",
  6978=>"111111010",
  6979=>"110010011",
  6980=>"100111011",
  6981=>"010010001",
  6982=>"001101101",
  6983=>"010101111",
  6984=>"011110011",
  6985=>"110001011",
  6986=>"110110100",
  6987=>"110111010",
  6988=>"100010100",
  6989=>"000000010",
  6990=>"110001101",
  6991=>"100001000",
  6992=>"000110111",
  6993=>"101111100",
  6994=>"000111011",
  6995=>"100011111",
  6996=>"001011101",
  6997=>"100110100",
  6998=>"011010011",
  6999=>"110110010",
  7000=>"000011010",
  7001=>"101110111",
  7002=>"111000011",
  7003=>"111110010",
  7004=>"001000101",
  7005=>"111110011",
  7006=>"111111011",
  7007=>"000101001",
  7008=>"011101010",
  7009=>"001110000",
  7010=>"100011000",
  7011=>"001110110",
  7012=>"001101101",
  7013=>"101101111",
  7014=>"101110010",
  7015=>"100110101",
  7016=>"110000101",
  7017=>"111000000",
  7018=>"010111100",
  7019=>"100010110",
  7020=>"110010111",
  7021=>"111111111",
  7022=>"010000101",
  7023=>"011010100",
  7024=>"111111000",
  7025=>"110111101",
  7026=>"000100110",
  7027=>"010110001",
  7028=>"011100100",
  7029=>"000000000",
  7030=>"011111011",
  7031=>"000100110",
  7032=>"011001000",
  7033=>"110001011",
  7034=>"011111011",
  7035=>"001110010",
  7036=>"000001000",
  7037=>"001011101",
  7038=>"000000101",
  7039=>"111110000",
  7040=>"010001001",
  7041=>"101110000",
  7042=>"000010110",
  7043=>"110110010",
  7044=>"001100111",
  7045=>"101001000",
  7046=>"001100001",
  7047=>"001100010",
  7048=>"111100101",
  7049=>"110111001",
  7050=>"101011001",
  7051=>"110101111",
  7052=>"111010001",
  7053=>"000111000",
  7054=>"000111110",
  7055=>"111100111",
  7056=>"101100000",
  7057=>"100101001",
  7058=>"101010101",
  7059=>"111100001",
  7060=>"101011111",
  7061=>"111010111",
  7062=>"011111000",
  7063=>"010101110",
  7064=>"011101011",
  7065=>"111010101",
  7066=>"101101001",
  7067=>"000111110",
  7068=>"001110001",
  7069=>"111011010",
  7070=>"010001101",
  7071=>"110100000",
  7072=>"000010010",
  7073=>"011000011",
  7074=>"011000000",
  7075=>"101000101",
  7076=>"001001110",
  7077=>"000111010",
  7078=>"100001001",
  7079=>"010001000",
  7080=>"000111111",
  7081=>"100100000",
  7082=>"011111011",
  7083=>"000100010",
  7084=>"101000100",
  7085=>"101000111",
  7086=>"111101110",
  7087=>"000010000",
  7088=>"011010111",
  7089=>"110100110",
  7090=>"100100010",
  7091=>"011110001",
  7092=>"011111010",
  7093=>"011000000",
  7094=>"011011111",
  7095=>"011001001",
  7096=>"101100111",
  7097=>"111100100",
  7098=>"111011010",
  7099=>"010100000",
  7100=>"101110011",
  7101=>"000101111",
  7102=>"010000001",
  7103=>"110100111",
  7104=>"011100010",
  7105=>"001111101",
  7106=>"111000111",
  7107=>"111110010",
  7108=>"000000000",
  7109=>"110001011",
  7110=>"101110100",
  7111=>"010110111",
  7112=>"111011001",
  7113=>"100101110",
  7114=>"101010001",
  7115=>"111011010",
  7116=>"010011111",
  7117=>"110111001",
  7118=>"101011110",
  7119=>"011111100",
  7120=>"001011001",
  7121=>"011000011",
  7122=>"111001010",
  7123=>"110000000",
  7124=>"011111111",
  7125=>"011010010",
  7126=>"100011000",
  7127=>"100001001",
  7128=>"110101011",
  7129=>"011011011",
  7130=>"001011000",
  7131=>"010111100",
  7132=>"111011011",
  7133=>"100101010",
  7134=>"001001100",
  7135=>"000010001",
  7136=>"001111010",
  7137=>"001001011",
  7138=>"101111001",
  7139=>"000001101",
  7140=>"101100011",
  7141=>"000000011",
  7142=>"010000011",
  7143=>"101100100",
  7144=>"101001001",
  7145=>"000010101",
  7146=>"000100111",
  7147=>"111000011",
  7148=>"000011101",
  7149=>"111010010",
  7150=>"100101110",
  7151=>"011110001",
  7152=>"100111001",
  7153=>"011110100",
  7154=>"001101100",
  7155=>"111101111",
  7156=>"110101011",
  7157=>"000010001",
  7158=>"000011011",
  7159=>"101111001",
  7160=>"111110000",
  7161=>"111111100",
  7162=>"101010110",
  7163=>"011000100",
  7164=>"101010101",
  7165=>"000110110",
  7166=>"110110000",
  7167=>"110111011",
  7168=>"000010011",
  7169=>"101100000",
  7170=>"110010101",
  7171=>"111000001",
  7172=>"110101010",
  7173=>"100011110",
  7174=>"101100011",
  7175=>"010011100",
  7176=>"110111000",
  7177=>"010101111",
  7178=>"000100111",
  7179=>"100010111",
  7180=>"001001010",
  7181=>"000010001",
  7182=>"100100100",
  7183=>"010010001",
  7184=>"111110111",
  7185=>"101010100",
  7186=>"011010110",
  7187=>"011100001",
  7188=>"101001011",
  7189=>"000001110",
  7190=>"011111011",
  7191=>"010000100",
  7192=>"111010011",
  7193=>"000010001",
  7194=>"100100101",
  7195=>"100001000",
  7196=>"011100010",
  7197=>"110010001",
  7198=>"011111110",
  7199=>"011000111",
  7200=>"000010001",
  7201=>"001111010",
  7202=>"111111101",
  7203=>"101000101",
  7204=>"010111110",
  7205=>"001110000",
  7206=>"010110101",
  7207=>"101100100",
  7208=>"011000011",
  7209=>"100110010",
  7210=>"101111010",
  7211=>"100100110",
  7212=>"100011111",
  7213=>"010011100",
  7214=>"000100101",
  7215=>"111011001",
  7216=>"000100001",
  7217=>"101010001",
  7218=>"111011011",
  7219=>"001111001",
  7220=>"010000101",
  7221=>"011001111",
  7222=>"111001000",
  7223=>"001010111",
  7224=>"011001001",
  7225=>"001001111",
  7226=>"000111001",
  7227=>"100000000",
  7228=>"110101001",
  7229=>"110010010",
  7230=>"100111101",
  7231=>"000011101",
  7232=>"101000110",
  7233=>"101000001",
  7234=>"101100101",
  7235=>"000001000",
  7236=>"001100100",
  7237=>"010010000",
  7238=>"001010110",
  7239=>"011100011",
  7240=>"100110001",
  7241=>"010110100",
  7242=>"011001011",
  7243=>"101010110",
  7244=>"110001101",
  7245=>"000011110",
  7246=>"100110000",
  7247=>"111001110",
  7248=>"101111110",
  7249=>"110001011",
  7250=>"101111100",
  7251=>"001111011",
  7252=>"011000110",
  7253=>"010101100",
  7254=>"010010000",
  7255=>"101111000",
  7256=>"111101000",
  7257=>"010101101",
  7258=>"010001010",
  7259=>"100000101",
  7260=>"001100001",
  7261=>"110001000",
  7262=>"010010110",
  7263=>"001111011",
  7264=>"011001001",
  7265=>"000010011",
  7266=>"010111101",
  7267=>"010010011",
  7268=>"101100011",
  7269=>"001111010",
  7270=>"101010100",
  7271=>"100101010",
  7272=>"100000000",
  7273=>"100011101",
  7274=>"111011001",
  7275=>"111101010",
  7276=>"000111011",
  7277=>"101101010",
  7278=>"001000111",
  7279=>"110000100",
  7280=>"010111100",
  7281=>"011111101",
  7282=>"001111100",
  7283=>"111011010",
  7284=>"100110110",
  7285=>"110110000",
  7286=>"010010010",
  7287=>"101110010",
  7288=>"110101110",
  7289=>"010100001",
  7290=>"011001001",
  7291=>"111010011",
  7292=>"100110010",
  7293=>"011001011",
  7294=>"100101011",
  7295=>"111010010",
  7296=>"111110100",
  7297=>"001000111",
  7298=>"001110101",
  7299=>"100100000",
  7300=>"110001111",
  7301=>"000101010",
  7302=>"101100001",
  7303=>"011101101",
  7304=>"000010001",
  7305=>"010101001",
  7306=>"111000111",
  7307=>"010010001",
  7308=>"110111100",
  7309=>"110001011",
  7310=>"010010000",
  7311=>"110111100",
  7312=>"011011111",
  7313=>"001010100",
  7314=>"000001010",
  7315=>"000010011",
  7316=>"001010001",
  7317=>"001100100",
  7318=>"110010101",
  7319=>"001110101",
  7320=>"101101000",
  7321=>"101010000",
  7322=>"011010011",
  7323=>"010000001",
  7324=>"001000100",
  7325=>"000110000",
  7326=>"111001000",
  7327=>"100111110",
  7328=>"100111001",
  7329=>"010001011",
  7330=>"100101110",
  7331=>"101100011",
  7332=>"111001011",
  7333=>"011111110",
  7334=>"011001100",
  7335=>"001011001",
  7336=>"000001010",
  7337=>"000001100",
  7338=>"101101001",
  7339=>"110001100",
  7340=>"111111111",
  7341=>"100001100",
  7342=>"110101111",
  7343=>"110101100",
  7344=>"010010111",
  7345=>"011011011",
  7346=>"111101110",
  7347=>"000100111",
  7348=>"001011000",
  7349=>"100101011",
  7350=>"001011111",
  7351=>"110101000",
  7352=>"000101101",
  7353=>"000011101",
  7354=>"110000110",
  7355=>"001001000",
  7356=>"010001110",
  7357=>"111010111",
  7358=>"110111000",
  7359=>"010110100",
  7360=>"110101110",
  7361=>"100011110",
  7362=>"100101111",
  7363=>"111001000",
  7364=>"111001011",
  7365=>"111001100",
  7366=>"110111101",
  7367=>"100101011",
  7368=>"010110000",
  7369=>"000010010",
  7370=>"000110001",
  7371=>"110010110",
  7372=>"110111001",
  7373=>"100100100",
  7374=>"000100011",
  7375=>"100110010",
  7376=>"100011001",
  7377=>"100001100",
  7378=>"111101101",
  7379=>"000001001",
  7380=>"111110110",
  7381=>"111101011",
  7382=>"010110001",
  7383=>"011001001",
  7384=>"100011100",
  7385=>"111011010",
  7386=>"101100011",
  7387=>"001000101",
  7388=>"100011001",
  7389=>"001101010",
  7390=>"010100110",
  7391=>"101111011",
  7392=>"000101110",
  7393=>"011101101",
  7394=>"001101111",
  7395=>"010110010",
  7396=>"010000010",
  7397=>"010001101",
  7398=>"010010100",
  7399=>"010111101",
  7400=>"100010101",
  7401=>"011100001",
  7402=>"100101111",
  7403=>"011101110",
  7404=>"100001010",
  7405=>"000011001",
  7406=>"001110111",
  7407=>"010010100",
  7408=>"101111010",
  7409=>"101101000",
  7410=>"010010000",
  7411=>"110011101",
  7412=>"110100011",
  7413=>"001111010",
  7414=>"110100000",
  7415=>"000110010",
  7416=>"100000111",
  7417=>"110111000",
  7418=>"111100100",
  7419=>"001001101",
  7420=>"000110101",
  7421=>"100011100",
  7422=>"001000110",
  7423=>"010011110",
  7424=>"010111111",
  7425=>"101010111",
  7426=>"111000110",
  7427=>"001010110",
  7428=>"001100100",
  7429=>"000111000",
  7430=>"001011000",
  7431=>"100001101",
  7432=>"000000001",
  7433=>"001010010",
  7434=>"011111110",
  7435=>"010001000",
  7436=>"010001011",
  7437=>"100000110",
  7438=>"111111011",
  7439=>"110000000",
  7440=>"001100100",
  7441=>"000011001",
  7442=>"100100010",
  7443=>"001101010",
  7444=>"110000000",
  7445=>"000101010",
  7446=>"101001111",
  7447=>"101111111",
  7448=>"000010111",
  7449=>"111111111",
  7450=>"001011011",
  7451=>"011000001",
  7452=>"100010011",
  7453=>"100001001",
  7454=>"101110010",
  7455=>"101001101",
  7456=>"000001110",
  7457=>"110111001",
  7458=>"011111000",
  7459=>"011000100",
  7460=>"110111100",
  7461=>"001010101",
  7462=>"110110010",
  7463=>"011111110",
  7464=>"100111010",
  7465=>"101100111",
  7466=>"111000110",
  7467=>"010001100",
  7468=>"110101101",
  7469=>"100110000",
  7470=>"010101110",
  7471=>"100111011",
  7472=>"100110100",
  7473=>"100010010",
  7474=>"001010011",
  7475=>"110110100",
  7476=>"100100100",
  7477=>"011010000",
  7478=>"000110011",
  7479=>"100011110",
  7480=>"011010000",
  7481=>"100101001",
  7482=>"000010000",
  7483=>"011000110",
  7484=>"110100110",
  7485=>"100101101",
  7486=>"011001001",
  7487=>"101110111",
  7488=>"110011101",
  7489=>"101000000",
  7490=>"001011100",
  7491=>"000111001",
  7492=>"101101001",
  7493=>"010101101",
  7494=>"010100100",
  7495=>"100011001",
  7496=>"100100010",
  7497=>"100100100",
  7498=>"100111010",
  7499=>"001010010",
  7500=>"100111010",
  7501=>"001101001",
  7502=>"101111111",
  7503=>"100010100",
  7504=>"010010100",
  7505=>"111111011",
  7506=>"100001110",
  7507=>"001110110",
  7508=>"011010100",
  7509=>"001010001",
  7510=>"011101010",
  7511=>"110110000",
  7512=>"000101100",
  7513=>"010110001",
  7514=>"011100001",
  7515=>"011101001",
  7516=>"011011111",
  7517=>"001101000",
  7518=>"000000011",
  7519=>"101000010",
  7520=>"011111100",
  7521=>"010000100",
  7522=>"000101111",
  7523=>"001000000",
  7524=>"111100001",
  7525=>"000011010",
  7526=>"000100111",
  7527=>"110111011",
  7528=>"010101101",
  7529=>"000110011",
  7530=>"101000010",
  7531=>"000010100",
  7532=>"010110011",
  7533=>"110001011",
  7534=>"100101000",
  7535=>"110100000",
  7536=>"001110001",
  7537=>"000101010",
  7538=>"000000101",
  7539=>"011011111",
  7540=>"001100010",
  7541=>"011001100",
  7542=>"001100110",
  7543=>"011110110",
  7544=>"101101110",
  7545=>"110001011",
  7546=>"100110011",
  7547=>"111100100",
  7548=>"101101011",
  7549=>"111111001",
  7550=>"111000011",
  7551=>"000010000",
  7552=>"110000001",
  7553=>"001110111",
  7554=>"100001110",
  7555=>"110011100",
  7556=>"000101100",
  7557=>"110000101",
  7558=>"110010100",
  7559=>"010011101",
  7560=>"001111000",
  7561=>"010011100",
  7562=>"111000110",
  7563=>"001101111",
  7564=>"010000101",
  7565=>"000001100",
  7566=>"111010100",
  7567=>"100110101",
  7568=>"110100100",
  7569=>"010000011",
  7570=>"100001110",
  7571=>"100000111",
  7572=>"111101010",
  7573=>"010011111",
  7574=>"011100010",
  7575=>"110001000",
  7576=>"101011110",
  7577=>"000111110",
  7578=>"010101001",
  7579=>"001000011",
  7580=>"101001101",
  7581=>"010101100",
  7582=>"010101111",
  7583=>"110001110",
  7584=>"100000000",
  7585=>"000001101",
  7586=>"000011100",
  7587=>"001011101",
  7588=>"111101100",
  7589=>"000000100",
  7590=>"100001010",
  7591=>"101100010",
  7592=>"001001110",
  7593=>"011101010",
  7594=>"100000101",
  7595=>"111010011",
  7596=>"110000111",
  7597=>"100011010",
  7598=>"100101010",
  7599=>"110011010",
  7600=>"111010111",
  7601=>"011100010",
  7602=>"101011010",
  7603=>"000010001",
  7604=>"010000100",
  7605=>"111001000",
  7606=>"110011010",
  7607=>"000100000",
  7608=>"001110011",
  7609=>"000011010",
  7610=>"000111101",
  7611=>"100011010",
  7612=>"100100110",
  7613=>"011100010",
  7614=>"111010000",
  7615=>"111111000",
  7616=>"010001010",
  7617=>"010111101",
  7618=>"101111110",
  7619=>"100100110",
  7620=>"100010011",
  7621=>"000111111",
  7622=>"000000111",
  7623=>"011010111",
  7624=>"110101110",
  7625=>"010011101",
  7626=>"000100111",
  7627=>"111101111",
  7628=>"001100010",
  7629=>"100011101",
  7630=>"001110000",
  7631=>"000111001",
  7632=>"110100011",
  7633=>"110111111",
  7634=>"100000101",
  7635=>"010100000",
  7636=>"100011111",
  7637=>"000100111",
  7638=>"001011101",
  7639=>"111000111",
  7640=>"001111001",
  7641=>"101011010",
  7642=>"101111001",
  7643=>"101111001",
  7644=>"110101000",
  7645=>"011001001",
  7646=>"111100011",
  7647=>"010111010",
  7648=>"100100011",
  7649=>"011011101",
  7650=>"011011011",
  7651=>"010011101",
  7652=>"111101100",
  7653=>"001001001",
  7654=>"110110101",
  7655=>"010011111",
  7656=>"100110101",
  7657=>"000001111",
  7658=>"010100001",
  7659=>"100111011",
  7660=>"101000111",
  7661=>"011011011",
  7662=>"100001110",
  7663=>"100011011",
  7664=>"111101111",
  7665=>"001011101",
  7666=>"001001000",
  7667=>"110111001",
  7668=>"000100111",
  7669=>"000000110",
  7670=>"111111011",
  7671=>"100100111",
  7672=>"000000000",
  7673=>"101011111",
  7674=>"100000111",
  7675=>"010110001",
  7676=>"110101101",
  7677=>"100011001",
  7678=>"100100010",
  7679=>"000000001",
  7680=>"111110011",
  7681=>"110011111",
  7682=>"111011010",
  7683=>"101100011",
  7684=>"110110110",
  7685=>"010011111",
  7686=>"111110000",
  7687=>"110000101",
  7688=>"010000101",
  7689=>"100000011",
  7690=>"000110101",
  7691=>"001101010",
  7692=>"001110110",
  7693=>"011011011",
  7694=>"100000000",
  7695=>"100100010",
  7696=>"011101000",
  7697=>"001000001",
  7698=>"011100010",
  7699=>"000100000",
  7700=>"100000010",
  7701=>"111000001",
  7702=>"000111110",
  7703=>"000001100",
  7704=>"101011111",
  7705=>"010111000",
  7706=>"101001000",
  7707=>"100101110",
  7708=>"000010010",
  7709=>"110010110",
  7710=>"111110011",
  7711=>"100001010",
  7712=>"010111110",
  7713=>"011101100",
  7714=>"000100101",
  7715=>"011101110",
  7716=>"111001000",
  7717=>"001100110",
  7718=>"010001100",
  7719=>"000100100",
  7720=>"001001111",
  7721=>"011111101",
  7722=>"000100100",
  7723=>"001010100",
  7724=>"010110100",
  7725=>"010000000",
  7726=>"110001000",
  7727=>"000100100",
  7728=>"101100001",
  7729=>"111111011",
  7730=>"000000111",
  7731=>"010010110",
  7732=>"011011000",
  7733=>"010010001",
  7734=>"110010100",
  7735=>"001111100",
  7736=>"000111110",
  7737=>"001110000",
  7738=>"101100111",
  7739=>"001000111",
  7740=>"111011110",
  7741=>"001011011",
  7742=>"000001010",
  7743=>"100011011",
  7744=>"110010100",
  7745=>"111110001",
  7746=>"000011000",
  7747=>"010101010",
  7748=>"100101111",
  7749=>"101000110",
  7750=>"011100001",
  7751=>"110001110",
  7752=>"001000010",
  7753=>"111101101",
  7754=>"000100000",
  7755=>"100011010",
  7756=>"011001001",
  7757=>"111000111",
  7758=>"110110101",
  7759=>"100101111",
  7760=>"010100110",
  7761=>"000000101",
  7762=>"101100010",
  7763=>"101010111",
  7764=>"100000010",
  7765=>"001000010",
  7766=>"010001010",
  7767=>"101001100",
  7768=>"000101100",
  7769=>"101001011",
  7770=>"101111001",
  7771=>"101100000",
  7772=>"110111101",
  7773=>"000000000",
  7774=>"111100101",
  7775=>"001001111",
  7776=>"011000011",
  7777=>"110010011",
  7778=>"011110110",
  7779=>"100001001",
  7780=>"110100011",
  7781=>"010000000",
  7782=>"111110110",
  7783=>"000010110",
  7784=>"010101001",
  7785=>"001011000",
  7786=>"000111010",
  7787=>"010110110",
  7788=>"001010110",
  7789=>"000110001",
  7790=>"101011000",
  7791=>"010100001",
  7792=>"101111010",
  7793=>"011000010",
  7794=>"111001010",
  7795=>"100010010",
  7796=>"110000011",
  7797=>"010111010",
  7798=>"001010010",
  7799=>"101011001",
  7800=>"111011011",
  7801=>"000001000",
  7802=>"100110110",
  7803=>"001010010",
  7804=>"111001101",
  7805=>"011111101",
  7806=>"110100111",
  7807=>"101110100",
  7808=>"001000010",
  7809=>"011111101",
  7810=>"001011111",
  7811=>"101010110",
  7812=>"011110111",
  7813=>"001111101",
  7814=>"011011101",
  7815=>"100100000",
  7816=>"011110010",
  7817=>"000010111",
  7818=>"011001100",
  7819=>"100001011",
  7820=>"100000000",
  7821=>"011000001",
  7822=>"011010100",
  7823=>"001000001",
  7824=>"110100110",
  7825=>"101101111",
  7826=>"101100101",
  7827=>"111001100",
  7828=>"011110100",
  7829=>"100011111",
  7830=>"000101110",
  7831=>"101111110",
  7832=>"101011011",
  7833=>"110101110",
  7834=>"111000101",
  7835=>"011110011",
  7836=>"011111101",
  7837=>"001010011",
  7838=>"110011110",
  7839=>"010111100",
  7840=>"001011111",
  7841=>"001110010",
  7842=>"011111110",
  7843=>"011100001",
  7844=>"111111011",
  7845=>"011111111",
  7846=>"000101101",
  7847=>"101001010",
  7848=>"010100010",
  7849=>"000111000",
  7850=>"010100110",
  7851=>"100000010",
  7852=>"000011100",
  7853=>"010110111",
  7854=>"011101001",
  7855=>"011011100",
  7856=>"001110010",
  7857=>"001110100",
  7858=>"011010100",
  7859=>"010101010",
  7860=>"110100000",
  7861=>"111010111",
  7862=>"010111101",
  7863=>"111001011",
  7864=>"101110100",
  7865=>"110101110",
  7866=>"101100001",
  7867=>"101000010",
  7868=>"100101000",
  7869=>"111010000",
  7870=>"111010000",
  7871=>"000001000",
  7872=>"000010111",
  7873=>"010110011",
  7874=>"010101100",
  7875=>"100110110",
  7876=>"110111101",
  7877=>"000110000",
  7878=>"111100011",
  7879=>"010010001",
  7880=>"000100001",
  7881=>"000100001",
  7882=>"001010101",
  7883=>"100111110",
  7884=>"011000011",
  7885=>"000110010",
  7886=>"010001100",
  7887=>"011101101",
  7888=>"111110100",
  7889=>"000001100",
  7890=>"000010010",
  7891=>"000100111",
  7892=>"011010000",
  7893=>"101011011",
  7894=>"000101001",
  7895=>"001100110",
  7896=>"010111110",
  7897=>"100010101",
  7898=>"010000101",
  7899=>"010000100",
  7900=>"010000100",
  7901=>"111100100",
  7902=>"001101011",
  7903=>"101111111",
  7904=>"001000010",
  7905=>"110011111",
  7906=>"010001010",
  7907=>"001110100",
  7908=>"000010111",
  7909=>"010010100",
  7910=>"001100110",
  7911=>"110010101",
  7912=>"101010110",
  7913=>"100010101",
  7914=>"010010011",
  7915=>"110101010",
  7916=>"101100111",
  7917=>"000010011",
  7918=>"001010111",
  7919=>"010101010",
  7920=>"111000001",
  7921=>"111000000",
  7922=>"101010001",
  7923=>"011011101",
  7924=>"010001001",
  7925=>"000101010",
  7926=>"110011111",
  7927=>"010010001",
  7928=>"001000100",
  7929=>"011101011",
  7930=>"011010000",
  7931=>"000100001",
  7932=>"101000001",
  7933=>"100001111",
  7934=>"011110110",
  7935=>"011000111",
  7936=>"011110000",
  7937=>"101011000",
  7938=>"111100101",
  7939=>"100000101",
  7940=>"010100111",
  7941=>"000110010",
  7942=>"001111000",
  7943=>"001000111",
  7944=>"111111111",
  7945=>"101001101",
  7946=>"010110101",
  7947=>"110001111",
  7948=>"110011110",
  7949=>"111100110",
  7950=>"101110110",
  7951=>"100101000",
  7952=>"110100000",
  7953=>"111010101",
  7954=>"100111101",
  7955=>"111011110",
  7956=>"100111111",
  7957=>"001011111",
  7958=>"110101110",
  7959=>"110100010",
  7960=>"011100110",
  7961=>"011000001",
  7962=>"111000110",
  7963=>"110111110",
  7964=>"100111110",
  7965=>"001010101",
  7966=>"010000100",
  7967=>"111100001",
  7968=>"111000101",
  7969=>"000001110",
  7970=>"100000000",
  7971=>"000010000",
  7972=>"000001001",
  7973=>"010011101",
  7974=>"101001111",
  7975=>"000000101",
  7976=>"111011001",
  7977=>"010100110",
  7978=>"110000010",
  7979=>"111100010",
  7980=>"000011001",
  7981=>"100111111",
  7982=>"001100011",
  7983=>"100001111",
  7984=>"010100101",
  7985=>"001000111",
  7986=>"000000101",
  7987=>"000000001",
  7988=>"100110010",
  7989=>"111010011",
  7990=>"100100001",
  7991=>"011001010",
  7992=>"101100000",
  7993=>"010100101",
  7994=>"100011000",
  7995=>"010001011",
  7996=>"001110101",
  7997=>"000110000",
  7998=>"010011101",
  7999=>"001001110",
  8000=>"110011010",
  8001=>"111110100",
  8002=>"110101001",
  8003=>"101010011",
  8004=>"100011001",
  8005=>"001101011",
  8006=>"000001100",
  8007=>"110010110",
  8008=>"010001101",
  8009=>"011011110",
  8010=>"001111100",
  8011=>"111101000",
  8012=>"001001111",
  8013=>"100100110",
  8014=>"000000001",
  8015=>"011011110",
  8016=>"111000000",
  8017=>"110011101",
  8018=>"100001010",
  8019=>"000101110",
  8020=>"100000000",
  8021=>"000110111",
  8022=>"101110011",
  8023=>"001000010",
  8024=>"000000100",
  8025=>"011111111",
  8026=>"111010011",
  8027=>"001111100",
  8028=>"011010111",
  8029=>"100010101",
  8030=>"001010111",
  8031=>"000100010",
  8032=>"101101101",
  8033=>"100101100",
  8034=>"111100101",
  8035=>"100011101",
  8036=>"101001110",
  8037=>"001001010",
  8038=>"010011111",
  8039=>"000000011",
  8040=>"011011001",
  8041=>"101111010",
  8042=>"100011001",
  8043=>"101000010",
  8044=>"010010011",
  8045=>"111000010",
  8046=>"000111100",
  8047=>"010010001",
  8048=>"000110001",
  8049=>"000001100",
  8050=>"101100101",
  8051=>"111100010",
  8052=>"010101010",
  8053=>"010001100",
  8054=>"110110100",
  8055=>"101101001",
  8056=>"101101001",
  8057=>"011011100",
  8058=>"011110001",
  8059=>"000000110",
  8060=>"000000010",
  8061=>"110011100",
  8062=>"011111111",
  8063=>"001110111",
  8064=>"000010011",
  8065=>"011110011",
  8066=>"000000110",
  8067=>"000100011",
  8068=>"011100100",
  8069=>"110011011",
  8070=>"111110111",
  8071=>"110110001",
  8072=>"011010011",
  8073=>"100011000",
  8074=>"011100000",
  8075=>"111011100",
  8076=>"110000100",
  8077=>"101010110",
  8078=>"011100001",
  8079=>"100101010",
  8080=>"000001001",
  8081=>"101010101",
  8082=>"000010011",
  8083=>"011000110",
  8084=>"110000101",
  8085=>"001100001",
  8086=>"110110010",
  8087=>"001011100",
  8088=>"111110111",
  8089=>"111000100",
  8090=>"001010000",
  8091=>"110010100",
  8092=>"111001010",
  8093=>"011110001",
  8094=>"110000111",
  8095=>"100001000",
  8096=>"100011101",
  8097=>"100111001",
  8098=>"000100111",
  8099=>"111000011",
  8100=>"000000000",
  8101=>"100001000",
  8102=>"101001000",
  8103=>"011011101",
  8104=>"010001100",
  8105=>"011110100",
  8106=>"101110100",
  8107=>"011010001",
  8108=>"101101100",
  8109=>"000111000",
  8110=>"101100000",
  8111=>"111001000",
  8112=>"111101000",
  8113=>"110000101",
  8114=>"101000100",
  8115=>"001010011",
  8116=>"111010010",
  8117=>"101001100",
  8118=>"100101110",
  8119=>"011011101",
  8120=>"000101000",
  8121=>"000010001",
  8122=>"100010011",
  8123=>"011110011",
  8124=>"111001101",
  8125=>"100110000",
  8126=>"001000110",
  8127=>"010110110",
  8128=>"001001111",
  8129=>"001011010",
  8130=>"101111111",
  8131=>"100111100",
  8132=>"000000001",
  8133=>"110011011",
  8134=>"111101001",
  8135=>"110100111",
  8136=>"000101000",
  8137=>"010111100",
  8138=>"000011110",
  8139=>"011110111",
  8140=>"100001000",
  8141=>"000000111",
  8142=>"000110010",
  8143=>"010000001",
  8144=>"011100011",
  8145=>"100011000",
  8146=>"100011011",
  8147=>"000101000",
  8148=>"101010000",
  8149=>"110001011",
  8150=>"111100100",
  8151=>"111100110",
  8152=>"100001010",
  8153=>"010010101",
  8154=>"110000010",
  8155=>"011000110",
  8156=>"011101110",
  8157=>"101000101",
  8158=>"101110001",
  8159=>"110100111",
  8160=>"011101111",
  8161=>"101101011",
  8162=>"100101100",
  8163=>"011101000",
  8164=>"011000000",
  8165=>"010101101",
  8166=>"111011111",
  8167=>"101100011",
  8168=>"010110011",
  8169=>"011110110",
  8170=>"110000010",
  8171=>"101101101",
  8172=>"110010111",
  8173=>"011100110",
  8174=>"010010001",
  8175=>"000110000",
  8176=>"100111000",
  8177=>"001101010",
  8178=>"011001111",
  8179=>"100110100",
  8180=>"100111101",
  8181=>"100010100",
  8182=>"110000110",
  8183=>"010001100",
  8184=>"001110001",
  8185=>"111110101",
  8186=>"011010111",
  8187=>"000110000",
  8188=>"000000111",
  8189=>"011001100",
  8190=>"000101011",
  8191=>"010001101",
  8192=>"101100111",
  8193=>"001001100",
  8194=>"000010110",
  8195=>"010000111",
  8196=>"001111101",
  8197=>"110110001",
  8198=>"010010100",
  8199=>"010001010",
  8200=>"010011001",
  8201=>"011010000",
  8202=>"110100000",
  8203=>"100110100",
  8204=>"101111111",
  8205=>"100100110",
  8206=>"000000001",
  8207=>"111100111",
  8208=>"001101110",
  8209=>"000100111",
  8210=>"111111110",
  8211=>"110110000",
  8212=>"001001110",
  8213=>"001001110",
  8214=>"110111111",
  8215=>"100000110",
  8216=>"110101101",
  8217=>"000111101",
  8218=>"101011000",
  8219=>"101001011",
  8220=>"100000000",
  8221=>"010000010",
  8222=>"000010001",
  8223=>"111100111",
  8224=>"101101110",
  8225=>"110010001",
  8226=>"100101111",
  8227=>"100101010",
  8228=>"010110110",
  8229=>"010011000",
  8230=>"000010100",
  8231=>"010010001",
  8232=>"010000110",
  8233=>"000000010",
  8234=>"110100000",
  8235=>"000110001",
  8236=>"001011100",
  8237=>"110101001",
  8238=>"100101001",
  8239=>"100101011",
  8240=>"111111101",
  8241=>"110110001",
  8242=>"100010101",
  8243=>"011110111",
  8244=>"000000100",
  8245=>"101011110",
  8246=>"001111011",
  8247=>"101001111",
  8248=>"101101111",
  8249=>"010100100",
  8250=>"011001110",
  8251=>"101111011",
  8252=>"101000111",
  8253=>"000010110",
  8254=>"100100110",
  8255=>"010110000",
  8256=>"111111101",
  8257=>"100010011",
  8258=>"110010111",
  8259=>"111111011",
  8260=>"001101111",
  8261=>"101000101",
  8262=>"100000000",
  8263=>"010000000",
  8264=>"010110111",
  8265=>"111000111",
  8266=>"111010111",
  8267=>"101001000",
  8268=>"110001111",
  8269=>"000110011",
  8270=>"110000000",
  8271=>"101100001",
  8272=>"100100010",
  8273=>"011000010",
  8274=>"101010010",
  8275=>"110010011",
  8276=>"111111001",
  8277=>"001001001",
  8278=>"000010000",
  8279=>"001001011",
  8280=>"111011110",
  8281=>"100001101",
  8282=>"111000100",
  8283=>"100011011",
  8284=>"011001111",
  8285=>"001001100",
  8286=>"000000101",
  8287=>"111101010",
  8288=>"100111101",
  8289=>"000001111",
  8290=>"111101111",
  8291=>"101001110",
  8292=>"011111001",
  8293=>"101001000",
  8294=>"010110000",
  8295=>"000011111",
  8296=>"110110100",
  8297=>"010110111",
  8298=>"001100110",
  8299=>"101001000",
  8300=>"011100111",
  8301=>"110110110",
  8302=>"101001010",
  8303=>"001000101",
  8304=>"110000001",
  8305=>"111111010",
  8306=>"111011101",
  8307=>"111000101",
  8308=>"100101000",
  8309=>"000001001",
  8310=>"011101000",
  8311=>"110100101",
  8312=>"001100110",
  8313=>"010010001",
  8314=>"111101010",
  8315=>"011001011",
  8316=>"000100110",
  8317=>"011010111",
  8318=>"011000110",
  8319=>"111100110",
  8320=>"010001110",
  8321=>"001100011",
  8322=>"000110100",
  8323=>"000000011",
  8324=>"000101000",
  8325=>"011000001",
  8326=>"110110001",
  8327=>"011100111",
  8328=>"100101000",
  8329=>"100111111",
  8330=>"011111011",
  8331=>"000000011",
  8332=>"000111100",
  8333=>"001010010",
  8334=>"101000110",
  8335=>"001011100",
  8336=>"111100111",
  8337=>"111101010",
  8338=>"110111100",
  8339=>"111010101",
  8340=>"010001011",
  8341=>"001011000",
  8342=>"001111000",
  8343=>"101100000",
  8344=>"110100110",
  8345=>"001110001",
  8346=>"100110111",
  8347=>"110000000",
  8348=>"011100011",
  8349=>"101111111",
  8350=>"111000111",
  8351=>"111001001",
  8352=>"011011101",
  8353=>"101110000",
  8354=>"011100011",
  8355=>"000100011",
  8356=>"011011101",
  8357=>"101011001",
  8358=>"110111111",
  8359=>"110101000",
  8360=>"001001001",
  8361=>"100001110",
  8362=>"001111101",
  8363=>"001111111",
  8364=>"000011001",
  8365=>"111001111",
  8366=>"010101101",
  8367=>"011001001",
  8368=>"001001110",
  8369=>"101110011",
  8370=>"011111101",
  8371=>"010011100",
  8372=>"111110000",
  8373=>"111100110",
  8374=>"010011011",
  8375=>"010000100",
  8376=>"110101001",
  8377=>"111100000",
  8378=>"100001000",
  8379=>"000100100",
  8380=>"111101101",
  8381=>"100001111",
  8382=>"000001111",
  8383=>"111000001",
  8384=>"011111010",
  8385=>"101100100",
  8386=>"111010111",
  8387=>"010111010",
  8388=>"101101001",
  8389=>"010000000",
  8390=>"101111100",
  8391=>"110011100",
  8392=>"010110101",
  8393=>"010000101",
  8394=>"010110111",
  8395=>"110111010",
  8396=>"011111110",
  8397=>"000000010",
  8398=>"011111000",
  8399=>"100111010",
  8400=>"001011011",
  8401=>"001101000",
  8402=>"001100001",
  8403=>"100100101",
  8404=>"010111110",
  8405=>"001101000",
  8406=>"000101110",
  8407=>"011100110",
  8408=>"011110111",
  8409=>"111110000",
  8410=>"000101001",
  8411=>"101100110",
  8412=>"011010010",
  8413=>"010001010",
  8414=>"000010110",
  8415=>"010111000",
  8416=>"101100010",
  8417=>"000100100",
  8418=>"001111101",
  8419=>"000100101",
  8420=>"110000111",
  8421=>"110111100",
  8422=>"111000000",
  8423=>"111111101",
  8424=>"100100101",
  8425=>"000110111",
  8426=>"111101101",
  8427=>"000000001",
  8428=>"011001101",
  8429=>"100010100",
  8430=>"101110000",
  8431=>"011101110",
  8432=>"011101010",
  8433=>"001111111",
  8434=>"000111010",
  8435=>"111011011",
  8436=>"010111011",
  8437=>"100101101",
  8438=>"110111111",
  8439=>"001100000",
  8440=>"010110111",
  8441=>"101011100",
  8442=>"010110010",
  8443=>"100001110",
  8444=>"001010001",
  8445=>"111010001",
  8446=>"110010010",
  8447=>"100011001",
  8448=>"011000111",
  8449=>"111110111",
  8450=>"010010010",
  8451=>"101000100",
  8452=>"000010011",
  8453=>"000010111",
  8454=>"101011100",
  8455=>"101001001",
  8456=>"010101000",
  8457=>"010111111",
  8458=>"000011111",
  8459=>"011000010",
  8460=>"011000111",
  8461=>"000000110",
  8462=>"001001101",
  8463=>"001011101",
  8464=>"001011000",
  8465=>"111100111",
  8466=>"001111111",
  8467=>"011010111",
  8468=>"000010001",
  8469=>"010001110",
  8470=>"111001100",
  8471=>"110000110",
  8472=>"011000110",
  8473=>"111010111",
  8474=>"010100100",
  8475=>"000100110",
  8476=>"000110001",
  8477=>"110100011",
  8478=>"011101110",
  8479=>"001000000",
  8480=>"010001110",
  8481=>"100011001",
  8482=>"001000101",
  8483=>"110011001",
  8484=>"001010001",
  8485=>"000000010",
  8486=>"101000010",
  8487=>"110010000",
  8488=>"010101100",
  8489=>"010100011",
  8490=>"001010001",
  8491=>"100111001",
  8492=>"000001001",
  8493=>"111111101",
  8494=>"011000101",
  8495=>"011010001",
  8496=>"100111001",
  8497=>"110101110",
  8498=>"100110010",
  8499=>"111101111",
  8500=>"110110110",
  8501=>"000110000",
  8502=>"110111111",
  8503=>"101111101",
  8504=>"111111110",
  8505=>"000111100",
  8506=>"000000011",
  8507=>"001111010",
  8508=>"110100000",
  8509=>"110111110",
  8510=>"100101101",
  8511=>"000010010",
  8512=>"110010001",
  8513=>"011110111",
  8514=>"011100000",
  8515=>"011111010",
  8516=>"100100011",
  8517=>"000100110",
  8518=>"011000001",
  8519=>"100001000",
  8520=>"001011000",
  8521=>"101011000",
  8522=>"100100000",
  8523=>"000000000",
  8524=>"000010011",
  8525=>"011110100",
  8526=>"111110000",
  8527=>"111011001",
  8528=>"011001101",
  8529=>"101000101",
  8530=>"100101111",
  8531=>"111101101",
  8532=>"100100000",
  8533=>"000110011",
  8534=>"101001001",
  8535=>"111010100",
  8536=>"101101000",
  8537=>"000101101",
  8538=>"010100111",
  8539=>"100000100",
  8540=>"011101111",
  8541=>"111011110",
  8542=>"111111111",
  8543=>"001100001",
  8544=>"000010100",
  8545=>"011100100",
  8546=>"111101101",
  8547=>"010111000",
  8548=>"000110011",
  8549=>"101011110",
  8550=>"110111001",
  8551=>"110100011",
  8552=>"101001001",
  8553=>"000000011",
  8554=>"000010010",
  8555=>"000000110",
  8556=>"100101010",
  8557=>"010010101",
  8558=>"101001010",
  8559=>"010111101",
  8560=>"000110110",
  8561=>"110100111",
  8562=>"010000011",
  8563=>"000010110",
  8564=>"101110001",
  8565=>"011010000",
  8566=>"010101111",
  8567=>"010010011",
  8568=>"110100110",
  8569=>"000100111",
  8570=>"011000010",
  8571=>"111111101",
  8572=>"011000000",
  8573=>"111111101",
  8574=>"000010000",
  8575=>"110110111",
  8576=>"111000110",
  8577=>"010011101",
  8578=>"000000101",
  8579=>"010001010",
  8580=>"101100110",
  8581=>"000111110",
  8582=>"000111010",
  8583=>"101101110",
  8584=>"011011110",
  8585=>"110101101",
  8586=>"100100111",
  8587=>"101100010",
  8588=>"111010011",
  8589=>"000100001",
  8590=>"000001110",
  8591=>"100000101",
  8592=>"111000100",
  8593=>"100000001",
  8594=>"001101100",
  8595=>"101111001",
  8596=>"001101010",
  8597=>"101100111",
  8598=>"110111000",
  8599=>"110100010",
  8600=>"000100110",
  8601=>"010100111",
  8602=>"001011101",
  8603=>"000101000",
  8604=>"100001111",
  8605=>"101000010",
  8606=>"101111010",
  8607=>"000010100",
  8608=>"000011011",
  8609=>"010001001",
  8610=>"101111111",
  8611=>"100000000",
  8612=>"010110100",
  8613=>"100111010",
  8614=>"001001010",
  8615=>"111110000",
  8616=>"000100110",
  8617=>"100110001",
  8618=>"110000001",
  8619=>"110101111",
  8620=>"101001010",
  8621=>"111010101",
  8622=>"000001111",
  8623=>"001101000",
  8624=>"110011001",
  8625=>"111101100",
  8626=>"000010101",
  8627=>"111110100",
  8628=>"100001001",
  8629=>"010101010",
  8630=>"100011010",
  8631=>"111101010",
  8632=>"110110011",
  8633=>"000101111",
  8634=>"000011000",
  8635=>"110011010",
  8636=>"110000101",
  8637=>"010000000",
  8638=>"101000000",
  8639=>"111011101",
  8640=>"000100110",
  8641=>"110111011",
  8642=>"000111010",
  8643=>"111001110",
  8644=>"101110011",
  8645=>"101101111",
  8646=>"111101111",
  8647=>"001001101",
  8648=>"000001110",
  8649=>"100101010",
  8650=>"111110111",
  8651=>"111011110",
  8652=>"101100100",
  8653=>"000111111",
  8654=>"100001110",
  8655=>"110101111",
  8656=>"001111100",
  8657=>"111111110",
  8658=>"110111100",
  8659=>"001001110",
  8660=>"011010111",
  8661=>"111100011",
  8662=>"110100000",
  8663=>"010011110",
  8664=>"110001011",
  8665=>"111001000",
  8666=>"100011001",
  8667=>"101101110",
  8668=>"111000000",
  8669=>"111110011",
  8670=>"000111001",
  8671=>"100110100",
  8672=>"111101000",
  8673=>"010011000",
  8674=>"110011111",
  8675=>"101100011",
  8676=>"011100101",
  8677=>"110110101",
  8678=>"011110001",
  8679=>"100010100",
  8680=>"000110001",
  8681=>"001001000",
  8682=>"010000100",
  8683=>"101011000",
  8684=>"101001000",
  8685=>"000000000",
  8686=>"111110001",
  8687=>"101000000",
  8688=>"001100001",
  8689=>"110100110",
  8690=>"000101001",
  8691=>"000111101",
  8692=>"110111010",
  8693=>"010010001",
  8694=>"010111000",
  8695=>"111110111",
  8696=>"111101101",
  8697=>"110010111",
  8698=>"110110001",
  8699=>"101111011",
  8700=>"001101110",
  8701=>"110100101",
  8702=>"010100110",
  8703=>"001110110",
  8704=>"000101110",
  8705=>"010111110",
  8706=>"001011101",
  8707=>"000110101",
  8708=>"101100000",
  8709=>"101101101",
  8710=>"111110101",
  8711=>"100110011",
  8712=>"111110010",
  8713=>"011101010",
  8714=>"111011001",
  8715=>"101010001",
  8716=>"111100110",
  8717=>"100111011",
  8718=>"000001100",
  8719=>"011101001",
  8720=>"111101010",
  8721=>"111110010",
  8722=>"111001010",
  8723=>"111000101",
  8724=>"001010001",
  8725=>"111000110",
  8726=>"111000110",
  8727=>"110011110",
  8728=>"101011111",
  8729=>"111110011",
  8730=>"011101101",
  8731=>"011101001",
  8732=>"001000010",
  8733=>"000000000",
  8734=>"110011001",
  8735=>"111101010",
  8736=>"000010101",
  8737=>"001010101",
  8738=>"111000110",
  8739=>"001110111",
  8740=>"110010010",
  8741=>"111010010",
  8742=>"111111100",
  8743=>"111111001",
  8744=>"101111111",
  8745=>"011100101",
  8746=>"111111111",
  8747=>"010001110",
  8748=>"101001111",
  8749=>"110100000",
  8750=>"011100000",
  8751=>"000011011",
  8752=>"111101111",
  8753=>"100010110",
  8754=>"000100111",
  8755=>"000000001",
  8756=>"101100001",
  8757=>"010101110",
  8758=>"110100011",
  8759=>"001011011",
  8760=>"111111110",
  8761=>"100111100",
  8762=>"000000010",
  8763=>"010001001",
  8764=>"100001001",
  8765=>"001100111",
  8766=>"011100101",
  8767=>"100100001",
  8768=>"111001011",
  8769=>"110100010",
  8770=>"111001011",
  8771=>"000011101",
  8772=>"111101111",
  8773=>"011100111",
  8774=>"000111110",
  8775=>"011000011",
  8776=>"110100010",
  8777=>"101000101",
  8778=>"011101001",
  8779=>"111010001",
  8780=>"000011000",
  8781=>"000001100",
  8782=>"110101101",
  8783=>"001100010",
  8784=>"010001000",
  8785=>"001010100",
  8786=>"000010001",
  8787=>"011011011",
  8788=>"110000110",
  8789=>"010001010",
  8790=>"111101100",
  8791=>"010100110",
  8792=>"011000111",
  8793=>"000000110",
  8794=>"000001100",
  8795=>"100001010",
  8796=>"100001101",
  8797=>"000000110",
  8798=>"111010111",
  8799=>"010110111",
  8800=>"010110001",
  8801=>"011110101",
  8802=>"101011000",
  8803=>"110000010",
  8804=>"110010110",
  8805=>"110101010",
  8806=>"001101011",
  8807=>"010001010",
  8808=>"000110111",
  8809=>"010101011",
  8810=>"101001111",
  8811=>"000111011",
  8812=>"000010111",
  8813=>"010001101",
  8814=>"111111011",
  8815=>"000011010",
  8816=>"101001111",
  8817=>"010111001",
  8818=>"111110111",
  8819=>"001111100",
  8820=>"010010011",
  8821=>"010011000",
  8822=>"000110000",
  8823=>"000000110",
  8824=>"011011101",
  8825=>"101000101",
  8826=>"111011000",
  8827=>"110101001",
  8828=>"000000011",
  8829=>"011100111",
  8830=>"101011011",
  8831=>"000101011",
  8832=>"101010011",
  8833=>"000000000",
  8834=>"111001111",
  8835=>"110110001",
  8836=>"001010001",
  8837=>"111111010",
  8838=>"111101110",
  8839=>"000110000",
  8840=>"110101101",
  8841=>"011000000",
  8842=>"010010011",
  8843=>"100111010",
  8844=>"001010101",
  8845=>"011010100",
  8846=>"111100100",
  8847=>"101000100",
  8848=>"100011101",
  8849=>"011010011",
  8850=>"101100001",
  8851=>"110111100",
  8852=>"001011001",
  8853=>"101110000",
  8854=>"001101010",
  8855=>"110000011",
  8856=>"001100001",
  8857=>"111100010",
  8858=>"010001110",
  8859=>"000000000",
  8860=>"001101101",
  8861=>"000000100",
  8862=>"001110111",
  8863=>"011101101",
  8864=>"010110110",
  8865=>"111011100",
  8866=>"000100110",
  8867=>"001011111",
  8868=>"011111110",
  8869=>"000111010",
  8870=>"110010011",
  8871=>"100001000",
  8872=>"010001111",
  8873=>"000110101",
  8874=>"001000011",
  8875=>"001001001",
  8876=>"100001010",
  8877=>"000101110",
  8878=>"101001000",
  8879=>"001110000",
  8880=>"000000001",
  8881=>"000000001",
  8882=>"111011111",
  8883=>"011101010",
  8884=>"110010101",
  8885=>"001100000",
  8886=>"100111011",
  8887=>"111101101",
  8888=>"010111111",
  8889=>"010100011",
  8890=>"110110000",
  8891=>"010000110",
  8892=>"111000111",
  8893=>"100100010",
  8894=>"001000010",
  8895=>"110000110",
  8896=>"000100001",
  8897=>"000101011",
  8898=>"101000001",
  8899=>"111100111",
  8900=>"011001110",
  8901=>"100101001",
  8902=>"001001110",
  8903=>"011111101",
  8904=>"110000000",
  8905=>"110010010",
  8906=>"010000001",
  8907=>"110001110",
  8908=>"010110100",
  8909=>"011101011",
  8910=>"011001011",
  8911=>"111111011",
  8912=>"111111111",
  8913=>"111011010",
  8914=>"110010010",
  8915=>"100000001",
  8916=>"100110101",
  8917=>"101011001",
  8918=>"100100011",
  8919=>"000011111",
  8920=>"101101110",
  8921=>"000011001",
  8922=>"011001001",
  8923=>"110001000",
  8924=>"100011110",
  8925=>"001000001",
  8926=>"101001110",
  8927=>"111111001",
  8928=>"010100011",
  8929=>"101010010",
  8930=>"101011111",
  8931=>"111100111",
  8932=>"001111001",
  8933=>"101001011",
  8934=>"101111011",
  8935=>"111011000",
  8936=>"000000111",
  8937=>"111011100",
  8938=>"000011001",
  8939=>"011001111",
  8940=>"000000110",
  8941=>"111011111",
  8942=>"101000010",
  8943=>"001111010",
  8944=>"110100011",
  8945=>"111111101",
  8946=>"101100010",
  8947=>"001110111",
  8948=>"100100001",
  8949=>"000000110",
  8950=>"000010101",
  8951=>"111011111",
  8952=>"001011010",
  8953=>"011100010",
  8954=>"011101111",
  8955=>"010111010",
  8956=>"000101001",
  8957=>"111010110",
  8958=>"101000100",
  8959=>"000100011",
  8960=>"000111001",
  8961=>"100010111",
  8962=>"110001011",
  8963=>"100000000",
  8964=>"010100010",
  8965=>"010011001",
  8966=>"001111000",
  8967=>"100101000",
  8968=>"100111001",
  8969=>"111100010",
  8970=>"000010111",
  8971=>"101011011",
  8972=>"010110110",
  8973=>"110100111",
  8974=>"001111111",
  8975=>"100100110",
  8976=>"101000011",
  8977=>"110110111",
  8978=>"101011101",
  8979=>"101000100",
  8980=>"000111010",
  8981=>"111011111",
  8982=>"111101101",
  8983=>"101000001",
  8984=>"101001111",
  8985=>"001000111",
  8986=>"000000000",
  8987=>"000001111",
  8988=>"000101001",
  8989=>"100011101",
  8990=>"101110000",
  8991=>"001001011",
  8992=>"001111000",
  8993=>"011100111",
  8994=>"000010001",
  8995=>"110111010",
  8996=>"101100000",
  8997=>"000010110",
  8998=>"011110000",
  8999=>"111001101",
  9000=>"111101011",
  9001=>"111101000",
  9002=>"001000001",
  9003=>"000011111",
  9004=>"011001010",
  9005=>"101011010",
  9006=>"000110010",
  9007=>"110101000",
  9008=>"010000111",
  9009=>"111110010",
  9010=>"000011000",
  9011=>"011000110",
  9012=>"100101111",
  9013=>"101001001",
  9014=>"010110000",
  9015=>"011101111",
  9016=>"101000000",
  9017=>"010100000",
  9018=>"000001100",
  9019=>"001010101",
  9020=>"010111111",
  9021=>"010001001",
  9022=>"100100101",
  9023=>"110011111",
  9024=>"010111101",
  9025=>"001011010",
  9026=>"011010001",
  9027=>"111110110",
  9028=>"110101101",
  9029=>"110011101",
  9030=>"001000110",
  9031=>"010101001",
  9032=>"010011010",
  9033=>"111001001",
  9034=>"101000010",
  9035=>"101011010",
  9036=>"110011101",
  9037=>"000100111",
  9038=>"101011110",
  9039=>"110111011",
  9040=>"101000011",
  9041=>"000001100",
  9042=>"001100001",
  9043=>"000100101",
  9044=>"001110010",
  9045=>"111000101",
  9046=>"001100001",
  9047=>"011010101",
  9048=>"011010111",
  9049=>"101010001",
  9050=>"111011110",
  9051=>"101100000",
  9052=>"011111111",
  9053=>"000101000",
  9054=>"111110010",
  9055=>"000101010",
  9056=>"001011011",
  9057=>"111100111",
  9058=>"101011110",
  9059=>"110110100",
  9060=>"110001111",
  9061=>"100101111",
  9062=>"000010100",
  9063=>"001100110",
  9064=>"000100111",
  9065=>"101111000",
  9066=>"010000110",
  9067=>"110011010",
  9068=>"110110000",
  9069=>"101010000",
  9070=>"111110111",
  9071=>"010110110",
  9072=>"011111000",
  9073=>"101000111",
  9074=>"100100011",
  9075=>"111001101",
  9076=>"000101010",
  9077=>"111101110",
  9078=>"101101000",
  9079=>"000101000",
  9080=>"101000111",
  9081=>"100101101",
  9082=>"111110101",
  9083=>"101000001",
  9084=>"111111111",
  9085=>"111100111",
  9086=>"111110011",
  9087=>"111101100",
  9088=>"000100010",
  9089=>"000000001",
  9090=>"011111011",
  9091=>"111010000",
  9092=>"110001101",
  9093=>"100110010",
  9094=>"101000110",
  9095=>"100010110",
  9096=>"001011100",
  9097=>"100110111",
  9098=>"000011100",
  9099=>"101010111",
  9100=>"001001101",
  9101=>"000100010",
  9102=>"000100100",
  9103=>"110101110",
  9104=>"000000100",
  9105=>"101011101",
  9106=>"000101010",
  9107=>"011000001",
  9108=>"010010010",
  9109=>"001000000",
  9110=>"000001011",
  9111=>"000011011",
  9112=>"111110110",
  9113=>"101011000",
  9114=>"000111101",
  9115=>"110001110",
  9116=>"000000101",
  9117=>"111010100",
  9118=>"101010011",
  9119=>"000111111",
  9120=>"110111000",
  9121=>"101010010",
  9122=>"101011111",
  9123=>"011010010",
  9124=>"000110000",
  9125=>"101100000",
  9126=>"110000100",
  9127=>"000010000",
  9128=>"111100111",
  9129=>"111111111",
  9130=>"011011111",
  9131=>"100001111",
  9132=>"010111111",
  9133=>"101100001",
  9134=>"111001101",
  9135=>"001001100",
  9136=>"011001000",
  9137=>"111110001",
  9138=>"111101101",
  9139=>"010100001",
  9140=>"110100000",
  9141=>"111110011",
  9142=>"011101011",
  9143=>"100011000",
  9144=>"000101010",
  9145=>"100001111",
  9146=>"011011010",
  9147=>"000110100",
  9148=>"110010111",
  9149=>"010011100",
  9150=>"111111000",
  9151=>"001001111",
  9152=>"000110110",
  9153=>"110100010",
  9154=>"110111100",
  9155=>"100010000",
  9156=>"000100000",
  9157=>"111001101",
  9158=>"011110110",
  9159=>"011011011",
  9160=>"000001101",
  9161=>"010101101",
  9162=>"001010100",
  9163=>"100100101",
  9164=>"101011001",
  9165=>"110010111",
  9166=>"011010010",
  9167=>"000001110",
  9168=>"100101111",
  9169=>"000100111",
  9170=>"101000101",
  9171=>"000110001",
  9172=>"000100010",
  9173=>"000000110",
  9174=>"000011111",
  9175=>"101100101",
  9176=>"000010011",
  9177=>"010010101",
  9178=>"010111110",
  9179=>"000000010",
  9180=>"110011101",
  9181=>"101111000",
  9182=>"101110001",
  9183=>"100100000",
  9184=>"111111100",
  9185=>"101001001",
  9186=>"101110011",
  9187=>"110010101",
  9188=>"101011101",
  9189=>"000010000",
  9190=>"001001001",
  9191=>"001011100",
  9192=>"000001111",
  9193=>"000111001",
  9194=>"010000000",
  9195=>"100010101",
  9196=>"010001000",
  9197=>"001011001",
  9198=>"111111001",
  9199=>"011101110",
  9200=>"010101001",
  9201=>"111001011",
  9202=>"101000001",
  9203=>"110110001",
  9204=>"111100000",
  9205=>"010010101",
  9206=>"001001101",
  9207=>"101001111",
  9208=>"000110011",
  9209=>"010010101",
  9210=>"001011110",
  9211=>"001010111",
  9212=>"001000001",
  9213=>"110000110",
  9214=>"001110101",
  9215=>"110101001",
  9216=>"001011110",
  9217=>"101110100",
  9218=>"010010000",
  9219=>"000001100",
  9220=>"111010110",
  9221=>"001000010",
  9222=>"110100001",
  9223=>"100110101",
  9224=>"000000101",
  9225=>"010000000",
  9226=>"000001001",
  9227=>"111001001",
  9228=>"101101101",
  9229=>"111110010",
  9230=>"101011101",
  9231=>"011111100",
  9232=>"011100101",
  9233=>"011110111",
  9234=>"001100001",
  9235=>"011011110",
  9236=>"010000111",
  9237=>"110111110",
  9238=>"111101110",
  9239=>"000001011",
  9240=>"001001101",
  9241=>"000100100",
  9242=>"110000011",
  9243=>"010101100",
  9244=>"010001000",
  9245=>"110000010",
  9246=>"110010110",
  9247=>"100011111",
  9248=>"001011110",
  9249=>"011100110",
  9250=>"010010001",
  9251=>"100110100",
  9252=>"001101110",
  9253=>"010010010",
  9254=>"100001110",
  9255=>"011001011",
  9256=>"100010000",
  9257=>"111110100",
  9258=>"010101010",
  9259=>"110101000",
  9260=>"111110101",
  9261=>"011001011",
  9262=>"000001000",
  9263=>"101001000",
  9264=>"000001100",
  9265=>"010010111",
  9266=>"011100110",
  9267=>"001011111",
  9268=>"000111100",
  9269=>"000100010",
  9270=>"000110000",
  9271=>"010011101",
  9272=>"001100100",
  9273=>"100111010",
  9274=>"110111111",
  9275=>"100110101",
  9276=>"101000010",
  9277=>"111001100",
  9278=>"010001000",
  9279=>"111111100",
  9280=>"111001111",
  9281=>"011110001",
  9282=>"111000000",
  9283=>"011010111",
  9284=>"110110110",
  9285=>"110011111",
  9286=>"001001000",
  9287=>"101110001",
  9288=>"010011111",
  9289=>"110000000",
  9290=>"011111001",
  9291=>"001011000",
  9292=>"001110001",
  9293=>"101000100",
  9294=>"101010010",
  9295=>"100010000",
  9296=>"010001110",
  9297=>"001010001",
  9298=>"001001100",
  9299=>"101010101",
  9300=>"110100010",
  9301=>"010011110",
  9302=>"100101110",
  9303=>"101110111",
  9304=>"000111001",
  9305=>"111101010",
  9306=>"101010111",
  9307=>"011110011",
  9308=>"010110101",
  9309=>"110101100",
  9310=>"111110110",
  9311=>"100100111",
  9312=>"110001000",
  9313=>"001000010",
  9314=>"000111011",
  9315=>"011111011",
  9316=>"100100110",
  9317=>"010101011",
  9318=>"110100001",
  9319=>"000010011",
  9320=>"010001101",
  9321=>"100010010",
  9322=>"111001001",
  9323=>"101001011",
  9324=>"010100000",
  9325=>"111101111",
  9326=>"100110000",
  9327=>"010001001",
  9328=>"100111110",
  9329=>"001011101",
  9330=>"110010001",
  9331=>"101011111",
  9332=>"111111111",
  9333=>"101001101",
  9334=>"101001111",
  9335=>"100000111",
  9336=>"110000110",
  9337=>"001000111",
  9338=>"010010000",
  9339=>"101011111",
  9340=>"011101000",
  9341=>"111001100",
  9342=>"110011000",
  9343=>"100001000",
  9344=>"110000010",
  9345=>"111011111",
  9346=>"110100111",
  9347=>"111010010",
  9348=>"100001101",
  9349=>"010001010",
  9350=>"010111011",
  9351=>"001101011",
  9352=>"101001101",
  9353=>"101111100",
  9354=>"100011111",
  9355=>"111010101",
  9356=>"100101110",
  9357=>"010101101",
  9358=>"000001110",
  9359=>"000001010",
  9360=>"101011101",
  9361=>"101011011",
  9362=>"101000111",
  9363=>"010111110",
  9364=>"001101101",
  9365=>"111001010",
  9366=>"001010011",
  9367=>"011110011",
  9368=>"001100001",
  9369=>"110111011",
  9370=>"110011000",
  9371=>"001100010",
  9372=>"110011101",
  9373=>"011100010",
  9374=>"111000000",
  9375=>"011011010",
  9376=>"111110111",
  9377=>"100100001",
  9378=>"011110000",
  9379=>"001000111",
  9380=>"000110011",
  9381=>"101000100",
  9382=>"000011011",
  9383=>"101001101",
  9384=>"001111010",
  9385=>"110101000",
  9386=>"110010011",
  9387=>"111110001",
  9388=>"101101001",
  9389=>"100010000",
  9390=>"111011000",
  9391=>"010001001",
  9392=>"001100111",
  9393=>"110100111",
  9394=>"010001101",
  9395=>"010011111",
  9396=>"101110011",
  9397=>"111001011",
  9398=>"100101110",
  9399=>"001000100",
  9400=>"111001101",
  9401=>"010111101",
  9402=>"000011101",
  9403=>"000011010",
  9404=>"100100000",
  9405=>"101100100",
  9406=>"000001100",
  9407=>"100100010",
  9408=>"111101000",
  9409=>"000010100",
  9410=>"111010101",
  9411=>"100010111",
  9412=>"001001010",
  9413=>"111111000",
  9414=>"010101101",
  9415=>"110110001",
  9416=>"011111000",
  9417=>"100111000",
  9418=>"110000100",
  9419=>"110111010",
  9420=>"111010111",
  9421=>"111111000",
  9422=>"111010000",
  9423=>"011111001",
  9424=>"011011110",
  9425=>"000101000",
  9426=>"111011011",
  9427=>"111000001",
  9428=>"111100100",
  9429=>"111010110",
  9430=>"010010100",
  9431=>"010100010",
  9432=>"011101100",
  9433=>"101110010",
  9434=>"111011100",
  9435=>"111001111",
  9436=>"000010010",
  9437=>"100100010",
  9438=>"010001011",
  9439=>"110101111",
  9440=>"010100011",
  9441=>"011001011",
  9442=>"111110110",
  9443=>"110101011",
  9444=>"000011010",
  9445=>"011011101",
  9446=>"000111111",
  9447=>"111000011",
  9448=>"011000111",
  9449=>"001110101",
  9450=>"100110010",
  9451=>"000101001",
  9452=>"010000011",
  9453=>"010010101",
  9454=>"101111111",
  9455=>"010000000",
  9456=>"110101100",
  9457=>"111111111",
  9458=>"001001110",
  9459=>"111100111",
  9460=>"111001100",
  9461=>"010101100",
  9462=>"000001000",
  9463=>"100011100",
  9464=>"010100010",
  9465=>"111011011",
  9466=>"011000100",
  9467=>"000011100",
  9468=>"101000100",
  9469=>"111011010",
  9470=>"010001110",
  9471=>"100100101",
  9472=>"111001011",
  9473=>"110000100",
  9474=>"101110000",
  9475=>"100011001",
  9476=>"001100110",
  9477=>"111000011",
  9478=>"101010001",
  9479=>"111111000",
  9480=>"101100100",
  9481=>"010011110",
  9482=>"000101010",
  9483=>"101011111",
  9484=>"010111110",
  9485=>"011111110",
  9486=>"110010010",
  9487=>"111110100",
  9488=>"000111100",
  9489=>"000000000",
  9490=>"111111101",
  9491=>"000111000",
  9492=>"110000110",
  9493=>"101100101",
  9494=>"110010111",
  9495=>"010010011",
  9496=>"000000001",
  9497=>"011010010",
  9498=>"110101000",
  9499=>"010001111",
  9500=>"010110111",
  9501=>"100000001",
  9502=>"100001110",
  9503=>"000011010",
  9504=>"010000011",
  9505=>"111011000",
  9506=>"011001111",
  9507=>"110000000",
  9508=>"111001111",
  9509=>"111111101",
  9510=>"000000000",
  9511=>"110000111",
  9512=>"100001011",
  9513=>"101110010",
  9514=>"001010111",
  9515=>"110011100",
  9516=>"001001110",
  9517=>"000101010",
  9518=>"100110111",
  9519=>"101101110",
  9520=>"110010000",
  9521=>"101010110",
  9522=>"101001101",
  9523=>"110001010",
  9524=>"101101111",
  9525=>"110111111",
  9526=>"111001010",
  9527=>"011111011",
  9528=>"000100111",
  9529=>"011100111",
  9530=>"100010011",
  9531=>"001001101",
  9532=>"101101011",
  9533=>"001010101",
  9534=>"010011100",
  9535=>"010010101",
  9536=>"010001100",
  9537=>"101110010",
  9538=>"100111111",
  9539=>"001011011",
  9540=>"100000011",
  9541=>"101111010",
  9542=>"001010011",
  9543=>"001001000",
  9544=>"110100000",
  9545=>"010111001",
  9546=>"111001101",
  9547=>"110011001",
  9548=>"100101001",
  9549=>"001101010",
  9550=>"000000001",
  9551=>"010100001",
  9552=>"111010010",
  9553=>"011000100",
  9554=>"110100101",
  9555=>"001100111",
  9556=>"101000011",
  9557=>"110110001",
  9558=>"101010000",
  9559=>"001001100",
  9560=>"010110010",
  9561=>"001110111",
  9562=>"111000100",
  9563=>"100000000",
  9564=>"111011110",
  9565=>"100000111",
  9566=>"011011100",
  9567=>"111010111",
  9568=>"111001011",
  9569=>"000100111",
  9570=>"000111111",
  9571=>"001100001",
  9572=>"110100001",
  9573=>"011100011",
  9574=>"100111001",
  9575=>"000101001",
  9576=>"001000001",
  9577=>"101001111",
  9578=>"001000000",
  9579=>"100011001",
  9580=>"100111011",
  9581=>"001101111",
  9582=>"100001110",
  9583=>"001000111",
  9584=>"100101100",
  9585=>"111011110",
  9586=>"011111100",
  9587=>"111111110",
  9588=>"000110000",
  9589=>"010001010",
  9590=>"010001100",
  9591=>"011101101",
  9592=>"000011010",
  9593=>"101001000",
  9594=>"110010001",
  9595=>"001000011",
  9596=>"001001001",
  9597=>"110110011",
  9598=>"100000001",
  9599=>"010010011",
  9600=>"010011010",
  9601=>"011000011",
  9602=>"111001010",
  9603=>"110010011",
  9604=>"101111111",
  9605=>"110001011",
  9606=>"010000110",
  9607=>"000110011",
  9608=>"110111100",
  9609=>"111010101",
  9610=>"100001001",
  9611=>"101111111",
  9612=>"001011010",
  9613=>"101100111",
  9614=>"000100000",
  9615=>"111010101",
  9616=>"000000011",
  9617=>"101100011",
  9618=>"100111100",
  9619=>"110101011",
  9620=>"111111100",
  9621=>"100010010",
  9622=>"010010110",
  9623=>"011011100",
  9624=>"111100011",
  9625=>"001100001",
  9626=>"000000001",
  9627=>"101011110",
  9628=>"011100110",
  9629=>"101101010",
  9630=>"111011010",
  9631=>"111001111",
  9632=>"010010000",
  9633=>"111001110",
  9634=>"011110111",
  9635=>"010011000",
  9636=>"100011001",
  9637=>"111000100",
  9638=>"110001111",
  9639=>"111010010",
  9640=>"010011110",
  9641=>"100000011",
  9642=>"010101111",
  9643=>"111111110",
  9644=>"100001000",
  9645=>"101010111",
  9646=>"001001100",
  9647=>"001110000",
  9648=>"011000011",
  9649=>"000111111",
  9650=>"010100100",
  9651=>"100001110",
  9652=>"011100001",
  9653=>"111100100",
  9654=>"111110001",
  9655=>"100000010",
  9656=>"000110010",
  9657=>"000100100",
  9658=>"100010101",
  9659=>"100001010",
  9660=>"000110111",
  9661=>"101001011",
  9662=>"101001000",
  9663=>"110000111",
  9664=>"100001110",
  9665=>"111010011",
  9666=>"001001000",
  9667=>"100001010",
  9668=>"010000111",
  9669=>"100000000",
  9670=>"111011111",
  9671=>"000101000",
  9672=>"011111000",
  9673=>"111011011",
  9674=>"101010010",
  9675=>"010110010",
  9676=>"111111010",
  9677=>"111100110",
  9678=>"111001011",
  9679=>"101010100",
  9680=>"010011010",
  9681=>"011101001",
  9682=>"011000101",
  9683=>"001010000",
  9684=>"101110001",
  9685=>"001001110",
  9686=>"000101000",
  9687=>"100100110",
  9688=>"001111111",
  9689=>"011111010",
  9690=>"100011111",
  9691=>"111110001",
  9692=>"001011101",
  9693=>"001101011",
  9694=>"100100100",
  9695=>"111111001",
  9696=>"011100110",
  9697=>"111011100",
  9698=>"110111101",
  9699=>"111010100",
  9700=>"100010111",
  9701=>"000001001",
  9702=>"111001010",
  9703=>"100010110",
  9704=>"101000011",
  9705=>"011011101",
  9706=>"011010101",
  9707=>"110111100",
  9708=>"111000000",
  9709=>"101100010",
  9710=>"100000101",
  9711=>"011010000",
  9712=>"111101001",
  9713=>"111111110",
  9714=>"110101111",
  9715=>"111000101",
  9716=>"100000010",
  9717=>"010010010",
  9718=>"111010001",
  9719=>"101110010",
  9720=>"010110111",
  9721=>"011010100",
  9722=>"000001001",
  9723=>"000101010",
  9724=>"011011100",
  9725=>"100000111",
  9726=>"111000111",
  9727=>"010100101",
  9728=>"011111110",
  9729=>"101011001",
  9730=>"110000110",
  9731=>"011110001",
  9732=>"110011001",
  9733=>"111101011",
  9734=>"101100010",
  9735=>"110110101",
  9736=>"100001111",
  9737=>"101110111",
  9738=>"000011001",
  9739=>"001010011",
  9740=>"010110000",
  9741=>"111010001",
  9742=>"000001011",
  9743=>"010100011",
  9744=>"100110101",
  9745=>"111110011",
  9746=>"111001101",
  9747=>"001001011",
  9748=>"010000010",
  9749=>"000011100",
  9750=>"000101011",
  9751=>"011010011",
  9752=>"010101100",
  9753=>"001101010",
  9754=>"101000000",
  9755=>"100010110",
  9756=>"001111111",
  9757=>"011100010",
  9758=>"101110110",
  9759=>"110010100",
  9760=>"011000011",
  9761=>"000110100",
  9762=>"001101110",
  9763=>"101111101",
  9764=>"101101100",
  9765=>"011000011",
  9766=>"100000000",
  9767=>"110011000",
  9768=>"100100110",
  9769=>"000100101",
  9770=>"001001110",
  9771=>"010100011",
  9772=>"001101110",
  9773=>"000011100",
  9774=>"011001110",
  9775=>"010101001",
  9776=>"001000100",
  9777=>"100010000",
  9778=>"100010011",
  9779=>"111101100",
  9780=>"011000011",
  9781=>"001111110",
  9782=>"001101101",
  9783=>"011111000",
  9784=>"101010111",
  9785=>"000111101",
  9786=>"000001101",
  9787=>"111100001",
  9788=>"000010000",
  9789=>"000110100",
  9790=>"110001000",
  9791=>"000110110",
  9792=>"001000101",
  9793=>"001011101",
  9794=>"001100000",
  9795=>"111000100",
  9796=>"000101111",
  9797=>"001010001",
  9798=>"001011011",
  9799=>"010110011",
  9800=>"110011000",
  9801=>"101011101",
  9802=>"000010000",
  9803=>"100111001",
  9804=>"101111011",
  9805=>"010111011",
  9806=>"001101111",
  9807=>"101110110",
  9808=>"110000001",
  9809=>"000110010",
  9810=>"011001000",
  9811=>"101100111",
  9812=>"111001011",
  9813=>"000100000",
  9814=>"011110010",
  9815=>"100010110",
  9816=>"101110010",
  9817=>"010111100",
  9818=>"100000000",
  9819=>"101111110",
  9820=>"101010010",
  9821=>"001000010",
  9822=>"111111101",
  9823=>"101011100",
  9824=>"011110000",
  9825=>"011101000",
  9826=>"000111010",
  9827=>"111000010",
  9828=>"001111110",
  9829=>"101101001",
  9830=>"100100110",
  9831=>"010010010",
  9832=>"100010111",
  9833=>"011000101",
  9834=>"110000010",
  9835=>"011110111",
  9836=>"000110011",
  9837=>"101001101",
  9838=>"110010101",
  9839=>"000000000",
  9840=>"100000101",
  9841=>"000001001",
  9842=>"010001000",
  9843=>"100001001",
  9844=>"100100000",
  9845=>"010101001",
  9846=>"111110110",
  9847=>"110010001",
  9848=>"100010110",
  9849=>"111110111",
  9850=>"001110000",
  9851=>"110111100",
  9852=>"110001100",
  9853=>"111100101",
  9854=>"100001011",
  9855=>"101001001",
  9856=>"010111110",
  9857=>"000101001",
  9858=>"010111000",
  9859=>"101111010",
  9860=>"010011111",
  9861=>"110011101",
  9862=>"111110010",
  9863=>"111111000",
  9864=>"100001111",
  9865=>"010000101",
  9866=>"011010010",
  9867=>"011101111",
  9868=>"000010111",
  9869=>"010000000",
  9870=>"110010001",
  9871=>"010101011",
  9872=>"010010000",
  9873=>"101000110",
  9874=>"110110000",
  9875=>"111111100",
  9876=>"011010111",
  9877=>"000001111",
  9878=>"110111101",
  9879=>"111111001",
  9880=>"001101101",
  9881=>"101000000",
  9882=>"000110110",
  9883=>"010000110",
  9884=>"110000111",
  9885=>"000110000",
  9886=>"000010100",
  9887=>"110001001",
  9888=>"010001011",
  9889=>"110111000",
  9890=>"010000110",
  9891=>"101010110",
  9892=>"010000100",
  9893=>"000111101",
  9894=>"100011000",
  9895=>"111000111",
  9896=>"001000101",
  9897=>"101000101",
  9898=>"000000100",
  9899=>"001000001",
  9900=>"010010000",
  9901=>"011110101",
  9902=>"011101010",
  9903=>"101001010",
  9904=>"111110011",
  9905=>"001001010",
  9906=>"000110011",
  9907=>"100011001",
  9908=>"111110010",
  9909=>"000100111",
  9910=>"101000100",
  9911=>"010000010",
  9912=>"111011011",
  9913=>"101000010",
  9914=>"110100011",
  9915=>"011010111",
  9916=>"000010000",
  9917=>"111101010",
  9918=>"011011100",
  9919=>"100110001",
  9920=>"001110011",
  9921=>"010001101",
  9922=>"101011010",
  9923=>"100011001",
  9924=>"110010011",
  9925=>"111001011",
  9926=>"101011101",
  9927=>"000101101",
  9928=>"000000011",
  9929=>"110101011",
  9930=>"101101011",
  9931=>"010110000",
  9932=>"001000101",
  9933=>"110010011",
  9934=>"100101111",
  9935=>"011110000",
  9936=>"010101011",
  9937=>"011101011",
  9938=>"010110110",
  9939=>"100101000",
  9940=>"101110011",
  9941=>"011100011",
  9942=>"010101100",
  9943=>"000101011",
  9944=>"001001001",
  9945=>"101010100",
  9946=>"010001001",
  9947=>"111011000",
  9948=>"101101001",
  9949=>"101000101",
  9950=>"010101000",
  9951=>"110111000",
  9952=>"111011011",
  9953=>"111111111",
  9954=>"100111101",
  9955=>"100100111",
  9956=>"001100111",
  9957=>"000011010",
  9958=>"010101000",
  9959=>"010111110",
  9960=>"111100010",
  9961=>"011001001",
  9962=>"100101101",
  9963=>"011101001",
  9964=>"100101101",
  9965=>"000100000",
  9966=>"011110101",
  9967=>"001110101",
  9968=>"100100100",
  9969=>"000101001",
  9970=>"011000000",
  9971=>"001011011",
  9972=>"111111010",
  9973=>"110000011",
  9974=>"111101111",
  9975=>"001111111",
  9976=>"010111011",
  9977=>"101011111",
  9978=>"100011110",
  9979=>"100011101",
  9980=>"110100100",
  9981=>"001000011",
  9982=>"000000000",
  9983=>"010000000",
  9984=>"001001010",
  9985=>"001000000",
  9986=>"101111111",
  9987=>"110010101",
  9988=>"101111101",
  9989=>"000000011",
  9990=>"111111110",
  9991=>"011001101",
  9992=>"010100111",
  9993=>"010101110",
  9994=>"110011101",
  9995=>"010011011",
  9996=>"100001101",
  9997=>"111110110",
  9998=>"110000101",
  9999=>"010111000",
  10000=>"110100000",
  10001=>"100111001",
  10002=>"001001100",
  10003=>"110110001",
  10004=>"110110110",
  10005=>"111011000",
  10006=>"111000101",
  10007=>"110101101",
  10008=>"010000000",
  10009=>"010011010",
  10010=>"010111101",
  10011=>"111001100",
  10012=>"001000000",
  10013=>"001001100",
  10014=>"010011001",
  10015=>"101000100",
  10016=>"000001111",
  10017=>"111011110",
  10018=>"011111111",
  10019=>"111111101",
  10020=>"111001000",
  10021=>"000111011",
  10022=>"011000110",
  10023=>"010001111",
  10024=>"010111100",
  10025=>"111001101",
  10026=>"010000000",
  10027=>"001001011",
  10028=>"010001000",
  10029=>"111110010",
  10030=>"000100111",
  10031=>"010100100",
  10032=>"111110001",
  10033=>"010011110",
  10034=>"101100001",
  10035=>"000100100",
  10036=>"101010100",
  10037=>"111110101",
  10038=>"110001110",
  10039=>"000111011",
  10040=>"011010000",
  10041=>"000101010",
  10042=>"101110010",
  10043=>"000010001",
  10044=>"001011110",
  10045=>"110111100",
  10046=>"010011101",
  10047=>"101110001",
  10048=>"100001010",
  10049=>"011010101",
  10050=>"111010010",
  10051=>"010111011",
  10052=>"001000010",
  10053=>"010101100",
  10054=>"100101011",
  10055=>"011101110",
  10056=>"110011111",
  10057=>"000101101",
  10058=>"111111111",
  10059=>"011011011",
  10060=>"100111000",
  10061=>"111000000",
  10062=>"101011010",
  10063=>"100000111",
  10064=>"000110010",
  10065=>"000011110",
  10066=>"011111101",
  10067=>"011000101",
  10068=>"111111000",
  10069=>"001011000",
  10070=>"000001010",
  10071=>"000010110",
  10072=>"001001011",
  10073=>"101000000",
  10074=>"010010110",
  10075=>"111100001",
  10076=>"010100001",
  10077=>"110011000",
  10078=>"000011001",
  10079=>"111010011",
  10080=>"100011110",
  10081=>"011000011",
  10082=>"101111111",
  10083=>"101111111",
  10084=>"110010000",
  10085=>"000100111",
  10086=>"000001011",
  10087=>"111001110",
  10088=>"110001101",
  10089=>"111100010",
  10090=>"010111100",
  10091=>"010111000",
  10092=>"110110110",
  10093=>"000101101",
  10094=>"111010010",
  10095=>"010000001",
  10096=>"101010001",
  10097=>"010101011",
  10098=>"111110011",
  10099=>"101100000",
  10100=>"110011100",
  10101=>"010000101",
  10102=>"111001110",
  10103=>"011100110",
  10104=>"010100010",
  10105=>"011010111",
  10106=>"010100010",
  10107=>"011001110",
  10108=>"101011111",
  10109=>"001110011",
  10110=>"011101111",
  10111=>"001001011",
  10112=>"000110010",
  10113=>"111101011",
  10114=>"100111100",
  10115=>"011110001",
  10116=>"001100110",
  10117=>"000010010",
  10118=>"000011110",
  10119=>"110101000",
  10120=>"111101001",
  10121=>"100010011",
  10122=>"000100000",
  10123=>"010100000",
  10124=>"010101000",
  10125=>"110001110",
  10126=>"001101011",
  10127=>"001110000",
  10128=>"011100110",
  10129=>"110011100",
  10130=>"001110101",
  10131=>"011111101",
  10132=>"001110111",
  10133=>"010011010",
  10134=>"101001000",
  10135=>"111011100",
  10136=>"010111001",
  10137=>"110001111",
  10138=>"110101011",
  10139=>"010111111",
  10140=>"111001011",
  10141=>"000010011",
  10142=>"001011100",
  10143=>"011001011",
  10144=>"011100110",
  10145=>"100010011",
  10146=>"001101101",
  10147=>"111111110",
  10148=>"000110101",
  10149=>"101111100",
  10150=>"010100101",
  10151=>"000101111",
  10152=>"001001011",
  10153=>"101011100",
  10154=>"110001101",
  10155=>"001101110",
  10156=>"110011000",
  10157=>"110001111",
  10158=>"110000101",
  10159=>"111100110",
  10160=>"011111000",
  10161=>"010001001",
  10162=>"001011110",
  10163=>"111001011",
  10164=>"111110110",
  10165=>"111001011",
  10166=>"101110000",
  10167=>"000111010",
  10168=>"000100000",
  10169=>"011000100",
  10170=>"110000110",
  10171=>"001010101",
  10172=>"010100000",
  10173=>"011010101",
  10174=>"100110101",
  10175=>"000100110",
  10176=>"101010000",
  10177=>"110011111",
  10178=>"100100111",
  10179=>"011011100",
  10180=>"111111110",
  10181=>"101101110",
  10182=>"011111100",
  10183=>"110010100",
  10184=>"000000011",
  10185=>"101101101",
  10186=>"001101111",
  10187=>"010001000",
  10188=>"100101100",
  10189=>"010000111",
  10190=>"110110100",
  10191=>"111111110",
  10192=>"000100000",
  10193=>"010001111",
  10194=>"110110001",
  10195=>"010001110",
  10196=>"101100010",
  10197=>"000010011",
  10198=>"111101000",
  10199=>"101010111",
  10200=>"010001100",
  10201=>"111111000",
  10202=>"000000100",
  10203=>"101100101",
  10204=>"010111110",
  10205=>"100101001",
  10206=>"100100111",
  10207=>"011111110",
  10208=>"111001101",
  10209=>"101110110",
  10210=>"101010010",
  10211=>"001101001",
  10212=>"101010000",
  10213=>"000011000",
  10214=>"011011000",
  10215=>"100010001",
  10216=>"111101111",
  10217=>"011010001",
  10218=>"000010110",
  10219=>"110110110",
  10220=>"001000111",
  10221=>"010010000",
  10222=>"101101000",
  10223=>"010100011",
  10224=>"000011011",
  10225=>"010111000",
  10226=>"010000111",
  10227=>"111001100",
  10228=>"000011111",
  10229=>"101101011",
  10230=>"011110110",
  10231=>"011110010",
  10232=>"101000000",
  10233=>"000010111",
  10234=>"001110111",
  10235=>"111010100",
  10236=>"011010111",
  10237=>"110101000",
  10238=>"010011100",
  10239=>"101000110",
  10240=>"111111010",
  10241=>"000000100",
  10242=>"100010101",
  10243=>"001001010",
  10244=>"100100011",
  10245=>"000010110",
  10246=>"010011111",
  10247=>"111111101",
  10248=>"011111101",
  10249=>"111000101",
  10250=>"011101100",
  10251=>"001001101",
  10252=>"111010011",
  10253=>"000000000",
  10254=>"111111001",
  10255=>"001101110",
  10256=>"010010101",
  10257=>"100011111",
  10258=>"000100100",
  10259=>"001100011",
  10260=>"111110110",
  10261=>"001001000",
  10262=>"010100110",
  10263=>"010101010",
  10264=>"100100111",
  10265=>"001001011",
  10266=>"110110100",
  10267=>"100111010",
  10268=>"101100000",
  10269=>"100111100",
  10270=>"001101111",
  10271=>"100110011",
  10272=>"001111001",
  10273=>"100001111",
  10274=>"111001001",
  10275=>"000010010",
  10276=>"011101000",
  10277=>"100011011",
  10278=>"010001011",
  10279=>"110101010",
  10280=>"011010001",
  10281=>"001010101",
  10282=>"101010110",
  10283=>"110010100",
  10284=>"110101010",
  10285=>"110101011",
  10286=>"110000001",
  10287=>"000001110",
  10288=>"000111000",
  10289=>"000011100",
  10290=>"101101111",
  10291=>"011101000",
  10292=>"101010100",
  10293=>"000111101",
  10294=>"010110000",
  10295=>"000100101",
  10296=>"111100000",
  10297=>"111001100",
  10298=>"100011110",
  10299=>"100100100",
  10300=>"000010000",
  10301=>"110111001",
  10302=>"111110100",
  10303=>"000001111",
  10304=>"111111000",
  10305=>"100110000",
  10306=>"000001011",
  10307=>"101101000",
  10308=>"001101011",
  10309=>"101100100",
  10310=>"100001011",
  10311=>"101100110",
  10312=>"011010011",
  10313=>"011101000",
  10314=>"101100101",
  10315=>"010100101",
  10316=>"000010011",
  10317=>"010000001",
  10318=>"011111011",
  10319=>"110010101",
  10320=>"000000001",
  10321=>"101111010",
  10322=>"101111010",
  10323=>"010000111",
  10324=>"110011111",
  10325=>"011011010",
  10326=>"110101000",
  10327=>"011001001",
  10328=>"010101111",
  10329=>"001011111",
  10330=>"111100001",
  10331=>"111011011",
  10332=>"011011101",
  10333=>"110001110",
  10334=>"001110001",
  10335=>"000010110",
  10336=>"000000010",
  10337=>"010110001",
  10338=>"010011010",
  10339=>"111100010",
  10340=>"000111100",
  10341=>"111111110",
  10342=>"000010011",
  10343=>"011111000",
  10344=>"101010110",
  10345=>"001001101",
  10346=>"011100011",
  10347=>"110010110",
  10348=>"010000111",
  10349=>"110110100",
  10350=>"000000001",
  10351=>"111101101",
  10352=>"100001100",
  10353=>"110000000",
  10354=>"011101011",
  10355=>"001110111",
  10356=>"100110111",
  10357=>"101000101",
  10358=>"110010000",
  10359=>"101101011",
  10360=>"110010101",
  10361=>"101010110",
  10362=>"011011100",
  10363=>"010100110",
  10364=>"000111111",
  10365=>"011011010",
  10366=>"000011100",
  10367=>"000011000",
  10368=>"000101000",
  10369=>"000101100",
  10370=>"111101101",
  10371=>"111110111",
  10372=>"011101011",
  10373=>"100011111",
  10374=>"110000010",
  10375=>"010001110",
  10376=>"010001011",
  10377=>"011100011",
  10378=>"010100001",
  10379=>"101000111",
  10380=>"111010111",
  10381=>"010100000",
  10382=>"101001000",
  10383=>"111100011",
  10384=>"110001010",
  10385=>"000110101",
  10386=>"001011010",
  10387=>"001111011",
  10388=>"100111110",
  10389=>"000000110",
  10390=>"000010001",
  10391=>"100001110",
  10392=>"010000000",
  10393=>"100010101",
  10394=>"000001101",
  10395=>"111101101",
  10396=>"010010101",
  10397=>"011000010",
  10398=>"101011011",
  10399=>"111011000",
  10400=>"110110111",
  10401=>"100011000",
  10402=>"110101011",
  10403=>"000110010",
  10404=>"100100010",
  10405=>"111010010",
  10406=>"000110000",
  10407=>"101010011",
  10408=>"110111111",
  10409=>"100011000",
  10410=>"010001000",
  10411=>"110010001",
  10412=>"011110011",
  10413=>"000011101",
  10414=>"011111110",
  10415=>"001001100",
  10416=>"000000000",
  10417=>"000000001",
  10418=>"001101000",
  10419=>"000101010",
  10420=>"101110111",
  10421=>"101100000",
  10422=>"011111100",
  10423=>"101110110",
  10424=>"110111001",
  10425=>"011100001",
  10426=>"101010011",
  10427=>"000010100",
  10428=>"010000111",
  10429=>"011110111",
  10430=>"111111001",
  10431=>"110101001",
  10432=>"101000001",
  10433=>"000000011",
  10434=>"000110100",
  10435=>"100010101",
  10436=>"000000111",
  10437=>"000000001",
  10438=>"000111001",
  10439=>"000001001",
  10440=>"011111011",
  10441=>"110100111",
  10442=>"010100111",
  10443=>"010000101",
  10444=>"001010000",
  10445=>"100101100",
  10446=>"001110000",
  10447=>"001001010",
  10448=>"101101100",
  10449=>"010111011",
  10450=>"101010000",
  10451=>"001111111",
  10452=>"001010010",
  10453=>"001010101",
  10454=>"011000000",
  10455=>"001110010",
  10456=>"101110110",
  10457=>"110100100",
  10458=>"010011011",
  10459=>"001010011",
  10460=>"001001101",
  10461=>"110011101",
  10462=>"000011101",
  10463=>"110101100",
  10464=>"001010110",
  10465=>"001010111",
  10466=>"010111101",
  10467=>"101101000",
  10468=>"101111011",
  10469=>"001011100",
  10470=>"001110010",
  10471=>"111011100",
  10472=>"110001010",
  10473=>"111001101",
  10474=>"000010001",
  10475=>"110001000",
  10476=>"000011110",
  10477=>"110110100",
  10478=>"100000110",
  10479=>"100000001",
  10480=>"111100101",
  10481=>"010010100",
  10482=>"000000100",
  10483=>"001001101",
  10484=>"100110110",
  10485=>"110001100",
  10486=>"000101001",
  10487=>"100010101",
  10488=>"101110011",
  10489=>"100100111",
  10490=>"110010101",
  10491=>"100010000",
  10492=>"101011100",
  10493=>"001011000",
  10494=>"111001110",
  10495=>"000111000",
  10496=>"011011001",
  10497=>"000010000",
  10498=>"100000110",
  10499=>"000111010",
  10500=>"000100011",
  10501=>"011110010",
  10502=>"111101100",
  10503=>"110010011",
  10504=>"000010110",
  10505=>"110000110",
  10506=>"010001001",
  10507=>"111100101",
  10508=>"101001101",
  10509=>"101011001",
  10510=>"011000111",
  10511=>"111110000",
  10512=>"111011011",
  10513=>"101110001",
  10514=>"010010010",
  10515=>"000010101",
  10516=>"111011100",
  10517=>"010000010",
  10518=>"111110001",
  10519=>"010011010",
  10520=>"011100001",
  10521=>"010001011",
  10522=>"101001110",
  10523=>"110000000",
  10524=>"100011011",
  10525=>"101010100",
  10526=>"111001001",
  10527=>"110100001",
  10528=>"011101101",
  10529=>"011010111",
  10530=>"000011001",
  10531=>"111010011",
  10532=>"111101000",
  10533=>"111001001",
  10534=>"101111111",
  10535=>"101111010",
  10536=>"110100010",
  10537=>"010011001",
  10538=>"111010001",
  10539=>"000000011",
  10540=>"000110111",
  10541=>"100010000",
  10542=>"001100010",
  10543=>"000111101",
  10544=>"100110000",
  10545=>"011101100",
  10546=>"010110101",
  10547=>"001100001",
  10548=>"100101000",
  10549=>"000001010",
  10550=>"111011101",
  10551=>"101110000",
  10552=>"001000001",
  10553=>"110001000",
  10554=>"101100100",
  10555=>"101000000",
  10556=>"010110010",
  10557=>"101001111",
  10558=>"010000001",
  10559=>"000011111",
  10560=>"111001110",
  10561=>"100111111",
  10562=>"000111111",
  10563=>"110101010",
  10564=>"011010100",
  10565=>"000100011",
  10566=>"010111110",
  10567=>"011111100",
  10568=>"010010011",
  10569=>"010010000",
  10570=>"001010010",
  10571=>"100100001",
  10572=>"111101101",
  10573=>"001000000",
  10574=>"011101000",
  10575=>"011100010",
  10576=>"110011000",
  10577=>"000111010",
  10578=>"010000111",
  10579=>"000001101",
  10580=>"101010010",
  10581=>"010011001",
  10582=>"011000000",
  10583=>"011100110",
  10584=>"001100011",
  10585=>"110010000",
  10586=>"001110001",
  10587=>"101101011",
  10588=>"100100110",
  10589=>"110111110",
  10590=>"111111011",
  10591=>"101111010",
  10592=>"111101001",
  10593=>"110010101",
  10594=>"010010000",
  10595=>"111100101",
  10596=>"001101101",
  10597=>"100111011",
  10598=>"001111110",
  10599=>"001110101",
  10600=>"100000011",
  10601=>"011111101",
  10602=>"000101100",
  10603=>"010101001",
  10604=>"001000100",
  10605=>"111111110",
  10606=>"000101000",
  10607=>"100001110",
  10608=>"001001010",
  10609=>"100111101",
  10610=>"101101010",
  10611=>"011101111",
  10612=>"010111101",
  10613=>"010111000",
  10614=>"111110100",
  10615=>"100101000",
  10616=>"110100011",
  10617=>"010000010",
  10618=>"101001101",
  10619=>"000000010",
  10620=>"000101001",
  10621=>"010111010",
  10622=>"100100101",
  10623=>"110011010",
  10624=>"001101010",
  10625=>"011011100",
  10626=>"100100111",
  10627=>"011011010",
  10628=>"011001101",
  10629=>"101110001",
  10630=>"001001111",
  10631=>"000010011",
  10632=>"011001001",
  10633=>"100110001",
  10634=>"011100011",
  10635=>"010010110",
  10636=>"101100011",
  10637=>"001001001",
  10638=>"110001101",
  10639=>"100000111",
  10640=>"100110111",
  10641=>"101010001",
  10642=>"101111010",
  10643=>"011110001",
  10644=>"100010100",
  10645=>"001011000",
  10646=>"100110111",
  10647=>"000010111",
  10648=>"001001010",
  10649=>"111010110",
  10650=>"110111100",
  10651=>"101100111",
  10652=>"010100110",
  10653=>"010101001",
  10654=>"110110010",
  10655=>"100011010",
  10656=>"100111110",
  10657=>"100110110",
  10658=>"001101000",
  10659=>"011100100",
  10660=>"001101011",
  10661=>"001000000",
  10662=>"111000111",
  10663=>"000011111",
  10664=>"100111111",
  10665=>"111000110",
  10666=>"001000010",
  10667=>"001100001",
  10668=>"010111000",
  10669=>"000101110",
  10670=>"000000011",
  10671=>"000001101",
  10672=>"101011011",
  10673=>"011111111",
  10674=>"011000000",
  10675=>"010011011",
  10676=>"101100010",
  10677=>"111111011",
  10678=>"001101010",
  10679=>"100110111",
  10680=>"101010000",
  10681=>"110010011",
  10682=>"110000100",
  10683=>"111111010",
  10684=>"010001110",
  10685=>"011010101",
  10686=>"110101100",
  10687=>"000110111",
  10688=>"111101010",
  10689=>"101001100",
  10690=>"010100110",
  10691=>"011101010",
  10692=>"111000010",
  10693=>"100110101",
  10694=>"010011010",
  10695=>"100010101",
  10696=>"000001010",
  10697=>"010100010",
  10698=>"011001101",
  10699=>"111111011",
  10700=>"100110110",
  10701=>"011010100",
  10702=>"100001010",
  10703=>"010110011",
  10704=>"001000100",
  10705=>"100011011",
  10706=>"000011001",
  10707=>"001000110",
  10708=>"010000100",
  10709=>"111110000",
  10710=>"011110101",
  10711=>"111001000",
  10712=>"101100100",
  10713=>"100011101",
  10714=>"011101101",
  10715=>"110100011",
  10716=>"110101100",
  10717=>"110010110",
  10718=>"001011001",
  10719=>"111010000",
  10720=>"000100000",
  10721=>"001110011",
  10722=>"100010010",
  10723=>"001010010",
  10724=>"010101110",
  10725=>"100010000",
  10726=>"101100011",
  10727=>"000110001",
  10728=>"111101100",
  10729=>"010111001",
  10730=>"010100000",
  10731=>"111000100",
  10732=>"011000101",
  10733=>"111011000",
  10734=>"011010111",
  10735=>"101001101",
  10736=>"010101111",
  10737=>"000010110",
  10738=>"100000011",
  10739=>"111111110",
  10740=>"001011001",
  10741=>"010110000",
  10742=>"010001000",
  10743=>"010001000",
  10744=>"011101001",
  10745=>"001011010",
  10746=>"000010000",
  10747=>"111110111",
  10748=>"011100110",
  10749=>"101110111",
  10750=>"110111000",
  10751=>"111001000",
  10752=>"001001000",
  10753=>"011101101",
  10754=>"111001100",
  10755=>"100010101",
  10756=>"111001010",
  10757=>"111000111",
  10758=>"000011010",
  10759=>"111110010",
  10760=>"010001111",
  10761=>"101100000",
  10762=>"111001110",
  10763=>"101000011",
  10764=>"101111110",
  10765=>"111110111",
  10766=>"111111110",
  10767=>"101101001",
  10768=>"010000101",
  10769=>"001100001",
  10770=>"111110110",
  10771=>"000001111",
  10772=>"101101000",
  10773=>"101110010",
  10774=>"101101010",
  10775=>"011010001",
  10776=>"110010100",
  10777=>"010000001",
  10778=>"101001110",
  10779=>"001011001",
  10780=>"110011001",
  10781=>"000101101",
  10782=>"101101111",
  10783=>"111001011",
  10784=>"001010110",
  10785=>"101111110",
  10786=>"011111111",
  10787=>"000100111",
  10788=>"111100110",
  10789=>"010101010",
  10790=>"110000011",
  10791=>"010000110",
  10792=>"010011000",
  10793=>"000111001",
  10794=>"101110111",
  10795=>"011011010",
  10796=>"001100101",
  10797=>"001110001",
  10798=>"101101110",
  10799=>"010101011",
  10800=>"000011001",
  10801=>"011011101",
  10802=>"010100101",
  10803=>"011001111",
  10804=>"011111010",
  10805=>"010010011",
  10806=>"101110010",
  10807=>"001100000",
  10808=>"000011111",
  10809=>"010111100",
  10810=>"110011000",
  10811=>"110011000",
  10812=>"101011000",
  10813=>"111010011",
  10814=>"101010010",
  10815=>"110011100",
  10816=>"110100111",
  10817=>"111011010",
  10818=>"100110010",
  10819=>"110101011",
  10820=>"011001111",
  10821=>"011111011",
  10822=>"111010111",
  10823=>"011000100",
  10824=>"100110101",
  10825=>"000010101",
  10826=>"011111011",
  10827=>"100100011",
  10828=>"000100110",
  10829=>"010100100",
  10830=>"010000000",
  10831=>"100100010",
  10832=>"111011111",
  10833=>"111110111",
  10834=>"001101100",
  10835=>"000011011",
  10836=>"101000100",
  10837=>"000100001",
  10838=>"000011000",
  10839=>"000011101",
  10840=>"000100101",
  10841=>"000110010",
  10842=>"100000000",
  10843=>"000010101",
  10844=>"111010101",
  10845=>"001001010",
  10846=>"101100001",
  10847=>"110110100",
  10848=>"001100111",
  10849=>"001011010",
  10850=>"011001011",
  10851=>"101110011",
  10852=>"100110000",
  10853=>"001101110",
  10854=>"101010011",
  10855=>"111111100",
  10856=>"011001110",
  10857=>"001000101",
  10858=>"010110011",
  10859=>"010110100",
  10860=>"011110110",
  10861=>"011110011",
  10862=>"100110101",
  10863=>"100011111",
  10864=>"001000100",
  10865=>"110111001",
  10866=>"001001000",
  10867=>"110111101",
  10868=>"000010101",
  10869=>"011110110",
  10870=>"000100110",
  10871=>"001001010",
  10872=>"101010000",
  10873=>"110101111",
  10874=>"110111011",
  10875=>"101001001",
  10876=>"011101111",
  10877=>"011000100",
  10878=>"110111111",
  10879=>"110001010",
  10880=>"111100001",
  10881=>"100011100",
  10882=>"001000001",
  10883=>"001000111",
  10884=>"011101111",
  10885=>"000100100",
  10886=>"010010010",
  10887=>"110101010",
  10888=>"011000001",
  10889=>"101110010",
  10890=>"100101101",
  10891=>"001110001",
  10892=>"100010101",
  10893=>"000101110",
  10894=>"100101111",
  10895=>"011001011",
  10896=>"101011111",
  10897=>"100101010",
  10898=>"001110111",
  10899=>"110010110",
  10900=>"011000001",
  10901=>"011010011",
  10902=>"000010001",
  10903=>"111110010",
  10904=>"000101001",
  10905=>"010000001",
  10906=>"111101011",
  10907=>"001101000",
  10908=>"000110010",
  10909=>"001000111",
  10910=>"110111010",
  10911=>"011011111",
  10912=>"101010000",
  10913=>"111011001",
  10914=>"001111010",
  10915=>"101100110",
  10916=>"110100101",
  10917=>"001010100",
  10918=>"001000100",
  10919=>"001000101",
  10920=>"111100010",
  10921=>"111001111",
  10922=>"101000110",
  10923=>"000000111",
  10924=>"001001100",
  10925=>"111010000",
  10926=>"100001010",
  10927=>"100001111",
  10928=>"111101101",
  10929=>"111011100",
  10930=>"110100111",
  10931=>"001010110",
  10932=>"111011011",
  10933=>"110000001",
  10934=>"110101100",
  10935=>"100011101",
  10936=>"001000011",
  10937=>"101001111",
  10938=>"100010011",
  10939=>"010100001",
  10940=>"100010000",
  10941=>"110011010",
  10942=>"110101101",
  10943=>"010100110",
  10944=>"111000011",
  10945=>"100010011",
  10946=>"001001011",
  10947=>"000000011",
  10948=>"000011011",
  10949=>"100001001",
  10950=>"101110011",
  10951=>"111111010",
  10952=>"100111011",
  10953=>"100111000",
  10954=>"000000000",
  10955=>"000001000",
  10956=>"101100111",
  10957=>"010001111",
  10958=>"111111110",
  10959=>"111111000",
  10960=>"011001000",
  10961=>"000001011",
  10962=>"011100011",
  10963=>"011011011",
  10964=>"100001001",
  10965=>"110001011",
  10966=>"100000011",
  10967=>"111111010",
  10968=>"111000101",
  10969=>"111101010",
  10970=>"111111010",
  10971=>"111011101",
  10972=>"110110001",
  10973=>"000000011",
  10974=>"010011001",
  10975=>"101111000",
  10976=>"001010101",
  10977=>"111011101",
  10978=>"101011100",
  10979=>"111000010",
  10980=>"101110000",
  10981=>"000111010",
  10982=>"011101011",
  10983=>"100011111",
  10984=>"101101011",
  10985=>"000000011",
  10986=>"111001111",
  10987=>"000110110",
  10988=>"111010110",
  10989=>"110101010",
  10990=>"001111100",
  10991=>"110000001",
  10992=>"000100111",
  10993=>"100101010",
  10994=>"011011100",
  10995=>"000011101",
  10996=>"010111000",
  10997=>"010111001",
  10998=>"000000010",
  10999=>"000010001",
  11000=>"110111001",
  11001=>"011110011",
  11002=>"100111011",
  11003=>"001011000",
  11004=>"001111110",
  11005=>"100111011",
  11006=>"010101100",
  11007=>"010110100",
  11008=>"001100011",
  11009=>"110000010",
  11010=>"100111100",
  11011=>"001101101",
  11012=>"101101011",
  11013=>"001000101",
  11014=>"000010101",
  11015=>"110111011",
  11016=>"111001011",
  11017=>"000010001",
  11018=>"100110000",
  11019=>"011000111",
  11020=>"110101101",
  11021=>"011011000",
  11022=>"001101000",
  11023=>"101101110",
  11024=>"010111010",
  11025=>"001110000",
  11026=>"011010011",
  11027=>"000001001",
  11028=>"010011001",
  11029=>"110110101",
  11030=>"000101000",
  11031=>"000000000",
  11032=>"000110110",
  11033=>"010000011",
  11034=>"000001110",
  11035=>"001001110",
  11036=>"010011111",
  11037=>"001001011",
  11038=>"111001110",
  11039=>"101001011",
  11040=>"011011011",
  11041=>"000110100",
  11042=>"011100011",
  11043=>"010100001",
  11044=>"001001001",
  11045=>"011101000",
  11046=>"101011100",
  11047=>"110111011",
  11048=>"010011101",
  11049=>"101011000",
  11050=>"011011000",
  11051=>"011001000",
  11052=>"100100000",
  11053=>"000100001",
  11054=>"010001000",
  11055=>"000101011",
  11056=>"100111110",
  11057=>"111101101",
  11058=>"101101101",
  11059=>"101000011",
  11060=>"100110000",
  11061=>"101110000",
  11062=>"000011110",
  11063=>"001110011",
  11064=>"010010001",
  11065=>"110110111",
  11066=>"011111111",
  11067=>"110111011",
  11068=>"001010000",
  11069=>"000000100",
  11070=>"011111111",
  11071=>"111100100",
  11072=>"000011110",
  11073=>"101101100",
  11074=>"000000010",
  11075=>"100101010",
  11076=>"101001100",
  11077=>"001101010",
  11078=>"001011110",
  11079=>"001100111",
  11080=>"000100000",
  11081=>"000000110",
  11082=>"110111101",
  11083=>"010100111",
  11084=>"000000111",
  11085=>"011010101",
  11086=>"001100110",
  11087=>"111111100",
  11088=>"010011100",
  11089=>"111111010",
  11090=>"011101000",
  11091=>"011100100",
  11092=>"010111111",
  11093=>"110101110",
  11094=>"010101011",
  11095=>"010000101",
  11096=>"111111111",
  11097=>"010010111",
  11098=>"010011100",
  11099=>"100111000",
  11100=>"100011001",
  11101=>"100111100",
  11102=>"110101001",
  11103=>"111000011",
  11104=>"001110000",
  11105=>"110111011",
  11106=>"011110010",
  11107=>"101010011",
  11108=>"110100001",
  11109=>"000110001",
  11110=>"111000011",
  11111=>"000000010",
  11112=>"001000101",
  11113=>"010100111",
  11114=>"010111111",
  11115=>"101101111",
  11116=>"100101000",
  11117=>"001100000",
  11118=>"110100001",
  11119=>"110111010",
  11120=>"011100001",
  11121=>"111111010",
  11122=>"000000000",
  11123=>"001101011",
  11124=>"110001011",
  11125=>"111000100",
  11126=>"011101011",
  11127=>"001010001",
  11128=>"100101101",
  11129=>"110001001",
  11130=>"110111001",
  11131=>"001000000",
  11132=>"000000001",
  11133=>"011111000",
  11134=>"000100100",
  11135=>"111101101",
  11136=>"000111101",
  11137=>"110011111",
  11138=>"100010110",
  11139=>"100001100",
  11140=>"001010000",
  11141=>"011011011",
  11142=>"010111000",
  11143=>"111000100",
  11144=>"110011111",
  11145=>"101110001",
  11146=>"101001101",
  11147=>"111110100",
  11148=>"110110111",
  11149=>"010110110",
  11150=>"000000100",
  11151=>"000010100",
  11152=>"101100100",
  11153=>"001110011",
  11154=>"111000110",
  11155=>"111011000",
  11156=>"100100100",
  11157=>"001101101",
  11158=>"110110010",
  11159=>"010001100",
  11160=>"110011010",
  11161=>"101110100",
  11162=>"011111101",
  11163=>"000101111",
  11164=>"011100101",
  11165=>"010001011",
  11166=>"101110111",
  11167=>"000110011",
  11168=>"100001010",
  11169=>"111010100",
  11170=>"001110110",
  11171=>"001110101",
  11172=>"111000100",
  11173=>"110110110",
  11174=>"001000001",
  11175=>"000001101",
  11176=>"001001001",
  11177=>"010010001",
  11178=>"001010011",
  11179=>"001000000",
  11180=>"110000000",
  11181=>"000110111",
  11182=>"110011011",
  11183=>"011111101",
  11184=>"000000001",
  11185=>"000010101",
  11186=>"011111111",
  11187=>"001010011",
  11188=>"111000111",
  11189=>"111110000",
  11190=>"001110111",
  11191=>"100011101",
  11192=>"000111111",
  11193=>"110001100",
  11194=>"000001101",
  11195=>"101100001",
  11196=>"101100101",
  11197=>"101111010",
  11198=>"100001010",
  11199=>"011111011",
  11200=>"011000010",
  11201=>"011001010",
  11202=>"111111111",
  11203=>"011101111",
  11204=>"010011110",
  11205=>"111111010",
  11206=>"101111100",
  11207=>"001001011",
  11208=>"000000000",
  11209=>"101001110",
  11210=>"101110000",
  11211=>"010110010",
  11212=>"000000001",
  11213=>"010111001",
  11214=>"010111100",
  11215=>"010111101",
  11216=>"001101110",
  11217=>"110001011",
  11218=>"010000110",
  11219=>"001101010",
  11220=>"001011001",
  11221=>"111011001",
  11222=>"000100001",
  11223=>"110111101",
  11224=>"001011110",
  11225=>"101011000",
  11226=>"100100100",
  11227=>"110011000",
  11228=>"100010011",
  11229=>"000101010",
  11230=>"010101101",
  11231=>"011110101",
  11232=>"011011010",
  11233=>"000010000",
  11234=>"000011101",
  11235=>"000101101",
  11236=>"010011001",
  11237=>"000110111",
  11238=>"110011110",
  11239=>"000110001",
  11240=>"000101000",
  11241=>"110110111",
  11242=>"111110111",
  11243=>"101111110",
  11244=>"010100111",
  11245=>"101110101",
  11246=>"100001000",
  11247=>"110100001",
  11248=>"000111011",
  11249=>"011000010",
  11250=>"110010111",
  11251=>"011101111",
  11252=>"101110111",
  11253=>"100000001",
  11254=>"010110010",
  11255=>"111001101",
  11256=>"010111111",
  11257=>"010001101",
  11258=>"011110000",
  11259=>"000100011",
  11260=>"110010010",
  11261=>"010000110",
  11262=>"000101001",
  11263=>"011011110",
  11264=>"000010110",
  11265=>"000011110",
  11266=>"010000011",
  11267=>"000011100",
  11268=>"101101011",
  11269=>"011001111",
  11270=>"010101001",
  11271=>"111011111",
  11272=>"110100010",
  11273=>"111010101",
  11274=>"011001100",
  11275=>"101110011",
  11276=>"010100101",
  11277=>"011101000",
  11278=>"100101011",
  11279=>"111000100",
  11280=>"111111101",
  11281=>"111101111",
  11282=>"011100001",
  11283=>"101010010",
  11284=>"111110000",
  11285=>"110111001",
  11286=>"011000111",
  11287=>"010001101",
  11288=>"100001010",
  11289=>"111000001",
  11290=>"000000001",
  11291=>"000100001",
  11292=>"110000110",
  11293=>"001110010",
  11294=>"001000101",
  11295=>"000101000",
  11296=>"000101100",
  11297=>"101011000",
  11298=>"111010010",
  11299=>"010100001",
  11300=>"101000001",
  11301=>"011001110",
  11302=>"010101110",
  11303=>"111111111",
  11304=>"100001011",
  11305=>"000010000",
  11306=>"010011101",
  11307=>"010000010",
  11308=>"000111010",
  11309=>"010111100",
  11310=>"111011110",
  11311=>"100000001",
  11312=>"101100000",
  11313=>"100010000",
  11314=>"100000000",
  11315=>"000001100",
  11316=>"001000001",
  11317=>"111010100",
  11318=>"011100010",
  11319=>"111111110",
  11320=>"011000011",
  11321=>"011110000",
  11322=>"101000011",
  11323=>"001011011",
  11324=>"001000101",
  11325=>"100011110",
  11326=>"000010011",
  11327=>"111111110",
  11328=>"101101100",
  11329=>"000101101",
  11330=>"011110101",
  11331=>"001000010",
  11332=>"110010100",
  11333=>"101100101",
  11334=>"100111101",
  11335=>"111101110",
  11336=>"100011100",
  11337=>"101101001",
  11338=>"010001110",
  11339=>"010000110",
  11340=>"111101100",
  11341=>"000111001",
  11342=>"011110101",
  11343=>"011010110",
  11344=>"001101101",
  11345=>"011011100",
  11346=>"011010100",
  11347=>"110100011",
  11348=>"000101101",
  11349=>"001001011",
  11350=>"111110011",
  11351=>"010110111",
  11352=>"100010011",
  11353=>"111111100",
  11354=>"001110110",
  11355=>"111000001",
  11356=>"000001110",
  11357=>"000111011",
  11358=>"011110100",
  11359=>"011100010",
  11360=>"001001110",
  11361=>"100011001",
  11362=>"101001111",
  11363=>"000111010",
  11364=>"000110000",
  11365=>"001111011",
  11366=>"111011011",
  11367=>"010110100",
  11368=>"001001100",
  11369=>"001100010",
  11370=>"011111100",
  11371=>"000111010",
  11372=>"100011111",
  11373=>"011111001",
  11374=>"101000000",
  11375=>"011001000",
  11376=>"001100000",
  11377=>"100001000",
  11378=>"011111111",
  11379=>"001100001",
  11380=>"111111001",
  11381=>"000011100",
  11382=>"110000111",
  11383=>"100100011",
  11384=>"110111100",
  11385=>"000110101",
  11386=>"011111011",
  11387=>"011100101",
  11388=>"001111101",
  11389=>"001111111",
  11390=>"101000001",
  11391=>"000011000",
  11392=>"001110110",
  11393=>"111010011",
  11394=>"010111111",
  11395=>"001100000",
  11396=>"010100110",
  11397=>"101010100",
  11398=>"010101111",
  11399=>"001000101",
  11400=>"001011001",
  11401=>"101011011",
  11402=>"101111000",
  11403=>"110000000",
  11404=>"010100100",
  11405=>"000000000",
  11406=>"101111001",
  11407=>"111000001",
  11408=>"101111101",
  11409=>"111100000",
  11410=>"110000001",
  11411=>"111001001",
  11412=>"111101001",
  11413=>"110110101",
  11414=>"010111010",
  11415=>"000100111",
  11416=>"100100011",
  11417=>"110010001",
  11418=>"011010000",
  11419=>"010110010",
  11420=>"001010010",
  11421=>"101101000",
  11422=>"111101001",
  11423=>"101001010",
  11424=>"010110110",
  11425=>"101111111",
  11426=>"011110011",
  11427=>"111011011",
  11428=>"010101100",
  11429=>"111000001",
  11430=>"001100000",
  11431=>"000110111",
  11432=>"001001001",
  11433=>"001000110",
  11434=>"001000101",
  11435=>"100001011",
  11436=>"110101111",
  11437=>"111011000",
  11438=>"010101010",
  11439=>"111101001",
  11440=>"011011111",
  11441=>"001101011",
  11442=>"100100010",
  11443=>"011100001",
  11444=>"011101100",
  11445=>"001111111",
  11446=>"001001111",
  11447=>"000110111",
  11448=>"101100100",
  11449=>"111101100",
  11450=>"110110111",
  11451=>"111111110",
  11452=>"001100100",
  11453=>"011000010",
  11454=>"000000111",
  11455=>"110101100",
  11456=>"110000111",
  11457=>"001100001",
  11458=>"010000001",
  11459=>"011000000",
  11460=>"001110001",
  11461=>"111111010",
  11462=>"000101001",
  11463=>"000110111",
  11464=>"100011010",
  11465=>"010001111",
  11466=>"000011010",
  11467=>"100000010",
  11468=>"101001101",
  11469=>"011011101",
  11470=>"000111100",
  11471=>"001000100",
  11472=>"010000100",
  11473=>"011111101",
  11474=>"001111011",
  11475=>"010100000",
  11476=>"101010100",
  11477=>"101000101",
  11478=>"111111110",
  11479=>"101100000",
  11480=>"101011010",
  11481=>"010001011",
  11482=>"010001001",
  11483=>"010111100",
  11484=>"000001110",
  11485=>"000101000",
  11486=>"101001101",
  11487=>"011111000",
  11488=>"100011000",
  11489=>"001101111",
  11490=>"011100000",
  11491=>"001111001",
  11492=>"111010110",
  11493=>"010111001",
  11494=>"111101001",
  11495=>"110101101",
  11496=>"100001011",
  11497=>"110110110",
  11498=>"101101011",
  11499=>"010110100",
  11500=>"101001011",
  11501=>"000101011",
  11502=>"111110100",
  11503=>"101010010",
  11504=>"000111011",
  11505=>"111110111",
  11506=>"100000111",
  11507=>"111001011",
  11508=>"100110001",
  11509=>"010011010",
  11510=>"011101011",
  11511=>"011000011",
  11512=>"001011011",
  11513=>"000010011",
  11514=>"110101100",
  11515=>"110100001",
  11516=>"010000111",
  11517=>"010110011",
  11518=>"001000000",
  11519=>"111101000",
  11520=>"101001100",
  11521=>"100001111",
  11522=>"000101100",
  11523=>"100111100",
  11524=>"010001101",
  11525=>"001001000",
  11526=>"110011101",
  11527=>"110111001",
  11528=>"110000000",
  11529=>"100000000",
  11530=>"001010000",
  11531=>"110100010",
  11532=>"011100000",
  11533=>"010001101",
  11534=>"010000100",
  11535=>"111011110",
  11536=>"011001101",
  11537=>"100101000",
  11538=>"011110111",
  11539=>"111010101",
  11540=>"010010001",
  11541=>"011111100",
  11542=>"011110110",
  11543=>"111110111",
  11544=>"101100011",
  11545=>"011011010",
  11546=>"001100010",
  11547=>"001000111",
  11548=>"111011101",
  11549=>"011001000",
  11550=>"101000010",
  11551=>"100101011",
  11552=>"100101011",
  11553=>"001010101",
  11554=>"110101010",
  11555=>"001000011",
  11556=>"100100000",
  11557=>"110011000",
  11558=>"010010001",
  11559=>"001101011",
  11560=>"101101101",
  11561=>"101110100",
  11562=>"000111111",
  11563=>"011110101",
  11564=>"000110111",
  11565=>"011110111",
  11566=>"000111010",
  11567=>"101011111",
  11568=>"101110000",
  11569=>"111000011",
  11570=>"000011000",
  11571=>"101100111",
  11572=>"001011010",
  11573=>"000000111",
  11574=>"110111101",
  11575=>"001001010",
  11576=>"001010000",
  11577=>"010010011",
  11578=>"100011101",
  11579=>"011000110",
  11580=>"000010001",
  11581=>"101010101",
  11582=>"100101110",
  11583=>"101101001",
  11584=>"011111111",
  11585=>"100000111",
  11586=>"000011011",
  11587=>"110000111",
  11588=>"011001011",
  11589=>"000111001",
  11590=>"000010001",
  11591=>"100011010",
  11592=>"000001100",
  11593=>"000101111",
  11594=>"110110101",
  11595=>"001100111",
  11596=>"001010110",
  11597=>"011111001",
  11598=>"011000000",
  11599=>"000110001",
  11600=>"010100110",
  11601=>"010110101",
  11602=>"100000110",
  11603=>"110100010",
  11604=>"001111111",
  11605=>"000101000",
  11606=>"111111011",
  11607=>"110000000",
  11608=>"101000000",
  11609=>"100111111",
  11610=>"000100001",
  11611=>"101101110",
  11612=>"110101101",
  11613=>"011110110",
  11614=>"111010010",
  11615=>"000101100",
  11616=>"010010100",
  11617=>"111111101",
  11618=>"000101111",
  11619=>"010101001",
  11620=>"011001101",
  11621=>"011101000",
  11622=>"100101101",
  11623=>"100010000",
  11624=>"011100001",
  11625=>"000001000",
  11626=>"111010000",
  11627=>"111010100",
  11628=>"001011110",
  11629=>"000100111",
  11630=>"110100000",
  11631=>"000011011",
  11632=>"110100011",
  11633=>"000010010",
  11634=>"011010100",
  11635=>"111001100",
  11636=>"100011001",
  11637=>"000100111",
  11638=>"111111110",
  11639=>"010101010",
  11640=>"111000100",
  11641=>"111100000",
  11642=>"010111011",
  11643=>"111011010",
  11644=>"100101100",
  11645=>"011010000",
  11646=>"010001011",
  11647=>"010000110",
  11648=>"101111101",
  11649=>"101001011",
  11650=>"101100111",
  11651=>"101010110",
  11652=>"100011011",
  11653=>"001011010",
  11654=>"111001101",
  11655=>"001011011",
  11656=>"111011011",
  11657=>"010001101",
  11658=>"101001110",
  11659=>"111011001",
  11660=>"101001100",
  11661=>"101111101",
  11662=>"000010000",
  11663=>"101111101",
  11664=>"000010100",
  11665=>"001011101",
  11666=>"101111011",
  11667=>"000000000",
  11668=>"100000000",
  11669=>"110000100",
  11670=>"101111010",
  11671=>"100110001",
  11672=>"100111001",
  11673=>"000111011",
  11674=>"000010111",
  11675=>"101001001",
  11676=>"101110100",
  11677=>"001110101",
  11678=>"111100000",
  11679=>"000100100",
  11680=>"110101101",
  11681=>"100110111",
  11682=>"111111111",
  11683=>"001011110",
  11684=>"111101001",
  11685=>"000101011",
  11686=>"011000010",
  11687=>"111000101",
  11688=>"111010000",
  11689=>"010110010",
  11690=>"011111001",
  11691=>"011010111",
  11692=>"100001000",
  11693=>"010111111",
  11694=>"101101110",
  11695=>"000010001",
  11696=>"000110101",
  11697=>"010011010",
  11698=>"001111101",
  11699=>"001010000",
  11700=>"111011011",
  11701=>"101110111",
  11702=>"011010011",
  11703=>"100001101",
  11704=>"001001000",
  11705=>"101111100",
  11706=>"100100001",
  11707=>"100010111",
  11708=>"100110111",
  11709=>"011010111",
  11710=>"100110101",
  11711=>"000101001",
  11712=>"010010011",
  11713=>"100000100",
  11714=>"000000101",
  11715=>"110011010",
  11716=>"010001000",
  11717=>"100001100",
  11718=>"000011011",
  11719=>"110010010",
  11720=>"000000010",
  11721=>"100110011",
  11722=>"101101101",
  11723=>"111001010",
  11724=>"011010111",
  11725=>"011011110",
  11726=>"000000110",
  11727=>"110010100",
  11728=>"011101101",
  11729=>"111101001",
  11730=>"001100000",
  11731=>"000000000",
  11732=>"100110100",
  11733=>"011010110",
  11734=>"110011001",
  11735=>"000110010",
  11736=>"001110001",
  11737=>"110110011",
  11738=>"101110001",
  11739=>"000111000",
  11740=>"000110110",
  11741=>"010011000",
  11742=>"010001110",
  11743=>"111011111",
  11744=>"000110001",
  11745=>"100110000",
  11746=>"101001100",
  11747=>"101000001",
  11748=>"001010111",
  11749=>"110110111",
  11750=>"110000011",
  11751=>"001110001",
  11752=>"010000001",
  11753=>"011011110",
  11754=>"011010010",
  11755=>"000111011",
  11756=>"001110000",
  11757=>"100111101",
  11758=>"011011000",
  11759=>"010110010",
  11760=>"100001010",
  11761=>"010111101",
  11762=>"010101111",
  11763=>"000000101",
  11764=>"000100100",
  11765=>"110101000",
  11766=>"101100110",
  11767=>"001111010",
  11768=>"000100101",
  11769=>"101101110",
  11770=>"010101010",
  11771=>"100011101",
  11772=>"000010010",
  11773=>"010011101",
  11774=>"001101100",
  11775=>"010111010",
  11776=>"100000011",
  11777=>"100111110",
  11778=>"100011111",
  11779=>"001011000",
  11780=>"101101001",
  11781=>"110100010",
  11782=>"101111111",
  11783=>"111100101",
  11784=>"001110101",
  11785=>"111111101",
  11786=>"111100100",
  11787=>"111001100",
  11788=>"000010101",
  11789=>"100010101",
  11790=>"101011101",
  11791=>"001110101",
  11792=>"111000111",
  11793=>"011001011",
  11794=>"101000011",
  11795=>"001101100",
  11796=>"001011111",
  11797=>"010000011",
  11798=>"001010010",
  11799=>"111111110",
  11800=>"110101110",
  11801=>"000011111",
  11802=>"110010101",
  11803=>"111110010",
  11804=>"100010011",
  11805=>"000000001",
  11806=>"000010110",
  11807=>"111010110",
  11808=>"001011101",
  11809=>"001100001",
  11810=>"001001010",
  11811=>"100001000",
  11812=>"001100101",
  11813=>"100111001",
  11814=>"000101101",
  11815=>"100110000",
  11816=>"010001000",
  11817=>"110111101",
  11818=>"001010011",
  11819=>"010110011",
  11820=>"000100111",
  11821=>"000010000",
  11822=>"100110010",
  11823=>"011000110",
  11824=>"110001111",
  11825=>"001010111",
  11826=>"000010001",
  11827=>"010110101",
  11828=>"111111101",
  11829=>"010001111",
  11830=>"010100101",
  11831=>"001101010",
  11832=>"101101011",
  11833=>"111111000",
  11834=>"000001111",
  11835=>"001110110",
  11836=>"011010111",
  11837=>"110101101",
  11838=>"111001011",
  11839=>"000011010",
  11840=>"011001111",
  11841=>"011101111",
  11842=>"011010001",
  11843=>"011110101",
  11844=>"010010110",
  11845=>"000010110",
  11846=>"100011001",
  11847=>"100000001",
  11848=>"011010111",
  11849=>"111110001",
  11850=>"000010011",
  11851=>"100111011",
  11852=>"000010011",
  11853=>"001001001",
  11854=>"101110000",
  11855=>"101110100",
  11856=>"101010110",
  11857=>"100100001",
  11858=>"001001011",
  11859=>"101100111",
  11860=>"101001111",
  11861=>"000011100",
  11862=>"100101001",
  11863=>"010011100",
  11864=>"011000011",
  11865=>"001000101",
  11866=>"001011110",
  11867=>"000000000",
  11868=>"110111010",
  11869=>"000101001",
  11870=>"111111000",
  11871=>"011101111",
  11872=>"110111011",
  11873=>"010011001",
  11874=>"000111110",
  11875=>"011000100",
  11876=>"111100001",
  11877=>"111000010",
  11878=>"000111000",
  11879=>"111101001",
  11880=>"101110100",
  11881=>"110001010",
  11882=>"000101011",
  11883=>"100001000",
  11884=>"111101011",
  11885=>"111100110",
  11886=>"100010100",
  11887=>"000101110",
  11888=>"001011101",
  11889=>"100111011",
  11890=>"111100101",
  11891=>"010000000",
  11892=>"011110011",
  11893=>"011100101",
  11894=>"011101011",
  11895=>"111111111",
  11896=>"000010001",
  11897=>"011011001",
  11898=>"000000010",
  11899=>"110010101",
  11900=>"110111000",
  11901=>"111100101",
  11902=>"000001101",
  11903=>"000100010",
  11904=>"101001011",
  11905=>"001110000",
  11906=>"001110011",
  11907=>"011111011",
  11908=>"001111101",
  11909=>"101100100",
  11910=>"111100010",
  11911=>"111110011",
  11912=>"000000010",
  11913=>"010110100",
  11914=>"100101110",
  11915=>"101001101",
  11916=>"001001100",
  11917=>"000111111",
  11918=>"000100011",
  11919=>"001000001",
  11920=>"100000000",
  11921=>"000100001",
  11922=>"000011010",
  11923=>"001110000",
  11924=>"110011011",
  11925=>"101010100",
  11926=>"001000101",
  11927=>"000111110",
  11928=>"101011011",
  11929=>"001001000",
  11930=>"100110101",
  11931=>"001001110",
  11932=>"100011001",
  11933=>"010111101",
  11934=>"110100001",
  11935=>"001001011",
  11936=>"101101110",
  11937=>"111110000",
  11938=>"101110011",
  11939=>"000100001",
  11940=>"001110101",
  11941=>"011111011",
  11942=>"011100000",
  11943=>"000011010",
  11944=>"101111000",
  11945=>"001010001",
  11946=>"001100000",
  11947=>"001010100",
  11948=>"000100010",
  11949=>"111110110",
  11950=>"001111000",
  11951=>"100111001",
  11952=>"000101001",
  11953=>"100011000",
  11954=>"000101010",
  11955=>"010001001",
  11956=>"011111010",
  11957=>"000011011",
  11958=>"011001000",
  11959=>"000111110",
  11960=>"011001100",
  11961=>"011111011",
  11962=>"001000000",
  11963=>"001101011",
  11964=>"100011010",
  11965=>"111001001",
  11966=>"010111001",
  11967=>"000111111",
  11968=>"011001010",
  11969=>"101110011",
  11970=>"011101000",
  11971=>"101011110",
  11972=>"010110110",
  11973=>"011001001",
  11974=>"101110111",
  11975=>"010100110",
  11976=>"010011010",
  11977=>"110101100",
  11978=>"110100110",
  11979=>"000001010",
  11980=>"010110011",
  11981=>"101011111",
  11982=>"101110011",
  11983=>"101000110",
  11984=>"111111111",
  11985=>"010000101",
  11986=>"001100000",
  11987=>"011111000",
  11988=>"000101010",
  11989=>"010011000",
  11990=>"010000000",
  11991=>"011011110",
  11992=>"110001111",
  11993=>"110101011",
  11994=>"000110001",
  11995=>"101010001",
  11996=>"111111101",
  11997=>"000011000",
  11998=>"101101011",
  11999=>"010000101",
  12000=>"000011110",
  12001=>"100111100",
  12002=>"001111000",
  12003=>"100100111",
  12004=>"000110011",
  12005=>"000000110",
  12006=>"000010001",
  12007=>"000111001",
  12008=>"101001110",
  12009=>"110000001",
  12010=>"101101000",
  12011=>"001110001",
  12012=>"000000000",
  12013=>"101001010",
  12014=>"000000000",
  12015=>"011101011",
  12016=>"000110001",
  12017=>"111111001",
  12018=>"001101101",
  12019=>"110001011",
  12020=>"100101110",
  12021=>"111001000",
  12022=>"111100110",
  12023=>"111010010",
  12024=>"110101100",
  12025=>"111100111",
  12026=>"101111100",
  12027=>"101001011",
  12028=>"000000100",
  12029=>"111100110",
  12030=>"100111110",
  12031=>"101000110",
  12032=>"101001001",
  12033=>"000100010",
  12034=>"010000011",
  12035=>"000111001",
  12036=>"000011111",
  12037=>"000100010",
  12038=>"100110010",
  12039=>"110101011",
  12040=>"110001100",
  12041=>"011111101",
  12042=>"110100001",
  12043=>"100110111",
  12044=>"010111100",
  12045=>"110011110",
  12046=>"100110010",
  12047=>"110101111",
  12048=>"101111001",
  12049=>"101011010",
  12050=>"101010010",
  12051=>"010101111",
  12052=>"101010010",
  12053=>"100110110",
  12054=>"101000001",
  12055=>"001111011",
  12056=>"011111001",
  12057=>"010000011",
  12058=>"100101011",
  12059=>"000010000",
  12060=>"001110010",
  12061=>"001000110",
  12062=>"000001110",
  12063=>"011101011",
  12064=>"011000000",
  12065=>"000100110",
  12066=>"011101111",
  12067=>"001001111",
  12068=>"011101111",
  12069=>"110000010",
  12070=>"011100110",
  12071=>"001001101",
  12072=>"011111001",
  12073=>"001000100",
  12074=>"101000101",
  12075=>"101001001",
  12076=>"000000101",
  12077=>"000110101",
  12078=>"110100111",
  12079=>"110010011",
  12080=>"111011111",
  12081=>"101001000",
  12082=>"010000000",
  12083=>"111000100",
  12084=>"111000001",
  12085=>"001000010",
  12086=>"110101011",
  12087=>"100000010",
  12088=>"111011100",
  12089=>"001110100",
  12090=>"101011001",
  12091=>"000010011",
  12092=>"000011111",
  12093=>"100001111",
  12094=>"001010101",
  12095=>"001100110",
  12096=>"001001101",
  12097=>"010000101",
  12098=>"100100001",
  12099=>"110100000",
  12100=>"001000101",
  12101=>"101101110",
  12102=>"001000011",
  12103=>"101101000",
  12104=>"011001101",
  12105=>"111000001",
  12106=>"111101111",
  12107=>"110101001",
  12108=>"000000000",
  12109=>"000011111",
  12110=>"010001010",
  12111=>"000101001",
  12112=>"001110011",
  12113=>"100010110",
  12114=>"100101001",
  12115=>"100011011",
  12116=>"011001011",
  12117=>"010101001",
  12118=>"100010100",
  12119=>"001000110",
  12120=>"010001100",
  12121=>"000010000",
  12122=>"100010110",
  12123=>"111101110",
  12124=>"111101011",
  12125=>"111001101",
  12126=>"001011011",
  12127=>"100000000",
  12128=>"111010110",
  12129=>"101001101",
  12130=>"100110111",
  12131=>"101011110",
  12132=>"111010100",
  12133=>"100011000",
  12134=>"000000101",
  12135=>"111111110",
  12136=>"001111100",
  12137=>"111010010",
  12138=>"010010000",
  12139=>"110000100",
  12140=>"101000000",
  12141=>"000000011",
  12142=>"111101110",
  12143=>"010101001",
  12144=>"000100111",
  12145=>"100000000",
  12146=>"100011110",
  12147=>"011001100",
  12148=>"111111000",
  12149=>"001001101",
  12150=>"101111111",
  12151=>"001001110",
  12152=>"111110001",
  12153=>"000110101",
  12154=>"000011110",
  12155=>"111001101",
  12156=>"110000001",
  12157=>"110001100",
  12158=>"100110110",
  12159=>"001001010",
  12160=>"100110100",
  12161=>"111001001",
  12162=>"011110110",
  12163=>"100100100",
  12164=>"000101000",
  12165=>"010000111",
  12166=>"111000000",
  12167=>"101000011",
  12168=>"010001100",
  12169=>"001101110",
  12170=>"100100000",
  12171=>"000011000",
  12172=>"010000001",
  12173=>"000011111",
  12174=>"011110101",
  12175=>"100110000",
  12176=>"010111001",
  12177=>"010100111",
  12178=>"001000000",
  12179=>"000100101",
  12180=>"000000000",
  12181=>"101000011",
  12182=>"011101011",
  12183=>"001010001",
  12184=>"111111000",
  12185=>"001001001",
  12186=>"001010110",
  12187=>"000010000",
  12188=>"000100111",
  12189=>"000001000",
  12190=>"000000011",
  12191=>"111000011",
  12192=>"100110010",
  12193=>"011101111",
  12194=>"110110110",
  12195=>"000101011",
  12196=>"010001001",
  12197=>"110110011",
  12198=>"001011110",
  12199=>"001111100",
  12200=>"000100100",
  12201=>"001000100",
  12202=>"111100101",
  12203=>"010111110",
  12204=>"000010011",
  12205=>"010100001",
  12206=>"111100100",
  12207=>"111100010",
  12208=>"111000011",
  12209=>"101001010",
  12210=>"011111001",
  12211=>"101000011",
  12212=>"101100110",
  12213=>"100001110",
  12214=>"111010001",
  12215=>"101100110",
  12216=>"100000000",
  12217=>"110011101",
  12218=>"110100100",
  12219=>"010111100",
  12220=>"110100100",
  12221=>"100001110",
  12222=>"100011110",
  12223=>"001001101",
  12224=>"010010010",
  12225=>"000010111",
  12226=>"000111110",
  12227=>"011010001",
  12228=>"111010111",
  12229=>"110010111",
  12230=>"111110100",
  12231=>"100001100",
  12232=>"100010000",
  12233=>"101011010",
  12234=>"111100110",
  12235=>"011001111",
  12236=>"000000010",
  12237=>"000100001",
  12238=>"111110101",
  12239=>"101000010",
  12240=>"110100111",
  12241=>"000111010",
  12242=>"101011101",
  12243=>"101010000",
  12244=>"110100110",
  12245=>"111100000",
  12246=>"000110000",
  12247=>"000000010",
  12248=>"011001001",
  12249=>"001101101",
  12250=>"011000111",
  12251=>"100001010",
  12252=>"110001000",
  12253=>"001000000",
  12254=>"110110011",
  12255=>"100110001",
  12256=>"110010100",
  12257=>"000110111",
  12258=>"001101011",
  12259=>"011000100",
  12260=>"000101010",
  12261=>"110010001",
  12262=>"010101110",
  12263=>"000111011",
  12264=>"001110000",
  12265=>"000010011",
  12266=>"100110000",
  12267=>"101101000",
  12268=>"000111011",
  12269=>"100011110",
  12270=>"000010010",
  12271=>"001010100",
  12272=>"110010001",
  12273=>"101011011",
  12274=>"000100001",
  12275=>"100100110",
  12276=>"111010001",
  12277=>"111001011",
  12278=>"100010101",
  12279=>"000110010",
  12280=>"010100000",
  12281=>"110001010",
  12282=>"111011001",
  12283=>"111110001",
  12284=>"110101010",
  12285=>"010101011",
  12286=>"000001100",
  12287=>"011101101",
  12288=>"110010011",
  12289=>"100101100",
  12290=>"110011011",
  12291=>"110100110",
  12292=>"001000000",
  12293=>"100110000",
  12294=>"101110101",
  12295=>"100001010",
  12296=>"000000100",
  12297=>"000010010",
  12298=>"000010101",
  12299=>"001001111",
  12300=>"111101101",
  12301=>"010000100",
  12302=>"001111111",
  12303=>"111011011",
  12304=>"000001011",
  12305=>"101100001",
  12306=>"110101110",
  12307=>"001011011",
  12308=>"101010000",
  12309=>"011111010",
  12310=>"000110011",
  12311=>"011100110",
  12312=>"111001100",
  12313=>"001010001",
  12314=>"000010111",
  12315=>"100111101",
  12316=>"011010011",
  12317=>"001000011",
  12318=>"110100000",
  12319=>"110010011",
  12320=>"011101000",
  12321=>"110111100",
  12322=>"000001101",
  12323=>"011110100",
  12324=>"110010101",
  12325=>"010101111",
  12326=>"110111111",
  12327=>"110100111",
  12328=>"101101001",
  12329=>"100110011",
  12330=>"111010001",
  12331=>"000000111",
  12332=>"011011011",
  12333=>"111111001",
  12334=>"100000100",
  12335=>"010100000",
  12336=>"000010101",
  12337=>"011000010",
  12338=>"110011001",
  12339=>"100111010",
  12340=>"101001000",
  12341=>"011101000",
  12342=>"111111100",
  12343=>"010101111",
  12344=>"010001000",
  12345=>"101011100",
  12346=>"001101110",
  12347=>"111011000",
  12348=>"110001001",
  12349=>"100011101",
  12350=>"111100000",
  12351=>"001001100",
  12352=>"011101000",
  12353=>"101010110",
  12354=>"101001110",
  12355=>"001100101",
  12356=>"000110011",
  12357=>"101101000",
  12358=>"011101100",
  12359=>"010101011",
  12360=>"001011100",
  12361=>"100000000",
  12362=>"000011110",
  12363=>"000110000",
  12364=>"001001111",
  12365=>"110011110",
  12366=>"011111000",
  12367=>"110101111",
  12368=>"111010111",
  12369=>"001110000",
  12370=>"111110111",
  12371=>"000001101",
  12372=>"111111010",
  12373=>"000010101",
  12374=>"100001111",
  12375=>"110001100",
  12376=>"011101101",
  12377=>"111000111",
  12378=>"100101000",
  12379=>"100101011",
  12380=>"001100100",
  12381=>"011100011",
  12382=>"111000000",
  12383=>"011010110",
  12384=>"010011011",
  12385=>"110011010",
  12386=>"000101001",
  12387=>"111010010",
  12388=>"101111101",
  12389=>"110111011",
  12390=>"100111111",
  12391=>"111100100",
  12392=>"111100001",
  12393=>"101000100",
  12394=>"001100010",
  12395=>"100010111",
  12396=>"111110001",
  12397=>"010001001",
  12398=>"111101101",
  12399=>"101110101",
  12400=>"111011111",
  12401=>"011011101",
  12402=>"101001110",
  12403=>"001100111",
  12404=>"110110101",
  12405=>"000010101",
  12406=>"000001100",
  12407=>"100111011",
  12408=>"001011011",
  12409=>"101010110",
  12410=>"011110011",
  12411=>"110101100",
  12412=>"001010011",
  12413=>"001111100",
  12414=>"010111010",
  12415=>"110111010",
  12416=>"100110000",
  12417=>"100000000",
  12418=>"011001100",
  12419=>"010010001",
  12420=>"110111010",
  12421=>"001110001",
  12422=>"111101010",
  12423=>"001101000",
  12424=>"101100110",
  12425=>"110000110",
  12426=>"100011110",
  12427=>"010111111",
  12428=>"000100011",
  12429=>"011110111",
  12430=>"111111011",
  12431=>"011011100",
  12432=>"010011111",
  12433=>"101110010",
  12434=>"111001110",
  12435=>"111010011",
  12436=>"000100110",
  12437=>"111111111",
  12438=>"011000000",
  12439=>"010001011",
  12440=>"010110011",
  12441=>"101110101",
  12442=>"000000100",
  12443=>"000110001",
  12444=>"010010000",
  12445=>"000101000",
  12446=>"010101111",
  12447=>"100011001",
  12448=>"000000010",
  12449=>"111001011",
  12450=>"011100101",
  12451=>"111000100",
  12452=>"011001011",
  12453=>"001101110",
  12454=>"110000010",
  12455=>"100100111",
  12456=>"000000101",
  12457=>"110101000",
  12458=>"011101000",
  12459=>"011101101",
  12460=>"000111011",
  12461=>"110100110",
  12462=>"001001001",
  12463=>"001001001",
  12464=>"000000100",
  12465=>"000000000",
  12466=>"010101111",
  12467=>"000000110",
  12468=>"010111010",
  12469=>"011001001",
  12470=>"010111010",
  12471=>"001011100",
  12472=>"111111111",
  12473=>"000000011",
  12474=>"100101100",
  12475=>"011000001",
  12476=>"010101100",
  12477=>"011111000",
  12478=>"000110001",
  12479=>"110001100",
  12480=>"110111110",
  12481=>"001110101",
  12482=>"011101111",
  12483=>"101101011",
  12484=>"001000001",
  12485=>"000101100",
  12486=>"101110110",
  12487=>"010010101",
  12488=>"101011011",
  12489=>"010000110",
  12490=>"001001001",
  12491=>"100011110",
  12492=>"111100110",
  12493=>"100110110",
  12494=>"101110110",
  12495=>"000000011",
  12496=>"000110111",
  12497=>"001101100",
  12498=>"111110001",
  12499=>"101110011",
  12500=>"010011001",
  12501=>"101111111",
  12502=>"101000010",
  12503=>"001110000",
  12504=>"100011011",
  12505=>"000100110",
  12506=>"100001101",
  12507=>"001000001",
  12508=>"111010000",
  12509=>"000101001",
  12510=>"000101001",
  12511=>"100101001",
  12512=>"000110000",
  12513=>"111101110",
  12514=>"100011100",
  12515=>"111010011",
  12516=>"010100000",
  12517=>"110100110",
  12518=>"111110000",
  12519=>"001011001",
  12520=>"111001011",
  12521=>"101101111",
  12522=>"111000001",
  12523=>"110001111",
  12524=>"000001011",
  12525=>"000110101",
  12526=>"001110111",
  12527=>"010000000",
  12528=>"110110110",
  12529=>"110010000",
  12530=>"101111000",
  12531=>"011111111",
  12532=>"100101110",
  12533=>"000001010",
  12534=>"011001010",
  12535=>"011000000",
  12536=>"001100110",
  12537=>"010110110",
  12538=>"001111000",
  12539=>"000000000",
  12540=>"000100110",
  12541=>"000010010",
  12542=>"100101000",
  12543=>"101001001",
  12544=>"111110000",
  12545=>"101101111",
  12546=>"101001100",
  12547=>"000100010",
  12548=>"110001011",
  12549=>"110111100",
  12550=>"111011010",
  12551=>"111111010",
  12552=>"111011111",
  12553=>"101101001",
  12554=>"001000001",
  12555=>"001011000",
  12556=>"100110111",
  12557=>"010001100",
  12558=>"100100010",
  12559=>"000010000",
  12560=>"101111111",
  12561=>"000011010",
  12562=>"110110110",
  12563=>"001001000",
  12564=>"001011001",
  12565=>"010000111",
  12566=>"011011011",
  12567=>"111011111",
  12568=>"101000110",
  12569=>"110111111",
  12570=>"000110101",
  12571=>"011110011",
  12572=>"101100011",
  12573=>"001111001",
  12574=>"011001011",
  12575=>"101001000",
  12576=>"010111011",
  12577=>"111101001",
  12578=>"011111010",
  12579=>"111011010",
  12580=>"010100010",
  12581=>"000111011",
  12582=>"001100100",
  12583=>"001111101",
  12584=>"100000001",
  12585=>"110001001",
  12586=>"100100101",
  12587=>"011110111",
  12588=>"001000011",
  12589=>"110110000",
  12590=>"001100100",
  12591=>"001001011",
  12592=>"010010101",
  12593=>"100010010",
  12594=>"111111000",
  12595=>"101010101",
  12596=>"110111110",
  12597=>"110100011",
  12598=>"011011001",
  12599=>"011000001",
  12600=>"011110100",
  12601=>"111111110",
  12602=>"010000111",
  12603=>"000000100",
  12604=>"000000001",
  12605=>"001111011",
  12606=>"011001110",
  12607=>"100110001",
  12608=>"010101110",
  12609=>"010000111",
  12610=>"001110110",
  12611=>"001111011",
  12612=>"101010011",
  12613=>"000111100",
  12614=>"101100000",
  12615=>"000001101",
  12616=>"010101010",
  12617=>"111001100",
  12618=>"000101110",
  12619=>"000000000",
  12620=>"000101100",
  12621=>"101100001",
  12622=>"100111001",
  12623=>"001110100",
  12624=>"111001000",
  12625=>"000111011",
  12626=>"110101111",
  12627=>"111001111",
  12628=>"011000011",
  12629=>"110000111",
  12630=>"100001100",
  12631=>"101010100",
  12632=>"001001100",
  12633=>"100111001",
  12634=>"000110001",
  12635=>"110101100",
  12636=>"110011011",
  12637=>"100000100",
  12638=>"110101110",
  12639=>"101100000",
  12640=>"110100100",
  12641=>"110110011",
  12642=>"000011101",
  12643=>"011111101",
  12644=>"111111000",
  12645=>"011110111",
  12646=>"010101100",
  12647=>"010110101",
  12648=>"010110111",
  12649=>"101001101",
  12650=>"110010111",
  12651=>"100111001",
  12652=>"000110111",
  12653=>"111111110",
  12654=>"110001101",
  12655=>"000000000",
  12656=>"010011110",
  12657=>"001010001",
  12658=>"011111111",
  12659=>"110010101",
  12660=>"110111100",
  12661=>"011101010",
  12662=>"111111011",
  12663=>"000110000",
  12664=>"101101001",
  12665=>"000001000",
  12666=>"101101000",
  12667=>"001100111",
  12668=>"101011100",
  12669=>"010100001",
  12670=>"110001011",
  12671=>"011100000",
  12672=>"000010101",
  12673=>"010011001",
  12674=>"101100101",
  12675=>"111001011",
  12676=>"100010111",
  12677=>"101000110",
  12678=>"011000100",
  12679=>"000000111",
  12680=>"001110000",
  12681=>"100001011",
  12682=>"001010010",
  12683=>"111101010",
  12684=>"011000111",
  12685=>"111000100",
  12686=>"000011000",
  12687=>"111010011",
  12688=>"000111011",
  12689=>"101110110",
  12690=>"100100110",
  12691=>"011111110",
  12692=>"000111100",
  12693=>"100100010",
  12694=>"011011100",
  12695=>"110000010",
  12696=>"000100000",
  12697=>"000111011",
  12698=>"111001010",
  12699=>"010011011",
  12700=>"011000111",
  12701=>"100010001",
  12702=>"101010101",
  12703=>"001000010",
  12704=>"110000010",
  12705=>"010100010",
  12706=>"100100011",
  12707=>"001000110",
  12708=>"111011010",
  12709=>"100100010",
  12710=>"101010001",
  12711=>"011110110",
  12712=>"001000000",
  12713=>"100110101",
  12714=>"100111111",
  12715=>"101111110",
  12716=>"100001100",
  12717=>"110111100",
  12718=>"011000101",
  12719=>"101110000",
  12720=>"110110000",
  12721=>"011100101",
  12722=>"000000110",
  12723=>"000110011",
  12724=>"001100001",
  12725=>"010001000",
  12726=>"000101010",
  12727=>"011000100",
  12728=>"110010010",
  12729=>"111111001",
  12730=>"101110111",
  12731=>"111100001",
  12732=>"100010011",
  12733=>"010100001",
  12734=>"011111011",
  12735=>"111000110",
  12736=>"001001010",
  12737=>"101000111",
  12738=>"101010001",
  12739=>"010101111",
  12740=>"101111111",
  12741=>"110110001",
  12742=>"101111010",
  12743=>"100110010",
  12744=>"100000001",
  12745=>"010001001",
  12746=>"010001101",
  12747=>"100011001",
  12748=>"100110101",
  12749=>"001101011",
  12750=>"110111111",
  12751=>"011001011",
  12752=>"101010001",
  12753=>"111100110",
  12754=>"001111100",
  12755=>"111010011",
  12756=>"100001111",
  12757=>"111011110",
  12758=>"111011100",
  12759=>"000010000",
  12760=>"000011010",
  12761=>"011011111",
  12762=>"010101101",
  12763=>"111011000",
  12764=>"110100100",
  12765=>"100101001",
  12766=>"110111011",
  12767=>"001101001",
  12768=>"101001000",
  12769=>"011000010",
  12770=>"000000100",
  12771=>"101000001",
  12772=>"010101100",
  12773=>"000010111",
  12774=>"111000011",
  12775=>"110010010",
  12776=>"011101011",
  12777=>"100101110",
  12778=>"111100000",
  12779=>"001111011",
  12780=>"011001110",
  12781=>"111000001",
  12782=>"101001001",
  12783=>"111000111",
  12784=>"010111010",
  12785=>"000110000",
  12786=>"001111000",
  12787=>"010111000",
  12788=>"111100010",
  12789=>"000111000",
  12790=>"010001110",
  12791=>"101111110",
  12792=>"110101010",
  12793=>"101011101",
  12794=>"111101001",
  12795=>"011000101",
  12796=>"111001111",
  12797=>"100000010",
  12798=>"001110000",
  12799=>"111000000",
  12800=>"010100111",
  12801=>"110000010",
  12802=>"100100111",
  12803=>"111010111",
  12804=>"010100010",
  12805=>"010000000",
  12806=>"110011001",
  12807=>"110111000",
  12808=>"111111100",
  12809=>"010000011",
  12810=>"111001001",
  12811=>"100001101",
  12812=>"001000000",
  12813=>"100110111",
  12814=>"000101101",
  12815=>"101001011",
  12816=>"111001101",
  12817=>"011101101",
  12818=>"100110111",
  12819=>"101010110",
  12820=>"111111011",
  12821=>"001011011",
  12822=>"101011000",
  12823=>"100001111",
  12824=>"011111111",
  12825=>"111000011",
  12826=>"100010111",
  12827=>"001011111",
  12828=>"100100100",
  12829=>"110100011",
  12830=>"111000111",
  12831=>"100000010",
  12832=>"010010101",
  12833=>"110100101",
  12834=>"001000011",
  12835=>"000100111",
  12836=>"110001101",
  12837=>"110000000",
  12838=>"001001100",
  12839=>"100101011",
  12840=>"010111011",
  12841=>"000010011",
  12842=>"000110101",
  12843=>"001100001",
  12844=>"111111101",
  12845=>"010011000",
  12846=>"010010111",
  12847=>"010001101",
  12848=>"011000100",
  12849=>"001111101",
  12850=>"100100111",
  12851=>"110001011",
  12852=>"110000110",
  12853=>"110000101",
  12854=>"010001000",
  12855=>"111100001",
  12856=>"101011100",
  12857=>"010100000",
  12858=>"001000001",
  12859=>"101111001",
  12860=>"011001101",
  12861=>"110010001",
  12862=>"100001011",
  12863=>"101001000",
  12864=>"000101011",
  12865=>"011110110",
  12866=>"011011100",
  12867=>"111100010",
  12868=>"111001110",
  12869=>"000000011",
  12870=>"000000000",
  12871=>"001011001",
  12872=>"100101110",
  12873=>"111101110",
  12874=>"000100110",
  12875=>"010111011",
  12876=>"100100001",
  12877=>"111100111",
  12878=>"011000100",
  12879=>"111100110",
  12880=>"010000010",
  12881=>"010110001",
  12882=>"000011000",
  12883=>"111000101",
  12884=>"111011011",
  12885=>"101000000",
  12886=>"100010100",
  12887=>"010110111",
  12888=>"001101100",
  12889=>"101001000",
  12890=>"011110010",
  12891=>"101001011",
  12892=>"101100100",
  12893=>"000100010",
  12894=>"011000111",
  12895=>"111110110",
  12896=>"101000100",
  12897=>"111011010",
  12898=>"011011100",
  12899=>"100011101",
  12900=>"111100110",
  12901=>"111111110",
  12902=>"011101001",
  12903=>"011111000",
  12904=>"101101101",
  12905=>"101110101",
  12906=>"001011010",
  12907=>"101001000",
  12908=>"110001100",
  12909=>"001110110",
  12910=>"010100001",
  12911=>"000000010",
  12912=>"101011100",
  12913=>"101010000",
  12914=>"101000100",
  12915=>"001100000",
  12916=>"011011001",
  12917=>"100110101",
  12918=>"000110000",
  12919=>"011111001",
  12920=>"101110110",
  12921=>"010000100",
  12922=>"111101010",
  12923=>"100100000",
  12924=>"001001110",
  12925=>"001000000",
  12926=>"111010101",
  12927=>"011101111",
  12928=>"100111000",
  12929=>"100001110",
  12930=>"100110111",
  12931=>"110110101",
  12932=>"010110101",
  12933=>"011110010",
  12934=>"101000001",
  12935=>"110101111",
  12936=>"000011111",
  12937=>"101110101",
  12938=>"010010010",
  12939=>"010101001",
  12940=>"000100000",
  12941=>"010000010",
  12942=>"010101101",
  12943=>"010100101",
  12944=>"110111111",
  12945=>"100011011",
  12946=>"101111011",
  12947=>"111011111",
  12948=>"001100001",
  12949=>"110011100",
  12950=>"110010100",
  12951=>"011010100",
  12952=>"111100100",
  12953=>"000101001",
  12954=>"111110110",
  12955=>"111011011",
  12956=>"000000110",
  12957=>"000111101",
  12958=>"000000010",
  12959=>"011010011",
  12960=>"101011000",
  12961=>"101000101",
  12962=>"100011100",
  12963=>"000101010",
  12964=>"111001000",
  12965=>"011111101",
  12966=>"100011110",
  12967=>"001101100",
  12968=>"111011010",
  12969=>"010111111",
  12970=>"000111001",
  12971=>"011000010",
  12972=>"101000011",
  12973=>"010100001",
  12974=>"110000011",
  12975=>"101001001",
  12976=>"011001100",
  12977=>"100101010",
  12978=>"111010010",
  12979=>"101101011",
  12980=>"101000010",
  12981=>"000010011",
  12982=>"010011101",
  12983=>"110011101",
  12984=>"011001001",
  12985=>"110011110",
  12986=>"010000011",
  12987=>"000110100",
  12988=>"010001101",
  12989=>"001000111",
  12990=>"001100000",
  12991=>"010101000",
  12992=>"110010101",
  12993=>"000100100",
  12994=>"101110001",
  12995=>"001001011",
  12996=>"111111110",
  12997=>"100001101",
  12998=>"001110111",
  12999=>"101000010",
  13000=>"010011111",
  13001=>"010111110",
  13002=>"111100010",
  13003=>"110011100",
  13004=>"011010011",
  13005=>"101100111",
  13006=>"110010010",
  13007=>"000001001",
  13008=>"011011111",
  13009=>"001110010",
  13010=>"000000111",
  13011=>"010001101",
  13012=>"101001101",
  13013=>"111010001",
  13014=>"011001011",
  13015=>"001011111",
  13016=>"000111001",
  13017=>"101111111",
  13018=>"000101111",
  13019=>"101001001",
  13020=>"111100010",
  13021=>"101100100",
  13022=>"111110110",
  13023=>"100011010",
  13024=>"110100111",
  13025=>"110111101",
  13026=>"110000110",
  13027=>"001111110",
  13028=>"000001001",
  13029=>"001100001",
  13030=>"100110010",
  13031=>"001010000",
  13032=>"010110110",
  13033=>"001111010",
  13034=>"101000100",
  13035=>"100011011",
  13036=>"101101101",
  13037=>"000001001",
  13038=>"001000100",
  13039=>"011001101",
  13040=>"111110000",
  13041=>"101001101",
  13042=>"010001001",
  13043=>"100000010",
  13044=>"110111011",
  13045=>"010111000",
  13046=>"000101111",
  13047=>"111011101",
  13048=>"010111111",
  13049=>"110000001",
  13050=>"000100001",
  13051=>"111110110",
  13052=>"111001010",
  13053=>"001100000",
  13054=>"000001011",
  13055=>"111111100",
  13056=>"111110110",
  13057=>"110101101",
  13058=>"101110110",
  13059=>"100011110",
  13060=>"000011111",
  13061=>"111110000",
  13062=>"111111001",
  13063=>"101001011",
  13064=>"000001011",
  13065=>"010010111",
  13066=>"111110101",
  13067=>"010001101",
  13068=>"110010110",
  13069=>"101001001",
  13070=>"011101010",
  13071=>"000100011",
  13072=>"000010001",
  13073=>"000101000",
  13074=>"011010101",
  13075=>"110101010",
  13076=>"101001110",
  13077=>"000111001",
  13078=>"111011011",
  13079=>"110000010",
  13080=>"100111000",
  13081=>"000000000",
  13082=>"111111101",
  13083=>"001100010",
  13084=>"101111001",
  13085=>"011000011",
  13086=>"011000010",
  13087=>"010100101",
  13088=>"011110101",
  13089=>"100110000",
  13090=>"100110001",
  13091=>"110101011",
  13092=>"000000010",
  13093=>"110001100",
  13094=>"110111101",
  13095=>"111010010",
  13096=>"101001010",
  13097=>"000000001",
  13098=>"111100100",
  13099=>"100001000",
  13100=>"111000101",
  13101=>"111011010",
  13102=>"100000001",
  13103=>"110101010",
  13104=>"010100011",
  13105=>"111111010",
  13106=>"111110011",
  13107=>"001000101",
  13108=>"110100010",
  13109=>"001010100",
  13110=>"110111000",
  13111=>"110011111",
  13112=>"101101100",
  13113=>"000010001",
  13114=>"000000101",
  13115=>"111011001",
  13116=>"100011111",
  13117=>"101110001",
  13118=>"011011110",
  13119=>"111111110",
  13120=>"110111110",
  13121=>"110010001",
  13122=>"011000010",
  13123=>"010011100",
  13124=>"000011101",
  13125=>"001011110",
  13126=>"010011001",
  13127=>"010010100",
  13128=>"000001101",
  13129=>"110101100",
  13130=>"110101101",
  13131=>"100010010",
  13132=>"011001001",
  13133=>"000110100",
  13134=>"000001100",
  13135=>"100000011",
  13136=>"111111111",
  13137=>"000100011",
  13138=>"000000011",
  13139=>"010100111",
  13140=>"100100010",
  13141=>"111000111",
  13142=>"111101100",
  13143=>"100111001",
  13144=>"111101111",
  13145=>"001000111",
  13146=>"101101001",
  13147=>"110101000",
  13148=>"101101000",
  13149=>"001010001",
  13150=>"001101001",
  13151=>"010000100",
  13152=>"111101010",
  13153=>"000001100",
  13154=>"110000111",
  13155=>"001100001",
  13156=>"000000101",
  13157=>"001000001",
  13158=>"011000100",
  13159=>"000110000",
  13160=>"101010001",
  13161=>"000000101",
  13162=>"101011110",
  13163=>"000111101",
  13164=>"101100000",
  13165=>"000000000",
  13166=>"010110001",
  13167=>"010010011",
  13168=>"011010010",
  13169=>"110000001",
  13170=>"010010001",
  13171=>"101011000",
  13172=>"001100100",
  13173=>"111100111",
  13174=>"111010000",
  13175=>"110101001",
  13176=>"000000011",
  13177=>"000010011",
  13178=>"111100000",
  13179=>"111110000",
  13180=>"010001111",
  13181=>"011100001",
  13182=>"001110001",
  13183=>"111110111",
  13184=>"110101110",
  13185=>"000100100",
  13186=>"101100101",
  13187=>"001010001",
  13188=>"001001000",
  13189=>"110101000",
  13190=>"111011111",
  13191=>"010101111",
  13192=>"001011101",
  13193=>"101011010",
  13194=>"000100000",
  13195=>"111011000",
  13196=>"111110010",
  13197=>"000011011",
  13198=>"010001010",
  13199=>"011110100",
  13200=>"011000001",
  13201=>"000000010",
  13202=>"000000110",
  13203=>"100000111",
  13204=>"011110001",
  13205=>"001011000",
  13206=>"100011111",
  13207=>"011111011",
  13208=>"111011101",
  13209=>"000010010",
  13210=>"111010110",
  13211=>"011000110",
  13212=>"001011000",
  13213=>"100101001",
  13214=>"100011110",
  13215=>"010101000",
  13216=>"011101110",
  13217=>"110011110",
  13218=>"010111110",
  13219=>"111110000",
  13220=>"110001101",
  13221=>"000110010",
  13222=>"100000100",
  13223=>"011100111",
  13224=>"100001011",
  13225=>"010011110",
  13226=>"010101101",
  13227=>"101110110",
  13228=>"111001101",
  13229=>"111101011",
  13230=>"111101001",
  13231=>"001110001",
  13232=>"010101000",
  13233=>"001010001",
  13234=>"011001111",
  13235=>"001001011",
  13236=>"000011000",
  13237=>"100100000",
  13238=>"001000100",
  13239=>"110110100",
  13240=>"100110001",
  13241=>"010101101",
  13242=>"100010101",
  13243=>"000010100",
  13244=>"100110010",
  13245=>"100100010",
  13246=>"001000001",
  13247=>"011110010",
  13248=>"100111010",
  13249=>"101001010",
  13250=>"010100100",
  13251=>"010100100",
  13252=>"000100011",
  13253=>"010000111",
  13254=>"010101111",
  13255=>"111011011",
  13256=>"000100000",
  13257=>"001101101",
  13258=>"101001001",
  13259=>"111101100",
  13260=>"101101101",
  13261=>"100010001",
  13262=>"100100010",
  13263=>"010110011",
  13264=>"101001111",
  13265=>"100110100",
  13266=>"110010001",
  13267=>"100011011",
  13268=>"111011100",
  13269=>"011001100",
  13270=>"111110110",
  13271=>"101100010",
  13272=>"111001010",
  13273=>"111000100",
  13274=>"100010100",
  13275=>"011010101",
  13276=>"111100000",
  13277=>"100101110",
  13278=>"001001100",
  13279=>"011100001",
  13280=>"111110001",
  13281=>"001100110",
  13282=>"011111001",
  13283=>"000001100",
  13284=>"001111110",
  13285=>"101011100",
  13286=>"000001011",
  13287=>"110000111",
  13288=>"011110111",
  13289=>"001010111",
  13290=>"111010010",
  13291=>"000000001",
  13292=>"001100111",
  13293=>"100110000",
  13294=>"111000011",
  13295=>"001001000",
  13296=>"000011101",
  13297=>"011000000",
  13298=>"110000111",
  13299=>"111101101",
  13300=>"000100110",
  13301=>"001000000",
  13302=>"101010000",
  13303=>"001000000",
  13304=>"000101100",
  13305=>"011011111",
  13306=>"100000101",
  13307=>"110101010",
  13308=>"001011111",
  13309=>"001111011",
  13310=>"110011111",
  13311=>"101101001",
  13312=>"110000010",
  13313=>"100111111",
  13314=>"110000100",
  13315=>"101101110",
  13316=>"000000110",
  13317=>"001101011",
  13318=>"101000111",
  13319=>"011011101",
  13320=>"011000001",
  13321=>"100111100",
  13322=>"011110000",
  13323=>"000000000",
  13324=>"111011001",
  13325=>"000001101",
  13326=>"010110000",
  13327=>"001010110",
  13328=>"100100101",
  13329=>"101010010",
  13330=>"110101111",
  13331=>"000010110",
  13332=>"101011001",
  13333=>"010001100",
  13334=>"111110001",
  13335=>"000100010",
  13336=>"101011101",
  13337=>"101111110",
  13338=>"111100111",
  13339=>"110001110",
  13340=>"000010100",
  13341=>"101011101",
  13342=>"100010010",
  13343=>"110100001",
  13344=>"100110110",
  13345=>"100101001",
  13346=>"000100100",
  13347=>"000110010",
  13348=>"001000110",
  13349=>"110011100",
  13350=>"100001001",
  13351=>"100010000",
  13352=>"110100000",
  13353=>"101100000",
  13354=>"111010111",
  13355=>"111001100",
  13356=>"101000000",
  13357=>"000101100",
  13358=>"110110101",
  13359=>"011111111",
  13360=>"101100100",
  13361=>"100100110",
  13362=>"100110001",
  13363=>"110100101",
  13364=>"101100000",
  13365=>"100100010",
  13366=>"010110111",
  13367=>"111110010",
  13368=>"010111011",
  13369=>"011101000",
  13370=>"111001010",
  13371=>"001011110",
  13372=>"111100000",
  13373=>"100111111",
  13374=>"011001000",
  13375=>"101011101",
  13376=>"101000011",
  13377=>"011011101",
  13378=>"110010011",
  13379=>"111100100",
  13380=>"110111011",
  13381=>"011101111",
  13382=>"110111100",
  13383=>"111010000",
  13384=>"011110110",
  13385=>"111101000",
  13386=>"011111010",
  13387=>"101101010",
  13388=>"011001011",
  13389=>"100111001",
  13390=>"100111011",
  13391=>"101100100",
  13392=>"110001010",
  13393=>"001011001",
  13394=>"010110100",
  13395=>"101010000",
  13396=>"000010101",
  13397=>"110111110",
  13398=>"101001101",
  13399=>"010010000",
  13400=>"100011001",
  13401=>"010110000",
  13402=>"001101010",
  13403=>"000110100",
  13404=>"100010111",
  13405=>"011111100",
  13406=>"110111000",
  13407=>"100011110",
  13408=>"101101000",
  13409=>"000100101",
  13410=>"110110110",
  13411=>"100001011",
  13412=>"100100001",
  13413=>"100111100",
  13414=>"001011001",
  13415=>"111111101",
  13416=>"101001100",
  13417=>"000001011",
  13418=>"001100010",
  13419=>"101000111",
  13420=>"000000110",
  13421=>"011011111",
  13422=>"000001100",
  13423=>"011001000",
  13424=>"011101001",
  13425=>"001110010",
  13426=>"000010000",
  13427=>"101010110",
  13428=>"101001000",
  13429=>"011010100",
  13430=>"001001001",
  13431=>"100000101",
  13432=>"011110011",
  13433=>"100010101",
  13434=>"111000110",
  13435=>"001111000",
  13436=>"001000001",
  13437=>"111000011",
  13438=>"101100001",
  13439=>"001010000",
  13440=>"110110111",
  13441=>"001110111",
  13442=>"000000011",
  13443=>"000001110",
  13444=>"101000000",
  13445=>"011011100",
  13446=>"101110110",
  13447=>"111100111",
  13448=>"110100001",
  13449=>"110111110",
  13450=>"001100111",
  13451=>"000101000",
  13452=>"010010000",
  13453=>"111010100",
  13454=>"011010010",
  13455=>"011000000",
  13456=>"111110011",
  13457=>"011101001",
  13458=>"111011001",
  13459=>"000100000",
  13460=>"101010000",
  13461=>"010011111",
  13462=>"011000100",
  13463=>"101111011",
  13464=>"011101000",
  13465=>"011101110",
  13466=>"110001001",
  13467=>"110101011",
  13468=>"101101100",
  13469=>"101100010",
  13470=>"110111101",
  13471=>"011010011",
  13472=>"100101101",
  13473=>"000000111",
  13474=>"110001010",
  13475=>"011110111",
  13476=>"011011100",
  13477=>"100111100",
  13478=>"010111011",
  13479=>"000011111",
  13480=>"000101011",
  13481=>"001111100",
  13482=>"101000101",
  13483=>"111000101",
  13484=>"000011111",
  13485=>"101110000",
  13486=>"000011000",
  13487=>"111101001",
  13488=>"001111001",
  13489=>"010001111",
  13490=>"010011100",
  13491=>"100101001",
  13492=>"100001010",
  13493=>"101101111",
  13494=>"110001100",
  13495=>"000011000",
  13496=>"101111010",
  13497=>"001101100",
  13498=>"110100010",
  13499=>"101011101",
  13500=>"110101101",
  13501=>"011000101",
  13502=>"000000001",
  13503=>"000100000",
  13504=>"110100011",
  13505=>"100100101",
  13506=>"000001101",
  13507=>"111101001",
  13508=>"011100101",
  13509=>"001000110",
  13510=>"100011110",
  13511=>"010011010",
  13512=>"010000011",
  13513=>"000111110",
  13514=>"111101110",
  13515=>"110101100",
  13516=>"011111011",
  13517=>"111100000",
  13518=>"010111101",
  13519=>"100101101",
  13520=>"001001101",
  13521=>"011101110",
  13522=>"010010001",
  13523=>"111001101",
  13524=>"001001011",
  13525=>"001010100",
  13526=>"010100101",
  13527=>"100110111",
  13528=>"000001011",
  13529=>"111111011",
  13530=>"111000001",
  13531=>"011001110",
  13532=>"010011111",
  13533=>"011010110",
  13534=>"000110110",
  13535=>"100110111",
  13536=>"110000111",
  13537=>"111111010",
  13538=>"000111110",
  13539=>"100010101",
  13540=>"000000100",
  13541=>"001101111",
  13542=>"000000010",
  13543=>"111011010",
  13544=>"100100100",
  13545=>"010111001",
  13546=>"111100101",
  13547=>"010111110",
  13548=>"100110110",
  13549=>"000001111",
  13550=>"110011111",
  13551=>"000101011",
  13552=>"000001111",
  13553=>"101010100",
  13554=>"011001110",
  13555=>"001100110",
  13556=>"101010001",
  13557=>"010011100",
  13558=>"010110111",
  13559=>"110001010",
  13560=>"000011001",
  13561=>"011010111",
  13562=>"101100000",
  13563=>"101011110",
  13564=>"010100010",
  13565=>"101100010",
  13566=>"011111111",
  13567=>"000000110",
  13568=>"001010010",
  13569=>"010010111",
  13570=>"101100110",
  13571=>"111111111",
  13572=>"110001111",
  13573=>"110111101",
  13574=>"110001101",
  13575=>"011111111",
  13576=>"110001110",
  13577=>"100100110",
  13578=>"100000101",
  13579=>"001000011",
  13580=>"011110110",
  13581=>"110010111",
  13582=>"010010011",
  13583=>"001000111",
  13584=>"010110101",
  13585=>"111101110",
  13586=>"111001010",
  13587=>"110110101",
  13588=>"111001001",
  13589=>"110101010",
  13590=>"001100000",
  13591=>"010101110",
  13592=>"000011110",
  13593=>"100110111",
  13594=>"010011010",
  13595=>"010000110",
  13596=>"100000001",
  13597=>"110101101",
  13598=>"111000011",
  13599=>"100101101",
  13600=>"011111001",
  13601=>"000010110",
  13602=>"000011011",
  13603=>"110111011",
  13604=>"011101001",
  13605=>"110110010",
  13606=>"101100111",
  13607=>"100110000",
  13608=>"110010111",
  13609=>"111100101",
  13610=>"111010110",
  13611=>"111010010",
  13612=>"111011000",
  13613=>"110100010",
  13614=>"100100001",
  13615=>"111100111",
  13616=>"100011110",
  13617=>"000010011",
  13618=>"000001100",
  13619=>"001110111",
  13620=>"111011000",
  13621=>"010111011",
  13622=>"111011001",
  13623=>"001000110",
  13624=>"010101101",
  13625=>"001000101",
  13626=>"100001011",
  13627=>"000100000",
  13628=>"110100000",
  13629=>"101110111",
  13630=>"101010111",
  13631=>"101001001",
  13632=>"110001011",
  13633=>"001010100",
  13634=>"101010000",
  13635=>"110101011",
  13636=>"101001011",
  13637=>"010110100",
  13638=>"001000001",
  13639=>"001001000",
  13640=>"001010001",
  13641=>"110101001",
  13642=>"101011110",
  13643=>"111101001",
  13644=>"110100100",
  13645=>"010000001",
  13646=>"000010101",
  13647=>"110011010",
  13648=>"010000000",
  13649=>"100101001",
  13650=>"110000111",
  13651=>"001000110",
  13652=>"101000100",
  13653=>"010101110",
  13654=>"100110001",
  13655=>"101111000",
  13656=>"011110110",
  13657=>"010110101",
  13658=>"010100000",
  13659=>"010111001",
  13660=>"010100111",
  13661=>"110110111",
  13662=>"111100011",
  13663=>"111100111",
  13664=>"111000101",
  13665=>"100000001",
  13666=>"000110101",
  13667=>"010011111",
  13668=>"110110000",
  13669=>"000101001",
  13670=>"111001100",
  13671=>"000011010",
  13672=>"010100101",
  13673=>"001101110",
  13674=>"111111111",
  13675=>"110111100",
  13676=>"000011110",
  13677=>"111000111",
  13678=>"111010000",
  13679=>"001010100",
  13680=>"001101100",
  13681=>"000011100",
  13682=>"111010101",
  13683=>"100011100",
  13684=>"111011011",
  13685=>"101000100",
  13686=>"001111010",
  13687=>"111110111",
  13688=>"011101110",
  13689=>"011011101",
  13690=>"111101000",
  13691=>"010110010",
  13692=>"010011100",
  13693=>"101111010",
  13694=>"101000000",
  13695=>"110101011",
  13696=>"110100001",
  13697=>"000100011",
  13698=>"000010110",
  13699=>"010001001",
  13700=>"011110011",
  13701=>"111011100",
  13702=>"111001011",
  13703=>"110000011",
  13704=>"011011110",
  13705=>"011100101",
  13706=>"000001011",
  13707=>"111011111",
  13708=>"100111001",
  13709=>"100101101",
  13710=>"100101101",
  13711=>"011000000",
  13712=>"011011100",
  13713=>"000011001",
  13714=>"011011101",
  13715=>"001011111",
  13716=>"100110000",
  13717=>"011011010",
  13718=>"000001010",
  13719=>"010111011",
  13720=>"110011110",
  13721=>"001101000",
  13722=>"010100111",
  13723=>"100011111",
  13724=>"111001111",
  13725=>"000110010",
  13726=>"000000010",
  13727=>"110000000",
  13728=>"011110011",
  13729=>"011111110",
  13730=>"000101101",
  13731=>"110011111",
  13732=>"011101011",
  13733=>"011010100",
  13734=>"001010000",
  13735=>"011101011",
  13736=>"111100010",
  13737=>"111101001",
  13738=>"111111111",
  13739=>"101010011",
  13740=>"100010110",
  13741=>"111110010",
  13742=>"000010101",
  13743=>"001011000",
  13744=>"111111001",
  13745=>"110001011",
  13746=>"011011101",
  13747=>"011101110",
  13748=>"100010110",
  13749=>"011000000",
  13750=>"101110100",
  13751=>"110110001",
  13752=>"001000101",
  13753=>"001001000",
  13754=>"011000010",
  13755=>"110100011",
  13756=>"111010000",
  13757=>"101000010",
  13758=>"000010000",
  13759=>"100010001",
  13760=>"100001111",
  13761=>"110010001",
  13762=>"111100001",
  13763=>"010000001",
  13764=>"110111011",
  13765=>"000011010",
  13766=>"011111001",
  13767=>"111101000",
  13768=>"000100011",
  13769=>"010010111",
  13770=>"010101111",
  13771=>"110100011",
  13772=>"100100101",
  13773=>"100100110",
  13774=>"000100110",
  13775=>"100100010",
  13776=>"011101001",
  13777=>"001110100",
  13778=>"100010011",
  13779=>"111010011",
  13780=>"110110000",
  13781=>"110100000",
  13782=>"000011100",
  13783=>"101100110",
  13784=>"000000001",
  13785=>"000000010",
  13786=>"001000010",
  13787=>"110110001",
  13788=>"010111000",
  13789=>"111011101",
  13790=>"111001001",
  13791=>"001101000",
  13792=>"011000001",
  13793=>"001000001",
  13794=>"101000000",
  13795=>"011110010",
  13796=>"011000000",
  13797=>"110010001",
  13798=>"010110000",
  13799=>"100011010",
  13800=>"011010011",
  13801=>"110001110",
  13802=>"001000101",
  13803=>"000100011",
  13804=>"111010100",
  13805=>"010000101",
  13806=>"101110101",
  13807=>"000100011",
  13808=>"111001001",
  13809=>"010110100",
  13810=>"000111000",
  13811=>"010111111",
  13812=>"111111100",
  13813=>"001001110",
  13814=>"001011010",
  13815=>"100111010",
  13816=>"111011101",
  13817=>"111010111",
  13818=>"100100011",
  13819=>"101111100",
  13820=>"000010111",
  13821=>"111111000",
  13822=>"101101001",
  13823=>"110010111",
  13824=>"111010001",
  13825=>"000010001",
  13826=>"011100111",
  13827=>"001110100",
  13828=>"010011001",
  13829=>"111011101",
  13830=>"101101000",
  13831=>"011010110",
  13832=>"001111101",
  13833=>"011010100",
  13834=>"111110110",
  13835=>"010010010",
  13836=>"000010001",
  13837=>"000110001",
  13838=>"001001010",
  13839=>"111010000",
  13840=>"110110001",
  13841=>"000011011",
  13842=>"100100101",
  13843=>"110111100",
  13844=>"001000101",
  13845=>"001110000",
  13846=>"111111100",
  13847=>"010001001",
  13848=>"010110100",
  13849=>"111001010",
  13850=>"000000110",
  13851=>"110001001",
  13852=>"011011110",
  13853=>"001000110",
  13854=>"010100110",
  13855=>"101101110",
  13856=>"111111000",
  13857=>"110001110",
  13858=>"101001111",
  13859=>"010010100",
  13860=>"111100100",
  13861=>"111111111",
  13862=>"111111010",
  13863=>"011100101",
  13864=>"100000101",
  13865=>"011000011",
  13866=>"011100101",
  13867=>"010101001",
  13868=>"000011000",
  13869=>"010010100",
  13870=>"101110000",
  13871=>"111111101",
  13872=>"100111011",
  13873=>"001001010",
  13874=>"001110011",
  13875=>"000100000",
  13876=>"001000010",
  13877=>"111011100",
  13878=>"111100000",
  13879=>"111101011",
  13880=>"111010010",
  13881=>"011101001",
  13882=>"000110011",
  13883=>"100111110",
  13884=>"000011010",
  13885=>"111100000",
  13886=>"111111011",
  13887=>"001111111",
  13888=>"101011010",
  13889=>"011001100",
  13890=>"100011001",
  13891=>"101011001",
  13892=>"000010010",
  13893=>"011110101",
  13894=>"001011101",
  13895=>"101000111",
  13896=>"101000011",
  13897=>"111010011",
  13898=>"111100100",
  13899=>"100111001",
  13900=>"101100101",
  13901=>"101101011",
  13902=>"110010110",
  13903=>"011110010",
  13904=>"111101100",
  13905=>"010111110",
  13906=>"001001101",
  13907=>"011110110",
  13908=>"110110111",
  13909=>"000110110",
  13910=>"110110000",
  13911=>"011110101",
  13912=>"111111010",
  13913=>"001101001",
  13914=>"101111110",
  13915=>"111011110",
  13916=>"111100011",
  13917=>"001110001",
  13918=>"110000111",
  13919=>"010011000",
  13920=>"010010101",
  13921=>"000001000",
  13922=>"110001111",
  13923=>"111101100",
  13924=>"000101011",
  13925=>"100010100",
  13926=>"001111111",
  13927=>"100111100",
  13928=>"001100101",
  13929=>"110000101",
  13930=>"000011100",
  13931=>"000101111",
  13932=>"100100101",
  13933=>"001010101",
  13934=>"010000101",
  13935=>"010010001",
  13936=>"101000001",
  13937=>"000001010",
  13938=>"111011100",
  13939=>"110000011",
  13940=>"000010011",
  13941=>"001100010",
  13942=>"110111010",
  13943=>"100000001",
  13944=>"111010010",
  13945=>"001011110",
  13946=>"100010011",
  13947=>"110111110",
  13948=>"110101110",
  13949=>"000010001",
  13950=>"101100110",
  13951=>"100111001",
  13952=>"000100100",
  13953=>"110011101",
  13954=>"001111110",
  13955=>"011011110",
  13956=>"011100010",
  13957=>"000111001",
  13958=>"111001001",
  13959=>"001000101",
  13960=>"010011111",
  13961=>"111011001",
  13962=>"100111010",
  13963=>"111110101",
  13964=>"110000001",
  13965=>"001110011",
  13966=>"010010100",
  13967=>"100110101",
  13968=>"011110111",
  13969=>"101101011",
  13970=>"101101101",
  13971=>"000101111",
  13972=>"111111000",
  13973=>"111011110",
  13974=>"000100000",
  13975=>"100110101",
  13976=>"111111000",
  13977=>"000100101",
  13978=>"000100000",
  13979=>"010000001",
  13980=>"000000001",
  13981=>"000001100",
  13982=>"110100000",
  13983=>"100011110",
  13984=>"111101110",
  13985=>"111100100",
  13986=>"111111111",
  13987=>"101001100",
  13988=>"111100011",
  13989=>"111100111",
  13990=>"100101100",
  13991=>"000010000",
  13992=>"100011101",
  13993=>"100001110",
  13994=>"001001000",
  13995=>"111000001",
  13996=>"100110000",
  13997=>"010110100",
  13998=>"101000101",
  13999=>"110110100",
  14000=>"110011000",
  14001=>"001110010",
  14002=>"111100111",
  14003=>"001001000",
  14004=>"001111001",
  14005=>"001100010",
  14006=>"010001101",
  14007=>"010100011",
  14008=>"111100010",
  14009=>"000010011",
  14010=>"010100110",
  14011=>"011011000",
  14012=>"111010111",
  14013=>"011110010",
  14014=>"010001011",
  14015=>"000011000",
  14016=>"011010110",
  14017=>"000000010",
  14018=>"001100100",
  14019=>"110011111",
  14020=>"110010011",
  14021=>"001101000",
  14022=>"001000001",
  14023=>"011111010",
  14024=>"100010101",
  14025=>"110111101",
  14026=>"111111100",
  14027=>"000011010",
  14028=>"011100100",
  14029=>"011110111",
  14030=>"001000001",
  14031=>"111000110",
  14032=>"011011101",
  14033=>"110100010",
  14034=>"101010111",
  14035=>"111110001",
  14036=>"011111000",
  14037=>"010100100",
  14038=>"000011101",
  14039=>"111101010",
  14040=>"001001101",
  14041=>"110100000",
  14042=>"001101111",
  14043=>"011101111",
  14044=>"000011111",
  14045=>"100000100",
  14046=>"011011110",
  14047=>"101110110",
  14048=>"011011010",
  14049=>"110000000",
  14050=>"101111101",
  14051=>"111110111",
  14052=>"100100010",
  14053=>"000001001",
  14054=>"011111010",
  14055=>"101000110",
  14056=>"011010000",
  14057=>"111110010",
  14058=>"001010000",
  14059=>"100100100",
  14060=>"001100010",
  14061=>"101100011",
  14062=>"101110110",
  14063=>"001010010",
  14064=>"100001010",
  14065=>"010100110",
  14066=>"111010110",
  14067=>"111010110",
  14068=>"010110111",
  14069=>"000010110",
  14070=>"001001001",
  14071=>"010100110",
  14072=>"001101110",
  14073=>"110011111",
  14074=>"001001011",
  14075=>"001000000",
  14076=>"010111110",
  14077=>"110000000",
  14078=>"010101110",
  14079=>"111010010",
  14080=>"110101010",
  14081=>"011110111",
  14082=>"100111111",
  14083=>"100010010",
  14084=>"011110000",
  14085=>"001100110",
  14086=>"100100001",
  14087=>"010101011",
  14088=>"100101111",
  14089=>"111110110",
  14090=>"111101111",
  14091=>"101111110",
  14092=>"000000111",
  14093=>"010010001",
  14094=>"000011111",
  14095=>"101010000",
  14096=>"000011111",
  14097=>"111011111",
  14098=>"110110010",
  14099=>"011001010",
  14100=>"011111011",
  14101=>"110000111",
  14102=>"101101111",
  14103=>"110100110",
  14104=>"001101010",
  14105=>"100100011",
  14106=>"000000100",
  14107=>"100101101",
  14108=>"110111000",
  14109=>"001110001",
  14110=>"010010111",
  14111=>"011101000",
  14112=>"000011010",
  14113=>"010010001",
  14114=>"111010011",
  14115=>"101000001",
  14116=>"101010101",
  14117=>"111101111",
  14118=>"110110111",
  14119=>"101100000",
  14120=>"011010100",
  14121=>"011110101",
  14122=>"011011000",
  14123=>"000110011",
  14124=>"010011011",
  14125=>"001000011",
  14126=>"001011110",
  14127=>"111111100",
  14128=>"101010001",
  14129=>"011011010",
  14130=>"001100010",
  14131=>"010011001",
  14132=>"100101010",
  14133=>"010101001",
  14134=>"011011100",
  14135=>"010000101",
  14136=>"011111101",
  14137=>"001101111",
  14138=>"011001110",
  14139=>"000111000",
  14140=>"111011010",
  14141=>"010111101",
  14142=>"011011010",
  14143=>"001010000",
  14144=>"010011110",
  14145=>"100100101",
  14146=>"111101010",
  14147=>"110110001",
  14148=>"111111001",
  14149=>"000010111",
  14150=>"000111011",
  14151=>"011011111",
  14152=>"111101001",
  14153=>"100000000",
  14154=>"001011100",
  14155=>"101011101",
  14156=>"001111000",
  14157=>"110101000",
  14158=>"010111000",
  14159=>"111111101",
  14160=>"101101011",
  14161=>"111001100",
  14162=>"010010101",
  14163=>"010001001",
  14164=>"110100011",
  14165=>"101001110",
  14166=>"010100010",
  14167=>"101110011",
  14168=>"010111100",
  14169=>"010100000",
  14170=>"100000010",
  14171=>"001111011",
  14172=>"101011111",
  14173=>"001100110",
  14174=>"000010001",
  14175=>"011101001",
  14176=>"100010111",
  14177=>"111111001",
  14178=>"011010000",
  14179=>"110001111",
  14180=>"100111010",
  14181=>"010111011",
  14182=>"001101101",
  14183=>"101000011",
  14184=>"000000001",
  14185=>"011110100",
  14186=>"001011111",
  14187=>"101010001",
  14188=>"000001101",
  14189=>"010000100",
  14190=>"100010001",
  14191=>"100111110",
  14192=>"110110110",
  14193=>"011101100",
  14194=>"111000111",
  14195=>"011000101",
  14196=>"011000010",
  14197=>"101011011",
  14198=>"001001010",
  14199=>"010010011",
  14200=>"010111111",
  14201=>"001000000",
  14202=>"100100110",
  14203=>"011000111",
  14204=>"001111100",
  14205=>"000011001",
  14206=>"101110100",
  14207=>"010101000",
  14208=>"001101010",
  14209=>"111101010",
  14210=>"000110101",
  14211=>"001101011",
  14212=>"001111011",
  14213=>"011000101",
  14214=>"011101101",
  14215=>"011011001",
  14216=>"000100111",
  14217=>"011001111",
  14218=>"001000110",
  14219=>"110101000",
  14220=>"100000010",
  14221=>"101000000",
  14222=>"111111001",
  14223=>"110110001",
  14224=>"000011000",
  14225=>"011100101",
  14226=>"000001010",
  14227=>"101001111",
  14228=>"010101110",
  14229=>"001011011",
  14230=>"101011100",
  14231=>"111010100",
  14232=>"000101010",
  14233=>"010110111",
  14234=>"111101010",
  14235=>"101011011",
  14236=>"101100100",
  14237=>"111101110",
  14238=>"101110100",
  14239=>"010000110",
  14240=>"010010010",
  14241=>"111111111",
  14242=>"010111100",
  14243=>"110001101",
  14244=>"100101111",
  14245=>"111100110",
  14246=>"000100110",
  14247=>"111001101",
  14248=>"011111011",
  14249=>"000011100",
  14250=>"111000000",
  14251=>"111011010",
  14252=>"110001110",
  14253=>"110110110",
  14254=>"101010110",
  14255=>"010000010",
  14256=>"110110011",
  14257=>"010110011",
  14258=>"101000001",
  14259=>"100110010",
  14260=>"000000001",
  14261=>"010011111",
  14262=>"100010100",
  14263=>"010000101",
  14264=>"001110000",
  14265=>"110100011",
  14266=>"100101110",
  14267=>"001101001",
  14268=>"011101011",
  14269=>"000011011",
  14270=>"011111100",
  14271=>"111000010",
  14272=>"110101100",
  14273=>"101011000",
  14274=>"011110000",
  14275=>"010100000",
  14276=>"101110101",
  14277=>"001111010",
  14278=>"101000111",
  14279=>"001111111",
  14280=>"000011000",
  14281=>"110110011",
  14282=>"001011110",
  14283=>"110100010",
  14284=>"011101000",
  14285=>"110101100",
  14286=>"110001001",
  14287=>"100111000",
  14288=>"101011001",
  14289=>"100110101",
  14290=>"000010111",
  14291=>"100100100",
  14292=>"000010010",
  14293=>"000101011",
  14294=>"000111111",
  14295=>"001111011",
  14296=>"010101010",
  14297=>"010101000",
  14298=>"110001011",
  14299=>"010100010",
  14300=>"010010100",
  14301=>"010100010",
  14302=>"010100010",
  14303=>"001101100",
  14304=>"111000000",
  14305=>"110110110",
  14306=>"110000000",
  14307=>"111010111",
  14308=>"101000000",
  14309=>"000101011",
  14310=>"001011111",
  14311=>"000101000",
  14312=>"101011111",
  14313=>"011001010",
  14314=>"111111010",
  14315=>"101001101",
  14316=>"011000111",
  14317=>"010110001",
  14318=>"000001001",
  14319=>"011101011",
  14320=>"111010011",
  14321=>"100111001",
  14322=>"101001000",
  14323=>"111110010",
  14324=>"001000011",
  14325=>"111110111",
  14326=>"000001011",
  14327=>"110101011",
  14328=>"010010101",
  14329=>"011101111",
  14330=>"111001101",
  14331=>"011000100",
  14332=>"001100111",
  14333=>"010011001",
  14334=>"110000100",
  14335=>"000000000",
  14336=>"000110001",
  14337=>"100101010",
  14338=>"011011110",
  14339=>"100001100",
  14340=>"011110011",
  14341=>"000011110",
  14342=>"101000001",
  14343=>"000100001",
  14344=>"000001110",
  14345=>"111000010",
  14346=>"000000010",
  14347=>"111110101",
  14348=>"101100111",
  14349=>"111001101",
  14350=>"001010001",
  14351=>"100011101",
  14352=>"001010100",
  14353=>"011111001",
  14354=>"110101010",
  14355=>"110110010",
  14356=>"000111011",
  14357=>"101100111",
  14358=>"010111101",
  14359=>"000011001",
  14360=>"000001111",
  14361=>"101011110",
  14362=>"110011110",
  14363=>"100101101",
  14364=>"100011101",
  14365=>"010001110",
  14366=>"100000010",
  14367=>"010001111",
  14368=>"111011001",
  14369=>"001110101",
  14370=>"010000111",
  14371=>"000101001",
  14372=>"111100100",
  14373=>"110101011",
  14374=>"001111101",
  14375=>"110010000",
  14376=>"000000000",
  14377=>"010110111",
  14378=>"110101100",
  14379=>"101001111",
  14380=>"111000010",
  14381=>"110101111",
  14382=>"111101100",
  14383=>"010011001",
  14384=>"000101110",
  14385=>"000011101",
  14386=>"110000011",
  14387=>"110101101",
  14388=>"110001000",
  14389=>"101111010",
  14390=>"000011000",
  14391=>"100110100",
  14392=>"001101000",
  14393=>"001001010",
  14394=>"001010100",
  14395=>"110011111",
  14396=>"001101110",
  14397=>"010010001",
  14398=>"110110110",
  14399=>"010111110",
  14400=>"101101110",
  14401=>"101101110",
  14402=>"011101101",
  14403=>"111100100",
  14404=>"100001101",
  14405=>"101001010",
  14406=>"010000001",
  14407=>"011110100",
  14408=>"000000011",
  14409=>"000010110",
  14410=>"101001110",
  14411=>"100011110",
  14412=>"011100001",
  14413=>"001111111",
  14414=>"111011111",
  14415=>"000000000",
  14416=>"101011001",
  14417=>"010010011",
  14418=>"111100110",
  14419=>"100011101",
  14420=>"101001010",
  14421=>"110001000",
  14422=>"010011111",
  14423=>"101100010",
  14424=>"101000011",
  14425=>"010000011",
  14426=>"111111100",
  14427=>"100001000",
  14428=>"011011101",
  14429=>"101001010",
  14430=>"000011110",
  14431=>"001000000",
  14432=>"100111001",
  14433=>"001010111",
  14434=>"010101011",
  14435=>"110111010",
  14436=>"001100101",
  14437=>"111100110",
  14438=>"001010110",
  14439=>"101111000",
  14440=>"000010100",
  14441=>"000010000",
  14442=>"100000101",
  14443=>"110100010",
  14444=>"001101011",
  14445=>"011100010",
  14446=>"101001101",
  14447=>"100011110",
  14448=>"110100001",
  14449=>"000011000",
  14450=>"000001001",
  14451=>"111011001",
  14452=>"110001010",
  14453=>"101101011",
  14454=>"011011101",
  14455=>"001000001",
  14456=>"100001101",
  14457=>"110010001",
  14458=>"001110100",
  14459=>"011101101",
  14460=>"000001001",
  14461=>"010010011",
  14462=>"010111000",
  14463=>"101100010",
  14464=>"001111111",
  14465=>"010000001",
  14466=>"101101111",
  14467=>"100000101",
  14468=>"011101101",
  14469=>"001000100",
  14470=>"110110111",
  14471=>"001011101",
  14472=>"001000000",
  14473=>"001100110",
  14474=>"011110001",
  14475=>"101011000",
  14476=>"101110111",
  14477=>"100001111",
  14478=>"111001010",
  14479=>"000111011",
  14480=>"101101101",
  14481=>"110010001",
  14482=>"011101010",
  14483=>"000110100",
  14484=>"101010000",
  14485=>"011000111",
  14486=>"100011010",
  14487=>"001111100",
  14488=>"001110000",
  14489=>"100011000",
  14490=>"001010110",
  14491=>"101110110",
  14492=>"100010000",
  14493=>"000000000",
  14494=>"101111111",
  14495=>"101100100",
  14496=>"011000011",
  14497=>"101101101",
  14498=>"000100111",
  14499=>"110110010",
  14500=>"111000010",
  14501=>"010111111",
  14502=>"001100111",
  14503=>"101010001",
  14504=>"001000111",
  14505=>"000010011",
  14506=>"010011011",
  14507=>"111001110",
  14508=>"001011000",
  14509=>"100111001",
  14510=>"100111001",
  14511=>"000001001",
  14512=>"111111101",
  14513=>"101100000",
  14514=>"110100001",
  14515=>"001001010",
  14516=>"110001001",
  14517=>"101101001",
  14518=>"001000010",
  14519=>"110010101",
  14520=>"010010011",
  14521=>"111010011",
  14522=>"101101011",
  14523=>"001111111",
  14524=>"110100111",
  14525=>"001000100",
  14526=>"001001000",
  14527=>"000100001",
  14528=>"001001000",
  14529=>"000011111",
  14530=>"100000010",
  14531=>"111100000",
  14532=>"101100011",
  14533=>"111101001",
  14534=>"010100110",
  14535=>"111011000",
  14536=>"010111110",
  14537=>"001011111",
  14538=>"011011001",
  14539=>"000000001",
  14540=>"011001111",
  14541=>"001001110",
  14542=>"010001101",
  14543=>"010110000",
  14544=>"000010011",
  14545=>"111101011",
  14546=>"100101001",
  14547=>"011100001",
  14548=>"100010011",
  14549=>"000111010",
  14550=>"011100110",
  14551=>"100111001",
  14552=>"111111011",
  14553=>"110110010",
  14554=>"110110101",
  14555=>"000001111",
  14556=>"010010010",
  14557=>"000111110",
  14558=>"100110110",
  14559=>"100010111",
  14560=>"100011000",
  14561=>"100100111",
  14562=>"010001100",
  14563=>"100010110",
  14564=>"011110100",
  14565=>"110101010",
  14566=>"011011111",
  14567=>"111001010",
  14568=>"000100111",
  14569=>"100101100",
  14570=>"100111000",
  14571=>"101111000",
  14572=>"100000100",
  14573=>"111101010",
  14574=>"001010111",
  14575=>"100001011",
  14576=>"001101100",
  14577=>"100100110",
  14578=>"111110010",
  14579=>"111010011",
  14580=>"011001000",
  14581=>"011010001",
  14582=>"111101111",
  14583=>"000100110",
  14584=>"110100111",
  14585=>"100110011",
  14586=>"000110001",
  14587=>"010001100",
  14588=>"110110110",
  14589=>"010111010",
  14590=>"110010111",
  14591=>"000111111",
  14592=>"000110101",
  14593=>"000000100",
  14594=>"111011111",
  14595=>"000011110",
  14596=>"011000110",
  14597=>"110010100",
  14598=>"011010000",
  14599=>"111000100",
  14600=>"100100000",
  14601=>"001110010",
  14602=>"110111001",
  14603=>"010110110",
  14604=>"010101010",
  14605=>"101100110",
  14606=>"110100001",
  14607=>"000110011",
  14608=>"001011110",
  14609=>"000100001",
  14610=>"001010110",
  14611=>"001000101",
  14612=>"011100010",
  14613=>"011101111",
  14614=>"000000000",
  14615=>"001010111",
  14616=>"110010011",
  14617=>"100101110",
  14618=>"011011001",
  14619=>"111010100",
  14620=>"001100011",
  14621=>"111010110",
  14622=>"110100001",
  14623=>"001111111",
  14624=>"000010110",
  14625=>"101000010",
  14626=>"010000011",
  14627=>"100100111",
  14628=>"110011110",
  14629=>"001111110",
  14630=>"011110010",
  14631=>"001101000",
  14632=>"111101111",
  14633=>"000110111",
  14634=>"011111111",
  14635=>"010101011",
  14636=>"011110101",
  14637=>"100111000",
  14638=>"000000010",
  14639=>"110101011",
  14640=>"110101100",
  14641=>"101011010",
  14642=>"011110011",
  14643=>"101101111",
  14644=>"010101110",
  14645=>"110100111",
  14646=>"011010100",
  14647=>"000010111",
  14648=>"100000000",
  14649=>"000011011",
  14650=>"110110011",
  14651=>"010001110",
  14652=>"100011000",
  14653=>"110011010",
  14654=>"010001001",
  14655=>"000001000",
  14656=>"110001001",
  14657=>"001110011",
  14658=>"000011011",
  14659=>"000100010",
  14660=>"101100111",
  14661=>"000011110",
  14662=>"000011001",
  14663=>"000100011",
  14664=>"010101000",
  14665=>"110001101",
  14666=>"001010101",
  14667=>"001100001",
  14668=>"100001110",
  14669=>"100001010",
  14670=>"000000111",
  14671=>"001110101",
  14672=>"110001000",
  14673=>"010000100",
  14674=>"111101101",
  14675=>"000100001",
  14676=>"111010000",
  14677=>"011111000",
  14678=>"000100000",
  14679=>"111100001",
  14680=>"111010010",
  14681=>"010000000",
  14682=>"001101001",
  14683=>"000000110",
  14684=>"001000111",
  14685=>"011100101",
  14686=>"011110100",
  14687=>"100110011",
  14688=>"100111101",
  14689=>"111011111",
  14690=>"101001011",
  14691=>"001000011",
  14692=>"001101001",
  14693=>"100010101",
  14694=>"001010110",
  14695=>"011110101",
  14696=>"111101011",
  14697=>"001110111",
  14698=>"111100110",
  14699=>"011110111",
  14700=>"010001000",
  14701=>"010000100",
  14702=>"000001111",
  14703=>"001110000",
  14704=>"101110011",
  14705=>"000010011",
  14706=>"111010011",
  14707=>"010100001",
  14708=>"101110111",
  14709=>"001000110",
  14710=>"111101111",
  14711=>"110101111",
  14712=>"111001000",
  14713=>"011111101",
  14714=>"011111010",
  14715=>"000011000",
  14716=>"010010101",
  14717=>"010011111",
  14718=>"000100001",
  14719=>"100010110",
  14720=>"110101100",
  14721=>"100011011",
  14722=>"110111110",
  14723=>"000001111",
  14724=>"010100111",
  14725=>"101000111",
  14726=>"111110101",
  14727=>"111110101",
  14728=>"101111011",
  14729=>"000011001",
  14730=>"000100011",
  14731=>"001110000",
  14732=>"100011110",
  14733=>"101110011",
  14734=>"000010001",
  14735=>"111110101",
  14736=>"011011010",
  14737=>"111011011",
  14738=>"001011100",
  14739=>"100100010",
  14740=>"001001001",
  14741=>"010100001",
  14742=>"001001111",
  14743=>"101000110",
  14744=>"101001000",
  14745=>"010001101",
  14746=>"001011011",
  14747=>"010011011",
  14748=>"001001010",
  14749=>"011000101",
  14750=>"001000100",
  14751=>"000000001",
  14752=>"110000100",
  14753=>"111000010",
  14754=>"010110101",
  14755=>"101001111",
  14756=>"001011010",
  14757=>"000101000",
  14758=>"001011000",
  14759=>"101000011",
  14760=>"001111110",
  14761=>"010001000",
  14762=>"110011011",
  14763=>"000100110",
  14764=>"101011000",
  14765=>"101000101",
  14766=>"000011110",
  14767=>"000010001",
  14768=>"001000100",
  14769=>"000101000",
  14770=>"001001111",
  14771=>"001000010",
  14772=>"111111000",
  14773=>"101111110",
  14774=>"000110101",
  14775=>"101010101",
  14776=>"000000000",
  14777=>"011000101",
  14778=>"000110011",
  14779=>"110000110",
  14780=>"001001010",
  14781=>"000100000",
  14782=>"010111000",
  14783=>"001101000",
  14784=>"001010110",
  14785=>"101011001",
  14786=>"000010001",
  14787=>"110111101",
  14788=>"110010010",
  14789=>"001011010",
  14790=>"110110111",
  14791=>"000011001",
  14792=>"001000011",
  14793=>"001010100",
  14794=>"111101101",
  14795=>"111110000",
  14796=>"001011100",
  14797=>"010010110",
  14798=>"111111000",
  14799=>"001010111",
  14800=>"010111011",
  14801=>"010110001",
  14802=>"011110010",
  14803=>"110111110",
  14804=>"000001100",
  14805=>"110110001",
  14806=>"011000110",
  14807=>"000110111",
  14808=>"111111000",
  14809=>"011010100",
  14810=>"011001000",
  14811=>"110001000",
  14812=>"101001101",
  14813=>"101001110",
  14814=>"100110011",
  14815=>"101010001",
  14816=>"111011011",
  14817=>"011001000",
  14818=>"110010010",
  14819=>"111010100",
  14820=>"001101010",
  14821=>"001010001",
  14822=>"111001111",
  14823=>"101101100",
  14824=>"111110100",
  14825=>"010110101",
  14826=>"110010011",
  14827=>"010101001",
  14828=>"010110010",
  14829=>"110000101",
  14830=>"010100010",
  14831=>"101110111",
  14832=>"011010111",
  14833=>"111111111",
  14834=>"111010100",
  14835=>"101101110",
  14836=>"100001000",
  14837=>"101100000",
  14838=>"100101100",
  14839=>"010110100",
  14840=>"000110010",
  14841=>"000000101",
  14842=>"011101100",
  14843=>"010101101",
  14844=>"110110101",
  14845=>"001100101",
  14846=>"011011100",
  14847=>"000100100",
  14848=>"010010111",
  14849=>"010011001",
  14850=>"000000110",
  14851=>"011000100",
  14852=>"000011000",
  14853=>"001111100",
  14854=>"011000001",
  14855=>"101001000",
  14856=>"111110111",
  14857=>"000001011",
  14858=>"100110011",
  14859=>"000101010",
  14860=>"101110010",
  14861=>"001001011",
  14862=>"110001001",
  14863=>"110001100",
  14864=>"010110011",
  14865=>"110000010",
  14866=>"001110001",
  14867=>"101000011",
  14868=>"101011010",
  14869=>"001101001",
  14870=>"110110111",
  14871=>"001111110",
  14872=>"110000100",
  14873=>"111110110",
  14874=>"101000100",
  14875=>"010110111",
  14876=>"011011100",
  14877=>"111010101",
  14878=>"101111100",
  14879=>"100010011",
  14880=>"101001101",
  14881=>"100001010",
  14882=>"110001010",
  14883=>"110010001",
  14884=>"111101101",
  14885=>"001000110",
  14886=>"000110110",
  14887=>"110111100",
  14888=>"001010000",
  14889=>"010100101",
  14890=>"110100001",
  14891=>"010000100",
  14892=>"011110101",
  14893=>"101010111",
  14894=>"011010100",
  14895=>"101000110",
  14896=>"001101111",
  14897=>"111101011",
  14898=>"101001000",
  14899=>"100000110",
  14900=>"101001110",
  14901=>"000000101",
  14902=>"110101001",
  14903=>"100101011",
  14904=>"011001101",
  14905=>"100011110",
  14906=>"011100000",
  14907=>"111100001",
  14908=>"000000110",
  14909=>"000100001",
  14910=>"100101101",
  14911=>"001011100",
  14912=>"111100010",
  14913=>"100011001",
  14914=>"110101100",
  14915=>"000100110",
  14916=>"100010000",
  14917=>"010001011",
  14918=>"101010110",
  14919=>"100010110",
  14920=>"001011011",
  14921=>"100011111",
  14922=>"111111111",
  14923=>"000011000",
  14924=>"000010111",
  14925=>"001001101",
  14926=>"011100010",
  14927=>"000101100",
  14928=>"110101101",
  14929=>"000001100",
  14930=>"001000000",
  14931=>"111100001",
  14932=>"110010110",
  14933=>"111110011",
  14934=>"001110011",
  14935=>"111111100",
  14936=>"100011011",
  14937=>"111101111",
  14938=>"001111100",
  14939=>"001111101",
  14940=>"101101001",
  14941=>"100101011",
  14942=>"110010000",
  14943=>"100001111",
  14944=>"000010110",
  14945=>"010111100",
  14946=>"001000000",
  14947=>"100110010",
  14948=>"100111011",
  14949=>"110110011",
  14950=>"001100001",
  14951=>"001100101",
  14952=>"100100101",
  14953=>"001110100",
  14954=>"011001111",
  14955=>"011100000",
  14956=>"010001000",
  14957=>"001101001",
  14958=>"100101110",
  14959=>"110000111",
  14960=>"010100110",
  14961=>"011111001",
  14962=>"001000110",
  14963=>"111101100",
  14964=>"100001000",
  14965=>"101011010",
  14966=>"011111101",
  14967=>"000100101",
  14968=>"000101110",
  14969=>"010101001",
  14970=>"111111001",
  14971=>"001011010",
  14972=>"001111100",
  14973=>"100000001",
  14974=>"000011111",
  14975=>"000000011",
  14976=>"100111000",
  14977=>"000011110",
  14978=>"000110111",
  14979=>"110110110",
  14980=>"111101011",
  14981=>"110000011",
  14982=>"101001010",
  14983=>"111110011",
  14984=>"011111111",
  14985=>"000111101",
  14986=>"100011111",
  14987=>"001100111",
  14988=>"111011100",
  14989=>"010011111",
  14990=>"110010011",
  14991=>"000000000",
  14992=>"001011101",
  14993=>"110010110",
  14994=>"000101001",
  14995=>"010101101",
  14996=>"000001100",
  14997=>"110010011",
  14998=>"110101111",
  14999=>"000011011",
  15000=>"010101001",
  15001=>"111100110",
  15002=>"100010100",
  15003=>"110101100",
  15004=>"110100010",
  15005=>"001110100",
  15006=>"001111111",
  15007=>"111100000",
  15008=>"011101100",
  15009=>"110000110",
  15010=>"010011110",
  15011=>"111000101",
  15012=>"111110001",
  15013=>"101011010",
  15014=>"101001100",
  15015=>"000110010",
  15016=>"101011011",
  15017=>"110011010",
  15018=>"111010101",
  15019=>"011101111",
  15020=>"000000010",
  15021=>"110011111",
  15022=>"110111010",
  15023=>"000010111",
  15024=>"000001000",
  15025=>"010101101",
  15026=>"000011110",
  15027=>"000110110",
  15028=>"101100011",
  15029=>"011100011",
  15030=>"101010001",
  15031=>"101011110",
  15032=>"111010111",
  15033=>"010000111",
  15034=>"011011001",
  15035=>"110111101",
  15036=>"000000000",
  15037=>"101001011",
  15038=>"011011110",
  15039=>"010000100",
  15040=>"110001000",
  15041=>"101111001",
  15042=>"111001011",
  15043=>"001100001",
  15044=>"100101100",
  15045=>"000000011",
  15046=>"110001010",
  15047=>"100111010",
  15048=>"000011101",
  15049=>"000110000",
  15050=>"000001101",
  15051=>"100101111",
  15052=>"011110000",
  15053=>"111110100",
  15054=>"011000110",
  15055=>"100001000",
  15056=>"011101110",
  15057=>"101000111",
  15058=>"110011111",
  15059=>"011100100",
  15060=>"000101110",
  15061=>"011111000",
  15062=>"110111011",
  15063=>"100111100",
  15064=>"101101100",
  15065=>"010101100",
  15066=>"100110011",
  15067=>"110000011",
  15068=>"000111010",
  15069=>"111111101",
  15070=>"100001101",
  15071=>"011100110",
  15072=>"101111000",
  15073=>"110011000",
  15074=>"010000110",
  15075=>"010000000",
  15076=>"100110001",
  15077=>"101101111",
  15078=>"101110111",
  15079=>"101011011",
  15080=>"000000000",
  15081=>"000011110",
  15082=>"001101000",
  15083=>"010001111",
  15084=>"101100100",
  15085=>"001100101",
  15086=>"110010001",
  15087=>"110010001",
  15088=>"011011010",
  15089=>"110011101",
  15090=>"101111100",
  15091=>"000110111",
  15092=>"100000001",
  15093=>"010110100",
  15094=>"011000001",
  15095=>"011011111",
  15096=>"111100111",
  15097=>"111001110",
  15098=>"010101101",
  15099=>"101000110",
  15100=>"110100100",
  15101=>"001001100",
  15102=>"111001001",
  15103=>"100010010",
  15104=>"100111101",
  15105=>"010000001",
  15106=>"010110111",
  15107=>"100100010",
  15108=>"110100010",
  15109=>"011011110",
  15110=>"010101100",
  15111=>"000100000",
  15112=>"011101011",
  15113=>"001010000",
  15114=>"100011100",
  15115=>"001110100",
  15116=>"111110001",
  15117=>"111100011",
  15118=>"000110010",
  15119=>"111001010",
  15120=>"001010111",
  15121=>"010101100",
  15122=>"110111111",
  15123=>"111011110",
  15124=>"111001011",
  15125=>"010100101",
  15126=>"111110010",
  15127=>"110001101",
  15128=>"111111100",
  15129=>"100111000",
  15130=>"000000000",
  15131=>"000010011",
  15132=>"110011001",
  15133=>"010101110",
  15134=>"000011000",
  15135=>"000000011",
  15136=>"011111101",
  15137=>"101101011",
  15138=>"011100001",
  15139=>"001011011",
  15140=>"110101000",
  15141=>"010110000",
  15142=>"000000101",
  15143=>"101000011",
  15144=>"001001001",
  15145=>"010001101",
  15146=>"110100011",
  15147=>"001101111",
  15148=>"011010000",
  15149=>"000010011",
  15150=>"101100100",
  15151=>"010001011",
  15152=>"010101001",
  15153=>"110000001",
  15154=>"100001010",
  15155=>"111001011",
  15156=>"110001110",
  15157=>"001011000",
  15158=>"001000110",
  15159=>"010000111",
  15160=>"011100000",
  15161=>"100101100",
  15162=>"001010000",
  15163=>"000011000",
  15164=>"110100001",
  15165=>"000000010",
  15166=>"001110100",
  15167=>"100110111",
  15168=>"011001000",
  15169=>"101010011",
  15170=>"001000111",
  15171=>"111001001",
  15172=>"101100110",
  15173=>"111100010",
  15174=>"001001111",
  15175=>"001100101",
  15176=>"100101110",
  15177=>"101100100",
  15178=>"000101100",
  15179=>"101000110",
  15180=>"100100100",
  15181=>"111000101",
  15182=>"010110100",
  15183=>"110011000",
  15184=>"010110110",
  15185=>"101100100",
  15186=>"000011100",
  15187=>"011100101",
  15188=>"101011111",
  15189=>"001100010",
  15190=>"100001100",
  15191=>"000000100",
  15192=>"101000000",
  15193=>"100100110",
  15194=>"100111011",
  15195=>"011010001",
  15196=>"111100010",
  15197=>"011000101",
  15198=>"001100110",
  15199=>"000010000",
  15200=>"010101110",
  15201=>"110101000",
  15202=>"110010100",
  15203=>"101000111",
  15204=>"010100100",
  15205=>"110101111",
  15206=>"111100011",
  15207=>"001100000",
  15208=>"000001101",
  15209=>"010010111",
  15210=>"000101010",
  15211=>"000100011",
  15212=>"010001100",
  15213=>"001101010",
  15214=>"001010010",
  15215=>"101101111",
  15216=>"000100100",
  15217=>"010011000",
  15218=>"000100111",
  15219=>"111000001",
  15220=>"010100100",
  15221=>"111111000",
  15222=>"110011011",
  15223=>"111101001",
  15224=>"000100101",
  15225=>"111100100",
  15226=>"000000010",
  15227=>"111100111",
  15228=>"110111000",
  15229=>"111001100",
  15230=>"111111100",
  15231=>"110111100",
  15232=>"100011101",
  15233=>"100100101",
  15234=>"001011110",
  15235=>"110101010",
  15236=>"000000000",
  15237=>"110000110",
  15238=>"110101111",
  15239=>"001100010",
  15240=>"000110100",
  15241=>"000111100",
  15242=>"001001001",
  15243=>"111101111",
  15244=>"001111110",
  15245=>"011101010",
  15246=>"111111000",
  15247=>"110101110",
  15248=>"000001011",
  15249=>"101010011",
  15250=>"011000000",
  15251=>"010010110",
  15252=>"010010001",
  15253=>"101000011",
  15254=>"101000100",
  15255=>"011001010",
  15256=>"000001110",
  15257=>"000100110",
  15258=>"010010010",
  15259=>"100010100",
  15260=>"111000000",
  15261=>"110111000",
  15262=>"010100010",
  15263=>"110101110",
  15264=>"110010010",
  15265=>"111000011",
  15266=>"111111100",
  15267=>"111111011",
  15268=>"000000100",
  15269=>"111111111",
  15270=>"001110011",
  15271=>"011001000",
  15272=>"000011111",
  15273=>"111001111",
  15274=>"000010110",
  15275=>"101101010",
  15276=>"100001001",
  15277=>"110011101",
  15278=>"100010001",
  15279=>"111001101",
  15280=>"010010000",
  15281=>"011111010",
  15282=>"101101101",
  15283=>"000110001",
  15284=>"110010011",
  15285=>"100001000",
  15286=>"100111111",
  15287=>"010011011",
  15288=>"001000111",
  15289=>"001001001",
  15290=>"100001000",
  15291=>"010110011",
  15292=>"000101100",
  15293=>"110000011",
  15294=>"000000000",
  15295=>"000111111",
  15296=>"111100100",
  15297=>"010110000",
  15298=>"100001111",
  15299=>"101110011",
  15300=>"000111111",
  15301=>"111010110",
  15302=>"111110101",
  15303=>"111010000",
  15304=>"000110101",
  15305=>"101110101",
  15306=>"010001000",
  15307=>"111100111",
  15308=>"111101011",
  15309=>"101101101",
  15310=>"000111001",
  15311=>"101011000",
  15312=>"011101101",
  15313=>"000011010",
  15314=>"011011111",
  15315=>"100101000",
  15316=>"110100000",
  15317=>"111110111",
  15318=>"111000010",
  15319=>"101000001",
  15320=>"101100001",
  15321=>"111111111",
  15322=>"100000111",
  15323=>"011111110",
  15324=>"000110111",
  15325=>"100010100",
  15326=>"011111110",
  15327=>"000100000",
  15328=>"110011001",
  15329=>"001111010",
  15330=>"101010000",
  15331=>"011011110",
  15332=>"010011000",
  15333=>"111101100",
  15334=>"100000010",
  15335=>"011000110",
  15336=>"001110111",
  15337=>"011101011",
  15338=>"111000101",
  15339=>"001110101",
  15340=>"010100010",
  15341=>"000100000",
  15342=>"111101100",
  15343=>"111101010",
  15344=>"000010010",
  15345=>"000110111",
  15346=>"011111101",
  15347=>"110101100",
  15348=>"011011111",
  15349=>"000110101",
  15350=>"100001111",
  15351=>"000111001",
  15352=>"000000100",
  15353=>"101110110",
  15354=>"000011101",
  15355=>"110010001",
  15356=>"010000011",
  15357=>"010111100",
  15358=>"111001001",
  15359=>"000000010",
  15360=>"010001011",
  15361=>"110101110",
  15362=>"011101011",
  15363=>"011111011",
  15364=>"101110111",
  15365=>"100001110",
  15366=>"011001010",
  15367=>"110111000",
  15368=>"101111100",
  15369=>"010100110",
  15370=>"011110011",
  15371=>"001101001",
  15372=>"010000111",
  15373=>"100101101",
  15374=>"001100000",
  15375=>"111001111",
  15376=>"101110010",
  15377=>"100101000",
  15378=>"110101001",
  15379=>"101101011",
  15380=>"011101011",
  15381=>"001000011",
  15382=>"101101111",
  15383=>"011001101",
  15384=>"101000100",
  15385=>"010000000",
  15386=>"011001111",
  15387=>"001000101",
  15388=>"000001010",
  15389=>"101110110",
  15390=>"011010010",
  15391=>"011110001",
  15392=>"100011110",
  15393=>"100010111",
  15394=>"111000100",
  15395=>"100011010",
  15396=>"000101000",
  15397=>"000001000",
  15398=>"110110010",
  15399=>"000111010",
  15400=>"000001111",
  15401=>"110111111",
  15402=>"010001011",
  15403=>"000001110",
  15404=>"000000011",
  15405=>"000011010",
  15406=>"001100100",
  15407=>"010111111",
  15408=>"100011010",
  15409=>"000001001",
  15410=>"110100000",
  15411=>"100010100",
  15412=>"000110001",
  15413=>"110000000",
  15414=>"001110000",
  15415=>"100011011",
  15416=>"111001110",
  15417=>"101111101",
  15418=>"010000001",
  15419=>"011000010",
  15420=>"100000110",
  15421=>"111010111",
  15422=>"010110010",
  15423=>"000111101",
  15424=>"101011001",
  15425=>"000001001",
  15426=>"001111011",
  15427=>"011101111",
  15428=>"000010111",
  15429=>"000011011",
  15430=>"110111011",
  15431=>"000000001",
  15432=>"111101110",
  15433=>"111010100",
  15434=>"101000010",
  15435=>"111111011",
  15436=>"001101110",
  15437=>"001111010",
  15438=>"101111111",
  15439=>"010010000",
  15440=>"100000111",
  15441=>"111001001",
  15442=>"100100110",
  15443=>"011101000",
  15444=>"101101100",
  15445=>"011001000",
  15446=>"010101101",
  15447=>"100101111",
  15448=>"000111110",
  15449=>"101111101",
  15450=>"011000110",
  15451=>"000111011",
  15452=>"001010101",
  15453=>"000001000",
  15454=>"011000100",
  15455=>"001101011",
  15456=>"001000011",
  15457=>"011001011",
  15458=>"101100110",
  15459=>"100011111",
  15460=>"011001111",
  15461=>"101011010",
  15462=>"000100111",
  15463=>"010000101",
  15464=>"000010100",
  15465=>"100111001",
  15466=>"010011011",
  15467=>"011110001",
  15468=>"111010010",
  15469=>"011100100",
  15470=>"111100000",
  15471=>"000000010",
  15472=>"001111001",
  15473=>"100110110",
  15474=>"100000101",
  15475=>"000110101",
  15476=>"001001011",
  15477=>"100100001",
  15478=>"011100101",
  15479=>"010101101",
  15480=>"011101111",
  15481=>"000111101",
  15482=>"000111110",
  15483=>"010000100",
  15484=>"000001000",
  15485=>"001101100",
  15486=>"110001000",
  15487=>"100010010",
  15488=>"101001101",
  15489=>"100011000",
  15490=>"010000100",
  15491=>"011111010",
  15492=>"001011000",
  15493=>"001100110",
  15494=>"110011101",
  15495=>"100011101",
  15496=>"010110001",
  15497=>"110011011",
  15498=>"001000000",
  15499=>"001000001",
  15500=>"010101101",
  15501=>"100001110",
  15502=>"001100001",
  15503=>"100101101",
  15504=>"100010011",
  15505=>"111111110",
  15506=>"000101110",
  15507=>"111101111",
  15508=>"000000001",
  15509=>"101000101",
  15510=>"000011010",
  15511=>"001101010",
  15512=>"111111011",
  15513=>"000110111",
  15514=>"100011101",
  15515=>"000100100",
  15516=>"010011010",
  15517=>"010000111",
  15518=>"000101000",
  15519=>"100110111",
  15520=>"101000001",
  15521=>"000001011",
  15522=>"101111110",
  15523=>"000110100",
  15524=>"000010011",
  15525=>"010001000",
  15526=>"110100100",
  15527=>"010110110",
  15528=>"001000011",
  15529=>"111101111",
  15530=>"010011101",
  15531=>"001101010",
  15532=>"010111100",
  15533=>"010111001",
  15534=>"001110100",
  15535=>"110010011",
  15536=>"011110100",
  15537=>"110010011",
  15538=>"000100101",
  15539=>"110001010",
  15540=>"001100000",
  15541=>"001000000",
  15542=>"001010100",
  15543=>"000001111",
  15544=>"011000001",
  15545=>"010100100",
  15546=>"110011111",
  15547=>"101010010",
  15548=>"101110100",
  15549=>"111111000",
  15550=>"011101010",
  15551=>"110000110",
  15552=>"001101000",
  15553=>"011111111",
  15554=>"110110011",
  15555=>"010111010",
  15556=>"001100011",
  15557=>"101010101",
  15558=>"011110010",
  15559=>"111001001",
  15560=>"111101011",
  15561=>"010010010",
  15562=>"011011101",
  15563=>"100100010",
  15564=>"010111011",
  15565=>"010000001",
  15566=>"011001111",
  15567=>"111000011",
  15568=>"111101011",
  15569=>"000001111",
  15570=>"101000100",
  15571=>"000001111",
  15572=>"001001101",
  15573=>"100001011",
  15574=>"111010111",
  15575=>"010000011",
  15576=>"110000101",
  15577=>"000011001",
  15578=>"100110000",
  15579=>"100101100",
  15580=>"100000110",
  15581=>"110001101",
  15582=>"111001111",
  15583=>"110100101",
  15584=>"001100001",
  15585=>"110011110",
  15586=>"000111101",
  15587=>"011111011",
  15588=>"101101010",
  15589=>"000011110",
  15590=>"011110010",
  15591=>"101000011",
  15592=>"010111101",
  15593=>"110001001",
  15594=>"001111101",
  15595=>"111011101",
  15596=>"010100010",
  15597=>"000111100",
  15598=>"011000011",
  15599=>"001101000",
  15600=>"010110101",
  15601=>"001100011",
  15602=>"000001100",
  15603=>"100110000",
  15604=>"000110101",
  15605=>"101001100",
  15606=>"000111010",
  15607=>"011001001",
  15608=>"011000110",
  15609=>"100111000",
  15610=>"000110110",
  15611=>"101010111",
  15612=>"111000101",
  15613=>"010101011",
  15614=>"011101000",
  15615=>"100101010",
  15616=>"000011011",
  15617=>"011101000",
  15618=>"001100011",
  15619=>"100101000",
  15620=>"111110110",
  15621=>"001001100",
  15622=>"011100100",
  15623=>"001101000",
  15624=>"111010101",
  15625=>"101100111",
  15626=>"110100101",
  15627=>"010101101",
  15628=>"111001011",
  15629=>"111001010",
  15630=>"010101101",
  15631=>"000001100",
  15632=>"111101111",
  15633=>"001000111",
  15634=>"010001011",
  15635=>"110111000",
  15636=>"111111001",
  15637=>"101011100",
  15638=>"010001111",
  15639=>"000100001",
  15640=>"010100100",
  15641=>"110100111",
  15642=>"100011100",
  15643=>"110111010",
  15644=>"010110111",
  15645=>"010100000",
  15646=>"001011111",
  15647=>"000001001",
  15648=>"101000100",
  15649=>"111011001",
  15650=>"110001111",
  15651=>"100111001",
  15652=>"110111111",
  15653=>"001111000",
  15654=>"010110000",
  15655=>"000100111",
  15656=>"101111111",
  15657=>"011111110",
  15658=>"000010100",
  15659=>"111100011",
  15660=>"000010111",
  15661=>"011111010",
  15662=>"010101010",
  15663=>"000010111",
  15664=>"010100111",
  15665=>"101100010",
  15666=>"101111101",
  15667=>"000101001",
  15668=>"011101100",
  15669=>"000010011",
  15670=>"001110100",
  15671=>"111010011",
  15672=>"010000101",
  15673=>"001000011",
  15674=>"011100011",
  15675=>"111110101",
  15676=>"010011010",
  15677=>"010101001",
  15678=>"000100001",
  15679=>"110010100",
  15680=>"111100010",
  15681=>"111100100",
  15682=>"111100000",
  15683=>"011010100",
  15684=>"010000110",
  15685=>"110011011",
  15686=>"010111100",
  15687=>"001110111",
  15688=>"101001001",
  15689=>"010001001",
  15690=>"010100110",
  15691=>"010011111",
  15692=>"111101100",
  15693=>"110101101",
  15694=>"011010101",
  15695=>"111101011",
  15696=>"001001010",
  15697=>"010100100",
  15698=>"100101010",
  15699=>"111011101",
  15700=>"111110011",
  15701=>"100111011",
  15702=>"110110100",
  15703=>"010010011",
  15704=>"000010000",
  15705=>"001101001",
  15706=>"101011100",
  15707=>"110100001",
  15708=>"000111100",
  15709=>"110011011",
  15710=>"100000100",
  15711=>"100111101",
  15712=>"111011100",
  15713=>"101000110",
  15714=>"000111100",
  15715=>"100000101",
  15716=>"011000110",
  15717=>"000000100",
  15718=>"000001101",
  15719=>"011011001",
  15720=>"001101100",
  15721=>"001010000",
  15722=>"010110010",
  15723=>"010000110",
  15724=>"110010010",
  15725=>"000000101",
  15726=>"011010010",
  15727=>"110001010",
  15728=>"110101010",
  15729=>"110011111",
  15730=>"100111000",
  15731=>"000110110",
  15732=>"001001010",
  15733=>"010100000",
  15734=>"010111111",
  15735=>"010101110",
  15736=>"010110111",
  15737=>"011000100",
  15738=>"111010101",
  15739=>"110101010",
  15740=>"010110000",
  15741=>"001101000",
  15742=>"101010111",
  15743=>"011100010",
  15744=>"000011011",
  15745=>"100010100",
  15746=>"110101010",
  15747=>"110100000",
  15748=>"011011111",
  15749=>"011011001",
  15750=>"010100100",
  15751=>"101110111",
  15752=>"111111011",
  15753=>"000110010",
  15754=>"000101100",
  15755=>"011111010",
  15756=>"001000010",
  15757=>"001110000",
  15758=>"101100001",
  15759=>"101101110",
  15760=>"101110001",
  15761=>"010001101",
  15762=>"010100011",
  15763=>"000000011",
  15764=>"010011000",
  15765=>"110100110",
  15766=>"000111111",
  15767=>"011000100",
  15768=>"111111001",
  15769=>"000101111",
  15770=>"111110010",
  15771=>"000011010",
  15772=>"010100100",
  15773=>"000011101",
  15774=>"101000001",
  15775=>"010010001",
  15776=>"101111011",
  15777=>"001100101",
  15778=>"111011011",
  15779=>"000011010",
  15780=>"000101010",
  15781=>"101010100",
  15782=>"111100100",
  15783=>"101101011",
  15784=>"101110010",
  15785=>"111110100",
  15786=>"100111110",
  15787=>"010001001",
  15788=>"000010101",
  15789=>"011100001",
  15790=>"110101001",
  15791=>"101100001",
  15792=>"001110111",
  15793=>"000100101",
  15794=>"000011011",
  15795=>"010001100",
  15796=>"100101110",
  15797=>"010000010",
  15798=>"110111000",
  15799=>"110110000",
  15800=>"000001010",
  15801=>"101000010",
  15802=>"000010010",
  15803=>"111100000",
  15804=>"001000110",
  15805=>"000000010",
  15806=>"101011111",
  15807=>"110101100",
  15808=>"101000010",
  15809=>"110110010",
  15810=>"111101101",
  15811=>"010110011",
  15812=>"010101010",
  15813=>"001110001",
  15814=>"011001010",
  15815=>"101011010",
  15816=>"011101011",
  15817=>"010000100",
  15818=>"000100100",
  15819=>"011011010",
  15820=>"011111011",
  15821=>"011100110",
  15822=>"001000000",
  15823=>"011010100",
  15824=>"010001110",
  15825=>"001010110",
  15826=>"101100101",
  15827=>"100000000",
  15828=>"001000011",
  15829=>"000111011",
  15830=>"010010011",
  15831=>"100101111",
  15832=>"011100010",
  15833=>"111101111",
  15834=>"100101101",
  15835=>"111010011",
  15836=>"010111000",
  15837=>"001101011",
  15838=>"011101111",
  15839=>"110000010",
  15840=>"000001001",
  15841=>"010010010",
  15842=>"100000100",
  15843=>"011001110",
  15844=>"010010100",
  15845=>"101010010",
  15846=>"001010000",
  15847=>"100010100",
  15848=>"110010111",
  15849=>"000011001",
  15850=>"110100000",
  15851=>"010010011",
  15852=>"111111101",
  15853=>"101110010",
  15854=>"111000000",
  15855=>"010001101",
  15856=>"110101110",
  15857=>"101001101",
  15858=>"111100100",
  15859=>"101110111",
  15860=>"010011010",
  15861=>"110100000",
  15862=>"000101011",
  15863=>"101101000",
  15864=>"110011010",
  15865=>"111101011",
  15866=>"100111101",
  15867=>"010011011",
  15868=>"000111010",
  15869=>"011011111",
  15870=>"000111111",
  15871=>"101001101",
  15872=>"000110110",
  15873=>"001000000",
  15874=>"100000101",
  15875=>"010100011",
  15876=>"000011011",
  15877=>"010111111",
  15878=>"001111100",
  15879=>"101010110",
  15880=>"011001110",
  15881=>"111000001",
  15882=>"110001100",
  15883=>"000010000",
  15884=>"100010010",
  15885=>"110010110",
  15886=>"010100100",
  15887=>"010111111",
  15888=>"100010100",
  15889=>"110000010",
  15890=>"111110011",
  15891=>"101000101",
  15892=>"110010010",
  15893=>"000110100",
  15894=>"001001000",
  15895=>"011011010",
  15896=>"000110010",
  15897=>"001010111",
  15898=>"111001101",
  15899=>"000010010",
  15900=>"011011001",
  15901=>"101111111",
  15902=>"011110000",
  15903=>"111011011",
  15904=>"011001111",
  15905=>"111010111",
  15906=>"111111010",
  15907=>"101011000",
  15908=>"100111011",
  15909=>"110111101",
  15910=>"000001011",
  15911=>"001001000",
  15912=>"000001000",
  15913=>"001010110",
  15914=>"001000011",
  15915=>"101000010",
  15916=>"010111000",
  15917=>"011000011",
  15918=>"110001111",
  15919=>"001001010",
  15920=>"110100110",
  15921=>"010101010",
  15922=>"100110100",
  15923=>"001001100",
  15924=>"001101000",
  15925=>"100001011",
  15926=>"000000010",
  15927=>"011011010",
  15928=>"010011111",
  15929=>"011001011",
  15930=>"001100010",
  15931=>"111001100",
  15932=>"111111000",
  15933=>"001101010",
  15934=>"011111011",
  15935=>"000000100",
  15936=>"101101100",
  15937=>"100010010",
  15938=>"101100001",
  15939=>"001001100",
  15940=>"111111011",
  15941=>"010010000",
  15942=>"111001010",
  15943=>"100001000",
  15944=>"100011111",
  15945=>"100011000",
  15946=>"001000000",
  15947=>"000111101",
  15948=>"111010000",
  15949=>"000000011",
  15950=>"011000110",
  15951=>"110101111",
  15952=>"000001010",
  15953=>"101001011",
  15954=>"101000001",
  15955=>"100101100",
  15956=>"010000010",
  15957=>"110000111",
  15958=>"001101001",
  15959=>"010011000",
  15960=>"101011000",
  15961=>"010101011",
  15962=>"001101010",
  15963=>"100111101",
  15964=>"001101101",
  15965=>"111110111",
  15966=>"001100000",
  15967=>"000100101",
  15968=>"000111010",
  15969=>"100100111",
  15970=>"101000010",
  15971=>"111001001",
  15972=>"000110011",
  15973=>"000100101",
  15974=>"110001111",
  15975=>"000011011",
  15976=>"101011100",
  15977=>"001110010",
  15978=>"110110110",
  15979=>"011100011",
  15980=>"000010100",
  15981=>"100001000",
  15982=>"101110001",
  15983=>"111100111",
  15984=>"110000001",
  15985=>"011100000",
  15986=>"111101001",
  15987=>"010001010",
  15988=>"101111000",
  15989=>"100110110",
  15990=>"101000111",
  15991=>"100111100",
  15992=>"010001101",
  15993=>"110000101",
  15994=>"111111000",
  15995=>"111110001",
  15996=>"111000010",
  15997=>"011111010",
  15998=>"100000001",
  15999=>"001010011",
  16000=>"000101001",
  16001=>"110010010",
  16002=>"011001011",
  16003=>"001011100",
  16004=>"010111101",
  16005=>"100010101",
  16006=>"101111001",
  16007=>"010000110",
  16008=>"000101000",
  16009=>"000111100",
  16010=>"011111000",
  16011=>"011100110",
  16012=>"011001101",
  16013=>"010110000",
  16014=>"000011011",
  16015=>"001101010",
  16016=>"010010000",
  16017=>"011010000",
  16018=>"101000000",
  16019=>"110010010",
  16020=>"100001011",
  16021=>"111001011",
  16022=>"011110000",
  16023=>"111000011",
  16024=>"011110111",
  16025=>"110000110",
  16026=>"100111101",
  16027=>"111110011",
  16028=>"000110000",
  16029=>"011001001",
  16030=>"010110000",
  16031=>"101001001",
  16032=>"000000010",
  16033=>"000100001",
  16034=>"000001011",
  16035=>"011000000",
  16036=>"100100001",
  16037=>"001010101",
  16038=>"000101101",
  16039=>"110000001",
  16040=>"111011010",
  16041=>"001001000",
  16042=>"011011010",
  16043=>"101110001",
  16044=>"001110110",
  16045=>"101101100",
  16046=>"110100101",
  16047=>"111100101",
  16048=>"011100000",
  16049=>"001010000",
  16050=>"110000010",
  16051=>"010000010",
  16052=>"010111110",
  16053=>"100001110",
  16054=>"101001011",
  16055=>"010100001",
  16056=>"111110011",
  16057=>"010010011",
  16058=>"100010011",
  16059=>"111000000",
  16060=>"110011101",
  16061=>"000111010",
  16062=>"111010010",
  16063=>"010111111",
  16064=>"011111011",
  16065=>"101011101",
  16066=>"000111111",
  16067=>"100100001",
  16068=>"010111010",
  16069=>"100001111",
  16070=>"110000011",
  16071=>"000000111",
  16072=>"100110000",
  16073=>"001010010",
  16074=>"100010111",
  16075=>"111001101",
  16076=>"110100101",
  16077=>"110000010",
  16078=>"110110000",
  16079=>"110110111",
  16080=>"111000101",
  16081=>"011010001",
  16082=>"001101011",
  16083=>"000111010",
  16084=>"000000010",
  16085=>"101100101",
  16086=>"100011100",
  16087=>"100011110",
  16088=>"001101011",
  16089=>"001111000",
  16090=>"101010111",
  16091=>"001010101",
  16092=>"000101000",
  16093=>"111011110",
  16094=>"111111101",
  16095=>"010001110",
  16096=>"001101011",
  16097=>"100000100",
  16098=>"111011101",
  16099=>"011101111",
  16100=>"110111101",
  16101=>"000111011",
  16102=>"110010010",
  16103=>"010111011",
  16104=>"110110111",
  16105=>"101111110",
  16106=>"010111001",
  16107=>"011010000",
  16108=>"001011000",
  16109=>"000101110",
  16110=>"100111010",
  16111=>"010000100",
  16112=>"011000000",
  16113=>"000000010",
  16114=>"111101100",
  16115=>"011110111",
  16116=>"101000010",
  16117=>"101011101",
  16118=>"101101000",
  16119=>"010000011",
  16120=>"011001001",
  16121=>"100110111",
  16122=>"110011011",
  16123=>"001100000",
  16124=>"010110110",
  16125=>"001001000",
  16126=>"000101011",
  16127=>"000000000",
  16128=>"000100101",
  16129=>"111011110",
  16130=>"101011110",
  16131=>"000010010",
  16132=>"001111100",
  16133=>"010000001",
  16134=>"010111101",
  16135=>"110011000",
  16136=>"111010000",
  16137=>"011111000",
  16138=>"111110010",
  16139=>"100101011",
  16140=>"011100100",
  16141=>"100100101",
  16142=>"101110000",
  16143=>"111111110",
  16144=>"010001100",
  16145=>"110100100",
  16146=>"111000000",
  16147=>"110111001",
  16148=>"010010011",
  16149=>"101000101",
  16150=>"011011011",
  16151=>"111111001",
  16152=>"010111110",
  16153=>"111010001",
  16154=>"100100010",
  16155=>"001100001",
  16156=>"110001110",
  16157=>"110111000",
  16158=>"001011010",
  16159=>"010110111",
  16160=>"010111111",
  16161=>"110101111",
  16162=>"111101010",
  16163=>"110001110",
  16164=>"011001011",
  16165=>"100110000",
  16166=>"110001100",
  16167=>"110001011",
  16168=>"011110001",
  16169=>"000000110",
  16170=>"111101100",
  16171=>"100011010",
  16172=>"001000011",
  16173=>"111100101",
  16174=>"111110010",
  16175=>"100000101",
  16176=>"110001000",
  16177=>"100010111",
  16178=>"011001010",
  16179=>"111001110",
  16180=>"101011011",
  16181=>"110101010",
  16182=>"110101011",
  16183=>"001000001",
  16184=>"011010001",
  16185=>"000010111",
  16186=>"000001110",
  16187=>"001101100",
  16188=>"010110000",
  16189=>"111010101",
  16190=>"111101000",
  16191=>"011110010",
  16192=>"111110110",
  16193=>"111000110",
  16194=>"001010100",
  16195=>"001011111",
  16196=>"010001111",
  16197=>"001110001",
  16198=>"001000000",
  16199=>"001111000",
  16200=>"111100101",
  16201=>"101011010",
  16202=>"101111110",
  16203=>"010010001",
  16204=>"011001010",
  16205=>"010011101",
  16206=>"111111001",
  16207=>"010101100",
  16208=>"001111000",
  16209=>"111001101",
  16210=>"011010011",
  16211=>"101111111",
  16212=>"111010111",
  16213=>"010101101",
  16214=>"011100101",
  16215=>"001110010",
  16216=>"011001111",
  16217=>"000001110",
  16218=>"111101011",
  16219=>"110101110",
  16220=>"101111111",
  16221=>"101010110",
  16222=>"010111010",
  16223=>"001010011",
  16224=>"110101000",
  16225=>"000110001",
  16226=>"010111111",
  16227=>"110111110",
  16228=>"001100011",
  16229=>"011100011",
  16230=>"011010100",
  16231=>"000110010",
  16232=>"110011011",
  16233=>"011000101",
  16234=>"110100111",
  16235=>"100101000",
  16236=>"100000001",
  16237=>"011000010",
  16238=>"000010011",
  16239=>"010010101",
  16240=>"101110010",
  16241=>"101100101",
  16242=>"011001000",
  16243=>"011011111",
  16244=>"011010011",
  16245=>"011010111",
  16246=>"001011001",
  16247=>"000101011",
  16248=>"111110011",
  16249=>"000110100",
  16250=>"100001010",
  16251=>"001110110",
  16252=>"111010110",
  16253=>"000010010",
  16254=>"100100100",
  16255=>"111110101",
  16256=>"001011000",
  16257=>"111100101",
  16258=>"111111111",
  16259=>"110111100",
  16260=>"000111101",
  16261=>"100000011",
  16262=>"001110101",
  16263=>"001010110",
  16264=>"101001110",
  16265=>"100100010",
  16266=>"011000110",
  16267=>"011111011",
  16268=>"000001111",
  16269=>"101001001",
  16270=>"000111101",
  16271=>"111011101",
  16272=>"111001110",
  16273=>"000110001",
  16274=>"010011001",
  16275=>"001010111",
  16276=>"110111111",
  16277=>"100110100",
  16278=>"010100110",
  16279=>"110101111",
  16280=>"100011101",
  16281=>"111101001",
  16282=>"110010011",
  16283=>"101111101",
  16284=>"111011110",
  16285=>"011111110",
  16286=>"011110101",
  16287=>"100010011",
  16288=>"110010111",
  16289=>"111000001",
  16290=>"010010011",
  16291=>"111010110",
  16292=>"111001001",
  16293=>"100110111",
  16294=>"100110011",
  16295=>"101111110",
  16296=>"011100010",
  16297=>"001100110",
  16298=>"010110101",
  16299=>"101100100",
  16300=>"000000011",
  16301=>"011110011",
  16302=>"010001001",
  16303=>"011111110",
  16304=>"000001001",
  16305=>"101000111",
  16306=>"011101110",
  16307=>"100100101",
  16308=>"111111110",
  16309=>"100111011",
  16310=>"001101111",
  16311=>"010011010",
  16312=>"110010110",
  16313=>"001100110",
  16314=>"110001001",
  16315=>"101001011",
  16316=>"111101101",
  16317=>"100000000",
  16318=>"000101100",
  16319=>"000000100",
  16320=>"111010110",
  16321=>"110110000",
  16322=>"000010000",
  16323=>"000010111",
  16324=>"100100100",
  16325=>"000011011",
  16326=>"001111000",
  16327=>"100001110",
  16328=>"010011110",
  16329=>"110000110",
  16330=>"000111100",
  16331=>"101111011",
  16332=>"111110011",
  16333=>"011111001",
  16334=>"000000001",
  16335=>"101001001",
  16336=>"100001101",
  16337=>"110111111",
  16338=>"011011010",
  16339=>"100010101",
  16340=>"001000011",
  16341=>"100110010",
  16342=>"010010000",
  16343=>"111111001",
  16344=>"000000111",
  16345=>"001100100",
  16346=>"111000000",
  16347=>"011001110",
  16348=>"110111011",
  16349=>"000100111",
  16350=>"010001000",
  16351=>"100010110",
  16352=>"011001011",
  16353=>"100011000",
  16354=>"000000110",
  16355=>"000011110",
  16356=>"101100100",
  16357=>"000110001",
  16358=>"111010001",
  16359=>"001011011",
  16360=>"110001101",
  16361=>"010010110",
  16362=>"000100010",
  16363=>"011001111",
  16364=>"100010010",
  16365=>"111100111",
  16366=>"000110011",
  16367=>"100111000",
  16368=>"010100110",
  16369=>"000010101",
  16370=>"011101001",
  16371=>"101000100",
  16372=>"111010000",
  16373=>"110101011",
  16374=>"001110001",
  16375=>"011011110",
  16376=>"010000110",
  16377=>"000100110",
  16378=>"100011111",
  16379=>"010111000",
  16380=>"010000000",
  16381=>"011010111",
  16382=>"111000010",
  16383=>"110001000",
  16384=>"010000111",
  16385=>"101110010",
  16386=>"011011111",
  16387=>"010011001",
  16388=>"110110000",
  16389=>"010010001",
  16390=>"011101011",
  16391=>"111111100",
  16392=>"010110101",
  16393=>"100000001",
  16394=>"111011100",
  16395=>"010001100",
  16396=>"111100111",
  16397=>"010001110",
  16398=>"000010100",
  16399=>"101101100",
  16400=>"101111111",
  16401=>"010011101",
  16402=>"101011111",
  16403=>"010110000",
  16404=>"101110000",
  16405=>"001111101",
  16406=>"011011000",
  16407=>"110100100",
  16408=>"111110110",
  16409=>"101110001",
  16410=>"111100001",
  16411=>"110101100",
  16412=>"000101010",
  16413=>"110110110",
  16414=>"011100111",
  16415=>"110100010",
  16416=>"000101011",
  16417=>"010110010",
  16418=>"110000100",
  16419=>"100011111",
  16420=>"010100011",
  16421=>"011011110",
  16422=>"111101011",
  16423=>"110000100",
  16424=>"101111010",
  16425=>"000101000",
  16426=>"101111010",
  16427=>"000111111",
  16428=>"011010110",
  16429=>"010111100",
  16430=>"011010110",
  16431=>"000100111",
  16432=>"000111000",
  16433=>"011110000",
  16434=>"111101010",
  16435=>"111110111",
  16436=>"110101111",
  16437=>"100001101",
  16438=>"111100010",
  16439=>"010011000",
  16440=>"011010010",
  16441=>"111100110",
  16442=>"101010011",
  16443=>"110000111",
  16444=>"111100101",
  16445=>"110010011",
  16446=>"100000101",
  16447=>"000001000",
  16448=>"010100101",
  16449=>"000001101",
  16450=>"111001110",
  16451=>"110100011",
  16452=>"111011100",
  16453=>"101101000",
  16454=>"001111111",
  16455=>"101011011",
  16456=>"110000010",
  16457=>"001011001",
  16458=>"010001010",
  16459=>"101001111",
  16460=>"101000111",
  16461=>"101100011",
  16462=>"111111110",
  16463=>"000001001",
  16464=>"011100100",
  16465=>"010001000",
  16466=>"100110000",
  16467=>"111110011",
  16468=>"110100101",
  16469=>"111101000",
  16470=>"001010010",
  16471=>"110101111",
  16472=>"110110100",
  16473=>"001010001",
  16474=>"001100010",
  16475=>"010111011",
  16476=>"011010001",
  16477=>"000011001",
  16478=>"100100101",
  16479=>"110010000",
  16480=>"000011011",
  16481=>"101011110",
  16482=>"100101010",
  16483=>"000001101",
  16484=>"110001101",
  16485=>"101000001",
  16486=>"101000000",
  16487=>"000010010",
  16488=>"001000101",
  16489=>"111101111",
  16490=>"100010010",
  16491=>"110011101",
  16492=>"011101001",
  16493=>"110010101",
  16494=>"111000110",
  16495=>"000111101",
  16496=>"111111111",
  16497=>"001101101",
  16498=>"000011000",
  16499=>"111000001",
  16500=>"010100100",
  16501=>"010010110",
  16502=>"001011000",
  16503=>"010010010",
  16504=>"110010000",
  16505=>"100010010",
  16506=>"110101001",
  16507=>"011110100",
  16508=>"111010000",
  16509=>"100110111",
  16510=>"100111101",
  16511=>"111100010",
  16512=>"110010010",
  16513=>"100010111",
  16514=>"000101100",
  16515=>"111111011",
  16516=>"110000010",
  16517=>"101110011",
  16518=>"101110111",
  16519=>"000111110",
  16520=>"001110000",
  16521=>"101011011",
  16522=>"101001111",
  16523=>"011101110",
  16524=>"111001101",
  16525=>"110001010",
  16526=>"100110000",
  16527=>"001101001",
  16528=>"111100111",
  16529=>"010111110",
  16530=>"111001111",
  16531=>"010011000",
  16532=>"100111011",
  16533=>"100001110",
  16534=>"101111011",
  16535=>"101101111",
  16536=>"101010000",
  16537=>"001011000",
  16538=>"000111000",
  16539=>"110001000",
  16540=>"110000000",
  16541=>"111111111",
  16542=>"110111001",
  16543=>"100101001",
  16544=>"100000110",
  16545=>"111000001",
  16546=>"100001101",
  16547=>"000001111",
  16548=>"001000001",
  16549=>"001000110",
  16550=>"000111101",
  16551=>"010001111",
  16552=>"000111000",
  16553=>"111011010",
  16554=>"111110011",
  16555=>"011111000",
  16556=>"011000011",
  16557=>"100001111",
  16558=>"000101101",
  16559=>"000111011",
  16560=>"010110010",
  16561=>"010110010",
  16562=>"000111110",
  16563=>"010010111",
  16564=>"111100000",
  16565=>"111011101",
  16566=>"000111101",
  16567=>"100110100",
  16568=>"111101001",
  16569=>"010001000",
  16570=>"010110011",
  16571=>"010011011",
  16572=>"110100110",
  16573=>"111000000",
  16574=>"001010010",
  16575=>"101101001",
  16576=>"001011101",
  16577=>"101010011",
  16578=>"000001111",
  16579=>"001001111",
  16580=>"101001011",
  16581=>"000111001",
  16582=>"001011011",
  16583=>"010001010",
  16584=>"111111011",
  16585=>"110000000",
  16586=>"111101101",
  16587=>"100101011",
  16588=>"010110000",
  16589=>"100011000",
  16590=>"100011101",
  16591=>"110001100",
  16592=>"111110000",
  16593=>"101001111",
  16594=>"111010000",
  16595=>"010111111",
  16596=>"011110010",
  16597=>"000101000",
  16598=>"000010101",
  16599=>"001000010",
  16600=>"101000010",
  16601=>"100010111",
  16602=>"101111100",
  16603=>"110100111",
  16604=>"111110001",
  16605=>"110011001",
  16606=>"001011110",
  16607=>"000101000",
  16608=>"111000111",
  16609=>"000110110",
  16610=>"100111001",
  16611=>"000001001",
  16612=>"100011100",
  16613=>"101010001",
  16614=>"100010000",
  16615=>"000011000",
  16616=>"110000011",
  16617=>"110001110",
  16618=>"101100001",
  16619=>"111100111",
  16620=>"010011001",
  16621=>"011011111",
  16622=>"110111100",
  16623=>"100100110",
  16624=>"101101011",
  16625=>"110101100",
  16626=>"100001010",
  16627=>"111111101",
  16628=>"001100010",
  16629=>"100001111",
  16630=>"001001100",
  16631=>"100000000",
  16632=>"000100101",
  16633=>"011100000",
  16634=>"110000010",
  16635=>"000101011",
  16636=>"000011000",
  16637=>"100100000",
  16638=>"010011011",
  16639=>"100111101",
  16640=>"111101101",
  16641=>"100000010",
  16642=>"101011010",
  16643=>"101010110",
  16644=>"001111010",
  16645=>"001000011",
  16646=>"000011000",
  16647=>"110010111",
  16648=>"000111011",
  16649=>"101111101",
  16650=>"010110100",
  16651=>"001010101",
  16652=>"001011000",
  16653=>"101111110",
  16654=>"111111110",
  16655=>"011111001",
  16656=>"111000110",
  16657=>"001101001",
  16658=>"110010011",
  16659=>"111110100",
  16660=>"101100100",
  16661=>"000000010",
  16662=>"110011101",
  16663=>"011010110",
  16664=>"011001101",
  16665=>"111100101",
  16666=>"100000011",
  16667=>"111111111",
  16668=>"111000111",
  16669=>"000001111",
  16670=>"111000111",
  16671=>"001001011",
  16672=>"110011001",
  16673=>"000010110",
  16674=>"100010001",
  16675=>"111001111",
  16676=>"111010111",
  16677=>"111100110",
  16678=>"111110010",
  16679=>"000001110",
  16680=>"000001111",
  16681=>"111101110",
  16682=>"001000100",
  16683=>"001100110",
  16684=>"110110000",
  16685=>"100100101",
  16686=>"101010011",
  16687=>"010101010",
  16688=>"010101100",
  16689=>"011111111",
  16690=>"000101100",
  16691=>"001000101",
  16692=>"110101110",
  16693=>"110011100",
  16694=>"100101011",
  16695=>"101111011",
  16696=>"101010000",
  16697=>"010100101",
  16698=>"000011000",
  16699=>"100100010",
  16700=>"111100001",
  16701=>"111100101",
  16702=>"110111001",
  16703=>"111111000",
  16704=>"110010100",
  16705=>"001010010",
  16706=>"111111100",
  16707=>"011011110",
  16708=>"111001000",
  16709=>"100101010",
  16710=>"000011000",
  16711=>"110000110",
  16712=>"010101101",
  16713=>"101111001",
  16714=>"101100000",
  16715=>"011101110",
  16716=>"010111110",
  16717=>"011000100",
  16718=>"111110101",
  16719=>"010000001",
  16720=>"010101000",
  16721=>"101110001",
  16722=>"111010101",
  16723=>"011001011",
  16724=>"000111000",
  16725=>"000001001",
  16726=>"111011011",
  16727=>"101101011",
  16728=>"100010111",
  16729=>"000001000",
  16730=>"100100001",
  16731=>"001101110",
  16732=>"000011010",
  16733=>"100001000",
  16734=>"011000111",
  16735=>"110001001",
  16736=>"001101001",
  16737=>"111111011",
  16738=>"100010010",
  16739=>"000010100",
  16740=>"111101011",
  16741=>"100010010",
  16742=>"100110011",
  16743=>"110101100",
  16744=>"001010011",
  16745=>"100111110",
  16746=>"000111000",
  16747=>"110000110",
  16748=>"010101000",
  16749=>"011001011",
  16750=>"010111011",
  16751=>"010111010",
  16752=>"000000000",
  16753=>"000110001",
  16754=>"101111001",
  16755=>"110111001",
  16756=>"001111100",
  16757=>"111101100",
  16758=>"000100000",
  16759=>"000111101",
  16760=>"011010101",
  16761=>"011010110",
  16762=>"100100000",
  16763=>"010111110",
  16764=>"100100010",
  16765=>"100110010",
  16766=>"100101101",
  16767=>"111100001",
  16768=>"111011001",
  16769=>"001101010",
  16770=>"000110011",
  16771=>"100100001",
  16772=>"001010111",
  16773=>"110111000",
  16774=>"001011101",
  16775=>"111100001",
  16776=>"101011011",
  16777=>"101001011",
  16778=>"001110101",
  16779=>"001010010",
  16780=>"100110111",
  16781=>"100110001",
  16782=>"110000010",
  16783=>"000011010",
  16784=>"000100101",
  16785=>"000010011",
  16786=>"010100001",
  16787=>"010101100",
  16788=>"000000000",
  16789=>"100011001",
  16790=>"111111001",
  16791=>"011001101",
  16792=>"000010110",
  16793=>"100111100",
  16794=>"010110000",
  16795=>"111110001",
  16796=>"101011001",
  16797=>"101111000",
  16798=>"000100000",
  16799=>"111011011",
  16800=>"111101101",
  16801=>"101011110",
  16802=>"000001011",
  16803=>"111010100",
  16804=>"101000110",
  16805=>"111001110",
  16806=>"010111111",
  16807=>"100101001",
  16808=>"100110011",
  16809=>"001011010",
  16810=>"000110000",
  16811=>"101010101",
  16812=>"011010100",
  16813=>"111111111",
  16814=>"110010010",
  16815=>"111010010",
  16816=>"010001100",
  16817=>"100001000",
  16818=>"110101001",
  16819=>"100010000",
  16820=>"111000000",
  16821=>"111111011",
  16822=>"000111001",
  16823=>"011001000",
  16824=>"001110111",
  16825=>"000100010",
  16826=>"000100110",
  16827=>"000110110",
  16828=>"111100101",
  16829=>"010110001",
  16830=>"110100101",
  16831=>"010010000",
  16832=>"010001100",
  16833=>"000010001",
  16834=>"000001011",
  16835=>"111101111",
  16836=>"001010100",
  16837=>"001111000",
  16838=>"011111111",
  16839=>"111001001",
  16840=>"001100001",
  16841=>"001010000",
  16842=>"100110110",
  16843=>"111011101",
  16844=>"100110000",
  16845=>"101001000",
  16846=>"000010001",
  16847=>"111110110",
  16848=>"100101001",
  16849=>"000010000",
  16850=>"010100100",
  16851=>"001010100",
  16852=>"000110100",
  16853=>"001110001",
  16854=>"110000011",
  16855=>"000111010",
  16856=>"000010011",
  16857=>"010011110",
  16858=>"011000011",
  16859=>"110011100",
  16860=>"001011000",
  16861=>"010011111",
  16862=>"011111111",
  16863=>"000110011",
  16864=>"101101010",
  16865=>"010010000",
  16866=>"001000000",
  16867=>"010010011",
  16868=>"110000001",
  16869=>"110111011",
  16870=>"101100110",
  16871=>"010100000",
  16872=>"010001011",
  16873=>"110001000",
  16874=>"101001111",
  16875=>"110000000",
  16876=>"001001100",
  16877=>"111111111",
  16878=>"011000101",
  16879=>"111100100",
  16880=>"010100100",
  16881=>"110111111",
  16882=>"101100001",
  16883=>"111101001",
  16884=>"110000010",
  16885=>"010010101",
  16886=>"000110001",
  16887=>"111101101",
  16888=>"111010000",
  16889=>"100001101",
  16890=>"110110111",
  16891=>"100101001",
  16892=>"000100000",
  16893=>"111110000",
  16894=>"000111101",
  16895=>"010101111",
  16896=>"111011100",
  16897=>"010010100",
  16898=>"111011001",
  16899=>"111000000",
  16900=>"101010111",
  16901=>"110010000",
  16902=>"101010101",
  16903=>"010011110",
  16904=>"101110000",
  16905=>"000110000",
  16906=>"010101000",
  16907=>"010010010",
  16908=>"010011011",
  16909=>"101101001",
  16910=>"111101000",
  16911=>"001100010",
  16912=>"101010010",
  16913=>"011111110",
  16914=>"100111001",
  16915=>"101101000",
  16916=>"111111110",
  16917=>"101000110",
  16918=>"110001101",
  16919=>"000101101",
  16920=>"000001011",
  16921=>"110110010",
  16922=>"111100000",
  16923=>"011110101",
  16924=>"111111000",
  16925=>"010110100",
  16926=>"100010111",
  16927=>"000110010",
  16928=>"111000011",
  16929=>"111010010",
  16930=>"011100100",
  16931=>"001001110",
  16932=>"000111111",
  16933=>"000000010",
  16934=>"101111010",
  16935=>"111000011",
  16936=>"111110000",
  16937=>"001110001",
  16938=>"011010100",
  16939=>"110001010",
  16940=>"010001110",
  16941=>"000111001",
  16942=>"100100110",
  16943=>"001111011",
  16944=>"111010011",
  16945=>"001001001",
  16946=>"000011010",
  16947=>"110010000",
  16948=>"001100100",
  16949=>"001011000",
  16950=>"001011110",
  16951=>"011001010",
  16952=>"010001001",
  16953=>"111111010",
  16954=>"110110100",
  16955=>"100111001",
  16956=>"001100101",
  16957=>"111101101",
  16958=>"101010011",
  16959=>"100100111",
  16960=>"010001110",
  16961=>"100101001",
  16962=>"001001011",
  16963=>"011110000",
  16964=>"111100010",
  16965=>"111000101",
  16966=>"100011100",
  16967=>"010111000",
  16968=>"111001011",
  16969=>"000110000",
  16970=>"011101010",
  16971=>"000000000",
  16972=>"010101000",
  16973=>"100100000",
  16974=>"110111001",
  16975=>"001000001",
  16976=>"001010001",
  16977=>"000100001",
  16978=>"101110010",
  16979=>"101001111",
  16980=>"001110101",
  16981=>"000100010",
  16982=>"100010111",
  16983=>"110111000",
  16984=>"111100010",
  16985=>"110111110",
  16986=>"101000111",
  16987=>"100111110",
  16988=>"110001101",
  16989=>"010011000",
  16990=>"001010000",
  16991=>"001000101",
  16992=>"000001111",
  16993=>"110110010",
  16994=>"101101011",
  16995=>"100010111",
  16996=>"000001111",
  16997=>"111101001",
  16998=>"001111110",
  16999=>"001110010",
  17000=>"000101000",
  17001=>"010011110",
  17002=>"011011001",
  17003=>"111000000",
  17004=>"111101100",
  17005=>"000100101",
  17006=>"110000000",
  17007=>"111010101",
  17008=>"000100001",
  17009=>"011000010",
  17010=>"001111000",
  17011=>"101111110",
  17012=>"111101101",
  17013=>"000111000",
  17014=>"011101010",
  17015=>"101100011",
  17016=>"111010000",
  17017=>"111100011",
  17018=>"011101000",
  17019=>"100011000",
  17020=>"001001001",
  17021=>"000001110",
  17022=>"110100110",
  17023=>"111010101",
  17024=>"110100111",
  17025=>"110100100",
  17026=>"101111010",
  17027=>"000011010",
  17028=>"000001001",
  17029=>"100100100",
  17030=>"011010110",
  17031=>"111111110",
  17032=>"100110111",
  17033=>"011010001",
  17034=>"000110101",
  17035=>"001010100",
  17036=>"101100000",
  17037=>"110110111",
  17038=>"111111111",
  17039=>"011111001",
  17040=>"000001111",
  17041=>"000001100",
  17042=>"000101110",
  17043=>"000011101",
  17044=>"000100000",
  17045=>"110011010",
  17046=>"000010101",
  17047=>"111001101",
  17048=>"001101000",
  17049=>"010110000",
  17050=>"001010011",
  17051=>"001010011",
  17052=>"111001001",
  17053=>"110110111",
  17054=>"100111101",
  17055=>"110010011",
  17056=>"001110110",
  17057=>"000100011",
  17058=>"101000111",
  17059=>"101101001",
  17060=>"101101111",
  17061=>"101000011",
  17062=>"000000111",
  17063=>"101000101",
  17064=>"000100011",
  17065=>"111001001",
  17066=>"101001110",
  17067=>"011101010",
  17068=>"011011111",
  17069=>"011100000",
  17070=>"111000110",
  17071=>"100111011",
  17072=>"101001001",
  17073=>"010100000",
  17074=>"000110111",
  17075=>"110010010",
  17076=>"101000001",
  17077=>"000001110",
  17078=>"010100011",
  17079=>"111111000",
  17080=>"100010101",
  17081=>"011110011",
  17082=>"010111010",
  17083=>"101011010",
  17084=>"010110011",
  17085=>"011000010",
  17086=>"000100001",
  17087=>"111010000",
  17088=>"110100000",
  17089=>"110100111",
  17090=>"010111001",
  17091=>"110000011",
  17092=>"000010010",
  17093=>"101101101",
  17094=>"011010111",
  17095=>"011101011",
  17096=>"110111111",
  17097=>"011001110",
  17098=>"110010010",
  17099=>"001111101",
  17100=>"000100000",
  17101=>"001011100",
  17102=>"101101000",
  17103=>"110001100",
  17104=>"011011000",
  17105=>"010111011",
  17106=>"111111110",
  17107=>"110101011",
  17108=>"111001011",
  17109=>"001111111",
  17110=>"100100000",
  17111=>"001101000",
  17112=>"001101100",
  17113=>"111000111",
  17114=>"101000110",
  17115=>"110011110",
  17116=>"001010010",
  17117=>"111001000",
  17118=>"000010010",
  17119=>"001000110",
  17120=>"100101111",
  17121=>"110110101",
  17122=>"100001110",
  17123=>"011011111",
  17124=>"000000110",
  17125=>"111101110",
  17126=>"111010100",
  17127=>"100001010",
  17128=>"000001010",
  17129=>"011110100",
  17130=>"010011100",
  17131=>"010010000",
  17132=>"010010110",
  17133=>"000000001",
  17134=>"000011001",
  17135=>"110011100",
  17136=>"100101100",
  17137=>"111111100",
  17138=>"110011101",
  17139=>"111101100",
  17140=>"000000000",
  17141=>"111111111",
  17142=>"010011111",
  17143=>"101110011",
  17144=>"111011010",
  17145=>"011111000",
  17146=>"101001101",
  17147=>"111100110",
  17148=>"001101000",
  17149=>"100001010",
  17150=>"111000110",
  17151=>"000001011",
  17152=>"110110001",
  17153=>"001100010",
  17154=>"000110111",
  17155=>"000110110",
  17156=>"010001010",
  17157=>"000100010",
  17158=>"001100001",
  17159=>"001010101",
  17160=>"001111101",
  17161=>"000011010",
  17162=>"011000101",
  17163=>"011010001",
  17164=>"001010111",
  17165=>"100100110",
  17166=>"110110110",
  17167=>"101100001",
  17168=>"100111111",
  17169=>"100100010",
  17170=>"111110100",
  17171=>"011100011",
  17172=>"010111011",
  17173=>"010010011",
  17174=>"001111101",
  17175=>"111010100",
  17176=>"001101001",
  17177=>"111000100",
  17178=>"111011100",
  17179=>"101111001",
  17180=>"111001100",
  17181=>"000111101",
  17182=>"100110000",
  17183=>"110011010",
  17184=>"000111000",
  17185=>"101001110",
  17186=>"010011000",
  17187=>"001011000",
  17188=>"000101011",
  17189=>"011011000",
  17190=>"000101010",
  17191=>"010100011",
  17192=>"010011111",
  17193=>"011010111",
  17194=>"011001111",
  17195=>"011100100",
  17196=>"111111000",
  17197=>"001101110",
  17198=>"100100110",
  17199=>"010010001",
  17200=>"101011110",
  17201=>"111110001",
  17202=>"101100000",
  17203=>"010001000",
  17204=>"100110111",
  17205=>"111100000",
  17206=>"101010101",
  17207=>"111001111",
  17208=>"110111100",
  17209=>"111100000",
  17210=>"110101010",
  17211=>"110001011",
  17212=>"000011001",
  17213=>"110001100",
  17214=>"111100001",
  17215=>"000011000",
  17216=>"101101101",
  17217=>"010001111",
  17218=>"111010101",
  17219=>"111100110",
  17220=>"001010111",
  17221=>"010111101",
  17222=>"001000000",
  17223=>"000111000",
  17224=>"111111101",
  17225=>"001000001",
  17226=>"000000101",
  17227=>"001100100",
  17228=>"110001011",
  17229=>"000110101",
  17230=>"010011001",
  17231=>"010101000",
  17232=>"101101101",
  17233=>"001000001",
  17234=>"100111100",
  17235=>"111101010",
  17236=>"011111011",
  17237=>"100100001",
  17238=>"010011101",
  17239=>"101011000",
  17240=>"110110100",
  17241=>"010000011",
  17242=>"011010111",
  17243=>"010111111",
  17244=>"111100011",
  17245=>"000000101",
  17246=>"111001000",
  17247=>"000111000",
  17248=>"000110000",
  17249=>"101011111",
  17250=>"000011110",
  17251=>"100000000",
  17252=>"100110011",
  17253=>"101010001",
  17254=>"011110010",
  17255=>"011101110",
  17256=>"111101001",
  17257=>"111000001",
  17258=>"011111000",
  17259=>"001000010",
  17260=>"101010110",
  17261=>"110101111",
  17262=>"101101100",
  17263=>"001101111",
  17264=>"110110000",
  17265=>"100000000",
  17266=>"011010111",
  17267=>"100001101",
  17268=>"111000000",
  17269=>"110011111",
  17270=>"000101100",
  17271=>"100000000",
  17272=>"011110111",
  17273=>"111100011",
  17274=>"000010000",
  17275=>"101011100",
  17276=>"000011000",
  17277=>"011100101",
  17278=>"010000100",
  17279=>"000010010",
  17280=>"000010010",
  17281=>"101000010",
  17282=>"100111000",
  17283=>"010101011",
  17284=>"100001110",
  17285=>"001010011",
  17286=>"110001011",
  17287=>"011101000",
  17288=>"101100110",
  17289=>"111111111",
  17290=>"000000001",
  17291=>"101111110",
  17292=>"011010100",
  17293=>"000010101",
  17294=>"101011011",
  17295=>"010011010",
  17296=>"100101101",
  17297=>"111011001",
  17298=>"111000000",
  17299=>"110000100",
  17300=>"111110001",
  17301=>"010000111",
  17302=>"111101011",
  17303=>"011011101",
  17304=>"001011011",
  17305=>"111110011",
  17306=>"000100011",
  17307=>"011110111",
  17308=>"001111001",
  17309=>"111101011",
  17310=>"101010010",
  17311=>"001000101",
  17312=>"101111001",
  17313=>"111111001",
  17314=>"000011000",
  17315=>"111011001",
  17316=>"101010100",
  17317=>"110001110",
  17318=>"000101100",
  17319=>"110000010",
  17320=>"111000000",
  17321=>"111011111",
  17322=>"010001010",
  17323=>"110001100",
  17324=>"011100010",
  17325=>"001010011",
  17326=>"000110110",
  17327=>"111111110",
  17328=>"011000001",
  17329=>"110010100",
  17330=>"101010110",
  17331=>"011001011",
  17332=>"001010010",
  17333=>"101110111",
  17334=>"010000010",
  17335=>"110000001",
  17336=>"001101011",
  17337=>"111010100",
  17338=>"101000010",
  17339=>"111101000",
  17340=>"111101011",
  17341=>"000101001",
  17342=>"110000100",
  17343=>"101100110",
  17344=>"000111101",
  17345=>"000001000",
  17346=>"001111001",
  17347=>"111111000",
  17348=>"010001001",
  17349=>"100000101",
  17350=>"010101101",
  17351=>"000101110",
  17352=>"000000001",
  17353=>"010010011",
  17354=>"010011011",
  17355=>"001111110",
  17356=>"101010110",
  17357=>"100101101",
  17358=>"010110100",
  17359=>"111100011",
  17360=>"010110001",
  17361=>"111100101",
  17362=>"001011000",
  17363=>"011001011",
  17364=>"100111011",
  17365=>"000111101",
  17366=>"110101100",
  17367=>"001000000",
  17368=>"001110011",
  17369=>"100001010",
  17370=>"000001000",
  17371=>"111110011",
  17372=>"110101001",
  17373=>"111110000",
  17374=>"000111010",
  17375=>"001100001",
  17376=>"101000000",
  17377=>"000111101",
  17378=>"000011010",
  17379=>"110000010",
  17380=>"101101000",
  17381=>"111000011",
  17382=>"000001110",
  17383=>"010110010",
  17384=>"110000000",
  17385=>"010101011",
  17386=>"101001010",
  17387=>"010111000",
  17388=>"000100000",
  17389=>"101111100",
  17390=>"001101110",
  17391=>"011111111",
  17392=>"100010110",
  17393=>"100110111",
  17394=>"001011111",
  17395=>"110100111",
  17396=>"111100000",
  17397=>"000000100",
  17398=>"111011000",
  17399=>"011010100",
  17400=>"011110001",
  17401=>"001001000",
  17402=>"111001000",
  17403=>"001001011",
  17404=>"100000011",
  17405=>"000000000",
  17406=>"000010001",
  17407=>"001101010",
  17408=>"011000010",
  17409=>"000101011",
  17410=>"111010111",
  17411=>"000010100",
  17412=>"110100001",
  17413=>"001010110",
  17414=>"110100011",
  17415=>"101010011",
  17416=>"111111111",
  17417=>"110010001",
  17418=>"110011011",
  17419=>"100101110",
  17420=>"100000101",
  17421=>"100010001",
  17422=>"101001110",
  17423=>"011100011",
  17424=>"001000000",
  17425=>"110010100",
  17426=>"111100101",
  17427=>"000111100",
  17428=>"111101111",
  17429=>"001101001",
  17430=>"101000110",
  17431=>"000001010",
  17432=>"110011001",
  17433=>"010011011",
  17434=>"100111001",
  17435=>"001010101",
  17436=>"000001110",
  17437=>"111010111",
  17438=>"111011101",
  17439=>"110101101",
  17440=>"110011111",
  17441=>"100111011",
  17442=>"011000001",
  17443=>"111011010",
  17444=>"011110000",
  17445=>"110111110",
  17446=>"001101100",
  17447=>"010001000",
  17448=>"101100110",
  17449=>"000110010",
  17450=>"000010101",
  17451=>"011100100",
  17452=>"110000000",
  17453=>"011110000",
  17454=>"110000001",
  17455=>"011110010",
  17456=>"111100010",
  17457=>"110100010",
  17458=>"010000101",
  17459=>"000110100",
  17460=>"101110010",
  17461=>"011100101",
  17462=>"001110101",
  17463=>"100011111",
  17464=>"100000100",
  17465=>"001100110",
  17466=>"110110011",
  17467=>"001001100",
  17468=>"110001101",
  17469=>"011100101",
  17470=>"111101011",
  17471=>"001001100",
  17472=>"000001100",
  17473=>"001100000",
  17474=>"010001101",
  17475=>"110101101",
  17476=>"101001110",
  17477=>"000001110",
  17478=>"010000000",
  17479=>"101111101",
  17480=>"001000011",
  17481=>"011000100",
  17482=>"001001000",
  17483=>"011011100",
  17484=>"011011101",
  17485=>"100101011",
  17486=>"010101001",
  17487=>"100001101",
  17488=>"111110110",
  17489=>"001101111",
  17490=>"000100100",
  17491=>"101011011",
  17492=>"000000010",
  17493=>"000001001",
  17494=>"001110110",
  17495=>"101001010",
  17496=>"000110111",
  17497=>"101001001",
  17498=>"001011000",
  17499=>"000010101",
  17500=>"100010011",
  17501=>"000000110",
  17502=>"000101010",
  17503=>"001101011",
  17504=>"101111010",
  17505=>"100000101",
  17506=>"000101101",
  17507=>"000011100",
  17508=>"111100000",
  17509=>"001111010",
  17510=>"111000001",
  17511=>"100011110",
  17512=>"110001101",
  17513=>"100111001",
  17514=>"000000001",
  17515=>"011010100",
  17516=>"101011101",
  17517=>"011110101",
  17518=>"001111111",
  17519=>"101000101",
  17520=>"010010010",
  17521=>"000100101",
  17522=>"011010100",
  17523=>"101110111",
  17524=>"010101000",
  17525=>"110000100",
  17526=>"000100010",
  17527=>"001011110",
  17528=>"100110011",
  17529=>"011010101",
  17530=>"011100010",
  17531=>"110100001",
  17532=>"000010101",
  17533=>"110110001",
  17534=>"100001010",
  17535=>"011001101",
  17536=>"100110101",
  17537=>"010111010",
  17538=>"011011101",
  17539=>"111000111",
  17540=>"110011100",
  17541=>"110101101",
  17542=>"001101101",
  17543=>"111001100",
  17544=>"100010010",
  17545=>"000011111",
  17546=>"100000000",
  17547=>"111001001",
  17548=>"101100001",
  17549=>"000010000",
  17550=>"110011011",
  17551=>"101110101",
  17552=>"100011011",
  17553=>"000011011",
  17554=>"111111110",
  17555=>"101110101",
  17556=>"110010010",
  17557=>"001110000",
  17558=>"101010100",
  17559=>"000110001",
  17560=>"111101001",
  17561=>"101001011",
  17562=>"000011101",
  17563=>"101100011",
  17564=>"001001100",
  17565=>"111000011",
  17566=>"010001011",
  17567=>"100011111",
  17568=>"111110111",
  17569=>"101100011",
  17570=>"010001111",
  17571=>"000000111",
  17572=>"100101001",
  17573=>"000000010",
  17574=>"001110010",
  17575=>"110011000",
  17576=>"111101011",
  17577=>"111111101",
  17578=>"111100011",
  17579=>"110011001",
  17580=>"000001110",
  17581=>"001010110",
  17582=>"001111001",
  17583=>"111011100",
  17584=>"111000100",
  17585=>"101100101",
  17586=>"100011111",
  17587=>"101110101",
  17588=>"110100101",
  17589=>"101101101",
  17590=>"000001111",
  17591=>"001000101",
  17592=>"110010000",
  17593=>"001010100",
  17594=>"010001111",
  17595=>"001001011",
  17596=>"110001001",
  17597=>"111001001",
  17598=>"100101111",
  17599=>"011100100",
  17600=>"011101001",
  17601=>"110101000",
  17602=>"010010110",
  17603=>"111010011",
  17604=>"100101000",
  17605=>"100101011",
  17606=>"001000101",
  17607=>"011101100",
  17608=>"100111010",
  17609=>"010100111",
  17610=>"110111110",
  17611=>"010001111",
  17612=>"100001000",
  17613=>"110000011",
  17614=>"000011011",
  17615=>"101000000",
  17616=>"010000110",
  17617=>"000101000",
  17618=>"010001011",
  17619=>"000001110",
  17620=>"110010110",
  17621=>"110001000",
  17622=>"101100101",
  17623=>"100010001",
  17624=>"011001101",
  17625=>"111000000",
  17626=>"001001101",
  17627=>"101111110",
  17628=>"011111100",
  17629=>"101110000",
  17630=>"000101110",
  17631=>"110101001",
  17632=>"100001110",
  17633=>"100000000",
  17634=>"101001010",
  17635=>"000101101",
  17636=>"001000101",
  17637=>"111111010",
  17638=>"010011001",
  17639=>"110101010",
  17640=>"000110111",
  17641=>"100000101",
  17642=>"000000000",
  17643=>"001011111",
  17644=>"110100110",
  17645=>"101100001",
  17646=>"011000000",
  17647=>"001101010",
  17648=>"011111001",
  17649=>"100011000",
  17650=>"000001001",
  17651=>"100101100",
  17652=>"111000011",
  17653=>"011000101",
  17654=>"010110011",
  17655=>"100001000",
  17656=>"011011011",
  17657=>"110010111",
  17658=>"111110100",
  17659=>"100110111",
  17660=>"001110101",
  17661=>"000100101",
  17662=>"100110011",
  17663=>"101001111",
  17664=>"111110011",
  17665=>"100000010",
  17666=>"111100100",
  17667=>"100000100",
  17668=>"011000010",
  17669=>"000111010",
  17670=>"000111100",
  17671=>"000001011",
  17672=>"011101010",
  17673=>"010000110",
  17674=>"111111101",
  17675=>"100010110",
  17676=>"001100100",
  17677=>"000011101",
  17678=>"011101001",
  17679=>"000110011",
  17680=>"100010011",
  17681=>"011111011",
  17682=>"001111000",
  17683=>"111000111",
  17684=>"011000011",
  17685=>"110100010",
  17686=>"110001010",
  17687=>"001111111",
  17688=>"010010100",
  17689=>"010000111",
  17690=>"111100111",
  17691=>"011011101",
  17692=>"001101010",
  17693=>"001110011",
  17694=>"100010010",
  17695=>"010110111",
  17696=>"000010100",
  17697=>"010100010",
  17698=>"101100100",
  17699=>"011010011",
  17700=>"110000001",
  17701=>"000101110",
  17702=>"010001001",
  17703=>"011100011",
  17704=>"011000100",
  17705=>"110101101",
  17706=>"110011110",
  17707=>"011010101",
  17708=>"001011001",
  17709=>"000111000",
  17710=>"101110000",
  17711=>"000000111",
  17712=>"010100110",
  17713=>"110110100",
  17714=>"011110110",
  17715=>"111010011",
  17716=>"111101000",
  17717=>"011001001",
  17718=>"011010001",
  17719=>"011110111",
  17720=>"011101000",
  17721=>"001010100",
  17722=>"100100001",
  17723=>"111000001",
  17724=>"000011110",
  17725=>"000001100",
  17726=>"100100000",
  17727=>"111010011",
  17728=>"111010011",
  17729=>"111111000",
  17730=>"001110000",
  17731=>"100001000",
  17732=>"110101010",
  17733=>"100000000",
  17734=>"110100111",
  17735=>"000110001",
  17736=>"101011000",
  17737=>"000101101",
  17738=>"101011000",
  17739=>"111111101",
  17740=>"111101110",
  17741=>"111101100",
  17742=>"001100110",
  17743=>"001100010",
  17744=>"010100010",
  17745=>"011000010",
  17746=>"001100001",
  17747=>"110000011",
  17748=>"110110100",
  17749=>"110100011",
  17750=>"101001101",
  17751=>"100000010",
  17752=>"110010000",
  17753=>"000101111",
  17754=>"001110100",
  17755=>"110100001",
  17756=>"101110101",
  17757=>"110010000",
  17758=>"000101000",
  17759=>"000111010",
  17760=>"011101111",
  17761=>"010000011",
  17762=>"111100000",
  17763=>"011111111",
  17764=>"000010010",
  17765=>"111011011",
  17766=>"000001001",
  17767=>"000001110",
  17768=>"110100111",
  17769=>"111001101",
  17770=>"001011100",
  17771=>"011011010",
  17772=>"010001100",
  17773=>"100011111",
  17774=>"001101100",
  17775=>"011100101",
  17776=>"100100000",
  17777=>"100011101",
  17778=>"000110100",
  17779=>"001110110",
  17780=>"011001110",
  17781=>"001000111",
  17782=>"100110001",
  17783=>"010100011",
  17784=>"000110110",
  17785=>"001010001",
  17786=>"011011100",
  17787=>"111111010",
  17788=>"011000101",
  17789=>"000110111",
  17790=>"101101011",
  17791=>"010101101",
  17792=>"100101111",
  17793=>"000111100",
  17794=>"010000010",
  17795=>"000111001",
  17796=>"100000000",
  17797=>"010000010",
  17798=>"011000110",
  17799=>"010010010",
  17800=>"100100110",
  17801=>"011000011",
  17802=>"100110011",
  17803=>"010101000",
  17804=>"001101001",
  17805=>"111101000",
  17806=>"010101000",
  17807=>"011101110",
  17808=>"001001111",
  17809=>"000000001",
  17810=>"010111011",
  17811=>"001011100",
  17812=>"010010110",
  17813=>"111101111",
  17814=>"001101011",
  17815=>"000110100",
  17816=>"011111101",
  17817=>"111111001",
  17818=>"010101011",
  17819=>"001110001",
  17820=>"000100010",
  17821=>"000000100",
  17822=>"100011110",
  17823=>"001001001",
  17824=>"111100000",
  17825=>"101101100",
  17826=>"010100001",
  17827=>"001001010",
  17828=>"001000110",
  17829=>"111111001",
  17830=>"110010011",
  17831=>"111001101",
  17832=>"011111001",
  17833=>"101111100",
  17834=>"000110010",
  17835=>"010001010",
  17836=>"010111001",
  17837=>"101001111",
  17838=>"101001101",
  17839=>"010010101",
  17840=>"110010101",
  17841=>"110111011",
  17842=>"100001011",
  17843=>"111101001",
  17844=>"101001110",
  17845=>"111101100",
  17846=>"100011000",
  17847=>"001101100",
  17848=>"011110011",
  17849=>"000100101",
  17850=>"110101001",
  17851=>"010001111",
  17852=>"011110111",
  17853=>"100101010",
  17854=>"000001010",
  17855=>"111110010",
  17856=>"111001001",
  17857=>"000001100",
  17858=>"000000110",
  17859=>"111100110",
  17860=>"010101001",
  17861=>"000111010",
  17862=>"010001001",
  17863=>"000010110",
  17864=>"001010000",
  17865=>"000000110",
  17866=>"011110001",
  17867=>"110101100",
  17868=>"110010000",
  17869=>"100111111",
  17870=>"101011111",
  17871=>"011011110",
  17872=>"111000101",
  17873=>"010101010",
  17874=>"001110101",
  17875=>"010110000",
  17876=>"011110111",
  17877=>"101000110",
  17878=>"000110000",
  17879=>"010111011",
  17880=>"100010110",
  17881=>"110011100",
  17882=>"011000111",
  17883=>"101110010",
  17884=>"110010011",
  17885=>"000110000",
  17886=>"010000100",
  17887=>"001111110",
  17888=>"111010101",
  17889=>"100011001",
  17890=>"110110100",
  17891=>"000010001",
  17892=>"000010000",
  17893=>"000000001",
  17894=>"101111101",
  17895=>"100010000",
  17896=>"100011110",
  17897=>"000111110",
  17898=>"000000010",
  17899=>"110111010",
  17900=>"110011000",
  17901=>"000001011",
  17902=>"110000000",
  17903=>"000101001",
  17904=>"110111100",
  17905=>"100101010",
  17906=>"000101100",
  17907=>"001001011",
  17908=>"111000001",
  17909=>"101111000",
  17910=>"010110011",
  17911=>"100000000",
  17912=>"111101000",
  17913=>"111110100",
  17914=>"000101101",
  17915=>"100111111",
  17916=>"011111110",
  17917=>"001010110",
  17918=>"000011111",
  17919=>"100011011",
  17920=>"101100010",
  17921=>"101011100",
  17922=>"110110111",
  17923=>"100011010",
  17924=>"101110010",
  17925=>"000100101",
  17926=>"101111001",
  17927=>"100111100",
  17928=>"100011001",
  17929=>"100110010",
  17930=>"010000000",
  17931=>"110010011",
  17932=>"000110010",
  17933=>"001100101",
  17934=>"000000100",
  17935=>"111110110",
  17936=>"011001010",
  17937=>"111101011",
  17938=>"000001010",
  17939=>"111100001",
  17940=>"110100101",
  17941=>"000101110",
  17942=>"100110100",
  17943=>"001101100",
  17944=>"100111000",
  17945=>"100010011",
  17946=>"010101001",
  17947=>"110110101",
  17948=>"000001000",
  17949=>"110001111",
  17950=>"001100001",
  17951=>"010110011",
  17952=>"101011001",
  17953=>"111111010",
  17954=>"010001010",
  17955=>"000010110",
  17956=>"011111011",
  17957=>"000110110",
  17958=>"010100000",
  17959=>"100010000",
  17960=>"100101010",
  17961=>"011101000",
  17962=>"101000011",
  17963=>"110010001",
  17964=>"100110111",
  17965=>"001110100",
  17966=>"110000110",
  17967=>"110101001",
  17968=>"111011100",
  17969=>"101001010",
  17970=>"101000111",
  17971=>"001001010",
  17972=>"110000000",
  17973=>"110110001",
  17974=>"110010000",
  17975=>"101100101",
  17976=>"011101110",
  17977=>"101111100",
  17978=>"011001011",
  17979=>"110001010",
  17980=>"101000011",
  17981=>"100011101",
  17982=>"111101111",
  17983=>"010010001",
  17984=>"000001100",
  17985=>"001010000",
  17986=>"010101011",
  17987=>"101011010",
  17988=>"000010110",
  17989=>"000100100",
  17990=>"100000011",
  17991=>"001000001",
  17992=>"101111000",
  17993=>"000011101",
  17994=>"001101001",
  17995=>"010010110",
  17996=>"111101110",
  17997=>"100101000",
  17998=>"111000011",
  17999=>"100100001",
  18000=>"000101010",
  18001=>"110100011",
  18002=>"111111011",
  18003=>"010001011",
  18004=>"101011010",
  18005=>"011101110",
  18006=>"000100001",
  18007=>"111111011",
  18008=>"100000101",
  18009=>"100000000",
  18010=>"001001110",
  18011=>"010010111",
  18012=>"110010010",
  18013=>"101101101",
  18014=>"000100110",
  18015=>"000101110",
  18016=>"010001100",
  18017=>"010001111",
  18018=>"100101101",
  18019=>"100000110",
  18020=>"011000000",
  18021=>"010101001",
  18022=>"000111010",
  18023=>"001111011",
  18024=>"000100101",
  18025=>"011010011",
  18026=>"011010001",
  18027=>"000111000",
  18028=>"100000110",
  18029=>"001000110",
  18030=>"010001010",
  18031=>"010001111",
  18032=>"110001100",
  18033=>"000010111",
  18034=>"001101001",
  18035=>"100100001",
  18036=>"110101000",
  18037=>"110100011",
  18038=>"110110011",
  18039=>"000101011",
  18040=>"101001111",
  18041=>"000111000",
  18042=>"011110010",
  18043=>"111010000",
  18044=>"111101001",
  18045=>"100111011",
  18046=>"100110101",
  18047=>"110110100",
  18048=>"000110110",
  18049=>"001101011",
  18050=>"000011000",
  18051=>"100111001",
  18052=>"111100100",
  18053=>"111000110",
  18054=>"101001110",
  18055=>"010010101",
  18056=>"101011001",
  18057=>"010001001",
  18058=>"001111110",
  18059=>"011111110",
  18060=>"101010111",
  18061=>"011010101",
  18062=>"101101100",
  18063=>"000110011",
  18064=>"011110000",
  18065=>"101011010",
  18066=>"110111110",
  18067=>"010001111",
  18068=>"001000010",
  18069=>"100100010",
  18070=>"111111011",
  18071=>"111010100",
  18072=>"100100000",
  18073=>"111101101",
  18074=>"001000000",
  18075=>"000111110",
  18076=>"110101000",
  18077=>"010101101",
  18078=>"100010000",
  18079=>"000001110",
  18080=>"100111011",
  18081=>"100101101",
  18082=>"111111101",
  18083=>"101110001",
  18084=>"110100001",
  18085=>"001110000",
  18086=>"011011100",
  18087=>"100000000",
  18088=>"011111110",
  18089=>"100000000",
  18090=>"101000111",
  18091=>"011110001",
  18092=>"011111000",
  18093=>"110011111",
  18094=>"010001100",
  18095=>"001111001",
  18096=>"001000111",
  18097=>"100011010",
  18098=>"010001000",
  18099=>"001110101",
  18100=>"010111001",
  18101=>"011010101",
  18102=>"000001101",
  18103=>"011110010",
  18104=>"000100001",
  18105=>"011110001",
  18106=>"010101111",
  18107=>"001001111",
  18108=>"111101101",
  18109=>"101101101",
  18110=>"110111001",
  18111=>"011011010",
  18112=>"010110011",
  18113=>"111001000",
  18114=>"101111101",
  18115=>"011011101",
  18116=>"101000011",
  18117=>"111000101",
  18118=>"110111101",
  18119=>"001000111",
  18120=>"111111001",
  18121=>"100111011",
  18122=>"001111111",
  18123=>"100000000",
  18124=>"100111110",
  18125=>"011010001",
  18126=>"101110000",
  18127=>"111101011",
  18128=>"110100100",
  18129=>"111111100",
  18130=>"001010010",
  18131=>"110001111",
  18132=>"010000101",
  18133=>"010100010",
  18134=>"111101111",
  18135=>"011110111",
  18136=>"011111101",
  18137=>"010110100",
  18138=>"000110001",
  18139=>"111010010",
  18140=>"001101010",
  18141=>"000000100",
  18142=>"100100100",
  18143=>"110001101",
  18144=>"011010101",
  18145=>"010010100",
  18146=>"000001000",
  18147=>"001110100",
  18148=>"110100011",
  18149=>"000101110",
  18150=>"100101000",
  18151=>"110110010",
  18152=>"011011101",
  18153=>"001111110",
  18154=>"110110010",
  18155=>"011011000",
  18156=>"111101110",
  18157=>"011111100",
  18158=>"101100110",
  18159=>"000100001",
  18160=>"111100100",
  18161=>"001011010",
  18162=>"110101111",
  18163=>"100111011",
  18164=>"000111111",
  18165=>"100011110",
  18166=>"000100010",
  18167=>"111100101",
  18168=>"011101001",
  18169=>"111010010",
  18170=>"011111101",
  18171=>"111101011",
  18172=>"110010111",
  18173=>"001011001",
  18174=>"110111101",
  18175=>"001010010",
  18176=>"110110000",
  18177=>"100101110",
  18178=>"101110001",
  18179=>"111011000",
  18180=>"110101001",
  18181=>"010101101",
  18182=>"101001000",
  18183=>"111010111",
  18184=>"011111000",
  18185=>"010101111",
  18186=>"100111110",
  18187=>"101001000",
  18188=>"100001100",
  18189=>"000010010",
  18190=>"000010001",
  18191=>"000100111",
  18192=>"100010100",
  18193=>"101011111",
  18194=>"101100101",
  18195=>"000011011",
  18196=>"111100111",
  18197=>"001110110",
  18198=>"111011011",
  18199=>"100000010",
  18200=>"010010110",
  18201=>"111001010",
  18202=>"100011001",
  18203=>"000010010",
  18204=>"100101111",
  18205=>"011101111",
  18206=>"001100001",
  18207=>"101110110",
  18208=>"011001010",
  18209=>"110000010",
  18210=>"011001101",
  18211=>"111101111",
  18212=>"010000110",
  18213=>"110111000",
  18214=>"010000011",
  18215=>"100010101",
  18216=>"010101101",
  18217=>"011101110",
  18218=>"011101111",
  18219=>"111011101",
  18220=>"000011001",
  18221=>"100101011",
  18222=>"111010100",
  18223=>"111101011",
  18224=>"110000001",
  18225=>"011111111",
  18226=>"100000110",
  18227=>"100011010",
  18228=>"101101100",
  18229=>"011010010",
  18230=>"000111100",
  18231=>"101001011",
  18232=>"101010010",
  18233=>"011110110",
  18234=>"000000001",
  18235=>"100001000",
  18236=>"100110010",
  18237=>"101110100",
  18238=>"000110101",
  18239=>"110001001",
  18240=>"000000100",
  18241=>"101001010",
  18242=>"111110111",
  18243=>"011100100",
  18244=>"111110110",
  18245=>"010011000",
  18246=>"010011100",
  18247=>"001110111",
  18248=>"100100010",
  18249=>"011101101",
  18250=>"110100010",
  18251=>"101010110",
  18252=>"001001111",
  18253=>"101000101",
  18254=>"010101111",
  18255=>"001011001",
  18256=>"100011000",
  18257=>"101110100",
  18258=>"001000101",
  18259=>"110100011",
  18260=>"000000111",
  18261=>"100001101",
  18262=>"010101010",
  18263=>"001000000",
  18264=>"001100111",
  18265=>"101100101",
  18266=>"100110000",
  18267=>"111110000",
  18268=>"010100111",
  18269=>"110111110",
  18270=>"011101101",
  18271=>"110111101",
  18272=>"011011000",
  18273=>"111001010",
  18274=>"001100101",
  18275=>"111101000",
  18276=>"011000000",
  18277=>"110001111",
  18278=>"011111000",
  18279=>"010011000",
  18280=>"100000000",
  18281=>"010000011",
  18282=>"001001010",
  18283=>"001101001",
  18284=>"010100100",
  18285=>"001101100",
  18286=>"010100011",
  18287=>"000010000",
  18288=>"011011001",
  18289=>"011011100",
  18290=>"010110111",
  18291=>"100001100",
  18292=>"110010000",
  18293=>"011011010",
  18294=>"110110111",
  18295=>"000101111",
  18296=>"001000110",
  18297=>"001100011",
  18298=>"011010010",
  18299=>"111111100",
  18300=>"001010100",
  18301=>"001010111",
  18302=>"101001111",
  18303=>"010010011",
  18304=>"000111011",
  18305=>"100101101",
  18306=>"110001000",
  18307=>"011000100",
  18308=>"011100001",
  18309=>"010001011",
  18310=>"011000000",
  18311=>"100100101",
  18312=>"011101100",
  18313=>"100111100",
  18314=>"100100001",
  18315=>"100100110",
  18316=>"010101110",
  18317=>"111011010",
  18318=>"000110101",
  18319=>"011100101",
  18320=>"101010100",
  18321=>"101110110",
  18322=>"000110001",
  18323=>"101100101",
  18324=>"010000000",
  18325=>"101110010",
  18326=>"111011011",
  18327=>"000000011",
  18328=>"101001100",
  18329=>"001011111",
  18330=>"010000100",
  18331=>"000100001",
  18332=>"000100110",
  18333=>"011001011",
  18334=>"000101101",
  18335=>"010000000",
  18336=>"010001001",
  18337=>"010001010",
  18338=>"010101000",
  18339=>"000110001",
  18340=>"100111111",
  18341=>"101101001",
  18342=>"101001000",
  18343=>"101000010",
  18344=>"111100000",
  18345=>"100101000",
  18346=>"011101001",
  18347=>"111110101",
  18348=>"111100001",
  18349=>"001000111",
  18350=>"100111000",
  18351=>"111000100",
  18352=>"010010000",
  18353=>"100000011",
  18354=>"101001101",
  18355=>"000111111",
  18356=>"110000000",
  18357=>"100001101",
  18358=>"001010001",
  18359=>"010100111",
  18360=>"001111100",
  18361=>"010111110",
  18362=>"101000100",
  18363=>"000000011",
  18364=>"010011111",
  18365=>"011011100",
  18366=>"110001010",
  18367=>"010011011",
  18368=>"111111010",
  18369=>"000000100",
  18370=>"001100110",
  18371=>"010001100",
  18372=>"110001111",
  18373=>"101010011",
  18374=>"001110100",
  18375=>"110101110",
  18376=>"110011111",
  18377=>"110101010",
  18378=>"110100001",
  18379=>"111010011",
  18380=>"100011000",
  18381=>"101001110",
  18382=>"010111011",
  18383=>"001111000",
  18384=>"111010010",
  18385=>"101011000",
  18386=>"010101011",
  18387=>"101010100",
  18388=>"100111100",
  18389=>"000010110",
  18390=>"000100100",
  18391=>"010010010",
  18392=>"000010101",
  18393=>"111111011",
  18394=>"010110101",
  18395=>"010011011",
  18396=>"011101111",
  18397=>"110011001",
  18398=>"000001101",
  18399=>"001000011",
  18400=>"111000110",
  18401=>"111101100",
  18402=>"100110000",
  18403=>"100101110",
  18404=>"101001101",
  18405=>"010111011",
  18406=>"001110011",
  18407=>"000001100",
  18408=>"010010100",
  18409=>"101011011",
  18410=>"010010110",
  18411=>"000101000",
  18412=>"001110000",
  18413=>"001100000",
  18414=>"010101011",
  18415=>"100000110",
  18416=>"101100101",
  18417=>"100100100",
  18418=>"100110111",
  18419=>"001101110",
  18420=>"000110111",
  18421=>"111011100",
  18422=>"000110110",
  18423=>"000010000",
  18424=>"100101001",
  18425=>"111001010",
  18426=>"101110011",
  18427=>"001110100",
  18428=>"101001111",
  18429=>"010101101",
  18430=>"101010001",
  18431=>"000110011",
  18432=>"100001100",
  18433=>"010011000",
  18434=>"011001010",
  18435=>"000000010",
  18436=>"010000111",
  18437=>"011010110",
  18438=>"000111011",
  18439=>"001001101",
  18440=>"110101000",
  18441=>"001111111",
  18442=>"000000010",
  18443=>"111111101",
  18444=>"100000000",
  18445=>"010000111",
  18446=>"111011100",
  18447=>"000111110",
  18448=>"000110001",
  18449=>"111010010",
  18450=>"101111110",
  18451=>"000101010",
  18452=>"000110001",
  18453=>"110111000",
  18454=>"101011010",
  18455=>"100101001",
  18456=>"000001111",
  18457=>"110000000",
  18458=>"110010011",
  18459=>"011101111",
  18460=>"010011010",
  18461=>"110111111",
  18462=>"010100111",
  18463=>"111001000",
  18464=>"001011000",
  18465=>"101001011",
  18466=>"111110110",
  18467=>"010011000",
  18468=>"010001011",
  18469=>"101110110",
  18470=>"101011111",
  18471=>"000001010",
  18472=>"110110101",
  18473=>"000000101",
  18474=>"010101010",
  18475=>"111011000",
  18476=>"111010000",
  18477=>"111101101",
  18478=>"000101110",
  18479=>"000010000",
  18480=>"000100001",
  18481=>"101110111",
  18482=>"100000110",
  18483=>"000111000",
  18484=>"100001111",
  18485=>"010111101",
  18486=>"110001001",
  18487=>"000010000",
  18488=>"000100011",
  18489=>"101101000",
  18490=>"000010001",
  18491=>"111011110",
  18492=>"111110001",
  18493=>"001010000",
  18494=>"010110001",
  18495=>"001101010",
  18496=>"001110010",
  18497=>"111110010",
  18498=>"000010100",
  18499=>"010110111",
  18500=>"111100000",
  18501=>"111110110",
  18502=>"110100100",
  18503=>"011010010",
  18504=>"101110000",
  18505=>"100111100",
  18506=>"101100000",
  18507=>"001101010",
  18508=>"001010111",
  18509=>"001011101",
  18510=>"011000010",
  18511=>"000110100",
  18512=>"010100100",
  18513=>"101000111",
  18514=>"000111110",
  18515=>"000100000",
  18516=>"101000101",
  18517=>"011110011",
  18518=>"100011110",
  18519=>"001100000",
  18520=>"101100101",
  18521=>"100101110",
  18522=>"101110000",
  18523=>"110000100",
  18524=>"011111001",
  18525=>"100010110",
  18526=>"100111010",
  18527=>"011111010",
  18528=>"111111111",
  18529=>"010100100",
  18530=>"111111001",
  18531=>"100010001",
  18532=>"101011001",
  18533=>"111000010",
  18534=>"101001101",
  18535=>"010111100",
  18536=>"110111011",
  18537=>"101010100",
  18538=>"000000000",
  18539=>"011000100",
  18540=>"100100000",
  18541=>"000011100",
  18542=>"110010110",
  18543=>"011111111",
  18544=>"001000010",
  18545=>"111010111",
  18546=>"111111001",
  18547=>"110111000",
  18548=>"101010001",
  18549=>"110111111",
  18550=>"011011100",
  18551=>"100001001",
  18552=>"111000110",
  18553=>"001100101",
  18554=>"010111010",
  18555=>"000101001",
  18556=>"110100010",
  18557=>"111000110",
  18558=>"000100111",
  18559=>"111000100",
  18560=>"000000010",
  18561=>"110011000",
  18562=>"100110101",
  18563=>"011111000",
  18564=>"111100010",
  18565=>"110101001",
  18566=>"110011001",
  18567=>"100111100",
  18568=>"001000111",
  18569=>"101000100",
  18570=>"000001010",
  18571=>"010011101",
  18572=>"011110100",
  18573=>"011001001",
  18574=>"111110010",
  18575=>"110100101",
  18576=>"000111110",
  18577=>"000010111",
  18578=>"001001111",
  18579=>"000010111",
  18580=>"011100110",
  18581=>"101101010",
  18582=>"011101001",
  18583=>"010000100",
  18584=>"001001110",
  18585=>"100100100",
  18586=>"101010110",
  18587=>"111011111",
  18588=>"111111101",
  18589=>"101011101",
  18590=>"111000010",
  18591=>"111100101",
  18592=>"000100110",
  18593=>"110110111",
  18594=>"101001010",
  18595=>"110111101",
  18596=>"000010111",
  18597=>"100011101",
  18598=>"001010100",
  18599=>"101001100",
  18600=>"100111111",
  18601=>"011111101",
  18602=>"001010100",
  18603=>"000010000",
  18604=>"110111010",
  18605=>"000111111",
  18606=>"111001011",
  18607=>"000111110",
  18608=>"000101011",
  18609=>"101000000",
  18610=>"001100100",
  18611=>"101001101",
  18612=>"111111111",
  18613=>"011100010",
  18614=>"111101000",
  18615=>"011000101",
  18616=>"111100010",
  18617=>"100000111",
  18618=>"001000011",
  18619=>"110001111",
  18620=>"110001001",
  18621=>"101110001",
  18622=>"011100100",
  18623=>"111001110",
  18624=>"100111000",
  18625=>"000001000",
  18626=>"010101011",
  18627=>"100010001",
  18628=>"111000101",
  18629=>"000000110",
  18630=>"101101101",
  18631=>"100001001",
  18632=>"111100011",
  18633=>"000100000",
  18634=>"000100111",
  18635=>"000000010",
  18636=>"101111000",
  18637=>"111111110",
  18638=>"001110001",
  18639=>"000001001",
  18640=>"001001000",
  18641=>"111010011",
  18642=>"010101010",
  18643=>"110111111",
  18644=>"110111111",
  18645=>"101111011",
  18646=>"010011001",
  18647=>"110111110",
  18648=>"011000001",
  18649=>"010111111",
  18650=>"000010100",
  18651=>"111100100",
  18652=>"011010001",
  18653=>"001111000",
  18654=>"101110111",
  18655=>"011010110",
  18656=>"101001000",
  18657=>"011101000",
  18658=>"111101011",
  18659=>"100001110",
  18660=>"010101011",
  18661=>"000000011",
  18662=>"101100010",
  18663=>"101101001",
  18664=>"111110111",
  18665=>"110011101",
  18666=>"001000000",
  18667=>"000110100",
  18668=>"101011000",
  18669=>"100101100",
  18670=>"000000100",
  18671=>"001111101",
  18672=>"111101011",
  18673=>"000010010",
  18674=>"010100011",
  18675=>"111011011",
  18676=>"111100110",
  18677=>"011001011",
  18678=>"000010001",
  18679=>"100100011",
  18680=>"001011111",
  18681=>"001100001",
  18682=>"011001011",
  18683=>"111000100",
  18684=>"110110011",
  18685=>"011010000",
  18686=>"000000000",
  18687=>"001110100",
  18688=>"001000010",
  18689=>"111011111",
  18690=>"100011100",
  18691=>"100011100",
  18692=>"010011100",
  18693=>"111000101",
  18694=>"110011010",
  18695=>"010110000",
  18696=>"110001111",
  18697=>"100011101",
  18698=>"011101001",
  18699=>"001001111",
  18700=>"010110000",
  18701=>"111110110",
  18702=>"010101010",
  18703=>"100100001",
  18704=>"101101100",
  18705=>"010000100",
  18706=>"110110000",
  18707=>"001011000",
  18708=>"100000010",
  18709=>"010000111",
  18710=>"111000101",
  18711=>"101000100",
  18712=>"001110101",
  18713=>"110000011",
  18714=>"000001111",
  18715=>"010001000",
  18716=>"110011111",
  18717=>"110101101",
  18718=>"000000100",
  18719=>"011010100",
  18720=>"000001001",
  18721=>"111101011",
  18722=>"010111001",
  18723=>"001000001",
  18724=>"101001000",
  18725=>"100101001",
  18726=>"100011001",
  18727=>"101010001",
  18728=>"001101100",
  18729=>"100111111",
  18730=>"111011001",
  18731=>"110010001",
  18732=>"011001111",
  18733=>"010000011",
  18734=>"111100110",
  18735=>"000001010",
  18736=>"100101100",
  18737=>"011100001",
  18738=>"000000010",
  18739=>"010011000",
  18740=>"001000111",
  18741=>"001101010",
  18742=>"100001111",
  18743=>"011111100",
  18744=>"101000000",
  18745=>"110000011",
  18746=>"000001001",
  18747=>"011010010",
  18748=>"111011111",
  18749=>"100101111",
  18750=>"111100101",
  18751=>"101110010",
  18752=>"101000110",
  18753=>"001101101",
  18754=>"000010110",
  18755=>"101010110",
  18756=>"111010010",
  18757=>"011101100",
  18758=>"011001001",
  18759=>"110100111",
  18760=>"111111011",
  18761=>"011001010",
  18762=>"011011000",
  18763=>"011011000",
  18764=>"111010000",
  18765=>"101001000",
  18766=>"111110110",
  18767=>"100010110",
  18768=>"110111110",
  18769=>"001010110",
  18770=>"000110110",
  18771=>"101111110",
  18772=>"001010101",
  18773=>"000110001",
  18774=>"000111000",
  18775=>"100111111",
  18776=>"110101110",
  18777=>"111101010",
  18778=>"101011010",
  18779=>"010100000",
  18780=>"111011111",
  18781=>"111001111",
  18782=>"011110011",
  18783=>"001011010",
  18784=>"011100101",
  18785=>"101110010",
  18786=>"010000010",
  18787=>"101001001",
  18788=>"110100010",
  18789=>"001011010",
  18790=>"001101110",
  18791=>"010001000",
  18792=>"100110101",
  18793=>"111101101",
  18794=>"110000101",
  18795=>"011010010",
  18796=>"000010111",
  18797=>"101110000",
  18798=>"011100111",
  18799=>"110010000",
  18800=>"001011111",
  18801=>"001011001",
  18802=>"011100101",
  18803=>"000010110",
  18804=>"100000011",
  18805=>"111101010",
  18806=>"011011010",
  18807=>"111110011",
  18808=>"010010000",
  18809=>"110101000",
  18810=>"100011011",
  18811=>"000010111",
  18812=>"010010000",
  18813=>"011101000",
  18814=>"010000100",
  18815=>"101001100",
  18816=>"000101000",
  18817=>"101001111",
  18818=>"011000010",
  18819=>"111001100",
  18820=>"101011110",
  18821=>"010011011",
  18822=>"001010101",
  18823=>"111000111",
  18824=>"111101100",
  18825=>"110110000",
  18826=>"000000010",
  18827=>"001010000",
  18828=>"000100110",
  18829=>"100000000",
  18830=>"010010110",
  18831=>"010001010",
  18832=>"110010111",
  18833=>"011111111",
  18834=>"011101111",
  18835=>"101101110",
  18836=>"000111100",
  18837=>"110111100",
  18838=>"000010111",
  18839=>"111011001",
  18840=>"001110111",
  18841=>"110010010",
  18842=>"111111100",
  18843=>"111101011",
  18844=>"110110110",
  18845=>"010010000",
  18846=>"010111011",
  18847=>"010110110",
  18848=>"101101010",
  18849=>"001001111",
  18850=>"010010011",
  18851=>"111111111",
  18852=>"100110101",
  18853=>"010001111",
  18854=>"110010111",
  18855=>"010011010",
  18856=>"100010000",
  18857=>"011000011",
  18858=>"101101101",
  18859=>"111000101",
  18860=>"100011101",
  18861=>"111110000",
  18862=>"101000001",
  18863=>"001001010",
  18864=>"111101011",
  18865=>"001111111",
  18866=>"000000000",
  18867=>"011000010",
  18868=>"000111000",
  18869=>"010001100",
  18870=>"011110101",
  18871=>"111010000",
  18872=>"111001001",
  18873=>"001100010",
  18874=>"100100100",
  18875=>"111010011",
  18876=>"000100010",
  18877=>"000001001",
  18878=>"101111100",
  18879=>"010010001",
  18880=>"001000100",
  18881=>"000000010",
  18882=>"111110100",
  18883=>"011111000",
  18884=>"101110111",
  18885=>"000101101",
  18886=>"001000000",
  18887=>"010000101",
  18888=>"111010110",
  18889=>"111011000",
  18890=>"111111101",
  18891=>"011011101",
  18892=>"000100111",
  18893=>"110000110",
  18894=>"010000101",
  18895=>"101001101",
  18896=>"010011000",
  18897=>"101101001",
  18898=>"001101111",
  18899=>"000010010",
  18900=>"000010011",
  18901=>"011110110",
  18902=>"011110011",
  18903=>"000011110",
  18904=>"000001111",
  18905=>"001010000",
  18906=>"100111111",
  18907=>"001111110",
  18908=>"111010100",
  18909=>"011001001",
  18910=>"100101000",
  18911=>"110000010",
  18912=>"111010000",
  18913=>"011111110",
  18914=>"110000011",
  18915=>"101100000",
  18916=>"011100011",
  18917=>"011101100",
  18918=>"011100001",
  18919=>"101111001",
  18920=>"011110100",
  18921=>"000000001",
  18922=>"011101101",
  18923=>"001011111",
  18924=>"000100011",
  18925=>"000011110",
  18926=>"100011000",
  18927=>"000110111",
  18928=>"000101001",
  18929=>"101001011",
  18930=>"010110100",
  18931=>"100000100",
  18932=>"111101101",
  18933=>"110011100",
  18934=>"001100111",
  18935=>"001110011",
  18936=>"111001011",
  18937=>"100110111",
  18938=>"100001100",
  18939=>"101011100",
  18940=>"001100111",
  18941=>"000011101",
  18942=>"011110000",
  18943=>"100111011",
  18944=>"111001001",
  18945=>"111001010",
  18946=>"011100000",
  18947=>"111001011",
  18948=>"010001011",
  18949=>"110000101",
  18950=>"101111110",
  18951=>"001100111",
  18952=>"110110010",
  18953=>"011101101",
  18954=>"010110011",
  18955=>"110110000",
  18956=>"100011110",
  18957=>"100011101",
  18958=>"011111010",
  18959=>"101001010",
  18960=>"011000010",
  18961=>"001010110",
  18962=>"100010011",
  18963=>"100101100",
  18964=>"111010100",
  18965=>"100010010",
  18966=>"100110111",
  18967=>"001101111",
  18968=>"001101100",
  18969=>"110101010",
  18970=>"000111110",
  18971=>"100010100",
  18972=>"100011111",
  18973=>"010101100",
  18974=>"100110100",
  18975=>"011111111",
  18976=>"101001111",
  18977=>"111110011",
  18978=>"111111000",
  18979=>"100110011",
  18980=>"110010110",
  18981=>"001010000",
  18982=>"111101110",
  18983=>"000110110",
  18984=>"001001011",
  18985=>"101000111",
  18986=>"111111101",
  18987=>"010001100",
  18988=>"011000011",
  18989=>"000001111",
  18990=>"111001101",
  18991=>"000111010",
  18992=>"011100000",
  18993=>"100100000",
  18994=>"101001010",
  18995=>"000101010",
  18996=>"111011001",
  18997=>"010100011",
  18998=>"011101001",
  18999=>"101000000",
  19000=>"010001110",
  19001=>"100111100",
  19002=>"100101000",
  19003=>"011100100",
  19004=>"110110111",
  19005=>"100000011",
  19006=>"101101001",
  19007=>"000110000",
  19008=>"101000000",
  19009=>"110000001",
  19010=>"011001000",
  19011=>"101110110",
  19012=>"000111000",
  19013=>"101010101",
  19014=>"111000100",
  19015=>"000110100",
  19016=>"110101000",
  19017=>"111000001",
  19018=>"000110000",
  19019=>"101110011",
  19020=>"110101000",
  19021=>"100011110",
  19022=>"011010000",
  19023=>"011001111",
  19024=>"111101111",
  19025=>"001001111",
  19026=>"000011101",
  19027=>"111111101",
  19028=>"110011101",
  19029=>"100111001",
  19030=>"011101010",
  19031=>"100110110",
  19032=>"111011111",
  19033=>"101001000",
  19034=>"001110110",
  19035=>"100111001",
  19036=>"111010111",
  19037=>"100100011",
  19038=>"101011010",
  19039=>"001111010",
  19040=>"011101100",
  19041=>"010110111",
  19042=>"010100010",
  19043=>"101111110",
  19044=>"101000000",
  19045=>"100001100",
  19046=>"111110110",
  19047=>"111010111",
  19048=>"001011001",
  19049=>"000000000",
  19050=>"000101100",
  19051=>"011111101",
  19052=>"001011010",
  19053=>"001101101",
  19054=>"001001010",
  19055=>"110001000",
  19056=>"000010101",
  19057=>"011001011",
  19058=>"101010101",
  19059=>"111111110",
  19060=>"000100101",
  19061=>"011000010",
  19062=>"111000010",
  19063=>"111101011",
  19064=>"110111100",
  19065=>"001001111",
  19066=>"111100101",
  19067=>"000001010",
  19068=>"110111111",
  19069=>"000001100",
  19070=>"001110110",
  19071=>"011101000",
  19072=>"101100101",
  19073=>"101001010",
  19074=>"111101111",
  19075=>"000010011",
  19076=>"100101100",
  19077=>"011101101",
  19078=>"000001111",
  19079=>"000100111",
  19080=>"011101111",
  19081=>"110100011",
  19082=>"101100101",
  19083=>"010111001",
  19084=>"111011101",
  19085=>"010011101",
  19086=>"110011111",
  19087=>"110011100",
  19088=>"111110101",
  19089=>"110011101",
  19090=>"110010001",
  19091=>"000111000",
  19092=>"000010000",
  19093=>"001110000",
  19094=>"010000110",
  19095=>"110101000",
  19096=>"111010111",
  19097=>"101110010",
  19098=>"101111011",
  19099=>"100010010",
  19100=>"000000101",
  19101=>"101000110",
  19102=>"110110010",
  19103=>"000101110",
  19104=>"000001100",
  19105=>"001111101",
  19106=>"111101010",
  19107=>"111100000",
  19108=>"010001011",
  19109=>"100001001",
  19110=>"101010110",
  19111=>"011001101",
  19112=>"000001011",
  19113=>"011010111",
  19114=>"001011101",
  19115=>"001010101",
  19116=>"000010111",
  19117=>"101110111",
  19118=>"010101101",
  19119=>"010101100",
  19120=>"101100001",
  19121=>"111101111",
  19122=>"011101010",
  19123=>"000101101",
  19124=>"110101011",
  19125=>"101011001",
  19126=>"000001100",
  19127=>"011000000",
  19128=>"011010000",
  19129=>"001111010",
  19130=>"010110001",
  19131=>"111011001",
  19132=>"001000001",
  19133=>"101010101",
  19134=>"100100100",
  19135=>"100111001",
  19136=>"100000011",
  19137=>"000011011",
  19138=>"110010101",
  19139=>"010100011",
  19140=>"110000000",
  19141=>"011100100",
  19142=>"010010111",
  19143=>"111001111",
  19144=>"100101110",
  19145=>"111110000",
  19146=>"000011010",
  19147=>"001011001",
  19148=>"001011101",
  19149=>"001001010",
  19150=>"100110000",
  19151=>"011111100",
  19152=>"001000111",
  19153=>"101001010",
  19154=>"101110100",
  19155=>"000101000",
  19156=>"111001100",
  19157=>"110001101",
  19158=>"010100010",
  19159=>"000010100",
  19160=>"100111101",
  19161=>"011001111",
  19162=>"001000100",
  19163=>"110111000",
  19164=>"001111111",
  19165=>"111101100",
  19166=>"100100011",
  19167=>"100000010",
  19168=>"100110110",
  19169=>"001101101",
  19170=>"001001010",
  19171=>"010010111",
  19172=>"001010000",
  19173=>"111101000",
  19174=>"000010001",
  19175=>"111111010",
  19176=>"110110000",
  19177=>"100111100",
  19178=>"111100010",
  19179=>"000011010",
  19180=>"010001111",
  19181=>"001101100",
  19182=>"101000101",
  19183=>"001100001",
  19184=>"001010010",
  19185=>"111101111",
  19186=>"100011011",
  19187=>"000101101",
  19188=>"011101000",
  19189=>"001000011",
  19190=>"001001100",
  19191=>"011000011",
  19192=>"101001000",
  19193=>"110100101",
  19194=>"001011111",
  19195=>"011001100",
  19196=>"111110100",
  19197=>"000111011",
  19198=>"111111011",
  19199=>"000011000",
  19200=>"000101010",
  19201=>"100110010",
  19202=>"101100111",
  19203=>"111111100",
  19204=>"111000011",
  19205=>"101111100",
  19206=>"100111000",
  19207=>"111010011",
  19208=>"001011111",
  19209=>"110100000",
  19210=>"100000000",
  19211=>"111111011",
  19212=>"001001000",
  19213=>"001110010",
  19214=>"011100011",
  19215=>"101011111",
  19216=>"001011101",
  19217=>"101010000",
  19218=>"110000100",
  19219=>"001001000",
  19220=>"001101001",
  19221=>"010010000",
  19222=>"111100000",
  19223=>"010011110",
  19224=>"101000111",
  19225=>"110001101",
  19226=>"110010100",
  19227=>"101111011",
  19228=>"010000000",
  19229=>"111110010",
  19230=>"111101010",
  19231=>"011000100",
  19232=>"000100000",
  19233=>"010001010",
  19234=>"001001101",
  19235=>"010000101",
  19236=>"011011101",
  19237=>"000000001",
  19238=>"110111111",
  19239=>"100101010",
  19240=>"100011101",
  19241=>"010001010",
  19242=>"111110100",
  19243=>"100100000",
  19244=>"100100001",
  19245=>"000000111",
  19246=>"111100000",
  19247=>"101111100",
  19248=>"011100111",
  19249=>"110000000",
  19250=>"111000111",
  19251=>"100100000",
  19252=>"111001000",
  19253=>"011100101",
  19254=>"001010011",
  19255=>"010100111",
  19256=>"000110110",
  19257=>"101011111",
  19258=>"001011100",
  19259=>"010101011",
  19260=>"001100111",
  19261=>"001110111",
  19262=>"010101010",
  19263=>"001110011",
  19264=>"100100000",
  19265=>"010001011",
  19266=>"001000000",
  19267=>"111000011",
  19268=>"000011001",
  19269=>"001000010",
  19270=>"001010001",
  19271=>"111011010",
  19272=>"010101100",
  19273=>"100010111",
  19274=>"001110000",
  19275=>"101001110",
  19276=>"000101100",
  19277=>"100010001",
  19278=>"111110101",
  19279=>"010001111",
  19280=>"100111110",
  19281=>"001001011",
  19282=>"001001101",
  19283=>"011000010",
  19284=>"111010110",
  19285=>"010101111",
  19286=>"000010110",
  19287=>"000101001",
  19288=>"111100011",
  19289=>"110111010",
  19290=>"001000000",
  19291=>"000100001",
  19292=>"000011011",
  19293=>"110110111",
  19294=>"111010110",
  19295=>"010010010",
  19296=>"001110111",
  19297=>"000101111",
  19298=>"100000111",
  19299=>"111100010",
  19300=>"111110110",
  19301=>"000000011",
  19302=>"100011101",
  19303=>"010000000",
  19304=>"101010010",
  19305=>"010101010",
  19306=>"111100010",
  19307=>"100011010",
  19308=>"101111110",
  19309=>"110011111",
  19310=>"111111011",
  19311=>"100101010",
  19312=>"111001001",
  19313=>"010010111",
  19314=>"011101111",
  19315=>"001100101",
  19316=>"010011010",
  19317=>"000010101",
  19318=>"000110000",
  19319=>"001000010",
  19320=>"110001000",
  19321=>"011011000",
  19322=>"011100111",
  19323=>"110010000",
  19324=>"101010111",
  19325=>"010101100",
  19326=>"111000110",
  19327=>"100011001",
  19328=>"011001001",
  19329=>"111111000",
  19330=>"101111000",
  19331=>"011100010",
  19332=>"000010110",
  19333=>"111111111",
  19334=>"001110111",
  19335=>"011110010",
  19336=>"111101010",
  19337=>"111111110",
  19338=>"111100111",
  19339=>"111100101",
  19340=>"010000110",
  19341=>"001101110",
  19342=>"001001101",
  19343=>"011010011",
  19344=>"111111001",
  19345=>"011010011",
  19346=>"001110011",
  19347=>"001111101",
  19348=>"111110001",
  19349=>"100001011",
  19350=>"111010001",
  19351=>"110001010",
  19352=>"000011100",
  19353=>"100011111",
  19354=>"100111101",
  19355=>"101011111",
  19356=>"100110111",
  19357=>"110001101",
  19358=>"101110101",
  19359=>"110100101",
  19360=>"101100011",
  19361=>"101011001",
  19362=>"000101010",
  19363=>"001000000",
  19364=>"001010001",
  19365=>"100100011",
  19366=>"001110000",
  19367=>"100011110",
  19368=>"011011000",
  19369=>"010000111",
  19370=>"101010011",
  19371=>"011111110",
  19372=>"010001111",
  19373=>"001001100",
  19374=>"010110101",
  19375=>"101000011",
  19376=>"100111001",
  19377=>"000101001",
  19378=>"010100001",
  19379=>"101100001",
  19380=>"111000110",
  19381=>"100001100",
  19382=>"010101001",
  19383=>"101011001",
  19384=>"111111111",
  19385=>"110111000",
  19386=>"010000010",
  19387=>"000110000",
  19388=>"000010011",
  19389=>"111001111",
  19390=>"101001010",
  19391=>"101000001",
  19392=>"111110010",
  19393=>"100100101",
  19394=>"000100101",
  19395=>"101100001",
  19396=>"101101101",
  19397=>"000111111",
  19398=>"001011100",
  19399=>"010001110",
  19400=>"110101011",
  19401=>"011100111",
  19402=>"110111000",
  19403=>"010001110",
  19404=>"001001000",
  19405=>"011000000",
  19406=>"011110101",
  19407=>"000111100",
  19408=>"000110001",
  19409=>"011110001",
  19410=>"010100001",
  19411=>"010100011",
  19412=>"101100010",
  19413=>"011101000",
  19414=>"010110111",
  19415=>"100111110",
  19416=>"010011010",
  19417=>"110111111",
  19418=>"110101110",
  19419=>"101100110",
  19420=>"101100110",
  19421=>"110011101",
  19422=>"100011110",
  19423=>"010010001",
  19424=>"111011000",
  19425=>"010010100",
  19426=>"000101010",
  19427=>"111100100",
  19428=>"000000000",
  19429=>"100111000",
  19430=>"111010001",
  19431=>"010000101",
  19432=>"101001000",
  19433=>"100100101",
  19434=>"000000010",
  19435=>"100011100",
  19436=>"000101111",
  19437=>"101001000",
  19438=>"111110000",
  19439=>"111001000",
  19440=>"111001001",
  19441=>"011101100",
  19442=>"000101001",
  19443=>"100000111",
  19444=>"111011000",
  19445=>"100101011",
  19446=>"010010001",
  19447=>"000000011",
  19448=>"010010110",
  19449=>"111011001",
  19450=>"100010001",
  19451=>"000010111",
  19452=>"111100000",
  19453=>"100000010",
  19454=>"111101110",
  19455=>"000111011",
  19456=>"010001110",
  19457=>"100000110",
  19458=>"011110101",
  19459=>"111110001",
  19460=>"110011011",
  19461=>"000111111",
  19462=>"110101001",
  19463=>"100001101",
  19464=>"000011001",
  19465=>"000010001",
  19466=>"010100110",
  19467=>"110001100",
  19468=>"000000010",
  19469=>"111110111",
  19470=>"011000110",
  19471=>"000111010",
  19472=>"101001111",
  19473=>"011010101",
  19474=>"000011101",
  19475=>"011101101",
  19476=>"000000110",
  19477=>"011110001",
  19478=>"101000101",
  19479=>"010000000",
  19480=>"100011101",
  19481=>"111001010",
  19482=>"110100110",
  19483=>"110000101",
  19484=>"010111100",
  19485=>"011100001",
  19486=>"010101111",
  19487=>"101111101",
  19488=>"011001000",
  19489=>"100100100",
  19490=>"010100111",
  19491=>"010110100",
  19492=>"010110101",
  19493=>"111001000",
  19494=>"010001010",
  19495=>"011101010",
  19496=>"101001001",
  19497=>"001000100",
  19498=>"000011000",
  19499=>"111000001",
  19500=>"110001011",
  19501=>"001100111",
  19502=>"100001101",
  19503=>"010100110",
  19504=>"011000110",
  19505=>"010010010",
  19506=>"011010011",
  19507=>"100101100",
  19508=>"101111100",
  19509=>"010001100",
  19510=>"101000111",
  19511=>"010000001",
  19512=>"100100100",
  19513=>"110011101",
  19514=>"001010100",
  19515=>"110100000",
  19516=>"000010110",
  19517=>"010000100",
  19518=>"001000111",
  19519=>"101001111",
  19520=>"111101011",
  19521=>"100000111",
  19522=>"001101001",
  19523=>"011110110",
  19524=>"110110010",
  19525=>"101000100",
  19526=>"000110000",
  19527=>"111001001",
  19528=>"100101000",
  19529=>"100010111",
  19530=>"000010010",
  19531=>"010001101",
  19532=>"110110111",
  19533=>"011111010",
  19534=>"011011100",
  19535=>"010010001",
  19536=>"010001101",
  19537=>"000000001",
  19538=>"011001110",
  19539=>"100110011",
  19540=>"011111101",
  19541=>"000010100",
  19542=>"111010100",
  19543=>"000111000",
  19544=>"101100101",
  19545=>"101001100",
  19546=>"011110101",
  19547=>"001100000",
  19548=>"101110010",
  19549=>"110101100",
  19550=>"111110111",
  19551=>"110000010",
  19552=>"011001001",
  19553=>"000001000",
  19554=>"111111110",
  19555=>"110111100",
  19556=>"110110101",
  19557=>"101110101",
  19558=>"001101101",
  19559=>"111010001",
  19560=>"000110010",
  19561=>"111100111",
  19562=>"011100110",
  19563=>"110101100",
  19564=>"010111110",
  19565=>"110001110",
  19566=>"000000100",
  19567=>"011101011",
  19568=>"101100001",
  19569=>"111011000",
  19570=>"010100101",
  19571=>"000001100",
  19572=>"101111001",
  19573=>"011101100",
  19574=>"110110110",
  19575=>"100101010",
  19576=>"001101111",
  19577=>"101111111",
  19578=>"100001010",
  19579=>"101001000",
  19580=>"011000111",
  19581=>"001000101",
  19582=>"110111101",
  19583=>"001010010",
  19584=>"110110000",
  19585=>"011100011",
  19586=>"100010011",
  19587=>"101010000",
  19588=>"111100011",
  19589=>"110001010",
  19590=>"110110010",
  19591=>"110100010",
  19592=>"001111000",
  19593=>"111001010",
  19594=>"111110001",
  19595=>"001011001",
  19596=>"011010111",
  19597=>"010111000",
  19598=>"101111011",
  19599=>"001100001",
  19600=>"100010001",
  19601=>"000100011",
  19602=>"011101111",
  19603=>"000110000",
  19604=>"101110000",
  19605=>"010010010",
  19606=>"001000000",
  19607=>"110111010",
  19608=>"000110000",
  19609=>"010011000",
  19610=>"101100111",
  19611=>"101110110",
  19612=>"000011101",
  19613=>"001110100",
  19614=>"000000100",
  19615=>"101100000",
  19616=>"000011111",
  19617=>"011101100",
  19618=>"011011011",
  19619=>"010111010",
  19620=>"110101110",
  19621=>"110111111",
  19622=>"111100100",
  19623=>"000101010",
  19624=>"101110101",
  19625=>"111001011",
  19626=>"101110100",
  19627=>"100110101",
  19628=>"100111000",
  19629=>"111011001",
  19630=>"011111101",
  19631=>"011111101",
  19632=>"101000001",
  19633=>"110000111",
  19634=>"100000101",
  19635=>"000000101",
  19636=>"001011011",
  19637=>"011100011",
  19638=>"011000010",
  19639=>"100011000",
  19640=>"100111010",
  19641=>"011011010",
  19642=>"001010100",
  19643=>"000100100",
  19644=>"101011011",
  19645=>"111101011",
  19646=>"101110111",
  19647=>"010000011",
  19648=>"011101001",
  19649=>"111001101",
  19650=>"001000001",
  19651=>"010010001",
  19652=>"100101010",
  19653=>"101100000",
  19654=>"101110110",
  19655=>"110101100",
  19656=>"001000111",
  19657=>"101100011",
  19658=>"101100000",
  19659=>"010000100",
  19660=>"101101110",
  19661=>"001110111",
  19662=>"001100101",
  19663=>"011111000",
  19664=>"001001101",
  19665=>"011101010",
  19666=>"100010000",
  19667=>"011011110",
  19668=>"111110001",
  19669=>"011010100",
  19670=>"100101110",
  19671=>"110111101",
  19672=>"111111110",
  19673=>"111101000",
  19674=>"011111010",
  19675=>"100000010",
  19676=>"000101111",
  19677=>"100110101",
  19678=>"001001011",
  19679=>"011100110",
  19680=>"000001110",
  19681=>"001010101",
  19682=>"010000010",
  19683=>"011100000",
  19684=>"010000001",
  19685=>"010100110",
  19686=>"000010111",
  19687=>"001101011",
  19688=>"010011010",
  19689=>"010110010",
  19690=>"011001110",
  19691=>"101100100",
  19692=>"111001010",
  19693=>"110001100",
  19694=>"100110011",
  19695=>"111101111",
  19696=>"111110110",
  19697=>"111100101",
  19698=>"011110010",
  19699=>"011111111",
  19700=>"100000001",
  19701=>"000000111",
  19702=>"101010000",
  19703=>"111010100",
  19704=>"110000100",
  19705=>"000101110",
  19706=>"111111110",
  19707=>"110010000",
  19708=>"101000001",
  19709=>"010010111",
  19710=>"001100001",
  19711=>"010000000",
  19712=>"011110010",
  19713=>"011111111",
  19714=>"000011101",
  19715=>"101011011",
  19716=>"101111000",
  19717=>"011000010",
  19718=>"111101011",
  19719=>"100110101",
  19720=>"011000000",
  19721=>"110111001",
  19722=>"111011111",
  19723=>"110010010",
  19724=>"111001100",
  19725=>"001001011",
  19726=>"100111101",
  19727=>"001001000",
  19728=>"000101110",
  19729=>"111011001",
  19730=>"101100010",
  19731=>"101101010",
  19732=>"000010101",
  19733=>"100001111",
  19734=>"000000010",
  19735=>"100011111",
  19736=>"101110110",
  19737=>"010110001",
  19738=>"100101001",
  19739=>"110011111",
  19740=>"001011010",
  19741=>"101011110",
  19742=>"000000110",
  19743=>"101010010",
  19744=>"000000110",
  19745=>"000110011",
  19746=>"110111111",
  19747=>"100011011",
  19748=>"100111010",
  19749=>"111000011",
  19750=>"101001100",
  19751=>"111011111",
  19752=>"100011110",
  19753=>"101000111",
  19754=>"100010101",
  19755=>"111011111",
  19756=>"011001001",
  19757=>"000001001",
  19758=>"010010100",
  19759=>"101000111",
  19760=>"010001101",
  19761=>"001111011",
  19762=>"111111110",
  19763=>"010001110",
  19764=>"000111101",
  19765=>"000100011",
  19766=>"001100101",
  19767=>"110101110",
  19768=>"111000100",
  19769=>"010111110",
  19770=>"000100010",
  19771=>"010111111",
  19772=>"111011000",
  19773=>"000001101",
  19774=>"110100111",
  19775=>"100100011",
  19776=>"000001011",
  19777=>"000100010",
  19778=>"010000101",
  19779=>"110010001",
  19780=>"010011100",
  19781=>"110111001",
  19782=>"111000100",
  19783=>"000001101",
  19784=>"010001000",
  19785=>"011000010",
  19786=>"010000001",
  19787=>"000010011",
  19788=>"100111010",
  19789=>"110010100",
  19790=>"011000000",
  19791=>"111011101",
  19792=>"111100010",
  19793=>"010011010",
  19794=>"101110101",
  19795=>"000001110",
  19796=>"010011001",
  19797=>"011001101",
  19798=>"110100100",
  19799=>"100000110",
  19800=>"000100011",
  19801=>"101000000",
  19802=>"011011111",
  19803=>"100101001",
  19804=>"001101110",
  19805=>"100010101",
  19806=>"111011100",
  19807=>"000110101",
  19808=>"010011111",
  19809=>"000011100",
  19810=>"111111110",
  19811=>"001101000",
  19812=>"111101101",
  19813=>"110111111",
  19814=>"001111110",
  19815=>"010000110",
  19816=>"100010111",
  19817=>"000011100",
  19818=>"011110111",
  19819=>"110100001",
  19820=>"001001010",
  19821=>"101111000",
  19822=>"110001001",
  19823=>"001011110",
  19824=>"001100101",
  19825=>"101000111",
  19826=>"010011110",
  19827=>"110100110",
  19828=>"001000100",
  19829=>"011110000",
  19830=>"100011101",
  19831=>"011101001",
  19832=>"000101001",
  19833=>"100100011",
  19834=>"000001111",
  19835=>"110000111",
  19836=>"101001101",
  19837=>"100000101",
  19838=>"000010101",
  19839=>"111000110",
  19840=>"110100110",
  19841=>"011101011",
  19842=>"111010101",
  19843=>"100111000",
  19844=>"000111111",
  19845=>"111101000",
  19846=>"100001100",
  19847=>"101000000",
  19848=>"000010100",
  19849=>"001010100",
  19850=>"000100101",
  19851=>"010010110",
  19852=>"011110011",
  19853=>"010011111",
  19854=>"101101100",
  19855=>"100011110",
  19856=>"100111101",
  19857=>"010011011",
  19858=>"100111000",
  19859=>"110100110",
  19860=>"110101001",
  19861=>"000010110",
  19862=>"110111101",
  19863=>"111101101",
  19864=>"001010010",
  19865=>"001001010",
  19866=>"011000011",
  19867=>"001001010",
  19868=>"011000001",
  19869=>"010110101",
  19870=>"100011010",
  19871=>"111101111",
  19872=>"010111001",
  19873=>"010110001",
  19874=>"101111110",
  19875=>"001011000",
  19876=>"001000000",
  19877=>"000010010",
  19878=>"111010101",
  19879=>"011111010",
  19880=>"110111101",
  19881=>"000001001",
  19882=>"001001110",
  19883=>"001000010",
  19884=>"000110101",
  19885=>"101010010",
  19886=>"101111101",
  19887=>"111010001",
  19888=>"001111101",
  19889=>"110000100",
  19890=>"011010101",
  19891=>"000001011",
  19892=>"001111000",
  19893=>"110000000",
  19894=>"110010101",
  19895=>"000111100",
  19896=>"001100000",
  19897=>"010000101",
  19898=>"100000001",
  19899=>"010111011",
  19900=>"110001001",
  19901=>"100110011",
  19902=>"000001101",
  19903=>"010001001",
  19904=>"010010000",
  19905=>"110111000",
  19906=>"110011001",
  19907=>"001011110",
  19908=>"001000110",
  19909=>"000010101",
  19910=>"010010010",
  19911=>"101110000",
  19912=>"110110011",
  19913=>"101110111",
  19914=>"111001100",
  19915=>"111001001",
  19916=>"011001001",
  19917=>"100110101",
  19918=>"111010010",
  19919=>"100101010",
  19920=>"001111001",
  19921=>"011010100",
  19922=>"000010100",
  19923=>"110111111",
  19924=>"111000000",
  19925=>"101101111",
  19926=>"000100111",
  19927=>"001111001",
  19928=>"101111110",
  19929=>"010011011",
  19930=>"001011001",
  19931=>"100010110",
  19932=>"100010011",
  19933=>"000011100",
  19934=>"101111111",
  19935=>"011100111",
  19936=>"101101100",
  19937=>"000110101",
  19938=>"111101000",
  19939=>"011000100",
  19940=>"001111001",
  19941=>"100010000",
  19942=>"111000001",
  19943=>"010100001",
  19944=>"001011000",
  19945=>"000101111",
  19946=>"000000010",
  19947=>"001000110",
  19948=>"101110110",
  19949=>"001010010",
  19950=>"010000101",
  19951=>"000101111",
  19952=>"000011000",
  19953=>"010101100",
  19954=>"101111110",
  19955=>"011000000",
  19956=>"000000000",
  19957=>"011011000",
  19958=>"010000010",
  19959=>"000100001",
  19960=>"011010000",
  19961=>"000100111",
  19962=>"010100110",
  19963=>"101001111",
  19964=>"010011111",
  19965=>"111010011",
  19966=>"101001101",
  19967=>"000010000",
  19968=>"011011001",
  19969=>"011000100",
  19970=>"001010111",
  19971=>"111001010",
  19972=>"010101100",
  19973=>"001001010",
  19974=>"000000100",
  19975=>"101100001",
  19976=>"000000001",
  19977=>"010100111",
  19978=>"010011011",
  19979=>"111111100",
  19980=>"011100001",
  19981=>"100001011",
  19982=>"110000000",
  19983=>"001001110",
  19984=>"110001001",
  19985=>"110001000",
  19986=>"011101101",
  19987=>"100010111",
  19988=>"001111101",
  19989=>"100010100",
  19990=>"001101001",
  19991=>"111011011",
  19992=>"111000101",
  19993=>"000101001",
  19994=>"011001101",
  19995=>"111000101",
  19996=>"110100011",
  19997=>"111111011",
  19998=>"000010000",
  19999=>"111010001",
  20000=>"111010001",
  20001=>"110011011",
  20002=>"101001011",
  20003=>"110111011",
  20004=>"001110010",
  20005=>"000101101",
  20006=>"110110100",
  20007=>"100010011",
  20008=>"101100100",
  20009=>"111100001",
  20010=>"100110100",
  20011=>"101000000",
  20012=>"100110010",
  20013=>"100101110",
  20014=>"011011000",
  20015=>"010101100",
  20016=>"011100010",
  20017=>"110110000",
  20018=>"101011000",
  20019=>"101001100",
  20020=>"000111010",
  20021=>"110011011",
  20022=>"100000100",
  20023=>"010101110",
  20024=>"011111111",
  20025=>"111010010",
  20026=>"110100010",
  20027=>"111011001",
  20028=>"001100110",
  20029=>"010001110",
  20030=>"010100001",
  20031=>"110010101",
  20032=>"101001010",
  20033=>"111111010",
  20034=>"111010111",
  20035=>"110101011",
  20036=>"100011101",
  20037=>"101111000",
  20038=>"110000100",
  20039=>"110000001",
  20040=>"001001111",
  20041=>"011110010",
  20042=>"011101100",
  20043=>"011100001",
  20044=>"010000101",
  20045=>"000001001",
  20046=>"000001001",
  20047=>"110010011",
  20048=>"111011000",
  20049=>"001010011",
  20050=>"000011001",
  20051=>"111101101",
  20052=>"010111100",
  20053=>"000000100",
  20054=>"010000110",
  20055=>"001110010",
  20056=>"010101010",
  20057=>"101010010",
  20058=>"110101111",
  20059=>"101001111",
  20060=>"000011111",
  20061=>"101100110",
  20062=>"101001000",
  20063=>"000010110",
  20064=>"010101111",
  20065=>"100110100",
  20066=>"101010010",
  20067=>"110110010",
  20068=>"001111011",
  20069=>"111001010",
  20070=>"000111011",
  20071=>"010000000",
  20072=>"010100111",
  20073=>"010101001",
  20074=>"000100110",
  20075=>"001100000",
  20076=>"011001010",
  20077=>"100000011",
  20078=>"010100001",
  20079=>"101110111",
  20080=>"101101101",
  20081=>"111011101",
  20082=>"011100000",
  20083=>"000011100",
  20084=>"000000011",
  20085=>"100010100",
  20086=>"011001000",
  20087=>"011100010",
  20088=>"010000000",
  20089=>"000100010",
  20090=>"010110111",
  20091=>"110000000",
  20092=>"111111010",
  20093=>"010001111",
  20094=>"100001010",
  20095=>"000110011",
  20096=>"010000011",
  20097=>"100001100",
  20098=>"000110110",
  20099=>"011011101",
  20100=>"000101111",
  20101=>"100000010",
  20102=>"100110110",
  20103=>"010011000",
  20104=>"000011111",
  20105=>"100010000",
  20106=>"111001001",
  20107=>"011001011",
  20108=>"101010000",
  20109=>"000001000",
  20110=>"011011011",
  20111=>"001101100",
  20112=>"100110010",
  20113=>"000101010",
  20114=>"110101011",
  20115=>"110100111",
  20116=>"001110001",
  20117=>"110000100",
  20118=>"000101100",
  20119=>"011000001",
  20120=>"001100011",
  20121=>"010101111",
  20122=>"110101110",
  20123=>"101111011",
  20124=>"010000110",
  20125=>"110011110",
  20126=>"000100001",
  20127=>"001110011",
  20128=>"011100100",
  20129=>"101111000",
  20130=>"010011111",
  20131=>"010101011",
  20132=>"000000000",
  20133=>"110000000",
  20134=>"100000110",
  20135=>"010001110",
  20136=>"011011110",
  20137=>"000001100",
  20138=>"100001010",
  20139=>"100011011",
  20140=>"111110000",
  20141=>"111101100",
  20142=>"111010011",
  20143=>"001010101",
  20144=>"000101010",
  20145=>"011010011",
  20146=>"101111011",
  20147=>"111110100",
  20148=>"001101010",
  20149=>"100010000",
  20150=>"011100010",
  20151=>"000011011",
  20152=>"011001101",
  20153=>"000000011",
  20154=>"000001111",
  20155=>"010100101",
  20156=>"100000111",
  20157=>"011000111",
  20158=>"110000100",
  20159=>"101111111",
  20160=>"000100111",
  20161=>"110011010",
  20162=>"100111001",
  20163=>"011010111",
  20164=>"111111100",
  20165=>"001000010",
  20166=>"111011101",
  20167=>"101100010",
  20168=>"100011101",
  20169=>"000000110",
  20170=>"011101010",
  20171=>"111111111",
  20172=>"111010001",
  20173=>"101101001",
  20174=>"010010100",
  20175=>"100001011",
  20176=>"110000111",
  20177=>"100010001",
  20178=>"100111101",
  20179=>"100110110",
  20180=>"011011101",
  20181=>"101111111",
  20182=>"100001100",
  20183=>"100000011",
  20184=>"001101010",
  20185=>"010001010",
  20186=>"101001001",
  20187=>"110110101",
  20188=>"110010000",
  20189=>"011110010",
  20190=>"001111111",
  20191=>"011110110",
  20192=>"101000001",
  20193=>"011110111",
  20194=>"101110001",
  20195=>"111011101",
  20196=>"100111001",
  20197=>"100101111",
  20198=>"111011111",
  20199=>"010001000",
  20200=>"011011001",
  20201=>"100110110",
  20202=>"111100001",
  20203=>"001011111",
  20204=>"100100111",
  20205=>"011000010",
  20206=>"100001010",
  20207=>"000100110",
  20208=>"110111101",
  20209=>"001011000",
  20210=>"101000000",
  20211=>"000100110",
  20212=>"010111010",
  20213=>"101000101",
  20214=>"000110010",
  20215=>"110011000",
  20216=>"000101101",
  20217=>"101110110",
  20218=>"010001011",
  20219=>"000101111",
  20220=>"011100011",
  20221=>"101100011",
  20222=>"010010001",
  20223=>"010001010",
  20224=>"101010001",
  20225=>"011010011",
  20226=>"111011111",
  20227=>"101011000",
  20228=>"100101001",
  20229=>"110000001",
  20230=>"010001110",
  20231=>"010010100",
  20232=>"110011110",
  20233=>"111111110",
  20234=>"000000110",
  20235=>"111001010",
  20236=>"010101010",
  20237=>"010100110",
  20238=>"001000011",
  20239=>"101010011",
  20240=>"101010001",
  20241=>"100101100",
  20242=>"010010110",
  20243=>"011010111",
  20244=>"010110001",
  20245=>"010001100",
  20246=>"010101000",
  20247=>"110110111",
  20248=>"010000011",
  20249=>"000100011",
  20250=>"101010111",
  20251=>"100100110",
  20252=>"111101000",
  20253=>"001100110",
  20254=>"001011000",
  20255=>"111110000",
  20256=>"011001001",
  20257=>"110100001",
  20258=>"010011010",
  20259=>"100001101",
  20260=>"101011101",
  20261=>"111110111",
  20262=>"110100000",
  20263=>"101111011",
  20264=>"110111000",
  20265=>"000001110",
  20266=>"101001101",
  20267=>"110111001",
  20268=>"011110100",
  20269=>"111111100",
  20270=>"011010001",
  20271=>"010110100",
  20272=>"111010110",
  20273=>"100110001",
  20274=>"010010011",
  20275=>"000000101",
  20276=>"000011111",
  20277=>"110111111",
  20278=>"111101011",
  20279=>"000010100",
  20280=>"100011100",
  20281=>"101010100",
  20282=>"010000000",
  20283=>"101111100",
  20284=>"011001111",
  20285=>"000001000",
  20286=>"000011110",
  20287=>"000100011",
  20288=>"100100110",
  20289=>"111111111",
  20290=>"001011100",
  20291=>"101000101",
  20292=>"001011110",
  20293=>"100101011",
  20294=>"101010101",
  20295=>"101001000",
  20296=>"100011001",
  20297=>"000100000",
  20298=>"001001111",
  20299=>"110010100",
  20300=>"010011100",
  20301=>"010101001",
  20302=>"101010101",
  20303=>"011010100",
  20304=>"000000100",
  20305=>"100000111",
  20306=>"111111101",
  20307=>"001001100",
  20308=>"101010010",
  20309=>"011011001",
  20310=>"000100011",
  20311=>"011011010",
  20312=>"001010001",
  20313=>"011111100",
  20314=>"110011001",
  20315=>"001111111",
  20316=>"101100011",
  20317=>"110011001",
  20318=>"000110101",
  20319=>"011001010",
  20320=>"110001000",
  20321=>"101000011",
  20322=>"110100100",
  20323=>"100101111",
  20324=>"100010001",
  20325=>"011011011",
  20326=>"000111110",
  20327=>"100001101",
  20328=>"000111101",
  20329=>"010001111",
  20330=>"010001000",
  20331=>"101110101",
  20332=>"110001101",
  20333=>"000110001",
  20334=>"100001010",
  20335=>"011011001",
  20336=>"111100110",
  20337=>"000010110",
  20338=>"110010101",
  20339=>"011001111",
  20340=>"011001000",
  20341=>"010101101",
  20342=>"001111011",
  20343=>"111001011",
  20344=>"100111100",
  20345=>"010001110",
  20346=>"111110000",
  20347=>"000000011",
  20348=>"000010110",
  20349=>"011001110",
  20350=>"001000100",
  20351=>"010011000",
  20352=>"010110001",
  20353=>"110001011",
  20354=>"111000100",
  20355=>"011010100",
  20356=>"100001110",
  20357=>"001111111",
  20358=>"101010110",
  20359=>"110101111",
  20360=>"101111111",
  20361=>"111001011",
  20362=>"101110111",
  20363=>"110000011",
  20364=>"010100000",
  20365=>"001110101",
  20366=>"100011100",
  20367=>"100101001",
  20368=>"000101101",
  20369=>"110110000",
  20370=>"010001000",
  20371=>"110101011",
  20372=>"010110111",
  20373=>"010010001",
  20374=>"000001001",
  20375=>"001100000",
  20376=>"011010000",
  20377=>"010110101",
  20378=>"111000000",
  20379=>"010110000",
  20380=>"001110110",
  20381=>"111000011",
  20382=>"001110000",
  20383=>"010101010",
  20384=>"101000101",
  20385=>"000010100",
  20386=>"001110110",
  20387=>"001001111",
  20388=>"110011100",
  20389=>"011000101",
  20390=>"101101110",
  20391=>"101111110",
  20392=>"011110000",
  20393=>"011011010",
  20394=>"100010011",
  20395=>"101010100",
  20396=>"010100111",
  20397=>"111111111",
  20398=>"000111100",
  20399=>"111001110",
  20400=>"101100000",
  20401=>"010110111",
  20402=>"100101100",
  20403=>"010100001",
  20404=>"111011001",
  20405=>"010011001",
  20406=>"001000001",
  20407=>"011110110",
  20408=>"010000001",
  20409=>"011110101",
  20410=>"111110010",
  20411=>"011001001",
  20412=>"110001011",
  20413=>"000100101",
  20414=>"011010100",
  20415=>"101100101",
  20416=>"110101101",
  20417=>"110101111",
  20418=>"100001111",
  20419=>"010110100",
  20420=>"100110110",
  20421=>"100010101",
  20422=>"001000110",
  20423=>"110110000",
  20424=>"011000010",
  20425=>"010110000",
  20426=>"101111011",
  20427=>"010101000",
  20428=>"100101111",
  20429=>"001011001",
  20430=>"111111111",
  20431=>"000110011",
  20432=>"111011000",
  20433=>"011000100",
  20434=>"011010011",
  20435=>"111100001",
  20436=>"111010011",
  20437=>"011111111",
  20438=>"101101001",
  20439=>"010000111",
  20440=>"011011110",
  20441=>"101101111",
  20442=>"000011011",
  20443=>"001000010",
  20444=>"100110010",
  20445=>"000110111",
  20446=>"110000101",
  20447=>"000101101",
  20448=>"011111010",
  20449=>"010000010",
  20450=>"111100011",
  20451=>"010110010",
  20452=>"111000001",
  20453=>"010100100",
  20454=>"101101000",
  20455=>"110101001",
  20456=>"001011111",
  20457=>"101100100",
  20458=>"000110101",
  20459=>"101000000",
  20460=>"111111111",
  20461=>"101110010",
  20462=>"111000010",
  20463=>"011010000",
  20464=>"001100100",
  20465=>"011000111",
  20466=>"010000111",
  20467=>"001100011",
  20468=>"010011000",
  20469=>"111001000",
  20470=>"101111010",
  20471=>"101111101",
  20472=>"101011101",
  20473=>"110100111",
  20474=>"001011100",
  20475=>"001101001",
  20476=>"100111100",
  20477=>"000110100",
  20478=>"011110110",
  20479=>"100101110",
  20480=>"011111000",
  20481=>"111100000",
  20482=>"111101011",
  20483=>"001100011",
  20484=>"001001100",
  20485=>"010000000",
  20486=>"000000101",
  20487=>"011111110",
  20488=>"100101110",
  20489=>"100000001",
  20490=>"100000100",
  20491=>"111111110",
  20492=>"110110011",
  20493=>"001011110",
  20494=>"100101110",
  20495=>"010110011",
  20496=>"011110101",
  20497=>"110111110",
  20498=>"100000101",
  20499=>"100110110",
  20500=>"100010111",
  20501=>"110101010",
  20502=>"000001111",
  20503=>"100101001",
  20504=>"000011000",
  20505=>"010011111",
  20506=>"101010110",
  20507=>"011001101",
  20508=>"010101011",
  20509=>"111000011",
  20510=>"001110001",
  20511=>"011111011",
  20512=>"011101110",
  20513=>"111100010",
  20514=>"100001011",
  20515=>"110110011",
  20516=>"100010100",
  20517=>"011111110",
  20518=>"100000110",
  20519=>"101000100",
  20520=>"111100111",
  20521=>"100101001",
  20522=>"001001011",
  20523=>"001011111",
  20524=>"111010110",
  20525=>"001011111",
  20526=>"110001001",
  20527=>"011010101",
  20528=>"110101001",
  20529=>"000010100",
  20530=>"110011110",
  20531=>"010000100",
  20532=>"111011010",
  20533=>"001110000",
  20534=>"100111011",
  20535=>"000011110",
  20536=>"101010100",
  20537=>"011101100",
  20538=>"000000000",
  20539=>"100010110",
  20540=>"011100011",
  20541=>"001001011",
  20542=>"110111110",
  20543=>"010010010",
  20544=>"111000101",
  20545=>"010011100",
  20546=>"111110010",
  20547=>"001001000",
  20548=>"000110100",
  20549=>"100001000",
  20550=>"010110101",
  20551=>"100111000",
  20552=>"011101011",
  20553=>"010001011",
  20554=>"100000110",
  20555=>"111000111",
  20556=>"100001001",
  20557=>"000001000",
  20558=>"111111011",
  20559=>"111011011",
  20560=>"100100110",
  20561=>"100100110",
  20562=>"101110101",
  20563=>"000001110",
  20564=>"100000000",
  20565=>"100011101",
  20566=>"000111011",
  20567=>"100100000",
  20568=>"100001110",
  20569=>"100100000",
  20570=>"001110011",
  20571=>"101110010",
  20572=>"100100001",
  20573=>"110110100",
  20574=>"001000101",
  20575=>"001100100",
  20576=>"000010001",
  20577=>"010011101",
  20578=>"010000111",
  20579=>"101100010",
  20580=>"010000011",
  20581=>"101111111",
  20582=>"000011010",
  20583=>"000111000",
  20584=>"111011101",
  20585=>"000110010",
  20586=>"110001000",
  20587=>"011000000",
  20588=>"100101100",
  20589=>"001101111",
  20590=>"000111011",
  20591=>"100110011",
  20592=>"111110101",
  20593=>"010101110",
  20594=>"010110010",
  20595=>"111000100",
  20596=>"011110000",
  20597=>"101101100",
  20598=>"001010110",
  20599=>"011100100",
  20600=>"101001010",
  20601=>"011000001",
  20602=>"001111001",
  20603=>"110110110",
  20604=>"100100100",
  20605=>"100001000",
  20606=>"101100111",
  20607=>"010100001",
  20608=>"011000111",
  20609=>"010111011",
  20610=>"000010111",
  20611=>"001111101",
  20612=>"000010001",
  20613=>"111010010",
  20614=>"011100000",
  20615=>"111001111",
  20616=>"110010001",
  20617=>"001000000",
  20618=>"111101011",
  20619=>"000110100",
  20620=>"111111010",
  20621=>"011100000",
  20622=>"111011001",
  20623=>"011010001",
  20624=>"000010000",
  20625=>"001010011",
  20626=>"101111111",
  20627=>"111110001",
  20628=>"100000110",
  20629=>"110000000",
  20630=>"011110101",
  20631=>"111001101",
  20632=>"100100111",
  20633=>"000001101",
  20634=>"110100111",
  20635=>"000010111",
  20636=>"100111000",
  20637=>"000100111",
  20638=>"100001000",
  20639=>"100011101",
  20640=>"011010110",
  20641=>"011101010",
  20642=>"101011011",
  20643=>"001110110",
  20644=>"110010111",
  20645=>"110000111",
  20646=>"011010111",
  20647=>"111011011",
  20648=>"010111110",
  20649=>"011001001",
  20650=>"000000000",
  20651=>"011111110",
  20652=>"110010001",
  20653=>"100110110",
  20654=>"001000010",
  20655=>"010111111",
  20656=>"011101110",
  20657=>"010101011",
  20658=>"111010001",
  20659=>"000100000",
  20660=>"000101110",
  20661=>"000100110",
  20662=>"100101000",
  20663=>"011101010",
  20664=>"101110010",
  20665=>"101101000",
  20666=>"001010010",
  20667=>"010011010",
  20668=>"001010001",
  20669=>"011110000",
  20670=>"101010010",
  20671=>"101001001",
  20672=>"111001110",
  20673=>"100110101",
  20674=>"001000110",
  20675=>"011000010",
  20676=>"110000100",
  20677=>"101001101",
  20678=>"100000101",
  20679=>"000101101",
  20680=>"010010100",
  20681=>"100010010",
  20682=>"011000011",
  20683=>"101111100",
  20684=>"100110101",
  20685=>"101111001",
  20686=>"001100111",
  20687=>"001001001",
  20688=>"011000000",
  20689=>"010011111",
  20690=>"110001000",
  20691=>"110110000",
  20692=>"101110010",
  20693=>"100011111",
  20694=>"101110010",
  20695=>"000111000",
  20696=>"110100111",
  20697=>"111010011",
  20698=>"111101010",
  20699=>"001100101",
  20700=>"100100111",
  20701=>"110110001",
  20702=>"100001100",
  20703=>"010010111",
  20704=>"100100011",
  20705=>"101100001",
  20706=>"011001100",
  20707=>"111110000",
  20708=>"100010000",
  20709=>"111011001",
  20710=>"011111000",
  20711=>"000111100",
  20712=>"101010000",
  20713=>"110010001",
  20714=>"101010111",
  20715=>"001100000",
  20716=>"110110100",
  20717=>"100101011",
  20718=>"000001011",
  20719=>"111101000",
  20720=>"010010111",
  20721=>"110100010",
  20722=>"100110001",
  20723=>"011011001",
  20724=>"000010011",
  20725=>"111011001",
  20726=>"100101000",
  20727=>"001001110",
  20728=>"110100001",
  20729=>"001011001",
  20730=>"111101010",
  20731=>"001101100",
  20732=>"111111011",
  20733=>"100110011",
  20734=>"100000111",
  20735=>"111010000",
  20736=>"110100111",
  20737=>"011111111",
  20738=>"011110011",
  20739=>"110111100",
  20740=>"100101001",
  20741=>"111110101",
  20742=>"011100010",
  20743=>"100101110",
  20744=>"100011111",
  20745=>"000100101",
  20746=>"100111010",
  20747=>"010010110",
  20748=>"011011010",
  20749=>"000110110",
  20750=>"110010001",
  20751=>"010101000",
  20752=>"011010011",
  20753=>"111111011",
  20754=>"011000000",
  20755=>"011100100",
  20756=>"111100001",
  20757=>"100111011",
  20758=>"101011011",
  20759=>"111101111",
  20760=>"100101010",
  20761=>"000111101",
  20762=>"100111001",
  20763=>"111110101",
  20764=>"110001011",
  20765=>"001111110",
  20766=>"110100101",
  20767=>"000100010",
  20768=>"001101101",
  20769=>"100100011",
  20770=>"011111011",
  20771=>"100111111",
  20772=>"101110010",
  20773=>"000001011",
  20774=>"111001100",
  20775=>"100111011",
  20776=>"100101100",
  20777=>"101100111",
  20778=>"011101011",
  20779=>"010011100",
  20780=>"000101011",
  20781=>"000101110",
  20782=>"101110011",
  20783=>"110001111",
  20784=>"000000000",
  20785=>"010011000",
  20786=>"100111110",
  20787=>"001100110",
  20788=>"000100011",
  20789=>"010001011",
  20790=>"111111000",
  20791=>"110110111",
  20792=>"000001000",
  20793=>"011010100",
  20794=>"101101101",
  20795=>"010100110",
  20796=>"011001010",
  20797=>"100010111",
  20798=>"111011000",
  20799=>"111001101",
  20800=>"010010110",
  20801=>"001101110",
  20802=>"100101001",
  20803=>"100010100",
  20804=>"000001000",
  20805=>"111101010",
  20806=>"010000111",
  20807=>"000000010",
  20808=>"010010010",
  20809=>"000000001",
  20810=>"111111100",
  20811=>"101010001",
  20812=>"100100000",
  20813=>"100000111",
  20814=>"101111000",
  20815=>"110010111",
  20816=>"101010000",
  20817=>"101111101",
  20818=>"101010000",
  20819=>"010111110",
  20820=>"101011101",
  20821=>"111110110",
  20822=>"001101000",
  20823=>"111000111",
  20824=>"110011111",
  20825=>"010011110",
  20826=>"010000011",
  20827=>"111001100",
  20828=>"011111000",
  20829=>"110000101",
  20830=>"110111100",
  20831=>"010010000",
  20832=>"110010000",
  20833=>"011110000",
  20834=>"000001001",
  20835=>"100000101",
  20836=>"001011010",
  20837=>"001101011",
  20838=>"000101001",
  20839=>"011010101",
  20840=>"011101111",
  20841=>"110000010",
  20842=>"010101001",
  20843=>"100110000",
  20844=>"101101010",
  20845=>"101101100",
  20846=>"100100011",
  20847=>"010010001",
  20848=>"011000001",
  20849=>"001000010",
  20850=>"110000111",
  20851=>"011000101",
  20852=>"110110010",
  20853=>"000110100",
  20854=>"011001101",
  20855=>"111110100",
  20856=>"000000110",
  20857=>"110110110",
  20858=>"000101111",
  20859=>"000011001",
  20860=>"111111101",
  20861=>"110011000",
  20862=>"011110000",
  20863=>"100101111",
  20864=>"111100010",
  20865=>"111000110",
  20866=>"010011101",
  20867=>"001001000",
  20868=>"100001101",
  20869=>"101110110",
  20870=>"011001100",
  20871=>"000000001",
  20872=>"111110001",
  20873=>"101110010",
  20874=>"011000110",
  20875=>"001110110",
  20876=>"011101010",
  20877=>"000110000",
  20878=>"011000000",
  20879=>"110111010",
  20880=>"010101010",
  20881=>"000000000",
  20882=>"010000100",
  20883=>"101111101",
  20884=>"011011100",
  20885=>"001010001",
  20886=>"101100100",
  20887=>"000001001",
  20888=>"111011101",
  20889=>"110100000",
  20890=>"111101000",
  20891=>"110110010",
  20892=>"010111000",
  20893=>"000001111",
  20894=>"010110101",
  20895=>"010010001",
  20896=>"000101101",
  20897=>"000010110",
  20898=>"100110011",
  20899=>"011110001",
  20900=>"100111101",
  20901=>"000010000",
  20902=>"101000000",
  20903=>"111000111",
  20904=>"010100000",
  20905=>"101100001",
  20906=>"000110001",
  20907=>"011000101",
  20908=>"001011001",
  20909=>"011010100",
  20910=>"011100110",
  20911=>"010110110",
  20912=>"011000011",
  20913=>"101111000",
  20914=>"100001100",
  20915=>"000100011",
  20916=>"110001000",
  20917=>"111011010",
  20918=>"111011100",
  20919=>"001100001",
  20920=>"000001011",
  20921=>"010010000",
  20922=>"110110110",
  20923=>"001000011",
  20924=>"010100011",
  20925=>"110110010",
  20926=>"011111011",
  20927=>"001001011",
  20928=>"101010110",
  20929=>"110101000",
  20930=>"000010111",
  20931=>"001111001",
  20932=>"100000011",
  20933=>"001100011",
  20934=>"101011101",
  20935=>"111010100",
  20936=>"110010001",
  20937=>"000011010",
  20938=>"101010110",
  20939=>"000011011",
  20940=>"110001001",
  20941=>"000001111",
  20942=>"011011100",
  20943=>"100000100",
  20944=>"111010111",
  20945=>"111010000",
  20946=>"111000010",
  20947=>"110001101",
  20948=>"011100011",
  20949=>"011011110",
  20950=>"100101001",
  20951=>"111010001",
  20952=>"011110110",
  20953=>"101110110",
  20954=>"111110100",
  20955=>"000110001",
  20956=>"110101111",
  20957=>"000010111",
  20958=>"110111110",
  20959=>"011110010",
  20960=>"110111010",
  20961=>"010000000",
  20962=>"000100000",
  20963=>"101000011",
  20964=>"110000001",
  20965=>"110110000",
  20966=>"111101010",
  20967=>"000011001",
  20968=>"100101111",
  20969=>"001111000",
  20970=>"110100110",
  20971=>"010111111",
  20972=>"000100100",
  20973=>"010100100",
  20974=>"111100010",
  20975=>"101010101",
  20976=>"000010011",
  20977=>"001100101",
  20978=>"010000001",
  20979=>"110010100",
  20980=>"101010010",
  20981=>"001000011",
  20982=>"111101111",
  20983=>"001000010",
  20984=>"111100101",
  20985=>"010111100",
  20986=>"101101110",
  20987=>"111101101",
  20988=>"000110111",
  20989=>"101101010",
  20990=>"000000000",
  20991=>"101101011",
  20992=>"010101111",
  20993=>"101110100",
  20994=>"100010000",
  20995=>"110111110",
  20996=>"010000100",
  20997=>"100000010",
  20998=>"111010000",
  20999=>"010001000",
  21000=>"000101001",
  21001=>"110100101",
  21002=>"111011101",
  21003=>"010001101",
  21004=>"101011111",
  21005=>"100101001",
  21006=>"110010101",
  21007=>"100011010",
  21008=>"010000110",
  21009=>"011010010",
  21010=>"101111000",
  21011=>"100010001",
  21012=>"110100101",
  21013=>"010011011",
  21014=>"010110111",
  21015=>"101011111",
  21016=>"000000010",
  21017=>"011111000",
  21018=>"001001100",
  21019=>"010000011",
  21020=>"111111011",
  21021=>"110001101",
  21022=>"101011010",
  21023=>"101011101",
  21024=>"101001001",
  21025=>"101011110",
  21026=>"101111101",
  21027=>"110110011",
  21028=>"010110110",
  21029=>"110000101",
  21030=>"111101110",
  21031=>"000000011",
  21032=>"110110111",
  21033=>"101100001",
  21034=>"001011111",
  21035=>"101011100",
  21036=>"101000111",
  21037=>"101101010",
  21038=>"100110001",
  21039=>"110110111",
  21040=>"000100101",
  21041=>"000101111",
  21042=>"111111111",
  21043=>"010110011",
  21044=>"101001101",
  21045=>"011111100",
  21046=>"100011111",
  21047=>"110000011",
  21048=>"101111011",
  21049=>"100001011",
  21050=>"000100101",
  21051=>"001100001",
  21052=>"000101100",
  21053=>"111001001",
  21054=>"100101111",
  21055=>"000000010",
  21056=>"000011010",
  21057=>"000000010",
  21058=>"000010011",
  21059=>"000111001",
  21060=>"101100000",
  21061=>"010100101",
  21062=>"000001100",
  21063=>"111000101",
  21064=>"100010000",
  21065=>"100101010",
  21066=>"010101011",
  21067=>"000000010",
  21068=>"101111001",
  21069=>"101100101",
  21070=>"110001000",
  21071=>"101001101",
  21072=>"001011000",
  21073=>"000010000",
  21074=>"101001001",
  21075=>"001100111",
  21076=>"010000100",
  21077=>"010101110",
  21078=>"011011010",
  21079=>"011111010",
  21080=>"111110011",
  21081=>"110111111",
  21082=>"000000001",
  21083=>"101111001",
  21084=>"010000000",
  21085=>"100100010",
  21086=>"101010000",
  21087=>"111000001",
  21088=>"010000101",
  21089=>"010000000",
  21090=>"111111111",
  21091=>"100101000",
  21092=>"111010110",
  21093=>"010001000",
  21094=>"011000101",
  21095=>"001001011",
  21096=>"000011110",
  21097=>"101110111",
  21098=>"001110101",
  21099=>"000111100",
  21100=>"100010111",
  21101=>"001101001",
  21102=>"111100111",
  21103=>"010100110",
  21104=>"011111000",
  21105=>"010110110",
  21106=>"110111110",
  21107=>"000011111",
  21108=>"111101000",
  21109=>"111111111",
  21110=>"111110001",
  21111=>"010110111",
  21112=>"011100101",
  21113=>"110100000",
  21114=>"110010100",
  21115=>"100111100",
  21116=>"100010011",
  21117=>"000110101",
  21118=>"100000001",
  21119=>"011011101",
  21120=>"000011000",
  21121=>"111010001",
  21122=>"100010001",
  21123=>"001000101",
  21124=>"010101011",
  21125=>"101100111",
  21126=>"110000001",
  21127=>"010011001",
  21128=>"010101111",
  21129=>"100100010",
  21130=>"101010011",
  21131=>"001100001",
  21132=>"110110011",
  21133=>"111101110",
  21134=>"110010011",
  21135=>"011011101",
  21136=>"110111010",
  21137=>"100010000",
  21138=>"100101110",
  21139=>"101000011",
  21140=>"001110010",
  21141=>"000100110",
  21142=>"100010100",
  21143=>"001010111",
  21144=>"110100100",
  21145=>"100111111",
  21146=>"111110110",
  21147=>"111111111",
  21148=>"010110001",
  21149=>"111100000",
  21150=>"010110001",
  21151=>"101101101",
  21152=>"101110000",
  21153=>"100010000",
  21154=>"111111101",
  21155=>"100000110",
  21156=>"000100011",
  21157=>"000110010",
  21158=>"011001001",
  21159=>"000001100",
  21160=>"101101011",
  21161=>"001000100",
  21162=>"110011100",
  21163=>"111011001",
  21164=>"011110011",
  21165=>"000011001",
  21166=>"101011101",
  21167=>"100001010",
  21168=>"001110000",
  21169=>"110110100",
  21170=>"010000011",
  21171=>"110000101",
  21172=>"010000011",
  21173=>"001111110",
  21174=>"011001010",
  21175=>"101000110",
  21176=>"110101100",
  21177=>"011011011",
  21178=>"010111010",
  21179=>"011101110",
  21180=>"110110100",
  21181=>"010110100",
  21182=>"100100111",
  21183=>"011000110",
  21184=>"101110000",
  21185=>"111110111",
  21186=>"101010000",
  21187=>"010111110",
  21188=>"100001001",
  21189=>"001010101",
  21190=>"000101101",
  21191=>"001101110",
  21192=>"110101100",
  21193=>"110100111",
  21194=>"111000010",
  21195=>"101000001",
  21196=>"101110101",
  21197=>"001110001",
  21198=>"001101000",
  21199=>"111011101",
  21200=>"000011110",
  21201=>"100001000",
  21202=>"101111000",
  21203=>"110101100",
  21204=>"001010101",
  21205=>"101011111",
  21206=>"010111000",
  21207=>"101001001",
  21208=>"001111101",
  21209=>"110000001",
  21210=>"100100100",
  21211=>"001001101",
  21212=>"101111100",
  21213=>"000001011",
  21214=>"100011110",
  21215=>"111001010",
  21216=>"101110000",
  21217=>"011000000",
  21218=>"100001110",
  21219=>"101111110",
  21220=>"101100101",
  21221=>"011111111",
  21222=>"000000010",
  21223=>"101000001",
  21224=>"001101110",
  21225=>"100001111",
  21226=>"011110100",
  21227=>"001101101",
  21228=>"101111100",
  21229=>"010101101",
  21230=>"110011110",
  21231=>"101111001",
  21232=>"101001000",
  21233=>"010011001",
  21234=>"010100101",
  21235=>"100000001",
  21236=>"101101101",
  21237=>"111001010",
  21238=>"100110111",
  21239=>"011111101",
  21240=>"001011001",
  21241=>"100100011",
  21242=>"011111100",
  21243=>"110101110",
  21244=>"111000100",
  21245=>"001011110",
  21246=>"010000101",
  21247=>"010011100",
  21248=>"111110100",
  21249=>"010101111",
  21250=>"011101101",
  21251=>"011100111",
  21252=>"101100011",
  21253=>"111110000",
  21254=>"001111011",
  21255=>"100010111",
  21256=>"110110001",
  21257=>"010000101",
  21258=>"010001001",
  21259=>"111011110",
  21260=>"111100110",
  21261=>"001000111",
  21262=>"001111101",
  21263=>"000010011",
  21264=>"000111010",
  21265=>"001100100",
  21266=>"010111000",
  21267=>"001010001",
  21268=>"010000001",
  21269=>"011001101",
  21270=>"001010010",
  21271=>"100000101",
  21272=>"000001010",
  21273=>"110001001",
  21274=>"101100011",
  21275=>"110101101",
  21276=>"101111001",
  21277=>"110110001",
  21278=>"010000000",
  21279=>"111101101",
  21280=>"101011010",
  21281=>"001101010",
  21282=>"100100100",
  21283=>"010101100",
  21284=>"010111110",
  21285=>"010100100",
  21286=>"110010100",
  21287=>"101010010",
  21288=>"111011001",
  21289=>"010101111",
  21290=>"101000101",
  21291=>"000101001",
  21292=>"100100111",
  21293=>"001000000",
  21294=>"000101000",
  21295=>"100101100",
  21296=>"010110110",
  21297=>"101100000",
  21298=>"100011101",
  21299=>"001001011",
  21300=>"111000001",
  21301=>"111111111",
  21302=>"000011011",
  21303=>"001110001",
  21304=>"100101110",
  21305=>"011100001",
  21306=>"011010110",
  21307=>"010110111",
  21308=>"111100110",
  21309=>"101100010",
  21310=>"111111100",
  21311=>"100011011",
  21312=>"001100101",
  21313=>"111000100",
  21314=>"011110100",
  21315=>"111100101",
  21316=>"101100101",
  21317=>"011011011",
  21318=>"000001000",
  21319=>"101001011",
  21320=>"111110100",
  21321=>"000111000",
  21322=>"101001101",
  21323=>"001100001",
  21324=>"110000001",
  21325=>"001000101",
  21326=>"111110011",
  21327=>"100000000",
  21328=>"101100101",
  21329=>"001111101",
  21330=>"000111001",
  21331=>"001000100",
  21332=>"110010010",
  21333=>"100111001",
  21334=>"101010111",
  21335=>"011000000",
  21336=>"100000000",
  21337=>"001110011",
  21338=>"010100000",
  21339=>"010111110",
  21340=>"000100110",
  21341=>"111001111",
  21342=>"010000011",
  21343=>"001110110",
  21344=>"100100110",
  21345=>"010011011",
  21346=>"001001100",
  21347=>"010010100",
  21348=>"100001110",
  21349=>"010010110",
  21350=>"011111110",
  21351=>"011111000",
  21352=>"011101101",
  21353=>"010110011",
  21354=>"110010100",
  21355=>"110000010",
  21356=>"110111001",
  21357=>"011000100",
  21358=>"100110011",
  21359=>"011000000",
  21360=>"011110001",
  21361=>"110100001",
  21362=>"001101111",
  21363=>"100001011",
  21364=>"001011000",
  21365=>"000011010",
  21366=>"100100010",
  21367=>"100110101",
  21368=>"000010100",
  21369=>"111110011",
  21370=>"010011001",
  21371=>"101000110",
  21372=>"010010001",
  21373=>"000101111",
  21374=>"101011100",
  21375=>"110101000",
  21376=>"010001110",
  21377=>"011000110",
  21378=>"100001001",
  21379=>"001010100",
  21380=>"110100101",
  21381=>"100101010",
  21382=>"100011001",
  21383=>"101011100",
  21384=>"111110101",
  21385=>"011001111",
  21386=>"010001110",
  21387=>"111011010",
  21388=>"101110011",
  21389=>"011100000",
  21390=>"001011001",
  21391=>"100111100",
  21392=>"100111001",
  21393=>"010110000",
  21394=>"000110001",
  21395=>"100101010",
  21396=>"111100011",
  21397=>"101101001",
  21398=>"000011011",
  21399=>"011010101",
  21400=>"000110111",
  21401=>"111001101",
  21402=>"000000111",
  21403=>"110110010",
  21404=>"010000111",
  21405=>"111011110",
  21406=>"011100000",
  21407=>"100011111",
  21408=>"001011000",
  21409=>"001001101",
  21410=>"000110111",
  21411=>"101110011",
  21412=>"100100100",
  21413=>"100111111",
  21414=>"101111000",
  21415=>"000001101",
  21416=>"100011000",
  21417=>"011110010",
  21418=>"001000111",
  21419=>"110100110",
  21420=>"001001000",
  21421=>"000100001",
  21422=>"100011000",
  21423=>"101100100",
  21424=>"000011000",
  21425=>"111000100",
  21426=>"010100100",
  21427=>"010100000",
  21428=>"000110010",
  21429=>"111111011",
  21430=>"100110111",
  21431=>"011100011",
  21432=>"101110100",
  21433=>"011001101",
  21434=>"100000010",
  21435=>"011101110",
  21436=>"101001100",
  21437=>"111011010",
  21438=>"101001101",
  21439=>"010111010",
  21440=>"011110000",
  21441=>"010010110",
  21442=>"001100000",
  21443=>"110111011",
  21444=>"111011010",
  21445=>"110001100",
  21446=>"000001011",
  21447=>"010100111",
  21448=>"001110111",
  21449=>"011011101",
  21450=>"111010111",
  21451=>"000110100",
  21452=>"001100010",
  21453=>"100100001",
  21454=>"011110010",
  21455=>"011110110",
  21456=>"100001010",
  21457=>"111101010",
  21458=>"101010001",
  21459=>"001001110",
  21460=>"100111100",
  21461=>"000100011",
  21462=>"011000111",
  21463=>"011101010",
  21464=>"001000001",
  21465=>"011111101",
  21466=>"010101000",
  21467=>"011110001",
  21468=>"110111011",
  21469=>"111011100",
  21470=>"110101110",
  21471=>"100110101",
  21472=>"101001001",
  21473=>"101111000",
  21474=>"101101011",
  21475=>"010001111",
  21476=>"110110001",
  21477=>"010000100",
  21478=>"110111100",
  21479=>"100000011",
  21480=>"010011010",
  21481=>"010011011",
  21482=>"000010001",
  21483=>"000011011",
  21484=>"001101100",
  21485=>"101100110",
  21486=>"000011000",
  21487=>"000111101",
  21488=>"000010001",
  21489=>"001010111",
  21490=>"001100110",
  21491=>"000001101",
  21492=>"100111111",
  21493=>"100001010",
  21494=>"111101010",
  21495=>"110011110",
  21496=>"000110001",
  21497=>"011000101",
  21498=>"100110001",
  21499=>"111001011",
  21500=>"000000100",
  21501=>"010101001",
  21502=>"011001111",
  21503=>"011001100",
  21504=>"111110111",
  21505=>"001110110",
  21506=>"111001010",
  21507=>"111110010",
  21508=>"111110111",
  21509=>"111000111",
  21510=>"001001000",
  21511=>"110111001",
  21512=>"101110011",
  21513=>"111110101",
  21514=>"000000111",
  21515=>"100110000",
  21516=>"111101000",
  21517=>"110111001",
  21518=>"100001010",
  21519=>"000101110",
  21520=>"000010100",
  21521=>"001110010",
  21522=>"101010100",
  21523=>"111111111",
  21524=>"110101010",
  21525=>"101101100",
  21526=>"110100110",
  21527=>"101010011",
  21528=>"100011111",
  21529=>"101101001",
  21530=>"000011100",
  21531=>"011000111",
  21532=>"010001110",
  21533=>"110000010",
  21534=>"110001000",
  21535=>"010001111",
  21536=>"001011111",
  21537=>"000000110",
  21538=>"011101100",
  21539=>"111011011",
  21540=>"101110001",
  21541=>"101010011",
  21542=>"101111101",
  21543=>"000100101",
  21544=>"000100010",
  21545=>"011101001",
  21546=>"010010101",
  21547=>"111110011",
  21548=>"100100101",
  21549=>"110011111",
  21550=>"110111000",
  21551=>"110000100",
  21552=>"010100110",
  21553=>"100000011",
  21554=>"100111010",
  21555=>"000001100",
  21556=>"001110110",
  21557=>"100110110",
  21558=>"001111000",
  21559=>"010000000",
  21560=>"000000010",
  21561=>"110100101",
  21562=>"001101011",
  21563=>"110100011",
  21564=>"101110010",
  21565=>"011111110",
  21566=>"011100001",
  21567=>"101110010",
  21568=>"000000000",
  21569=>"100101000",
  21570=>"000001011",
  21571=>"001110111",
  21572=>"000110111",
  21573=>"111011101",
  21574=>"001111100",
  21575=>"000111001",
  21576=>"000000000",
  21577=>"000010000",
  21578=>"101100111",
  21579=>"100010110",
  21580=>"000000001",
  21581=>"110110100",
  21582=>"100110101",
  21583=>"011000100",
  21584=>"110101100",
  21585=>"000010110",
  21586=>"000000110",
  21587=>"101000001",
  21588=>"011001111",
  21589=>"011011110",
  21590=>"110101110",
  21591=>"100001001",
  21592=>"101001101",
  21593=>"111000001",
  21594=>"111110100",
  21595=>"111100010",
  21596=>"011110111",
  21597=>"100100111",
  21598=>"010100100",
  21599=>"110011111",
  21600=>"110111101",
  21601=>"111100100",
  21602=>"111010000",
  21603=>"000001010",
  21604=>"011110010",
  21605=>"111111010",
  21606=>"100111011",
  21607=>"101001101",
  21608=>"010011100",
  21609=>"010001100",
  21610=>"000001000",
  21611=>"111011010",
  21612=>"110011010",
  21613=>"110011101",
  21614=>"100010100",
  21615=>"100101110",
  21616=>"110001010",
  21617=>"101010011",
  21618=>"010010100",
  21619=>"101101101",
  21620=>"101000010",
  21621=>"011011011",
  21622=>"001111111",
  21623=>"100100000",
  21624=>"000000010",
  21625=>"011101101",
  21626=>"111111101",
  21627=>"010001110",
  21628=>"100010111",
  21629=>"000111101",
  21630=>"110000111",
  21631=>"000101001",
  21632=>"101011000",
  21633=>"100110110",
  21634=>"110110000",
  21635=>"000110010",
  21636=>"010111100",
  21637=>"100001010",
  21638=>"000101000",
  21639=>"010001010",
  21640=>"111011111",
  21641=>"001001100",
  21642=>"001000001",
  21643=>"001110100",
  21644=>"001111010",
  21645=>"010101000",
  21646=>"010111111",
  21647=>"101110101",
  21648=>"110010100",
  21649=>"011011111",
  21650=>"110010111",
  21651=>"110011111",
  21652=>"000111010",
  21653=>"101010010",
  21654=>"001010011",
  21655=>"111100100",
  21656=>"100100010",
  21657=>"011000011",
  21658=>"101111011",
  21659=>"011100010",
  21660=>"111000011",
  21661=>"000110000",
  21662=>"111110110",
  21663=>"110000110",
  21664=>"000111111",
  21665=>"101000110",
  21666=>"001000000",
  21667=>"100001110",
  21668=>"110011011",
  21669=>"100101111",
  21670=>"110100010",
  21671=>"100110011",
  21672=>"010001000",
  21673=>"111011001",
  21674=>"000111110",
  21675=>"110001100",
  21676=>"110101110",
  21677=>"000011110",
  21678=>"000010101",
  21679=>"010101100",
  21680=>"011011101",
  21681=>"001010111",
  21682=>"101000010",
  21683=>"010101111",
  21684=>"111000111",
  21685=>"001111000",
  21686=>"010001100",
  21687=>"011101101",
  21688=>"100100000",
  21689=>"111101100",
  21690=>"100101101",
  21691=>"000001011",
  21692=>"010110000",
  21693=>"000001000",
  21694=>"011010010",
  21695=>"100101010",
  21696=>"001001101",
  21697=>"011111110",
  21698=>"100001100",
  21699=>"001000110",
  21700=>"101111001",
  21701=>"001101100",
  21702=>"000000101",
  21703=>"100000010",
  21704=>"101001010",
  21705=>"011001011",
  21706=>"110001101",
  21707=>"101101010",
  21708=>"011111000",
  21709=>"110111001",
  21710=>"110101100",
  21711=>"011001001",
  21712=>"011010010",
  21713=>"110110010",
  21714=>"101110100",
  21715=>"010011001",
  21716=>"010111000",
  21717=>"011101110",
  21718=>"001111001",
  21719=>"001110101",
  21720=>"100111110",
  21721=>"001100000",
  21722=>"011111100",
  21723=>"110100001",
  21724=>"010001010",
  21725=>"001100001",
  21726=>"010111010",
  21727=>"000100000",
  21728=>"100000101",
  21729=>"110111101",
  21730=>"001101101",
  21731=>"000100000",
  21732=>"001100111",
  21733=>"101010100",
  21734=>"101001011",
  21735=>"110011111",
  21736=>"100001011",
  21737=>"010101001",
  21738=>"110000010",
  21739=>"000100011",
  21740=>"000010000",
  21741=>"011100011",
  21742=>"111010011",
  21743=>"111000101",
  21744=>"010011011",
  21745=>"111010011",
  21746=>"111000111",
  21747=>"011111000",
  21748=>"100110001",
  21749=>"000011110",
  21750=>"011101111",
  21751=>"100010110",
  21752=>"000111011",
  21753=>"110100101",
  21754=>"001111111",
  21755=>"100100001",
  21756=>"011101001",
  21757=>"100010111",
  21758=>"011101000",
  21759=>"011010111",
  21760=>"000010001",
  21761=>"100110011",
  21762=>"011011011",
  21763=>"010000000",
  21764=>"010001110",
  21765=>"100000011",
  21766=>"111111011",
  21767=>"100110011",
  21768=>"000011101",
  21769=>"100100010",
  21770=>"011001000",
  21771=>"011110001",
  21772=>"110100001",
  21773=>"011011110",
  21774=>"000110100",
  21775=>"110000101",
  21776=>"111000100",
  21777=>"110100011",
  21778=>"100100011",
  21779=>"010111010",
  21780=>"010000101",
  21781=>"101111011",
  21782=>"001111001",
  21783=>"011010101",
  21784=>"011110000",
  21785=>"101101000",
  21786=>"011111101",
  21787=>"111110101",
  21788=>"000000001",
  21789=>"001000100",
  21790=>"111011101",
  21791=>"001001100",
  21792=>"001111110",
  21793=>"010111010",
  21794=>"010100101",
  21795=>"000001100",
  21796=>"110101110",
  21797=>"110101111",
  21798=>"101111110",
  21799=>"010101101",
  21800=>"101000010",
  21801=>"101100011",
  21802=>"111011001",
  21803=>"110110011",
  21804=>"011011011",
  21805=>"111010000",
  21806=>"010010001",
  21807=>"100100011",
  21808=>"100011000",
  21809=>"000001000",
  21810=>"111101110",
  21811=>"000110000",
  21812=>"001111110",
  21813=>"000111110",
  21814=>"010010111",
  21815=>"000111000",
  21816=>"010001100",
  21817=>"100110001",
  21818=>"010011100",
  21819=>"011000011",
  21820=>"100111010",
  21821=>"111010001",
  21822=>"010001001",
  21823=>"100000000",
  21824=>"010001011",
  21825=>"011011001",
  21826=>"000011001",
  21827=>"010101110",
  21828=>"011001011",
  21829=>"111100101",
  21830=>"110010000",
  21831=>"010011000",
  21832=>"101000110",
  21833=>"111100000",
  21834=>"010101001",
  21835=>"011100000",
  21836=>"101000110",
  21837=>"011001110",
  21838=>"101010000",
  21839=>"110110110",
  21840=>"110000010",
  21841=>"011010101",
  21842=>"000111000",
  21843=>"011101101",
  21844=>"100001010",
  21845=>"010100100",
  21846=>"101100100",
  21847=>"101100000",
  21848=>"101101101",
  21849=>"001010011",
  21850=>"001000010",
  21851=>"110111101",
  21852=>"100100110",
  21853=>"011001111",
  21854=>"010010111",
  21855=>"000010001",
  21856=>"111101111",
  21857=>"010100001",
  21858=>"100101101",
  21859=>"001000111",
  21860=>"011111011",
  21861=>"010010010",
  21862=>"010101001",
  21863=>"011100101",
  21864=>"000100101",
  21865=>"111011101",
  21866=>"011111011",
  21867=>"001000100",
  21868=>"010110111",
  21869=>"010111000",
  21870=>"000011000",
  21871=>"010111111",
  21872=>"001110001",
  21873=>"000110010",
  21874=>"100100111",
  21875=>"111111011",
  21876=>"000000111",
  21877=>"001111110",
  21878=>"010101101",
  21879=>"101011011",
  21880=>"110111000",
  21881=>"100101100",
  21882=>"010001100",
  21883=>"011110001",
  21884=>"111001000",
  21885=>"110101011",
  21886=>"000000000",
  21887=>"101001001",
  21888=>"001000000",
  21889=>"000000001",
  21890=>"001010100",
  21891=>"011110100",
  21892=>"001000101",
  21893=>"111100000",
  21894=>"000101000",
  21895=>"010101010",
  21896=>"011000011",
  21897=>"100110100",
  21898=>"110100011",
  21899=>"011010100",
  21900=>"111000010",
  21901=>"000010000",
  21902=>"010101000",
  21903=>"101001001",
  21904=>"100111001",
  21905=>"010100000",
  21906=>"110000001",
  21907=>"110011110",
  21908=>"001111101",
  21909=>"010000100",
  21910=>"000000101",
  21911=>"000100110",
  21912=>"111000000",
  21913=>"011010100",
  21914=>"111101000",
  21915=>"010011100",
  21916=>"001100011",
  21917=>"100001000",
  21918=>"111010011",
  21919=>"010000110",
  21920=>"100110111",
  21921=>"001111000",
  21922=>"100001100",
  21923=>"101010011",
  21924=>"101111111",
  21925=>"001011100",
  21926=>"111111011",
  21927=>"000001011",
  21928=>"000111100",
  21929=>"111101110",
  21930=>"000011110",
  21931=>"101001000",
  21932=>"111011100",
  21933=>"101011010",
  21934=>"010000011",
  21935=>"101110011",
  21936=>"010000011",
  21937=>"101001110",
  21938=>"110000101",
  21939=>"001101010",
  21940=>"111110001",
  21941=>"010011100",
  21942=>"110111111",
  21943=>"000010000",
  21944=>"100010011",
  21945=>"001011000",
  21946=>"011101110",
  21947=>"001010111",
  21948=>"101101010",
  21949=>"011011001",
  21950=>"101001111",
  21951=>"101011010",
  21952=>"111011100",
  21953=>"111111111",
  21954=>"001011101",
  21955=>"110000101",
  21956=>"110101010",
  21957=>"101101011",
  21958=>"001100101",
  21959=>"100110001",
  21960=>"011011110",
  21961=>"100001100",
  21962=>"010011110",
  21963=>"011101100",
  21964=>"001101100",
  21965=>"110100110",
  21966=>"111011001",
  21967=>"100010010",
  21968=>"001000111",
  21969=>"011000001",
  21970=>"000001000",
  21971=>"101000100",
  21972=>"011000101",
  21973=>"101110010",
  21974=>"101110111",
  21975=>"111011011",
  21976=>"111010011",
  21977=>"011101101",
  21978=>"110011001",
  21979=>"001110011",
  21980=>"010000000",
  21981=>"010100110",
  21982=>"010010110",
  21983=>"111101000",
  21984=>"110110000",
  21985=>"100111011",
  21986=>"000100100",
  21987=>"001111101",
  21988=>"111000100",
  21989=>"001010101",
  21990=>"011100011",
  21991=>"111000010",
  21992=>"101011111",
  21993=>"111011010",
  21994=>"001101110",
  21995=>"011100010",
  21996=>"001100100",
  21997=>"110110000",
  21998=>"001000011",
  21999=>"001110110",
  22000=>"101011000",
  22001=>"111111010",
  22002=>"000011100",
  22003=>"110100100",
  22004=>"010001001",
  22005=>"011011100",
  22006=>"011100101",
  22007=>"001000110",
  22008=>"101000110",
  22009=>"100010100",
  22010=>"001001101",
  22011=>"111011110",
  22012=>"011000111",
  22013=>"110010110",
  22014=>"011011000",
  22015=>"000111010",
  22016=>"011100000",
  22017=>"111001111",
  22018=>"100101010",
  22019=>"111110111",
  22020=>"011000000",
  22021=>"001001110",
  22022=>"110111011",
  22023=>"000000000",
  22024=>"011000000",
  22025=>"000010100",
  22026=>"001000000",
  22027=>"111110100",
  22028=>"100000110",
  22029=>"100111101",
  22030=>"000011111",
  22031=>"010111111",
  22032=>"001000100",
  22033=>"110000000",
  22034=>"011110101",
  22035=>"001000011",
  22036=>"001111101",
  22037=>"010110010",
  22038=>"010100000",
  22039=>"111101001",
  22040=>"001110101",
  22041=>"001001101",
  22042=>"010001011",
  22043=>"000000001",
  22044=>"101110111",
  22045=>"110101101",
  22046=>"011110001",
  22047=>"110100111",
  22048=>"111000000",
  22049=>"101000011",
  22050=>"100111100",
  22051=>"100110011",
  22052=>"101011111",
  22053=>"101011101",
  22054=>"010010000",
  22055=>"101100001",
  22056=>"011111010",
  22057=>"010001000",
  22058=>"111000010",
  22059=>"101100001",
  22060=>"111111001",
  22061=>"101011101",
  22062=>"101010010",
  22063=>"100100110",
  22064=>"010110100",
  22065=>"010011010",
  22066=>"000010111",
  22067=>"101101000",
  22068=>"000110110",
  22069=>"010011101",
  22070=>"000100101",
  22071=>"000110001",
  22072=>"101111101",
  22073=>"010000100",
  22074=>"010111000",
  22075=>"101011011",
  22076=>"111101111",
  22077=>"001110000",
  22078=>"110110101",
  22079=>"001000001",
  22080=>"110101100",
  22081=>"011101011",
  22082=>"011010110",
  22083=>"010110110",
  22084=>"001100101",
  22085=>"000100111",
  22086=>"110000000",
  22087=>"100000010",
  22088=>"110101000",
  22089=>"010000110",
  22090=>"001001000",
  22091=>"010010100",
  22092=>"110010011",
  22093=>"100101100",
  22094=>"001100011",
  22095=>"011000000",
  22096=>"110001000",
  22097=>"000001000",
  22098=>"000100100",
  22099=>"011000111",
  22100=>"001110101",
  22101=>"001100100",
  22102=>"001101000",
  22103=>"110100101",
  22104=>"001011000",
  22105=>"011101001",
  22106=>"011110111",
  22107=>"101101010",
  22108=>"001000011",
  22109=>"000101001",
  22110=>"000011100",
  22111=>"111011000",
  22112=>"111110101",
  22113=>"101011100",
  22114=>"011011010",
  22115=>"011010011",
  22116=>"001110101",
  22117=>"101001100",
  22118=>"010111010",
  22119=>"100000000",
  22120=>"011001001",
  22121=>"100001011",
  22122=>"100011001",
  22123=>"101001110",
  22124=>"011111111",
  22125=>"110011111",
  22126=>"001110101",
  22127=>"100111101",
  22128=>"000101111",
  22129=>"100001000",
  22130=>"001111010",
  22131=>"001101101",
  22132=>"100011110",
  22133=>"011101001",
  22134=>"101011000",
  22135=>"100101000",
  22136=>"101001111",
  22137=>"100000110",
  22138=>"111110110",
  22139=>"111101100",
  22140=>"000010001",
  22141=>"100011100",
  22142=>"111100011",
  22143=>"010001101",
  22144=>"110110111",
  22145=>"111000100",
  22146=>"110100111",
  22147=>"000110111",
  22148=>"111110001",
  22149=>"111010111",
  22150=>"100011101",
  22151=>"000001111",
  22152=>"101010111",
  22153=>"010101010",
  22154=>"111111110",
  22155=>"011001111",
  22156=>"000100010",
  22157=>"000011001",
  22158=>"001011010",
  22159=>"011111111",
  22160=>"101001001",
  22161=>"010010110",
  22162=>"011010010",
  22163=>"001100000",
  22164=>"001010011",
  22165=>"110100110",
  22166=>"111100110",
  22167=>"100011111",
  22168=>"100110010",
  22169=>"111101101",
  22170=>"101100001",
  22171=>"101001111",
  22172=>"011001110",
  22173=>"001111001",
  22174=>"111101011",
  22175=>"010110100",
  22176=>"011000011",
  22177=>"111101011",
  22178=>"010000000",
  22179=>"011100100",
  22180=>"100111011",
  22181=>"010100010",
  22182=>"000111001",
  22183=>"110110010",
  22184=>"101010101",
  22185=>"110000111",
  22186=>"001011010",
  22187=>"011111000",
  22188=>"111010100",
  22189=>"100011010",
  22190=>"000000011",
  22191=>"100010111",
  22192=>"110100001",
  22193=>"111111000",
  22194=>"010100111",
  22195=>"010001011",
  22196=>"110100001",
  22197=>"101101000",
  22198=>"001101101",
  22199=>"110100111",
  22200=>"111111000",
  22201=>"010011001",
  22202=>"101111101",
  22203=>"100000011",
  22204=>"100001110",
  22205=>"001110101",
  22206=>"000100101",
  22207=>"011101000",
  22208=>"000100010",
  22209=>"101101111",
  22210=>"011000010",
  22211=>"000100110",
  22212=>"100111001",
  22213=>"101011011",
  22214=>"001011001",
  22215=>"100110110",
  22216=>"000010110",
  22217=>"110001101",
  22218=>"000010110",
  22219=>"001001011",
  22220=>"010000101",
  22221=>"111111001",
  22222=>"111111111",
  22223=>"001010100",
  22224=>"001010000",
  22225=>"011111011",
  22226=>"010101101",
  22227=>"111101100",
  22228=>"011000101",
  22229=>"111000100",
  22230=>"010100000",
  22231=>"011100111",
  22232=>"000100000",
  22233=>"001000100",
  22234=>"011111011",
  22235=>"011000100",
  22236=>"010111000",
  22237=>"010011101",
  22238=>"001111101",
  22239=>"010010000",
  22240=>"100001001",
  22241=>"000101101",
  22242=>"001101100",
  22243=>"101100001",
  22244=>"010110010",
  22245=>"101011011",
  22246=>"100001100",
  22247=>"001101101",
  22248=>"100101011",
  22249=>"101111110",
  22250=>"110010000",
  22251=>"111000111",
  22252=>"110000100",
  22253=>"000001100",
  22254=>"010110101",
  22255=>"111001110",
  22256=>"111001011",
  22257=>"010010011",
  22258=>"001111101",
  22259=>"000101000",
  22260=>"010111001",
  22261=>"011011011",
  22262=>"011100101",
  22263=>"100000000",
  22264=>"001011111",
  22265=>"101001001",
  22266=>"101100001",
  22267=>"101110110",
  22268=>"110000010",
  22269=>"101010000",
  22270=>"110001000",
  22271=>"111100011",
  22272=>"010010000",
  22273=>"011010000",
  22274=>"000110111",
  22275=>"011101100",
  22276=>"010011111",
  22277=>"101000111",
  22278=>"111101111",
  22279=>"000011110",
  22280=>"000101001",
  22281=>"011011001",
  22282=>"110101110",
  22283=>"000100011",
  22284=>"111111100",
  22285=>"101001101",
  22286=>"100110000",
  22287=>"110001010",
  22288=>"100011001",
  22289=>"110001000",
  22290=>"001110001",
  22291=>"100101000",
  22292=>"001000001",
  22293=>"010100110",
  22294=>"101011111",
  22295=>"000100001",
  22296=>"111111111",
  22297=>"001001100",
  22298=>"000000001",
  22299=>"111001011",
  22300=>"100100100",
  22301=>"001111010",
  22302=>"100111110",
  22303=>"101011000",
  22304=>"101111111",
  22305=>"010010100",
  22306=>"000000010",
  22307=>"100011110",
  22308=>"100000110",
  22309=>"000010000",
  22310=>"000111011",
  22311=>"000111001",
  22312=>"010011101",
  22313=>"111111011",
  22314=>"110111110",
  22315=>"010000111",
  22316=>"110011001",
  22317=>"100101010",
  22318=>"111000100",
  22319=>"101101010",
  22320=>"101011010",
  22321=>"000001111",
  22322=>"000100001",
  22323=>"001101001",
  22324=>"011101101",
  22325=>"010000111",
  22326=>"100100011",
  22327=>"010001110",
  22328=>"000010111",
  22329=>"111111101",
  22330=>"010100100",
  22331=>"110100000",
  22332=>"010000100",
  22333=>"011000111",
  22334=>"011111101",
  22335=>"000100110",
  22336=>"000100000",
  22337=>"100001110",
  22338=>"110111100",
  22339=>"011001110",
  22340=>"100011001",
  22341=>"001010101",
  22342=>"100000110",
  22343=>"100010100",
  22344=>"011011100",
  22345=>"100100101",
  22346=>"100000000",
  22347=>"110001101",
  22348=>"011010100",
  22349=>"001101000",
  22350=>"000000100",
  22351=>"010000010",
  22352=>"001111111",
  22353=>"011010000",
  22354=>"101011111",
  22355=>"011000101",
  22356=>"111000110",
  22357=>"001001000",
  22358=>"100100000",
  22359=>"101110100",
  22360=>"101000100",
  22361=>"011101111",
  22362=>"000111011",
  22363=>"111100110",
  22364=>"000110011",
  22365=>"101111000",
  22366=>"111111011",
  22367=>"000000010",
  22368=>"111110001",
  22369=>"111000111",
  22370=>"000101010",
  22371=>"110011001",
  22372=>"000001010",
  22373=>"000010111",
  22374=>"010111110",
  22375=>"111000111",
  22376=>"000111110",
  22377=>"000111111",
  22378=>"100100111",
  22379=>"101001110",
  22380=>"010111100",
  22381=>"000010101",
  22382=>"111001000",
  22383=>"100001111",
  22384=>"001110110",
  22385=>"101100100",
  22386=>"110010001",
  22387=>"100011000",
  22388=>"010001111",
  22389=>"110000001",
  22390=>"110000010",
  22391=>"010010100",
  22392=>"110110110",
  22393=>"101111010",
  22394=>"101110110",
  22395=>"011111000",
  22396=>"010110111",
  22397=>"010011100",
  22398=>"000101010",
  22399=>"010110110",
  22400=>"110101001",
  22401=>"111001011",
  22402=>"001010100",
  22403=>"111001000",
  22404=>"001110001",
  22405=>"100001010",
  22406=>"000000011",
  22407=>"111010101",
  22408=>"010110001",
  22409=>"001111001",
  22410=>"101110010",
  22411=>"001001000",
  22412=>"111111101",
  22413=>"011011100",
  22414=>"010001010",
  22415=>"001100100",
  22416=>"001000100",
  22417=>"101000111",
  22418=>"101101110",
  22419=>"010011101",
  22420=>"100100100",
  22421=>"110000001",
  22422=>"010010011",
  22423=>"110001111",
  22424=>"101101101",
  22425=>"011011010",
  22426=>"100000000",
  22427=>"100010011",
  22428=>"111110010",
  22429=>"100111001",
  22430=>"010010001",
  22431=>"100011000",
  22432=>"111101011",
  22433=>"110001000",
  22434=>"110111101",
  22435=>"100000100",
  22436=>"111001010",
  22437=>"111101010",
  22438=>"011100001",
  22439=>"100010101",
  22440=>"011100110",
  22441=>"101000101",
  22442=>"001110001",
  22443=>"000010110",
  22444=>"100100101",
  22445=>"111100100",
  22446=>"100100101",
  22447=>"100011011",
  22448=>"101000001",
  22449=>"001101110",
  22450=>"111111011",
  22451=>"100001110",
  22452=>"010101111",
  22453=>"001101010",
  22454=>"010010111",
  22455=>"111010101",
  22456=>"011011010",
  22457=>"111001001",
  22458=>"101000101",
  22459=>"011000010",
  22460=>"010010010",
  22461=>"000110010",
  22462=>"110110001",
  22463=>"100100000",
  22464=>"001010001",
  22465=>"111001110",
  22466=>"100001100",
  22467=>"011010010",
  22468=>"000100101",
  22469=>"010111110",
  22470=>"110110011",
  22471=>"101101101",
  22472=>"110010101",
  22473=>"111100000",
  22474=>"000000100",
  22475=>"000001010",
  22476=>"001101111",
  22477=>"000000000",
  22478=>"101110000",
  22479=>"010111111",
  22480=>"011011010",
  22481=>"001011110",
  22482=>"101000000",
  22483=>"111011100",
  22484=>"001010010",
  22485=>"000100000",
  22486=>"101111101",
  22487=>"010001000",
  22488=>"000111101",
  22489=>"101010010",
  22490=>"100010110",
  22491=>"111011111",
  22492=>"111001011",
  22493=>"111101110",
  22494=>"110001100",
  22495=>"100011110",
  22496=>"011011000",
  22497=>"010111101",
  22498=>"100100001",
  22499=>"110001001",
  22500=>"110000010",
  22501=>"001111011",
  22502=>"010010110",
  22503=>"101010000",
  22504=>"110110010",
  22505=>"111101011",
  22506=>"010000010",
  22507=>"101010100",
  22508=>"100100111",
  22509=>"111001111",
  22510=>"000111000",
  22511=>"111010011",
  22512=>"000110110",
  22513=>"110110000",
  22514=>"110010010",
  22515=>"001100010",
  22516=>"010111100",
  22517=>"110100011",
  22518=>"000101000",
  22519=>"001011001",
  22520=>"010011110",
  22521=>"110000000",
  22522=>"101010101",
  22523=>"111011010",
  22524=>"011101111",
  22525=>"111110010",
  22526=>"010100101",
  22527=>"001010101",
  22528=>"111111111",
  22529=>"010101000",
  22530=>"010000101",
  22531=>"001111111",
  22532=>"100011110",
  22533=>"000010110",
  22534=>"110111100",
  22535=>"010000010",
  22536=>"101010011",
  22537=>"000100011",
  22538=>"101010011",
  22539=>"101001100",
  22540=>"111110001",
  22541=>"111100000",
  22542=>"110100011",
  22543=>"101100100",
  22544=>"010010000",
  22545=>"101100011",
  22546=>"100111011",
  22547=>"100111010",
  22548=>"110100001",
  22549=>"101010110",
  22550=>"100001010",
  22551=>"000110101",
  22552=>"011000011",
  22553=>"111001101",
  22554=>"111011000",
  22555=>"001110111",
  22556=>"101100001",
  22557=>"011101100",
  22558=>"001110010",
  22559=>"011111101",
  22560=>"100101100",
  22561=>"010101000",
  22562=>"100110111",
  22563=>"101101100",
  22564=>"111111101",
  22565=>"000010110",
  22566=>"110000111",
  22567=>"101010100",
  22568=>"001011011",
  22569=>"100000011",
  22570=>"100000110",
  22571=>"001110000",
  22572=>"011011111",
  22573=>"010101100",
  22574=>"001000001",
  22575=>"010011010",
  22576=>"111110010",
  22577=>"111100101",
  22578=>"101000111",
  22579=>"010010100",
  22580=>"011101101",
  22581=>"100100001",
  22582=>"101000110",
  22583=>"001001010",
  22584=>"000101011",
  22585=>"100110111",
  22586=>"110100101",
  22587=>"101110111",
  22588=>"010010111",
  22589=>"101011111",
  22590=>"101110000",
  22591=>"011101110",
  22592=>"000100110",
  22593=>"001100101",
  22594=>"000010100",
  22595=>"000100101",
  22596=>"011010011",
  22597=>"101001000",
  22598=>"001110001",
  22599=>"001000010",
  22600=>"001101110",
  22601=>"101111110",
  22602=>"011110011",
  22603=>"100000110",
  22604=>"101101000",
  22605=>"100000101",
  22606=>"111111110",
  22607=>"001001010",
  22608=>"010111010",
  22609=>"111100011",
  22610=>"110000110",
  22611=>"111101010",
  22612=>"110000011",
  22613=>"111110011",
  22614=>"010000010",
  22615=>"100000000",
  22616=>"011011100",
  22617=>"010101010",
  22618=>"000010000",
  22619=>"111110100",
  22620=>"001100111",
  22621=>"000011000",
  22622=>"111101001",
  22623=>"111101000",
  22624=>"111110001",
  22625=>"111001101",
  22626=>"111000011",
  22627=>"001000100",
  22628=>"111101100",
  22629=>"000011000",
  22630=>"000100101",
  22631=>"100000101",
  22632=>"111111101",
  22633=>"101110010",
  22634=>"001100101",
  22635=>"000000110",
  22636=>"110101000",
  22637=>"100111110",
  22638=>"010100011",
  22639=>"111101111",
  22640=>"100001000",
  22641=>"010011110",
  22642=>"110101010",
  22643=>"111110010",
  22644=>"111100100",
  22645=>"110100010",
  22646=>"000000011",
  22647=>"010100000",
  22648=>"001000011",
  22649=>"001100000",
  22650=>"011101010",
  22651=>"101101100",
  22652=>"001110101",
  22653=>"100101101",
  22654=>"111001111",
  22655=>"110110111",
  22656=>"001101100",
  22657=>"101000100",
  22658=>"000001010",
  22659=>"010001010",
  22660=>"000011101",
  22661=>"110110110",
  22662=>"100010010",
  22663=>"011010100",
  22664=>"000011011",
  22665=>"110100001",
  22666=>"011011101",
  22667=>"011001111",
  22668=>"101110011",
  22669=>"011011010",
  22670=>"100110010",
  22671=>"010000001",
  22672=>"000010001",
  22673=>"101001111",
  22674=>"110000110",
  22675=>"110101000",
  22676=>"000000010",
  22677=>"110000111",
  22678=>"000000100",
  22679=>"110101000",
  22680=>"100011100",
  22681=>"101000101",
  22682=>"111000101",
  22683=>"101001111",
  22684=>"000010000",
  22685=>"010010110",
  22686=>"001110000",
  22687=>"011000100",
  22688=>"010000101",
  22689=>"101001101",
  22690=>"001111001",
  22691=>"100101110",
  22692=>"000001101",
  22693=>"001000010",
  22694=>"011111001",
  22695=>"101110010",
  22696=>"110100101",
  22697=>"011111111",
  22698=>"010001100",
  22699=>"110110001",
  22700=>"100111001",
  22701=>"010101010",
  22702=>"111001000",
  22703=>"101010100",
  22704=>"011011110",
  22705=>"011110011",
  22706=>"010010000",
  22707=>"011111110",
  22708=>"001011010",
  22709=>"111001101",
  22710=>"101011000",
  22711=>"011111001",
  22712=>"101101111",
  22713=>"100001110",
  22714=>"110000000",
  22715=>"110111111",
  22716=>"000101100",
  22717=>"001111000",
  22718=>"010101110",
  22719=>"110101011",
  22720=>"111111110",
  22721=>"011010100",
  22722=>"100111100",
  22723=>"101100000",
  22724=>"110011000",
  22725=>"111101101",
  22726=>"101110110",
  22727=>"110111011",
  22728=>"000100101",
  22729=>"001010010",
  22730=>"000100100",
  22731=>"111110011",
  22732=>"011101100",
  22733=>"110101011",
  22734=>"111110101",
  22735=>"100000101",
  22736=>"110011111",
  22737=>"101110011",
  22738=>"001100001",
  22739=>"011101001",
  22740=>"100100010",
  22741=>"010111011",
  22742=>"110000000",
  22743=>"100011111",
  22744=>"111010000",
  22745=>"110101010",
  22746=>"000010100",
  22747=>"101011110",
  22748=>"001111110",
  22749=>"111110001",
  22750=>"111101100",
  22751=>"000110100",
  22752=>"000000001",
  22753=>"101011111",
  22754=>"101010101",
  22755=>"100001100",
  22756=>"111001001",
  22757=>"000001011",
  22758=>"110000000",
  22759=>"000111001",
  22760=>"000001011",
  22761=>"111100111",
  22762=>"010001110",
  22763=>"010001001",
  22764=>"101101011",
  22765=>"000110100",
  22766=>"010100010",
  22767=>"100100000",
  22768=>"111110010",
  22769=>"111100011",
  22770=>"001000010",
  22771=>"000101001",
  22772=>"100000010",
  22773=>"110100000",
  22774=>"110111000",
  22775=>"010101001",
  22776=>"001011111",
  22777=>"100011001",
  22778=>"011011111",
  22779=>"010101111",
  22780=>"000110001",
  22781=>"110011111",
  22782=>"001001100",
  22783=>"111011011",
  22784=>"011000011",
  22785=>"011001010",
  22786=>"010011101",
  22787=>"001010111",
  22788=>"000110000",
  22789=>"101110110",
  22790=>"100110110",
  22791=>"010111111",
  22792=>"011110001",
  22793=>"000111100",
  22794=>"000000100",
  22795=>"000101011",
  22796=>"001001100",
  22797=>"011101101",
  22798=>"101100111",
  22799=>"000111110",
  22800=>"110010100",
  22801=>"010010000",
  22802=>"100010111",
  22803=>"101111010",
  22804=>"100010001",
  22805=>"010000100",
  22806=>"110100110",
  22807=>"011010110",
  22808=>"110110110",
  22809=>"100000010",
  22810=>"110110011",
  22811=>"100100011",
  22812=>"010100110",
  22813=>"010101111",
  22814=>"001011011",
  22815=>"111010110",
  22816=>"100110110",
  22817=>"000011010",
  22818=>"000011001",
  22819=>"011101011",
  22820=>"010100100",
  22821=>"011001011",
  22822=>"011000101",
  22823=>"101010001",
  22824=>"101111000",
  22825=>"010101000",
  22826=>"100011000",
  22827=>"000111000",
  22828=>"011000010",
  22829=>"001011001",
  22830=>"000011101",
  22831=>"010110010",
  22832=>"000100010",
  22833=>"001111000",
  22834=>"000101001",
  22835=>"000111110",
  22836=>"010101010",
  22837=>"010011110",
  22838=>"100101011",
  22839=>"110000010",
  22840=>"001001001",
  22841=>"001011001",
  22842=>"011011011",
  22843=>"001110101",
  22844=>"000000110",
  22845=>"100110011",
  22846=>"000000110",
  22847=>"011000011",
  22848=>"010000010",
  22849=>"010111111",
  22850=>"111010001",
  22851=>"000010001",
  22852=>"001100101",
  22853=>"010101111",
  22854=>"011100001",
  22855=>"111011000",
  22856=>"011111011",
  22857=>"000100100",
  22858=>"110111010",
  22859=>"000100010",
  22860=>"110011110",
  22861=>"110010001",
  22862=>"011111011",
  22863=>"001111100",
  22864=>"100101001",
  22865=>"111010101",
  22866=>"111111001",
  22867=>"110000111",
  22868=>"111000000",
  22869=>"111100111",
  22870=>"001111100",
  22871=>"011111110",
  22872=>"001000111",
  22873=>"000111011",
  22874=>"001101100",
  22875=>"110111001",
  22876=>"111010111",
  22877=>"111111011",
  22878=>"100011001",
  22879=>"000111101",
  22880=>"000100010",
  22881=>"010110011",
  22882=>"110111101",
  22883=>"001000100",
  22884=>"100010000",
  22885=>"111100001",
  22886=>"110100010",
  22887=>"000001110",
  22888=>"000011010",
  22889=>"011000001",
  22890=>"010111101",
  22891=>"100011010",
  22892=>"010100000",
  22893=>"011110001",
  22894=>"100111000",
  22895=>"001001000",
  22896=>"000100111",
  22897=>"011010110",
  22898=>"110111110",
  22899=>"101111000",
  22900=>"011101100",
  22901=>"011001110",
  22902=>"000000110",
  22903=>"011101100",
  22904=>"001001011",
  22905=>"101000010",
  22906=>"111101010",
  22907=>"100101110",
  22908=>"011010010",
  22909=>"111101101",
  22910=>"101001000",
  22911=>"011010100",
  22912=>"101000111",
  22913=>"001010100",
  22914=>"110111010",
  22915=>"111110111",
  22916=>"011111010",
  22917=>"111100111",
  22918=>"111010111",
  22919=>"000111010",
  22920=>"100000010",
  22921=>"011011100",
  22922=>"101000110",
  22923=>"101000111",
  22924=>"110001001",
  22925=>"111111010",
  22926=>"111100111",
  22927=>"000110111",
  22928=>"110010001",
  22929=>"011000001",
  22930=>"100000011",
  22931=>"101011010",
  22932=>"101100000",
  22933=>"101011111",
  22934=>"000001010",
  22935=>"100000010",
  22936=>"010110111",
  22937=>"001010000",
  22938=>"100001001",
  22939=>"111100100",
  22940=>"110100111",
  22941=>"001111110",
  22942=>"111100010",
  22943=>"101100101",
  22944=>"010001111",
  22945=>"100000000",
  22946=>"110011101",
  22947=>"110011111",
  22948=>"001100000",
  22949=>"101000001",
  22950=>"011111011",
  22951=>"011010100",
  22952=>"111000100",
  22953=>"000010000",
  22954=>"000011010",
  22955=>"011100110",
  22956=>"110000000",
  22957=>"100101000",
  22958=>"110000101",
  22959=>"001110100",
  22960=>"000101001",
  22961=>"100011000",
  22962=>"010010100",
  22963=>"100011100",
  22964=>"101001101",
  22965=>"111101100",
  22966=>"001101100",
  22967=>"101110000",
  22968=>"011001101",
  22969=>"100011101",
  22970=>"100000010",
  22971=>"000110011",
  22972=>"110100100",
  22973=>"000001001",
  22974=>"101111101",
  22975=>"010000000",
  22976=>"111110100",
  22977=>"010101010",
  22978=>"011001101",
  22979=>"101011000",
  22980=>"101101011",
  22981=>"011101001",
  22982=>"111100111",
  22983=>"110100010",
  22984=>"010010111",
  22985=>"111010001",
  22986=>"011000101",
  22987=>"011010110",
  22988=>"010111100",
  22989=>"100110001",
  22990=>"111000100",
  22991=>"000000011",
  22992=>"101110010",
  22993=>"010100000",
  22994=>"101101011",
  22995=>"011111101",
  22996=>"000011111",
  22997=>"101001111",
  22998=>"000100001",
  22999=>"100001010",
  23000=>"001100010",
  23001=>"100100000",
  23002=>"101001000",
  23003=>"101000001",
  23004=>"000000111",
  23005=>"111001110",
  23006=>"100001001",
  23007=>"001010111",
  23008=>"000000000",
  23009=>"000000101",
  23010=>"111010000",
  23011=>"000001001",
  23012=>"000010011",
  23013=>"101010010",
  23014=>"000111011",
  23015=>"000110010",
  23016=>"100001100",
  23017=>"000001100",
  23018=>"000100100",
  23019=>"010001101",
  23020=>"100001110",
  23021=>"000101111",
  23022=>"010001110",
  23023=>"010101100",
  23024=>"000001101",
  23025=>"000000110",
  23026=>"100101011",
  23027=>"000000111",
  23028=>"000010101",
  23029=>"110011001",
  23030=>"100100000",
  23031=>"011000011",
  23032=>"001111010",
  23033=>"100101100",
  23034=>"000110110",
  23035=>"110100100",
  23036=>"000010100",
  23037=>"010000011",
  23038=>"101001010",
  23039=>"111111110",
  23040=>"001101111",
  23041=>"100011001",
  23042=>"101100001",
  23043=>"001001110",
  23044=>"011111000",
  23045=>"111100111",
  23046=>"101111011",
  23047=>"000010000",
  23048=>"111111000",
  23049=>"011110011",
  23050=>"000001100",
  23051=>"100100011",
  23052=>"010001011",
  23053=>"010000001",
  23054=>"001010110",
  23055=>"000110100",
  23056=>"101010111",
  23057=>"001100110",
  23058=>"110010000",
  23059=>"000010010",
  23060=>"110010000",
  23061=>"010011011",
  23062=>"101101000",
  23063=>"100111001",
  23064=>"000100011",
  23065=>"011010001",
  23066=>"001100001",
  23067=>"001100000",
  23068=>"001011100",
  23069=>"111010010",
  23070=>"010010011",
  23071=>"010101101",
  23072=>"111110001",
  23073=>"110110100",
  23074=>"100010010",
  23075=>"000110011",
  23076=>"100011111",
  23077=>"001000010",
  23078=>"101110000",
  23079=>"010000000",
  23080=>"101000010",
  23081=>"001010011",
  23082=>"010110100",
  23083=>"001100111",
  23084=>"111110100",
  23085=>"101101010",
  23086=>"010111001",
  23087=>"110101101",
  23088=>"111100001",
  23089=>"100000111",
  23090=>"000100001",
  23091=>"001100101",
  23092=>"011110010",
  23093=>"000000001",
  23094=>"101000001",
  23095=>"110111111",
  23096=>"110111011",
  23097=>"100011000",
  23098=>"010101110",
  23099=>"111001100",
  23100=>"000010100",
  23101=>"101110011",
  23102=>"000110100",
  23103=>"011101100",
  23104=>"010001111",
  23105=>"001100000",
  23106=>"000000100",
  23107=>"010110001",
  23108=>"111101010",
  23109=>"111111111",
  23110=>"100111001",
  23111=>"001101011",
  23112=>"100110001",
  23113=>"100111110",
  23114=>"100001000",
  23115=>"111101010",
  23116=>"001001111",
  23117=>"110100011",
  23118=>"011011111",
  23119=>"111011111",
  23120=>"001001010",
  23121=>"101001001",
  23122=>"100101000",
  23123=>"000010011",
  23124=>"110001110",
  23125=>"101110111",
  23126=>"100110100",
  23127=>"101101111",
  23128=>"110101111",
  23129=>"010100001",
  23130=>"101010011",
  23131=>"101000110",
  23132=>"000011000",
  23133=>"110000000",
  23134=>"001101110",
  23135=>"100000010",
  23136=>"110000100",
  23137=>"000100110",
  23138=>"101000001",
  23139=>"100100000",
  23140=>"101101010",
  23141=>"111000000",
  23142=>"000111011",
  23143=>"010000110",
  23144=>"100111110",
  23145=>"100000001",
  23146=>"000010110",
  23147=>"110111110",
  23148=>"000101110",
  23149=>"000001101",
  23150=>"100110110",
  23151=>"110001000",
  23152=>"101101000",
  23153=>"010001000",
  23154=>"110011001",
  23155=>"101101101",
  23156=>"000011110",
  23157=>"111101010",
  23158=>"100000000",
  23159=>"110101110",
  23160=>"111100000",
  23161=>"101110001",
  23162=>"101101001",
  23163=>"010111111",
  23164=>"001001011",
  23165=>"001000100",
  23166=>"100010011",
  23167=>"111111101",
  23168=>"001011010",
  23169=>"010001101",
  23170=>"111100101",
  23171=>"000001001",
  23172=>"110011100",
  23173=>"011000101",
  23174=>"101110011",
  23175=>"000100001",
  23176=>"001010011",
  23177=>"001100110",
  23178=>"010100010",
  23179=>"001100111",
  23180=>"111111111",
  23181=>"001110101",
  23182=>"111011111",
  23183=>"000000110",
  23184=>"001101011",
  23185=>"110111111",
  23186=>"010011111",
  23187=>"101110100",
  23188=>"010101010",
  23189=>"000101100",
  23190=>"011010001",
  23191=>"011000001",
  23192=>"000000001",
  23193=>"110100111",
  23194=>"111111001",
  23195=>"110010001",
  23196=>"011011000",
  23197=>"001010011",
  23198=>"111101101",
  23199=>"001011100",
  23200=>"001010001",
  23201=>"110011111",
  23202=>"010001001",
  23203=>"111000111",
  23204=>"001110010",
  23205=>"011010011",
  23206=>"011000000",
  23207=>"000100010",
  23208=>"110111010",
  23209=>"000111110",
  23210=>"000001010",
  23211=>"000010000",
  23212=>"010110110",
  23213=>"101110011",
  23214=>"011001111",
  23215=>"001011000",
  23216=>"000110010",
  23217=>"111101111",
  23218=>"000100011",
  23219=>"000100100",
  23220=>"110110000",
  23221=>"111000101",
  23222=>"111111110",
  23223=>"000111101",
  23224=>"100110101",
  23225=>"111011000",
  23226=>"111101111",
  23227=>"001000100",
  23228=>"111010011",
  23229=>"101101111",
  23230=>"101000001",
  23231=>"010110101",
  23232=>"000111011",
  23233=>"011000110",
  23234=>"000100100",
  23235=>"100101011",
  23236=>"111000001",
  23237=>"110100101",
  23238=>"000100010",
  23239=>"111101001",
  23240=>"001011111",
  23241=>"001101111",
  23242=>"001001110",
  23243=>"100010000",
  23244=>"010000000",
  23245=>"010000100",
  23246=>"000111011",
  23247=>"101001011",
  23248=>"011001011",
  23249=>"110100010",
  23250=>"101011010",
  23251=>"111100110",
  23252=>"110001000",
  23253=>"111101101",
  23254=>"111110000",
  23255=>"010100111",
  23256=>"000011010",
  23257=>"001010111",
  23258=>"000100010",
  23259=>"100010000",
  23260=>"101110110",
  23261=>"101110001",
  23262=>"001010110",
  23263=>"100101101",
  23264=>"101100101",
  23265=>"000001110",
  23266=>"100100011",
  23267=>"001100001",
  23268=>"100100010",
  23269=>"101000101",
  23270=>"011111000",
  23271=>"110100000",
  23272=>"101100100",
  23273=>"001100001",
  23274=>"010010111",
  23275=>"010001100",
  23276=>"111011100",
  23277=>"010011000",
  23278=>"011111011",
  23279=>"010001011",
  23280=>"110111011",
  23281=>"101000000",
  23282=>"110111110",
  23283=>"110010110",
  23284=>"010010000",
  23285=>"101100001",
  23286=>"001111001",
  23287=>"010000010",
  23288=>"010011101",
  23289=>"000000100",
  23290=>"100000110",
  23291=>"110001000",
  23292=>"000011010",
  23293=>"010100011",
  23294=>"000011100",
  23295=>"101100111",
  23296=>"111000001",
  23297=>"000000011",
  23298=>"000110001",
  23299=>"101000101",
  23300=>"001111101",
  23301=>"100111100",
  23302=>"010011111",
  23303=>"111010000",
  23304=>"100001110",
  23305=>"100010110",
  23306=>"110000010",
  23307=>"001010000",
  23308=>"001110100",
  23309=>"110001100",
  23310=>"010010100",
  23311=>"110110110",
  23312=>"111110100",
  23313=>"010101101",
  23314=>"011011011",
  23315=>"010101010",
  23316=>"000110100",
  23317=>"001111110",
  23318=>"000100010",
  23319=>"011100011",
  23320=>"111101100",
  23321=>"011100101",
  23322=>"100001101",
  23323=>"101110000",
  23324=>"011111111",
  23325=>"101000101",
  23326=>"001101110",
  23327=>"111011001",
  23328=>"110000001",
  23329=>"100100000",
  23330=>"100010101",
  23331=>"001010001",
  23332=>"000010000",
  23333=>"000100101",
  23334=>"001111111",
  23335=>"011110111",
  23336=>"010000100",
  23337=>"001101111",
  23338=>"111010001",
  23339=>"000000011",
  23340=>"101111111",
  23341=>"001000001",
  23342=>"011101101",
  23343=>"110000001",
  23344=>"111101100",
  23345=>"111111010",
  23346=>"101000111",
  23347=>"110101000",
  23348=>"111000000",
  23349=>"000001001",
  23350=>"110001000",
  23351=>"101110011",
  23352=>"100001101",
  23353=>"000000011",
  23354=>"001110100",
  23355=>"010110000",
  23356=>"101010101",
  23357=>"101110101",
  23358=>"000100000",
  23359=>"001111001",
  23360=>"111010001",
  23361=>"011111010",
  23362=>"010111000",
  23363=>"011100111",
  23364=>"010100101",
  23365=>"100111001",
  23366=>"111011110",
  23367=>"010111010",
  23368=>"010101000",
  23369=>"111001111",
  23370=>"011110000",
  23371=>"011010111",
  23372=>"111010001",
  23373=>"110011011",
  23374=>"010101001",
  23375=>"110010010",
  23376=>"111110010",
  23377=>"011101111",
  23378=>"001001010",
  23379=>"101010001",
  23380=>"111111001",
  23381=>"111110111",
  23382=>"000101001",
  23383=>"110101010",
  23384=>"100110101",
  23385=>"111111110",
  23386=>"010111100",
  23387=>"001101001",
  23388=>"111000010",
  23389=>"011000000",
  23390=>"010000000",
  23391=>"011100110",
  23392=>"011010010",
  23393=>"101100111",
  23394=>"100101001",
  23395=>"000110000",
  23396=>"110010111",
  23397=>"101001111",
  23398=>"111001101",
  23399=>"111000000",
  23400=>"011000001",
  23401=>"111100101",
  23402=>"001000001",
  23403=>"001101010",
  23404=>"110010111",
  23405=>"010100100",
  23406=>"101110110",
  23407=>"011011110",
  23408=>"000111101",
  23409=>"010111100",
  23410=>"110110101",
  23411=>"000000111",
  23412=>"010001000",
  23413=>"010110100",
  23414=>"101001101",
  23415=>"111101111",
  23416=>"011101010",
  23417=>"110001111",
  23418=>"001001111",
  23419=>"000110110",
  23420=>"000001101",
  23421=>"111101100",
  23422=>"000001101",
  23423=>"111110110",
  23424=>"011001101",
  23425=>"110010100",
  23426=>"010011101",
  23427=>"011001010",
  23428=>"100001101",
  23429=>"011001000",
  23430=>"100100011",
  23431=>"010000010",
  23432=>"011111101",
  23433=>"001110000",
  23434=>"110001000",
  23435=>"000100101",
  23436=>"000000110",
  23437=>"001100110",
  23438=>"100000000",
  23439=>"001011010",
  23440=>"010110011",
  23441=>"101000001",
  23442=>"100010110",
  23443=>"101111001",
  23444=>"001000100",
  23445=>"100111110",
  23446=>"011001001",
  23447=>"100011010",
  23448=>"111111000",
  23449=>"010101001",
  23450=>"010111110",
  23451=>"111100000",
  23452=>"010010010",
  23453=>"001000011",
  23454=>"110100101",
  23455=>"010011101",
  23456=>"111011010",
  23457=>"011011110",
  23458=>"000010001",
  23459=>"100111000",
  23460=>"000010001",
  23461=>"100110011",
  23462=>"010010110",
  23463=>"111111111",
  23464=>"011000101",
  23465=>"000100110",
  23466=>"000110011",
  23467=>"111001000",
  23468=>"001110111",
  23469=>"111111001",
  23470=>"000001001",
  23471=>"000000000",
  23472=>"011100011",
  23473=>"100011001",
  23474=>"000100011",
  23475=>"010011110",
  23476=>"110110001",
  23477=>"101010011",
  23478=>"110100111",
  23479=>"100100101",
  23480=>"100111000",
  23481=>"111011101",
  23482=>"010011000",
  23483=>"000001010",
  23484=>"111101110",
  23485=>"010100110",
  23486=>"010000100",
  23487=>"111010110",
  23488=>"000000010",
  23489=>"111101110",
  23490=>"011111000",
  23491=>"000111001",
  23492=>"111111101",
  23493=>"111101111",
  23494=>"100011110",
  23495=>"000110011",
  23496=>"111001100",
  23497=>"011000000",
  23498=>"100010110",
  23499=>"111000000",
  23500=>"000000000",
  23501=>"010010111",
  23502=>"111000111",
  23503=>"000100001",
  23504=>"000100111",
  23505=>"001010011",
  23506=>"000010000",
  23507=>"101100011",
  23508=>"001100111",
  23509=>"111001100",
  23510=>"011111000",
  23511=>"111010110",
  23512=>"101101011",
  23513=>"001110001",
  23514=>"010010011",
  23515=>"010111101",
  23516=>"010110000",
  23517=>"100110010",
  23518=>"000101001",
  23519=>"110101010",
  23520=>"001010101",
  23521=>"001001000",
  23522=>"000111111",
  23523=>"110010110",
  23524=>"100101110",
  23525=>"110101010",
  23526=>"110011111",
  23527=>"000001100",
  23528=>"000100110",
  23529=>"100011110",
  23530=>"110000001",
  23531=>"000011101",
  23532=>"111000101",
  23533=>"000010101",
  23534=>"010111001",
  23535=>"100110111",
  23536=>"010110000",
  23537=>"110010111",
  23538=>"010111111",
  23539=>"010010011",
  23540=>"110011011",
  23541=>"110110110",
  23542=>"001110000",
  23543=>"101101110",
  23544=>"010001000",
  23545=>"011000000",
  23546=>"110000111",
  23547=>"100010000",
  23548=>"101101110",
  23549=>"011010010",
  23550=>"110000110",
  23551=>"110110111",
  23552=>"010111111",
  23553=>"110101111",
  23554=>"100100011",
  23555=>"101000010",
  23556=>"111100110",
  23557=>"101110110",
  23558=>"000011000",
  23559=>"110000000",
  23560=>"100110100",
  23561=>"101011000",
  23562=>"101100001",
  23563=>"010101101",
  23564=>"000000100",
  23565=>"010011101",
  23566=>"010010100",
  23567=>"001100101",
  23568=>"000011011",
  23569=>"110111101",
  23570=>"011110000",
  23571=>"011101101",
  23572=>"100000110",
  23573=>"010111110",
  23574=>"100010110",
  23575=>"000001010",
  23576=>"100000000",
  23577=>"000101100",
  23578=>"000111101",
  23579=>"100110001",
  23580=>"010011101",
  23581=>"100100111",
  23582=>"110010110",
  23583=>"010000001",
  23584=>"000000011",
  23585=>"011100010",
  23586=>"111101101",
  23587=>"110100001",
  23588=>"110010110",
  23589=>"111101010",
  23590=>"110010011",
  23591=>"111100101",
  23592=>"101000000",
  23593=>"111101010",
  23594=>"101000110",
  23595=>"011111000",
  23596=>"110111100",
  23597=>"010000000",
  23598=>"010111111",
  23599=>"001110111",
  23600=>"100111001",
  23601=>"101111000",
  23602=>"110001001",
  23603=>"100000101",
  23604=>"010110011",
  23605=>"110010101",
  23606=>"000000010",
  23607=>"101000000",
  23608=>"111100110",
  23609=>"111010101",
  23610=>"100011010",
  23611=>"000011000",
  23612=>"000101111",
  23613=>"001100010",
  23614=>"000010110",
  23615=>"011000000",
  23616=>"101000010",
  23617=>"111110011",
  23618=>"111111010",
  23619=>"011111000",
  23620=>"011110110",
  23621=>"011100011",
  23622=>"101001111",
  23623=>"100111111",
  23624=>"101010101",
  23625=>"111101101",
  23626=>"111100011",
  23627=>"100001101",
  23628=>"001100010",
  23629=>"010101100",
  23630=>"100010000",
  23631=>"101111111",
  23632=>"101101111",
  23633=>"110111111",
  23634=>"101100011",
  23635=>"000011001",
  23636=>"101000001",
  23637=>"000111111",
  23638=>"001011100",
  23639=>"001100110",
  23640=>"100010110",
  23641=>"101100011",
  23642=>"101000110",
  23643=>"101010001",
  23644=>"000111010",
  23645=>"111001110",
  23646=>"010100110",
  23647=>"110101110",
  23648=>"100110111",
  23649=>"001110011",
  23650=>"110100010",
  23651=>"111111111",
  23652=>"000111100",
  23653=>"111100101",
  23654=>"100011000",
  23655=>"110110111",
  23656=>"101100110",
  23657=>"011100010",
  23658=>"100100110",
  23659=>"111100000",
  23660=>"100001000",
  23661=>"100001101",
  23662=>"111110101",
  23663=>"110000110",
  23664=>"010001000",
  23665=>"100110011",
  23666=>"000101110",
  23667=>"001100010",
  23668=>"110010000",
  23669=>"111100110",
  23670=>"110110111",
  23671=>"101001010",
  23672=>"101011001",
  23673=>"011100100",
  23674=>"101110001",
  23675=>"110000110",
  23676=>"110010100",
  23677=>"101111001",
  23678=>"111001111",
  23679=>"111101101",
  23680=>"111001001",
  23681=>"010000001",
  23682=>"000100001",
  23683=>"001001010",
  23684=>"010001100",
  23685=>"111110000",
  23686=>"111111111",
  23687=>"000010011",
  23688=>"111110000",
  23689=>"010110001",
  23690=>"010011101",
  23691=>"111000011",
  23692=>"011101101",
  23693=>"000010010",
  23694=>"100011100",
  23695=>"101001110",
  23696=>"110010110",
  23697=>"101101011",
  23698=>"000001001",
  23699=>"110001000",
  23700=>"000000000",
  23701=>"001100100",
  23702=>"111100000",
  23703=>"011110000",
  23704=>"101001100",
  23705=>"101010101",
  23706=>"110011011",
  23707=>"011110011",
  23708=>"110100111",
  23709=>"110001011",
  23710=>"110110100",
  23711=>"000101000",
  23712=>"010001000",
  23713=>"111010100",
  23714=>"101000000",
  23715=>"101000011",
  23716=>"000000001",
  23717=>"100000001",
  23718=>"000111000",
  23719=>"101111001",
  23720=>"011100110",
  23721=>"010100010",
  23722=>"100000011",
  23723=>"100101100",
  23724=>"001001011",
  23725=>"101101001",
  23726=>"000011011",
  23727=>"100010111",
  23728=>"101011111",
  23729=>"011000101",
  23730=>"010011011",
  23731=>"010000101",
  23732=>"101010010",
  23733=>"110011010",
  23734=>"111101001",
  23735=>"101010100",
  23736=>"001100010",
  23737=>"101001000",
  23738=>"110011000",
  23739=>"111011101",
  23740=>"010000001",
  23741=>"010001101",
  23742=>"001010000",
  23743=>"010000110",
  23744=>"111101101",
  23745=>"100101110",
  23746=>"100011000",
  23747=>"101001001",
  23748=>"100010101",
  23749=>"010101100",
  23750=>"011011000",
  23751=>"001011000",
  23752=>"111111101",
  23753=>"101110010",
  23754=>"000000000",
  23755=>"101001111",
  23756=>"011010111",
  23757=>"100001010",
  23758=>"101001111",
  23759=>"000101101",
  23760=>"111111110",
  23761=>"101100001",
  23762=>"000011101",
  23763=>"101101000",
  23764=>"100111111",
  23765=>"111100001",
  23766=>"000110101",
  23767=>"000110010",
  23768=>"100000001",
  23769=>"111110101",
  23770=>"110000001",
  23771=>"001101000",
  23772=>"100011000",
  23773=>"101011100",
  23774=>"000010110",
  23775=>"111110011",
  23776=>"000000010",
  23777=>"000011000",
  23778=>"010100111",
  23779=>"101000010",
  23780=>"100001101",
  23781=>"010111000",
  23782=>"011000010",
  23783=>"001000001",
  23784=>"101001001",
  23785=>"011101110",
  23786=>"010000000",
  23787=>"011000001",
  23788=>"110010000",
  23789=>"010101110",
  23790=>"110110010",
  23791=>"101010110",
  23792=>"100001001",
  23793=>"011010100",
  23794=>"111001101",
  23795=>"110010011",
  23796=>"010011111",
  23797=>"010011011",
  23798=>"110111010",
  23799=>"101000000",
  23800=>"000101110",
  23801=>"101000011",
  23802=>"000100010",
  23803=>"000000000",
  23804=>"100000100",
  23805=>"010000011",
  23806=>"111111111",
  23807=>"011110110",
  23808=>"101100011",
  23809=>"011110000",
  23810=>"011110001",
  23811=>"101111011",
  23812=>"111011110",
  23813=>"000110101",
  23814=>"001111001",
  23815=>"000000100",
  23816=>"001000001",
  23817=>"111011011",
  23818=>"001110010",
  23819=>"011000011",
  23820=>"100010000",
  23821=>"001100111",
  23822=>"100010101",
  23823=>"100010000",
  23824=>"010111111",
  23825=>"111101101",
  23826=>"000010111",
  23827=>"000000110",
  23828=>"011010101",
  23829=>"100000010",
  23830=>"111110100",
  23831=>"000011011",
  23832=>"101000000",
  23833=>"110101011",
  23834=>"010010010",
  23835=>"011010010",
  23836=>"001111101",
  23837=>"001010101",
  23838=>"011101001",
  23839=>"001000011",
  23840=>"010101010",
  23841=>"000000100",
  23842=>"000010011",
  23843=>"011010011",
  23844=>"000110001",
  23845=>"100111011",
  23846=>"111101001",
  23847=>"110001110",
  23848=>"101110111",
  23849=>"111110101",
  23850=>"110001011",
  23851=>"000111000",
  23852=>"100101101",
  23853=>"000101111",
  23854=>"100100010",
  23855=>"100001000",
  23856=>"000001010",
  23857=>"010000101",
  23858=>"101101110",
  23859=>"000010011",
  23860=>"101000001",
  23861=>"110011100",
  23862=>"101100011",
  23863=>"010010111",
  23864=>"010000111",
  23865=>"111110111",
  23866=>"010000101",
  23867=>"000000011",
  23868=>"101100110",
  23869=>"101001100",
  23870=>"001110011",
  23871=>"111101011",
  23872=>"101101010",
  23873=>"011011010",
  23874=>"111010000",
  23875=>"100100111",
  23876=>"101101000",
  23877=>"011111111",
  23878=>"101101100",
  23879=>"000000110",
  23880=>"111011111",
  23881=>"010000001",
  23882=>"001011011",
  23883=>"000001001",
  23884=>"110110101",
  23885=>"110110111",
  23886=>"010101011",
  23887=>"110111100",
  23888=>"001111110",
  23889=>"000000100",
  23890=>"000000011",
  23891=>"101101000",
  23892=>"100000001",
  23893=>"101111011",
  23894=>"011110101",
  23895=>"000101111",
  23896=>"011000101",
  23897=>"101100001",
  23898=>"011000000",
  23899=>"111100001",
  23900=>"001011110",
  23901=>"011101100",
  23902=>"100010110",
  23903=>"111101001",
  23904=>"100101101",
  23905=>"000011100",
  23906=>"000010011",
  23907=>"001111011",
  23908=>"110010100",
  23909=>"110101101",
  23910=>"000001100",
  23911=>"100001100",
  23912=>"100110010",
  23913=>"100111000",
  23914=>"111000010",
  23915=>"111001111",
  23916=>"110011111",
  23917=>"011111111",
  23918=>"101001001",
  23919=>"101001011",
  23920=>"000110110",
  23921=>"001000101",
  23922=>"110100000",
  23923=>"100010110",
  23924=>"001110000",
  23925=>"101000010",
  23926=>"111001001",
  23927=>"100101111",
  23928=>"001111011",
  23929=>"001110010",
  23930=>"001100001",
  23931=>"110001100",
  23932=>"111101010",
  23933=>"110000000",
  23934=>"101000010",
  23935=>"010011101",
  23936=>"011101101",
  23937=>"000110011",
  23938=>"111001100",
  23939=>"110111001",
  23940=>"001001001",
  23941=>"000000110",
  23942=>"000000110",
  23943=>"111011110",
  23944=>"000000100",
  23945=>"111011101",
  23946=>"101010111",
  23947=>"001000011",
  23948=>"110000111",
  23949=>"101100000",
  23950=>"110100011",
  23951=>"001100101",
  23952=>"011001110",
  23953=>"000010000",
  23954=>"100101001",
  23955=>"101001100",
  23956=>"101011101",
  23957=>"110010101",
  23958=>"010111011",
  23959=>"010110001",
  23960=>"110001100",
  23961=>"011101000",
  23962=>"000010001",
  23963=>"011001010",
  23964=>"011111111",
  23965=>"011100100",
  23966=>"100011001",
  23967=>"000100011",
  23968=>"110010110",
  23969=>"111111010",
  23970=>"100110000",
  23971=>"000010010",
  23972=>"110100000",
  23973=>"101000011",
  23974=>"001100110",
  23975=>"101111000",
  23976=>"010111111",
  23977=>"100111000",
  23978=>"001000001",
  23979=>"000010111",
  23980=>"000000000",
  23981=>"010010011",
  23982=>"011011100",
  23983=>"101110011",
  23984=>"111100000",
  23985=>"111011011",
  23986=>"101101111",
  23987=>"010110100",
  23988=>"000011110",
  23989=>"011000010",
  23990=>"100111110",
  23991=>"101000001",
  23992=>"111000011",
  23993=>"000001011",
  23994=>"000100100",
  23995=>"011111111",
  23996=>"011101010",
  23997=>"011100001",
  23998=>"100001000",
  23999=>"011010111",
  24000=>"100100100",
  24001=>"101001001",
  24002=>"111011111",
  24003=>"010100110",
  24004=>"111001111",
  24005=>"100010011",
  24006=>"101100011",
  24007=>"011100011",
  24008=>"010000100",
  24009=>"101110110",
  24010=>"100001000",
  24011=>"010111001",
  24012=>"011110110",
  24013=>"100010000",
  24014=>"101010111",
  24015=>"100101111",
  24016=>"100001001",
  24017=>"111011111",
  24018=>"111100100",
  24019=>"110111111",
  24020=>"011110011",
  24021=>"000000011",
  24022=>"011111010",
  24023=>"101111000",
  24024=>"011010000",
  24025=>"010001100",
  24026=>"110101110",
  24027=>"011100000",
  24028=>"101100100",
  24029=>"110101111",
  24030=>"001010101",
  24031=>"010100000",
  24032=>"001111111",
  24033=>"001000111",
  24034=>"111100111",
  24035=>"010100010",
  24036=>"010011100",
  24037=>"101011000",
  24038=>"110110110",
  24039=>"101100000",
  24040=>"000000110",
  24041=>"000110001",
  24042=>"001011011",
  24043=>"010000111",
  24044=>"100010110",
  24045=>"111100111",
  24046=>"110011100",
  24047=>"111110110",
  24048=>"001011111",
  24049=>"010111001",
  24050=>"111010111",
  24051=>"001001111",
  24052=>"100000100",
  24053=>"101011011",
  24054=>"111011100",
  24055=>"111011100",
  24056=>"110011010",
  24057=>"100011001",
  24058=>"001011111",
  24059=>"110000111",
  24060=>"000001011",
  24061=>"001101101",
  24062=>"111110111",
  24063=>"110001011",
  24064=>"110000000",
  24065=>"111010111",
  24066=>"110001110",
  24067=>"011111000",
  24068=>"111110111",
  24069=>"001011001",
  24070=>"011100011",
  24071=>"110101100",
  24072=>"100100110",
  24073=>"100110001",
  24074=>"111001000",
  24075=>"010010000",
  24076=>"110011011",
  24077=>"000000010",
  24078=>"000000000",
  24079=>"001101011",
  24080=>"010101010",
  24081=>"000100101",
  24082=>"101101001",
  24083=>"100000100",
  24084=>"001010111",
  24085=>"001001110",
  24086=>"010011101",
  24087=>"110001111",
  24088=>"000000011",
  24089=>"100010111",
  24090=>"001001101",
  24091=>"111111110",
  24092=>"011110011",
  24093=>"000110110",
  24094=>"001000101",
  24095=>"001101001",
  24096=>"101100001",
  24097=>"000110011",
  24098=>"100100101",
  24099=>"101000111",
  24100=>"110000111",
  24101=>"011101110",
  24102=>"011111111",
  24103=>"011101111",
  24104=>"001011100",
  24105=>"110101100",
  24106=>"000000010",
  24107=>"110000101",
  24108=>"100111000",
  24109=>"010110111",
  24110=>"001110100",
  24111=>"011111110",
  24112=>"111001000",
  24113=>"110000111",
  24114=>"110010011",
  24115=>"111010111",
  24116=>"000000100",
  24117=>"101100101",
  24118=>"111001000",
  24119=>"111101110",
  24120=>"100011111",
  24121=>"101011001",
  24122=>"000100011",
  24123=>"000000010",
  24124=>"000000010",
  24125=>"000001001",
  24126=>"100011010",
  24127=>"110100100",
  24128=>"010111011",
  24129=>"111110001",
  24130=>"110000111",
  24131=>"111011001",
  24132=>"100000011",
  24133=>"110011000",
  24134=>"000011110",
  24135=>"100111111",
  24136=>"000010010",
  24137=>"100001011",
  24138=>"011001111",
  24139=>"000011000",
  24140=>"000101111",
  24141=>"101100001",
  24142=>"101010110",
  24143=>"000100010",
  24144=>"110111000",
  24145=>"101001010",
  24146=>"011010010",
  24147=>"000101010",
  24148=>"001111000",
  24149=>"100100011",
  24150=>"101000000",
  24151=>"010111001",
  24152=>"111001100",
  24153=>"111010011",
  24154=>"000101111",
  24155=>"011000000",
  24156=>"111100000",
  24157=>"001001000",
  24158=>"001110000",
  24159=>"100100011",
  24160=>"110101011",
  24161=>"000010011",
  24162=>"101100011",
  24163=>"111010001",
  24164=>"010001101",
  24165=>"110101100",
  24166=>"011001000",
  24167=>"101101011",
  24168=>"001101000",
  24169=>"010010001",
  24170=>"101001100",
  24171=>"001101010",
  24172=>"000101101",
  24173=>"101000111",
  24174=>"001111001",
  24175=>"011011100",
  24176=>"100011010",
  24177=>"011000001",
  24178=>"100101111",
  24179=>"100100000",
  24180=>"010101000",
  24181=>"000000000",
  24182=>"011000000",
  24183=>"111110001",
  24184=>"100000001",
  24185=>"001011000",
  24186=>"101000101",
  24187=>"000000001",
  24188=>"110010010",
  24189=>"001011111",
  24190=>"110100100",
  24191=>"001110100",
  24192=>"010111000",
  24193=>"110110100",
  24194=>"101110011",
  24195=>"110010001",
  24196=>"111001000",
  24197=>"001101010",
  24198=>"101010100",
  24199=>"000100100",
  24200=>"101011100",
  24201=>"101000100",
  24202=>"001101101",
  24203=>"000111010",
  24204=>"111100100",
  24205=>"011011111",
  24206=>"011011001",
  24207=>"001100001",
  24208=>"000101001",
  24209=>"110011000",
  24210=>"011111101",
  24211=>"111101000",
  24212=>"000010100",
  24213=>"100001100",
  24214=>"010011000",
  24215=>"000000100",
  24216=>"101111011",
  24217=>"100100001",
  24218=>"010011101",
  24219=>"010110001",
  24220=>"001100100",
  24221=>"100100101",
  24222=>"000001010",
  24223=>"011010100",
  24224=>"100100011",
  24225=>"011001000",
  24226=>"011001100",
  24227=>"011011101",
  24228=>"010111000",
  24229=>"000010010",
  24230=>"011010101",
  24231=>"001110000",
  24232=>"110000111",
  24233=>"000100010",
  24234=>"001110010",
  24235=>"011110010",
  24236=>"001010000",
  24237=>"101000100",
  24238=>"011001100",
  24239=>"110101111",
  24240=>"001000011",
  24241=>"011001001",
  24242=>"000100100",
  24243=>"011010011",
  24244=>"001101001",
  24245=>"010000000",
  24246=>"111000110",
  24247=>"011111101",
  24248=>"000010010",
  24249=>"111101101",
  24250=>"100001101",
  24251=>"011000000",
  24252=>"100010110",
  24253=>"100000000",
  24254=>"101000001",
  24255=>"011001111",
  24256=>"000111001",
  24257=>"010111000",
  24258=>"010110010",
  24259=>"011000001",
  24260=>"010010110",
  24261=>"000000110",
  24262=>"101011010",
  24263=>"000001011",
  24264=>"100011001",
  24265=>"111110101",
  24266=>"000010010",
  24267=>"110100111",
  24268=>"111001001",
  24269=>"001010100",
  24270=>"100001110",
  24271=>"111100100",
  24272=>"100001110",
  24273=>"010000010",
  24274=>"011100000",
  24275=>"100101000",
  24276=>"110001000",
  24277=>"110101110",
  24278=>"110001011",
  24279=>"101111111",
  24280=>"100000111",
  24281=>"011010111",
  24282=>"001010100",
  24283=>"000001000",
  24284=>"011111100",
  24285=>"000000000",
  24286=>"100011110",
  24287=>"111101101",
  24288=>"101001011",
  24289=>"111011100",
  24290=>"100111010",
  24291=>"011111110",
  24292=>"110110001",
  24293=>"010000010",
  24294=>"101001110",
  24295=>"111101111",
  24296=>"001110001",
  24297=>"011011011",
  24298=>"001010001",
  24299=>"000001101",
  24300=>"001001110",
  24301=>"110000001",
  24302=>"011100000",
  24303=>"010000001",
  24304=>"100000110",
  24305=>"111100110",
  24306=>"000110010",
  24307=>"010010001",
  24308=>"010111001",
  24309=>"111000101",
  24310=>"000110111",
  24311=>"101011000",
  24312=>"011011000",
  24313=>"010101001",
  24314=>"001001001",
  24315=>"100110011",
  24316=>"101001110",
  24317=>"100000100",
  24318=>"111001010",
  24319=>"110010011",
  24320=>"000000000",
  24321=>"101010101",
  24322=>"111101110",
  24323=>"110001111",
  24324=>"110101100",
  24325=>"010110110",
  24326=>"011011100",
  24327=>"001010110",
  24328=>"011111010",
  24329=>"001001010",
  24330=>"100110100",
  24331=>"111000111",
  24332=>"111101011",
  24333=>"100001000",
  24334=>"100010100",
  24335=>"000011111",
  24336=>"010011010",
  24337=>"111010010",
  24338=>"111101111",
  24339=>"100111110",
  24340=>"110100100",
  24341=>"010010000",
  24342=>"001100110",
  24343=>"111100000",
  24344=>"100001110",
  24345=>"011011001",
  24346=>"101110101",
  24347=>"010100110",
  24348=>"010111101",
  24349=>"110001111",
  24350=>"000011000",
  24351=>"001011010",
  24352=>"000111011",
  24353=>"011100100",
  24354=>"111101111",
  24355=>"111111010",
  24356=>"110101101",
  24357=>"000010111",
  24358=>"100010100",
  24359=>"101000101",
  24360=>"111001111",
  24361=>"000000010",
  24362=>"110010111",
  24363=>"001111101",
  24364=>"000001010",
  24365=>"001100100",
  24366=>"011000110",
  24367=>"110000101",
  24368=>"100000110",
  24369=>"010100000",
  24370=>"100000110",
  24371=>"010001001",
  24372=>"111111001",
  24373=>"100001101",
  24374=>"000111110",
  24375=>"101010000",
  24376=>"111101101",
  24377=>"010011100",
  24378=>"111100110",
  24379=>"110011001",
  24380=>"010011100",
  24381=>"010000001",
  24382=>"010010010",
  24383=>"101101101",
  24384=>"000101110",
  24385=>"000110001",
  24386=>"001001010",
  24387=>"111101111",
  24388=>"110101001",
  24389=>"111010101",
  24390=>"000100010",
  24391=>"110111010",
  24392=>"010101100",
  24393=>"000111011",
  24394=>"011011110",
  24395=>"100001000",
  24396=>"001101001",
  24397=>"100010010",
  24398=>"101010000",
  24399=>"011100011",
  24400=>"011100011",
  24401=>"111110101",
  24402=>"110110100",
  24403=>"000110100",
  24404=>"010100110",
  24405=>"100100000",
  24406=>"000001100",
  24407=>"000110010",
  24408=>"011011100",
  24409=>"011110101",
  24410=>"001001001",
  24411=>"001000001",
  24412=>"000110101",
  24413=>"010101111",
  24414=>"100101011",
  24415=>"100101110",
  24416=>"000100001",
  24417=>"110110101",
  24418=>"010111001",
  24419=>"111001110",
  24420=>"100010101",
  24421=>"110010100",
  24422=>"101001001",
  24423=>"001001010",
  24424=>"011010101",
  24425=>"100010100",
  24426=>"011001101",
  24427=>"010101101",
  24428=>"010010010",
  24429=>"000101110",
  24430=>"010000010",
  24431=>"011001000",
  24432=>"000010110",
  24433=>"110000010",
  24434=>"100100100",
  24435=>"101101100",
  24436=>"000111111",
  24437=>"101011000",
  24438=>"000110011",
  24439=>"110110001",
  24440=>"101101000",
  24441=>"011010001",
  24442=>"011100001",
  24443=>"100010001",
  24444=>"110100011",
  24445=>"011010111",
  24446=>"110001010",
  24447=>"111111111",
  24448=>"111001001",
  24449=>"110100011",
  24450=>"101000111",
  24451=>"001010110",
  24452=>"101000101",
  24453=>"011110000",
  24454=>"011000101",
  24455=>"001101011",
  24456=>"100110111",
  24457=>"101111010",
  24458=>"111110010",
  24459=>"111111100",
  24460=>"101111100",
  24461=>"110001101",
  24462=>"000110101",
  24463=>"001000111",
  24464=>"111101011",
  24465=>"001111000",
  24466=>"000000000",
  24467=>"000001111",
  24468=>"001100001",
  24469=>"010100101",
  24470=>"000111011",
  24471=>"011001010",
  24472=>"010101000",
  24473=>"111111111",
  24474=>"110010010",
  24475=>"110000000",
  24476=>"100100111",
  24477=>"100111100",
  24478=>"000000100",
  24479=>"110101011",
  24480=>"000111111",
  24481=>"000110000",
  24482=>"111001001",
  24483=>"000001000",
  24484=>"000011011",
  24485=>"100011010",
  24486=>"011111010",
  24487=>"111011110",
  24488=>"000010001",
  24489=>"000000101",
  24490=>"101100001",
  24491=>"111000001",
  24492=>"111010001",
  24493=>"000110111",
  24494=>"011010001",
  24495=>"010001001",
  24496=>"011010011",
  24497=>"110100110",
  24498=>"010100100",
  24499=>"101111000",
  24500=>"101001100",
  24501=>"100010000",
  24502=>"101100111",
  24503=>"010100100",
  24504=>"101010011",
  24505=>"000011011",
  24506=>"101111111",
  24507=>"000100100",
  24508=>"010001101",
  24509=>"010011010",
  24510=>"010100010",
  24511=>"000000000",
  24512=>"111001111",
  24513=>"000100100",
  24514=>"101010011",
  24515=>"110010010",
  24516=>"100000101",
  24517=>"000000011",
  24518=>"010010111",
  24519=>"110010100",
  24520=>"001000000",
  24521=>"111001101",
  24522=>"111011010",
  24523=>"100011011",
  24524=>"011110010",
  24525=>"001000100",
  24526=>"111000011",
  24527=>"110010011",
  24528=>"101111001",
  24529=>"000010011",
  24530=>"000111001",
  24531=>"000100001",
  24532=>"000000000",
  24533=>"010000100",
  24534=>"000001000",
  24535=>"001011100",
  24536=>"111001001",
  24537=>"111011110",
  24538=>"000011000",
  24539=>"111110000",
  24540=>"111000100",
  24541=>"100111010",
  24542=>"110100010",
  24543=>"000101010",
  24544=>"000100011",
  24545=>"111110000",
  24546=>"110111101",
  24547=>"111110010",
  24548=>"111101111",
  24549=>"011010001",
  24550=>"000011101",
  24551=>"010000011",
  24552=>"010100111",
  24553=>"111111010",
  24554=>"111110001",
  24555=>"000000011",
  24556=>"110000101",
  24557=>"101000110",
  24558=>"110001101",
  24559=>"111100111",
  24560=>"001111101",
  24561=>"101000101",
  24562=>"011010110",
  24563=>"011111111",
  24564=>"001011110",
  24565=>"011111000",
  24566=>"000101111",
  24567=>"011110110",
  24568=>"110110110",
  24569=>"000010011",
  24570=>"101010110",
  24571=>"100111111",
  24572=>"010010000",
  24573=>"110000101",
  24574=>"101001011",
  24575=>"010111101",
  24576=>"000011110",
  24577=>"000101010",
  24578=>"001101111",
  24579=>"111100010",
  24580=>"100111000",
  24581=>"011000000",
  24582=>"101001011",
  24583=>"101111000",
  24584=>"011110000",
  24585=>"101111100",
  24586=>"110000110",
  24587=>"101011101",
  24588=>"000001101",
  24589=>"110100110",
  24590=>"010010110",
  24591=>"110010101",
  24592=>"101111010",
  24593=>"011111100",
  24594=>"110101011",
  24595=>"101001011",
  24596=>"011010111",
  24597=>"110010010",
  24598=>"111110010",
  24599=>"101101001",
  24600=>"110111110",
  24601=>"001000110",
  24602=>"011010000",
  24603=>"111000101",
  24604=>"011000000",
  24605=>"111001101",
  24606=>"110001110",
  24607=>"000001111",
  24608=>"001001001",
  24609=>"100111100",
  24610=>"011110110",
  24611=>"110110101",
  24612=>"001101111",
  24613=>"001110100",
  24614=>"100000111",
  24615=>"001110010",
  24616=>"001101011",
  24617=>"100001111",
  24618=>"111111011",
  24619=>"010001011",
  24620=>"110111110",
  24621=>"001010101",
  24622=>"000110000",
  24623=>"101111111",
  24624=>"000111111",
  24625=>"101010101",
  24626=>"011101101",
  24627=>"011000100",
  24628=>"111000010",
  24629=>"010000010",
  24630=>"001011110",
  24631=>"010001010",
  24632=>"010100010",
  24633=>"001100111",
  24634=>"001000111",
  24635=>"100010111",
  24636=>"010000000",
  24637=>"110100010",
  24638=>"110010010",
  24639=>"001010111",
  24640=>"101010001",
  24641=>"011001101",
  24642=>"001011101",
  24643=>"010110010",
  24644=>"100100110",
  24645=>"101000000",
  24646=>"010100111",
  24647=>"100101101",
  24648=>"010110100",
  24649=>"001001011",
  24650=>"001011111",
  24651=>"011111000",
  24652=>"100001101",
  24653=>"111101101",
  24654=>"011010010",
  24655=>"010001001",
  24656=>"100011011",
  24657=>"110111101",
  24658=>"100100010",
  24659=>"001011001",
  24660=>"100111111",
  24661=>"001010100",
  24662=>"000101010",
  24663=>"000110000",
  24664=>"010000111",
  24665=>"110010101",
  24666=>"110111010",
  24667=>"110001000",
  24668=>"001000010",
  24669=>"101110011",
  24670=>"110100000",
  24671=>"000000011",
  24672=>"100100001",
  24673=>"100010110",
  24674=>"111010101",
  24675=>"001110101",
  24676=>"011001101",
  24677=>"110001111",
  24678=>"001000001",
  24679=>"011011111",
  24680=>"101100101",
  24681=>"101101010",
  24682=>"000011011",
  24683=>"110110100",
  24684=>"111011100",
  24685=>"111100001",
  24686=>"111101110",
  24687=>"100100000",
  24688=>"000001101",
  24689=>"000011101",
  24690=>"101101111",
  24691=>"101101011",
  24692=>"010011110",
  24693=>"011001000",
  24694=>"110000001",
  24695=>"011110111",
  24696=>"111100011",
  24697=>"110101110",
  24698=>"011110011",
  24699=>"011010010",
  24700=>"111111111",
  24701=>"000001101",
  24702=>"110011010",
  24703=>"100000001",
  24704=>"010011110",
  24705=>"000000011",
  24706=>"001100011",
  24707=>"001101100",
  24708=>"000010111",
  24709=>"001011110",
  24710=>"010111010",
  24711=>"000101100",
  24712=>"000110011",
  24713=>"000100101",
  24714=>"110011001",
  24715=>"101100001",
  24716=>"010011110",
  24717=>"111100111",
  24718=>"110100000",
  24719=>"001010100",
  24720=>"110101010",
  24721=>"011011110",
  24722=>"101010010",
  24723=>"110110100",
  24724=>"111100100",
  24725=>"011111000",
  24726=>"100001111",
  24727=>"010100010",
  24728=>"100111110",
  24729=>"011010100",
  24730=>"001101011",
  24731=>"011000100",
  24732=>"010110000",
  24733=>"010100000",
  24734=>"100101100",
  24735=>"101100010",
  24736=>"101101011",
  24737=>"011101101",
  24738=>"110110101",
  24739=>"010101011",
  24740=>"110101000",
  24741=>"010011010",
  24742=>"010100010",
  24743=>"100000111",
  24744=>"101110110",
  24745=>"001000001",
  24746=>"011111000",
  24747=>"000011100",
  24748=>"000110011",
  24749=>"110101001",
  24750=>"001010101",
  24751=>"011101110",
  24752=>"000110100",
  24753=>"101001011",
  24754=>"001111111",
  24755=>"101001101",
  24756=>"111110011",
  24757=>"001100000",
  24758=>"001100100",
  24759=>"111011000",
  24760=>"000000001",
  24761=>"001100000",
  24762=>"000110001",
  24763=>"101000011",
  24764=>"110000011",
  24765=>"011010110",
  24766=>"110011011",
  24767=>"100011111",
  24768=>"111001001",
  24769=>"010000111",
  24770=>"001110011",
  24771=>"111111011",
  24772=>"001000011",
  24773=>"010110010",
  24774=>"001011110",
  24775=>"100000111",
  24776=>"001100010",
  24777=>"010000000",
  24778=>"000001111",
  24779=>"111110010",
  24780=>"001110000",
  24781=>"011111100",
  24782=>"010001111",
  24783=>"010101101",
  24784=>"001111000",
  24785=>"010000101",
  24786=>"000110010",
  24787=>"011111100",
  24788=>"100010101",
  24789=>"000110001",
  24790=>"011100001",
  24791=>"011110001",
  24792=>"011000011",
  24793=>"000011001",
  24794=>"011011010",
  24795=>"000000000",
  24796=>"110100101",
  24797=>"110001101",
  24798=>"000011110",
  24799=>"100010011",
  24800=>"100001101",
  24801=>"100100101",
  24802=>"111110010",
  24803=>"100011001",
  24804=>"000110100",
  24805=>"010010110",
  24806=>"011000101",
  24807=>"110111110",
  24808=>"100010011",
  24809=>"010000010",
  24810=>"010001101",
  24811=>"000001001",
  24812=>"111011101",
  24813=>"100011010",
  24814=>"000101011",
  24815=>"000111000",
  24816=>"111100011",
  24817=>"001000110",
  24818=>"001100111",
  24819=>"101100100",
  24820=>"101101000",
  24821=>"101111100",
  24822=>"100010011",
  24823=>"001001010",
  24824=>"000001010",
  24825=>"011011011",
  24826=>"000000111",
  24827=>"100010011",
  24828=>"101100001",
  24829=>"000110111",
  24830=>"010011100",
  24831=>"101011101",
  24832=>"110100111",
  24833=>"001000111",
  24834=>"010000000",
  24835=>"111110101",
  24836=>"100111101",
  24837=>"111100010",
  24838=>"111111100",
  24839=>"101101011",
  24840=>"100000011",
  24841=>"000010111",
  24842=>"010110010",
  24843=>"100011001",
  24844=>"111011110",
  24845=>"000101000",
  24846=>"100110010",
  24847=>"100100111",
  24848=>"000001100",
  24849=>"000110011",
  24850=>"111011101",
  24851=>"010110101",
  24852=>"000001101",
  24853=>"011010000",
  24854=>"000000001",
  24855=>"110100011",
  24856=>"000110001",
  24857=>"100000101",
  24858=>"001100011",
  24859=>"000100101",
  24860=>"111011010",
  24861=>"110011110",
  24862=>"011101000",
  24863=>"100001000",
  24864=>"000001010",
  24865=>"000011010",
  24866=>"010000011",
  24867=>"011011100",
  24868=>"011110101",
  24869=>"101001001",
  24870=>"010010100",
  24871=>"110101101",
  24872=>"101100000",
  24873=>"101110110",
  24874=>"000001111",
  24875=>"101000010",
  24876=>"000101010",
  24877=>"110111001",
  24878=>"101001110",
  24879=>"001100001",
  24880=>"100101101",
  24881=>"111001111",
  24882=>"101101110",
  24883=>"011111010",
  24884=>"000111100",
  24885=>"001000000",
  24886=>"100000001",
  24887=>"101100110",
  24888=>"111101000",
  24889=>"110010000",
  24890=>"001101111",
  24891=>"011000110",
  24892=>"110100011",
  24893=>"101011111",
  24894=>"100001110",
  24895=>"010101100",
  24896=>"011001000",
  24897=>"011010001",
  24898=>"101101110",
  24899=>"010010010",
  24900=>"111010010",
  24901=>"001011001",
  24902=>"111100010",
  24903=>"010110110",
  24904=>"100011100",
  24905=>"000110000",
  24906=>"110110111",
  24907=>"101001100",
  24908=>"001001001",
  24909=>"010010110",
  24910=>"101101010",
  24911=>"011111011",
  24912=>"111011100",
  24913=>"110101111",
  24914=>"011100010",
  24915=>"111000110",
  24916=>"010011010",
  24917=>"101111101",
  24918=>"001000001",
  24919=>"101110101",
  24920=>"100100111",
  24921=>"110111011",
  24922=>"001000000",
  24923=>"010001000",
  24924=>"010001000",
  24925=>"110010011",
  24926=>"001111000",
  24927=>"000000001",
  24928=>"111000000",
  24929=>"011000010",
  24930=>"000000100",
  24931=>"100100100",
  24932=>"011000011",
  24933=>"011111000",
  24934=>"011010100",
  24935=>"101001101",
  24936=>"010010111",
  24937=>"100111101",
  24938=>"111000010",
  24939=>"100100110",
  24940=>"101110110",
  24941=>"100010010",
  24942=>"011100000",
  24943=>"010010010",
  24944=>"101011101",
  24945=>"100100111",
  24946=>"111111100",
  24947=>"110000100",
  24948=>"111101100",
  24949=>"011110100",
  24950=>"111010011",
  24951=>"110110000",
  24952=>"000000101",
  24953=>"000111111",
  24954=>"010110011",
  24955=>"010100101",
  24956=>"101100101",
  24957=>"111001110",
  24958=>"101000011",
  24959=>"111000101",
  24960=>"100110000",
  24961=>"110100011",
  24962=>"111100011",
  24963=>"101111101",
  24964=>"111100101",
  24965=>"111110101",
  24966=>"010111010",
  24967=>"100000010",
  24968=>"001000010",
  24969=>"110010101",
  24970=>"100000110",
  24971=>"010000010",
  24972=>"110011111",
  24973=>"101000000",
  24974=>"001111110",
  24975=>"001101100",
  24976=>"111111011",
  24977=>"100100101",
  24978=>"101101011",
  24979=>"111011100",
  24980=>"010000011",
  24981=>"110000100",
  24982=>"110010010",
  24983=>"110100100",
  24984=>"001011011",
  24985=>"110000100",
  24986=>"110111011",
  24987=>"001010011",
  24988=>"101010010",
  24989=>"100100110",
  24990=>"100001000",
  24991=>"110000111",
  24992=>"111110011",
  24993=>"101001011",
  24994=>"100111100",
  24995=>"100000010",
  24996=>"001110010",
  24997=>"111101100",
  24998=>"101001100",
  24999=>"110110100",
  25000=>"101100111",
  25001=>"010110010",
  25002=>"110110000",
  25003=>"011010011",
  25004=>"101110100",
  25005=>"011101000",
  25006=>"000110100",
  25007=>"101001100",
  25008=>"001000000",
  25009=>"111101010",
  25010=>"101101111",
  25011=>"000111001",
  25012=>"001100001",
  25013=>"101001010",
  25014=>"111110110",
  25015=>"110001110",
  25016=>"101101001",
  25017=>"111000100",
  25018=>"011000001",
  25019=>"101101001",
  25020=>"010110101",
  25021=>"000000100",
  25022=>"111000101",
  25023=>"100001000",
  25024=>"110110001",
  25025=>"000011011",
  25026=>"111010111",
  25027=>"101001011",
  25028=>"101001010",
  25029=>"100110101",
  25030=>"001111110",
  25031=>"010000100",
  25032=>"000000000",
  25033=>"101101111",
  25034=>"011010001",
  25035=>"010101100",
  25036=>"101111111",
  25037=>"111000100",
  25038=>"000111001",
  25039=>"101011001",
  25040=>"100110000",
  25041=>"010101110",
  25042=>"001001000",
  25043=>"110100011",
  25044=>"001011111",
  25045=>"111001111",
  25046=>"111000001",
  25047=>"001001010",
  25048=>"110001000",
  25049=>"111100111",
  25050=>"010100011",
  25051=>"011001000",
  25052=>"001100000",
  25053=>"111111110",
  25054=>"001100110",
  25055=>"000111011",
  25056=>"111111111",
  25057=>"110110011",
  25058=>"100110100",
  25059=>"001010110",
  25060=>"110000110",
  25061=>"100011100",
  25062=>"000001111",
  25063=>"001101101",
  25064=>"001000011",
  25065=>"100011111",
  25066=>"010011111",
  25067=>"010000010",
  25068=>"001100001",
  25069=>"110001001",
  25070=>"101100110",
  25071=>"010011010",
  25072=>"011001011",
  25073=>"000000010",
  25074=>"111011011",
  25075=>"001010011",
  25076=>"100011101",
  25077=>"010000011",
  25078=>"111001110",
  25079=>"010101011",
  25080=>"100111010",
  25081=>"101001110",
  25082=>"111010111",
  25083=>"000010101",
  25084=>"011101010",
  25085=>"011000011",
  25086=>"100011110",
  25087=>"101100000",
  25088=>"011000111",
  25089=>"010100101",
  25090=>"001011100",
  25091=>"100011101",
  25092=>"000100110",
  25093=>"011111111",
  25094=>"101101000",
  25095=>"001101111",
  25096=>"110110110",
  25097=>"000101101",
  25098=>"100110110",
  25099=>"010110000",
  25100=>"000110011",
  25101=>"100110111",
  25102=>"000000100",
  25103=>"101110101",
  25104=>"000101101",
  25105=>"000001111",
  25106=>"001011011",
  25107=>"011110011",
  25108=>"111001101",
  25109=>"100010100",
  25110=>"100111110",
  25111=>"110001111",
  25112=>"110100110",
  25113=>"010110111",
  25114=>"000010100",
  25115=>"100011001",
  25116=>"110100100",
  25117=>"011001101",
  25118=>"110000011",
  25119=>"100010010",
  25120=>"110110000",
  25121=>"011010011",
  25122=>"011001000",
  25123=>"010101001",
  25124=>"010111010",
  25125=>"000001110",
  25126=>"110011000",
  25127=>"110011011",
  25128=>"010101101",
  25129=>"110010010",
  25130=>"011010000",
  25131=>"111010000",
  25132=>"100100101",
  25133=>"001010110",
  25134=>"001100011",
  25135=>"010100011",
  25136=>"010001000",
  25137=>"000001111",
  25138=>"110110100",
  25139=>"010000010",
  25140=>"111011111",
  25141=>"000101011",
  25142=>"000110111",
  25143=>"000000010",
  25144=>"101101000",
  25145=>"001100000",
  25146=>"100000111",
  25147=>"000011111",
  25148=>"010111110",
  25149=>"110000010",
  25150=>"110011001",
  25151=>"000011111",
  25152=>"100100111",
  25153=>"011100000",
  25154=>"100000010",
  25155=>"111110100",
  25156=>"101000001",
  25157=>"100111010",
  25158=>"111110100",
  25159=>"111000111",
  25160=>"001001100",
  25161=>"111100110",
  25162=>"000101010",
  25163=>"101000110",
  25164=>"000001101",
  25165=>"111110000",
  25166=>"011100000",
  25167=>"101110000",
  25168=>"010100000",
  25169=>"111110100",
  25170=>"011100001",
  25171=>"101100000",
  25172=>"011100000",
  25173=>"110011011",
  25174=>"011000001",
  25175=>"011100111",
  25176=>"111100010",
  25177=>"111111110",
  25178=>"001110101",
  25179=>"011000001",
  25180=>"111100101",
  25181=>"001001010",
  25182=>"111011100",
  25183=>"001011110",
  25184=>"110101001",
  25185=>"011000101",
  25186=>"101000110",
  25187=>"111101001",
  25188=>"110101000",
  25189=>"101101101",
  25190=>"100110111",
  25191=>"111011000",
  25192=>"010110000",
  25193=>"010111010",
  25194=>"011100110",
  25195=>"000010101",
  25196=>"100011111",
  25197=>"000010001",
  25198=>"100100000",
  25199=>"000101001",
  25200=>"101100011",
  25201=>"110010000",
  25202=>"111100001",
  25203=>"000100111",
  25204=>"100010011",
  25205=>"000100101",
  25206=>"011000100",
  25207=>"111000011",
  25208=>"010001100",
  25209=>"000101110",
  25210=>"110110111",
  25211=>"100101010",
  25212=>"001011110",
  25213=>"001101000",
  25214=>"110010001",
  25215=>"011110111",
  25216=>"000011011",
  25217=>"111011111",
  25218=>"100101010",
  25219=>"110001111",
  25220=>"110110111",
  25221=>"000100001",
  25222=>"111000001",
  25223=>"111111100",
  25224=>"110110111",
  25225=>"011011110",
  25226=>"000000111",
  25227=>"100001001",
  25228=>"101000000",
  25229=>"110001101",
  25230=>"111111010",
  25231=>"110101111",
  25232=>"011110010",
  25233=>"110110110",
  25234=>"010011101",
  25235=>"011010111",
  25236=>"110010000",
  25237=>"111000011",
  25238=>"110011001",
  25239=>"010010011",
  25240=>"000100001",
  25241=>"000000010",
  25242=>"010100001",
  25243=>"011000011",
  25244=>"101000110",
  25245=>"100100000",
  25246=>"000010000",
  25247=>"110000011",
  25248=>"001011010",
  25249=>"111101011",
  25250=>"011000001",
  25251=>"110100000",
  25252=>"110101010",
  25253=>"001001110",
  25254=>"101010100",
  25255=>"110100010",
  25256=>"001001000",
  25257=>"001010111",
  25258=>"110100000",
  25259=>"100000100",
  25260=>"111010011",
  25261=>"011100010",
  25262=>"000010100",
  25263=>"000011011",
  25264=>"010000010",
  25265=>"101101111",
  25266=>"111010000",
  25267=>"010100110",
  25268=>"001010010",
  25269=>"000001110",
  25270=>"010000010",
  25271=>"011010001",
  25272=>"011111101",
  25273=>"110100000",
  25274=>"001011010",
  25275=>"001000010",
  25276=>"010000111",
  25277=>"100010001",
  25278=>"110001110",
  25279=>"000001100",
  25280=>"010110011",
  25281=>"010001110",
  25282=>"001101101",
  25283=>"110111100",
  25284=>"100111110",
  25285=>"111110111",
  25286=>"011011010",
  25287=>"000101110",
  25288=>"111111001",
  25289=>"010111101",
  25290=>"000110111",
  25291=>"111111010",
  25292=>"010101001",
  25293=>"011100010",
  25294=>"111000000",
  25295=>"111110001",
  25296=>"011110110",
  25297=>"010010001",
  25298=>"111100001",
  25299=>"000101001",
  25300=>"010110000",
  25301=>"000000010",
  25302=>"011110101",
  25303=>"001011010",
  25304=>"111110110",
  25305=>"000111110",
  25306=>"111011000",
  25307=>"110001101",
  25308=>"110001001",
  25309=>"110010000",
  25310=>"000111100",
  25311=>"010010111",
  25312=>"001100100",
  25313=>"000001101",
  25314=>"111101011",
  25315=>"001101011",
  25316=>"001101011",
  25317=>"000101110",
  25318=>"011101010",
  25319=>"011000101",
  25320=>"001000000",
  25321=>"010000000",
  25322=>"010011010",
  25323=>"000111010",
  25324=>"001101111",
  25325=>"111000010",
  25326=>"011011010",
  25327=>"010100110",
  25328=>"011101011",
  25329=>"110111111",
  25330=>"010110111",
  25331=>"000001000",
  25332=>"010011010",
  25333=>"101010110",
  25334=>"111010111",
  25335=>"101010010",
  25336=>"101010000",
  25337=>"011000011",
  25338=>"001001100",
  25339=>"101000001",
  25340=>"000011000",
  25341=>"001010110",
  25342=>"111011101",
  25343=>"000011001",
  25344=>"111100101",
  25345=>"001111010",
  25346=>"110111000",
  25347=>"100000010",
  25348=>"111111111",
  25349=>"010000000",
  25350=>"000100001",
  25351=>"001100010",
  25352=>"001111100",
  25353=>"010001010",
  25354=>"010101011",
  25355=>"001101110",
  25356=>"000010100",
  25357=>"001100101",
  25358=>"000011001",
  25359=>"101000110",
  25360=>"100011010",
  25361=>"100011100",
  25362=>"111100010",
  25363=>"101001011",
  25364=>"000000110",
  25365=>"010001111",
  25366=>"111001100",
  25367=>"111100110",
  25368=>"001010000",
  25369=>"010011000",
  25370=>"000100111",
  25371=>"110101011",
  25372=>"111011001",
  25373=>"001001001",
  25374=>"110100110",
  25375=>"001110010",
  25376=>"100111011",
  25377=>"101110101",
  25378=>"110011101",
  25379=>"110111001",
  25380=>"110100010",
  25381=>"100101101",
  25382=>"110000011",
  25383=>"010111001",
  25384=>"100101011",
  25385=>"100111101",
  25386=>"101111010",
  25387=>"110010111",
  25388=>"111111110",
  25389=>"001000111",
  25390=>"010010010",
  25391=>"101001101",
  25392=>"100010011",
  25393=>"010100101",
  25394=>"011110101",
  25395=>"001011010",
  25396=>"111100010",
  25397=>"001000010",
  25398=>"010111100",
  25399=>"010001100",
  25400=>"001010110",
  25401=>"010101101",
  25402=>"011001010",
  25403=>"010011010",
  25404=>"110010001",
  25405=>"101000010",
  25406=>"100011001",
  25407=>"011110110",
  25408=>"001111000",
  25409=>"110000000",
  25410=>"101011101",
  25411=>"000000100",
  25412=>"111100111",
  25413=>"000101100",
  25414=>"000100001",
  25415=>"001010110",
  25416=>"000110011",
  25417=>"001111110",
  25418=>"001001011",
  25419=>"111110110",
  25420=>"011100101",
  25421=>"111101000",
  25422=>"010100100",
  25423=>"101001100",
  25424=>"110100101",
  25425=>"001010101",
  25426=>"010010011",
  25427=>"000101011",
  25428=>"001000001",
  25429=>"110100110",
  25430=>"011001111",
  25431=>"011010001",
  25432=>"110110101",
  25433=>"100110111",
  25434=>"001010000",
  25435=>"000101110",
  25436=>"100001000",
  25437=>"111111000",
  25438=>"100110010",
  25439=>"001000011",
  25440=>"100101111",
  25441=>"001010111",
  25442=>"100001010",
  25443=>"011010110",
  25444=>"001110100",
  25445=>"010010000",
  25446=>"001000110",
  25447=>"111010011",
  25448=>"011001000",
  25449=>"100001110",
  25450=>"000001100",
  25451=>"111111000",
  25452=>"000100000",
  25453=>"000001000",
  25454=>"101110000",
  25455=>"011110100",
  25456=>"111111100",
  25457=>"010010010",
  25458=>"000111001",
  25459=>"001101011",
  25460=>"001110100",
  25461=>"010000010",
  25462=>"000111101",
  25463=>"110101110",
  25464=>"010011001",
  25465=>"110111011",
  25466=>"101111011",
  25467=>"100111111",
  25468=>"000000100",
  25469=>"111010101",
  25470=>"101101110",
  25471=>"110111010",
  25472=>"110001101",
  25473=>"001010101",
  25474=>"110011001",
  25475=>"010100100",
  25476=>"001011011",
  25477=>"111000000",
  25478=>"000101110",
  25479=>"000010010",
  25480=>"100011111",
  25481=>"000000011",
  25482=>"010011100",
  25483=>"000110101",
  25484=>"011011011",
  25485=>"100001100",
  25486=>"000000000",
  25487=>"111010111",
  25488=>"001110000",
  25489=>"110000001",
  25490=>"000000101",
  25491=>"111101100",
  25492=>"101011011",
  25493=>"000001110",
  25494=>"010010101",
  25495=>"011101000",
  25496=>"010100000",
  25497=>"001001101",
  25498=>"110101011",
  25499=>"100101000",
  25500=>"110110010",
  25501=>"001100010",
  25502=>"110001110",
  25503=>"011000001",
  25504=>"011011010",
  25505=>"110011000",
  25506=>"011000101",
  25507=>"111001001",
  25508=>"011000010",
  25509=>"011111011",
  25510=>"101001010",
  25511=>"001001110",
  25512=>"000101100",
  25513=>"011100111",
  25514=>"101111110",
  25515=>"111011010",
  25516=>"100101101",
  25517=>"001000001",
  25518=>"111111110",
  25519=>"010101100",
  25520=>"101010111",
  25521=>"011111111",
  25522=>"010101111",
  25523=>"001110001",
  25524=>"101001101",
  25525=>"111100010",
  25526=>"011100100",
  25527=>"110000011",
  25528=>"111111010",
  25529=>"000001110",
  25530=>"100000011",
  25531=>"110111101",
  25532=>"001001101",
  25533=>"100101111",
  25534=>"010110100",
  25535=>"110000101",
  25536=>"100011100",
  25537=>"001000011",
  25538=>"010100011",
  25539=>"010100111",
  25540=>"000111011",
  25541=>"001001100",
  25542=>"100100100",
  25543=>"010111010",
  25544=>"100100111",
  25545=>"100000001",
  25546=>"011101110",
  25547=>"000110111",
  25548=>"011001000",
  25549=>"111100100",
  25550=>"001111111",
  25551=>"100101010",
  25552=>"010011101",
  25553=>"010100010",
  25554=>"100001110",
  25555=>"110110101",
  25556=>"100001001",
  25557=>"011001010",
  25558=>"110111001",
  25559=>"100110111",
  25560=>"111110101",
  25561=>"101111110",
  25562=>"000001010",
  25563=>"110000001",
  25564=>"111000010",
  25565=>"101100010",
  25566=>"000110101",
  25567=>"100011101",
  25568=>"101000110",
  25569=>"001001100",
  25570=>"101101111",
  25571=>"001001000",
  25572=>"000110001",
  25573=>"111010100",
  25574=>"111010100",
  25575=>"111111100",
  25576=>"111000001",
  25577=>"000001001",
  25578=>"010110011",
  25579=>"000110111",
  25580=>"010011001",
  25581=>"101101110",
  25582=>"101100110",
  25583=>"011111010",
  25584=>"100011111",
  25585=>"101101110",
  25586=>"111001001",
  25587=>"101111001",
  25588=>"110100000",
  25589=>"000100110",
  25590=>"010101101",
  25591=>"011101110",
  25592=>"101110000",
  25593=>"011010011",
  25594=>"110001011",
  25595=>"101111110",
  25596=>"010000011",
  25597=>"111111111",
  25598=>"010010110",
  25599=>"100010110",
  25600=>"101111110",
  25601=>"101011011",
  25602=>"110101110",
  25603=>"111000101",
  25604=>"011101010",
  25605=>"010110101",
  25606=>"000101100",
  25607=>"010101110",
  25608=>"101111000",
  25609=>"001111000",
  25610=>"010000111",
  25611=>"110000101",
  25612=>"101101100",
  25613=>"101111111",
  25614=>"011111011",
  25615=>"111000010",
  25616=>"010101100",
  25617=>"011101110",
  25618=>"011001011",
  25619=>"011110011",
  25620=>"000100100",
  25621=>"010000011",
  25622=>"110001111",
  25623=>"110001001",
  25624=>"010010100",
  25625=>"110001101",
  25626=>"011110111",
  25627=>"111110100",
  25628=>"111011000",
  25629=>"110100001",
  25630=>"101010000",
  25631=>"110010011",
  25632=>"110011111",
  25633=>"101101110",
  25634=>"101101000",
  25635=>"011011001",
  25636=>"010010110",
  25637=>"000100100",
  25638=>"001101000",
  25639=>"011111111",
  25640=>"001000000",
  25641=>"110111101",
  25642=>"110101111",
  25643=>"001010011",
  25644=>"001110110",
  25645=>"000010010",
  25646=>"000001110",
  25647=>"100011000",
  25648=>"001000110",
  25649=>"011001100",
  25650=>"110111000",
  25651=>"101001010",
  25652=>"011011010",
  25653=>"000010011",
  25654=>"011011110",
  25655=>"011110101",
  25656=>"110101110",
  25657=>"010100111",
  25658=>"110101111",
  25659=>"110000101",
  25660=>"100001100",
  25661=>"110001101",
  25662=>"111011111",
  25663=>"100010101",
  25664=>"111000010",
  25665=>"111001100",
  25666=>"010000110",
  25667=>"110000001",
  25668=>"011100110",
  25669=>"011010111",
  25670=>"001000111",
  25671=>"010101101",
  25672=>"110011100",
  25673=>"010101000",
  25674=>"101001001",
  25675=>"111111011",
  25676=>"110001101",
  25677=>"110100101",
  25678=>"011111111",
  25679=>"111111101",
  25680=>"110101010",
  25681=>"111011000",
  25682=>"101001111",
  25683=>"111000001",
  25684=>"001111001",
  25685=>"101101110",
  25686=>"000011100",
  25687=>"010100010",
  25688=>"010111111",
  25689=>"001110110",
  25690=>"100100000",
  25691=>"101101100",
  25692=>"000100110",
  25693=>"111000010",
  25694=>"000111110",
  25695=>"010011111",
  25696=>"001000000",
  25697=>"111111000",
  25698=>"001010000",
  25699=>"000110101",
  25700=>"100011001",
  25701=>"101000101",
  25702=>"110110111",
  25703=>"100000100",
  25704=>"111011010",
  25705=>"011010000",
  25706=>"101000010",
  25707=>"101010011",
  25708=>"001000111",
  25709=>"110101101",
  25710=>"110010010",
  25711=>"110010001",
  25712=>"010010010",
  25713=>"100000000",
  25714=>"110010000",
  25715=>"000000010",
  25716=>"001110001",
  25717=>"010110111",
  25718=>"001010011",
  25719=>"110100110",
  25720=>"101101100",
  25721=>"100101000",
  25722=>"110100010",
  25723=>"100100010",
  25724=>"100000100",
  25725=>"011110110",
  25726=>"101100100",
  25727=>"100001111",
  25728=>"010111010",
  25729=>"100100110",
  25730=>"110011010",
  25731=>"110111100",
  25732=>"010001111",
  25733=>"000000101",
  25734=>"111100110",
  25735=>"000100110",
  25736=>"110011100",
  25737=>"111000010",
  25738=>"100010111",
  25739=>"101111100",
  25740=>"110000101",
  25741=>"010110100",
  25742=>"001001111",
  25743=>"011000010",
  25744=>"010001100",
  25745=>"000000111",
  25746=>"100110001",
  25747=>"101100011",
  25748=>"010111111",
  25749=>"000111000",
  25750=>"010100100",
  25751=>"100011001",
  25752=>"110111110",
  25753=>"111110010",
  25754=>"111100011",
  25755=>"001001011",
  25756=>"111000110",
  25757=>"000011001",
  25758=>"000001011",
  25759=>"011100010",
  25760=>"001101100",
  25761=>"001011101",
  25762=>"110011101",
  25763=>"110011010",
  25764=>"110111011",
  25765=>"111000101",
  25766=>"000000101",
  25767=>"000101011",
  25768=>"001100110",
  25769=>"100110011",
  25770=>"001010111",
  25771=>"000001111",
  25772=>"101001100",
  25773=>"100010110",
  25774=>"000100011",
  25775=>"101000111",
  25776=>"100011000",
  25777=>"100001010",
  25778=>"111110001",
  25779=>"110111111",
  25780=>"001101011",
  25781=>"101011001",
  25782=>"011011100",
  25783=>"010110111",
  25784=>"011011011",
  25785=>"010100000",
  25786=>"111111110",
  25787=>"000000111",
  25788=>"010010000",
  25789=>"000101101",
  25790=>"001001001",
  25791=>"111000100",
  25792=>"110100010",
  25793=>"010010010",
  25794=>"000101011",
  25795=>"100101001",
  25796=>"111111110",
  25797=>"000101101",
  25798=>"001000100",
  25799=>"101110111",
  25800=>"111010010",
  25801=>"001010101",
  25802=>"101011101",
  25803=>"010111100",
  25804=>"100111010",
  25805=>"001101000",
  25806=>"101101100",
  25807=>"001101000",
  25808=>"001000100",
  25809=>"101101110",
  25810=>"111101101",
  25811=>"000110110",
  25812=>"100011111",
  25813=>"101110001",
  25814=>"010101110",
  25815=>"000001110",
  25816=>"011110000",
  25817=>"110010110",
  25818=>"110111100",
  25819=>"000000001",
  25820=>"110111001",
  25821=>"110001100",
  25822=>"000110001",
  25823=>"110010001",
  25824=>"000111010",
  25825=>"111000111",
  25826=>"111110101",
  25827=>"010011011",
  25828=>"011010010",
  25829=>"011101100",
  25830=>"111000000",
  25831=>"101010110",
  25832=>"001010001",
  25833=>"111101001",
  25834=>"110101011",
  25835=>"101101111",
  25836=>"010011101",
  25837=>"111110100",
  25838=>"101000001",
  25839=>"001111000",
  25840=>"000100011",
  25841=>"011110110",
  25842=>"000100101",
  25843=>"000001100",
  25844=>"011111110",
  25845=>"011011010",
  25846=>"000111110",
  25847=>"111010000",
  25848=>"101111110",
  25849=>"100101000",
  25850=>"111000110",
  25851=>"111110100",
  25852=>"110100001",
  25853=>"100010010",
  25854=>"100000101",
  25855=>"010011000",
  25856=>"100111011",
  25857=>"010100100",
  25858=>"100100001",
  25859=>"011000001",
  25860=>"100011010",
  25861=>"010101000",
  25862=>"111110011",
  25863=>"010010110",
  25864=>"011000000",
  25865=>"111010101",
  25866=>"000000001",
  25867=>"111111110",
  25868=>"100110000",
  25869=>"010110001",
  25870=>"001001110",
  25871=>"110100010",
  25872=>"000100100",
  25873=>"000100110",
  25874=>"000110111",
  25875=>"110100001",
  25876=>"101101110",
  25877=>"111110011",
  25878=>"101011111",
  25879=>"000110100",
  25880=>"101110110",
  25881=>"000110110",
  25882=>"011111111",
  25883=>"100010110",
  25884=>"000010100",
  25885=>"011001010",
  25886=>"010101111",
  25887=>"000111101",
  25888=>"111110101",
  25889=>"000100110",
  25890=>"001010100",
  25891=>"100000101",
  25892=>"110000111",
  25893=>"111010001",
  25894=>"000110110",
  25895=>"110100010",
  25896=>"010101010",
  25897=>"011011000",
  25898=>"000101000",
  25899=>"101101000",
  25900=>"011111010",
  25901=>"011101110",
  25902=>"100100101",
  25903=>"111110010",
  25904=>"110011100",
  25905=>"110101100",
  25906=>"101101010",
  25907=>"111010010",
  25908=>"101010111",
  25909=>"110100111",
  25910=>"000100000",
  25911=>"011000010",
  25912=>"011000000",
  25913=>"000000011",
  25914=>"100101111",
  25915=>"000000001",
  25916=>"010000101",
  25917=>"010000001",
  25918=>"001000100",
  25919=>"111101010",
  25920=>"111000101",
  25921=>"000110100",
  25922=>"111111101",
  25923=>"011111101",
  25924=>"010101100",
  25925=>"010110001",
  25926=>"010011000",
  25927=>"001111111",
  25928=>"111110001",
  25929=>"011000000",
  25930=>"011110101",
  25931=>"011111110",
  25932=>"010101100",
  25933=>"010000101",
  25934=>"111001000",
  25935=>"111110010",
  25936=>"011011101",
  25937=>"101011101",
  25938=>"111111010",
  25939=>"110011011",
  25940=>"000000010",
  25941=>"101110010",
  25942=>"111010100",
  25943=>"110111111",
  25944=>"010001000",
  25945=>"100000001",
  25946=>"001000110",
  25947=>"001001110",
  25948=>"110011011",
  25949=>"000110101",
  25950=>"001010000",
  25951=>"100010111",
  25952=>"001001100",
  25953=>"101101110",
  25954=>"111011100",
  25955=>"100001011",
  25956=>"101010110",
  25957=>"001001001",
  25958=>"001100010",
  25959=>"001011001",
  25960=>"010111111",
  25961=>"111111001",
  25962=>"111100010",
  25963=>"001010100",
  25964=>"001110000",
  25965=>"011010100",
  25966=>"011000011",
  25967=>"000101101",
  25968=>"001011100",
  25969=>"010010010",
  25970=>"111001100",
  25971=>"011110111",
  25972=>"010011101",
  25973=>"011101001",
  25974=>"010000011",
  25975=>"001000010",
  25976=>"011010100",
  25977=>"011111111",
  25978=>"110101100",
  25979=>"110111101",
  25980=>"100001101",
  25981=>"011011011",
  25982=>"010011111",
  25983=>"111001000",
  25984=>"000000000",
  25985=>"000000000",
  25986=>"110101010",
  25987=>"001101110",
  25988=>"001101110",
  25989=>"010000110",
  25990=>"100001111",
  25991=>"110100110",
  25992=>"100000111",
  25993=>"110011111",
  25994=>"111000100",
  25995=>"001010110",
  25996=>"010101001",
  25997=>"110100000",
  25998=>"111111111",
  25999=>"011011010",
  26000=>"000111010",
  26001=>"010110000",
  26002=>"000101011",
  26003=>"101001101",
  26004=>"100011000",
  26005=>"111100000",
  26006=>"110100111",
  26007=>"011001111",
  26008=>"001110101",
  26009=>"100111110",
  26010=>"011100011",
  26011=>"010111101",
  26012=>"010010001",
  26013=>"011010101",
  26014=>"010000000",
  26015=>"011000001",
  26016=>"110111010",
  26017=>"111000001",
  26018=>"011101001",
  26019=>"100101111",
  26020=>"000100100",
  26021=>"110000000",
  26022=>"110001101",
  26023=>"011000100",
  26024=>"001011111",
  26025=>"011110101",
  26026=>"101010011",
  26027=>"011011000",
  26028=>"110000111",
  26029=>"000100011",
  26030=>"101010000",
  26031=>"000110100",
  26032=>"001100000",
  26033=>"000100010",
  26034=>"001000001",
  26035=>"100100000",
  26036=>"100001000",
  26037=>"011111100",
  26038=>"010010011",
  26039=>"001111010",
  26040=>"011101011",
  26041=>"111000000",
  26042=>"011001101",
  26043=>"111001110",
  26044=>"010001010",
  26045=>"101111010",
  26046=>"011101011",
  26047=>"100000001",
  26048=>"111111000",
  26049=>"011010110",
  26050=>"000100011",
  26051=>"001000001",
  26052=>"100001111",
  26053=>"111111110",
  26054=>"010111110",
  26055=>"110011000",
  26056=>"100001000",
  26057=>"101001000",
  26058=>"001000000",
  26059=>"011011000",
  26060=>"101111100",
  26061=>"111111000",
  26062=>"001001110",
  26063=>"100001101",
  26064=>"101101010",
  26065=>"100001110",
  26066=>"011100110",
  26067=>"001110110",
  26068=>"010110110",
  26069=>"010101110",
  26070=>"111010111",
  26071=>"111010101",
  26072=>"011101111",
  26073=>"011010010",
  26074=>"001110001",
  26075=>"001001110",
  26076=>"110011100",
  26077=>"001001000",
  26078=>"101110011",
  26079=>"001010001",
  26080=>"000100111",
  26081=>"001111101",
  26082=>"110101001",
  26083=>"001000001",
  26084=>"110001101",
  26085=>"110001011",
  26086=>"000111110",
  26087=>"101010010",
  26088=>"010100110",
  26089=>"000101100",
  26090=>"111110010",
  26091=>"100001100",
  26092=>"101010101",
  26093=>"101111001",
  26094=>"101111110",
  26095=>"110100010",
  26096=>"110001000",
  26097=>"110101001",
  26098=>"001010111",
  26099=>"001001110",
  26100=>"000001110",
  26101=>"001000110",
  26102=>"000110011",
  26103=>"101101001",
  26104=>"001100100",
  26105=>"101001000",
  26106=>"101100000",
  26107=>"001000010",
  26108=>"111100110",
  26109=>"110001100",
  26110=>"100001010",
  26111=>"000010001",
  26112=>"010110011",
  26113=>"111010011",
  26114=>"011000010",
  26115=>"111101010",
  26116=>"010011010",
  26117=>"000100010",
  26118=>"111011101",
  26119=>"000010100",
  26120=>"111110010",
  26121=>"110000000",
  26122=>"100010000",
  26123=>"001111011",
  26124=>"011000011",
  26125=>"010010000",
  26126=>"101011110",
  26127=>"001011011",
  26128=>"110001000",
  26129=>"111001100",
  26130=>"011010000",
  26131=>"111001011",
  26132=>"010111111",
  26133=>"001001001",
  26134=>"101011001",
  26135=>"100101011",
  26136=>"110101011",
  26137=>"000001001",
  26138=>"111000100",
  26139=>"000000110",
  26140=>"110111111",
  26141=>"110001011",
  26142=>"001110011",
  26143=>"000001010",
  26144=>"000001111",
  26145=>"101011100",
  26146=>"001111110",
  26147=>"000110111",
  26148=>"110100011",
  26149=>"100011101",
  26150=>"100110011",
  26151=>"010100100",
  26152=>"001101100",
  26153=>"110011000",
  26154=>"010110011",
  26155=>"111111110",
  26156=>"000000101",
  26157=>"000111011",
  26158=>"001110111",
  26159=>"011010100",
  26160=>"001100001",
  26161=>"011100011",
  26162=>"111100010",
  26163=>"011011000",
  26164=>"011110010",
  26165=>"100011011",
  26166=>"011100111",
  26167=>"010011010",
  26168=>"110100010",
  26169=>"100110010",
  26170=>"110100110",
  26171=>"110011000",
  26172=>"100010011",
  26173=>"101100000",
  26174=>"000000000",
  26175=>"000101111",
  26176=>"010001101",
  26177=>"111001111",
  26178=>"000011000",
  26179=>"010101111",
  26180=>"000101011",
  26181=>"001010011",
  26182=>"001010101",
  26183=>"010111010",
  26184=>"111100111",
  26185=>"110111011",
  26186=>"010111010",
  26187=>"010110010",
  26188=>"001000010",
  26189=>"110100101",
  26190=>"101010110",
  26191=>"010101111",
  26192=>"001101011",
  26193=>"011010010",
  26194=>"001111010",
  26195=>"101010011",
  26196=>"010100011",
  26197=>"111001101",
  26198=>"000111001",
  26199=>"100010000",
  26200=>"010011011",
  26201=>"110101000",
  26202=>"101011111",
  26203=>"100010000",
  26204=>"000101011",
  26205=>"110100000",
  26206=>"000010111",
  26207=>"101100100",
  26208=>"101010010",
  26209=>"010010001",
  26210=>"011110110",
  26211=>"111001111",
  26212=>"001011011",
  26213=>"111101000",
  26214=>"111110011",
  26215=>"010111100",
  26216=>"111001011",
  26217=>"101111111",
  26218=>"000110011",
  26219=>"111011101",
  26220=>"100010010",
  26221=>"101111111",
  26222=>"010011011",
  26223=>"001000011",
  26224=>"011110100",
  26225=>"101001011",
  26226=>"000001000",
  26227=>"001001101",
  26228=>"011000011",
  26229=>"010101001",
  26230=>"011011010",
  26231=>"000100100",
  26232=>"101001100",
  26233=>"011110101",
  26234=>"011110110",
  26235=>"010110101",
  26236=>"111100011",
  26237=>"010001000",
  26238=>"000101000",
  26239=>"010100010",
  26240=>"000011111",
  26241=>"100011100",
  26242=>"110010110",
  26243=>"101100001",
  26244=>"101111110",
  26245=>"101001010",
  26246=>"000110110",
  26247=>"111011011",
  26248=>"100001100",
  26249=>"001001001",
  26250=>"001111111",
  26251=>"111010010",
  26252=>"011100000",
  26253=>"001001110",
  26254=>"000111110",
  26255=>"100001010",
  26256=>"000110010",
  26257=>"000111010",
  26258=>"100000011",
  26259=>"011000111",
  26260=>"000101101",
  26261=>"011110010",
  26262=>"110011001",
  26263=>"010111001",
  26264=>"010101110",
  26265=>"101011001",
  26266=>"000001111",
  26267=>"011101110",
  26268=>"111110111",
  26269=>"000010011",
  26270=>"010010110",
  26271=>"010001000",
  26272=>"110000001",
  26273=>"100000111",
  26274=>"101011101",
  26275=>"011101001",
  26276=>"011110101",
  26277=>"110110110",
  26278=>"000010111",
  26279=>"000110110",
  26280=>"110110111",
  26281=>"011011011",
  26282=>"110101101",
  26283=>"011010100",
  26284=>"100001101",
  26285=>"110000000",
  26286=>"010101001",
  26287=>"100000110",
  26288=>"011101001",
  26289=>"010111100",
  26290=>"110011011",
  26291=>"111011110",
  26292=>"010001010",
  26293=>"000110001",
  26294=>"111100011",
  26295=>"001010011",
  26296=>"010011000",
  26297=>"101001111",
  26298=>"100101010",
  26299=>"010001011",
  26300=>"101011000",
  26301=>"110110001",
  26302=>"100100000",
  26303=>"101001110",
  26304=>"100100110",
  26305=>"101010000",
  26306=>"110101000",
  26307=>"001110010",
  26308=>"010110011",
  26309=>"001110111",
  26310=>"101111101",
  26311=>"110001011",
  26312=>"011110011",
  26313=>"011110111",
  26314=>"110001101",
  26315=>"000010000",
  26316=>"000000100",
  26317=>"000011001",
  26318=>"010111010",
  26319=>"011111000",
  26320=>"111101001",
  26321=>"110110111",
  26322=>"011100010",
  26323=>"100011011",
  26324=>"010100100",
  26325=>"000101000",
  26326=>"000100110",
  26327=>"111010101",
  26328=>"000000000",
  26329=>"000011101",
  26330=>"100011100",
  26331=>"001110110",
  26332=>"101000101",
  26333=>"111111111",
  26334=>"000010101",
  26335=>"000101110",
  26336=>"000000111",
  26337=>"111100111",
  26338=>"100111011",
  26339=>"100011110",
  26340=>"111111111",
  26341=>"110111000",
  26342=>"101001101",
  26343=>"110110110",
  26344=>"001011010",
  26345=>"011000010",
  26346=>"011100010",
  26347=>"111001101",
  26348=>"111001010",
  26349=>"001000011",
  26350=>"100100110",
  26351=>"001001011",
  26352=>"101111111",
  26353=>"101011000",
  26354=>"101110110",
  26355=>"010111000",
  26356=>"110000101",
  26357=>"111001100",
  26358=>"100000001",
  26359=>"011000010",
  26360=>"101100001",
  26361=>"100100101",
  26362=>"111000001",
  26363=>"111110000",
  26364=>"001100110",
  26365=>"011110000",
  26366=>"111100000",
  26367=>"010011101",
  26368=>"111010100",
  26369=>"010011000",
  26370=>"100110001",
  26371=>"010011101",
  26372=>"011011000",
  26373=>"111110111",
  26374=>"001101011",
  26375=>"001111111",
  26376=>"001110100",
  26377=>"100010010",
  26378=>"010010100",
  26379=>"101010000",
  26380=>"101111111",
  26381=>"100011011",
  26382=>"010010010",
  26383=>"101111011",
  26384=>"111011110",
  26385=>"000000011",
  26386=>"111101011",
  26387=>"010111100",
  26388=>"110011000",
  26389=>"001101011",
  26390=>"001101000",
  26391=>"011010010",
  26392=>"010110010",
  26393=>"100101001",
  26394=>"011111010",
  26395=>"000011000",
  26396=>"100001100",
  26397=>"110110101",
  26398=>"001100111",
  26399=>"001110000",
  26400=>"110111001",
  26401=>"001111111",
  26402=>"000010000",
  26403=>"010000101",
  26404=>"100001001",
  26405=>"010111010",
  26406=>"110100000",
  26407=>"011101010",
  26408=>"011100111",
  26409=>"101111011",
  26410=>"010011111",
  26411=>"101101011",
  26412=>"110001010",
  26413=>"000011001",
  26414=>"110100001",
  26415=>"000101010",
  26416=>"110001000",
  26417=>"100000101",
  26418=>"010111000",
  26419=>"111011011",
  26420=>"110111110",
  26421=>"111111010",
  26422=>"010010010",
  26423=>"010011010",
  26424=>"010010010",
  26425=>"111010000",
  26426=>"000110011",
  26427=>"100001011",
  26428=>"010000001",
  26429=>"111000001",
  26430=>"001100100",
  26431=>"101010101",
  26432=>"100100101",
  26433=>"100100110",
  26434=>"111100101",
  26435=>"110000111",
  26436=>"011111110",
  26437=>"001101111",
  26438=>"110000100",
  26439=>"101100001",
  26440=>"101001001",
  26441=>"000010001",
  26442=>"110110000",
  26443=>"000000001",
  26444=>"001110100",
  26445=>"001110101",
  26446=>"011111110",
  26447=>"110111111",
  26448=>"101000101",
  26449=>"100101001",
  26450=>"001100011",
  26451=>"100101110",
  26452=>"001001010",
  26453=>"001011110",
  26454=>"011000010",
  26455=>"001000000",
  26456=>"010001101",
  26457=>"110111110",
  26458=>"001011000",
  26459=>"001101100",
  26460=>"101111000",
  26461=>"000000001",
  26462=>"010100111",
  26463=>"010101101",
  26464=>"010100010",
  26465=>"000110101",
  26466=>"001110101",
  26467=>"010001000",
  26468=>"000000011",
  26469=>"000001100",
  26470=>"011111001",
  26471=>"111110000",
  26472=>"100111101",
  26473=>"001101001",
  26474=>"100101101",
  26475=>"111000001",
  26476=>"000010011",
  26477=>"100100011",
  26478=>"001101111",
  26479=>"110100100",
  26480=>"100000001",
  26481=>"100100100",
  26482=>"011101110",
  26483=>"000101101",
  26484=>"010110000",
  26485=>"111101010",
  26486=>"010000010",
  26487=>"011000010",
  26488=>"001111111",
  26489=>"101000001",
  26490=>"011110010",
  26491=>"000111010",
  26492=>"100110010",
  26493=>"001100100",
  26494=>"000101011",
  26495=>"100100110",
  26496=>"000000001",
  26497=>"110011111",
  26498=>"011001001",
  26499=>"111101011",
  26500=>"000000100",
  26501=>"000100001",
  26502=>"001001100",
  26503=>"101001111",
  26504=>"111111111",
  26505=>"101000010",
  26506=>"001000001",
  26507=>"111110011",
  26508=>"100011011",
  26509=>"100001000",
  26510=>"000100010",
  26511=>"001010100",
  26512=>"101000000",
  26513=>"001111111",
  26514=>"011001001",
  26515=>"001000000",
  26516=>"101110010",
  26517=>"100100110",
  26518=>"100011111",
  26519=>"010111011",
  26520=>"110100011",
  26521=>"001011101",
  26522=>"100000111",
  26523=>"101010100",
  26524=>"100110001",
  26525=>"101011000",
  26526=>"101000011",
  26527=>"000000010",
  26528=>"100011111",
  26529=>"001010010",
  26530=>"111100100",
  26531=>"100000100",
  26532=>"000100101",
  26533=>"111001001",
  26534=>"010111111",
  26535=>"010110011",
  26536=>"101101111",
  26537=>"001011100",
  26538=>"000011010",
  26539=>"001000011",
  26540=>"100100000",
  26541=>"001001000",
  26542=>"110011001",
  26543=>"001010000",
  26544=>"011001100",
  26545=>"111010000",
  26546=>"000110110",
  26547=>"000110001",
  26548=>"001010110",
  26549=>"000001000",
  26550=>"111111001",
  26551=>"100111001",
  26552=>"101111010",
  26553=>"011110011",
  26554=>"010111001",
  26555=>"010100011",
  26556=>"000100011",
  26557=>"100100110",
  26558=>"101100110",
  26559=>"000100011",
  26560=>"011001110",
  26561=>"111001000",
  26562=>"011000110",
  26563=>"000010101",
  26564=>"110110100",
  26565=>"101100111",
  26566=>"100011100",
  26567=>"110010011",
  26568=>"111100101",
  26569=>"000110000",
  26570=>"111111010",
  26571=>"010001000",
  26572=>"010100110",
  26573=>"011110010",
  26574=>"000110101",
  26575=>"110110010",
  26576=>"101111100",
  26577=>"000010110",
  26578=>"000100010",
  26579=>"001011011",
  26580=>"101011111",
  26581=>"000001101",
  26582=>"010011010",
  26583=>"111010110",
  26584=>"010010000",
  26585=>"101001111",
  26586=>"011111001",
  26587=>"010110010",
  26588=>"111011100",
  26589=>"001011000",
  26590=>"100000011",
  26591=>"101111000",
  26592=>"110100100",
  26593=>"000001111",
  26594=>"101111011",
  26595=>"011011111",
  26596=>"111011000",
  26597=>"011011111",
  26598=>"100101111",
  26599=>"101100111",
  26600=>"111111010",
  26601=>"011111110",
  26602=>"101011100",
  26603=>"011101100",
  26604=>"010010011",
  26605=>"000011101",
  26606=>"100000011",
  26607=>"011011101",
  26608=>"110010100",
  26609=>"010010011",
  26610=>"111110101",
  26611=>"000111101",
  26612=>"011011110",
  26613=>"001101011",
  26614=>"100110101",
  26615=>"101101010",
  26616=>"000110010",
  26617=>"000110101",
  26618=>"000110111",
  26619=>"101110110",
  26620=>"100111111",
  26621=>"000000100",
  26622=>"101111011",
  26623=>"100100011",
  26624=>"010010100",
  26625=>"010010010",
  26626=>"010011101",
  26627=>"111110000",
  26628=>"101010010",
  26629=>"101011010",
  26630=>"001110110",
  26631=>"101001101",
  26632=>"010001111",
  26633=>"010110000",
  26634=>"100000100",
  26635=>"111010111",
  26636=>"110011010",
  26637=>"110111111",
  26638=>"011100010",
  26639=>"011010010",
  26640=>"001111001",
  26641=>"101010000",
  26642=>"100110110",
  26643=>"110000010",
  26644=>"011110001",
  26645=>"101011011",
  26646=>"101010001",
  26647=>"100110001",
  26648=>"110010110",
  26649=>"101111101",
  26650=>"011100001",
  26651=>"110101101",
  26652=>"100011111",
  26653=>"101100010",
  26654=>"110001000",
  26655=>"010110010",
  26656=>"001000100",
  26657=>"100010000",
  26658=>"001001100",
  26659=>"100001000",
  26660=>"000001101",
  26661=>"101011010",
  26662=>"111001001",
  26663=>"000010000",
  26664=>"001100111",
  26665=>"010111010",
  26666=>"101101110",
  26667=>"000001011",
  26668=>"010011110",
  26669=>"110111101",
  26670=>"111100010",
  26671=>"010001101",
  26672=>"100010001",
  26673=>"111001101",
  26674=>"011001111",
  26675=>"000100001",
  26676=>"000101010",
  26677=>"100110010",
  26678=>"101000100",
  26679=>"100101111",
  26680=>"100101111",
  26681=>"100010011",
  26682=>"111101000",
  26683=>"010000101",
  26684=>"100100000",
  26685=>"010001111",
  26686=>"101101000",
  26687=>"000111011",
  26688=>"111110111",
  26689=>"001011001",
  26690=>"100011000",
  26691=>"011011011",
  26692=>"000011010",
  26693=>"001000111",
  26694=>"010011001",
  26695=>"000011010",
  26696=>"001101111",
  26697=>"110101011",
  26698=>"111001101",
  26699=>"000100001",
  26700=>"100000100",
  26701=>"011101100",
  26702=>"001110101",
  26703=>"111100111",
  26704=>"110110010",
  26705=>"001111110",
  26706=>"111011001",
  26707=>"100011001",
  26708=>"111101110",
  26709=>"101101010",
  26710=>"011101111",
  26711=>"110100000",
  26712=>"111001000",
  26713=>"000001010",
  26714=>"011101101",
  26715=>"000100111",
  26716=>"101101110",
  26717=>"110001010",
  26718=>"111110101",
  26719=>"110000001",
  26720=>"000000100",
  26721=>"001110010",
  26722=>"000100011",
  26723=>"100110100",
  26724=>"111110100",
  26725=>"001011010",
  26726=>"101100110",
  26727=>"000100111",
  26728=>"110111101",
  26729=>"101100010",
  26730=>"110010100",
  26731=>"010110001",
  26732=>"001110111",
  26733=>"110001011",
  26734=>"110010111",
  26735=>"010011011",
  26736=>"110001101",
  26737=>"110000101",
  26738=>"111100011",
  26739=>"001110000",
  26740=>"111111111",
  26741=>"011001101",
  26742=>"111111111",
  26743=>"111001000",
  26744=>"100111000",
  26745=>"010110001",
  26746=>"010010101",
  26747=>"011110000",
  26748=>"111010111",
  26749=>"100100010",
  26750=>"100011000",
  26751=>"101000000",
  26752=>"001101001",
  26753=>"001100111",
  26754=>"101010001",
  26755=>"110110110",
  26756=>"101010010",
  26757=>"001101111",
  26758=>"110100110",
  26759=>"101110000",
  26760=>"001011000",
  26761=>"001100010",
  26762=>"000001011",
  26763=>"111111110",
  26764=>"100111001",
  26765=>"110111011",
  26766=>"101100110",
  26767=>"110100001",
  26768=>"000110011",
  26769=>"001001110",
  26770=>"101000111",
  26771=>"101100100",
  26772=>"111101100",
  26773=>"011111101",
  26774=>"001010101",
  26775=>"000001010",
  26776=>"000011111",
  26777=>"100100000",
  26778=>"101011011",
  26779=>"001010010",
  26780=>"011111000",
  26781=>"011101010",
  26782=>"100110010",
  26783=>"111001001",
  26784=>"001000101",
  26785=>"101100010",
  26786=>"100100111",
  26787=>"000101110",
  26788=>"101001011",
  26789=>"000101101",
  26790=>"010010001",
  26791=>"100000100",
  26792=>"110110011",
  26793=>"101000111",
  26794=>"111111101",
  26795=>"100011011",
  26796=>"100001011",
  26797=>"111101001",
  26798=>"011000011",
  26799=>"110011100",
  26800=>"110100111",
  26801=>"111010010",
  26802=>"011011110",
  26803=>"100100000",
  26804=>"110001010",
  26805=>"101111010",
  26806=>"110000001",
  26807=>"001111110",
  26808=>"101100100",
  26809=>"010000100",
  26810=>"001110000",
  26811=>"000010011",
  26812=>"000111001",
  26813=>"011110111",
  26814=>"001101111",
  26815=>"110110000",
  26816=>"000010010",
  26817=>"111010100",
  26818=>"110011111",
  26819=>"011010100",
  26820=>"111000001",
  26821=>"000001111",
  26822=>"000110111",
  26823=>"111011111",
  26824=>"011010000",
  26825=>"001100011",
  26826=>"011111110",
  26827=>"001011011",
  26828=>"110110111",
  26829=>"110110111",
  26830=>"100111100",
  26831=>"001001001",
  26832=>"010010001",
  26833=>"100001010",
  26834=>"011001000",
  26835=>"101010110",
  26836=>"001100010",
  26837=>"000101011",
  26838=>"110011101",
  26839=>"001100100",
  26840=>"000110100",
  26841=>"001000101",
  26842=>"001101011",
  26843=>"011110111",
  26844=>"001111101",
  26845=>"011111111",
  26846=>"000010001",
  26847=>"110001001",
  26848=>"111100010",
  26849=>"101110001",
  26850=>"101000111",
  26851=>"111011111",
  26852=>"010011100",
  26853=>"000111101",
  26854=>"110000001",
  26855=>"100000001",
  26856=>"100001101",
  26857=>"011010101",
  26858=>"000100011",
  26859=>"011010000",
  26860=>"111000100",
  26861=>"000101100",
  26862=>"000000110",
  26863=>"110111011",
  26864=>"110010001",
  26865=>"001000110",
  26866=>"000001101",
  26867=>"001010010",
  26868=>"100100111",
  26869=>"110010001",
  26870=>"011100000",
  26871=>"111110111",
  26872=>"100001011",
  26873=>"001000000",
  26874=>"011010010",
  26875=>"111001010",
  26876=>"101010111",
  26877=>"010010111",
  26878=>"101110111",
  26879=>"101011010",
  26880=>"010001001",
  26881=>"001001110",
  26882=>"010011111",
  26883=>"111100101",
  26884=>"101001010",
  26885=>"110011000",
  26886=>"010000100",
  26887=>"101010100",
  26888=>"100101111",
  26889=>"101011100",
  26890=>"111000110",
  26891=>"100111010",
  26892=>"010101111",
  26893=>"000111000",
  26894=>"101100100",
  26895=>"101000001",
  26896=>"101011111",
  26897=>"111101110",
  26898=>"010111110",
  26899=>"001111001",
  26900=>"110000100",
  26901=>"100111001",
  26902=>"101001101",
  26903=>"111001110",
  26904=>"001101110",
  26905=>"101100001",
  26906=>"100111111",
  26907=>"011101010",
  26908=>"010110000",
  26909=>"110000000",
  26910=>"110101011",
  26911=>"000010000",
  26912=>"110101000",
  26913=>"111100001",
  26914=>"101011110",
  26915=>"000010101",
  26916=>"110001100",
  26917=>"000101110",
  26918=>"000111000",
  26919=>"111010111",
  26920=>"000010110",
  26921=>"101010010",
  26922=>"100010100",
  26923=>"011001011",
  26924=>"110001001",
  26925=>"000000000",
  26926=>"111111001",
  26927=>"101010110",
  26928=>"101000000",
  26929=>"101000010",
  26930=>"000000101",
  26931=>"001110100",
  26932=>"010000111",
  26933=>"001011110",
  26934=>"010111001",
  26935=>"000001000",
  26936=>"110110110",
  26937=>"001000100",
  26938=>"010011011",
  26939=>"000111101",
  26940=>"000000000",
  26941=>"101110000",
  26942=>"011000011",
  26943=>"010111101",
  26944=>"000011000",
  26945=>"111000001",
  26946=>"011010001",
  26947=>"011101011",
  26948=>"110100110",
  26949=>"000111011",
  26950=>"001001010",
  26951=>"001011010",
  26952=>"000100000",
  26953=>"111010000",
  26954=>"010010011",
  26955=>"000001001",
  26956=>"100100111",
  26957=>"011101000",
  26958=>"000000011",
  26959=>"111110000",
  26960=>"011001001",
  26961=>"111010010",
  26962=>"101101100",
  26963=>"100110001",
  26964=>"010111110",
  26965=>"101000110",
  26966=>"110000100",
  26967=>"111110000",
  26968=>"111000011",
  26969=>"010011110",
  26970=>"000001010",
  26971=>"001101100",
  26972=>"000101110",
  26973=>"000011011",
  26974=>"100011011",
  26975=>"101000011",
  26976=>"110111111",
  26977=>"000001100",
  26978=>"001100101",
  26979=>"100110111",
  26980=>"101111010",
  26981=>"100101001",
  26982=>"010111000",
  26983=>"110111100",
  26984=>"110100001",
  26985=>"011001011",
  26986=>"010110101",
  26987=>"010010110",
  26988=>"111100101",
  26989=>"101101001",
  26990=>"000011101",
  26991=>"110010110",
  26992=>"000110010",
  26993=>"110001100",
  26994=>"000110111",
  26995=>"101101001",
  26996=>"000101110",
  26997=>"001100000",
  26998=>"001010011",
  26999=>"011100010",
  27000=>"000011100",
  27001=>"100000110",
  27002=>"101111101",
  27003=>"010100110",
  27004=>"011010111",
  27005=>"110011010",
  27006=>"111010111",
  27007=>"111011110",
  27008=>"100001001",
  27009=>"101100000",
  27010=>"111110111",
  27011=>"000101111",
  27012=>"100011101",
  27013=>"100011100",
  27014=>"011110011",
  27015=>"100110101",
  27016=>"011010001",
  27017=>"110010011",
  27018=>"010011001",
  27019=>"001011011",
  27020=>"010010010",
  27021=>"011101011",
  27022=>"011111101",
  27023=>"100011111",
  27024=>"100111100",
  27025=>"100001001",
  27026=>"111000001",
  27027=>"011111111",
  27028=>"101111011",
  27029=>"011111100",
  27030=>"010110001",
  27031=>"000110010",
  27032=>"010000010",
  27033=>"110110010",
  27034=>"111011111",
  27035=>"101111111",
  27036=>"110110010",
  27037=>"101110010",
  27038=>"101010101",
  27039=>"111000100",
  27040=>"110100010",
  27041=>"101100111",
  27042=>"111101100",
  27043=>"000000000",
  27044=>"011010001",
  27045=>"111011011",
  27046=>"011000010",
  27047=>"010011001",
  27048=>"000011110",
  27049=>"010000100",
  27050=>"000000101",
  27051=>"111000101",
  27052=>"000000111",
  27053=>"100010011",
  27054=>"100011000",
  27055=>"000010101",
  27056=>"011111001",
  27057=>"010100010",
  27058=>"000011111",
  27059=>"011000111",
  27060=>"100010111",
  27061=>"011101101",
  27062=>"111100001",
  27063=>"110100110",
  27064=>"001101111",
  27065=>"110000010",
  27066=>"001110101",
  27067=>"010111111",
  27068=>"001011010",
  27069=>"111000100",
  27070=>"001100001",
  27071=>"110110010",
  27072=>"010000001",
  27073=>"001001010",
  27074=>"110011101",
  27075=>"010011101",
  27076=>"000000010",
  27077=>"101110110",
  27078=>"100000000",
  27079=>"010000011",
  27080=>"101000011",
  27081=>"111110011",
  27082=>"111101001",
  27083=>"000011001",
  27084=>"011011000",
  27085=>"011000111",
  27086=>"110010111",
  27087=>"000011010",
  27088=>"101001111",
  27089=>"001111100",
  27090=>"110100101",
  27091=>"101101000",
  27092=>"101101010",
  27093=>"101101101",
  27094=>"010000000",
  27095=>"001001000",
  27096=>"000101101",
  27097=>"000011010",
  27098=>"110010011",
  27099=>"101000000",
  27100=>"110101110",
  27101=>"011101011",
  27102=>"111010110",
  27103=>"110000101",
  27104=>"010101100",
  27105=>"111100001",
  27106=>"101100001",
  27107=>"111111111",
  27108=>"010100000",
  27109=>"111001111",
  27110=>"100000010",
  27111=>"101111011",
  27112=>"001000011",
  27113=>"011111000",
  27114=>"001101010",
  27115=>"000000010",
  27116=>"111000111",
  27117=>"111000110",
  27118=>"100000101",
  27119=>"000010000",
  27120=>"100010000",
  27121=>"111111010",
  27122=>"111011010",
  27123=>"101101011",
  27124=>"000011011",
  27125=>"000011101",
  27126=>"011101100",
  27127=>"100111100",
  27128=>"000000111",
  27129=>"101000101",
  27130=>"100001010",
  27131=>"010101011",
  27132=>"101011110",
  27133=>"000101001",
  27134=>"001010011",
  27135=>"111100100",
  27136=>"001001101",
  27137=>"110101001",
  27138=>"110100001",
  27139=>"000101111",
  27140=>"010011000",
  27141=>"110110101",
  27142=>"011011010",
  27143=>"110111111",
  27144=>"001010101",
  27145=>"011010100",
  27146=>"100101101",
  27147=>"100000000",
  27148=>"001001001",
  27149=>"000011010",
  27150=>"100011110",
  27151=>"010100010",
  27152=>"111011101",
  27153=>"110101110",
  27154=>"011001001",
  27155=>"101101111",
  27156=>"111001010",
  27157=>"010011000",
  27158=>"110101101",
  27159=>"111000110",
  27160=>"100001011",
  27161=>"011000110",
  27162=>"010000110",
  27163=>"010010111",
  27164=>"100001110",
  27165=>"001000100",
  27166=>"101001010",
  27167=>"110010000",
  27168=>"000000000",
  27169=>"101100100",
  27170=>"011000110",
  27171=>"011110101",
  27172=>"111011001",
  27173=>"000011000",
  27174=>"101000111",
  27175=>"000111000",
  27176=>"101101100",
  27177=>"011101010",
  27178=>"001011100",
  27179=>"000001110",
  27180=>"100001110",
  27181=>"000001000",
  27182=>"110011100",
  27183=>"000111111",
  27184=>"011010100",
  27185=>"101100010",
  27186=>"010101110",
  27187=>"000011100",
  27188=>"010111010",
  27189=>"101001101",
  27190=>"111000010",
  27191=>"110110011",
  27192=>"111111110",
  27193=>"010000100",
  27194=>"010001001",
  27195=>"010010101",
  27196=>"111100111",
  27197=>"000111111",
  27198=>"000001110",
  27199=>"000110100",
  27200=>"101000010",
  27201=>"011000011",
  27202=>"010010010",
  27203=>"100000001",
  27204=>"110111110",
  27205=>"010011001",
  27206=>"011000011",
  27207=>"011101010",
  27208=>"001011001",
  27209=>"010000101",
  27210=>"001110011",
  27211=>"100100010",
  27212=>"000111010",
  27213=>"000000000",
  27214=>"010010111",
  27215=>"000011000",
  27216=>"000011100",
  27217=>"011101111",
  27218=>"011001000",
  27219=>"011010001",
  27220=>"010001011",
  27221=>"010101100",
  27222=>"011111111",
  27223=>"010101010",
  27224=>"100101000",
  27225=>"111000010",
  27226=>"010110110",
  27227=>"110110111",
  27228=>"111100000",
  27229=>"110000101",
  27230=>"000000100",
  27231=>"111010011",
  27232=>"100011100",
  27233=>"001110010",
  27234=>"110100111",
  27235=>"101101110",
  27236=>"111110011",
  27237=>"111110101",
  27238=>"001101111",
  27239=>"000100011",
  27240=>"100110001",
  27241=>"101000101",
  27242=>"110100010",
  27243=>"000001000",
  27244=>"000001101",
  27245=>"010000000",
  27246=>"100011110",
  27247=>"000101011",
  27248=>"110111001",
  27249=>"001000110",
  27250=>"111101110",
  27251=>"011111010",
  27252=>"110001010",
  27253=>"000011001",
  27254=>"100001000",
  27255=>"101100000",
  27256=>"110111111",
  27257=>"110010110",
  27258=>"101110110",
  27259=>"101100011",
  27260=>"100001010",
  27261=>"100000110",
  27262=>"000010110",
  27263=>"010101110",
  27264=>"101110000",
  27265=>"100101100",
  27266=>"101000111",
  27267=>"000101110",
  27268=>"001111111",
  27269=>"000100010",
  27270=>"000110101",
  27271=>"111101011",
  27272=>"011000111",
  27273=>"110110111",
  27274=>"000010011",
  27275=>"001111011",
  27276=>"110001101",
  27277=>"100111111",
  27278=>"001011000",
  27279=>"110110101",
  27280=>"110011110",
  27281=>"100111000",
  27282=>"001110101",
  27283=>"100110110",
  27284=>"001100011",
  27285=>"101000101",
  27286=>"010010001",
  27287=>"111110001",
  27288=>"001101111",
  27289=>"101100100",
  27290=>"010110001",
  27291=>"100001001",
  27292=>"000100001",
  27293=>"110001011",
  27294=>"001010101",
  27295=>"001000000",
  27296=>"010010011",
  27297=>"011101100",
  27298=>"100111001",
  27299=>"111001101",
  27300=>"010101011",
  27301=>"111011100",
  27302=>"010000110",
  27303=>"011111011",
  27304=>"011101000",
  27305=>"011000101",
  27306=>"011000001",
  27307=>"100101000",
  27308=>"110010100",
  27309=>"100000001",
  27310=>"011100001",
  27311=>"111100000",
  27312=>"000010100",
  27313=>"001110110",
  27314=>"110011111",
  27315=>"010001111",
  27316=>"001110101",
  27317=>"010010111",
  27318=>"000110010",
  27319=>"101000011",
  27320=>"001011010",
  27321=>"100111011",
  27322=>"010011001",
  27323=>"001111100",
  27324=>"110000101",
  27325=>"000010000",
  27326=>"000010010",
  27327=>"001100111",
  27328=>"000111010",
  27329=>"111101111",
  27330=>"000001010",
  27331=>"101110100",
  27332=>"010101001",
  27333=>"010110101",
  27334=>"100111100",
  27335=>"000101110",
  27336=>"010010110",
  27337=>"010101001",
  27338=>"100100011",
  27339=>"000010000",
  27340=>"110101010",
  27341=>"000010011",
  27342=>"111110110",
  27343=>"100010000",
  27344=>"000000000",
  27345=>"001001110",
  27346=>"000001101",
  27347=>"100011010",
  27348=>"110110001",
  27349=>"110001001",
  27350=>"010111110",
  27351=>"000110101",
  27352=>"011101001",
  27353=>"110010011",
  27354=>"001110010",
  27355=>"011111111",
  27356=>"101101100",
  27357=>"111000000",
  27358=>"101100000",
  27359=>"001111001",
  27360=>"101010011",
  27361=>"101110110",
  27362=>"011111011",
  27363=>"011100100",
  27364=>"111011111",
  27365=>"101000010",
  27366=>"011100111",
  27367=>"110100101",
  27368=>"110000100",
  27369=>"100010100",
  27370=>"010111010",
  27371=>"101011011",
  27372=>"100101010",
  27373=>"010100111",
  27374=>"100111010",
  27375=>"000011110",
  27376=>"110101111",
  27377=>"011101001",
  27378=>"101111100",
  27379=>"000001000",
  27380=>"001101101",
  27381=>"101110011",
  27382=>"100000101",
  27383=>"111110110",
  27384=>"010000010",
  27385=>"001011001",
  27386=>"000010001",
  27387=>"011100001",
  27388=>"100011011",
  27389=>"011001100",
  27390=>"101100000",
  27391=>"101011110",
  27392=>"010001000",
  27393=>"010010110",
  27394=>"000010110",
  27395=>"100000011",
  27396=>"011011101",
  27397=>"010000111",
  27398=>"000001111",
  27399=>"111000010",
  27400=>"101000011",
  27401=>"000011101",
  27402=>"011000101",
  27403=>"000010001",
  27404=>"001010011",
  27405=>"111111000",
  27406=>"110001110",
  27407=>"011101001",
  27408=>"000110111",
  27409=>"011011000",
  27410=>"111011101",
  27411=>"110001100",
  27412=>"110111110",
  27413=>"101100111",
  27414=>"011000111",
  27415=>"101000010",
  27416=>"110110011",
  27417=>"001010110",
  27418=>"001000110",
  27419=>"010000001",
  27420=>"101110011",
  27421=>"011101101",
  27422=>"000000011",
  27423=>"001100111",
  27424=>"001110100",
  27425=>"011011110",
  27426=>"111010001",
  27427=>"001110110",
  27428=>"010100101",
  27429=>"010100011",
  27430=>"010011010",
  27431=>"101101001",
  27432=>"011000011",
  27433=>"101100110",
  27434=>"101111010",
  27435=>"111010010",
  27436=>"000000011",
  27437=>"000001010",
  27438=>"000000100",
  27439=>"010011111",
  27440=>"100110101",
  27441=>"000001111",
  27442=>"110111101",
  27443=>"010011110",
  27444=>"110001100",
  27445=>"100011011",
  27446=>"101010100",
  27447=>"010100010",
  27448=>"101010000",
  27449=>"100100000",
  27450=>"001110101",
  27451=>"100010101",
  27452=>"101000000",
  27453=>"111001010",
  27454=>"011001111",
  27455=>"111101101",
  27456=>"100000110",
  27457=>"111001101",
  27458=>"011110010",
  27459=>"100101101",
  27460=>"000010000",
  27461=>"101101010",
  27462=>"100110101",
  27463=>"100000100",
  27464=>"110011100",
  27465=>"000010101",
  27466=>"100011111",
  27467=>"111111110",
  27468=>"010111111",
  27469=>"111101010",
  27470=>"001111111",
  27471=>"000000111",
  27472=>"111011100",
  27473=>"001110110",
  27474=>"011000010",
  27475=>"111100001",
  27476=>"010000010",
  27477=>"011001001",
  27478=>"011110110",
  27479=>"111001101",
  27480=>"011000010",
  27481=>"100100110",
  27482=>"100110111",
  27483=>"011010101",
  27484=>"001101011",
  27485=>"101101001",
  27486=>"011101101",
  27487=>"001100100",
  27488=>"000000101",
  27489=>"101011011",
  27490=>"101110001",
  27491=>"101000011",
  27492=>"011100111",
  27493=>"011010001",
  27494=>"011100100",
  27495=>"010111110",
  27496=>"100010001",
  27497=>"001101101",
  27498=>"110011011",
  27499=>"001011001",
  27500=>"011010011",
  27501=>"101101011",
  27502=>"010101110",
  27503=>"001010000",
  27504=>"001100000",
  27505=>"010110010",
  27506=>"101010011",
  27507=>"000101110",
  27508=>"010111010",
  27509=>"100000101",
  27510=>"111111100",
  27511=>"000101100",
  27512=>"100000010",
  27513=>"001001011",
  27514=>"010001011",
  27515=>"010010011",
  27516=>"000101011",
  27517=>"010110000",
  27518=>"110101010",
  27519=>"100010111",
  27520=>"011100100",
  27521=>"100001000",
  27522=>"000010000",
  27523=>"110011010",
  27524=>"010001100",
  27525=>"000001010",
  27526=>"111000000",
  27527=>"000001111",
  27528=>"000011110",
  27529=>"000101110",
  27530=>"100110001",
  27531=>"111100011",
  27532=>"101110110",
  27533=>"111110100",
  27534=>"001100111",
  27535=>"111110010",
  27536=>"010101010",
  27537=>"111111011",
  27538=>"111111111",
  27539=>"000011101",
  27540=>"110100001",
  27541=>"001111100",
  27542=>"100100000",
  27543=>"101100001",
  27544=>"111110010",
  27545=>"000010010",
  27546=>"111110000",
  27547=>"010001010",
  27548=>"011001011",
  27549=>"100010101",
  27550=>"110001000",
  27551=>"011101010",
  27552=>"011011001",
  27553=>"110001111",
  27554=>"110101111",
  27555=>"111111101",
  27556=>"110000011",
  27557=>"101100111",
  27558=>"100110111",
  27559=>"001111000",
  27560=>"110101001",
  27561=>"001111011",
  27562=>"100011000",
  27563=>"111001000",
  27564=>"100000011",
  27565=>"010001101",
  27566=>"000101000",
  27567=>"001111010",
  27568=>"110100100",
  27569=>"011001000",
  27570=>"000001110",
  27571=>"001011101",
  27572=>"111001101",
  27573=>"111111111",
  27574=>"000111010",
  27575=>"101101100",
  27576=>"101011000",
  27577=>"100001110",
  27578=>"001000010",
  27579=>"111110001",
  27580=>"010110010",
  27581=>"100010100",
  27582=>"100111000",
  27583=>"111100100",
  27584=>"100110100",
  27585=>"110001000",
  27586=>"111111001",
  27587=>"110100110",
  27588=>"000100001",
  27589=>"101101101",
  27590=>"011100111",
  27591=>"110001001",
  27592=>"000000100",
  27593=>"010100110",
  27594=>"000111010",
  27595=>"111111110",
  27596=>"010101000",
  27597=>"001001001",
  27598=>"001000010",
  27599=>"000001000",
  27600=>"000000000",
  27601=>"110111111",
  27602=>"100001001",
  27603=>"101101011",
  27604=>"010111110",
  27605=>"100110010",
  27606=>"010001000",
  27607=>"100110100",
  27608=>"001000111",
  27609=>"100100011",
  27610=>"011110000",
  27611=>"011000110",
  27612=>"000011111",
  27613=>"101001000",
  27614=>"001101111",
  27615=>"000110100",
  27616=>"010000100",
  27617=>"101111011",
  27618=>"000001111",
  27619=>"010000100",
  27620=>"100010011",
  27621=>"111101011",
  27622=>"000100001",
  27623=>"110111111",
  27624=>"010000101",
  27625=>"101101000",
  27626=>"100000010",
  27627=>"111011000",
  27628=>"010001100",
  27629=>"110111101",
  27630=>"101100011",
  27631=>"001100100",
  27632=>"110101111",
  27633=>"010000101",
  27634=>"000111011",
  27635=>"010101010",
  27636=>"011000001",
  27637=>"101000000",
  27638=>"000111111",
  27639=>"101101101",
  27640=>"000100111",
  27641=>"000100101",
  27642=>"101101000",
  27643=>"011010011",
  27644=>"000100001",
  27645=>"010000111",
  27646=>"101100000",
  27647=>"111010011",
  27648=>"111100011",
  27649=>"111100010",
  27650=>"110101101",
  27651=>"110110010",
  27652=>"011000001",
  27653=>"010101110",
  27654=>"000100110",
  27655=>"110001000",
  27656=>"010111000",
  27657=>"111101101",
  27658=>"011110100",
  27659=>"101110110",
  27660=>"100100010",
  27661=>"010010110",
  27662=>"000101010",
  27663=>"110110001",
  27664=>"010100100",
  27665=>"001111111",
  27666=>"000100111",
  27667=>"010111010",
  27668=>"111111101",
  27669=>"000001101",
  27670=>"111111111",
  27671=>"101110110",
  27672=>"111101000",
  27673=>"010101101",
  27674=>"110001000",
  27675=>"101000110",
  27676=>"101110101",
  27677=>"111111000",
  27678=>"100100110",
  27679=>"000100011",
  27680=>"110000101",
  27681=>"010101100",
  27682=>"101000000",
  27683=>"010001100",
  27684=>"110111100",
  27685=>"100100111",
  27686=>"100101010",
  27687=>"101010110",
  27688=>"111101110",
  27689=>"000111111",
  27690=>"011111011",
  27691=>"000001010",
  27692=>"101010011",
  27693=>"010000001",
  27694=>"011001011",
  27695=>"111110110",
  27696=>"001000111",
  27697=>"101111011",
  27698=>"001010110",
  27699=>"001011100",
  27700=>"011110100",
  27701=>"001010110",
  27702=>"011001011",
  27703=>"001010010",
  27704=>"110101100",
  27705=>"100001110",
  27706=>"111110000",
  27707=>"101000000",
  27708=>"011111111",
  27709=>"010011001",
  27710=>"101100111",
  27711=>"000000101",
  27712=>"101101111",
  27713=>"111010100",
  27714=>"100000110",
  27715=>"100100110",
  27716=>"111001110",
  27717=>"101001010",
  27718=>"001100100",
  27719=>"101010010",
  27720=>"100000001",
  27721=>"110011110",
  27722=>"110101110",
  27723=>"111010010",
  27724=>"111000100",
  27725=>"011110100",
  27726=>"000011011",
  27727=>"101010000",
  27728=>"111111000",
  27729=>"001101111",
  27730=>"100000100",
  27731=>"010100011",
  27732=>"110001100",
  27733=>"111010000",
  27734=>"011000110",
  27735=>"001111001",
  27736=>"101111101",
  27737=>"111011101",
  27738=>"000010010",
  27739=>"010011001",
  27740=>"110110001",
  27741=>"000100010",
  27742=>"111001100",
  27743=>"001100011",
  27744=>"001001111",
  27745=>"100010110",
  27746=>"100110000",
  27747=>"000010000",
  27748=>"110010110",
  27749=>"011100000",
  27750=>"011011011",
  27751=>"011101011",
  27752=>"110100111",
  27753=>"111101111",
  27754=>"110001010",
  27755=>"100010110",
  27756=>"000011010",
  27757=>"111100110",
  27758=>"110000000",
  27759=>"111101100",
  27760=>"100001110",
  27761=>"111010010",
  27762=>"001100000",
  27763=>"001110110",
  27764=>"110100001",
  27765=>"011000010",
  27766=>"100001110",
  27767=>"110011100",
  27768=>"000010110",
  27769=>"110000101",
  27770=>"101001110",
  27771=>"100111111",
  27772=>"110010110",
  27773=>"011000110",
  27774=>"100100011",
  27775=>"011010000",
  27776=>"001110111",
  27777=>"110001000",
  27778=>"010011101",
  27779=>"001011000",
  27780=>"011011110",
  27781=>"111100110",
  27782=>"000100100",
  27783=>"110100110",
  27784=>"100110000",
  27785=>"111101000",
  27786=>"010110110",
  27787=>"100011110",
  27788=>"110000010",
  27789=>"100010101",
  27790=>"110011000",
  27791=>"110101110",
  27792=>"110100001",
  27793=>"011011010",
  27794=>"110011000",
  27795=>"011100101",
  27796=>"110101000",
  27797=>"000000111",
  27798=>"100110100",
  27799=>"111111101",
  27800=>"111010100",
  27801=>"110110101",
  27802=>"100001011",
  27803=>"000101100",
  27804=>"010110111",
  27805=>"010111011",
  27806=>"100101101",
  27807=>"110000111",
  27808=>"111110010",
  27809=>"110011101",
  27810=>"100110110",
  27811=>"101100101",
  27812=>"111100011",
  27813=>"111100011",
  27814=>"011010010",
  27815=>"101100001",
  27816=>"010111110",
  27817=>"000111001",
  27818=>"000100111",
  27819=>"110001100",
  27820=>"101101011",
  27821=>"001110111",
  27822=>"000110110",
  27823=>"101010010",
  27824=>"110011000",
  27825=>"100011111",
  27826=>"010001101",
  27827=>"000000111",
  27828=>"010101001",
  27829=>"100111101",
  27830=>"000001010",
  27831=>"001000101",
  27832=>"110111111",
  27833=>"000010010",
  27834=>"011000111",
  27835=>"010001011",
  27836=>"100100101",
  27837=>"011001100",
  27838=>"101010011",
  27839=>"010110111",
  27840=>"110011001",
  27841=>"010001110",
  27842=>"000100010",
  27843=>"101100001",
  27844=>"010011110",
  27845=>"011000010",
  27846=>"100111001",
  27847=>"010000110",
  27848=>"001001001",
  27849=>"001111101",
  27850=>"101010111",
  27851=>"001011010",
  27852=>"001111100",
  27853=>"101011100",
  27854=>"111111010",
  27855=>"000100001",
  27856=>"110000100",
  27857=>"100001010",
  27858=>"000110111",
  27859=>"111011101",
  27860=>"000111110",
  27861=>"101001010",
  27862=>"111011011",
  27863=>"110000101",
  27864=>"000010011",
  27865=>"101010101",
  27866=>"100110101",
  27867=>"111101011",
  27868=>"010011111",
  27869=>"110111111",
  27870=>"001001110",
  27871=>"101001111",
  27872=>"001100010",
  27873=>"010110111",
  27874=>"110101110",
  27875=>"111111010",
  27876=>"001000100",
  27877=>"000111010",
  27878=>"110000010",
  27879=>"010000111",
  27880=>"011011011",
  27881=>"011110101",
  27882=>"001101100",
  27883=>"001101100",
  27884=>"101000010",
  27885=>"010010100",
  27886=>"001001001",
  27887=>"010101011",
  27888=>"000100100",
  27889=>"101001101",
  27890=>"111010110",
  27891=>"001110000",
  27892=>"101101010",
  27893=>"000110001",
  27894=>"011111111",
  27895=>"010110000",
  27896=>"110100110",
  27897=>"000001000",
  27898=>"000101001",
  27899=>"000101100",
  27900=>"001010001",
  27901=>"001101100",
  27902=>"001011011",
  27903=>"010000000",
  27904=>"010010111",
  27905=>"100011001",
  27906=>"000110100",
  27907=>"011010010",
  27908=>"111101111",
  27909=>"011010010",
  27910=>"001111000",
  27911=>"111100101",
  27912=>"111001001",
  27913=>"000001001",
  27914=>"000010011",
  27915=>"000010011",
  27916=>"101000000",
  27917=>"001110011",
  27918=>"010101010",
  27919=>"110011111",
  27920=>"001000001",
  27921=>"010010011",
  27922=>"010101010",
  27923=>"110110101",
  27924=>"111110010",
  27925=>"001011110",
  27926=>"010010111",
  27927=>"100101010",
  27928=>"110101001",
  27929=>"000101111",
  27930=>"100110010",
  27931=>"101011011",
  27932=>"000110100",
  27933=>"000010010",
  27934=>"011000010",
  27935=>"011101010",
  27936=>"111111101",
  27937=>"100110101",
  27938=>"000010100",
  27939=>"110001110",
  27940=>"110000100",
  27941=>"100101100",
  27942=>"001101101",
  27943=>"101111000",
  27944=>"110110001",
  27945=>"101010000",
  27946=>"100001000",
  27947=>"011100001",
  27948=>"110001010",
  27949=>"010011110",
  27950=>"010010000",
  27951=>"011010101",
  27952=>"101110011",
  27953=>"100001111",
  27954=>"100000110",
  27955=>"010011010",
  27956=>"101000101",
  27957=>"000100001",
  27958=>"000110100",
  27959=>"010111101",
  27960=>"010110000",
  27961=>"001011110",
  27962=>"101011000",
  27963=>"111000010",
  27964=>"000100011",
  27965=>"000011011",
  27966=>"100011111",
  27967=>"101010111",
  27968=>"100100010",
  27969=>"110010110",
  27970=>"000100100",
  27971=>"111011010",
  27972=>"111010001",
  27973=>"010101111",
  27974=>"010001011",
  27975=>"001101000",
  27976=>"111001111",
  27977=>"011010000",
  27978=>"000111100",
  27979=>"000100110",
  27980=>"010001101",
  27981=>"011110011",
  27982=>"110111001",
  27983=>"000101111",
  27984=>"000111001",
  27985=>"010010111",
  27986=>"011001110",
  27987=>"101011111",
  27988=>"100011001",
  27989=>"010000101",
  27990=>"110001110",
  27991=>"110100111",
  27992=>"010000001",
  27993=>"000100110",
  27994=>"000101100",
  27995=>"010100100",
  27996=>"001011001",
  27997=>"000110011",
  27998=>"011010011",
  27999=>"001111010",
  28000=>"111100011",
  28001=>"011110000",
  28002=>"110001000",
  28003=>"100000110",
  28004=>"100100001",
  28005=>"110111000",
  28006=>"000001100",
  28007=>"000100111",
  28008=>"100111111",
  28009=>"110000100",
  28010=>"111101111",
  28011=>"111101111",
  28012=>"110010110",
  28013=>"110000110",
  28014=>"101100010",
  28015=>"000100101",
  28016=>"101100011",
  28017=>"000110100",
  28018=>"010111110",
  28019=>"101100001",
  28020=>"100000000",
  28021=>"011000010",
  28022=>"001000001",
  28023=>"101101000",
  28024=>"110000000",
  28025=>"110101110",
  28026=>"000101110",
  28027=>"001110011",
  28028=>"110000000",
  28029=>"001000111",
  28030=>"111111100",
  28031=>"010000000",
  28032=>"011100110",
  28033=>"110001110",
  28034=>"001110111",
  28035=>"110110000",
  28036=>"111100000",
  28037=>"000111100",
  28038=>"100100111",
  28039=>"111110001",
  28040=>"010001110",
  28041=>"101011001",
  28042=>"011111111",
  28043=>"111001101",
  28044=>"011110111",
  28045=>"010000011",
  28046=>"000000100",
  28047=>"011011100",
  28048=>"101010110",
  28049=>"100101001",
  28050=>"001111010",
  28051=>"110111000",
  28052=>"111010000",
  28053=>"110110110",
  28054=>"010010111",
  28055=>"101001100",
  28056=>"111011100",
  28057=>"010110101",
  28058=>"110011011",
  28059=>"000101010",
  28060=>"100100011",
  28061=>"000001100",
  28062=>"000001010",
  28063=>"101000111",
  28064=>"000010110",
  28065=>"000010010",
  28066=>"111010000",
  28067=>"000010100",
  28068=>"000001100",
  28069=>"000000001",
  28070=>"000111110",
  28071=>"010111001",
  28072=>"010101101",
  28073=>"100110100",
  28074=>"000100000",
  28075=>"100010100",
  28076=>"100101110",
  28077=>"010000000",
  28078=>"101110001",
  28079=>"010110000",
  28080=>"100011011",
  28081=>"111110000",
  28082=>"110100111",
  28083=>"000111110",
  28084=>"001001010",
  28085=>"101110110",
  28086=>"010010010",
  28087=>"100000001",
  28088=>"110001001",
  28089=>"110101001",
  28090=>"100000110",
  28091=>"011111101",
  28092=>"001110011",
  28093=>"010101010",
  28094=>"111111010",
  28095=>"100001010",
  28096=>"101101101",
  28097=>"010010011",
  28098=>"110110000",
  28099=>"100001011",
  28100=>"101110000",
  28101=>"001110010",
  28102=>"111101111",
  28103=>"110101010",
  28104=>"111110010",
  28105=>"111100001",
  28106=>"110111110",
  28107=>"111111101",
  28108=>"110100001",
  28109=>"100001110",
  28110=>"111101101",
  28111=>"000001100",
  28112=>"110001111",
  28113=>"000100010",
  28114=>"001010011",
  28115=>"001000010",
  28116=>"101100101",
  28117=>"010111011",
  28118=>"000101101",
  28119=>"110100111",
  28120=>"010011100",
  28121=>"010001111",
  28122=>"000010011",
  28123=>"001100000",
  28124=>"110011101",
  28125=>"111000001",
  28126=>"011000110",
  28127=>"100011000",
  28128=>"000110101",
  28129=>"110100000",
  28130=>"100110000",
  28131=>"100011011",
  28132=>"101011110",
  28133=>"100001001",
  28134=>"001000100",
  28135=>"010001001",
  28136=>"011011010",
  28137=>"011101110",
  28138=>"000000100",
  28139=>"110010101",
  28140=>"110110110",
  28141=>"100101101",
  28142=>"000000110",
  28143=>"010001011",
  28144=>"000101101",
  28145=>"000010111",
  28146=>"001010110",
  28147=>"000011001",
  28148=>"101000111",
  28149=>"011111110",
  28150=>"000110111",
  28151=>"100110011",
  28152=>"001000000",
  28153=>"000101110",
  28154=>"010100010",
  28155=>"001010001",
  28156=>"000110100",
  28157=>"101100101",
  28158=>"100010101",
  28159=>"100011110",
  28160=>"101011101",
  28161=>"101010001",
  28162=>"010000010",
  28163=>"101110001",
  28164=>"011101101",
  28165=>"111110111",
  28166=>"011011001",
  28167=>"011110111",
  28168=>"110011010",
  28169=>"101101010",
  28170=>"100000111",
  28171=>"001100100",
  28172=>"011100101",
  28173=>"001001101",
  28174=>"011110010",
  28175=>"111001000",
  28176=>"010101110",
  28177=>"011111110",
  28178=>"100110111",
  28179=>"010000100",
  28180=>"000110111",
  28181=>"000011110",
  28182=>"100001101",
  28183=>"100011110",
  28184=>"100000110",
  28185=>"001000000",
  28186=>"011001011",
  28187=>"000100101",
  28188=>"000011100",
  28189=>"000011000",
  28190=>"010111001",
  28191=>"010011100",
  28192=>"100001001",
  28193=>"111101010",
  28194=>"100100011",
  28195=>"111111010",
  28196=>"101111010",
  28197=>"011011111",
  28198=>"010110011",
  28199=>"010111000",
  28200=>"010111001",
  28201=>"101010110",
  28202=>"101110100",
  28203=>"001111111",
  28204=>"111110011",
  28205=>"000100111",
  28206=>"011110110",
  28207=>"101001010",
  28208=>"010101100",
  28209=>"111111111",
  28210=>"100100000",
  28211=>"010111100",
  28212=>"000011010",
  28213=>"101001101",
  28214=>"010101110",
  28215=>"101101101",
  28216=>"000111101",
  28217=>"111111101",
  28218=>"110000110",
  28219=>"100011101",
  28220=>"011000101",
  28221=>"000011100",
  28222=>"110111010",
  28223=>"101110011",
  28224=>"111111101",
  28225=>"001111010",
  28226=>"100100010",
  28227=>"111010000",
  28228=>"010101101",
  28229=>"000011010",
  28230=>"100110100",
  28231=>"111011101",
  28232=>"000010110",
  28233=>"010100100",
  28234=>"111011010",
  28235=>"111111110",
  28236=>"001001010",
  28237=>"110010010",
  28238=>"101110101",
  28239=>"010011001",
  28240=>"011010010",
  28241=>"100100111",
  28242=>"001001111",
  28243=>"010010101",
  28244=>"101000001",
  28245=>"000101100",
  28246=>"101010100",
  28247=>"111110111",
  28248=>"101111111",
  28249=>"000111101",
  28250=>"000111111",
  28251=>"011111110",
  28252=>"100010000",
  28253=>"110000010",
  28254=>"010111111",
  28255=>"110101010",
  28256=>"010000000",
  28257=>"000011011",
  28258=>"011100011",
  28259=>"111100110",
  28260=>"110011011",
  28261=>"011110110",
  28262=>"010110010",
  28263=>"100000101",
  28264=>"000001001",
  28265=>"001101110",
  28266=>"100001010",
  28267=>"011100011",
  28268=>"110101010",
  28269=>"011010110",
  28270=>"100010011",
  28271=>"110010100",
  28272=>"111101000",
  28273=>"101000001",
  28274=>"111000011",
  28275=>"010101111",
  28276=>"000111111",
  28277=>"100010110",
  28278=>"100000111",
  28279=>"000010100",
  28280=>"010011110",
  28281=>"010011111",
  28282=>"000111001",
  28283=>"110000111",
  28284=>"111100100",
  28285=>"000010110",
  28286=>"010000111",
  28287=>"001010100",
  28288=>"000010010",
  28289=>"111011100",
  28290=>"001000100",
  28291=>"001101111",
  28292=>"000001001",
  28293=>"111110110",
  28294=>"011011010",
  28295=>"000101011",
  28296=>"000010100",
  28297=>"000111001",
  28298=>"000001101",
  28299=>"001111111",
  28300=>"110001010",
  28301=>"110110101",
  28302=>"001010000",
  28303=>"000100100",
  28304=>"001101101",
  28305=>"001110101",
  28306=>"001101110",
  28307=>"011000010",
  28308=>"101111000",
  28309=>"000001010",
  28310=>"111111101",
  28311=>"000100011",
  28312=>"100110000",
  28313=>"110101101",
  28314=>"011101000",
  28315=>"111000010",
  28316=>"111111010",
  28317=>"000100100",
  28318=>"000010000",
  28319=>"011001000",
  28320=>"101001000",
  28321=>"000000101",
  28322=>"001000011",
  28323=>"110011010",
  28324=>"101100001",
  28325=>"101100011",
  28326=>"111101010",
  28327=>"110010000",
  28328=>"000110000",
  28329=>"101100111",
  28330=>"111011000",
  28331=>"100000000",
  28332=>"110001000",
  28333=>"101011010",
  28334=>"101000000",
  28335=>"011100011",
  28336=>"010010001",
  28337=>"100011001",
  28338=>"001110111",
  28339=>"111101110",
  28340=>"110010100",
  28341=>"010101100",
  28342=>"010010100",
  28343=>"001011001",
  28344=>"101110011",
  28345=>"101010110",
  28346=>"001101111",
  28347=>"011100101",
  28348=>"000101110",
  28349=>"011110010",
  28350=>"101111100",
  28351=>"101000101",
  28352=>"110100110",
  28353=>"111011000",
  28354=>"111010110",
  28355=>"011101011",
  28356=>"000000010",
  28357=>"011011010",
  28358=>"010101010",
  28359=>"110001110",
  28360=>"011010000",
  28361=>"110110010",
  28362=>"010001010",
  28363=>"001011010",
  28364=>"011111110",
  28365=>"110111101",
  28366=>"101110101",
  28367=>"000010000",
  28368=>"111101100",
  28369=>"000011011",
  28370=>"111001100",
  28371=>"101100001",
  28372=>"101011001",
  28373=>"000110100",
  28374=>"101100011",
  28375=>"101001000",
  28376=>"010111011",
  28377=>"111110111",
  28378=>"100001111",
  28379=>"110011111",
  28380=>"110110010",
  28381=>"001100011",
  28382=>"011110010",
  28383=>"000110000",
  28384=>"001110111",
  28385=>"111110011",
  28386=>"001100110",
  28387=>"100011011",
  28388=>"000000110",
  28389=>"011000100",
  28390=>"011010000",
  28391=>"101011000",
  28392=>"110101100",
  28393=>"100100111",
  28394=>"101010101",
  28395=>"111101110",
  28396=>"100000000",
  28397=>"010000010",
  28398=>"011000001",
  28399=>"001000100",
  28400=>"100110011",
  28401=>"110010100",
  28402=>"101001100",
  28403=>"000011010",
  28404=>"011110000",
  28405=>"001101110",
  28406=>"011011001",
  28407=>"101011110",
  28408=>"011101011",
  28409=>"001110011",
  28410=>"000000101",
  28411=>"000101000",
  28412=>"011010101",
  28413=>"111101101",
  28414=>"100110110",
  28415=>"101001111",
  28416=>"001111011",
  28417=>"001000011",
  28418=>"110010011",
  28419=>"111101100",
  28420=>"010110101",
  28421=>"110101110",
  28422=>"000001110",
  28423=>"000101100",
  28424=>"010101010",
  28425=>"011000110",
  28426=>"111111110",
  28427=>"010111010",
  28428=>"001010011",
  28429=>"010101011",
  28430=>"010011001",
  28431=>"111110011",
  28432=>"111000101",
  28433=>"010011110",
  28434=>"101110001",
  28435=>"000100001",
  28436=>"010111000",
  28437=>"100011100",
  28438=>"000110011",
  28439=>"101111010",
  28440=>"000110000",
  28441=>"000001001",
  28442=>"000101111",
  28443=>"011011001",
  28444=>"111111101",
  28445=>"011110010",
  28446=>"101110000",
  28447=>"011111001",
  28448=>"001010010",
  28449=>"011110000",
  28450=>"110000011",
  28451=>"000010100",
  28452=>"001110001",
  28453=>"010010100",
  28454=>"100111011",
  28455=>"001110001",
  28456=>"010011000",
  28457=>"101101000",
  28458=>"111111000",
  28459=>"000001001",
  28460=>"111001101",
  28461=>"000110011",
  28462=>"011110110",
  28463=>"111011111",
  28464=>"101111011",
  28465=>"101100111",
  28466=>"100000100",
  28467=>"100001011",
  28468=>"000110111",
  28469=>"101000000",
  28470=>"011110110",
  28471=>"000010010",
  28472=>"111110000",
  28473=>"100010000",
  28474=>"000111101",
  28475=>"010010011",
  28476=>"011000100",
  28477=>"000011000",
  28478=>"011111100",
  28479=>"101010001",
  28480=>"101110000",
  28481=>"111111110",
  28482=>"000001011",
  28483=>"100010010",
  28484=>"010011001",
  28485=>"000001111",
  28486=>"100011101",
  28487=>"100110010",
  28488=>"010101010",
  28489=>"110100011",
  28490=>"110100101",
  28491=>"000001001",
  28492=>"011001000",
  28493=>"100101111",
  28494=>"100000110",
  28495=>"111110001",
  28496=>"011100110",
  28497=>"000001100",
  28498=>"000100011",
  28499=>"000111000",
  28500=>"100010010",
  28501=>"101011001",
  28502=>"001000000",
  28503=>"111101011",
  28504=>"010110101",
  28505=>"110011011",
  28506=>"100110011",
  28507=>"010100100",
  28508=>"010001100",
  28509=>"110111111",
  28510=>"100000100",
  28511=>"010001111",
  28512=>"010011111",
  28513=>"101001000",
  28514=>"000110111",
  28515=>"100011101",
  28516=>"111110010",
  28517=>"101110001",
  28518=>"101000001",
  28519=>"100001110",
  28520=>"110000100",
  28521=>"011101101",
  28522=>"110101001",
  28523=>"000001100",
  28524=>"001001111",
  28525=>"000001010",
  28526=>"010011000",
  28527=>"100000101",
  28528=>"011000000",
  28529=>"010101001",
  28530=>"110000010",
  28531=>"100110010",
  28532=>"001000000",
  28533=>"000100101",
  28534=>"010001111",
  28535=>"101011110",
  28536=>"000010100",
  28537=>"011010011",
  28538=>"001101100",
  28539=>"001000111",
  28540=>"000001000",
  28541=>"100101011",
  28542=>"011001010",
  28543=>"001000011",
  28544=>"000100101",
  28545=>"010010100",
  28546=>"111100110",
  28547=>"000011100",
  28548=>"101010100",
  28549=>"100001101",
  28550=>"100001000",
  28551=>"101100111",
  28552=>"001001101",
  28553=>"100101111",
  28554=>"000110110",
  28555=>"000010001",
  28556=>"010010001",
  28557=>"010110010",
  28558=>"110110010",
  28559=>"101111110",
  28560=>"011101010",
  28561=>"101111110",
  28562=>"000000001",
  28563=>"100100000",
  28564=>"000110011",
  28565=>"100101110",
  28566=>"011101110",
  28567=>"101001011",
  28568=>"010000101",
  28569=>"000111000",
  28570=>"101000100",
  28571=>"000111000",
  28572=>"111000011",
  28573=>"101101101",
  28574=>"110101000",
  28575=>"001010000",
  28576=>"010110010",
  28577=>"011010110",
  28578=>"010001000",
  28579=>"011011011",
  28580=>"010100010",
  28581=>"101001111",
  28582=>"000111101",
  28583=>"001111101",
  28584=>"000010101",
  28585=>"000000001",
  28586=>"001010000",
  28587=>"111101000",
  28588=>"101011100",
  28589=>"000001010",
  28590=>"000000001",
  28591=>"101001101",
  28592=>"101100011",
  28593=>"001111001",
  28594=>"101000100",
  28595=>"101101100",
  28596=>"100001111",
  28597=>"100010010",
  28598=>"011010100",
  28599=>"110110011",
  28600=>"011111110",
  28601=>"010101111",
  28602=>"001101111",
  28603=>"001101101",
  28604=>"010000010",
  28605=>"101010011",
  28606=>"101101110",
  28607=>"110100110",
  28608=>"010011011",
  28609=>"100011100",
  28610=>"111100110",
  28611=>"010011100",
  28612=>"110000110",
  28613=>"001100011",
  28614=>"010010000",
  28615=>"000110111",
  28616=>"110001110",
  28617=>"000111001",
  28618=>"110100011",
  28619=>"000000100",
  28620=>"000010001",
  28621=>"010000000",
  28622=>"000101010",
  28623=>"101111001",
  28624=>"010000110",
  28625=>"111001110",
  28626=>"101110010",
  28627=>"000110011",
  28628=>"001101011",
  28629=>"011100010",
  28630=>"100100001",
  28631=>"000101100",
  28632=>"110101010",
  28633=>"000010111",
  28634=>"111000110",
  28635=>"101100001",
  28636=>"110010000",
  28637=>"010000110",
  28638=>"010101001",
  28639=>"100001000",
  28640=>"111010011",
  28641=>"011110111",
  28642=>"111110010",
  28643=>"101000100",
  28644=>"001110100",
  28645=>"001111110",
  28646=>"110011011",
  28647=>"011011000",
  28648=>"110001011",
  28649=>"100100111",
  28650=>"111000010",
  28651=>"000100000",
  28652=>"110011100",
  28653=>"111110011",
  28654=>"100100011",
  28655=>"001111000",
  28656=>"010010011",
  28657=>"001011010",
  28658=>"010000101",
  28659=>"010100101",
  28660=>"000100000",
  28661=>"000101100",
  28662=>"101111101",
  28663=>"100101001",
  28664=>"111110100",
  28665=>"111011001",
  28666=>"100000010",
  28667=>"011101011",
  28668=>"100100001",
  28669=>"010100110",
  28670=>"000001000",
  28671=>"001100010",
  28672=>"001000000",
  28673=>"100000001",
  28674=>"000101001",
  28675=>"110101100",
  28676=>"011010011",
  28677=>"100100001",
  28678=>"100110110",
  28679=>"100010101",
  28680=>"111110111",
  28681=>"001010000",
  28682=>"001010010",
  28683=>"011011001",
  28684=>"001101001",
  28685=>"011001011",
  28686=>"110000101",
  28687=>"100001001",
  28688=>"100010100",
  28689=>"110011100",
  28690=>"010000010",
  28691=>"100111000",
  28692=>"010000010",
  28693=>"110110011",
  28694=>"101100001",
  28695=>"001001100",
  28696=>"000100111",
  28697=>"011011010",
  28698=>"010001110",
  28699=>"101010000",
  28700=>"110000000",
  28701=>"001000001",
  28702=>"101000011",
  28703=>"110111011",
  28704=>"010011000",
  28705=>"101000010",
  28706=>"011001000",
  28707=>"010000110",
  28708=>"000011100",
  28709=>"001111110",
  28710=>"101011011",
  28711=>"101101000",
  28712=>"111111000",
  28713=>"011001100",
  28714=>"011000100",
  28715=>"101011100",
  28716=>"110110000",
  28717=>"011001001",
  28718=>"000010110",
  28719=>"101010010",
  28720=>"000100100",
  28721=>"011001111",
  28722=>"100101011",
  28723=>"110100101",
  28724=>"111000000",
  28725=>"111110100",
  28726=>"001100011",
  28727=>"111011011",
  28728=>"011011000",
  28729=>"001111110",
  28730=>"001110110",
  28731=>"101011001",
  28732=>"100010100",
  28733=>"011010001",
  28734=>"111110101",
  28735=>"001100101",
  28736=>"001010010",
  28737=>"000001001",
  28738=>"001000101",
  28739=>"000100101",
  28740=>"100001000",
  28741=>"011110111",
  28742=>"111011100",
  28743=>"010010001",
  28744=>"011100101",
  28745=>"111110000",
  28746=>"100000000",
  28747=>"000001100",
  28748=>"010010101",
  28749=>"010010011",
  28750=>"101110011",
  28751=>"110001001",
  28752=>"000000001",
  28753=>"001110111",
  28754=>"111111111",
  28755=>"000001110",
  28756=>"110100101",
  28757=>"110110001",
  28758=>"011001010",
  28759=>"111100011",
  28760=>"011011100",
  28761=>"010001100",
  28762=>"111110010",
  28763=>"110011000",
  28764=>"110101111",
  28765=>"110111101",
  28766=>"010101111",
  28767=>"111101011",
  28768=>"100111011",
  28769=>"100011100",
  28770=>"111001010",
  28771=>"111010110",
  28772=>"011101110",
  28773=>"001100110",
  28774=>"110101010",
  28775=>"100111110",
  28776=>"010100011",
  28777=>"010100110",
  28778=>"000000010",
  28779=>"101000000",
  28780=>"000000100",
  28781=>"111101001",
  28782=>"111111111",
  28783=>"100001010",
  28784=>"101111010",
  28785=>"111100000",
  28786=>"001101010",
  28787=>"000110100",
  28788=>"011111110",
  28789=>"010100101",
  28790=>"000100111",
  28791=>"100000001",
  28792=>"110000111",
  28793=>"101001010",
  28794=>"010011110",
  28795=>"010110000",
  28796=>"111001100",
  28797=>"110101001",
  28798=>"100100010",
  28799=>"010111111",
  28800=>"110101001",
  28801=>"100101000",
  28802=>"111110101",
  28803=>"011001100",
  28804=>"000001110",
  28805=>"011000111",
  28806=>"011101001",
  28807=>"000100100",
  28808=>"111111001",
  28809=>"001000000",
  28810=>"111111101",
  28811=>"100010011",
  28812=>"100110010",
  28813=>"011110101",
  28814=>"000000100",
  28815=>"101010111",
  28816=>"110010100",
  28817=>"000100000",
  28818=>"001011011",
  28819=>"000110001",
  28820=>"100100001",
  28821=>"100000110",
  28822=>"001001101",
  28823=>"000000111",
  28824=>"011100011",
  28825=>"101001010",
  28826=>"100111011",
  28827=>"000000000",
  28828=>"001000010",
  28829=>"101010001",
  28830=>"101111000",
  28831=>"100011000",
  28832=>"101100101",
  28833=>"001100001",
  28834=>"011010011",
  28835=>"011000100",
  28836=>"101000000",
  28837=>"001000100",
  28838=>"010111100",
  28839=>"110010101",
  28840=>"101000001",
  28841=>"110001001",
  28842=>"000000101",
  28843=>"000100111",
  28844=>"101100101",
  28845=>"000010110",
  28846=>"111111111",
  28847=>"100010001",
  28848=>"111100111",
  28849=>"111111000",
  28850=>"011111001",
  28851=>"101000100",
  28852=>"011011000",
  28853=>"110110110",
  28854=>"110000011",
  28855=>"110110001",
  28856=>"000111011",
  28857=>"101101111",
  28858=>"011001000",
  28859=>"010011010",
  28860=>"010101001",
  28861=>"001010111",
  28862=>"001100000",
  28863=>"100000000",
  28864=>"100101000",
  28865=>"100010011",
  28866=>"110110000",
  28867=>"000101011",
  28868=>"101011100",
  28869=>"010110111",
  28870=>"010000010",
  28871=>"100001010",
  28872=>"001101100",
  28873=>"011000010",
  28874=>"011100011",
  28875=>"001000000",
  28876=>"101100001",
  28877=>"101010111",
  28878=>"011001010",
  28879=>"000010110",
  28880=>"011110001",
  28881=>"111110000",
  28882=>"011001100",
  28883=>"101001001",
  28884=>"001101010",
  28885=>"101101100",
  28886=>"000111101",
  28887=>"001000101",
  28888=>"111011001",
  28889=>"100110000",
  28890=>"100011111",
  28891=>"010101011",
  28892=>"111110100",
  28893=>"111001000",
  28894=>"110110100",
  28895=>"110011000",
  28896=>"011011001",
  28897=>"100001100",
  28898=>"110010111",
  28899=>"000110101",
  28900=>"001000011",
  28901=>"100010101",
  28902=>"111101101",
  28903=>"001100000",
  28904=>"011111001",
  28905=>"010101000",
  28906=>"111101111",
  28907=>"100101101",
  28908=>"001001000",
  28909=>"000011111",
  28910=>"001001100",
  28911=>"000010001",
  28912=>"101110000",
  28913=>"101110001",
  28914=>"011011110",
  28915=>"000011010",
  28916=>"011111000",
  28917=>"111111001",
  28918=>"101101000",
  28919=>"111111111",
  28920=>"010111010",
  28921=>"111111110",
  28922=>"011010000",
  28923=>"111101011",
  28924=>"100010011",
  28925=>"000000000",
  28926=>"101111111",
  28927=>"010110000",
  28928=>"001001110",
  28929=>"011001010",
  28930=>"100000100",
  28931=>"001110101",
  28932=>"000000100",
  28933=>"010111011",
  28934=>"110000110",
  28935=>"101001111",
  28936=>"100001010",
  28937=>"010010001",
  28938=>"110110011",
  28939=>"110010011",
  28940=>"010010010",
  28941=>"010001111",
  28942=>"101110111",
  28943=>"101100011",
  28944=>"010101111",
  28945=>"101001111",
  28946=>"000101000",
  28947=>"101111111",
  28948=>"000011001",
  28949=>"011100001",
  28950=>"011101110",
  28951=>"010010000",
  28952=>"110110110",
  28953=>"110000111",
  28954=>"111110110",
  28955=>"100101101",
  28956=>"010000110",
  28957=>"100001101",
  28958=>"110111001",
  28959=>"001000010",
  28960=>"000000010",
  28961=>"011111011",
  28962=>"001000010",
  28963=>"110011000",
  28964=>"111001011",
  28965=>"011110011",
  28966=>"111100110",
  28967=>"111110110",
  28968=>"110110101",
  28969=>"111001111",
  28970=>"110010101",
  28971=>"001110000",
  28972=>"000001110",
  28973=>"011011100",
  28974=>"011101101",
  28975=>"000111101",
  28976=>"010000000",
  28977=>"000100001",
  28978=>"011101011",
  28979=>"001010001",
  28980=>"110000100",
  28981=>"011111011",
  28982=>"000101111",
  28983=>"110100110",
  28984=>"100001010",
  28985=>"100101001",
  28986=>"110110101",
  28987=>"110010111",
  28988=>"000111100",
  28989=>"000001010",
  28990=>"111101001",
  28991=>"010001111",
  28992=>"111100101",
  28993=>"111001011",
  28994=>"100000100",
  28995=>"000111111",
  28996=>"011000000",
  28997=>"110000111",
  28998=>"001110111",
  28999=>"010010100",
  29000=>"001011100",
  29001=>"011101100",
  29002=>"110101001",
  29003=>"001100011",
  29004=>"000001000",
  29005=>"010111101",
  29006=>"100110000",
  29007=>"011010001",
  29008=>"000011011",
  29009=>"001111000",
  29010=>"001110010",
  29011=>"101000000",
  29012=>"011110010",
  29013=>"011001100",
  29014=>"101111000",
  29015=>"101111010",
  29016=>"100101001",
  29017=>"101001101",
  29018=>"101110110",
  29019=>"001111001",
  29020=>"010001011",
  29021=>"110000100",
  29022=>"001010001",
  29023=>"110100011",
  29024=>"101110101",
  29025=>"001100010",
  29026=>"111000101",
  29027=>"111101001",
  29028=>"110000101",
  29029=>"010001010",
  29030=>"101000000",
  29031=>"001000001",
  29032=>"010000001",
  29033=>"010101110",
  29034=>"001100010",
  29035=>"000110010",
  29036=>"111110010",
  29037=>"011101001",
  29038=>"010110110",
  29039=>"110001100",
  29040=>"111011100",
  29041=>"111010010",
  29042=>"100100010",
  29043=>"101100111",
  29044=>"101101101",
  29045=>"110001000",
  29046=>"001100001",
  29047=>"110111111",
  29048=>"100101000",
  29049=>"111000111",
  29050=>"100010000",
  29051=>"100100100",
  29052=>"101000001",
  29053=>"110011101",
  29054=>"110001001",
  29055=>"001110100",
  29056=>"000111000",
  29057=>"000011110",
  29058=>"010000000",
  29059=>"010111011",
  29060=>"001111001",
  29061=>"010010001",
  29062=>"101100000",
  29063=>"000011011",
  29064=>"011110000",
  29065=>"110000100",
  29066=>"100000000",
  29067=>"011111000",
  29068=>"110000100",
  29069=>"011010101",
  29070=>"011011101",
  29071=>"010110010",
  29072=>"000110100",
  29073=>"100001110",
  29074=>"000001000",
  29075=>"110111011",
  29076=>"101100100",
  29077=>"001101110",
  29078=>"101010000",
  29079=>"111001001",
  29080=>"111101110",
  29081=>"011000100",
  29082=>"011010101",
  29083=>"110100000",
  29084=>"110100101",
  29085=>"000000100",
  29086=>"100011011",
  29087=>"110011100",
  29088=>"111111001",
  29089=>"000011101",
  29090=>"111001000",
  29091=>"010000100",
  29092=>"100001110",
  29093=>"100111111",
  29094=>"101111011",
  29095=>"001001010",
  29096=>"101110010",
  29097=>"111101010",
  29098=>"111101111",
  29099=>"100110110",
  29100=>"101010110",
  29101=>"100110010",
  29102=>"110100010",
  29103=>"110000010",
  29104=>"111001111",
  29105=>"100001011",
  29106=>"111000011",
  29107=>"001110100",
  29108=>"010010101",
  29109=>"010010010",
  29110=>"100100010",
  29111=>"100000000",
  29112=>"111000011",
  29113=>"111100100",
  29114=>"000001101",
  29115=>"011001101",
  29116=>"111001111",
  29117=>"110001001",
  29118=>"100101000",
  29119=>"011100011",
  29120=>"110110111",
  29121=>"111111101",
  29122=>"110110111",
  29123=>"110111010",
  29124=>"111001110",
  29125=>"100011110",
  29126=>"001001011",
  29127=>"001100100",
  29128=>"000011001",
  29129=>"100011000",
  29130=>"011111011",
  29131=>"000110100",
  29132=>"001001000",
  29133=>"011010010",
  29134=>"011101111",
  29135=>"111100111",
  29136=>"100001111",
  29137=>"110100010",
  29138=>"011000001",
  29139=>"000111010",
  29140=>"011101001",
  29141=>"111001100",
  29142=>"001011101",
  29143=>"000011010",
  29144=>"001010100",
  29145=>"100011110",
  29146=>"011100010",
  29147=>"101001101",
  29148=>"100100000",
  29149=>"001001101",
  29150=>"001001101",
  29151=>"110101101",
  29152=>"001001110",
  29153=>"011011100",
  29154=>"100011000",
  29155=>"100101101",
  29156=>"000111000",
  29157=>"011001001",
  29158=>"111110101",
  29159=>"111000001",
  29160=>"101111111",
  29161=>"010000110",
  29162=>"001000101",
  29163=>"011110101",
  29164=>"111000000",
  29165=>"100101110",
  29166=>"011110101",
  29167=>"001101101",
  29168=>"011100101",
  29169=>"010111111",
  29170=>"001110111",
  29171=>"101011000",
  29172=>"011100110",
  29173=>"111000011",
  29174=>"010100101",
  29175=>"100111000",
  29176=>"000100101",
  29177=>"110110100",
  29178=>"001110101",
  29179=>"111000110",
  29180=>"100001111",
  29181=>"000110011",
  29182=>"000001110",
  29183=>"011111111",
  29184=>"110001100",
  29185=>"101110110",
  29186=>"110111101",
  29187=>"001110001",
  29188=>"110001101",
  29189=>"001101111",
  29190=>"111001011",
  29191=>"100111101",
  29192=>"010011101",
  29193=>"001101111",
  29194=>"111111111",
  29195=>"101010110",
  29196=>"011000100",
  29197=>"000011101",
  29198=>"111111010",
  29199=>"110000000",
  29200=>"001111000",
  29201=>"111000000",
  29202=>"111011101",
  29203=>"101010010",
  29204=>"110111000",
  29205=>"110101111",
  29206=>"011111111",
  29207=>"010010001",
  29208=>"011000100",
  29209=>"110011111",
  29210=>"101011110",
  29211=>"110000001",
  29212=>"001100010",
  29213=>"111000111",
  29214=>"010000110",
  29215=>"101011110",
  29216=>"000001100",
  29217=>"000101000",
  29218=>"000100110",
  29219=>"111101001",
  29220=>"010011111",
  29221=>"110101001",
  29222=>"100100101",
  29223=>"111110111",
  29224=>"111000001",
  29225=>"000100111",
  29226=>"010101001",
  29227=>"001001101",
  29228=>"010111001",
  29229=>"001101101",
  29230=>"001010000",
  29231=>"111110010",
  29232=>"111101011",
  29233=>"101010010",
  29234=>"000110110",
  29235=>"010001101",
  29236=>"011010001",
  29237=>"001010011",
  29238=>"001000011",
  29239=>"111001010",
  29240=>"010111000",
  29241=>"000001110",
  29242=>"000101110",
  29243=>"010001000",
  29244=>"011101111",
  29245=>"000101100",
  29246=>"111101111",
  29247=>"101001001",
  29248=>"010000111",
  29249=>"100100110",
  29250=>"010000101",
  29251=>"001001010",
  29252=>"111111101",
  29253=>"011110100",
  29254=>"010011001",
  29255=>"000011100",
  29256=>"000000100",
  29257=>"010001101",
  29258=>"001000000",
  29259=>"000100101",
  29260=>"101001011",
  29261=>"001001010",
  29262=>"000000111",
  29263=>"010110110",
  29264=>"010101101",
  29265=>"000000111",
  29266=>"011010011",
  29267=>"101000010",
  29268=>"101001010",
  29269=>"111010110",
  29270=>"000010111",
  29271=>"011111000",
  29272=>"000011010",
  29273=>"110100001",
  29274=>"100100000",
  29275=>"111011011",
  29276=>"010110000",
  29277=>"101111110",
  29278=>"111111111",
  29279=>"010100001",
  29280=>"110010100",
  29281=>"110111010",
  29282=>"111101001",
  29283=>"010001101",
  29284=>"010101100",
  29285=>"000100110",
  29286=>"101011010",
  29287=>"011010011",
  29288=>"101011001",
  29289=>"001101110",
  29290=>"000111011",
  29291=>"010000110",
  29292=>"001001000",
  29293=>"101110100",
  29294=>"100001001",
  29295=>"100110101",
  29296=>"000000011",
  29297=>"010101110",
  29298=>"100001010",
  29299=>"000010010",
  29300=>"000000010",
  29301=>"110000010",
  29302=>"000001000",
  29303=>"110010000",
  29304=>"010110001",
  29305=>"010101110",
  29306=>"111001001",
  29307=>"110111111",
  29308=>"011101000",
  29309=>"111110010",
  29310=>"000101111",
  29311=>"111011010",
  29312=>"110100101",
  29313=>"000101000",
  29314=>"101111100",
  29315=>"001001110",
  29316=>"100011111",
  29317=>"110011100",
  29318=>"001101111",
  29319=>"011101111",
  29320=>"001000101",
  29321=>"000111011",
  29322=>"101010100",
  29323=>"111100011",
  29324=>"000010001",
  29325=>"101111100",
  29326=>"011110001",
  29327=>"110111100",
  29328=>"010010001",
  29329=>"111001000",
  29330=>"100101011",
  29331=>"111111111",
  29332=>"100101100",
  29333=>"101001111",
  29334=>"011001000",
  29335=>"110011111",
  29336=>"110101011",
  29337=>"100101110",
  29338=>"010001111",
  29339=>"100111111",
  29340=>"110111011",
  29341=>"101000000",
  29342=>"000110001",
  29343=>"111011110",
  29344=>"010010111",
  29345=>"001100101",
  29346=>"100101011",
  29347=>"100010011",
  29348=>"011011001",
  29349=>"000001111",
  29350=>"011100110",
  29351=>"100111101",
  29352=>"001011000",
  29353=>"111000010",
  29354=>"110110100",
  29355=>"010100100",
  29356=>"101101001",
  29357=>"000000001",
  29358=>"110000100",
  29359=>"001100010",
  29360=>"100011110",
  29361=>"101011101",
  29362=>"100000010",
  29363=>"010100000",
  29364=>"101001001",
  29365=>"011110100",
  29366=>"100000010",
  29367=>"010010011",
  29368=>"001101100",
  29369=>"110011000",
  29370=>"011111111",
  29371=>"001101100",
  29372=>"010100010",
  29373=>"110101100",
  29374=>"110000101",
  29375=>"111101010",
  29376=>"001011111",
  29377=>"001101110",
  29378=>"000001000",
  29379=>"101001111",
  29380=>"101101110",
  29381=>"111100101",
  29382=>"111100101",
  29383=>"101111110",
  29384=>"100111100",
  29385=>"010101100",
  29386=>"100100010",
  29387=>"111001000",
  29388=>"111110011",
  29389=>"000000101",
  29390=>"100001100",
  29391=>"000000100",
  29392=>"001110011",
  29393=>"100010011",
  29394=>"111110011",
  29395=>"000111100",
  29396=>"100110101",
  29397=>"111101100",
  29398=>"000110001",
  29399=>"010100100",
  29400=>"010100101",
  29401=>"001100100",
  29402=>"001010001",
  29403=>"110010110",
  29404=>"111111000",
  29405=>"011011101",
  29406=>"001011010",
  29407=>"100100011",
  29408=>"000111111",
  29409=>"111000101",
  29410=>"000111110",
  29411=>"001001010",
  29412=>"000001101",
  29413=>"100111001",
  29414=>"000000011",
  29415=>"010110110",
  29416=>"111010100",
  29417=>"011100100",
  29418=>"011111001",
  29419=>"010110110",
  29420=>"110010111",
  29421=>"001110100",
  29422=>"110100011",
  29423=>"111110001",
  29424=>"110101100",
  29425=>"000010110",
  29426=>"010000101",
  29427=>"001111011",
  29428=>"111111010",
  29429=>"111011110",
  29430=>"110011010",
  29431=>"111000000",
  29432=>"010101110",
  29433=>"010100111",
  29434=>"010101010",
  29435=>"110111000",
  29436=>"110001110",
  29437=>"111111000",
  29438=>"111110010",
  29439=>"010110100",
  29440=>"110111001",
  29441=>"010000100",
  29442=>"010100101",
  29443=>"101111111",
  29444=>"110101100",
  29445=>"001000101",
  29446=>"111010001",
  29447=>"001111000",
  29448=>"101001010",
  29449=>"011001111",
  29450=>"000000000",
  29451=>"101100001",
  29452=>"101010111",
  29453=>"010010011",
  29454=>"101000110",
  29455=>"111011111",
  29456=>"011000100",
  29457=>"011010110",
  29458=>"000000101",
  29459=>"101100010",
  29460=>"111111110",
  29461=>"111110100",
  29462=>"001110101",
  29463=>"111000100",
  29464=>"110011001",
  29465=>"000100100",
  29466=>"111101011",
  29467=>"111110100",
  29468=>"110100011",
  29469=>"011100001",
  29470=>"101011001",
  29471=>"100110011",
  29472=>"110001010",
  29473=>"111001110",
  29474=>"101100000",
  29475=>"001100011",
  29476=>"010110011",
  29477=>"110001000",
  29478=>"000011110",
  29479=>"001111000",
  29480=>"000001001",
  29481=>"000001101",
  29482=>"100100100",
  29483=>"110111111",
  29484=>"100001010",
  29485=>"011101001",
  29486=>"101111010",
  29487=>"100111000",
  29488=>"110110000",
  29489=>"001100111",
  29490=>"100110111",
  29491=>"100111011",
  29492=>"111110110",
  29493=>"100110100",
  29494=>"100110100",
  29495=>"110001000",
  29496=>"110001110",
  29497=>"011111101",
  29498=>"010001110",
  29499=>"010101000",
  29500=>"001101011",
  29501=>"111011011",
  29502=>"010011000",
  29503=>"111001010",
  29504=>"011000101",
  29505=>"001100101",
  29506=>"110010110",
  29507=>"111000101",
  29508=>"001110111",
  29509=>"100000100",
  29510=>"101001100",
  29511=>"000101100",
  29512=>"111000101",
  29513=>"000001000",
  29514=>"101101000",
  29515=>"000100111",
  29516=>"101101101",
  29517=>"100100001",
  29518=>"100110111",
  29519=>"000100011",
  29520=>"010101101",
  29521=>"010000011",
  29522=>"011011101",
  29523=>"111111011",
  29524=>"101111111",
  29525=>"010010101",
  29526=>"001011110",
  29527=>"011111101",
  29528=>"000000000",
  29529=>"101010011",
  29530=>"110100001",
  29531=>"001011111",
  29532=>"100010110",
  29533=>"011101000",
  29534=>"110000101",
  29535=>"111111110",
  29536=>"011011111",
  29537=>"110101010",
  29538=>"010011011",
  29539=>"110110100",
  29540=>"111110111",
  29541=>"011011011",
  29542=>"001000011",
  29543=>"111111110",
  29544=>"100011000",
  29545=>"000010110",
  29546=>"010111110",
  29547=>"000011111",
  29548=>"010100111",
  29549=>"100000000",
  29550=>"101001111",
  29551=>"010101100",
  29552=>"110100011",
  29553=>"110110111",
  29554=>"001001100",
  29555=>"110011000",
  29556=>"001011111",
  29557=>"000111100",
  29558=>"110100010",
  29559=>"101011011",
  29560=>"000111100",
  29561=>"110101000",
  29562=>"101100000",
  29563=>"011111000",
  29564=>"110100100",
  29565=>"110001111",
  29566=>"000101101",
  29567=>"100011111",
  29568=>"011110010",
  29569=>"111010100",
  29570=>"000001111",
  29571=>"111110001",
  29572=>"000010000",
  29573=>"111100011",
  29574=>"101000111",
  29575=>"000100010",
  29576=>"101010110",
  29577=>"001110000",
  29578=>"001001110",
  29579=>"100000010",
  29580=>"110010010",
  29581=>"011001101",
  29582=>"111110011",
  29583=>"101111111",
  29584=>"110100001",
  29585=>"101110111",
  29586=>"111001001",
  29587=>"111101111",
  29588=>"111011001",
  29589=>"001001010",
  29590=>"110100010",
  29591=>"011101111",
  29592=>"011010001",
  29593=>"100101110",
  29594=>"011000011",
  29595=>"011000011",
  29596=>"010010111",
  29597=>"110110000",
  29598=>"100001110",
  29599=>"001011001",
  29600=>"111111001",
  29601=>"011100100",
  29602=>"110100110",
  29603=>"110011110",
  29604=>"011000011",
  29605=>"011011100",
  29606=>"101111110",
  29607=>"110001101",
  29608=>"111100111",
  29609=>"000111111",
  29610=>"000111111",
  29611=>"110111001",
  29612=>"111101111",
  29613=>"000000110",
  29614=>"110001010",
  29615=>"101100101",
  29616=>"000011000",
  29617=>"011001111",
  29618=>"011111110",
  29619=>"000011111",
  29620=>"010000111",
  29621=>"001011111",
  29622=>"010000000",
  29623=>"001011101",
  29624=>"001100101",
  29625=>"011110101",
  29626=>"010000011",
  29627=>"100100100",
  29628=>"111001111",
  29629=>"011101111",
  29630=>"010011101",
  29631=>"110100100",
  29632=>"001111101",
  29633=>"000011111",
  29634=>"010000000",
  29635=>"110111010",
  29636=>"111100011",
  29637=>"010000100",
  29638=>"101100010",
  29639=>"110111110",
  29640=>"110110100",
  29641=>"001011110",
  29642=>"011011011",
  29643=>"000011101",
  29644=>"101000110",
  29645=>"101001110",
  29646=>"100100100",
  29647=>"110111011",
  29648=>"010011010",
  29649=>"010110100",
  29650=>"011011000",
  29651=>"000011001",
  29652=>"001000000",
  29653=>"000000101",
  29654=>"111110110",
  29655=>"000001100",
  29656=>"001011100",
  29657=>"111100111",
  29658=>"011001100",
  29659=>"001101111",
  29660=>"110000101",
  29661=>"001000111",
  29662=>"101111010",
  29663=>"110011110",
  29664=>"000101111",
  29665=>"000011001",
  29666=>"011101101",
  29667=>"100101100",
  29668=>"111111000",
  29669=>"110111001",
  29670=>"010110001",
  29671=>"111010100",
  29672=>"000100111",
  29673=>"011011010",
  29674=>"101001100",
  29675=>"011001100",
  29676=>"010110110",
  29677=>"111111010",
  29678=>"110111101",
  29679=>"101001000",
  29680=>"110101110",
  29681=>"111100101",
  29682=>"110110111",
  29683=>"000100000",
  29684=>"111111010",
  29685=>"100100101",
  29686=>"011011111",
  29687=>"011011001",
  29688=>"010000101",
  29689=>"011010001",
  29690=>"001000011",
  29691=>"011110001",
  29692=>"001100000",
  29693=>"011101001",
  29694=>"010010111",
  29695=>"111010000",
  29696=>"111100000",
  29697=>"010001011",
  29698=>"000001010",
  29699=>"111101110",
  29700=>"000101100",
  29701=>"111000011",
  29702=>"100010100",
  29703=>"000101110",
  29704=>"110000101",
  29705=>"011111010",
  29706=>"000101010",
  29707=>"100111001",
  29708=>"110001010",
  29709=>"110001111",
  29710=>"110110010",
  29711=>"111010101",
  29712=>"111101111",
  29713=>"000000001",
  29714=>"100010000",
  29715=>"100010111",
  29716=>"010001101",
  29717=>"111111101",
  29718=>"101010000",
  29719=>"101000110",
  29720=>"100000001",
  29721=>"101000001",
  29722=>"101100011",
  29723=>"100110000",
  29724=>"010011110",
  29725=>"100111101",
  29726=>"110010010",
  29727=>"111000101",
  29728=>"001001111",
  29729=>"000000111",
  29730=>"010010010",
  29731=>"111110100",
  29732=>"000011111",
  29733=>"110110000",
  29734=>"001100110",
  29735=>"001001011",
  29736=>"000110011",
  29737=>"000110111",
  29738=>"110110101",
  29739=>"000110110",
  29740=>"111110110",
  29741=>"111101110",
  29742=>"000111110",
  29743=>"001010100",
  29744=>"101111101",
  29745=>"111111010",
  29746=>"001000011",
  29747=>"000101000",
  29748=>"100000000",
  29749=>"011110001",
  29750=>"100011100",
  29751=>"111111010",
  29752=>"001100010",
  29753=>"100111011",
  29754=>"001001110",
  29755=>"111100111",
  29756=>"101011101",
  29757=>"110011011",
  29758=>"010000000",
  29759=>"010010001",
  29760=>"000111001",
  29761=>"101000010",
  29762=>"010000110",
  29763=>"101101000",
  29764=>"001100111",
  29765=>"011000010",
  29766=>"100000101",
  29767=>"101010110",
  29768=>"100001100",
  29769=>"010011100",
  29770=>"000010011",
  29771=>"000101110",
  29772=>"001001111",
  29773=>"101101111",
  29774=>"101111101",
  29775=>"010000000",
  29776=>"110000010",
  29777=>"010010000",
  29778=>"010000011",
  29779=>"101101111",
  29780=>"001111010",
  29781=>"000100000",
  29782=>"011011101",
  29783=>"111001010",
  29784=>"111101000",
  29785=>"100110011",
  29786=>"101101110",
  29787=>"001011011",
  29788=>"011010101",
  29789=>"100001001",
  29790=>"011000010",
  29791=>"111101100",
  29792=>"110000011",
  29793=>"001100010",
  29794=>"100000010",
  29795=>"100001110",
  29796=>"101100001",
  29797=>"001000011",
  29798=>"011010010",
  29799=>"000010110",
  29800=>"110101100",
  29801=>"000011011",
  29802=>"000010001",
  29803=>"011111101",
  29804=>"001110101",
  29805=>"111100101",
  29806=>"000100111",
  29807=>"111001111",
  29808=>"111000000",
  29809=>"011001100",
  29810=>"001110010",
  29811=>"000100111",
  29812=>"001111010",
  29813=>"100011010",
  29814=>"001100011",
  29815=>"010010100",
  29816=>"100101000",
  29817=>"100110010",
  29818=>"100101010",
  29819=>"100001010",
  29820=>"110001001",
  29821=>"110101001",
  29822=>"110111010",
  29823=>"011001111",
  29824=>"001000111",
  29825=>"111010111",
  29826=>"110101111",
  29827=>"101010100",
  29828=>"000010101",
  29829=>"000010110",
  29830=>"101010110",
  29831=>"011101101",
  29832=>"111101101",
  29833=>"111001111",
  29834=>"010110110",
  29835=>"000101111",
  29836=>"010000010",
  29837=>"011101101",
  29838=>"111001101",
  29839=>"110100111",
  29840=>"001110111",
  29841=>"101010001",
  29842=>"111111001",
  29843=>"101000111",
  29844=>"010101001",
  29845=>"101000101",
  29846=>"010000100",
  29847=>"001101111",
  29848=>"001010111",
  29849=>"010011010",
  29850=>"011111011",
  29851=>"000000000",
  29852=>"000111011",
  29853=>"110000101",
  29854=>"001111010",
  29855=>"101000111",
  29856=>"000111011",
  29857=>"001100011",
  29858=>"001101000",
  29859=>"100001010",
  29860=>"011101101",
  29861=>"101110110",
  29862=>"011110110",
  29863=>"000100000",
  29864=>"010010001",
  29865=>"010101100",
  29866=>"110000001",
  29867=>"011100001",
  29868=>"111101011",
  29869=>"111101110",
  29870=>"110000001",
  29871=>"011001011",
  29872=>"110010000",
  29873=>"010110000",
  29874=>"101011010",
  29875=>"001011000",
  29876=>"001111010",
  29877=>"101000000",
  29878=>"100100111",
  29879=>"001111000",
  29880=>"011101001",
  29881=>"000100001",
  29882=>"000110111",
  29883=>"000001111",
  29884=>"000011010",
  29885=>"110001110",
  29886=>"111100000",
  29887=>"100100010",
  29888=>"000010100",
  29889=>"000111011",
  29890=>"010010011",
  29891=>"100001000",
  29892=>"011101111",
  29893=>"001011000",
  29894=>"101011001",
  29895=>"101011000",
  29896=>"011100101",
  29897=>"000110001",
  29898=>"100101010",
  29899=>"011011011",
  29900=>"110011010",
  29901=>"011010000",
  29902=>"111011000",
  29903=>"100111110",
  29904=>"111111111",
  29905=>"101100101",
  29906=>"000101111",
  29907=>"010101001",
  29908=>"101001001",
  29909=>"100010000",
  29910=>"000010100",
  29911=>"111010110",
  29912=>"001010011",
  29913=>"000110000",
  29914=>"111001101",
  29915=>"110100000",
  29916=>"111010011",
  29917=>"101010111",
  29918=>"000101000",
  29919=>"011001001",
  29920=>"011011111",
  29921=>"000010111",
  29922=>"111101001",
  29923=>"110100110",
  29924=>"010100110",
  29925=>"100110100",
  29926=>"011101000",
  29927=>"010001000",
  29928=>"111100100",
  29929=>"011101101",
  29930=>"000101110",
  29931=>"110111111",
  29932=>"001001011",
  29933=>"001011100",
  29934=>"100100101",
  29935=>"110001110",
  29936=>"011110101",
  29937=>"110001001",
  29938=>"000010011",
  29939=>"010011011",
  29940=>"011001110",
  29941=>"010100100",
  29942=>"011000000",
  29943=>"000111111",
  29944=>"000100100",
  29945=>"001011001",
  29946=>"110111110",
  29947=>"100000011",
  29948=>"000101100",
  29949=>"011000000",
  29950=>"100011001",
  29951=>"001001111",
  29952=>"010101010",
  29953=>"111111011",
  29954=>"110111011",
  29955=>"001100001",
  29956=>"000011100",
  29957=>"110000111",
  29958=>"010000100",
  29959=>"001001001",
  29960=>"100001000",
  29961=>"101101011",
  29962=>"001110110",
  29963=>"001011000",
  29964=>"011111100",
  29965=>"011010010",
  29966=>"010110000",
  29967=>"000010110",
  29968=>"001110010",
  29969=>"100001011",
  29970=>"111110110",
  29971=>"111001000",
  29972=>"100101100",
  29973=>"111101101",
  29974=>"111110110",
  29975=>"000100000",
  29976=>"000010110",
  29977=>"111101001",
  29978=>"010000001",
  29979=>"010110010",
  29980=>"110011001",
  29981=>"100010110",
  29982=>"100110001",
  29983=>"101010010",
  29984=>"100110100",
  29985=>"101001110",
  29986=>"101101101",
  29987=>"000000000",
  29988=>"101101001",
  29989=>"100111111",
  29990=>"000001100",
  29991=>"111001101",
  29992=>"100110110",
  29993=>"101010101",
  29994=>"110011111",
  29995=>"011000011",
  29996=>"110101111",
  29997=>"011101101",
  29998=>"000000010",
  29999=>"101110011",
  30000=>"101100111",
  30001=>"011111000",
  30002=>"011101011",
  30003=>"011011010",
  30004=>"000101100",
  30005=>"100000011",
  30006=>"110100001",
  30007=>"011001010",
  30008=>"111111111",
  30009=>"010100110",
  30010=>"101100010",
  30011=>"001000001",
  30012=>"100011101",
  30013=>"001001000",
  30014=>"111011101",
  30015=>"011111111",
  30016=>"011010000",
  30017=>"111101111",
  30018=>"111110001",
  30019=>"001001010",
  30020=>"011110010",
  30021=>"010100000",
  30022=>"000001000",
  30023=>"101011101",
  30024=>"011110100",
  30025=>"010001101",
  30026=>"101100101",
  30027=>"101101011",
  30028=>"010011011",
  30029=>"011100100",
  30030=>"001111100",
  30031=>"110011010",
  30032=>"100011000",
  30033=>"100101111",
  30034=>"110101001",
  30035=>"111001000",
  30036=>"000000101",
  30037=>"000101111",
  30038=>"111010111",
  30039=>"000001111",
  30040=>"001000101",
  30041=>"001011010",
  30042=>"110000011",
  30043=>"100100111",
  30044=>"011000101",
  30045=>"001011010",
  30046=>"000111111",
  30047=>"001010010",
  30048=>"011011101",
  30049=>"011110100",
  30050=>"000101110",
  30051=>"000000011",
  30052=>"001010110",
  30053=>"000111100",
  30054=>"001110011",
  30055=>"001110011",
  30056=>"111100011",
  30057=>"000100000",
  30058=>"110111011",
  30059=>"011000110",
  30060=>"010010110",
  30061=>"111011000",
  30062=>"001000001",
  30063=>"101111101",
  30064=>"100101110",
  30065=>"011101010",
  30066=>"000001100",
  30067=>"110001000",
  30068=>"001101001",
  30069=>"011011110",
  30070=>"010011100",
  30071=>"011101010",
  30072=>"111011110",
  30073=>"111111100",
  30074=>"111100100",
  30075=>"110001100",
  30076=>"000000000",
  30077=>"110100101",
  30078=>"000101000",
  30079=>"111011010",
  30080=>"010110011",
  30081=>"111010111",
  30082=>"111100001",
  30083=>"100110011",
  30084=>"010100101",
  30085=>"110001111",
  30086=>"110101101",
  30087=>"100001110",
  30088=>"100100100",
  30089=>"011011101",
  30090=>"011110101",
  30091=>"101000111",
  30092=>"011010001",
  30093=>"111001111",
  30094=>"010011011",
  30095=>"111010101",
  30096=>"100000010",
  30097=>"110011000",
  30098=>"000110011",
  30099=>"001100111",
  30100=>"110110101",
  30101=>"101011110",
  30102=>"110101011",
  30103=>"000100010",
  30104=>"110111010",
  30105=>"000100100",
  30106=>"010111011",
  30107=>"101110100",
  30108=>"111101010",
  30109=>"000101000",
  30110=>"111001110",
  30111=>"011010101",
  30112=>"100110111",
  30113=>"110001111",
  30114=>"101101000",
  30115=>"000011101",
  30116=>"011101100",
  30117=>"101101011",
  30118=>"011110001",
  30119=>"110111111",
  30120=>"000000111",
  30121=>"001111110",
  30122=>"110000101",
  30123=>"111100101",
  30124=>"010101100",
  30125=>"010111100",
  30126=>"111100011",
  30127=>"110011110",
  30128=>"110111101",
  30129=>"010110000",
  30130=>"100000000",
  30131=>"111101110",
  30132=>"100110001",
  30133=>"010101001",
  30134=>"010101011",
  30135=>"011001001",
  30136=>"000101000",
  30137=>"110100111",
  30138=>"111110011",
  30139=>"010001011",
  30140=>"000011111",
  30141=>"011100101",
  30142=>"100011111",
  30143=>"001001011",
  30144=>"001001101",
  30145=>"010111100",
  30146=>"110101101",
  30147=>"000011100",
  30148=>"000100100",
  30149=>"000010000",
  30150=>"101000001",
  30151=>"001101101",
  30152=>"010001101",
  30153=>"001001100",
  30154=>"101110100",
  30155=>"100000010",
  30156=>"111010100",
  30157=>"101000011",
  30158=>"010000011",
  30159=>"110011011",
  30160=>"010110101",
  30161=>"101001110",
  30162=>"101011000",
  30163=>"000000011",
  30164=>"011100000",
  30165=>"011011011",
  30166=>"111000001",
  30167=>"000010010",
  30168=>"011001011",
  30169=>"010110110",
  30170=>"100000110",
  30171=>"111111101",
  30172=>"000010010",
  30173=>"001001110",
  30174=>"001011101",
  30175=>"111110110",
  30176=>"110101111",
  30177=>"100001100",
  30178=>"101011100",
  30179=>"011011110",
  30180=>"111001111",
  30181=>"000010010",
  30182=>"111001000",
  30183=>"000001110",
  30184=>"000010010",
  30185=>"100011001",
  30186=>"100000001",
  30187=>"001000101",
  30188=>"011101111",
  30189=>"111100111",
  30190=>"001000110",
  30191=>"001110001",
  30192=>"110100101",
  30193=>"100001110",
  30194=>"010111000",
  30195=>"001000010",
  30196=>"100101001",
  30197=>"100001010",
  30198=>"111000011",
  30199=>"100101001",
  30200=>"110000110",
  30201=>"111011100",
  30202=>"101000100",
  30203=>"110100110",
  30204=>"110011011",
  30205=>"100001111",
  30206=>"001000001",
  30207=>"010010001",
  30208=>"000101101",
  30209=>"010011000",
  30210=>"100001101",
  30211=>"000110100",
  30212=>"010010000",
  30213=>"000011001",
  30214=>"010001110",
  30215=>"100000001",
  30216=>"111110111",
  30217=>"101101110",
  30218=>"011001111",
  30219=>"110100000",
  30220=>"100111100",
  30221=>"101110111",
  30222=>"000010111",
  30223=>"001001111",
  30224=>"010100001",
  30225=>"011100111",
  30226=>"110110010",
  30227=>"010101010",
  30228=>"000010101",
  30229=>"101001010",
  30230=>"111001001",
  30231=>"000111110",
  30232=>"011001110",
  30233=>"101111101",
  30234=>"001111101",
  30235=>"000100011",
  30236=>"100011011",
  30237=>"100101000",
  30238=>"101111010",
  30239=>"001110001",
  30240=>"100010111",
  30241=>"100111111",
  30242=>"000100011",
  30243=>"100110001",
  30244=>"101101001",
  30245=>"101000011",
  30246=>"010111101",
  30247=>"111110010",
  30248=>"011011011",
  30249=>"111000101",
  30250=>"000111101",
  30251=>"001011100",
  30252=>"111101101",
  30253=>"000000000",
  30254=>"111011110",
  30255=>"111110010",
  30256=>"101110001",
  30257=>"110001100",
  30258=>"001011101",
  30259=>"110011000",
  30260=>"010010010",
  30261=>"001111001",
  30262=>"111010100",
  30263=>"100000101",
  30264=>"111011101",
  30265=>"001101110",
  30266=>"000001100",
  30267=>"001101011",
  30268=>"001010011",
  30269=>"110010100",
  30270=>"001001111",
  30271=>"100010011",
  30272=>"111010011",
  30273=>"001101001",
  30274=>"101110111",
  30275=>"001101110",
  30276=>"010000011",
  30277=>"010010000",
  30278=>"000001001",
  30279=>"100000000",
  30280=>"101101110",
  30281=>"010111101",
  30282=>"001010000",
  30283=>"111000011",
  30284=>"110010001",
  30285=>"010100010",
  30286=>"101000111",
  30287=>"111000101",
  30288=>"110110110",
  30289=>"001110100",
  30290=>"111011100",
  30291=>"000100001",
  30292=>"000101111",
  30293=>"001001111",
  30294=>"111110011",
  30295=>"011011000",
  30296=>"011100010",
  30297=>"010111100",
  30298=>"010101101",
  30299=>"110010111",
  30300=>"110000011",
  30301=>"011110100",
  30302=>"000001011",
  30303=>"100001110",
  30304=>"100111001",
  30305=>"110000111",
  30306=>"100011010",
  30307=>"100101111",
  30308=>"000100011",
  30309=>"000110101",
  30310=>"000111111",
  30311=>"001010000",
  30312=>"001111110",
  30313=>"011100010",
  30314=>"101111010",
  30315=>"001110010",
  30316=>"011011011",
  30317=>"110101101",
  30318=>"111111110",
  30319=>"011010011",
  30320=>"110001000",
  30321=>"100111111",
  30322=>"100010010",
  30323=>"100010001",
  30324=>"000000011",
  30325=>"010111000",
  30326=>"000000111",
  30327=>"000001011",
  30328=>"101111111",
  30329=>"000110100",
  30330=>"000110111",
  30331=>"000010111",
  30332=>"100011011",
  30333=>"011110101",
  30334=>"010111010",
  30335=>"101110110",
  30336=>"111110011",
  30337=>"011111011",
  30338=>"111011101",
  30339=>"000011101",
  30340=>"101100100",
  30341=>"101101101",
  30342=>"101111111",
  30343=>"100101001",
  30344=>"001100000",
  30345=>"010001100",
  30346=>"000010101",
  30347=>"101110101",
  30348=>"000100000",
  30349=>"100110111",
  30350=>"010111010",
  30351=>"110010111",
  30352=>"011001000",
  30353=>"110100111",
  30354=>"010100011",
  30355=>"000101111",
  30356=>"001111000",
  30357=>"001011101",
  30358=>"111100111",
  30359=>"100010001",
  30360=>"000010111",
  30361=>"100001011",
  30362=>"011100010",
  30363=>"000011011",
  30364=>"010011111",
  30365=>"111110011",
  30366=>"110111000",
  30367=>"001111000",
  30368=>"011001110",
  30369=>"111101101",
  30370=>"111011100",
  30371=>"010100101",
  30372=>"010010001",
  30373=>"101011110",
  30374=>"111001111",
  30375=>"010011101",
  30376=>"000000011",
  30377=>"111000011",
  30378=>"000100011",
  30379=>"101000001",
  30380=>"000000101",
  30381=>"000101000",
  30382=>"001100100",
  30383=>"011101000",
  30384=>"000101111",
  30385=>"010100110",
  30386=>"010110000",
  30387=>"001011100",
  30388=>"000010010",
  30389=>"101111100",
  30390=>"001111011",
  30391=>"101011011",
  30392=>"010010001",
  30393=>"111110011",
  30394=>"110010111",
  30395=>"100010000",
  30396=>"011111010",
  30397=>"001000010",
  30398=>"000010101",
  30399=>"100010001",
  30400=>"110101100",
  30401=>"111100100",
  30402=>"100100001",
  30403=>"011001000",
  30404=>"011101111",
  30405=>"100010010",
  30406=>"111010011",
  30407=>"011101110",
  30408=>"000101010",
  30409=>"011110010",
  30410=>"000001111",
  30411=>"101011000",
  30412=>"111111110",
  30413=>"110101101",
  30414=>"101101101",
  30415=>"001010100",
  30416=>"101011110",
  30417=>"110111111",
  30418=>"111001011",
  30419=>"000101101",
  30420=>"000100111",
  30421=>"000000010",
  30422=>"111101001",
  30423=>"111000000",
  30424=>"000111010",
  30425=>"111111111",
  30426=>"011111000",
  30427=>"110010011",
  30428=>"101101110",
  30429=>"001011001",
  30430=>"110100000",
  30431=>"001010001",
  30432=>"111101111",
  30433=>"110001000",
  30434=>"111101100",
  30435=>"100000111",
  30436=>"010101000",
  30437=>"001010010",
  30438=>"101000010",
  30439=>"100011100",
  30440=>"000101111",
  30441=>"110010011",
  30442=>"000111000",
  30443=>"011001101",
  30444=>"000110100",
  30445=>"001110001",
  30446=>"100101110",
  30447=>"100101001",
  30448=>"110011000",
  30449=>"001010010",
  30450=>"011000010",
  30451=>"000100001",
  30452=>"000111011",
  30453=>"010111101",
  30454=>"101101001",
  30455=>"110000111",
  30456=>"011101110",
  30457=>"100111011",
  30458=>"001011001",
  30459=>"010000010",
  30460=>"110000110",
  30461=>"100001101",
  30462=>"010011010",
  30463=>"011110111",
  30464=>"011100000",
  30465=>"100011010",
  30466=>"100011001",
  30467=>"100010000",
  30468=>"011010001",
  30469=>"111101010",
  30470=>"001111001",
  30471=>"110000101",
  30472=>"011110011",
  30473=>"100111001",
  30474=>"010101000",
  30475=>"001001101",
  30476=>"101001110",
  30477=>"101011001",
  30478=>"000000111",
  30479=>"101011001",
  30480=>"001011110",
  30481=>"000000000",
  30482=>"000100011",
  30483=>"011110111",
  30484=>"001001000",
  30485=>"111000011",
  30486=>"101011001",
  30487=>"011101111",
  30488=>"010011111",
  30489=>"000011010",
  30490=>"100010110",
  30491=>"001101110",
  30492=>"110000001",
  30493=>"011001100",
  30494=>"010101010",
  30495=>"111011101",
  30496=>"100111010",
  30497=>"110001011",
  30498=>"001001000",
  30499=>"111001100",
  30500=>"010000010",
  30501=>"010000110",
  30502=>"001100011",
  30503=>"101011011",
  30504=>"010110101",
  30505=>"110000100",
  30506=>"000010111",
  30507=>"000010100",
  30508=>"110011000",
  30509=>"111000001",
  30510=>"000010011",
  30511=>"101111111",
  30512=>"001110111",
  30513=>"101010101",
  30514=>"101000001",
  30515=>"011001101",
  30516=>"110001010",
  30517=>"001010011",
  30518=>"011000101",
  30519=>"101010000",
  30520=>"101001101",
  30521=>"000111000",
  30522=>"100000000",
  30523=>"110000110",
  30524=>"111111100",
  30525=>"111100100",
  30526=>"101010101",
  30527=>"111011110",
  30528=>"111000101",
  30529=>"011011001",
  30530=>"000100001",
  30531=>"000111011",
  30532=>"110011001",
  30533=>"001010101",
  30534=>"110010000",
  30535=>"011100100",
  30536=>"110101100",
  30537=>"011000010",
  30538=>"110111111",
  30539=>"011010000",
  30540=>"001110111",
  30541=>"000000010",
  30542=>"001101111",
  30543=>"000000000",
  30544=>"101000100",
  30545=>"110110101",
  30546=>"101000011",
  30547=>"111101110",
  30548=>"001001011",
  30549=>"110101011",
  30550=>"010000001",
  30551=>"100001101",
  30552=>"011101000",
  30553=>"111111001",
  30554=>"101001101",
  30555=>"100111000",
  30556=>"110111111",
  30557=>"111101010",
  30558=>"100010011",
  30559=>"100011010",
  30560=>"101100001",
  30561=>"000011000",
  30562=>"010110010",
  30563=>"011000101",
  30564=>"000111111",
  30565=>"111110001",
  30566=>"011110100",
  30567=>"100101111",
  30568=>"011100100",
  30569=>"000001101",
  30570=>"100000010",
  30571=>"001110001",
  30572=>"001111011",
  30573=>"010111111",
  30574=>"011000011",
  30575=>"110001000",
  30576=>"000111010",
  30577=>"101101011",
  30578=>"111111101",
  30579=>"000111100",
  30580=>"101000001",
  30581=>"111111000",
  30582=>"100110010",
  30583=>"110101101",
  30584=>"101100100",
  30585=>"001001000",
  30586=>"001010110",
  30587=>"011010011",
  30588=>"111000110",
  30589=>"101101100",
  30590=>"001100111",
  30591=>"110110010",
  30592=>"111101011",
  30593=>"011111110",
  30594=>"011010100",
  30595=>"111001001",
  30596=>"110110010",
  30597=>"100110000",
  30598=>"011010001",
  30599=>"101000101",
  30600=>"101001100",
  30601=>"111010110",
  30602=>"001110010",
  30603=>"000000010",
  30604=>"001100011",
  30605=>"101001111",
  30606=>"111000010",
  30607=>"011001100",
  30608=>"000000101",
  30609=>"110111011",
  30610=>"000111010",
  30611=>"011010000",
  30612=>"100110100",
  30613=>"011111000",
  30614=>"100110010",
  30615=>"110100110",
  30616=>"010011111",
  30617=>"000001010",
  30618=>"000101101",
  30619=>"110010100",
  30620=>"001010100",
  30621=>"111101111",
  30622=>"010110010",
  30623=>"010001110",
  30624=>"100101110",
  30625=>"101110001",
  30626=>"100100011",
  30627=>"111000100",
  30628=>"000010011",
  30629=>"000010011",
  30630=>"110011111",
  30631=>"010000010",
  30632=>"111101101",
  30633=>"110000011",
  30634=>"000100010",
  30635=>"110111101",
  30636=>"010110011",
  30637=>"001000001",
  30638=>"000000011",
  30639=>"101101100",
  30640=>"110000000",
  30641=>"110101001",
  30642=>"000011010",
  30643=>"100010010",
  30644=>"000010010",
  30645=>"110000110",
  30646=>"011010111",
  30647=>"100011111",
  30648=>"010010100",
  30649=>"111011000",
  30650=>"010010001",
  30651=>"011111000",
  30652=>"000000011",
  30653=>"011101000",
  30654=>"111001101",
  30655=>"001110101",
  30656=>"101101111",
  30657=>"000010000",
  30658=>"111001111",
  30659=>"010111011",
  30660=>"000100000",
  30661=>"011110011",
  30662=>"110110101",
  30663=>"001000000",
  30664=>"101010101",
  30665=>"001100000",
  30666=>"011001101",
  30667=>"101100011",
  30668=>"110111111",
  30669=>"110101001",
  30670=>"100111110",
  30671=>"100111001",
  30672=>"100110110",
  30673=>"101101101",
  30674=>"111110111",
  30675=>"110000011",
  30676=>"111001110",
  30677=>"000011011",
  30678=>"010011011",
  30679=>"001000101",
  30680=>"110111111",
  30681=>"110000001",
  30682=>"111100000",
  30683=>"011101011",
  30684=>"111101001",
  30685=>"110010111",
  30686=>"000100000",
  30687=>"100101010",
  30688=>"110101101",
  30689=>"101010111",
  30690=>"001101111",
  30691=>"101000011",
  30692=>"011011101",
  30693=>"000010101",
  30694=>"101011101",
  30695=>"001110111",
  30696=>"100000100",
  30697=>"001011101",
  30698=>"001000101",
  30699=>"010101000",
  30700=>"101001010",
  30701=>"001111100",
  30702=>"110000101",
  30703=>"100111111",
  30704=>"001011111",
  30705=>"111101001",
  30706=>"111001101",
  30707=>"110100011",
  30708=>"110001101",
  30709=>"111001000",
  30710=>"000101110",
  30711=>"110011100",
  30712=>"000010111",
  30713=>"011111111",
  30714=>"001110101",
  30715=>"010010000",
  30716=>"010100011",
  30717=>"010101110",
  30718=>"000011101",
  30719=>"001010101",
  30720=>"001100001",
  30721=>"100001010",
  30722=>"001010110",
  30723=>"111011110",
  30724=>"001111010",
  30725=>"101010011",
  30726=>"111111101",
  30727=>"000000000",
  30728=>"000001010",
  30729=>"011101010",
  30730=>"000001111",
  30731=>"100111010",
  30732=>"111001010",
  30733=>"001100111",
  30734=>"011001000",
  30735=>"000000000",
  30736=>"000011011",
  30737=>"101001110",
  30738=>"100001001",
  30739=>"110010000",
  30740=>"101110101",
  30741=>"000100001",
  30742=>"110111011",
  30743=>"000000010",
  30744=>"111011110",
  30745=>"110010010",
  30746=>"010000010",
  30747=>"001110010",
  30748=>"001000100",
  30749=>"010001100",
  30750=>"011101001",
  30751=>"111110000",
  30752=>"101011001",
  30753=>"010001100",
  30754=>"110001001",
  30755=>"001100010",
  30756=>"111101101",
  30757=>"000101110",
  30758=>"010101111",
  30759=>"000110000",
  30760=>"101110100",
  30761=>"010100100",
  30762=>"000100110",
  30763=>"011110111",
  30764=>"001000111",
  30765=>"101011011",
  30766=>"101001000",
  30767=>"011111100",
  30768=>"010111010",
  30769=>"001100110",
  30770=>"000000001",
  30771=>"010110001",
  30772=>"111010010",
  30773=>"000001110",
  30774=>"000000101",
  30775=>"101111100",
  30776=>"110111001",
  30777=>"011101010",
  30778=>"001101101",
  30779=>"111100001",
  30780=>"011001011",
  30781=>"010001010",
  30782=>"110000001",
  30783=>"100111110",
  30784=>"101101011",
  30785=>"011000011",
  30786=>"001011000",
  30787=>"100100101",
  30788=>"110011000",
  30789=>"000010111",
  30790=>"010111010",
  30791=>"001110101",
  30792=>"000111011",
  30793=>"101101111",
  30794=>"100101001",
  30795=>"011001111",
  30796=>"000001001",
  30797=>"111001100",
  30798=>"010100001",
  30799=>"100010000",
  30800=>"111101110",
  30801=>"000111011",
  30802=>"010110000",
  30803=>"011000101",
  30804=>"001011100",
  30805=>"000010111",
  30806=>"000010010",
  30807=>"111100001",
  30808=>"011011001",
  30809=>"010001010",
  30810=>"100000110",
  30811=>"100100000",
  30812=>"110100010",
  30813=>"101000100",
  30814=>"100000011",
  30815=>"111111000",
  30816=>"000100101",
  30817=>"100010100",
  30818=>"010000101",
  30819=>"010001101",
  30820=>"010110000",
  30821=>"010110001",
  30822=>"010100010",
  30823=>"100110110",
  30824=>"010000000",
  30825=>"101011001",
  30826=>"011100000",
  30827=>"101101010",
  30828=>"000001111",
  30829=>"101011010",
  30830=>"100010101",
  30831=>"011001100",
  30832=>"100000010",
  30833=>"101001101",
  30834=>"011111110",
  30835=>"100000001",
  30836=>"111011100",
  30837=>"110010010",
  30838=>"110101010",
  30839=>"010010110",
  30840=>"111110001",
  30841=>"111110111",
  30842=>"001111011",
  30843=>"110000101",
  30844=>"111100011",
  30845=>"010111000",
  30846=>"011010010",
  30847=>"000010000",
  30848=>"100010000",
  30849=>"011001100",
  30850=>"110001100",
  30851=>"001110101",
  30852=>"100000000",
  30853=>"101011000",
  30854=>"001001011",
  30855=>"000000011",
  30856=>"010110110",
  30857=>"111111111",
  30858=>"011110010",
  30859=>"011101010",
  30860=>"110110000",
  30861=>"011100011",
  30862=>"111111101",
  30863=>"001010000",
  30864=>"010100011",
  30865=>"000010111",
  30866=>"000001000",
  30867=>"011001111",
  30868=>"011010011",
  30869=>"011100100",
  30870=>"011011001",
  30871=>"000111111",
  30872=>"101100001",
  30873=>"000101111",
  30874=>"101101000",
  30875=>"010100011",
  30876=>"110000011",
  30877=>"100100010",
  30878=>"100101100",
  30879=>"001101101",
  30880=>"111010101",
  30881=>"100101010",
  30882=>"100011111",
  30883=>"000000011",
  30884=>"001010110",
  30885=>"111110111",
  30886=>"111110100",
  30887=>"001110111",
  30888=>"110000111",
  30889=>"011111001",
  30890=>"100000010",
  30891=>"010001000",
  30892=>"110011110",
  30893=>"001001001",
  30894=>"111110011",
  30895=>"000000000",
  30896=>"010101111",
  30897=>"010101100",
  30898=>"100100111",
  30899=>"010010101",
  30900=>"000111101",
  30901=>"000100010",
  30902=>"000011111",
  30903=>"010010011",
  30904=>"010000000",
  30905=>"110000010",
  30906=>"110001101",
  30907=>"001011010",
  30908=>"101010010",
  30909=>"111100100",
  30910=>"001000010",
  30911=>"100110001",
  30912=>"101110111",
  30913=>"101000011",
  30914=>"110111000",
  30915=>"011001010",
  30916=>"000001011",
  30917=>"010001100",
  30918=>"001111101",
  30919=>"001110001",
  30920=>"110101100",
  30921=>"101011101",
  30922=>"010001001",
  30923=>"101100010",
  30924=>"101011110",
  30925=>"111101110",
  30926=>"100001001",
  30927=>"000100010",
  30928=>"010101100",
  30929=>"010010101",
  30930=>"100011000",
  30931=>"001011011",
  30932=>"011101000",
  30933=>"001011001",
  30934=>"111011100",
  30935=>"001011011",
  30936=>"011101001",
  30937=>"001100000",
  30938=>"000111001",
  30939=>"100100000",
  30940=>"010111101",
  30941=>"000001100",
  30942=>"111011100",
  30943=>"110101100",
  30944=>"010010101",
  30945=>"000110001",
  30946=>"010000010",
  30947=>"111100110",
  30948=>"101011111",
  30949=>"101000110",
  30950=>"100011111",
  30951=>"110110001",
  30952=>"111001111",
  30953=>"001100010",
  30954=>"100101101",
  30955=>"011001101",
  30956=>"000011001",
  30957=>"111000000",
  30958=>"001011111",
  30959=>"010101100",
  30960=>"111111010",
  30961=>"000111110",
  30962=>"010001000",
  30963=>"000010000",
  30964=>"100111000",
  30965=>"100100101",
  30966=>"111010000",
  30967=>"100001010",
  30968=>"111001000",
  30969=>"101000100",
  30970=>"010111111",
  30971=>"010000111",
  30972=>"000000110",
  30973=>"001010001",
  30974=>"101111000",
  30975=>"000011011",
  30976=>"010101001",
  30977=>"110110001",
  30978=>"100011010",
  30979=>"000110010",
  30980=>"101110110",
  30981=>"010011101",
  30982=>"010111111",
  30983=>"110001100",
  30984=>"010011001",
  30985=>"011100001",
  30986=>"110011101",
  30987=>"011100001",
  30988=>"101011010",
  30989=>"010010001",
  30990=>"001111100",
  30991=>"010100110",
  30992=>"101101100",
  30993=>"111111110",
  30994=>"001110111",
  30995=>"101111000",
  30996=>"000000010",
  30997=>"011010111",
  30998=>"000001110",
  30999=>"100000110",
  31000=>"110010100",
  31001=>"011010110",
  31002=>"110110111",
  31003=>"010100001",
  31004=>"000010110",
  31005=>"011111110",
  31006=>"010101010",
  31007=>"001001011",
  31008=>"000001111",
  31009=>"011100101",
  31010=>"101111011",
  31011=>"000111001",
  31012=>"011111110",
  31013=>"000101110",
  31014=>"001011010",
  31015=>"011110111",
  31016=>"100011110",
  31017=>"000111010",
  31018=>"111001110",
  31019=>"101110010",
  31020=>"011001011",
  31021=>"100110011",
  31022=>"101100111",
  31023=>"000011111",
  31024=>"101011111",
  31025=>"100011111",
  31026=>"001010001",
  31027=>"000011001",
  31028=>"100110010",
  31029=>"000100100",
  31030=>"110000110",
  31031=>"010111000",
  31032=>"101101111",
  31033=>"111001001",
  31034=>"100101001",
  31035=>"111000010",
  31036=>"001101100",
  31037=>"011000001",
  31038=>"001100101",
  31039=>"000110101",
  31040=>"000001000",
  31041=>"110001001",
  31042=>"010111010",
  31043=>"001001110",
  31044=>"001110000",
  31045=>"001000001",
  31046=>"100010001",
  31047=>"011010110",
  31048=>"010100001",
  31049=>"100100000",
  31050=>"011011110",
  31051=>"011001001",
  31052=>"111110110",
  31053=>"011100000",
  31054=>"010000000",
  31055=>"011110111",
  31056=>"111110110",
  31057=>"001111110",
  31058=>"101000001",
  31059=>"111000000",
  31060=>"100000010",
  31061=>"100001101",
  31062=>"011101010",
  31063=>"100001001",
  31064=>"101000000",
  31065=>"001101111",
  31066=>"001101101",
  31067=>"011000000",
  31068=>"011111011",
  31069=>"001111111",
  31070=>"000011011",
  31071=>"000011110",
  31072=>"100101000",
  31073=>"011000011",
  31074=>"011101100",
  31075=>"100001011",
  31076=>"101110111",
  31077=>"100100000",
  31078=>"101011111",
  31079=>"101001000",
  31080=>"100101011",
  31081=>"010110010",
  31082=>"100100010",
  31083=>"000001111",
  31084=>"001000110",
  31085=>"011110000",
  31086=>"000110000",
  31087=>"101111011",
  31088=>"011111111",
  31089=>"110101110",
  31090=>"011110000",
  31091=>"101110101",
  31092=>"010011000",
  31093=>"101011000",
  31094=>"000101111",
  31095=>"000010111",
  31096=>"110110111",
  31097=>"101000110",
  31098=>"101110100",
  31099=>"111111110",
  31100=>"010000110",
  31101=>"000001010",
  31102=>"100100111",
  31103=>"011100101",
  31104=>"000101101",
  31105=>"011010100",
  31106=>"110111011",
  31107=>"101000000",
  31108=>"111101010",
  31109=>"000101001",
  31110=>"000001000",
  31111=>"011110000",
  31112=>"010000110",
  31113=>"101110110",
  31114=>"110110001",
  31115=>"110011000",
  31116=>"010001110",
  31117=>"110101001",
  31118=>"001000000",
  31119=>"010000101",
  31120=>"101001011",
  31121=>"000101110",
  31122=>"101000001",
  31123=>"100000000",
  31124=>"110001110",
  31125=>"101111100",
  31126=>"000111101",
  31127=>"000100000",
  31128=>"110001001",
  31129=>"000011010",
  31130=>"000001011",
  31131=>"000101110",
  31132=>"010011111",
  31133=>"000111001",
  31134=>"111110011",
  31135=>"011111100",
  31136=>"100001001",
  31137=>"001100100",
  31138=>"111000010",
  31139=>"101001101",
  31140=>"011111010",
  31141=>"000100011",
  31142=>"110111010",
  31143=>"001111110",
  31144=>"000101011",
  31145=>"010100111",
  31146=>"001110111",
  31147=>"111111001",
  31148=>"100011100",
  31149=>"110100100",
  31150=>"110000100",
  31151=>"011000110",
  31152=>"101100101",
  31153=>"010100101",
  31154=>"011100100",
  31155=>"101100000",
  31156=>"011010101",
  31157=>"011111110",
  31158=>"001101100",
  31159=>"100010000",
  31160=>"101100000",
  31161=>"011000000",
  31162=>"100011110",
  31163=>"000000001",
  31164=>"110011000",
  31165=>"111001111",
  31166=>"001110110",
  31167=>"000000011",
  31168=>"010000001",
  31169=>"100000110",
  31170=>"111010110",
  31171=>"100100010",
  31172=>"011110000",
  31173=>"010010101",
  31174=>"101111010",
  31175=>"001000001",
  31176=>"000100000",
  31177=>"101001000",
  31178=>"111110011",
  31179=>"000101010",
  31180=>"100101011",
  31181=>"111110101",
  31182=>"101000001",
  31183=>"000110011",
  31184=>"111011100",
  31185=>"011010010",
  31186=>"000011111",
  31187=>"110110010",
  31188=>"110000101",
  31189=>"100011000",
  31190=>"010110111",
  31191=>"110010110",
  31192=>"011000111",
  31193=>"001001110",
  31194=>"111111111",
  31195=>"101000111",
  31196=>"101111101",
  31197=>"011110111",
  31198=>"011110111",
  31199=>"111111000",
  31200=>"111010000",
  31201=>"010000111",
  31202=>"101100010",
  31203=>"010110000",
  31204=>"101011111",
  31205=>"000000100",
  31206=>"010110001",
  31207=>"110100111",
  31208=>"001110111",
  31209=>"010101111",
  31210=>"101100111",
  31211=>"000001100",
  31212=>"000001000",
  31213=>"011010010",
  31214=>"100110111",
  31215=>"101111010",
  31216=>"010010101",
  31217=>"111001010",
  31218=>"011000111",
  31219=>"100000001",
  31220=>"000011010",
  31221=>"001100110",
  31222=>"111101101",
  31223=>"110100010",
  31224=>"001000010",
  31225=>"100011101",
  31226=>"000000010",
  31227=>"000001001",
  31228=>"010101100",
  31229=>"011101000",
  31230=>"000110010",
  31231=>"111000110",
  31232=>"010110011",
  31233=>"001000011",
  31234=>"000110010",
  31235=>"000000101",
  31236=>"001111110",
  31237=>"100010101",
  31238=>"101010110",
  31239=>"010010010",
  31240=>"000010101",
  31241=>"000000011",
  31242=>"111100110",
  31243=>"010010000",
  31244=>"101100111",
  31245=>"110111000",
  31246=>"110010000",
  31247=>"110001101",
  31248=>"001111000",
  31249=>"000001101",
  31250=>"010001010",
  31251=>"011011111",
  31252=>"011010111",
  31253=>"011001000",
  31254=>"011100000",
  31255=>"001110100",
  31256=>"100111111",
  31257=>"100000110",
  31258=>"010001110",
  31259=>"010010001",
  31260=>"001000000",
  31261=>"000001100",
  31262=>"110111000",
  31263=>"010011010",
  31264=>"000010101",
  31265=>"101111111",
  31266=>"001100111",
  31267=>"101100010",
  31268=>"101011111",
  31269=>"101011100",
  31270=>"000010010",
  31271=>"010101001",
  31272=>"100110010",
  31273=>"011011111",
  31274=>"100101111",
  31275=>"100010000",
  31276=>"010010100",
  31277=>"100010111",
  31278=>"010000000",
  31279=>"001001110",
  31280=>"101111101",
  31281=>"110001100",
  31282=>"011011000",
  31283=>"111010010",
  31284=>"000100000",
  31285=>"001111010",
  31286=>"010010011",
  31287=>"100001100",
  31288=>"111011100",
  31289=>"011011100",
  31290=>"110100110",
  31291=>"101111001",
  31292=>"011110100",
  31293=>"000001110",
  31294=>"111001101",
  31295=>"111101101",
  31296=>"111110010",
  31297=>"101011100",
  31298=>"101000011",
  31299=>"100001101",
  31300=>"100000100",
  31301=>"100111101",
  31302=>"001011000",
  31303=>"100111111",
  31304=>"110100000",
  31305=>"010010010",
  31306=>"101110010",
  31307=>"100100101",
  31308=>"010010110",
  31309=>"101001111",
  31310=>"101111010",
  31311=>"100110101",
  31312=>"111010100",
  31313=>"100111111",
  31314=>"010111100",
  31315=>"111111011",
  31316=>"111011111",
  31317=>"100001011",
  31318=>"001001011",
  31319=>"001111010",
  31320=>"101100100",
  31321=>"110010101",
  31322=>"111011100",
  31323=>"000101111",
  31324=>"101101111",
  31325=>"010100000",
  31326=>"101001000",
  31327=>"101000010",
  31328=>"011001000",
  31329=>"111111111",
  31330=>"100011001",
  31331=>"101101111",
  31332=>"111110001",
  31333=>"000000100",
  31334=>"110111110",
  31335=>"001001010",
  31336=>"000000001",
  31337=>"110100011",
  31338=>"100011101",
  31339=>"100101001",
  31340=>"100111110",
  31341=>"101011000",
  31342=>"010110001",
  31343=>"110100110",
  31344=>"100100111",
  31345=>"000001000",
  31346=>"111101111",
  31347=>"010010110",
  31348=>"101111111",
  31349=>"100001011",
  31350=>"111001011",
  31351=>"000011000",
  31352=>"100111111",
  31353=>"001011001",
  31354=>"100111111",
  31355=>"110011100",
  31356=>"010000001",
  31357=>"100001100",
  31358=>"101011000",
  31359=>"111001011",
  31360=>"010011000",
  31361=>"100110010",
  31362=>"001100000",
  31363=>"110110110",
  31364=>"110100100",
  31365=>"010000000",
  31366=>"101010101",
  31367=>"100110001",
  31368=>"100100110",
  31369=>"000100100",
  31370=>"100110010",
  31371=>"110101101",
  31372=>"111001001",
  31373=>"000000100",
  31374=>"111101110",
  31375=>"100001001",
  31376=>"110100011",
  31377=>"101110100",
  31378=>"101110011",
  31379=>"001111011",
  31380=>"000010010",
  31381=>"010110111",
  31382=>"011111111",
  31383=>"010101111",
  31384=>"001011000",
  31385=>"011001111",
  31386=>"100000010",
  31387=>"110111110",
  31388=>"010110110",
  31389=>"010100111",
  31390=>"110010101",
  31391=>"101100010",
  31392=>"101100011",
  31393=>"111001110",
  31394=>"011001110",
  31395=>"001010010",
  31396=>"111100001",
  31397=>"101000011",
  31398=>"001011010",
  31399=>"000000110",
  31400=>"111111010",
  31401=>"110011101",
  31402=>"001000101",
  31403=>"000000000",
  31404=>"010010011",
  31405=>"010101010",
  31406=>"010111001",
  31407=>"100011010",
  31408=>"000001111",
  31409=>"100111001",
  31410=>"111000100",
  31411=>"110101011",
  31412=>"110111010",
  31413=>"011110101",
  31414=>"110011100",
  31415=>"001100100",
  31416=>"010110011",
  31417=>"001101111",
  31418=>"101100001",
  31419=>"110101101",
  31420=>"101100110",
  31421=>"111000110",
  31422=>"011001010",
  31423=>"010110100",
  31424=>"110101110",
  31425=>"110010011",
  31426=>"100100000",
  31427=>"010000001",
  31428=>"101010000",
  31429=>"100100000",
  31430=>"001110010",
  31431=>"101101011",
  31432=>"010110110",
  31433=>"100011110",
  31434=>"000110111",
  31435=>"100110111",
  31436=>"100000010",
  31437=>"111011011",
  31438=>"111001011",
  31439=>"000011111",
  31440=>"100100110",
  31441=>"111000000",
  31442=>"011100000",
  31443=>"000101011",
  31444=>"010000011",
  31445=>"110111111",
  31446=>"100011011",
  31447=>"011000100",
  31448=>"001000110",
  31449=>"010010110",
  31450=>"011100010",
  31451=>"011101111",
  31452=>"011000111",
  31453=>"000010001",
  31454=>"111000000",
  31455=>"101011100",
  31456=>"011100111",
  31457=>"110000101",
  31458=>"011100111",
  31459=>"000110110",
  31460=>"101101010",
  31461=>"101010000",
  31462=>"100111111",
  31463=>"100001001",
  31464=>"100101110",
  31465=>"111000011",
  31466=>"011101000",
  31467=>"101001100",
  31468=>"011011011",
  31469=>"000001111",
  31470=>"110011110",
  31471=>"110111000",
  31472=>"000111011",
  31473=>"110110000",
  31474=>"111001000",
  31475=>"100011010",
  31476=>"000100010",
  31477=>"110111110",
  31478=>"001110110",
  31479=>"110110010",
  31480=>"010010011",
  31481=>"011101011",
  31482=>"111101110",
  31483=>"101001011",
  31484=>"000011001",
  31485=>"011100010",
  31486=>"010101111",
  31487=>"011001000",
  31488=>"011011011",
  31489=>"001000100",
  31490=>"100011111",
  31491=>"100011101",
  31492=>"101001000",
  31493=>"100000010",
  31494=>"101100100",
  31495=>"101111000",
  31496=>"100110010",
  31497=>"111010001",
  31498=>"000110001",
  31499=>"101000111",
  31500=>"000000001",
  31501=>"110010101",
  31502=>"100101011",
  31503=>"101011110",
  31504=>"001110001",
  31505=>"010011000",
  31506=>"111001111",
  31507=>"100001100",
  31508=>"101000100",
  31509=>"010010010",
  31510=>"011110011",
  31511=>"101110101",
  31512=>"011001110",
  31513=>"011011010",
  31514=>"011001101",
  31515=>"111001010",
  31516=>"111111101",
  31517=>"000001001",
  31518=>"000111101",
  31519=>"100001110",
  31520=>"100111101",
  31521=>"100110110",
  31522=>"110011111",
  31523=>"010101011",
  31524=>"101100011",
  31525=>"001010110",
  31526=>"001110000",
  31527=>"010101000",
  31528=>"000010001",
  31529=>"111100100",
  31530=>"101010001",
  31531=>"111100111",
  31532=>"011011011",
  31533=>"101110111",
  31534=>"111000000",
  31535=>"001001010",
  31536=>"110000011",
  31537=>"011101111",
  31538=>"010000001",
  31539=>"000101101",
  31540=>"001011010",
  31541=>"111110110",
  31542=>"101100110",
  31543=>"001010101",
  31544=>"101110101",
  31545=>"101000010",
  31546=>"001010011",
  31547=>"000010010",
  31548=>"001011001",
  31549=>"000101111",
  31550=>"100101010",
  31551=>"110000110",
  31552=>"111101001",
  31553=>"010011100",
  31554=>"110000000",
  31555=>"001111000",
  31556=>"110010001",
  31557=>"100010010",
  31558=>"001101001",
  31559=>"010001111",
  31560=>"111011111",
  31561=>"110001010",
  31562=>"100111000",
  31563=>"010100001",
  31564=>"111011111",
  31565=>"010011111",
  31566=>"111101000",
  31567=>"010000101",
  31568=>"001001111",
  31569=>"100000011",
  31570=>"100000111",
  31571=>"010111101",
  31572=>"011010100",
  31573=>"100100011",
  31574=>"101000110",
  31575=>"000000100",
  31576=>"000001010",
  31577=>"000011100",
  31578=>"011100100",
  31579=>"101101011",
  31580=>"111010110",
  31581=>"010011001",
  31582=>"001110011",
  31583=>"100100110",
  31584=>"100001001",
  31585=>"111100111",
  31586=>"110011010",
  31587=>"000000101",
  31588=>"111111101",
  31589=>"010111011",
  31590=>"010001011",
  31591=>"000110110",
  31592=>"111011010",
  31593=>"010010000",
  31594=>"110101001",
  31595=>"110110110",
  31596=>"101111101",
  31597=>"101001111",
  31598=>"001011110",
  31599=>"000011100",
  31600=>"101001010",
  31601=>"100110000",
  31602=>"011000101",
  31603=>"000110001",
  31604=>"001011101",
  31605=>"111111101",
  31606=>"110110100",
  31607=>"000011100",
  31608=>"111100101",
  31609=>"111111100",
  31610=>"111000000",
  31611=>"000101010",
  31612=>"000000010",
  31613=>"100000100",
  31614=>"111100000",
  31615=>"110001111",
  31616=>"010111111",
  31617=>"100001100",
  31618=>"001000000",
  31619=>"001111010",
  31620=>"111100110",
  31621=>"111111011",
  31622=>"001101000",
  31623=>"100101100",
  31624=>"111010101",
  31625=>"010001010",
  31626=>"100101100",
  31627=>"111110101",
  31628=>"100010101",
  31629=>"001000110",
  31630=>"011101010",
  31631=>"001011110",
  31632=>"000111001",
  31633=>"011100000",
  31634=>"000101000",
  31635=>"101000111",
  31636=>"100110101",
  31637=>"100011101",
  31638=>"010001011",
  31639=>"101110101",
  31640=>"110000110",
  31641=>"010000110",
  31642=>"101111000",
  31643=>"001001011",
  31644=>"001101000",
  31645=>"011110111",
  31646=>"000010010",
  31647=>"111110100",
  31648=>"001110000",
  31649=>"111000100",
  31650=>"110011001",
  31651=>"111000110",
  31652=>"001111001",
  31653=>"110110111",
  31654=>"101111010",
  31655=>"010100010",
  31656=>"100010001",
  31657=>"100001111",
  31658=>"010110110",
  31659=>"011011101",
  31660=>"110011101",
  31661=>"111001110",
  31662=>"111110011",
  31663=>"000111100",
  31664=>"101010000",
  31665=>"110011111",
  31666=>"010010000",
  31667=>"100001111",
  31668=>"011111010",
  31669=>"111011011",
  31670=>"111110001",
  31671=>"101001000",
  31672=>"000110111",
  31673=>"001111111",
  31674=>"010101011",
  31675=>"100010100",
  31676=>"100110111",
  31677=>"000101000",
  31678=>"110101110",
  31679=>"011001111",
  31680=>"101100001",
  31681=>"111101100",
  31682=>"001001110",
  31683=>"001100101",
  31684=>"001100101",
  31685=>"101000001",
  31686=>"000011010",
  31687=>"000100100",
  31688=>"001100010",
  31689=>"101001110",
  31690=>"010000101",
  31691=>"101000010",
  31692=>"010110011",
  31693=>"000010001",
  31694=>"010010000",
  31695=>"000011010",
  31696=>"000001111",
  31697=>"011101001",
  31698=>"011010100",
  31699=>"101110100",
  31700=>"000001100",
  31701=>"100010011",
  31702=>"110011011",
  31703=>"000100001",
  31704=>"001010111",
  31705=>"001001101",
  31706=>"011010010",
  31707=>"100001011",
  31708=>"001111011",
  31709=>"100011111",
  31710=>"101011010",
  31711=>"111000001",
  31712=>"100111000",
  31713=>"111111010",
  31714=>"000000100",
  31715=>"100000110",
  31716=>"000110011",
  31717=>"011101100",
  31718=>"000010100",
  31719=>"100010001",
  31720=>"010000010",
  31721=>"111011011",
  31722=>"101000100",
  31723=>"000110100",
  31724=>"000000000",
  31725=>"000000101",
  31726=>"100101000",
  31727=>"101000110",
  31728=>"101100010",
  31729=>"101101110",
  31730=>"001010000",
  31731=>"011100100",
  31732=>"110011101",
  31733=>"111001111",
  31734=>"101001000",
  31735=>"011000111",
  31736=>"000001100",
  31737=>"101101100",
  31738=>"011011011",
  31739=>"100111100",
  31740=>"001010010",
  31741=>"001110000",
  31742=>"100011101",
  31743=>"011111011",
  31744=>"000100001",
  31745=>"111110000",
  31746=>"010000011",
  31747=>"110000010",
  31748=>"101101110",
  31749=>"100100010",
  31750=>"110010001",
  31751=>"000001111",
  31752=>"101101111",
  31753=>"001001010",
  31754=>"111010110",
  31755=>"010000100",
  31756=>"100111000",
  31757=>"101010110",
  31758=>"011111101",
  31759=>"011100011",
  31760=>"110110000",
  31761=>"000001011",
  31762=>"101111111",
  31763=>"100101001",
  31764=>"011011001",
  31765=>"001100001",
  31766=>"010010111",
  31767=>"110000111",
  31768=>"000000001",
  31769=>"001010110",
  31770=>"010101001",
  31771=>"001011001",
  31772=>"111010000",
  31773=>"110011010",
  31774=>"111101001",
  31775=>"101010001",
  31776=>"101011011",
  31777=>"011010010",
  31778=>"110001000",
  31779=>"011011011",
  31780=>"111011101",
  31781=>"101001111",
  31782=>"001101010",
  31783=>"010101001",
  31784=>"100010001",
  31785=>"000110110",
  31786=>"011100111",
  31787=>"100100110",
  31788=>"111111011",
  31789=>"101111111",
  31790=>"100001101",
  31791=>"100111011",
  31792=>"010011110",
  31793=>"001111000",
  31794=>"110000001",
  31795=>"111011100",
  31796=>"111100101",
  31797=>"100101000",
  31798=>"111010010",
  31799=>"110000000",
  31800=>"000001011",
  31801=>"100010111",
  31802=>"000010100",
  31803=>"111010110",
  31804=>"001001000",
  31805=>"001101011",
  31806=>"000101000",
  31807=>"100000100",
  31808=>"011011010",
  31809=>"000101011",
  31810=>"111001010",
  31811=>"101010001",
  31812=>"000000000",
  31813=>"000001001",
  31814=>"011100011",
  31815=>"011000001",
  31816=>"001010000",
  31817=>"010001111",
  31818=>"100110100",
  31819=>"111001011",
  31820=>"001000110",
  31821=>"100000101",
  31822=>"110011000",
  31823=>"000111010",
  31824=>"011110110",
  31825=>"101101101",
  31826=>"110110111",
  31827=>"001101010",
  31828=>"110111001",
  31829=>"101110111",
  31830=>"101111110",
  31831=>"010101100",
  31832=>"110111000",
  31833=>"000011101",
  31834=>"100010000",
  31835=>"111111010",
  31836=>"111000100",
  31837=>"101100101",
  31838=>"000100101",
  31839=>"001001111",
  31840=>"110010100",
  31841=>"101000001",
  31842=>"011011010",
  31843=>"000100101",
  31844=>"101110000",
  31845=>"101010110",
  31846=>"101100000",
  31847=>"011111111",
  31848=>"000100010",
  31849=>"001010011",
  31850=>"011110111",
  31851=>"011011000",
  31852=>"111101111",
  31853=>"010101101",
  31854=>"111111000",
  31855=>"011001101",
  31856=>"101001011",
  31857=>"101000110",
  31858=>"111110100",
  31859=>"111011111",
  31860=>"101111001",
  31861=>"100110000",
  31862=>"000110011",
  31863=>"101100010",
  31864=>"100111010",
  31865=>"010101110",
  31866=>"101100010",
  31867=>"010111010",
  31868=>"110101010",
  31869=>"000010000",
  31870=>"110100001",
  31871=>"101000001",
  31872=>"000011111",
  31873=>"111000010",
  31874=>"000011111",
  31875=>"001001010",
  31876=>"101101001",
  31877=>"011001100",
  31878=>"001111101",
  31879=>"001001010",
  31880=>"001010100",
  31881=>"010101000",
  31882=>"001001101",
  31883=>"111101000",
  31884=>"111000101",
  31885=>"111011110",
  31886=>"011001101",
  31887=>"111010010",
  31888=>"011111110",
  31889=>"110101100",
  31890=>"011001101",
  31891=>"101111101",
  31892=>"111000101",
  31893=>"011101110",
  31894=>"001101000",
  31895=>"110101110",
  31896=>"100000111",
  31897=>"000011001",
  31898=>"110111110",
  31899=>"101101000",
  31900=>"100011010",
  31901=>"001000000",
  31902=>"000100001",
  31903=>"101100100",
  31904=>"000110011",
  31905=>"100001101",
  31906=>"000000000",
  31907=>"100011000",
  31908=>"011010011",
  31909=>"101100101",
  31910=>"011000101",
  31911=>"001000100",
  31912=>"101000011",
  31913=>"101101111",
  31914=>"111010001",
  31915=>"111100110",
  31916=>"110110101",
  31917=>"110101111",
  31918=>"010111100",
  31919=>"101111010",
  31920=>"101011111",
  31921=>"101001011",
  31922=>"001111111",
  31923=>"000111011",
  31924=>"110100000",
  31925=>"010000000",
  31926=>"010000010",
  31927=>"100011001",
  31928=>"110110010",
  31929=>"111100000",
  31930=>"110100100",
  31931=>"101010111",
  31932=>"011101011",
  31933=>"000101001",
  31934=>"101110100",
  31935=>"000011010",
  31936=>"011000001",
  31937=>"001110110",
  31938=>"100000010",
  31939=>"101011111",
  31940=>"010101100",
  31941=>"110111001",
  31942=>"101100001",
  31943=>"000000010",
  31944=>"101001001",
  31945=>"101101111",
  31946=>"010110011",
  31947=>"100001100",
  31948=>"000000101",
  31949=>"011010111",
  31950=>"101110111",
  31951=>"111100101",
  31952=>"010100100",
  31953=>"111111110",
  31954=>"100001111",
  31955=>"111000101",
  31956=>"011011000",
  31957=>"110011010",
  31958=>"010111101",
  31959=>"011100001",
  31960=>"001000010",
  31961=>"001100100",
  31962=>"110010000",
  31963=>"101100011",
  31964=>"100110110",
  31965=>"000000100",
  31966=>"111001111",
  31967=>"111011001",
  31968=>"100011101",
  31969=>"100111110",
  31970=>"011001110",
  31971=>"001011110",
  31972=>"000000101",
  31973=>"011101100",
  31974=>"010000001",
  31975=>"101000111",
  31976=>"101011111",
  31977=>"101011010",
  31978=>"010010000",
  31979=>"011100110",
  31980=>"111110111",
  31981=>"001011100",
  31982=>"101100000",
  31983=>"100000010",
  31984=>"111010111",
  31985=>"011000001",
  31986=>"010111111",
  31987=>"101111111",
  31988=>"110110111",
  31989=>"101111010",
  31990=>"100100011",
  31991=>"011110000",
  31992=>"001001100",
  31993=>"000110111",
  31994=>"111100011",
  31995=>"111101111",
  31996=>"100010000",
  31997=>"111001101",
  31998=>"001110001",
  31999=>"001001001",
  32000=>"011010011",
  32001=>"111110010",
  32002=>"101000111",
  32003=>"111001111",
  32004=>"010110101",
  32005=>"011001010",
  32006=>"001100111",
  32007=>"000100001",
  32008=>"010011001",
  32009=>"100010111",
  32010=>"010000001",
  32011=>"000010000",
  32012=>"100101001",
  32013=>"001110111",
  32014=>"011100000",
  32015=>"111101011",
  32016=>"000100101",
  32017=>"101000011",
  32018=>"001010111",
  32019=>"001101000",
  32020=>"010011101",
  32021=>"000101011",
  32022=>"101001100",
  32023=>"101110011",
  32024=>"111010111",
  32025=>"100010000",
  32026=>"011001100",
  32027=>"000110101",
  32028=>"001111111",
  32029=>"000100011",
  32030=>"011111011",
  32031=>"011011101",
  32032=>"001100001",
  32033=>"011000110",
  32034=>"100000001",
  32035=>"000101000",
  32036=>"101010000",
  32037=>"100000010",
  32038=>"011001110",
  32039=>"001111001",
  32040=>"001100000",
  32041=>"001111011",
  32042=>"010100110",
  32043=>"100011011",
  32044=>"010111000",
  32045=>"110101011",
  32046=>"111111001",
  32047=>"100111101",
  32048=>"001101101",
  32049=>"100011000",
  32050=>"100001000",
  32051=>"001110100",
  32052=>"000010100",
  32053=>"000001100",
  32054=>"100010101",
  32055=>"100010111",
  32056=>"000010101",
  32057=>"010010111",
  32058=>"010110001",
  32059=>"111101111",
  32060=>"111111110",
  32061=>"000110011",
  32062=>"011001011",
  32063=>"000000011",
  32064=>"000000111",
  32065=>"110001010",
  32066=>"111101111",
  32067=>"111010101",
  32068=>"000110100",
  32069=>"111001001",
  32070=>"010000111",
  32071=>"000110000",
  32072=>"001000001",
  32073=>"000100001",
  32074=>"000001101",
  32075=>"001110000",
  32076=>"111011111",
  32077=>"110000110",
  32078=>"101001011",
  32079=>"011001100",
  32080=>"111101111",
  32081=>"111101100",
  32082=>"101101111",
  32083=>"000001010",
  32084=>"100100010",
  32085=>"011110100",
  32086=>"011010001",
  32087=>"010100100",
  32088=>"011100010",
  32089=>"111110100",
  32090=>"001110100",
  32091=>"111010111",
  32092=>"011010100",
  32093=>"001101101",
  32094=>"111111000",
  32095=>"111011000",
  32096=>"001101000",
  32097=>"100010011",
  32098=>"100001011",
  32099=>"100010111",
  32100=>"111010010",
  32101=>"101110111",
  32102=>"110010110",
  32103=>"111110010",
  32104=>"100110101",
  32105=>"100000010",
  32106=>"101001010",
  32107=>"100100101",
  32108=>"011110011",
  32109=>"100101111",
  32110=>"001010110",
  32111=>"111110011",
  32112=>"111001110",
  32113=>"010111111",
  32114=>"001100001",
  32115=>"010010100",
  32116=>"110101010",
  32117=>"010111000",
  32118=>"010001100",
  32119=>"001001101",
  32120=>"000110111",
  32121=>"111101111",
  32122=>"110011001",
  32123=>"111000011",
  32124=>"000000111",
  32125=>"011010011",
  32126=>"101111101",
  32127=>"100101001",
  32128=>"000001000",
  32129=>"010011010",
  32130=>"100001000",
  32131=>"110101110",
  32132=>"100000110",
  32133=>"011000100",
  32134=>"111110000",
  32135=>"100110001",
  32136=>"110000100",
  32137=>"001101010",
  32138=>"000110010",
  32139=>"000000100",
  32140=>"101001010",
  32141=>"010100011",
  32142=>"011001100",
  32143=>"001001101",
  32144=>"011001001",
  32145=>"100110000",
  32146=>"011010100",
  32147=>"111100011",
  32148=>"101000111",
  32149=>"011000010",
  32150=>"011110011",
  32151=>"101111111",
  32152=>"100001011",
  32153=>"100000011",
  32154=>"100010100",
  32155=>"111010101",
  32156=>"101001101",
  32157=>"011101111",
  32158=>"010101111",
  32159=>"101001001",
  32160=>"101101110",
  32161=>"011001111",
  32162=>"001100010",
  32163=>"011110100",
  32164=>"011000001",
  32165=>"000111110",
  32166=>"000100101",
  32167=>"101111111",
  32168=>"000101000",
  32169=>"000100101",
  32170=>"011001000",
  32171=>"100100101",
  32172=>"010100011",
  32173=>"001110001",
  32174=>"010000000",
  32175=>"111111101",
  32176=>"000100000",
  32177=>"010011000",
  32178=>"000110001",
  32179=>"111101011",
  32180=>"100011111",
  32181=>"101100100",
  32182=>"100101101",
  32183=>"011001110",
  32184=>"100011010",
  32185=>"000000101",
  32186=>"010101110",
  32187=>"001001111",
  32188=>"000000010",
  32189=>"111111101",
  32190=>"110110101",
  32191=>"101001000",
  32192=>"000110001",
  32193=>"111010100",
  32194=>"000110000",
  32195=>"000110111",
  32196=>"101010000",
  32197=>"101100010",
  32198=>"100000000",
  32199=>"001101001",
  32200=>"000000000",
  32201=>"000001001",
  32202=>"110110011",
  32203=>"111010001",
  32204=>"111111000",
  32205=>"000100000",
  32206=>"010001011",
  32207=>"011000110",
  32208=>"000001000",
  32209=>"010111100",
  32210=>"101011011",
  32211=>"010000101",
  32212=>"010111111",
  32213=>"111100101",
  32214=>"000011001",
  32215=>"010000010",
  32216=>"101100000",
  32217=>"111011011",
  32218=>"001001110",
  32219=>"110100000",
  32220=>"111100001",
  32221=>"000011011",
  32222=>"100000000",
  32223=>"011010100",
  32224=>"001010010",
  32225=>"010011011",
  32226=>"110011110",
  32227=>"000110011",
  32228=>"001000001",
  32229=>"111101100",
  32230=>"101000001",
  32231=>"111001101",
  32232=>"010011101",
  32233=>"100110101",
  32234=>"101011100",
  32235=>"000000100",
  32236=>"000000000",
  32237=>"110001010",
  32238=>"010000100",
  32239=>"001101011",
  32240=>"001011110",
  32241=>"101000110",
  32242=>"101011000",
  32243=>"010100101",
  32244=>"101000000",
  32245=>"111100110",
  32246=>"101001010",
  32247=>"011001011",
  32248=>"010101100",
  32249=>"010110110",
  32250=>"010101000",
  32251=>"011111111",
  32252=>"101101111",
  32253=>"001001111",
  32254=>"100101101",
  32255=>"110110101",
  32256=>"100010010",
  32257=>"111000010",
  32258=>"000000111",
  32259=>"010101000",
  32260=>"101111000",
  32261=>"011110010",
  32262=>"000001111",
  32263=>"010110000",
  32264=>"111100000",
  32265=>"101001001",
  32266=>"111101110",
  32267=>"010011010",
  32268=>"101001101",
  32269=>"000010100",
  32270=>"000111101",
  32271=>"100010010",
  32272=>"011100001",
  32273=>"001110101",
  32274=>"100011110",
  32275=>"010111011",
  32276=>"010000001",
  32277=>"001011111",
  32278=>"001000011",
  32279=>"010000000",
  32280=>"101011010",
  32281=>"001101111",
  32282=>"000100001",
  32283=>"001011000",
  32284=>"100001000",
  32285=>"010010111",
  32286=>"111000111",
  32287=>"111100010",
  32288=>"011110110",
  32289=>"000010010",
  32290=>"001000000",
  32291=>"001000101",
  32292=>"000100110",
  32293=>"100101010",
  32294=>"110000010",
  32295=>"010000100",
  32296=>"000111111",
  32297=>"101111101",
  32298=>"001010100",
  32299=>"101110100",
  32300=>"101011001",
  32301=>"101111011",
  32302=>"001010101",
  32303=>"000010001",
  32304=>"100001010",
  32305=>"010111110",
  32306=>"100000100",
  32307=>"100111001",
  32308=>"110110100",
  32309=>"010110001",
  32310=>"001110111",
  32311=>"010001100",
  32312=>"011001101",
  32313=>"000110100",
  32314=>"101110000",
  32315=>"001100111",
  32316=>"111111111",
  32317=>"111110111",
  32318=>"110000011",
  32319=>"010000011",
  32320=>"000100010",
  32321=>"100000110",
  32322=>"010101010",
  32323=>"001101101",
  32324=>"001010001",
  32325=>"001001011",
  32326=>"001001100",
  32327=>"100111110",
  32328=>"011101010",
  32329=>"100100010",
  32330=>"100100000",
  32331=>"101001100",
  32332=>"111101110",
  32333=>"101010011",
  32334=>"100000001",
  32335=>"000011110",
  32336=>"100000100",
  32337=>"000000001",
  32338=>"100110110",
  32339=>"001100100",
  32340=>"000001110",
  32341=>"111110011",
  32342=>"111100100",
  32343=>"011010101",
  32344=>"111111000",
  32345=>"001011110",
  32346=>"010011101",
  32347=>"101010000",
  32348=>"010001011",
  32349=>"110010010",
  32350=>"011011101",
  32351=>"000000100",
  32352=>"101001100",
  32353=>"010111011",
  32354=>"011101011",
  32355=>"010101001",
  32356=>"100100111",
  32357=>"111011100",
  32358=>"111110001",
  32359=>"011101010",
  32360=>"010000010",
  32361=>"101110110",
  32362=>"000100000",
  32363=>"000011100",
  32364=>"001100001",
  32365=>"111111011",
  32366=>"011100110",
  32367=>"110110101",
  32368=>"100110011",
  32369=>"010000010",
  32370=>"101110110",
  32371=>"000101000",
  32372=>"001001110",
  32373=>"101010011",
  32374=>"010001010",
  32375=>"010100010",
  32376=>"010000010",
  32377=>"011101011",
  32378=>"000000010",
  32379=>"001111000",
  32380=>"001001000",
  32381=>"011111101",
  32382=>"100011110",
  32383=>"010001010",
  32384=>"001010100",
  32385=>"000101000",
  32386=>"110001011",
  32387=>"010001100",
  32388=>"010001101",
  32389=>"000100000",
  32390=>"111101001",
  32391=>"000111111",
  32392=>"111100001",
  32393=>"000000010",
  32394=>"011001001",
  32395=>"001101001",
  32396=>"100111110",
  32397=>"000010110",
  32398=>"010111000",
  32399=>"100100101",
  32400=>"011101100",
  32401=>"101111000",
  32402=>"010000000",
  32403=>"110110000",
  32404=>"111100100",
  32405=>"010111000",
  32406=>"010110010",
  32407=>"111100110",
  32408=>"100111001",
  32409=>"011111010",
  32410=>"001110010",
  32411=>"100101101",
  32412=>"110001011",
  32413=>"011000000",
  32414=>"010101010",
  32415=>"010100110",
  32416=>"111111110",
  32417=>"010000111",
  32418=>"001000110",
  32419=>"100010110",
  32420=>"111111101",
  32421=>"101101111",
  32422=>"001000101",
  32423=>"101110111",
  32424=>"000110111",
  32425=>"000011011",
  32426=>"011000111",
  32427=>"100111100",
  32428=>"000110011",
  32429=>"111110100",
  32430=>"111101010",
  32431=>"111010010",
  32432=>"000000010",
  32433=>"110111010",
  32434=>"110000011",
  32435=>"001000010",
  32436=>"110101010",
  32437=>"001100111",
  32438=>"111101100",
  32439=>"111010111",
  32440=>"011111101",
  32441=>"100100010",
  32442=>"110111011",
  32443=>"100011101",
  32444=>"010010010",
  32445=>"100011010",
  32446=>"011101100",
  32447=>"100000000",
  32448=>"111000111",
  32449=>"001000001",
  32450=>"110010111",
  32451=>"101110101",
  32452=>"100000101",
  32453=>"100100101",
  32454=>"000110011",
  32455=>"111110111",
  32456=>"001000000",
  32457=>"010000000",
  32458=>"010000010",
  32459=>"010101101",
  32460=>"111111111",
  32461=>"000000100",
  32462=>"110010110",
  32463=>"011011010",
  32464=>"011110111",
  32465=>"100001111",
  32466=>"000010110",
  32467=>"011111011",
  32468=>"000101001",
  32469=>"111011110",
  32470=>"110000011",
  32471=>"001011010",
  32472=>"010011011",
  32473=>"110111001",
  32474=>"000111110",
  32475=>"111110011",
  32476=>"000110110",
  32477=>"110111000",
  32478=>"100011100",
  32479=>"001010100",
  32480=>"000001111",
  32481=>"001001101",
  32482=>"000100100",
  32483=>"100001101",
  32484=>"111110100",
  32485=>"101111110",
  32486=>"011101010",
  32487=>"110100101",
  32488=>"010011100",
  32489=>"110111001",
  32490=>"001000011",
  32491=>"010010111",
  32492=>"001111110",
  32493=>"111111001",
  32494=>"011100001",
  32495=>"000010000",
  32496=>"101110001",
  32497=>"011111111",
  32498=>"111110001",
  32499=>"100110011",
  32500=>"010001110",
  32501=>"101100101",
  32502=>"011001111",
  32503=>"110100110",
  32504=>"000111101",
  32505=>"010111001",
  32506=>"000000011",
  32507=>"000101101",
  32508=>"111101101",
  32509=>"011111111",
  32510=>"000110010",
  32511=>"110100010",
  32512=>"101111101",
  32513=>"111110011",
  32514=>"011010001",
  32515=>"110100001",
  32516=>"011010000",
  32517=>"111011111",
  32518=>"000111010",
  32519=>"000110110",
  32520=>"010101100",
  32521=>"001000001",
  32522=>"001011100",
  32523=>"000000000",
  32524=>"010100001",
  32525=>"001100011",
  32526=>"010110111",
  32527=>"101010000",
  32528=>"111100111",
  32529=>"100010001",
  32530=>"101001111",
  32531=>"011100001",
  32532=>"110011110",
  32533=>"001110110",
  32534=>"011010101",
  32535=>"010111001",
  32536=>"101001001",
  32537=>"011100000",
  32538=>"111000100",
  32539=>"110000011",
  32540=>"101100111",
  32541=>"101101010",
  32542=>"110001100",
  32543=>"110011101",
  32544=>"010101001",
  32545=>"011110010",
  32546=>"001101011",
  32547=>"001010110",
  32548=>"111111010",
  32549=>"010101111",
  32550=>"110011100",
  32551=>"001011100",
  32552=>"101011010",
  32553=>"000001101",
  32554=>"111100100",
  32555=>"011111111",
  32556=>"000110101",
  32557=>"111101001",
  32558=>"010000110",
  32559=>"110100111",
  32560=>"011101111",
  32561=>"001000011",
  32562=>"001010000",
  32563=>"100011010",
  32564=>"101000001",
  32565=>"111101001",
  32566=>"110111010",
  32567=>"111001010",
  32568=>"100110000",
  32569=>"011101000",
  32570=>"000000001",
  32571=>"111111001",
  32572=>"010111010",
  32573=>"110000010",
  32574=>"010100101",
  32575=>"010101111",
  32576=>"100100100",
  32577=>"001011110",
  32578=>"100100100",
  32579=>"110010100",
  32580=>"101001011",
  32581=>"100101001",
  32582=>"111111011",
  32583=>"011100011",
  32584=>"111110010",
  32585=>"000010011",
  32586=>"011100101",
  32587=>"100110011",
  32588=>"011101000",
  32589=>"100010010",
  32590=>"001001101",
  32591=>"110111010",
  32592=>"100011001",
  32593=>"000111010",
  32594=>"000000010",
  32595=>"010110111",
  32596=>"110001111",
  32597=>"110111101",
  32598=>"000100111",
  32599=>"111110000",
  32600=>"110000110",
  32601=>"110011100",
  32602=>"110110011",
  32603=>"001101101",
  32604=>"010101000",
  32605=>"101000000",
  32606=>"111111100",
  32607=>"011101111",
  32608=>"110011000",
  32609=>"000100000",
  32610=>"111100000",
  32611=>"100000100",
  32612=>"010101111",
  32613=>"010100000",
  32614=>"101000010",
  32615=>"101111111",
  32616=>"111010111",
  32617=>"111110110",
  32618=>"001110000",
  32619=>"111110010",
  32620=>"001111110",
  32621=>"101101110",
  32622=>"100100111",
  32623=>"111001111",
  32624=>"000111010",
  32625=>"000100000",
  32626=>"000110110",
  32627=>"111100010",
  32628=>"000010111",
  32629=>"100000110",
  32630=>"011001100",
  32631=>"000000000",
  32632=>"000010101",
  32633=>"111101100",
  32634=>"010111110",
  32635=>"101111001",
  32636=>"100111010",
  32637=>"000100011",
  32638=>"111011111",
  32639=>"100010100",
  32640=>"110000100",
  32641=>"000001001",
  32642=>"000010100",
  32643=>"100010110",
  32644=>"100011101",
  32645=>"000010110",
  32646=>"000100100",
  32647=>"110010100",
  32648=>"010001000",
  32649=>"011001110",
  32650=>"010010100",
  32651=>"111001101",
  32652=>"000110100",
  32653=>"110101011",
  32654=>"001101111",
  32655=>"101110111",
  32656=>"000001000",
  32657=>"001100101",
  32658=>"110000001",
  32659=>"000000001",
  32660=>"011110010",
  32661=>"100000000",
  32662=>"010000111",
  32663=>"010101110",
  32664=>"110001111",
  32665=>"100101001",
  32666=>"110111111",
  32667=>"000101011",
  32668=>"100101111",
  32669=>"110111011",
  32670=>"010001100",
  32671=>"101100111",
  32672=>"111110100",
  32673=>"100100010",
  32674=>"110100111",
  32675=>"100000111",
  32676=>"000000111",
  32677=>"110111100",
  32678=>"001111010",
  32679=>"101100000",
  32680=>"010000000",
  32681=>"001011001",
  32682=>"101010111",
  32683=>"011101000",
  32684=>"001010001",
  32685=>"011110110",
  32686=>"110011011",
  32687=>"000100010",
  32688=>"101101000",
  32689=>"000110100",
  32690=>"101100100",
  32691=>"111100100",
  32692=>"101111001",
  32693=>"001110011",
  32694=>"110101100",
  32695=>"110110001",
  32696=>"000011001",
  32697=>"000001011",
  32698=>"001001100",
  32699=>"010011001",
  32700=>"101011110",
  32701=>"001101111",
  32702=>"010011001",
  32703=>"111110011",
  32704=>"101100000",
  32705=>"000011010",
  32706=>"011111110",
  32707=>"000110111",
  32708=>"000100001",
  32709=>"111011101",
  32710=>"010000100",
  32711=>"011000000",
  32712=>"111000001",
  32713=>"100001000",
  32714=>"111001111",
  32715=>"111010001",
  32716=>"100010101",
  32717=>"011001110",
  32718=>"011011010",
  32719=>"010000000",
  32720=>"101100001",
  32721=>"100111110",
  32722=>"000110000",
  32723=>"101101010",
  32724=>"101111110",
  32725=>"001010111",
  32726=>"111010011",
  32727=>"010001001",
  32728=>"110111111",
  32729=>"100100101",
  32730=>"101101111",
  32731=>"100001010",
  32732=>"110111101",
  32733=>"100000011",
  32734=>"011111010",
  32735=>"100001011",
  32736=>"110111110",
  32737=>"001101101",
  32738=>"001011011",
  32739=>"001000011",
  32740=>"110011010",
  32741=>"000010000",
  32742=>"011001011",
  32743=>"011011111",
  32744=>"110111011",
  32745=>"100010101",
  32746=>"000000011",
  32747=>"100010111",
  32748=>"111010011",
  32749=>"001010001",
  32750=>"100001100",
  32751=>"001111011",
  32752=>"010011011",
  32753=>"001011001",
  32754=>"111001000",
  32755=>"101000100",
  32756=>"110000100",
  32757=>"111110010",
  32758=>"111110110",
  32759=>"001000011",
  32760=>"100000001",
  32761=>"000111001",
  32762=>"010000011",
  32763=>"100100011",
  32764=>"111001110",
  32765=>"111010100",
  32766=>"110001101",
  32767=>"011000000",
  32768=>"101000100",
  32769=>"110011100",
  32770=>"000101011",
  32771=>"110100110",
  32772=>"000001110",
  32773=>"000011101",
  32774=>"010001100",
  32775=>"101000011",
  32776=>"000111010",
  32777=>"101010101",
  32778=>"110111110",
  32779=>"110111111",
  32780=>"000101110",
  32781=>"001000111",
  32782=>"011010010",
  32783=>"110000010",
  32784=>"110010000",
  32785=>"111110101",
  32786=>"001000000",
  32787=>"010111111",
  32788=>"001000110",
  32789=>"111001110",
  32790=>"011101101",
  32791=>"000000000",
  32792=>"000101101",
  32793=>"101101111",
  32794=>"100010110",
  32795=>"011100000",
  32796=>"111101001",
  32797=>"110100100",
  32798=>"000000001",
  32799=>"001010001",
  32800=>"111011111",
  32801=>"000011101",
  32802=>"101101000",
  32803=>"100010101",
  32804=>"010111001",
  32805=>"001011110",
  32806=>"001010101",
  32807=>"110101101",
  32808=>"001110000",
  32809=>"001011101",
  32810=>"101101011",
  32811=>"001110110",
  32812=>"000110011",
  32813=>"001110110",
  32814=>"010010010",
  32815=>"110111100",
  32816=>"100110011",
  32817=>"001110101",
  32818=>"001110101",
  32819=>"001110111",
  32820=>"100101011",
  32821=>"111100010",
  32822=>"011010000",
  32823=>"010010011",
  32824=>"011111101",
  32825=>"100001010",
  32826=>"010101110",
  32827=>"111111111",
  32828=>"001000101",
  32829=>"111011001",
  32830=>"111111100",
  32831=>"001000001",
  32832=>"000010110",
  32833=>"001000000",
  32834=>"011001000",
  32835=>"100001110",
  32836=>"001110011",
  32837=>"101001011",
  32838=>"000010110",
  32839=>"110000111",
  32840=>"100011001",
  32841=>"011001001",
  32842=>"011100100",
  32843=>"000010000",
  32844=>"100110000",
  32845=>"001110001",
  32846=>"001110111",
  32847=>"010111001",
  32848=>"011010001",
  32849=>"100110001",
  32850=>"111111110",
  32851=>"110001000",
  32852=>"101010000",
  32853=>"010110111",
  32854=>"001000001",
  32855=>"110000001",
  32856=>"000011110",
  32857=>"111110000",
  32858=>"111000101",
  32859=>"000100000",
  32860=>"110011111",
  32861=>"100000101",
  32862=>"001110001",
  32863=>"001001110",
  32864=>"001000000",
  32865=>"101001010",
  32866=>"110111000",
  32867=>"000100110",
  32868=>"100111000",
  32869=>"101000010",
  32870=>"001010001",
  32871=>"110111100",
  32872=>"011100110",
  32873=>"000101000",
  32874=>"110010111",
  32875=>"001000001",
  32876=>"000000100",
  32877=>"011101011",
  32878=>"000101100",
  32879=>"101000111",
  32880=>"011101011",
  32881=>"111001101",
  32882=>"010111001",
  32883=>"011100110",
  32884=>"000010110",
  32885=>"101001110",
  32886=>"010000000",
  32887=>"011100111",
  32888=>"001101110",
  32889=>"111001001",
  32890=>"001011000",
  32891=>"011100001",
  32892=>"011010010",
  32893=>"101110101",
  32894=>"000001000",
  32895=>"010000101",
  32896=>"100011001",
  32897=>"101011101",
  32898=>"001000100",
  32899=>"100110010",
  32900=>"101000011",
  32901=>"100111101",
  32902=>"001000111",
  32903=>"001111001",
  32904=>"010010001",
  32905=>"100101001",
  32906=>"011001011",
  32907=>"100111110",
  32908=>"100101111",
  32909=>"100001100",
  32910=>"101001001",
  32911=>"100100010",
  32912=>"111100111",
  32913=>"111100111",
  32914=>"010110110",
  32915=>"000100100",
  32916=>"010011110",
  32917=>"111011100",
  32918=>"100010000",
  32919=>"010110110",
  32920=>"110110110",
  32921=>"010111011",
  32922=>"001011000",
  32923=>"010000001",
  32924=>"111100000",
  32925=>"001110011",
  32926=>"100001011",
  32927=>"100101010",
  32928=>"100101101",
  32929=>"111110111",
  32930=>"000011101",
  32931=>"011101001",
  32932=>"000111100",
  32933=>"001010101",
  32934=>"010000111",
  32935=>"000001010",
  32936=>"000010000",
  32937=>"010001101",
  32938=>"111001111",
  32939=>"011110100",
  32940=>"000010110",
  32941=>"000010101",
  32942=>"100110010",
  32943=>"000111001",
  32944=>"011001101",
  32945=>"000110010",
  32946=>"001110001",
  32947=>"000101011",
  32948=>"110110111",
  32949=>"001010101",
  32950=>"101110111",
  32951=>"111110100",
  32952=>"001101111",
  32953=>"111011000",
  32954=>"101001011",
  32955=>"110111011",
  32956=>"110001010",
  32957=>"100011001",
  32958=>"010110101",
  32959=>"011110011",
  32960=>"100010000",
  32961=>"001011101",
  32962=>"110111000",
  32963=>"111101111",
  32964=>"110101010",
  32965=>"000001100",
  32966=>"001010010",
  32967=>"110101101",
  32968=>"000000111",
  32969=>"101000100",
  32970=>"001101101",
  32971=>"010001110",
  32972=>"111101001",
  32973=>"100110101",
  32974=>"011001101",
  32975=>"011111010",
  32976=>"110111100",
  32977=>"111010010",
  32978=>"100010110",
  32979=>"110011111",
  32980=>"000110010",
  32981=>"110011001",
  32982=>"110111111",
  32983=>"101010110",
  32984=>"011011100",
  32985=>"001101110",
  32986=>"000000000",
  32987=>"001001000",
  32988=>"001100111",
  32989=>"011000000",
  32990=>"110011110",
  32991=>"010110111",
  32992=>"100000110",
  32993=>"001110011",
  32994=>"010001001",
  32995=>"010101001",
  32996=>"011101101",
  32997=>"111100101",
  32998=>"100010100",
  32999=>"011000111",
  33000=>"111010000",
  33001=>"110111000",
  33002=>"011101111",
  33003=>"110000110",
  33004=>"011000000",
  33005=>"010000001",
  33006=>"000001010",
  33007=>"111011110",
  33008=>"000000010",
  33009=>"010001000",
  33010=>"001001010",
  33011=>"011010110",
  33012=>"101011111",
  33013=>"111100100",
  33014=>"010011010",
  33015=>"010110111",
  33016=>"001111011",
  33017=>"001010100",
  33018=>"001101110",
  33019=>"101101011",
  33020=>"110011111",
  33021=>"000010011",
  33022=>"111110101",
  33023=>"000011111",
  33024=>"110111101",
  33025=>"001000001",
  33026=>"011010011",
  33027=>"111011101",
  33028=>"011000000",
  33029=>"001110111",
  33030=>"111000001",
  33031=>"010111010",
  33032=>"101101110",
  33033=>"001100011",
  33034=>"101111101",
  33035=>"000000100",
  33036=>"100101011",
  33037=>"111000011",
  33038=>"001100111",
  33039=>"001101100",
  33040=>"010000011",
  33041=>"001110100",
  33042=>"110111011",
  33043=>"000110101",
  33044=>"101111011",
  33045=>"000011000",
  33046=>"101110000",
  33047=>"000001000",
  33048=>"111001101",
  33049=>"000000010",
  33050=>"100100010",
  33051=>"001000010",
  33052=>"000110100",
  33053=>"010100001",
  33054=>"111011101",
  33055=>"000101101",
  33056=>"000111010",
  33057=>"101110111",
  33058=>"011000101",
  33059=>"111110110",
  33060=>"011000111",
  33061=>"001000001",
  33062=>"001111101",
  33063=>"010011100",
  33064=>"100100001",
  33065=>"000110111",
  33066=>"011110010",
  33067=>"001001001",
  33068=>"110011001",
  33069=>"000000100",
  33070=>"010101100",
  33071=>"000011111",
  33072=>"100111010",
  33073=>"001101101",
  33074=>"111111110",
  33075=>"100000111",
  33076=>"111110100",
  33077=>"101010100",
  33078=>"001011000",
  33079=>"001001101",
  33080=>"010011001",
  33081=>"010101000",
  33082=>"011000010",
  33083=>"101111100",
  33084=>"000000000",
  33085=>"001000011",
  33086=>"110011100",
  33087=>"001011100",
  33088=>"110011001",
  33089=>"110010111",
  33090=>"000110010",
  33091=>"100110011",
  33092=>"010011110",
  33093=>"101110100",
  33094=>"101000011",
  33095=>"101111000",
  33096=>"100001110",
  33097=>"101000010",
  33098=>"000010111",
  33099=>"011100010",
  33100=>"111000110",
  33101=>"100000000",
  33102=>"001111110",
  33103=>"111001110",
  33104=>"100000101",
  33105=>"100110110",
  33106=>"000000001",
  33107=>"000001110",
  33108=>"000110010",
  33109=>"101111110",
  33110=>"101101000",
  33111=>"010010110",
  33112=>"001010100",
  33113=>"110010010",
  33114=>"010000100",
  33115=>"100101110",
  33116=>"100001011",
  33117=>"110111100",
  33118=>"011101000",
  33119=>"001000101",
  33120=>"110000011",
  33121=>"010101010",
  33122=>"111100000",
  33123=>"101001111",
  33124=>"111100110",
  33125=>"110010110",
  33126=>"100001111",
  33127=>"100000001",
  33128=>"100010110",
  33129=>"111010110",
  33130=>"001101110",
  33131=>"000000110",
  33132=>"000001000",
  33133=>"010001101",
  33134=>"110101000",
  33135=>"000100100",
  33136=>"001110110",
  33137=>"111000011",
  33138=>"001111110",
  33139=>"111010111",
  33140=>"011111000",
  33141=>"001011000",
  33142=>"000001100",
  33143=>"000101011",
  33144=>"001000010",
  33145=>"011001000",
  33146=>"001101100",
  33147=>"100000101",
  33148=>"000010110",
  33149=>"110111110",
  33150=>"011111111",
  33151=>"110011000",
  33152=>"100111011",
  33153=>"000010000",
  33154=>"011111101",
  33155=>"111111001",
  33156=>"111100110",
  33157=>"010010000",
  33158=>"111100011",
  33159=>"001001011",
  33160=>"000001100",
  33161=>"011111111",
  33162=>"001001101",
  33163=>"110011000",
  33164=>"011110101",
  33165=>"000000000",
  33166=>"000111011",
  33167=>"110111100",
  33168=>"111000101",
  33169=>"010000000",
  33170=>"100001000",
  33171=>"010010011",
  33172=>"010100000",
  33173=>"000001111",
  33174=>"100001110",
  33175=>"010110110",
  33176=>"011101111",
  33177=>"101100100",
  33178=>"010111000",
  33179=>"010110000",
  33180=>"111111000",
  33181=>"100110100",
  33182=>"001100110",
  33183=>"011111101",
  33184=>"100110011",
  33185=>"101001000",
  33186=>"010100011",
  33187=>"011000101",
  33188=>"000100101",
  33189=>"111111001",
  33190=>"011000100",
  33191=>"111001100",
  33192=>"110011001",
  33193=>"100110011",
  33194=>"011111001",
  33195=>"111111101",
  33196=>"100101010",
  33197=>"110011010",
  33198=>"111001010",
  33199=>"110111111",
  33200=>"111110110",
  33201=>"100000010",
  33202=>"100011111",
  33203=>"000010010",
  33204=>"110101010",
  33205=>"110110010",
  33206=>"001110010",
  33207=>"001111111",
  33208=>"101110111",
  33209=>"010010110",
  33210=>"100101001",
  33211=>"000110110",
  33212=>"111110010",
  33213=>"110110111",
  33214=>"001100000",
  33215=>"111110000",
  33216=>"110001000",
  33217=>"100010111",
  33218=>"110100011",
  33219=>"000011010",
  33220=>"000010010",
  33221=>"001101000",
  33222=>"110110101",
  33223=>"111000111",
  33224=>"111100101",
  33225=>"010100101",
  33226=>"111110111",
  33227=>"010110111",
  33228=>"101010100",
  33229=>"100010000",
  33230=>"101001000",
  33231=>"111000111",
  33232=>"000000000",
  33233=>"111010010",
  33234=>"100100001",
  33235=>"100101111",
  33236=>"001111111",
  33237=>"101000110",
  33238=>"101101111",
  33239=>"101010000",
  33240=>"010001010",
  33241=>"111100011",
  33242=>"110101011",
  33243=>"001111000",
  33244=>"001010010",
  33245=>"110010101",
  33246=>"011001101",
  33247=>"100101101",
  33248=>"100010100",
  33249=>"010100100",
  33250=>"101011101",
  33251=>"100011101",
  33252=>"001000000",
  33253=>"101011011",
  33254=>"010001010",
  33255=>"111001110",
  33256=>"100010110",
  33257=>"101011111",
  33258=>"010000000",
  33259=>"011001011",
  33260=>"111100111",
  33261=>"000000111",
  33262=>"101001101",
  33263=>"110101100",
  33264=>"101001000",
  33265=>"101111100",
  33266=>"100010011",
  33267=>"011001010",
  33268=>"101011011",
  33269=>"001001001",
  33270=>"110011100",
  33271=>"101000101",
  33272=>"000000110",
  33273=>"100010000",
  33274=>"010010010",
  33275=>"111011110",
  33276=>"111010110",
  33277=>"100100011",
  33278=>"001110001",
  33279=>"011000110",
  33280=>"000100100",
  33281=>"100111011",
  33282=>"101101011",
  33283=>"000000010",
  33284=>"111000101",
  33285=>"001101011",
  33286=>"011100110",
  33287=>"100011001",
  33288=>"011001011",
  33289=>"000100111",
  33290=>"010110110",
  33291=>"000100100",
  33292=>"010110010",
  33293=>"000101110",
  33294=>"000110010",
  33295=>"100001111",
  33296=>"110000111",
  33297=>"111000100",
  33298=>"000110100",
  33299=>"111010110",
  33300=>"000000110",
  33301=>"011110101",
  33302=>"000000000",
  33303=>"001111010",
  33304=>"000111110",
  33305=>"100110110",
  33306=>"010000000",
  33307=>"101010010",
  33308=>"001110111",
  33309=>"001000011",
  33310=>"001010100",
  33311=>"011111111",
  33312=>"101101011",
  33313=>"000000000",
  33314=>"101110101",
  33315=>"000010111",
  33316=>"011100011",
  33317=>"100001101",
  33318=>"110100010",
  33319=>"101010011",
  33320=>"111100011",
  33321=>"001101000",
  33322=>"101110101",
  33323=>"010100111",
  33324=>"010111010",
  33325=>"010000000",
  33326=>"010111010",
  33327=>"111011101",
  33328=>"011001001",
  33329=>"100000000",
  33330=>"010001010",
  33331=>"001000100",
  33332=>"010011010",
  33333=>"101100101",
  33334=>"000110011",
  33335=>"001101010",
  33336=>"101111100",
  33337=>"100101000",
  33338=>"110011011",
  33339=>"010110000",
  33340=>"111101000",
  33341=>"000010000",
  33342=>"100001100",
  33343=>"001110110",
  33344=>"000111000",
  33345=>"011011111",
  33346=>"011000110",
  33347=>"110010100",
  33348=>"000010101",
  33349=>"011011011",
  33350=>"011000110",
  33351=>"110111000",
  33352=>"011001010",
  33353=>"111101111",
  33354=>"011001010",
  33355=>"001111111",
  33356=>"100000001",
  33357=>"111110110",
  33358=>"000010101",
  33359=>"000001110",
  33360=>"110111011",
  33361=>"001100011",
  33362=>"001010001",
  33363=>"011010001",
  33364=>"000011111",
  33365=>"010001011",
  33366=>"111110010",
  33367=>"101110100",
  33368=>"111001010",
  33369=>"001011010",
  33370=>"110101110",
  33371=>"111110111",
  33372=>"100100110",
  33373=>"010000010",
  33374=>"100010110",
  33375=>"001000011",
  33376=>"000010001",
  33377=>"010010010",
  33378=>"010111101",
  33379=>"111101110",
  33380=>"000000001",
  33381=>"110010111",
  33382=>"001000110",
  33383=>"100010000",
  33384=>"011000100",
  33385=>"110101001",
  33386=>"100010010",
  33387=>"101001011",
  33388=>"101011101",
  33389=>"000100011",
  33390=>"101101010",
  33391=>"111011000",
  33392=>"101101100",
  33393=>"001100110",
  33394=>"011011101",
  33395=>"101001110",
  33396=>"011111111",
  33397=>"111011000",
  33398=>"100111110",
  33399=>"010101011",
  33400=>"001011111",
  33401=>"111010101",
  33402=>"111101111",
  33403=>"101101001",
  33404=>"000110100",
  33405=>"111110101",
  33406=>"000001110",
  33407=>"101101011",
  33408=>"110011010",
  33409=>"101010101",
  33410=>"000011100",
  33411=>"100100111",
  33412=>"011000111",
  33413=>"001111001",
  33414=>"100010111",
  33415=>"111101110",
  33416=>"001000001",
  33417=>"100110100",
  33418=>"111111111",
  33419=>"101010111",
  33420=>"010111111",
  33421=>"010010011",
  33422=>"000001100",
  33423=>"001001001",
  33424=>"000100000",
  33425=>"000101001",
  33426=>"100100100",
  33427=>"001011111",
  33428=>"100011001",
  33429=>"010100110",
  33430=>"001110011",
  33431=>"111100000",
  33432=>"101100100",
  33433=>"001000011",
  33434=>"011010001",
  33435=>"000010110",
  33436=>"100000110",
  33437=>"011100000",
  33438=>"111011000",
  33439=>"101101000",
  33440=>"101001101",
  33441=>"100101000",
  33442=>"011001101",
  33443=>"000110010",
  33444=>"001001000",
  33445=>"111100011",
  33446=>"000000011",
  33447=>"001000110",
  33448=>"110111001",
  33449=>"010110111",
  33450=>"101110011",
  33451=>"101110100",
  33452=>"000000000",
  33453=>"110000011",
  33454=>"001011101",
  33455=>"110101111",
  33456=>"111111001",
  33457=>"001011110",
  33458=>"000000001",
  33459=>"111111110",
  33460=>"110111100",
  33461=>"010001100",
  33462=>"001000111",
  33463=>"101000001",
  33464=>"001011111",
  33465=>"100011111",
  33466=>"101100001",
  33467=>"010010001",
  33468=>"111111111",
  33469=>"100100000",
  33470=>"000000011",
  33471=>"111111010",
  33472=>"001111100",
  33473=>"111011101",
  33474=>"110110001",
  33475=>"101001110",
  33476=>"100110011",
  33477=>"111001100",
  33478=>"100000011",
  33479=>"011100101",
  33480=>"011100000",
  33481=>"010010100",
  33482=>"000101010",
  33483=>"000010010",
  33484=>"101111000",
  33485=>"010101101",
  33486=>"100100001",
  33487=>"000110111",
  33488=>"011001110",
  33489=>"000000101",
  33490=>"110100100",
  33491=>"000101101",
  33492=>"111100000",
  33493=>"001010001",
  33494=>"000101100",
  33495=>"100000010",
  33496=>"111111001",
  33497=>"110110001",
  33498=>"110100010",
  33499=>"010100011",
  33500=>"000000001",
  33501=>"100101110",
  33502=>"101000011",
  33503=>"011001101",
  33504=>"011000010",
  33505=>"000000011",
  33506=>"100010010",
  33507=>"011111101",
  33508=>"111111001",
  33509=>"101011100",
  33510=>"001111101",
  33511=>"111110100",
  33512=>"010000111",
  33513=>"111110111",
  33514=>"001101110",
  33515=>"010010000",
  33516=>"000100100",
  33517=>"001101100",
  33518=>"100001011",
  33519=>"000001000",
  33520=>"010110011",
  33521=>"000011011",
  33522=>"001110011",
  33523=>"000010110",
  33524=>"010101011",
  33525=>"100101000",
  33526=>"001001110",
  33527=>"111011101",
  33528=>"100000111",
  33529=>"011100010",
  33530=>"101011110",
  33531=>"001000110",
  33532=>"000110010",
  33533=>"110111110",
  33534=>"111111000",
  33535=>"000010111",
  33536=>"100000101",
  33537=>"000011101",
  33538=>"111111011",
  33539=>"000000011",
  33540=>"000010001",
  33541=>"000111101",
  33542=>"010100001",
  33543=>"111100100",
  33544=>"110110010",
  33545=>"111111011",
  33546=>"010011101",
  33547=>"010011111",
  33548=>"110001001",
  33549=>"001010011",
  33550=>"110110110",
  33551=>"001000101",
  33552=>"100111110",
  33553=>"010010001",
  33554=>"111100110",
  33555=>"001011000",
  33556=>"101011100",
  33557=>"101101101",
  33558=>"110001000",
  33559=>"100001110",
  33560=>"101011110",
  33561=>"001001001",
  33562=>"001100110",
  33563=>"010010111",
  33564=>"110100101",
  33565=>"000001100",
  33566=>"011101110",
  33567=>"100110010",
  33568=>"100111111",
  33569=>"011010010",
  33570=>"000000100",
  33571=>"111000000",
  33572=>"011001111",
  33573=>"000001001",
  33574=>"000000001",
  33575=>"110111100",
  33576=>"100010111",
  33577=>"010001011",
  33578=>"100110100",
  33579=>"100011001",
  33580=>"011101111",
  33581=>"000000001",
  33582=>"000101001",
  33583=>"101111000",
  33584=>"101101010",
  33585=>"001110000",
  33586=>"101001010",
  33587=>"101110111",
  33588=>"111001000",
  33589=>"111100110",
  33590=>"010000100",
  33591=>"001101011",
  33592=>"100001101",
  33593=>"010100100",
  33594=>"000111111",
  33595=>"110011101",
  33596=>"011000100",
  33597=>"110101111",
  33598=>"111001111",
  33599=>"100111001",
  33600=>"110011001",
  33601=>"100010001",
  33602=>"010111001",
  33603=>"111011010",
  33604=>"101100010",
  33605=>"110001110",
  33606=>"100110001",
  33607=>"011111100",
  33608=>"110101100",
  33609=>"101101011",
  33610=>"001000110",
  33611=>"000011011",
  33612=>"110101011",
  33613=>"010010111",
  33614=>"111111111",
  33615=>"101010100",
  33616=>"011101000",
  33617=>"100011111",
  33618=>"000010100",
  33619=>"110010010",
  33620=>"101000000",
  33621=>"001110000",
  33622=>"000100101",
  33623=>"001000100",
  33624=>"001011011",
  33625=>"110000010",
  33626=>"011110000",
  33627=>"010100010",
  33628=>"001011001",
  33629=>"011100110",
  33630=>"101011001",
  33631=>"010010010",
  33632=>"000000100",
  33633=>"000100001",
  33634=>"011101001",
  33635=>"111111110",
  33636=>"010001001",
  33637=>"101000101",
  33638=>"101000010",
  33639=>"100100101",
  33640=>"000010000",
  33641=>"100111101",
  33642=>"101000001",
  33643=>"011010000",
  33644=>"011011011",
  33645=>"101110000",
  33646=>"100111110",
  33647=>"111011100",
  33648=>"100000000",
  33649=>"000001111",
  33650=>"101001011",
  33651=>"111001010",
  33652=>"000101110",
  33653=>"001000111",
  33654=>"010011000",
  33655=>"011011110",
  33656=>"000010011",
  33657=>"100010100",
  33658=>"000001001",
  33659=>"100111000",
  33660=>"000100001",
  33661=>"111100010",
  33662=>"101111100",
  33663=>"011110110",
  33664=>"111100100",
  33665=>"100010101",
  33666=>"100001111",
  33667=>"000001100",
  33668=>"101010100",
  33669=>"101110001",
  33670=>"001101001",
  33671=>"000110100",
  33672=>"100000110",
  33673=>"000100111",
  33674=>"101101101",
  33675=>"000000100",
  33676=>"010010011",
  33677=>"111010101",
  33678=>"111100101",
  33679=>"001110110",
  33680=>"111011110",
  33681=>"001101010",
  33682=>"110111011",
  33683=>"011110001",
  33684=>"010001110",
  33685=>"101110011",
  33686=>"001100010",
  33687=>"100111100",
  33688=>"111111111",
  33689=>"011111011",
  33690=>"000100111",
  33691=>"110111111",
  33692=>"100000100",
  33693=>"001000010",
  33694=>"001110010",
  33695=>"011001110",
  33696=>"010001010",
  33697=>"011001011",
  33698=>"100111000",
  33699=>"000000010",
  33700=>"001110101",
  33701=>"111111111",
  33702=>"101000111",
  33703=>"110000011",
  33704=>"110100010",
  33705=>"010100111",
  33706=>"110101110",
  33707=>"001101011",
  33708=>"111110100",
  33709=>"011110101",
  33710=>"100101101",
  33711=>"000011111",
  33712=>"001001001",
  33713=>"110110111",
  33714=>"001011111",
  33715=>"100000011",
  33716=>"011111010",
  33717=>"111100011",
  33718=>"111010101",
  33719=>"011110111",
  33720=>"011001000",
  33721=>"001011000",
  33722=>"000101101",
  33723=>"010001010",
  33724=>"000011001",
  33725=>"100010010",
  33726=>"111101110",
  33727=>"100001100",
  33728=>"000101110",
  33729=>"001110111",
  33730=>"000000000",
  33731=>"100001100",
  33732=>"000101111",
  33733=>"110011101",
  33734=>"110111111",
  33735=>"001011101",
  33736=>"101000000",
  33737=>"100111100",
  33738=>"001100101",
  33739=>"000000010",
  33740=>"100010010",
  33741=>"001011011",
  33742=>"111100101",
  33743=>"000110110",
  33744=>"001000110",
  33745=>"101110001",
  33746=>"000000110",
  33747=>"011011100",
  33748=>"010000000",
  33749=>"101011001",
  33750=>"001100000",
  33751=>"100100111",
  33752=>"011000111",
  33753=>"000010110",
  33754=>"001010001",
  33755=>"000100111",
  33756=>"111110110",
  33757=>"101011011",
  33758=>"010100011",
  33759=>"111110001",
  33760=>"111110001",
  33761=>"000000010",
  33762=>"100111000",
  33763=>"101001110",
  33764=>"100001111",
  33765=>"111011110",
  33766=>"000110110",
  33767=>"010001111",
  33768=>"010000101",
  33769=>"101101100",
  33770=>"010001000",
  33771=>"011011001",
  33772=>"110010110",
  33773=>"000100100",
  33774=>"111111100",
  33775=>"011001010",
  33776=>"010000011",
  33777=>"011010100",
  33778=>"101110111",
  33779=>"000000110",
  33780=>"100010001",
  33781=>"100001001",
  33782=>"000000111",
  33783=>"100010100",
  33784=>"110110101",
  33785=>"100011111",
  33786=>"001101001",
  33787=>"011001000",
  33788=>"100110110",
  33789=>"111010100",
  33790=>"000000111",
  33791=>"001001011",
  33792=>"111100101",
  33793=>"100001101",
  33794=>"110101100",
  33795=>"111011011",
  33796=>"010010011",
  33797=>"001101001",
  33798=>"010000010",
  33799=>"100101111",
  33800=>"010100111",
  33801=>"101101100",
  33802=>"011111100",
  33803=>"111011011",
  33804=>"100010001",
  33805=>"110111111",
  33806=>"100000101",
  33807=>"000011000",
  33808=>"101010100",
  33809=>"101111111",
  33810=>"110100101",
  33811=>"111100111",
  33812=>"010000110",
  33813=>"110111101",
  33814=>"000011010",
  33815=>"010111111",
  33816=>"011111110",
  33817=>"000001000",
  33818=>"111110101",
  33819=>"101111000",
  33820=>"111100001",
  33821=>"110101100",
  33822=>"101110101",
  33823=>"010101001",
  33824=>"100011011",
  33825=>"001001011",
  33826=>"011101001",
  33827=>"110101011",
  33828=>"100101111",
  33829=>"010010111",
  33830=>"011011111",
  33831=>"011111000",
  33832=>"011000100",
  33833=>"001111000",
  33834=>"110111000",
  33835=>"010000000",
  33836=>"011111111",
  33837=>"101010001",
  33838=>"010111001",
  33839=>"000111001",
  33840=>"001111111",
  33841=>"010101011",
  33842=>"010101000",
  33843=>"001001111",
  33844=>"010010011",
  33845=>"010010010",
  33846=>"110010111",
  33847=>"111101100",
  33848=>"100100011",
  33849=>"011110010",
  33850=>"110101011",
  33851=>"101110011",
  33852=>"011000010",
  33853=>"110101100",
  33854=>"101001011",
  33855=>"101100000",
  33856=>"100011010",
  33857=>"110101010",
  33858=>"001010101",
  33859=>"011100111",
  33860=>"111000110",
  33861=>"000011010",
  33862=>"000011010",
  33863=>"010101001",
  33864=>"011000001",
  33865=>"111000101",
  33866=>"000101100",
  33867=>"011000001",
  33868=>"010010100",
  33869=>"011110001",
  33870=>"101011001",
  33871=>"000111000",
  33872=>"000000001",
  33873=>"000100100",
  33874=>"100001100",
  33875=>"001101010",
  33876=>"010001001",
  33877=>"100110010",
  33878=>"110110011",
  33879=>"010000000",
  33880=>"011111110",
  33881=>"110001000",
  33882=>"110110101",
  33883=>"011011110",
  33884=>"001000010",
  33885=>"000000111",
  33886=>"110011001",
  33887=>"111101010",
  33888=>"110010001",
  33889=>"000010001",
  33890=>"111001101",
  33891=>"001101100",
  33892=>"011101001",
  33893=>"010001101",
  33894=>"111000001",
  33895=>"101011000",
  33896=>"011001001",
  33897=>"000011100",
  33898=>"001001010",
  33899=>"011001101",
  33900=>"111010111",
  33901=>"011100010",
  33902=>"011101000",
  33903=>"000010100",
  33904=>"110100101",
  33905=>"110011011",
  33906=>"110110010",
  33907=>"000110111",
  33908=>"001100100",
  33909=>"101001011",
  33910=>"100110000",
  33911=>"000101111",
  33912=>"010001011",
  33913=>"101011111",
  33914=>"011110011",
  33915=>"101100100",
  33916=>"011100011",
  33917=>"010110111",
  33918=>"110011001",
  33919=>"010000000",
  33920=>"000011111",
  33921=>"101111000",
  33922=>"001101011",
  33923=>"111001101",
  33924=>"010000000",
  33925=>"100000111",
  33926=>"100010010",
  33927=>"000110001",
  33928=>"000111000",
  33929=>"101110101",
  33930=>"111011101",
  33931=>"111100010",
  33932=>"000010010",
  33933=>"000001101",
  33934=>"100101101",
  33935=>"101101011",
  33936=>"000001111",
  33937=>"001001011",
  33938=>"011010101",
  33939=>"001011100",
  33940=>"011000100",
  33941=>"011011010",
  33942=>"001011001",
  33943=>"010011110",
  33944=>"110111110",
  33945=>"000010110",
  33946=>"101100100",
  33947=>"000101000",
  33948=>"111011100",
  33949=>"111011101",
  33950=>"010010000",
  33951=>"101000101",
  33952=>"111111000",
  33953=>"111101100",
  33954=>"010101011",
  33955=>"100010001",
  33956=>"010110010",
  33957=>"111011001",
  33958=>"111100110",
  33959=>"110110101",
  33960=>"110011010",
  33961=>"001000011",
  33962=>"100100010",
  33963=>"111000101",
  33964=>"010110011",
  33965=>"100001110",
  33966=>"000000111",
  33967=>"100011111",
  33968=>"110010001",
  33969=>"110010001",
  33970=>"111111110",
  33971=>"100010101",
  33972=>"101001101",
  33973=>"011101111",
  33974=>"011101111",
  33975=>"111110001",
  33976=>"101000001",
  33977=>"001010010",
  33978=>"001101110",
  33979=>"001101011",
  33980=>"111000110",
  33981=>"111010011",
  33982=>"110011011",
  33983=>"111111100",
  33984=>"011011001",
  33985=>"111000110",
  33986=>"111110000",
  33987=>"110010101",
  33988=>"100101110",
  33989=>"110001100",
  33990=>"001000100",
  33991=>"100100110",
  33992=>"110001000",
  33993=>"000101000",
  33994=>"110101000",
  33995=>"000111010",
  33996=>"010010100",
  33997=>"110100000",
  33998=>"011001101",
  33999=>"111111101",
  34000=>"011111100",
  34001=>"100110001",
  34002=>"011101000",
  34003=>"111011011",
  34004=>"110101000",
  34005=>"001000001",
  34006=>"110111010",
  34007=>"101010011",
  34008=>"011000000",
  34009=>"011011010",
  34010=>"110100111",
  34011=>"001100111",
  34012=>"110000001",
  34013=>"100101000",
  34014=>"011110000",
  34015=>"100111000",
  34016=>"000111010",
  34017=>"111010010",
  34018=>"001100110",
  34019=>"110100000",
  34020=>"001001000",
  34021=>"100100100",
  34022=>"000010011",
  34023=>"101100100",
  34024=>"110000011",
  34025=>"111010110",
  34026=>"101100010",
  34027=>"100100100",
  34028=>"010001000",
  34029=>"010011011",
  34030=>"001011101",
  34031=>"100001011",
  34032=>"110111101",
  34033=>"000000101",
  34034=>"010101001",
  34035=>"111111111",
  34036=>"100011111",
  34037=>"100101101",
  34038=>"000011111",
  34039=>"001100011",
  34040=>"111101101",
  34041=>"001000010",
  34042=>"111100000",
  34043=>"000001110",
  34044=>"000010001",
  34045=>"000000110",
  34046=>"000011101",
  34047=>"111110101",
  34048=>"000100011",
  34049=>"011010111",
  34050=>"001011111",
  34051=>"101101100",
  34052=>"000101111",
  34053=>"000011011",
  34054=>"010101000",
  34055=>"010101101",
  34056=>"011000010",
  34057=>"100001110",
  34058=>"000000101",
  34059=>"001011111",
  34060=>"011011101",
  34061=>"111101000",
  34062=>"010001100",
  34063=>"001001111",
  34064=>"011001111",
  34065=>"010101100",
  34066=>"100100110",
  34067=>"011101101",
  34068=>"010100110",
  34069=>"111001010",
  34070=>"100111111",
  34071=>"111001111",
  34072=>"111010111",
  34073=>"010011110",
  34074=>"010101101",
  34075=>"010111010",
  34076=>"001111011",
  34077=>"101110110",
  34078=>"111010001",
  34079=>"100011111",
  34080=>"111011100",
  34081=>"001000100",
  34082=>"001100010",
  34083=>"011001111",
  34084=>"010111101",
  34085=>"111110011",
  34086=>"100111110",
  34087=>"001011011",
  34088=>"001110110",
  34089=>"100100011",
  34090=>"011001011",
  34091=>"110010111",
  34092=>"001000010",
  34093=>"011010101",
  34094=>"100001011",
  34095=>"000010110",
  34096=>"100110100",
  34097=>"000011011",
  34098=>"001100001",
  34099=>"001100101",
  34100=>"000010011",
  34101=>"111101010",
  34102=>"111000010",
  34103=>"010010011",
  34104=>"001001100",
  34105=>"100100110",
  34106=>"110111010",
  34107=>"100111011",
  34108=>"111001110",
  34109=>"111001000",
  34110=>"010100101",
  34111=>"000101001",
  34112=>"001010011",
  34113=>"001000001",
  34114=>"111000110",
  34115=>"011001101",
  34116=>"000101000",
  34117=>"100110100",
  34118=>"110100100",
  34119=>"001100000",
  34120=>"010110000",
  34121=>"011101001",
  34122=>"110000101",
  34123=>"100011000",
  34124=>"101110111",
  34125=>"001110101",
  34126=>"001000000",
  34127=>"000111011",
  34128=>"100011001",
  34129=>"101011111",
  34130=>"001000110",
  34131=>"000010001",
  34132=>"000110010",
  34133=>"010100101",
  34134=>"011000011",
  34135=>"100100110",
  34136=>"100101100",
  34137=>"001001111",
  34138=>"101111110",
  34139=>"010000011",
  34140=>"010000101",
  34141=>"011011111",
  34142=>"010111111",
  34143=>"000100010",
  34144=>"101110010",
  34145=>"111100110",
  34146=>"001000000",
  34147=>"100001110",
  34148=>"000110000",
  34149=>"111100111",
  34150=>"110001010",
  34151=>"100000110",
  34152=>"101110101",
  34153=>"000010011",
  34154=>"001001110",
  34155=>"111100001",
  34156=>"101111010",
  34157=>"110110100",
  34158=>"111100110",
  34159=>"100100111",
  34160=>"000011001",
  34161=>"100011001",
  34162=>"001110000",
  34163=>"111011001",
  34164=>"011010011",
  34165=>"100110100",
  34166=>"000111111",
  34167=>"100001000",
  34168=>"000000011",
  34169=>"100110010",
  34170=>"000100000",
  34171=>"100001100",
  34172=>"011000010",
  34173=>"111000000",
  34174=>"001000011",
  34175=>"111110110",
  34176=>"000010000",
  34177=>"100010101",
  34178=>"000111111",
  34179=>"110011010",
  34180=>"101111010",
  34181=>"110000000",
  34182=>"010111010",
  34183=>"100111010",
  34184=>"110000100",
  34185=>"011100100",
  34186=>"101100011",
  34187=>"111010011",
  34188=>"000010110",
  34189=>"000001100",
  34190=>"101110010",
  34191=>"000011001",
  34192=>"000111011",
  34193=>"111100010",
  34194=>"010010010",
  34195=>"110101110",
  34196=>"100100010",
  34197=>"000110111",
  34198=>"010010100",
  34199=>"010100110",
  34200=>"000111100",
  34201=>"100100110",
  34202=>"111100111",
  34203=>"010011000",
  34204=>"011110101",
  34205=>"010001000",
  34206=>"101000111",
  34207=>"001111100",
  34208=>"101011110",
  34209=>"000010001",
  34210=>"110011010",
  34211=>"110000110",
  34212=>"010110110",
  34213=>"010000000",
  34214=>"010101000",
  34215=>"101111101",
  34216=>"011001001",
  34217=>"010101010",
  34218=>"110111101",
  34219=>"111111110",
  34220=>"000000101",
  34221=>"101111010",
  34222=>"011100100",
  34223=>"110100011",
  34224=>"000001100",
  34225=>"100011100",
  34226=>"000010000",
  34227=>"100011110",
  34228=>"010001000",
  34229=>"000011100",
  34230=>"110001010",
  34231=>"010001100",
  34232=>"001000101",
  34233=>"110111110",
  34234=>"001000110",
  34235=>"111111101",
  34236=>"101110101",
  34237=>"101101000",
  34238=>"110011111",
  34239=>"001101010",
  34240=>"110101001",
  34241=>"000001000",
  34242=>"011101001",
  34243=>"011111000",
  34244=>"111111111",
  34245=>"000101011",
  34246=>"001011100",
  34247=>"100010001",
  34248=>"011001011",
  34249=>"011001000",
  34250=>"100111010",
  34251=>"000110000",
  34252=>"011101101",
  34253=>"100100010",
  34254=>"110111110",
  34255=>"001000000",
  34256=>"011000000",
  34257=>"001011001",
  34258=>"000001011",
  34259=>"110110111",
  34260=>"111101000",
  34261=>"001101010",
  34262=>"111101001",
  34263=>"000100101",
  34264=>"010010100",
  34265=>"111111011",
  34266=>"111000101",
  34267=>"111000100",
  34268=>"111001101",
  34269=>"110011110",
  34270=>"110011001",
  34271=>"110110111",
  34272=>"101010111",
  34273=>"111110101",
  34274=>"001000001",
  34275=>"110011011",
  34276=>"011100110",
  34277=>"100011001",
  34278=>"110111111",
  34279=>"110000000",
  34280=>"111100101",
  34281=>"110101111",
  34282=>"110000100",
  34283=>"101110100",
  34284=>"001010101",
  34285=>"000011111",
  34286=>"110001111",
  34287=>"100101100",
  34288=>"001110111",
  34289=>"101110000",
  34290=>"111111011",
  34291=>"101011000",
  34292=>"001011111",
  34293=>"111001100",
  34294=>"101100010",
  34295=>"111101101",
  34296=>"110011100",
  34297=>"100111110",
  34298=>"111010111",
  34299=>"111000000",
  34300=>"000010100",
  34301=>"111111110",
  34302=>"010101011",
  34303=>"111110101",
  34304=>"110111101",
  34305=>"000101100",
  34306=>"001100010",
  34307=>"111010001",
  34308=>"000100011",
  34309=>"101100000",
  34310=>"110001100",
  34311=>"111111011",
  34312=>"011011111",
  34313=>"001100100",
  34314=>"111111011",
  34315=>"111100000",
  34316=>"000100010",
  34317=>"011110110",
  34318=>"101100010",
  34319=>"001010010",
  34320=>"111001111",
  34321=>"011011001",
  34322=>"111010001",
  34323=>"010101100",
  34324=>"011101000",
  34325=>"111100110",
  34326=>"011000111",
  34327=>"010100110",
  34328=>"010011100",
  34329=>"011001001",
  34330=>"010000000",
  34331=>"010110110",
  34332=>"111111101",
  34333=>"010000001",
  34334=>"111000100",
  34335=>"001011010",
  34336=>"101000100",
  34337=>"011010100",
  34338=>"001001011",
  34339=>"110100000",
  34340=>"111101100",
  34341=>"111001110",
  34342=>"110000101",
  34343=>"111000001",
  34344=>"111011111",
  34345=>"111010001",
  34346=>"000100101",
  34347=>"010110011",
  34348=>"011111011",
  34349=>"110100000",
  34350=>"010000111",
  34351=>"101101100",
  34352=>"010011000",
  34353=>"010010101",
  34354=>"010001100",
  34355=>"111101101",
  34356=>"101110010",
  34357=>"010000001",
  34358=>"001111010",
  34359=>"000101100",
  34360=>"110000111",
  34361=>"101100111",
  34362=>"001010101",
  34363=>"110011110",
  34364=>"011001010",
  34365=>"101010011",
  34366=>"011001010",
  34367=>"100011110",
  34368=>"100111100",
  34369=>"000101100",
  34370=>"010111110",
  34371=>"110010010",
  34372=>"100100100",
  34373=>"111010000",
  34374=>"100010001",
  34375=>"100110011",
  34376=>"101101001",
  34377=>"110110110",
  34378=>"111101111",
  34379=>"110001001",
  34380=>"001110111",
  34381=>"000000110",
  34382=>"110010011",
  34383=>"001101111",
  34384=>"010011111",
  34385=>"001111100",
  34386=>"001100000",
  34387=>"000001001",
  34388=>"110001001",
  34389=>"101100100",
  34390=>"011001100",
  34391=>"101111100",
  34392=>"110101100",
  34393=>"100101110",
  34394=>"110100010",
  34395=>"011000111",
  34396=>"001010010",
  34397=>"110101100",
  34398=>"011111011",
  34399=>"011110100",
  34400=>"010101110",
  34401=>"010011000",
  34402=>"100011010",
  34403=>"011010001",
  34404=>"001010000",
  34405=>"001100100",
  34406=>"100001111",
  34407=>"000101000",
  34408=>"110010110",
  34409=>"011001010",
  34410=>"011110010",
  34411=>"100100010",
  34412=>"010011010",
  34413=>"001001000",
  34414=>"000111010",
  34415=>"100011010",
  34416=>"000010101",
  34417=>"000111011",
  34418=>"011001111",
  34419=>"011100001",
  34420=>"101000100",
  34421=>"101001010",
  34422=>"011111011",
  34423=>"001011010",
  34424=>"010101110",
  34425=>"010010100",
  34426=>"110110111",
  34427=>"011110011",
  34428=>"100000010",
  34429=>"101001010",
  34430=>"001000101",
  34431=>"001001110",
  34432=>"011010010",
  34433=>"101000110",
  34434=>"111101001",
  34435=>"000000111",
  34436=>"101001101",
  34437=>"011110000",
  34438=>"111111000",
  34439=>"010110011",
  34440=>"111111000",
  34441=>"001101011",
  34442=>"111101010",
  34443=>"100011011",
  34444=>"011000000",
  34445=>"000110000",
  34446=>"110010010",
  34447=>"001100011",
  34448=>"101000010",
  34449=>"001101110",
  34450=>"110110110",
  34451=>"001011100",
  34452=>"110001101",
  34453=>"010010010",
  34454=>"000100000",
  34455=>"001100100",
  34456=>"011011000",
  34457=>"110100011",
  34458=>"100011100",
  34459=>"101100000",
  34460=>"110100000",
  34461=>"000010110",
  34462=>"010111001",
  34463=>"100111010",
  34464=>"010100110",
  34465=>"010011110",
  34466=>"000111111",
  34467=>"100110011",
  34468=>"001010010",
  34469=>"010011010",
  34470=>"010111010",
  34471=>"101110001",
  34472=>"111010010",
  34473=>"110011101",
  34474=>"011100010",
  34475=>"110011011",
  34476=>"111010011",
  34477=>"010111101",
  34478=>"110010000",
  34479=>"011101000",
  34480=>"010011011",
  34481=>"001001001",
  34482=>"101000101",
  34483=>"111110000",
  34484=>"011111010",
  34485=>"100101100",
  34486=>"001111011",
  34487=>"000001001",
  34488=>"010000000",
  34489=>"101100001",
  34490=>"010111101",
  34491=>"101000101",
  34492=>"110000000",
  34493=>"011110011",
  34494=>"100101010",
  34495=>"111111010",
  34496=>"001100001",
  34497=>"000000100",
  34498=>"110011000",
  34499=>"110100001",
  34500=>"001001110",
  34501=>"010011110",
  34502=>"011111111",
  34503=>"011110100",
  34504=>"000001000",
  34505=>"010100001",
  34506=>"100000101",
  34507=>"111001001",
  34508=>"111010100",
  34509=>"111001110",
  34510=>"000100100",
  34511=>"101101010",
  34512=>"101111101",
  34513=>"001001110",
  34514=>"110011100",
  34515=>"011001000",
  34516=>"111101011",
  34517=>"011001110",
  34518=>"001000111",
  34519=>"111010100",
  34520=>"101100011",
  34521=>"000001010",
  34522=>"011001110",
  34523=>"100001010",
  34524=>"101101000",
  34525=>"010001000",
  34526=>"111010101",
  34527=>"001001110",
  34528=>"101100110",
  34529=>"110010110",
  34530=>"000000111",
  34531=>"000111011",
  34532=>"000101000",
  34533=>"000000110",
  34534=>"001110000",
  34535=>"101110000",
  34536=>"101011000",
  34537=>"110111111",
  34538=>"010000000",
  34539=>"001100001",
  34540=>"001101111",
  34541=>"010110100",
  34542=>"100111001",
  34543=>"111010000",
  34544=>"110001101",
  34545=>"101110011",
  34546=>"001000110",
  34547=>"110110010",
  34548=>"100111110",
  34549=>"101111010",
  34550=>"100100001",
  34551=>"001101001",
  34552=>"111111100",
  34553=>"011110000",
  34554=>"011101000",
  34555=>"000101001",
  34556=>"011001010",
  34557=>"011100111",
  34558=>"111111111",
  34559=>"111011001",
  34560=>"101101011",
  34561=>"110000000",
  34562=>"010011011",
  34563=>"110100001",
  34564=>"111100011",
  34565=>"011101100",
  34566=>"100001010",
  34567=>"110111110",
  34568=>"011101110",
  34569=>"010101111",
  34570=>"000100010",
  34571=>"011001011",
  34572=>"000010000",
  34573=>"110101001",
  34574=>"001101101",
  34575=>"011110011",
  34576=>"000100111",
  34577=>"101101000",
  34578=>"111000010",
  34579=>"001000001",
  34580=>"011111100",
  34581=>"010010100",
  34582=>"000000001",
  34583=>"011101100",
  34584=>"010011000",
  34585=>"100101101",
  34586=>"100111010",
  34587=>"100101001",
  34588=>"111000010",
  34589=>"110111100",
  34590=>"101101010",
  34591=>"110110110",
  34592=>"100110011",
  34593=>"111110110",
  34594=>"111101001",
  34595=>"110110010",
  34596=>"111011110",
  34597=>"000000011",
  34598=>"001111111",
  34599=>"000000001",
  34600=>"100101001",
  34601=>"001100101",
  34602=>"111001001",
  34603=>"010001001",
  34604=>"000011110",
  34605=>"011101101",
  34606=>"011001001",
  34607=>"101110111",
  34608=>"110010110",
  34609=>"000100100",
  34610=>"010011101",
  34611=>"000010100",
  34612=>"111101011",
  34613=>"010111110",
  34614=>"110111101",
  34615=>"011011001",
  34616=>"110101011",
  34617=>"111011010",
  34618=>"011100111",
  34619=>"010111011",
  34620=>"010110111",
  34621=>"000100000",
  34622=>"011001010",
  34623=>"010111010",
  34624=>"000110001",
  34625=>"010100110",
  34626=>"001000000",
  34627=>"000111000",
  34628=>"100010100",
  34629=>"100101101",
  34630=>"010100100",
  34631=>"000110000",
  34632=>"001101000",
  34633=>"110101110",
  34634=>"010100010",
  34635=>"001110010",
  34636=>"010011100",
  34637=>"101111000",
  34638=>"001110001",
  34639=>"010010111",
  34640=>"100100100",
  34641=>"000011101",
  34642=>"111101111",
  34643=>"000001011",
  34644=>"010000111",
  34645=>"000001011",
  34646=>"100111111",
  34647=>"101001110",
  34648=>"011101011",
  34649=>"100101010",
  34650=>"110100110",
  34651=>"000101001",
  34652=>"110111101",
  34653=>"101011011",
  34654=>"001010101",
  34655=>"010111000",
  34656=>"000010000",
  34657=>"101000010",
  34658=>"011010001",
  34659=>"010000110",
  34660=>"110001011",
  34661=>"011100101",
  34662=>"010010000",
  34663=>"011110111",
  34664=>"001001011",
  34665=>"010011101",
  34666=>"101110000",
  34667=>"010010100",
  34668=>"000000010",
  34669=>"000110010",
  34670=>"101100100",
  34671=>"010110011",
  34672=>"001101001",
  34673=>"110101101",
  34674=>"101101011",
  34675=>"111000010",
  34676=>"101110100",
  34677=>"000011111",
  34678=>"111101011",
  34679=>"111111000",
  34680=>"101001111",
  34681=>"001000000",
  34682=>"110000001",
  34683=>"100110111",
  34684=>"100001001",
  34685=>"011100001",
  34686=>"010000001",
  34687=>"111111001",
  34688=>"000011001",
  34689=>"010111110",
  34690=>"000000011",
  34691=>"001000001",
  34692=>"100101111",
  34693=>"110101101",
  34694=>"101111110",
  34695=>"001011001",
  34696=>"101001111",
  34697=>"111010011",
  34698=>"011000000",
  34699=>"111110100",
  34700=>"000111101",
  34701=>"100100111",
  34702=>"110111011",
  34703=>"001110101",
  34704=>"011011100",
  34705=>"111000010",
  34706=>"000010011",
  34707=>"011111101",
  34708=>"011011010",
  34709=>"100110101",
  34710=>"001111101",
  34711=>"110000011",
  34712=>"010001001",
  34713=>"101110001",
  34714=>"000101010",
  34715=>"001100011",
  34716=>"001110111",
  34717=>"111110100",
  34718=>"111111100",
  34719=>"101001001",
  34720=>"000101010",
  34721=>"101111110",
  34722=>"111110101",
  34723=>"000010000",
  34724=>"111000001",
  34725=>"010110010",
  34726=>"000110110",
  34727=>"100000101",
  34728=>"101111000",
  34729=>"111110101",
  34730=>"101101011",
  34731=>"001100001",
  34732=>"100000110",
  34733=>"011101000",
  34734=>"101100110",
  34735=>"100101101",
  34736=>"101101010",
  34737=>"000100011",
  34738=>"000101101",
  34739=>"101111001",
  34740=>"001011100",
  34741=>"101010000",
  34742=>"001001010",
  34743=>"010011100",
  34744=>"110101110",
  34745=>"100000110",
  34746=>"011011101",
  34747=>"011100101",
  34748=>"110110010",
  34749=>"001111011",
  34750=>"111011110",
  34751=>"000111010",
  34752=>"001110001",
  34753=>"001100100",
  34754=>"001000000",
  34755=>"001100011",
  34756=>"101110011",
  34757=>"101111110",
  34758=>"010011011",
  34759=>"001010011",
  34760=>"010101100",
  34761=>"000101000",
  34762=>"110100000",
  34763=>"101110011",
  34764=>"110000100",
  34765=>"000111100",
  34766=>"010001111",
  34767=>"001010001",
  34768=>"111101000",
  34769=>"111100001",
  34770=>"001011111",
  34771=>"110001100",
  34772=>"000100100",
  34773=>"111111010",
  34774=>"001101111",
  34775=>"100111011",
  34776=>"000000110",
  34777=>"100100001",
  34778=>"111110010",
  34779=>"111100111",
  34780=>"010100111",
  34781=>"001001100",
  34782=>"100000000",
  34783=>"010101010",
  34784=>"110001011",
  34785=>"101000100",
  34786=>"110010111",
  34787=>"001100111",
  34788=>"000100100",
  34789=>"101100110",
  34790=>"000100001",
  34791=>"011111111",
  34792=>"100110010",
  34793=>"010000101",
  34794=>"010111011",
  34795=>"101000111",
  34796=>"101111111",
  34797=>"100100101",
  34798=>"101101010",
  34799=>"001001100",
  34800=>"000001110",
  34801=>"111100000",
  34802=>"001011011",
  34803=>"010101001",
  34804=>"001100011",
  34805=>"001111111",
  34806=>"101100000",
  34807=>"101000000",
  34808=>"111001100",
  34809=>"110010001",
  34810=>"000100011",
  34811=>"100011111",
  34812=>"011111110",
  34813=>"000101110",
  34814=>"000001000",
  34815=>"111100111",
  34816=>"101010101",
  34817=>"100111010",
  34818=>"101100111",
  34819=>"000001000",
  34820=>"011001100",
  34821=>"101101011",
  34822=>"111111000",
  34823=>"000000011",
  34824=>"010101000",
  34825=>"111111001",
  34826=>"001011011",
  34827=>"010100010",
  34828=>"011000000",
  34829=>"111011010",
  34830=>"100110010",
  34831=>"101011010",
  34832=>"101100011",
  34833=>"011011101",
  34834=>"111111110",
  34835=>"011100000",
  34836=>"010011101",
  34837=>"100111011",
  34838=>"100100011",
  34839=>"001000000",
  34840=>"011110001",
  34841=>"000011111",
  34842=>"001111110",
  34843=>"010001110",
  34844=>"110101011",
  34845=>"100000000",
  34846=>"100010010",
  34847=>"010011000",
  34848=>"111001100",
  34849=>"001101111",
  34850=>"010011001",
  34851=>"000001011",
  34852=>"011101111",
  34853=>"010100011",
  34854=>"100001001",
  34855=>"001111101",
  34856=>"001111101",
  34857=>"100110011",
  34858=>"101110111",
  34859=>"101000001",
  34860=>"100001010",
  34861=>"000001001",
  34862=>"001100110",
  34863=>"111111001",
  34864=>"111010111",
  34865=>"001101100",
  34866=>"111111000",
  34867=>"101100101",
  34868=>"011100011",
  34869=>"001001110",
  34870=>"100101011",
  34871=>"000011011",
  34872=>"101000111",
  34873=>"001011111",
  34874=>"111011001",
  34875=>"000101100",
  34876=>"001100010",
  34877=>"010000100",
  34878=>"100001001",
  34879=>"111001010",
  34880=>"000110110",
  34881=>"010000010",
  34882=>"011011001",
  34883=>"001110001",
  34884=>"111111100",
  34885=>"010000101",
  34886=>"100111000",
  34887=>"001000110",
  34888=>"010100100",
  34889=>"101111110",
  34890=>"010110000",
  34891=>"110100111",
  34892=>"111100010",
  34893=>"011000110",
  34894=>"000110011",
  34895=>"101010110",
  34896=>"100000110",
  34897=>"110010000",
  34898=>"111000100",
  34899=>"101000101",
  34900=>"111011110",
  34901=>"010001000",
  34902=>"001001011",
  34903=>"000000111",
  34904=>"001000010",
  34905=>"011110000",
  34906=>"101110011",
  34907=>"000001111",
  34908=>"010000001",
  34909=>"101100111",
  34910=>"100001000",
  34911=>"101101010",
  34912=>"000110110",
  34913=>"111001101",
  34914=>"000000000",
  34915=>"100001011",
  34916=>"000101011",
  34917=>"110101110",
  34918=>"111011111",
  34919=>"001010001",
  34920=>"000010010",
  34921=>"011111011",
  34922=>"101011010",
  34923=>"110010100",
  34924=>"101110101",
  34925=>"101001101",
  34926=>"111001011",
  34927=>"001100001",
  34928=>"111000100",
  34929=>"000010101",
  34930=>"100011010",
  34931=>"000010000",
  34932=>"011111011",
  34933=>"011100000",
  34934=>"001001111",
  34935=>"101001100",
  34936=>"100100100",
  34937=>"011010010",
  34938=>"101111000",
  34939=>"001001110",
  34940=>"111010011",
  34941=>"000001111",
  34942=>"111001111",
  34943=>"001100111",
  34944=>"111111011",
  34945=>"110000011",
  34946=>"000000001",
  34947=>"001110000",
  34948=>"000001110",
  34949=>"001101110",
  34950=>"011000111",
  34951=>"000001010",
  34952=>"011011010",
  34953=>"101000001",
  34954=>"000000101",
  34955=>"111110101",
  34956=>"101100000",
  34957=>"111101010",
  34958=>"011000111",
  34959=>"110110010",
  34960=>"101011100",
  34961=>"110101001",
  34962=>"011000000",
  34963=>"101011011",
  34964=>"010001110",
  34965=>"100100010",
  34966=>"000101011",
  34967=>"100001110",
  34968=>"100100001",
  34969=>"011110001",
  34970=>"101000100",
  34971=>"100011011",
  34972=>"011100110",
  34973=>"111010001",
  34974=>"101010000",
  34975=>"101101001",
  34976=>"010110001",
  34977=>"110010010",
  34978=>"010000010",
  34979=>"101111000",
  34980=>"011100000",
  34981=>"010001000",
  34982=>"111110001",
  34983=>"111011100",
  34984=>"100010000",
  34985=>"011011000",
  34986=>"101011100",
  34987=>"111111110",
  34988=>"001101110",
  34989=>"010001001",
  34990=>"001000010",
  34991=>"010011001",
  34992=>"010110000",
  34993=>"000110010",
  34994=>"000011000",
  34995=>"101111011",
  34996=>"101100011",
  34997=>"101000011",
  34998=>"101001101",
  34999=>"100001101",
  35000=>"011000100",
  35001=>"110111011",
  35002=>"011100000",
  35003=>"111111010",
  35004=>"001101010",
  35005=>"101000111",
  35006=>"000010100",
  35007=>"001110011",
  35008=>"110100111",
  35009=>"001001011",
  35010=>"001100110",
  35011=>"010111100",
  35012=>"001100111",
  35013=>"010101001",
  35014=>"111010101",
  35015=>"000110010",
  35016=>"101000111",
  35017=>"000001011",
  35018=>"100111111",
  35019=>"101101100",
  35020=>"110100001",
  35021=>"100111101",
  35022=>"000011101",
  35023=>"110101101",
  35024=>"010100010",
  35025=>"011101000",
  35026=>"101101100",
  35027=>"100111110",
  35028=>"011110100",
  35029=>"010001001",
  35030=>"100100011",
  35031=>"010001001",
  35032=>"110001000",
  35033=>"110101101",
  35034=>"010110001",
  35035=>"011101000",
  35036=>"011000101",
  35037=>"110000110",
  35038=>"011100010",
  35039=>"001100011",
  35040=>"111101001",
  35041=>"101101010",
  35042=>"001111100",
  35043=>"001100010",
  35044=>"011101010",
  35045=>"111100011",
  35046=>"100000100",
  35047=>"011110111",
  35048=>"100100010",
  35049=>"110111110",
  35050=>"001111000",
  35051=>"010100000",
  35052=>"111101110",
  35053=>"100101100",
  35054=>"001101000",
  35055=>"000111101",
  35056=>"011100101",
  35057=>"101001100",
  35058=>"001110111",
  35059=>"100010011",
  35060=>"010000101",
  35061=>"100010100",
  35062=>"101110100",
  35063=>"000110100",
  35064=>"011110011",
  35065=>"000100100",
  35066=>"111010101",
  35067=>"100000000",
  35068=>"000010011",
  35069=>"101100001",
  35070=>"011011100",
  35071=>"100011111",
  35072=>"100010011",
  35073=>"001011101",
  35074=>"111100001",
  35075=>"001001111",
  35076=>"010001001",
  35077=>"001100111",
  35078=>"100110100",
  35079=>"111011100",
  35080=>"010001001",
  35081=>"011010011",
  35082=>"111111101",
  35083=>"100110100",
  35084=>"101010010",
  35085=>"001100100",
  35086=>"111101111",
  35087=>"110001110",
  35088=>"110100111",
  35089=>"101011010",
  35090=>"010010111",
  35091=>"011100110",
  35092=>"100001001",
  35093=>"011010000",
  35094=>"010001110",
  35095=>"101101001",
  35096=>"110111000",
  35097=>"111100101",
  35098=>"101100000",
  35099=>"000010001",
  35100=>"110010010",
  35101=>"110001010",
  35102=>"000001100",
  35103=>"000001011",
  35104=>"001000100",
  35105=>"110100001",
  35106=>"001010011",
  35107=>"010100100",
  35108=>"001111011",
  35109=>"100001000",
  35110=>"111001110",
  35111=>"111111111",
  35112=>"011001011",
  35113=>"100011001",
  35114=>"011000000",
  35115=>"100011110",
  35116=>"110010001",
  35117=>"001001010",
  35118=>"010000011",
  35119=>"010100110",
  35120=>"100100101",
  35121=>"110100101",
  35122=>"010010111",
  35123=>"001010110",
  35124=>"101111001",
  35125=>"111111010",
  35126=>"111101111",
  35127=>"100001100",
  35128=>"001100101",
  35129=>"010101111",
  35130=>"110011100",
  35131=>"010100110",
  35132=>"111000110",
  35133=>"100110000",
  35134=>"110011010",
  35135=>"000111111",
  35136=>"101001011",
  35137=>"101101100",
  35138=>"000010110",
  35139=>"100000101",
  35140=>"110101111",
  35141=>"010101111",
  35142=>"000001100",
  35143=>"001100011",
  35144=>"100111000",
  35145=>"101110000",
  35146=>"011010100",
  35147=>"000101011",
  35148=>"010011100",
  35149=>"001000011",
  35150=>"010110111",
  35151=>"110110011",
  35152=>"111011111",
  35153=>"011001010",
  35154=>"100000101",
  35155=>"001001011",
  35156=>"111010010",
  35157=>"001110100",
  35158=>"100111100",
  35159=>"111000110",
  35160=>"101000111",
  35161=>"110000001",
  35162=>"000111101",
  35163=>"111010111",
  35164=>"111000001",
  35165=>"000000001",
  35166=>"111111110",
  35167=>"001110101",
  35168=>"001111110",
  35169=>"101000000",
  35170=>"000101101",
  35171=>"111010011",
  35172=>"001000010",
  35173=>"100110111",
  35174=>"001110110",
  35175=>"010000001",
  35176=>"011001101",
  35177=>"000111010",
  35178=>"100010000",
  35179=>"101111111",
  35180=>"111011101",
  35181=>"110111101",
  35182=>"011000101",
  35183=>"001010100",
  35184=>"001011000",
  35185=>"101000011",
  35186=>"000010100",
  35187=>"010001000",
  35188=>"101000111",
  35189=>"010101010",
  35190=>"000101000",
  35191=>"100000111",
  35192=>"000110110",
  35193=>"111001000",
  35194=>"000011100",
  35195=>"111001010",
  35196=>"001101001",
  35197=>"000110110",
  35198=>"100110010",
  35199=>"001101100",
  35200=>"010011000",
  35201=>"001100111",
  35202=>"001001000",
  35203=>"111000101",
  35204=>"010100010",
  35205=>"000000111",
  35206=>"111111111",
  35207=>"100101111",
  35208=>"000001010",
  35209=>"101110100",
  35210=>"100011000",
  35211=>"100000101",
  35212=>"010111110",
  35213=>"000110110",
  35214=>"000001001",
  35215=>"100010101",
  35216=>"010101110",
  35217=>"000011111",
  35218=>"000110000",
  35219=>"011100010",
  35220=>"010110011",
  35221=>"111011011",
  35222=>"111111010",
  35223=>"100111001",
  35224=>"001010001",
  35225=>"000101111",
  35226=>"000010111",
  35227=>"010100100",
  35228=>"111010100",
  35229=>"110000111",
  35230=>"100100110",
  35231=>"001011100",
  35232=>"100000011",
  35233=>"010010000",
  35234=>"000101110",
  35235=>"010010010",
  35236=>"111001111",
  35237=>"010000100",
  35238=>"010111010",
  35239=>"000101000",
  35240=>"000100011",
  35241=>"101110011",
  35242=>"101011001",
  35243=>"000110011",
  35244=>"111100110",
  35245=>"111111000",
  35246=>"111110010",
  35247=>"011001000",
  35248=>"011010000",
  35249=>"000001011",
  35250=>"011101011",
  35251=>"011001000",
  35252=>"110011001",
  35253=>"000110100",
  35254=>"000110100",
  35255=>"000100001",
  35256=>"111010111",
  35257=>"000101100",
  35258=>"110000101",
  35259=>"101000010",
  35260=>"100110111",
  35261=>"010010111",
  35262=>"111011111",
  35263=>"001111101",
  35264=>"011000010",
  35265=>"001110011",
  35266=>"011101100",
  35267=>"101001100",
  35268=>"001010000",
  35269=>"100110001",
  35270=>"111001000",
  35271=>"100100101",
  35272=>"010000111",
  35273=>"010010110",
  35274=>"101011010",
  35275=>"111100011",
  35276=>"110010011",
  35277=>"011111001",
  35278=>"001000100",
  35279=>"000110000",
  35280=>"010000011",
  35281=>"000001100",
  35282=>"100001100",
  35283=>"100001010",
  35284=>"000000001",
  35285=>"000001000",
  35286=>"100000001",
  35287=>"001001001",
  35288=>"110011001",
  35289=>"100000001",
  35290=>"111110101",
  35291=>"010010101",
  35292=>"000101001",
  35293=>"011011010",
  35294=>"010000011",
  35295=>"110010111",
  35296=>"011101100",
  35297=>"001011011",
  35298=>"111101111",
  35299=>"110010110",
  35300=>"001001011",
  35301=>"100110010",
  35302=>"001101010",
  35303=>"000000111",
  35304=>"101011000",
  35305=>"110000111",
  35306=>"000000011",
  35307=>"111101010",
  35308=>"001011011",
  35309=>"111001000",
  35310=>"011101010",
  35311=>"001100110",
  35312=>"000011010",
  35313=>"101010011",
  35314=>"111101110",
  35315=>"101110101",
  35316=>"100001100",
  35317=>"001101110",
  35318=>"001100100",
  35319=>"100100101",
  35320=>"111010010",
  35321=>"100110110",
  35322=>"000011001",
  35323=>"100101101",
  35324=>"101001101",
  35325=>"111011101",
  35326=>"110111101",
  35327=>"011001110",
  35328=>"100001001",
  35329=>"000101000",
  35330=>"110101101",
  35331=>"101000100",
  35332=>"110110110",
  35333=>"011001001",
  35334=>"000011111",
  35335=>"110000011",
  35336=>"001101110",
  35337=>"000000101",
  35338=>"111100101",
  35339=>"000111110",
  35340=>"001010100",
  35341=>"000010001",
  35342=>"110011111",
  35343=>"100011011",
  35344=>"011010100",
  35345=>"000110111",
  35346=>"010000000",
  35347=>"111111001",
  35348=>"011101011",
  35349=>"010000001",
  35350=>"010011001",
  35351=>"111111001",
  35352=>"111001100",
  35353=>"011111010",
  35354=>"000111001",
  35355=>"000101110",
  35356=>"010110100",
  35357=>"010010111",
  35358=>"110001101",
  35359=>"111111100",
  35360=>"001000010",
  35361=>"111101111",
  35362=>"001011100",
  35363=>"001001010",
  35364=>"101111011",
  35365=>"000101111",
  35366=>"110000110",
  35367=>"111110100",
  35368=>"011010111",
  35369=>"100110100",
  35370=>"011011010",
  35371=>"100110111",
  35372=>"110011101",
  35373=>"111101100",
  35374=>"111100001",
  35375=>"111111100",
  35376=>"110010110",
  35377=>"110001000",
  35378=>"111010000",
  35379=>"110000011",
  35380=>"100001000",
  35381=>"000110000",
  35382=>"100100111",
  35383=>"100010100",
  35384=>"111100000",
  35385=>"000111000",
  35386=>"101001111",
  35387=>"010110001",
  35388=>"010001010",
  35389=>"011010010",
  35390=>"011010000",
  35391=>"100010110",
  35392=>"111111100",
  35393=>"110010010",
  35394=>"101111011",
  35395=>"011100111",
  35396=>"010111011",
  35397=>"001111001",
  35398=>"001010100",
  35399=>"100111011",
  35400=>"111111000",
  35401=>"011000100",
  35402=>"001111111",
  35403=>"100001101",
  35404=>"000110010",
  35405=>"001111000",
  35406=>"000111100",
  35407=>"111010000",
  35408=>"010111001",
  35409=>"001111100",
  35410=>"111101000",
  35411=>"110110100",
  35412=>"011010111",
  35413=>"100001000",
  35414=>"110100011",
  35415=>"110111111",
  35416=>"111110111",
  35417=>"110111010",
  35418=>"001011010",
  35419=>"000000110",
  35420=>"001000001",
  35421=>"110101101",
  35422=>"111111001",
  35423=>"100101101",
  35424=>"011110000",
  35425=>"001010010",
  35426=>"100111110",
  35427=>"101000000",
  35428=>"011100010",
  35429=>"100010001",
  35430=>"000001010",
  35431=>"011101111",
  35432=>"100001011",
  35433=>"010001101",
  35434=>"100011010",
  35435=>"101100001",
  35436=>"110000110",
  35437=>"111100110",
  35438=>"111101101",
  35439=>"000101011",
  35440=>"000000000",
  35441=>"001111011",
  35442=>"001100000",
  35443=>"110111011",
  35444=>"001010010",
  35445=>"011101101",
  35446=>"000101111",
  35447=>"000111100",
  35448=>"010010010",
  35449=>"110000010",
  35450=>"010101110",
  35451=>"010110111",
  35452=>"101010000",
  35453=>"110010110",
  35454=>"100001000",
  35455=>"010010110",
  35456=>"000101101",
  35457=>"111010010",
  35458=>"101000000",
  35459=>"000111111",
  35460=>"011001010",
  35461=>"000100000",
  35462=>"100110000",
  35463=>"110101111",
  35464=>"000101011",
  35465=>"011100100",
  35466=>"010110101",
  35467=>"111001101",
  35468=>"001100101",
  35469=>"000000111",
  35470=>"101101000",
  35471=>"100100000",
  35472=>"101001101",
  35473=>"011110100",
  35474=>"011011100",
  35475=>"111000110",
  35476=>"011010101",
  35477=>"000011100",
  35478=>"100001000",
  35479=>"011111011",
  35480=>"010110101",
  35481=>"000101001",
  35482=>"010000011",
  35483=>"100010000",
  35484=>"110100000",
  35485=>"101111111",
  35486=>"111001100",
  35487=>"011011101",
  35488=>"110101010",
  35489=>"111100011",
  35490=>"110000111",
  35491=>"011011110",
  35492=>"011010101",
  35493=>"101101111",
  35494=>"110110001",
  35495=>"000001000",
  35496=>"011000011",
  35497=>"111010100",
  35498=>"010101000",
  35499=>"010101110",
  35500=>"010001111",
  35501=>"110010010",
  35502=>"001100010",
  35503=>"111010011",
  35504=>"010010010",
  35505=>"100100000",
  35506=>"100101101",
  35507=>"001010110",
  35508=>"101001000",
  35509=>"000110111",
  35510=>"111010010",
  35511=>"110100111",
  35512=>"111101111",
  35513=>"010110101",
  35514=>"101100111",
  35515=>"100100000",
  35516=>"000101001",
  35517=>"001000000",
  35518=>"110111100",
  35519=>"100010011",
  35520=>"001110000",
  35521=>"110110100",
  35522=>"110111111",
  35523=>"010100010",
  35524=>"110000001",
  35525=>"100111001",
  35526=>"000110000",
  35527=>"110101000",
  35528=>"000000101",
  35529=>"000101000",
  35530=>"100010110",
  35531=>"000001110",
  35532=>"100110001",
  35533=>"111000111",
  35534=>"100110001",
  35535=>"010011000",
  35536=>"101101101",
  35537=>"110111010",
  35538=>"010110001",
  35539=>"100101101",
  35540=>"011101000",
  35541=>"000011111",
  35542=>"011000001",
  35543=>"100010011",
  35544=>"010100100",
  35545=>"111011000",
  35546=>"111011111",
  35547=>"100100010",
  35548=>"001001001",
  35549=>"010000000",
  35550=>"011111000",
  35551=>"011010000",
  35552=>"000010011",
  35553=>"101001111",
  35554=>"101101111",
  35555=>"111001100",
  35556=>"110010000",
  35557=>"000110111",
  35558=>"000001010",
  35559=>"100100101",
  35560=>"100010001",
  35561=>"000110100",
  35562=>"100100011",
  35563=>"010011011",
  35564=>"010001000",
  35565=>"001111101",
  35566=>"011110101",
  35567=>"101011011",
  35568=>"100000111",
  35569=>"110111011",
  35570=>"001011011",
  35571=>"100111110",
  35572=>"100101111",
  35573=>"111101111",
  35574=>"010111000",
  35575=>"010011101",
  35576=>"101010100",
  35577=>"011100000",
  35578=>"110010000",
  35579=>"010000111",
  35580=>"110010111",
  35581=>"001111100",
  35582=>"000010000",
  35583=>"100111011",
  35584=>"111001001",
  35585=>"101000100",
  35586=>"011111111",
  35587=>"001000110",
  35588=>"101010000",
  35589=>"101111101",
  35590=>"000010101",
  35591=>"001110100",
  35592=>"100010011",
  35593=>"110010001",
  35594=>"101101101",
  35595=>"001110000",
  35596=>"000001011",
  35597=>"101110110",
  35598=>"000010010",
  35599=>"011100110",
  35600=>"001111001",
  35601=>"000001111",
  35602=>"111000111",
  35603=>"100001001",
  35604=>"010110001",
  35605=>"110100110",
  35606=>"011101010",
  35607=>"001100100",
  35608=>"011110011",
  35609=>"111100101",
  35610=>"011111001",
  35611=>"100001101",
  35612=>"001111100",
  35613=>"010100111",
  35614=>"010000000",
  35615=>"101101101",
  35616=>"111111011",
  35617=>"100010101",
  35618=>"100000101",
  35619=>"001010010",
  35620=>"101110101",
  35621=>"011111111",
  35622=>"110100110",
  35623=>"010010010",
  35624=>"010011100",
  35625=>"000101001",
  35626=>"000001111",
  35627=>"110110011",
  35628=>"110000011",
  35629=>"110100011",
  35630=>"001100000",
  35631=>"000000100",
  35632=>"000000000",
  35633=>"110101011",
  35634=>"111010100",
  35635=>"111000001",
  35636=>"000101011",
  35637=>"101100100",
  35638=>"110010111",
  35639=>"001110010",
  35640=>"110110000",
  35641=>"110010110",
  35642=>"010101010",
  35643=>"000001011",
  35644=>"101111101",
  35645=>"011010100",
  35646=>"000010101",
  35647=>"111001001",
  35648=>"010100011",
  35649=>"101111000",
  35650=>"110110011",
  35651=>"111001111",
  35652=>"100101100",
  35653=>"111010111",
  35654=>"100111111",
  35655=>"000000011",
  35656=>"100001111",
  35657=>"111101000",
  35658=>"000001000",
  35659=>"101110010",
  35660=>"111011100",
  35661=>"111101001",
  35662=>"110001100",
  35663=>"000110001",
  35664=>"001010110",
  35665=>"010010010",
  35666=>"010110010",
  35667=>"011101000",
  35668=>"100010111",
  35669=>"101000100",
  35670=>"000010001",
  35671=>"000100011",
  35672=>"001111100",
  35673=>"110111000",
  35674=>"101101100",
  35675=>"100101101",
  35676=>"111010000",
  35677=>"111011100",
  35678=>"111011110",
  35679=>"000100101",
  35680=>"010011001",
  35681=>"101001101",
  35682=>"110110011",
  35683=>"010110000",
  35684=>"100100110",
  35685=>"010001011",
  35686=>"101000000",
  35687=>"100100110",
  35688=>"000011110",
  35689=>"100010101",
  35690=>"111100000",
  35691=>"110001001",
  35692=>"011001001",
  35693=>"001010011",
  35694=>"001101001",
  35695=>"010110100",
  35696=>"001001101",
  35697=>"001110100",
  35698=>"100011100",
  35699=>"111000100",
  35700=>"100000100",
  35701=>"101011010",
  35702=>"011101000",
  35703=>"001010110",
  35704=>"011011110",
  35705=>"100001000",
  35706=>"000010000",
  35707=>"010101011",
  35708=>"000000000",
  35709=>"101100010",
  35710=>"010010110",
  35711=>"011001001",
  35712=>"101101010",
  35713=>"111101011",
  35714=>"000111010",
  35715=>"000000110",
  35716=>"100010011",
  35717=>"100001101",
  35718=>"011001001",
  35719=>"000001100",
  35720=>"100000111",
  35721=>"101000001",
  35722=>"110110010",
  35723=>"011110010",
  35724=>"011111101",
  35725=>"001000011",
  35726=>"001100001",
  35727=>"101101100",
  35728=>"010001001",
  35729=>"010011110",
  35730=>"000010000",
  35731=>"101111100",
  35732=>"001111010",
  35733=>"001011001",
  35734=>"100010010",
  35735=>"100100101",
  35736=>"001010110",
  35737=>"100110000",
  35738=>"111110100",
  35739=>"001000101",
  35740=>"000000010",
  35741=>"011000011",
  35742=>"010001101",
  35743=>"000001100",
  35744=>"000111100",
  35745=>"011001101",
  35746=>"000000111",
  35747=>"010101100",
  35748=>"011010011",
  35749=>"000111110",
  35750=>"000101100",
  35751=>"010100111",
  35752=>"001000011",
  35753=>"010001000",
  35754=>"010010100",
  35755=>"111101001",
  35756=>"011001101",
  35757=>"100011010",
  35758=>"000101011",
  35759=>"010100110",
  35760=>"110101100",
  35761=>"111001110",
  35762=>"001101001",
  35763=>"001010010",
  35764=>"010101100",
  35765=>"110010111",
  35766=>"010000000",
  35767=>"001110100",
  35768=>"101101000",
  35769=>"100000010",
  35770=>"110101101",
  35771=>"001110010",
  35772=>"010101110",
  35773=>"101011011",
  35774=>"000100100",
  35775=>"101011100",
  35776=>"000010001",
  35777=>"101110011",
  35778=>"001001011",
  35779=>"001010000",
  35780=>"100000000",
  35781=>"000111100",
  35782=>"001100110",
  35783=>"100111000",
  35784=>"001100110",
  35785=>"000001000",
  35786=>"111110001",
  35787=>"111000110",
  35788=>"010001110",
  35789=>"110100000",
  35790=>"101100100",
  35791=>"100001000",
  35792=>"101111110",
  35793=>"000000101",
  35794=>"011111111",
  35795=>"100001101",
  35796=>"110101101",
  35797=>"001101100",
  35798=>"000100001",
  35799=>"101000001",
  35800=>"110100111",
  35801=>"000100001",
  35802=>"011101110",
  35803=>"000100110",
  35804=>"011000001",
  35805=>"101010111",
  35806=>"001101101",
  35807=>"111011111",
  35808=>"010101110",
  35809=>"000010101",
  35810=>"000001100",
  35811=>"000000101",
  35812=>"010000000",
  35813=>"111111000",
  35814=>"010101011",
  35815=>"000001001",
  35816=>"111101000",
  35817=>"011001111",
  35818=>"111101100",
  35819=>"110101000",
  35820=>"011101111",
  35821=>"001001010",
  35822=>"000000010",
  35823=>"000010000",
  35824=>"000000000",
  35825=>"111001111",
  35826=>"001000100",
  35827=>"000110101",
  35828=>"100000110",
  35829=>"001010000",
  35830=>"100000000",
  35831=>"100001100",
  35832=>"101010000",
  35833=>"101110001",
  35834=>"001010100",
  35835=>"100100100",
  35836=>"011101000",
  35837=>"000111100",
  35838=>"110000001",
  35839=>"010111010",
  35840=>"010001100",
  35841=>"010110011",
  35842=>"100101101",
  35843=>"101110011",
  35844=>"111000111",
  35845=>"101101110",
  35846=>"110111010",
  35847=>"010101001",
  35848=>"111111011",
  35849=>"011010101",
  35850=>"100110100",
  35851=>"011011101",
  35852=>"100100011",
  35853=>"100010000",
  35854=>"001100110",
  35855=>"000101010",
  35856=>"100111110",
  35857=>"011000110",
  35858=>"101000101",
  35859=>"110111001",
  35860=>"100000000",
  35861=>"001111100",
  35862=>"010111011",
  35863=>"001101010",
  35864=>"001111001",
  35865=>"001001000",
  35866=>"111010101",
  35867=>"100111000",
  35868=>"100000011",
  35869=>"001010011",
  35870=>"010100011",
  35871=>"110110001",
  35872=>"111001001",
  35873=>"101010100",
  35874=>"110100101",
  35875=>"000010100",
  35876=>"101110011",
  35877=>"010111110",
  35878=>"000011001",
  35879=>"101001110",
  35880=>"000011000",
  35881=>"001100000",
  35882=>"110000110",
  35883=>"110110011",
  35884=>"101001111",
  35885=>"001010001",
  35886=>"100001011",
  35887=>"010110111",
  35888=>"111011001",
  35889=>"010011110",
  35890=>"000000000",
  35891=>"100111011",
  35892=>"111001000",
  35893=>"100000001",
  35894=>"100101010",
  35895=>"111111100",
  35896=>"000100110",
  35897=>"101001101",
  35898=>"001001110",
  35899=>"000011100",
  35900=>"010111000",
  35901=>"010001111",
  35902=>"011000101",
  35903=>"000110001",
  35904=>"111111000",
  35905=>"001001111",
  35906=>"000011010",
  35907=>"011010011",
  35908=>"010000001",
  35909=>"111101101",
  35910=>"000110010",
  35911=>"001001010",
  35912=>"010110000",
  35913=>"000111000",
  35914=>"110010011",
  35915=>"000000001",
  35916=>"000110100",
  35917=>"110111011",
  35918=>"110010111",
  35919=>"100001000",
  35920=>"101101000",
  35921=>"101010100",
  35922=>"000000001",
  35923=>"011101110",
  35924=>"011010000",
  35925=>"000010010",
  35926=>"001000011",
  35927=>"000000101",
  35928=>"010011101",
  35929=>"101001001",
  35930=>"100001010",
  35931=>"000000011",
  35932=>"111110000",
  35933=>"101100000",
  35934=>"111000000",
  35935=>"111001000",
  35936=>"100001111",
  35937=>"010111010",
  35938=>"010110111",
  35939=>"001111011",
  35940=>"111101101",
  35941=>"010010111",
  35942=>"001111001",
  35943=>"001011101",
  35944=>"010001101",
  35945=>"101011001",
  35946=>"000110001",
  35947=>"000101011",
  35948=>"010101111",
  35949=>"010011010",
  35950=>"100000101",
  35951=>"001111101",
  35952=>"100000000",
  35953=>"111000110",
  35954=>"101110001",
  35955=>"000110101",
  35956=>"000101100",
  35957=>"101010110",
  35958=>"001101101",
  35959=>"011100111",
  35960=>"101101101",
  35961=>"001000100",
  35962=>"101101101",
  35963=>"111000000",
  35964=>"100100101",
  35965=>"111010111",
  35966=>"001000101",
  35967=>"000000000",
  35968=>"111000101",
  35969=>"101010100",
  35970=>"001000001",
  35971=>"001011000",
  35972=>"011010100",
  35973=>"100000111",
  35974=>"001111110",
  35975=>"110100100",
  35976=>"000110101",
  35977=>"000000011",
  35978=>"111100000",
  35979=>"110001011",
  35980=>"101001110",
  35981=>"000001111",
  35982=>"101001101",
  35983=>"110001010",
  35984=>"001010010",
  35985=>"100100001",
  35986=>"010011101",
  35987=>"001000011",
  35988=>"000100110",
  35989=>"001010001",
  35990=>"001010111",
  35991=>"100000110",
  35992=>"011100000",
  35993=>"010101101",
  35994=>"000011000",
  35995=>"111111111",
  35996=>"100111011",
  35997=>"110000110",
  35998=>"110110000",
  35999=>"011110101",
  36000=>"101100110",
  36001=>"010001011",
  36002=>"100101000",
  36003=>"000011110",
  36004=>"111111011",
  36005=>"001011010",
  36006=>"111111010",
  36007=>"011000001",
  36008=>"111110000",
  36009=>"001110010",
  36010=>"000100011",
  36011=>"001001011",
  36012=>"001001010",
  36013=>"100001110",
  36014=>"100000110",
  36015=>"011101010",
  36016=>"000000101",
  36017=>"000110110",
  36018=>"111001000",
  36019=>"011000100",
  36020=>"101011100",
  36021=>"010010000",
  36022=>"100101110",
  36023=>"001001100",
  36024=>"101001000",
  36025=>"011101000",
  36026=>"000101011",
  36027=>"100000101",
  36028=>"001010100",
  36029=>"111011010",
  36030=>"100111100",
  36031=>"110010000",
  36032=>"001101101",
  36033=>"001001111",
  36034=>"110111111",
  36035=>"000000011",
  36036=>"001110100",
  36037=>"101110111",
  36038=>"111011110",
  36039=>"100100110",
  36040=>"111011100",
  36041=>"000011101",
  36042=>"110110100",
  36043=>"011110011",
  36044=>"110000000",
  36045=>"101001101",
  36046=>"000010001",
  36047=>"111101001",
  36048=>"110101011",
  36049=>"001110011",
  36050=>"000111000",
  36051=>"000011000",
  36052=>"010101110",
  36053=>"110101110",
  36054=>"000001101",
  36055=>"110010110",
  36056=>"000000100",
  36057=>"111100000",
  36058=>"100001101",
  36059=>"110111010",
  36060=>"001010000",
  36061=>"001011000",
  36062=>"101110000",
  36063=>"101010101",
  36064=>"111010110",
  36065=>"100111110",
  36066=>"011111111",
  36067=>"111010010",
  36068=>"010100000",
  36069=>"111111100",
  36070=>"100011001",
  36071=>"111100011",
  36072=>"001111110",
  36073=>"011001010",
  36074=>"011111011",
  36075=>"111100101",
  36076=>"111001000",
  36077=>"111011010",
  36078=>"111100101",
  36079=>"100101011",
  36080=>"010001110",
  36081=>"101101001",
  36082=>"111100101",
  36083=>"100010111",
  36084=>"000111101",
  36085=>"111011000",
  36086=>"000000011",
  36087=>"100011010",
  36088=>"000011101",
  36089=>"100100000",
  36090=>"000101000",
  36091=>"000100100",
  36092=>"001001010",
  36093=>"101001001",
  36094=>"010010100",
  36095=>"000100101",
  36096=>"111101101",
  36097=>"110011000",
  36098=>"001010010",
  36099=>"101011110",
  36100=>"000000010",
  36101=>"110001000",
  36102=>"001110011",
  36103=>"001010110",
  36104=>"111111011",
  36105=>"110010100",
  36106=>"000001100",
  36107=>"001111010",
  36108=>"010010010",
  36109=>"111101101",
  36110=>"110101100",
  36111=>"000100001",
  36112=>"001111011",
  36113=>"010010110",
  36114=>"001001111",
  36115=>"101100100",
  36116=>"100010110",
  36117=>"101110101",
  36118=>"010000001",
  36119=>"011000100",
  36120=>"111100101",
  36121=>"010011110",
  36122=>"010000100",
  36123=>"000001010",
  36124=>"110111101",
  36125=>"001101001",
  36126=>"110110100",
  36127=>"110100101",
  36128=>"101110001",
  36129=>"110101111",
  36130=>"011100011",
  36131=>"011110101",
  36132=>"110111001",
  36133=>"101110001",
  36134=>"101101100",
  36135=>"111011010",
  36136=>"111110001",
  36137=>"111110001",
  36138=>"111101001",
  36139=>"000000010",
  36140=>"000000000",
  36141=>"011011111",
  36142=>"110010001",
  36143=>"001110010",
  36144=>"010001101",
  36145=>"011011001",
  36146=>"101100011",
  36147=>"011010000",
  36148=>"011100100",
  36149=>"000000010",
  36150=>"111101010",
  36151=>"001001101",
  36152=>"000001000",
  36153=>"010000010",
  36154=>"111101000",
  36155=>"110100100",
  36156=>"100011001",
  36157=>"100110010",
  36158=>"100011011",
  36159=>"000000111",
  36160=>"100010101",
  36161=>"111011111",
  36162=>"011110011",
  36163=>"001011110",
  36164=>"001000100",
  36165=>"001101000",
  36166=>"100010000",
  36167=>"010111010",
  36168=>"011011001",
  36169=>"010011001",
  36170=>"110001010",
  36171=>"000000000",
  36172=>"111111110",
  36173=>"011011001",
  36174=>"000100011",
  36175=>"011010000",
  36176=>"111101101",
  36177=>"111011110",
  36178=>"110011000",
  36179=>"100011111",
  36180=>"100001111",
  36181=>"100100110",
  36182=>"100101000",
  36183=>"000110001",
  36184=>"110101000",
  36185=>"000000110",
  36186=>"101000100",
  36187=>"000000110",
  36188=>"101110111",
  36189=>"110001010",
  36190=>"110111100",
  36191=>"110000011",
  36192=>"001100010",
  36193=>"101110000",
  36194=>"100110100",
  36195=>"000111110",
  36196=>"110100100",
  36197=>"000100000",
  36198=>"000001101",
  36199=>"010111100",
  36200=>"100111011",
  36201=>"111110000",
  36202=>"000100111",
  36203=>"110101100",
  36204=>"001010100",
  36205=>"110011111",
  36206=>"101000010",
  36207=>"010110000",
  36208=>"011111000",
  36209=>"110100011",
  36210=>"001110011",
  36211=>"000110010",
  36212=>"100000011",
  36213=>"101101011",
  36214=>"100011101",
  36215=>"110010001",
  36216=>"110011001",
  36217=>"101101000",
  36218=>"111111111",
  36219=>"000111001",
  36220=>"001100110",
  36221=>"100000011",
  36222=>"100111111",
  36223=>"101001100",
  36224=>"111000010",
  36225=>"011000101",
  36226=>"011001111",
  36227=>"100100101",
  36228=>"100001110",
  36229=>"100110000",
  36230=>"010011110",
  36231=>"101001000",
  36232=>"000100010",
  36233=>"000110110",
  36234=>"101100101",
  36235=>"100110100",
  36236=>"000100000",
  36237=>"100101000",
  36238=>"111100100",
  36239=>"011010110",
  36240=>"001110110",
  36241=>"000100111",
  36242=>"100011001",
  36243=>"100101000",
  36244=>"010010110",
  36245=>"100111101",
  36246=>"001111010",
  36247=>"110000011",
  36248=>"111001111",
  36249=>"100000000",
  36250=>"110010110",
  36251=>"100111001",
  36252=>"010001000",
  36253=>"101001010",
  36254=>"000011111",
  36255=>"011110011",
  36256=>"000111110",
  36257=>"001010100",
  36258=>"011110110",
  36259=>"000100011",
  36260=>"101000000",
  36261=>"000000000",
  36262=>"111101000",
  36263=>"101101001",
  36264=>"000101011",
  36265=>"000110000",
  36266=>"000001111",
  36267=>"000000101",
  36268=>"100111100",
  36269=>"001001001",
  36270=>"101111100",
  36271=>"111111010",
  36272=>"101001100",
  36273=>"101010010",
  36274=>"101000110",
  36275=>"000101000",
  36276=>"100110100",
  36277=>"101010100",
  36278=>"111100010",
  36279=>"101011111",
  36280=>"011111111",
  36281=>"001110000",
  36282=>"100001111",
  36283=>"100011000",
  36284=>"011101010",
  36285=>"101000100",
  36286=>"010000010",
  36287=>"000101110",
  36288=>"110000111",
  36289=>"001001000",
  36290=>"110100010",
  36291=>"000011001",
  36292=>"100000010",
  36293=>"110111111",
  36294=>"011010010",
  36295=>"100000110",
  36296=>"111011011",
  36297=>"010011110",
  36298=>"100110000",
  36299=>"001101000",
  36300=>"101011010",
  36301=>"001000101",
  36302=>"100000101",
  36303=>"101100111",
  36304=>"100101110",
  36305=>"000011010",
  36306=>"110001100",
  36307=>"101010100",
  36308=>"111100011",
  36309=>"111010011",
  36310=>"010000011",
  36311=>"010101111",
  36312=>"110000100",
  36313=>"001001000",
  36314=>"010011000",
  36315=>"011101010",
  36316=>"110100101",
  36317=>"100101101",
  36318=>"110111111",
  36319=>"110110110",
  36320=>"001100110",
  36321=>"111000011",
  36322=>"000110000",
  36323=>"001110000",
  36324=>"101010100",
  36325=>"110100001",
  36326=>"100111010",
  36327=>"101111111",
  36328=>"100010001",
  36329=>"111110110",
  36330=>"011001001",
  36331=>"011000001",
  36332=>"110001011",
  36333=>"101111101",
  36334=>"110001000",
  36335=>"011111100",
  36336=>"101011010",
  36337=>"111101111",
  36338=>"001011000",
  36339=>"001000000",
  36340=>"001100110",
  36341=>"001110101",
  36342=>"010111000",
  36343=>"101101100",
  36344=>"101100001",
  36345=>"111011111",
  36346=>"111100001",
  36347=>"000001110",
  36348=>"100000011",
  36349=>"000110111",
  36350=>"111010010",
  36351=>"110011101",
  36352=>"110101111",
  36353=>"110100011",
  36354=>"011101010",
  36355=>"101100100",
  36356=>"000000011",
  36357=>"011011000",
  36358=>"111011101",
  36359=>"010101011",
  36360=>"010000111",
  36361=>"110101100",
  36362=>"000100001",
  36363=>"000010110",
  36364=>"010101000",
  36365=>"111000111",
  36366=>"101000011",
  36367=>"111011110",
  36368=>"010110111",
  36369=>"101001010",
  36370=>"000001011",
  36371=>"101010100",
  36372=>"000111001",
  36373=>"000010111",
  36374=>"110010110",
  36375=>"000111101",
  36376=>"111010101",
  36377=>"001111101",
  36378=>"010011100",
  36379=>"001100111",
  36380=>"101100000",
  36381=>"101000110",
  36382=>"001110010",
  36383=>"111110101",
  36384=>"110010001",
  36385=>"010000000",
  36386=>"001100110",
  36387=>"100100111",
  36388=>"011101011",
  36389=>"100111111",
  36390=>"001001110",
  36391=>"111011011",
  36392=>"100110101",
  36393=>"011011111",
  36394=>"101100010",
  36395=>"011110101",
  36396=>"001000100",
  36397=>"001110001",
  36398=>"100100110",
  36399=>"111011001",
  36400=>"110111111",
  36401=>"010100000",
  36402=>"100101001",
  36403=>"111101011",
  36404=>"111010000",
  36405=>"010001000",
  36406=>"101000010",
  36407=>"110011010",
  36408=>"010101111",
  36409=>"101011111",
  36410=>"100010001",
  36411=>"000111111",
  36412=>"010011010",
  36413=>"000000000",
  36414=>"110010001",
  36415=>"010000100",
  36416=>"111100000",
  36417=>"011110011",
  36418=>"000101110",
  36419=>"101000111",
  36420=>"110000111",
  36421=>"101111101",
  36422=>"110011110",
  36423=>"111011110",
  36424=>"000010011",
  36425=>"000110010",
  36426=>"110100101",
  36427=>"110100010",
  36428=>"111111111",
  36429=>"001100101",
  36430=>"101111111",
  36431=>"111010110",
  36432=>"100011100",
  36433=>"011111101",
  36434=>"011010101",
  36435=>"010001010",
  36436=>"010000000",
  36437=>"010000100",
  36438=>"000100001",
  36439=>"110000011",
  36440=>"101101011",
  36441=>"100100001",
  36442=>"000100000",
  36443=>"100000011",
  36444=>"110101100",
  36445=>"000010000",
  36446=>"011011100",
  36447=>"111101001",
  36448=>"100100000",
  36449=>"110000011",
  36450=>"101111011",
  36451=>"000001000",
  36452=>"100111001",
  36453=>"000010100",
  36454=>"111111000",
  36455=>"001101100",
  36456=>"010000000",
  36457=>"011010000",
  36458=>"100111000",
  36459=>"111000100",
  36460=>"001001000",
  36461=>"000101000",
  36462=>"011110110",
  36463=>"101011110",
  36464=>"000100000",
  36465=>"111000111",
  36466=>"001010011",
  36467=>"111111000",
  36468=>"111110100",
  36469=>"111111000",
  36470=>"100101001",
  36471=>"100110011",
  36472=>"001101000",
  36473=>"101000010",
  36474=>"001001111",
  36475=>"101010010",
  36476=>"101000100",
  36477=>"110000100",
  36478=>"110101011",
  36479=>"010101111",
  36480=>"110011111",
  36481=>"110011110",
  36482=>"001011110",
  36483=>"101001110",
  36484=>"001000000",
  36485=>"001000000",
  36486=>"101110101",
  36487=>"011001000",
  36488=>"001110100",
  36489=>"101101110",
  36490=>"101110010",
  36491=>"011000001",
  36492=>"011100000",
  36493=>"010111000",
  36494=>"110010110",
  36495=>"100111100",
  36496=>"110110001",
  36497=>"110011011",
  36498=>"000000101",
  36499=>"110110010",
  36500=>"000100001",
  36501=>"110001110",
  36502=>"100110011",
  36503=>"011010111",
  36504=>"101010100",
  36505=>"111100100",
  36506=>"011011101",
  36507=>"001011111",
  36508=>"111000001",
  36509=>"000101001",
  36510=>"000100101",
  36511=>"011011001",
  36512=>"101101110",
  36513=>"100100001",
  36514=>"111101101",
  36515=>"000110101",
  36516=>"101111000",
  36517=>"000010010",
  36518=>"000001001",
  36519=>"010000001",
  36520=>"011100010",
  36521=>"000100000",
  36522=>"001011010",
  36523=>"001010000",
  36524=>"001011000",
  36525=>"110001001",
  36526=>"101000101",
  36527=>"010100001",
  36528=>"010010010",
  36529=>"010000111",
  36530=>"110100010",
  36531=>"000100001",
  36532=>"001101100",
  36533=>"001110111",
  36534=>"110111010",
  36535=>"000010000",
  36536=>"101101001",
  36537=>"110010110",
  36538=>"010000100",
  36539=>"010001111",
  36540=>"101111110",
  36541=>"101001001",
  36542=>"100100010",
  36543=>"011101110",
  36544=>"110011010",
  36545=>"101010111",
  36546=>"100100101",
  36547=>"101010111",
  36548=>"000111010",
  36549=>"011100000",
  36550=>"100000000",
  36551=>"000000011",
  36552=>"111000011",
  36553=>"000010100",
  36554=>"001011010",
  36555=>"000000100",
  36556=>"010010000",
  36557=>"110011111",
  36558=>"101011110",
  36559=>"111010101",
  36560=>"101101000",
  36561=>"100010101",
  36562=>"101100000",
  36563=>"010010000",
  36564=>"111001111",
  36565=>"100100010",
  36566=>"000110111",
  36567=>"000111010",
  36568=>"101010000",
  36569=>"010100011",
  36570=>"001001011",
  36571=>"011011001",
  36572=>"000101111",
  36573=>"111101111",
  36574=>"101010100",
  36575=>"000011000",
  36576=>"010010000",
  36577=>"000010111",
  36578=>"011100101",
  36579=>"111011010",
  36580=>"101110111",
  36581=>"111101111",
  36582=>"100000000",
  36583=>"010001010",
  36584=>"000010001",
  36585=>"101110111",
  36586=>"110001010",
  36587=>"111000110",
  36588=>"010100000",
  36589=>"000111111",
  36590=>"101100100",
  36591=>"000011111",
  36592=>"000100100",
  36593=>"100110010",
  36594=>"001100111",
  36595=>"111111011",
  36596=>"100100010",
  36597=>"011100101",
  36598=>"101110011",
  36599=>"111101001",
  36600=>"011101011",
  36601=>"101000010",
  36602=>"001001101",
  36603=>"100111001",
  36604=>"110001011",
  36605=>"011111000",
  36606=>"010000011",
  36607=>"110011100",
  36608=>"111100010",
  36609=>"010000010",
  36610=>"010110100",
  36611=>"000101001",
  36612=>"110010011",
  36613=>"101001110",
  36614=>"001001010",
  36615=>"101101011",
  36616=>"101010110",
  36617=>"001111011",
  36618=>"111010101",
  36619=>"000010101",
  36620=>"011000011",
  36621=>"111101100",
  36622=>"010101111",
  36623=>"011011111",
  36624=>"001010111",
  36625=>"001001100",
  36626=>"011011000",
  36627=>"011101001",
  36628=>"100001011",
  36629=>"001011001",
  36630=>"011011011",
  36631=>"100110001",
  36632=>"100101100",
  36633=>"001000011",
  36634=>"110000100",
  36635=>"110101110",
  36636=>"010101010",
  36637=>"010011110",
  36638=>"100000000",
  36639=>"011110110",
  36640=>"110001001",
  36641=>"111010111",
  36642=>"101011101",
  36643=>"100011010",
  36644=>"010010110",
  36645=>"001100110",
  36646=>"011011010",
  36647=>"011011010",
  36648=>"110111110",
  36649=>"000011100",
  36650=>"001001000",
  36651=>"010011001",
  36652=>"110011001",
  36653=>"001001010",
  36654=>"100000000",
  36655=>"010110000",
  36656=>"100000010",
  36657=>"000011101",
  36658=>"010100010",
  36659=>"100001010",
  36660=>"111100100",
  36661=>"010000100",
  36662=>"110000100",
  36663=>"000001000",
  36664=>"010100100",
  36665=>"111110101",
  36666=>"010100111",
  36667=>"011101011",
  36668=>"010100100",
  36669=>"000101010",
  36670=>"000100000",
  36671=>"010111110",
  36672=>"001000001",
  36673=>"001010100",
  36674=>"011110011",
  36675=>"011110011",
  36676=>"001001100",
  36677=>"111101000",
  36678=>"101000010",
  36679=>"000110010",
  36680=>"000010010",
  36681=>"111000111",
  36682=>"011111100",
  36683=>"100010100",
  36684=>"011101110",
  36685=>"110101010",
  36686=>"011110110",
  36687=>"101010010",
  36688=>"000100000",
  36689=>"000111100",
  36690=>"101000100",
  36691=>"010010101",
  36692=>"010111110",
  36693=>"110111010",
  36694=>"111110100",
  36695=>"000011101",
  36696=>"010000011",
  36697=>"101110110",
  36698=>"111011010",
  36699=>"010010010",
  36700=>"000011110",
  36701=>"011000101",
  36702=>"101111110",
  36703=>"000000001",
  36704=>"011000100",
  36705=>"001010110",
  36706=>"001010000",
  36707=>"111111001",
  36708=>"110100100",
  36709=>"101011000",
  36710=>"010001110",
  36711=>"101110011",
  36712=>"001001000",
  36713=>"001001000",
  36714=>"000110101",
  36715=>"011111011",
  36716=>"101001101",
  36717=>"010010001",
  36718=>"000000100",
  36719=>"001001101",
  36720=>"110101101",
  36721=>"010011110",
  36722=>"110111010",
  36723=>"010010001",
  36724=>"010101001",
  36725=>"001010110",
  36726=>"110101000",
  36727=>"000001111",
  36728=>"000010101",
  36729=>"001011001",
  36730=>"101010101",
  36731=>"011100101",
  36732=>"000100000",
  36733=>"100101111",
  36734=>"000111110",
  36735=>"110110111",
  36736=>"111110001",
  36737=>"011100101",
  36738=>"111010101",
  36739=>"000010110",
  36740=>"010010100",
  36741=>"100111011",
  36742=>"010101000",
  36743=>"110101101",
  36744=>"110100000",
  36745=>"000101101",
  36746=>"111101100",
  36747=>"100000001",
  36748=>"101011000",
  36749=>"001110100",
  36750=>"001111100",
  36751=>"110101010",
  36752=>"110100011",
  36753=>"110100110",
  36754=>"100110110",
  36755=>"000010110",
  36756=>"101111111",
  36757=>"100011100",
  36758=>"110000010",
  36759=>"011000010",
  36760=>"111001110",
  36761=>"000100111",
  36762=>"110111100",
  36763=>"110101010",
  36764=>"001010000",
  36765=>"001111010",
  36766=>"111000001",
  36767=>"111111101",
  36768=>"010100101",
  36769=>"001000010",
  36770=>"000100001",
  36771=>"001000011",
  36772=>"100110001",
  36773=>"100001100",
  36774=>"100010000",
  36775=>"000100111",
  36776=>"001011010",
  36777=>"001000110",
  36778=>"001101111",
  36779=>"011011101",
  36780=>"101010000",
  36781=>"101101001",
  36782=>"111011110",
  36783=>"110011000",
  36784=>"001001010",
  36785=>"111111111",
  36786=>"100001101",
  36787=>"001000110",
  36788=>"100101110",
  36789=>"100101011",
  36790=>"000110111",
  36791=>"111101001",
  36792=>"101110010",
  36793=>"110010000",
  36794=>"110111010",
  36795=>"010000100",
  36796=>"011110100",
  36797=>"000000010",
  36798=>"001010110",
  36799=>"011010100",
  36800=>"000001110",
  36801=>"001001111",
  36802=>"000101101",
  36803=>"100010101",
  36804=>"100110111",
  36805=>"111011011",
  36806=>"000101000",
  36807=>"110010101",
  36808=>"011000100",
  36809=>"111110110",
  36810=>"110100011",
  36811=>"100101010",
  36812=>"000000011",
  36813=>"000000100",
  36814=>"000110100",
  36815=>"110101001",
  36816=>"000010100",
  36817=>"110010010",
  36818=>"010011000",
  36819=>"010111011",
  36820=>"001110100",
  36821=>"100010001",
  36822=>"101010010",
  36823=>"000111000",
  36824=>"101010000",
  36825=>"000101101",
  36826=>"010000100",
  36827=>"011001001",
  36828=>"011000010",
  36829=>"011101010",
  36830=>"100101000",
  36831=>"001110110",
  36832=>"101110010",
  36833=>"011110111",
  36834=>"111110101",
  36835=>"001110100",
  36836=>"010000101",
  36837=>"000111111",
  36838=>"101101101",
  36839=>"000101101",
  36840=>"000100010",
  36841=>"010010011",
  36842=>"001111100",
  36843=>"100100001",
  36844=>"111010011",
  36845=>"101100101",
  36846=>"100110111",
  36847=>"010011100",
  36848=>"100100001",
  36849=>"111001001",
  36850=>"000000110",
  36851=>"000101111",
  36852=>"001011010",
  36853=>"001111000",
  36854=>"100111101",
  36855=>"011001011",
  36856=>"011011011",
  36857=>"100010011",
  36858=>"011101000",
  36859=>"111010000",
  36860=>"000100010",
  36861=>"001001111",
  36862=>"111111010",
  36863=>"010110111",
  36864=>"010001001",
  36865=>"101011001",
  36866=>"100011011",
  36867=>"111011011",
  36868=>"100110101",
  36869=>"111010010",
  36870=>"101111100",
  36871=>"011001001",
  36872=>"001101111",
  36873=>"100100110",
  36874=>"001010001",
  36875=>"000100101",
  36876=>"011101000",
  36877=>"111100000",
  36878=>"000010111",
  36879=>"001101101",
  36880=>"001011011",
  36881=>"100111111",
  36882=>"000000100",
  36883=>"011010001",
  36884=>"101101111",
  36885=>"110000101",
  36886=>"101001111",
  36887=>"101101001",
  36888=>"000010000",
  36889=>"111111111",
  36890=>"000111100",
  36891=>"011101011",
  36892=>"010100000",
  36893=>"111110110",
  36894=>"111001101",
  36895=>"000011100",
  36896=>"010100010",
  36897=>"111111001",
  36898=>"110000000",
  36899=>"001000010",
  36900=>"000010001",
  36901=>"101101110",
  36902=>"000101111",
  36903=>"111001100",
  36904=>"101001000",
  36905=>"001011100",
  36906=>"000010100",
  36907=>"100010101",
  36908=>"111010100",
  36909=>"111111001",
  36910=>"000110001",
  36911=>"010110110",
  36912=>"010001101",
  36913=>"110110101",
  36914=>"111101001",
  36915=>"001000111",
  36916=>"110111111",
  36917=>"100111110",
  36918=>"010010000",
  36919=>"000001110",
  36920=>"101100110",
  36921=>"101110100",
  36922=>"001111111",
  36923=>"100100110",
  36924=>"111100000",
  36925=>"110111111",
  36926=>"000010100",
  36927=>"111010001",
  36928=>"011100110",
  36929=>"100111110",
  36930=>"100000010",
  36931=>"011001011",
  36932=>"111000010",
  36933=>"110011111",
  36934=>"010100010",
  36935=>"110001010",
  36936=>"000101101",
  36937=>"011000111",
  36938=>"111110101",
  36939=>"100111111",
  36940=>"100110010",
  36941=>"000001101",
  36942=>"001000111",
  36943=>"010010000",
  36944=>"100011000",
  36945=>"001001001",
  36946=>"001111000",
  36947=>"111110010",
  36948=>"110111000",
  36949=>"011110111",
  36950=>"000111000",
  36951=>"100101000",
  36952=>"111110111",
  36953=>"100111110",
  36954=>"101000000",
  36955=>"001011011",
  36956=>"100000101",
  36957=>"001010000",
  36958=>"010111100",
  36959=>"000101010",
  36960=>"000010100",
  36961=>"101000000",
  36962=>"100101000",
  36963=>"101110011",
  36964=>"000000111",
  36965=>"011000111",
  36966=>"101111010",
  36967=>"011110111",
  36968=>"111000011",
  36969=>"000111110",
  36970=>"101111111",
  36971=>"000000100",
  36972=>"111100000",
  36973=>"111001011",
  36974=>"000011101",
  36975=>"110110110",
  36976=>"111101101",
  36977=>"010111000",
  36978=>"111100100",
  36979=>"000010110",
  36980=>"011110011",
  36981=>"111100100",
  36982=>"001000000",
  36983=>"100101110",
  36984=>"100111111",
  36985=>"011011111",
  36986=>"100010011",
  36987=>"101001001",
  36988=>"110001100",
  36989=>"010011000",
  36990=>"111111011",
  36991=>"001110011",
  36992=>"110011111",
  36993=>"001110101",
  36994=>"111011101",
  36995=>"001000011",
  36996=>"001010010",
  36997=>"110000101",
  36998=>"000000111",
  36999=>"010001001",
  37000=>"001010111",
  37001=>"101111101",
  37002=>"010100110",
  37003=>"000110111",
  37004=>"100101010",
  37005=>"001111111",
  37006=>"111000001",
  37007=>"010110000",
  37008=>"100011000",
  37009=>"101101000",
  37010=>"100011110",
  37011=>"111011011",
  37012=>"101000000",
  37013=>"111101010",
  37014=>"111001100",
  37015=>"001101101",
  37016=>"110110111",
  37017=>"001100100",
  37018=>"000111111",
  37019=>"010001100",
  37020=>"111100001",
  37021=>"000111111",
  37022=>"110000111",
  37023=>"000110100",
  37024=>"111111100",
  37025=>"101111111",
  37026=>"011011011",
  37027=>"001100010",
  37028=>"111100111",
  37029=>"011010011",
  37030=>"001100110",
  37031=>"010111111",
  37032=>"101000000",
  37033=>"010010111",
  37034=>"001101110",
  37035=>"101111000",
  37036=>"100010010",
  37037=>"100000001",
  37038=>"010100000",
  37039=>"000000000",
  37040=>"111100011",
  37041=>"001111100",
  37042=>"101011111",
  37043=>"000001111",
  37044=>"101100101",
  37045=>"111110011",
  37046=>"000101001",
  37047=>"101101110",
  37048=>"111110011",
  37049=>"101001101",
  37050=>"000010111",
  37051=>"100011101",
  37052=>"001111110",
  37053=>"000110100",
  37054=>"001011100",
  37055=>"110111111",
  37056=>"010111110",
  37057=>"000000010",
  37058=>"110110001",
  37059=>"101011100",
  37060=>"111010000",
  37061=>"000111111",
  37062=>"110110101",
  37063=>"010110101",
  37064=>"110001011",
  37065=>"011111101",
  37066=>"001000001",
  37067=>"011010010",
  37068=>"110101100",
  37069=>"001101000",
  37070=>"011010010",
  37071=>"101001010",
  37072=>"000100100",
  37073=>"101000001",
  37074=>"101111101",
  37075=>"111001001",
  37076=>"111010111",
  37077=>"001111011",
  37078=>"000101000",
  37079=>"010110111",
  37080=>"111011110",
  37081=>"101100111",
  37082=>"100111111",
  37083=>"100100000",
  37084=>"101011111",
  37085=>"001000011",
  37086=>"011111001",
  37087=>"000000001",
  37088=>"101111110",
  37089=>"101111100",
  37090=>"101110100",
  37091=>"101100011",
  37092=>"001011000",
  37093=>"100101110",
  37094=>"100011111",
  37095=>"110111001",
  37096=>"000010111",
  37097=>"000111001",
  37098=>"110110111",
  37099=>"111010101",
  37100=>"010000010",
  37101=>"010110001",
  37102=>"001011110",
  37103=>"010101001",
  37104=>"111100100",
  37105=>"100110110",
  37106=>"100100111",
  37107=>"111001110",
  37108=>"010011100",
  37109=>"110100010",
  37110=>"001010100",
  37111=>"100101010",
  37112=>"101110110",
  37113=>"110000000",
  37114=>"101000101",
  37115=>"000111011",
  37116=>"110100011",
  37117=>"110001110",
  37118=>"010001111",
  37119=>"001100000",
  37120=>"010001001",
  37121=>"011000000",
  37122=>"110000001",
  37123=>"000111111",
  37124=>"101111001",
  37125=>"011111100",
  37126=>"000111100",
  37127=>"101000010",
  37128=>"101011000",
  37129=>"001000011",
  37130=>"111101000",
  37131=>"111001110",
  37132=>"000001011",
  37133=>"111111111",
  37134=>"101011000",
  37135=>"110100011",
  37136=>"110100001",
  37137=>"010010101",
  37138=>"011111110",
  37139=>"100100111",
  37140=>"101001000",
  37141=>"001001111",
  37142=>"000000001",
  37143=>"111011000",
  37144=>"111001100",
  37145=>"111000111",
  37146=>"011111111",
  37147=>"011010011",
  37148=>"100100111",
  37149=>"000100111",
  37150=>"111000010",
  37151=>"000010001",
  37152=>"000100001",
  37153=>"000010111",
  37154=>"111001110",
  37155=>"001011110",
  37156=>"110100000",
  37157=>"111010111",
  37158=>"010000000",
  37159=>"111011011",
  37160=>"110001011",
  37161=>"010000110",
  37162=>"011110010",
  37163=>"001100001",
  37164=>"111101101",
  37165=>"001100110",
  37166=>"001000010",
  37167=>"011010010",
  37168=>"111101010",
  37169=>"100110100",
  37170=>"001110111",
  37171=>"001101011",
  37172=>"001000000",
  37173=>"010001100",
  37174=>"100000110",
  37175=>"010110100",
  37176=>"011011101",
  37177=>"110010011",
  37178=>"011101110",
  37179=>"111011101",
  37180=>"011111110",
  37181=>"000111011",
  37182=>"101001000",
  37183=>"010001100",
  37184=>"101110110",
  37185=>"111110100",
  37186=>"001010101",
  37187=>"101110101",
  37188=>"000001111",
  37189=>"000110100",
  37190=>"010000100",
  37191=>"001101001",
  37192=>"101110111",
  37193=>"111101011",
  37194=>"101100010",
  37195=>"011000101",
  37196=>"101111011",
  37197=>"010110111",
  37198=>"010001000",
  37199=>"001011100",
  37200=>"010010001",
  37201=>"111100000",
  37202=>"011011101",
  37203=>"101010010",
  37204=>"001011100",
  37205=>"001100110",
  37206=>"100100001",
  37207=>"001110011",
  37208=>"101110111",
  37209=>"110001011",
  37210=>"110101010",
  37211=>"111010111",
  37212=>"111110110",
  37213=>"100110101",
  37214=>"010110101",
  37215=>"010010101",
  37216=>"101011001",
  37217=>"100011111",
  37218=>"111011011",
  37219=>"000000100",
  37220=>"111110011",
  37221=>"110101100",
  37222=>"101000000",
  37223=>"000011010",
  37224=>"011010000",
  37225=>"110001100",
  37226=>"111100011",
  37227=>"011111011",
  37228=>"111110111",
  37229=>"000101101",
  37230=>"011010101",
  37231=>"000110111",
  37232=>"001111001",
  37233=>"110100011",
  37234=>"100011011",
  37235=>"000000000",
  37236=>"100100011",
  37237=>"000011110",
  37238=>"000110000",
  37239=>"101110010",
  37240=>"010110110",
  37241=>"001000101",
  37242=>"001000101",
  37243=>"100010001",
  37244=>"101111101",
  37245=>"011110110",
  37246=>"110111010",
  37247=>"001001100",
  37248=>"000101111",
  37249=>"110101000",
  37250=>"110000000",
  37251=>"001011011",
  37252=>"011101101",
  37253=>"100001100",
  37254=>"110101000",
  37255=>"010001111",
  37256=>"011010110",
  37257=>"000000100",
  37258=>"001011111",
  37259=>"011110101",
  37260=>"100111000",
  37261=>"110011100",
  37262=>"110001101",
  37263=>"111000000",
  37264=>"010111111",
  37265=>"010001010",
  37266=>"000111110",
  37267=>"111011001",
  37268=>"111010001",
  37269=>"000010001",
  37270=>"001110001",
  37271=>"001100010",
  37272=>"110011010",
  37273=>"101111111",
  37274=>"101110010",
  37275=>"101011000",
  37276=>"010110111",
  37277=>"010111111",
  37278=>"111111001",
  37279=>"010000010",
  37280=>"100000101",
  37281=>"000100010",
  37282=>"000100110",
  37283=>"100111100",
  37284=>"011000100",
  37285=>"100001000",
  37286=>"001110111",
  37287=>"010001001",
  37288=>"101100000",
  37289=>"111101010",
  37290=>"001110000",
  37291=>"011001111",
  37292=>"010111001",
  37293=>"111010100",
  37294=>"010001000",
  37295=>"101101110",
  37296=>"011011010",
  37297=>"000001111",
  37298=>"111110100",
  37299=>"111101011",
  37300=>"011001111",
  37301=>"011110111",
  37302=>"000010011",
  37303=>"100100011",
  37304=>"101100000",
  37305=>"000001011",
  37306=>"010011001",
  37307=>"111011100",
  37308=>"000011100",
  37309=>"111001111",
  37310=>"000011100",
  37311=>"110101001",
  37312=>"100000111",
  37313=>"110010011",
  37314=>"010001110",
  37315=>"110011111",
  37316=>"111011001",
  37317=>"010011100",
  37318=>"111101011",
  37319=>"101101111",
  37320=>"001100101",
  37321=>"111111111",
  37322=>"011010111",
  37323=>"000100000",
  37324=>"010011101",
  37325=>"110001000",
  37326=>"101011100",
  37327=>"010010011",
  37328=>"111000110",
  37329=>"001110101",
  37330=>"110101001",
  37331=>"011111101",
  37332=>"111110010",
  37333=>"010000101",
  37334=>"001101000",
  37335=>"110111101",
  37336=>"110100011",
  37337=>"000100001",
  37338=>"010011000",
  37339=>"101011111",
  37340=>"111001111",
  37341=>"000000010",
  37342=>"011101111",
  37343=>"010010110",
  37344=>"011000101",
  37345=>"101010101",
  37346=>"001010101",
  37347=>"111110110",
  37348=>"111110011",
  37349=>"101011100",
  37350=>"010100100",
  37351=>"101000011",
  37352=>"010011110",
  37353=>"010111010",
  37354=>"001001011",
  37355=>"110110110",
  37356=>"001101011",
  37357=>"000111011",
  37358=>"110101001",
  37359=>"101111111",
  37360=>"010110101",
  37361=>"000100001",
  37362=>"001111111",
  37363=>"011101111",
  37364=>"010111011",
  37365=>"011010011",
  37366=>"000110000",
  37367=>"100111111",
  37368=>"010001101",
  37369=>"010010001",
  37370=>"010000111",
  37371=>"000011001",
  37372=>"000111011",
  37373=>"001011001",
  37374=>"011000000",
  37375=>"010001101",
  37376=>"100100100",
  37377=>"110110101",
  37378=>"001001011",
  37379=>"000110011",
  37380=>"100101011",
  37381=>"110001010",
  37382=>"101100101",
  37383=>"000111001",
  37384=>"011011010",
  37385=>"101101110",
  37386=>"110110111",
  37387=>"110111110",
  37388=>"001011111",
  37389=>"111111101",
  37390=>"111111100",
  37391=>"000101101",
  37392=>"000111010",
  37393=>"100000010",
  37394=>"001111001",
  37395=>"100011101",
  37396=>"110101011",
  37397=>"101001011",
  37398=>"111111000",
  37399=>"110011100",
  37400=>"010110110",
  37401=>"000000101",
  37402=>"101011111",
  37403=>"000111110",
  37404=>"110000011",
  37405=>"001000001",
  37406=>"110011000",
  37407=>"011001110",
  37408=>"001101100",
  37409=>"110101111",
  37410=>"110100111",
  37411=>"100101101",
  37412=>"110111101",
  37413=>"101111111",
  37414=>"100111010",
  37415=>"100000111",
  37416=>"010010101",
  37417=>"000101011",
  37418=>"001011100",
  37419=>"111111110",
  37420=>"101110010",
  37421=>"111101100",
  37422=>"100101000",
  37423=>"000001001",
  37424=>"000110000",
  37425=>"110101001",
  37426=>"110011110",
  37427=>"000100000",
  37428=>"010011101",
  37429=>"000001100",
  37430=>"110101100",
  37431=>"001000111",
  37432=>"001110000",
  37433=>"001011111",
  37434=>"110110101",
  37435=>"100110111",
  37436=>"110010100",
  37437=>"101110110",
  37438=>"010001101",
  37439=>"100100110",
  37440=>"010001011",
  37441=>"110100001",
  37442=>"011111111",
  37443=>"101000111",
  37444=>"011010110",
  37445=>"111111010",
  37446=>"100000011",
  37447=>"000001001",
  37448=>"000100010",
  37449=>"101110001",
  37450=>"110000101",
  37451=>"010101011",
  37452=>"111111111",
  37453=>"110111110",
  37454=>"010101111",
  37455=>"100110101",
  37456=>"101011010",
  37457=>"000010100",
  37458=>"100010010",
  37459=>"111001101",
  37460=>"010011010",
  37461=>"100101110",
  37462=>"010101000",
  37463=>"010110001",
  37464=>"111010111",
  37465=>"101001000",
  37466=>"000010110",
  37467=>"110111010",
  37468=>"001011101",
  37469=>"000011111",
  37470=>"111101110",
  37471=>"110010101",
  37472=>"010100001",
  37473=>"001110111",
  37474=>"011110110",
  37475=>"100110111",
  37476=>"001001011",
  37477=>"111011010",
  37478=>"111100001",
  37479=>"101001111",
  37480=>"111110110",
  37481=>"001100101",
  37482=>"100100000",
  37483=>"101100110",
  37484=>"100011001",
  37485=>"111000011",
  37486=>"100101001",
  37487=>"110100100",
  37488=>"110011010",
  37489=>"101110000",
  37490=>"110111000",
  37491=>"100010110",
  37492=>"000010011",
  37493=>"110111100",
  37494=>"111010111",
  37495=>"101000001",
  37496=>"110001011",
  37497=>"011001001",
  37498=>"110010011",
  37499=>"111001101",
  37500=>"110110000",
  37501=>"001100111",
  37502=>"010100001",
  37503=>"010101000",
  37504=>"011110110",
  37505=>"101000111",
  37506=>"001111110",
  37507=>"110101000",
  37508=>"001101010",
  37509=>"110111100",
  37510=>"100111110",
  37511=>"000111000",
  37512=>"000001001",
  37513=>"100011001",
  37514=>"010010101",
  37515=>"111110111",
  37516=>"111011111",
  37517=>"011110100",
  37518=>"111100100",
  37519=>"001011100",
  37520=>"110111011",
  37521=>"101100011",
  37522=>"101111111",
  37523=>"110111101",
  37524=>"111011101",
  37525=>"100011010",
  37526=>"010001010",
  37527=>"011101011",
  37528=>"100100010",
  37529=>"100001001",
  37530=>"001110101",
  37531=>"010110100",
  37532=>"000010111",
  37533=>"001110011",
  37534=>"100110100",
  37535=>"001101111",
  37536=>"001100111",
  37537=>"000001010",
  37538=>"101011100",
  37539=>"111010010",
  37540=>"000011111",
  37541=>"001010111",
  37542=>"111011011",
  37543=>"000000011",
  37544=>"111100101",
  37545=>"111101001",
  37546=>"101000010",
  37547=>"101101011",
  37548=>"000011101",
  37549=>"100101110",
  37550=>"010100100",
  37551=>"000011001",
  37552=>"001111000",
  37553=>"111001010",
  37554=>"011110011",
  37555=>"100000101",
  37556=>"101100100",
  37557=>"110101010",
  37558=>"110110101",
  37559=>"111000001",
  37560=>"100011011",
  37561=>"101010100",
  37562=>"000010001",
  37563=>"010000000",
  37564=>"011011001",
  37565=>"100110010",
  37566=>"010110111",
  37567=>"000010101",
  37568=>"100110111",
  37569=>"110110111",
  37570=>"101110101",
  37571=>"100100100",
  37572=>"001111011",
  37573=>"000001010",
  37574=>"111000100",
  37575=>"111011011",
  37576=>"110001101",
  37577=>"110101110",
  37578=>"100100100",
  37579=>"001011111",
  37580=>"001011111",
  37581=>"111101101",
  37582=>"011000001",
  37583=>"000111001",
  37584=>"111001111",
  37585=>"010111100",
  37586=>"100111001",
  37587=>"101101101",
  37588=>"100100101",
  37589=>"111110111",
  37590=>"110111000",
  37591=>"101010001",
  37592=>"011001011",
  37593=>"010010101",
  37594=>"101100001",
  37595=>"111001111",
  37596=>"101001010",
  37597=>"000001101",
  37598=>"000100010",
  37599=>"100110111",
  37600=>"001011101",
  37601=>"000011011",
  37602=>"101001111",
  37603=>"100101110",
  37604=>"001011000",
  37605=>"000100000",
  37606=>"010111001",
  37607=>"001101011",
  37608=>"001101100",
  37609=>"010000110",
  37610=>"011011111",
  37611=>"010000110",
  37612=>"011010100",
  37613=>"110011000",
  37614=>"011101111",
  37615=>"101000011",
  37616=>"011111111",
  37617=>"110010000",
  37618=>"101100011",
  37619=>"011111100",
  37620=>"011111011",
  37621=>"111010000",
  37622=>"111010010",
  37623=>"111111110",
  37624=>"011110111",
  37625=>"110011101",
  37626=>"110111000",
  37627=>"100101111",
  37628=>"111110110",
  37629=>"111110011",
  37630=>"110010011",
  37631=>"000110100",
  37632=>"100111010",
  37633=>"110111011",
  37634=>"001010101",
  37635=>"111010001",
  37636=>"111011010",
  37637=>"011101000",
  37638=>"110011010",
  37639=>"010011100",
  37640=>"110001101",
  37641=>"010001100",
  37642=>"001101010",
  37643=>"011101111",
  37644=>"000001011",
  37645=>"110111110",
  37646=>"000001010",
  37647=>"011001010",
  37648=>"101100010",
  37649=>"000111011",
  37650=>"001001101",
  37651=>"110110011",
  37652=>"111010001",
  37653=>"111111001",
  37654=>"010001010",
  37655=>"101001000",
  37656=>"001001010",
  37657=>"110100010",
  37658=>"111011001",
  37659=>"111010111",
  37660=>"100100010",
  37661=>"010110100",
  37662=>"001000000",
  37663=>"111011011",
  37664=>"011111001",
  37665=>"110101011",
  37666=>"110001001",
  37667=>"000011110",
  37668=>"011111001",
  37669=>"101111101",
  37670=>"100010111",
  37671=>"001110000",
  37672=>"100110101",
  37673=>"100011001",
  37674=>"000010100",
  37675=>"011010101",
  37676=>"111001111",
  37677=>"111100110",
  37678=>"001111010",
  37679=>"000010001",
  37680=>"000100100",
  37681=>"011000011",
  37682=>"111111111",
  37683=>"111001110",
  37684=>"111010001",
  37685=>"100010101",
  37686=>"101000010",
  37687=>"010000111",
  37688=>"001111000",
  37689=>"000101010",
  37690=>"111100010",
  37691=>"001011011",
  37692=>"011111000",
  37693=>"000000000",
  37694=>"100111101",
  37695=>"110011001",
  37696=>"101000110",
  37697=>"100011011",
  37698=>"001110100",
  37699=>"000111000",
  37700=>"011110001",
  37701=>"010111101",
  37702=>"101001001",
  37703=>"000100101",
  37704=>"110110011",
  37705=>"010101000",
  37706=>"011011001",
  37707=>"000011111",
  37708=>"110111010",
  37709=>"101011110",
  37710=>"010010010",
  37711=>"001111010",
  37712=>"000001011",
  37713=>"111001111",
  37714=>"111011111",
  37715=>"110001110",
  37716=>"010111001",
  37717=>"001101011",
  37718=>"000100000",
  37719=>"011111111",
  37720=>"001110101",
  37721=>"110011111",
  37722=>"101011101",
  37723=>"101100001",
  37724=>"101001011",
  37725=>"101111100",
  37726=>"000011000",
  37727=>"011101110",
  37728=>"111111011",
  37729=>"011011011",
  37730=>"000101010",
  37731=>"000000101",
  37732=>"111010101",
  37733=>"001001011",
  37734=>"001010101",
  37735=>"110101011",
  37736=>"000011111",
  37737=>"111111001",
  37738=>"011111101",
  37739=>"110110000",
  37740=>"111001001",
  37741=>"011110111",
  37742=>"010001000",
  37743=>"100100110",
  37744=>"000101000",
  37745=>"110111110",
  37746=>"000101011",
  37747=>"111111111",
  37748=>"100101011",
  37749=>"111101011",
  37750=>"001010100",
  37751=>"101010010",
  37752=>"110011101",
  37753=>"011001000",
  37754=>"101110101",
  37755=>"001111100",
  37756=>"011111111",
  37757=>"111000011",
  37758=>"011001111",
  37759=>"010000010",
  37760=>"011001011",
  37761=>"011100100",
  37762=>"100110100",
  37763=>"000011010",
  37764=>"111101011",
  37765=>"111100011",
  37766=>"001110011",
  37767=>"101011001",
  37768=>"111000001",
  37769=>"111001011",
  37770=>"011011110",
  37771=>"001010100",
  37772=>"111000100",
  37773=>"100000010",
  37774=>"100010110",
  37775=>"000100100",
  37776=>"001100001",
  37777=>"110100101",
  37778=>"001011001",
  37779=>"100001101",
  37780=>"100011000",
  37781=>"000001000",
  37782=>"000010010",
  37783=>"010001110",
  37784=>"011001100",
  37785=>"001001011",
  37786=>"101011111",
  37787=>"101010101",
  37788=>"101110010",
  37789=>"010010110",
  37790=>"000101001",
  37791=>"110100000",
  37792=>"101111111",
  37793=>"011111111",
  37794=>"101011100",
  37795=>"110011110",
  37796=>"100011011",
  37797=>"100100100",
  37798=>"010011111",
  37799=>"011010110",
  37800=>"010111011",
  37801=>"101100111",
  37802=>"101000111",
  37803=>"011011101",
  37804=>"010000111",
  37805=>"000001110",
  37806=>"011110111",
  37807=>"100001101",
  37808=>"100010100",
  37809=>"101100100",
  37810=>"100111101",
  37811=>"110111110",
  37812=>"011000000",
  37813=>"111010010",
  37814=>"110110101",
  37815=>"001101011",
  37816=>"001110001",
  37817=>"101100010",
  37818=>"110101011",
  37819=>"011001111",
  37820=>"011101111",
  37821=>"001010100",
  37822=>"010000100",
  37823=>"010011110",
  37824=>"011110000",
  37825=>"110001011",
  37826=>"110111001",
  37827=>"011000000",
  37828=>"010000100",
  37829=>"110101101",
  37830=>"011011011",
  37831=>"110101011",
  37832=>"101110001",
  37833=>"111001100",
  37834=>"011000011",
  37835=>"000100000",
  37836=>"100010001",
  37837=>"110001001",
  37838=>"011111110",
  37839=>"000111001",
  37840=>"001100111",
  37841=>"001001000",
  37842=>"101011111",
  37843=>"101111101",
  37844=>"001011100",
  37845=>"000101000",
  37846=>"000010110",
  37847=>"010101100",
  37848=>"000111001",
  37849=>"111000001",
  37850=>"001000000",
  37851=>"111011001",
  37852=>"100001001",
  37853=>"110010101",
  37854=>"100010101",
  37855=>"101100111",
  37856=>"010001100",
  37857=>"111011001",
  37858=>"001110000",
  37859=>"111001111",
  37860=>"000110011",
  37861=>"100110110",
  37862=>"101110101",
  37863=>"010010011",
  37864=>"111110111",
  37865=>"010010110",
  37866=>"100011111",
  37867=>"100110110",
  37868=>"111111000",
  37869=>"101110110",
  37870=>"100101111",
  37871=>"110101101",
  37872=>"101010101",
  37873=>"101000100",
  37874=>"110011110",
  37875=>"100001000",
  37876=>"001010111",
  37877=>"011101000",
  37878=>"000110010",
  37879=>"000111111",
  37880=>"111010000",
  37881=>"010100111",
  37882=>"111100001",
  37883=>"101010000",
  37884=>"010011000",
  37885=>"110100100",
  37886=>"110110100",
  37887=>"011010010",
  37888=>"000110111",
  37889=>"100011000",
  37890=>"000101010",
  37891=>"110110000",
  37892=>"001010000",
  37893=>"100011101",
  37894=>"110001011",
  37895=>"010110100",
  37896=>"000001101",
  37897=>"101011110",
  37898=>"111111111",
  37899=>"100000011",
  37900=>"101011101",
  37901=>"111111011",
  37902=>"100011000",
  37903=>"110101010",
  37904=>"000100001",
  37905=>"000001101",
  37906=>"111010000",
  37907=>"100100001",
  37908=>"101010001",
  37909=>"101010000",
  37910=>"100011010",
  37911=>"101011101",
  37912=>"001100011",
  37913=>"100110010",
  37914=>"100010110",
  37915=>"111011000",
  37916=>"011001000",
  37917=>"100000101",
  37918=>"001111000",
  37919=>"000011110",
  37920=>"101111000",
  37921=>"011000001",
  37922=>"110111011",
  37923=>"001001101",
  37924=>"001111001",
  37925=>"010001000",
  37926=>"111111111",
  37927=>"001110000",
  37928=>"001111010",
  37929=>"101011101",
  37930=>"100101101",
  37931=>"111001010",
  37932=>"000111000",
  37933=>"101010101",
  37934=>"010110000",
  37935=>"100100000",
  37936=>"111111001",
  37937=>"110100100",
  37938=>"110001001",
  37939=>"011000001",
  37940=>"111111011",
  37941=>"110111110",
  37942=>"010100010",
  37943=>"001000000",
  37944=>"111010110",
  37945=>"110111011",
  37946=>"001110001",
  37947=>"110101111",
  37948=>"000111010",
  37949=>"100110010",
  37950=>"100011011",
  37951=>"011101100",
  37952=>"101100001",
  37953=>"000001100",
  37954=>"011101111",
  37955=>"010000000",
  37956=>"000111100",
  37957=>"001100111",
  37958=>"000000000",
  37959=>"110001100",
  37960=>"111101010",
  37961=>"000010111",
  37962=>"110111010",
  37963=>"100000011",
  37964=>"000001001",
  37965=>"000100101",
  37966=>"101010000",
  37967=>"101000110",
  37968=>"111000100",
  37969=>"101111011",
  37970=>"111111100",
  37971=>"111001010",
  37972=>"000100010",
  37973=>"111110011",
  37974=>"011000111",
  37975=>"011010010",
  37976=>"101100101",
  37977=>"011111000",
  37978=>"111111011",
  37979=>"110010000",
  37980=>"101001110",
  37981=>"111010110",
  37982=>"111001000",
  37983=>"111001110",
  37984=>"000101001",
  37985=>"101110111",
  37986=>"111111111",
  37987=>"111000110",
  37988=>"111011110",
  37989=>"001101011",
  37990=>"110111110",
  37991=>"101110010",
  37992=>"111100110",
  37993=>"100011010",
  37994=>"111110010",
  37995=>"111111011",
  37996=>"111101010",
  37997=>"110101111",
  37998=>"110010000",
  37999=>"111101101",
  38000=>"110100100",
  38001=>"111111010",
  38002=>"011110101",
  38003=>"010111001",
  38004=>"010111011",
  38005=>"011101000",
  38006=>"111111101",
  38007=>"000010011",
  38008=>"000100001",
  38009=>"101000111",
  38010=>"000010010",
  38011=>"110111111",
  38012=>"000110100",
  38013=>"100111101",
  38014=>"110101111",
  38015=>"011011011",
  38016=>"101011010",
  38017=>"101010000",
  38018=>"111000110",
  38019=>"011101111",
  38020=>"010010001",
  38021=>"100011110",
  38022=>"110101110",
  38023=>"111111100",
  38024=>"000011000",
  38025=>"010001101",
  38026=>"111100111",
  38027=>"001000110",
  38028=>"010011100",
  38029=>"110001001",
  38030=>"111001010",
  38031=>"111100010",
  38032=>"100110101",
  38033=>"100010100",
  38034=>"111100001",
  38035=>"100101010",
  38036=>"110100111",
  38037=>"101110111",
  38038=>"010111111",
  38039=>"000011100",
  38040=>"001100100",
  38041=>"011011000",
  38042=>"000110010",
  38043=>"001001001",
  38044=>"011110111",
  38045=>"100010011",
  38046=>"011011100",
  38047=>"110100011",
  38048=>"011001100",
  38049=>"100011101",
  38050=>"101111001",
  38051=>"011000011",
  38052=>"100100110",
  38053=>"111110111",
  38054=>"110001001",
  38055=>"001000010",
  38056=>"101100100",
  38057=>"000011001",
  38058=>"100101011",
  38059=>"110110101",
  38060=>"100000000",
  38061=>"000001111",
  38062=>"101110101",
  38063=>"000010000",
  38064=>"001111110",
  38065=>"000000110",
  38066=>"101111110",
  38067=>"011001101",
  38068=>"100110110",
  38069=>"100001110",
  38070=>"111111000",
  38071=>"001111010",
  38072=>"111011000",
  38073=>"001001011",
  38074=>"011101000",
  38075=>"000101001",
  38076=>"011011000",
  38077=>"001110001",
  38078=>"101000100",
  38079=>"001111101",
  38080=>"010101110",
  38081=>"110111010",
  38082=>"101101111",
  38083=>"110100110",
  38084=>"001100110",
  38085=>"101111010",
  38086=>"100111111",
  38087=>"001011000",
  38088=>"101101000",
  38089=>"001001011",
  38090=>"001001111",
  38091=>"110101111",
  38092=>"001100100",
  38093=>"101001000",
  38094=>"000110010",
  38095=>"001001001",
  38096=>"001011001",
  38097=>"100101100",
  38098=>"011000101",
  38099=>"100110111",
  38100=>"111111110",
  38101=>"000101111",
  38102=>"110001000",
  38103=>"100001111",
  38104=>"110000111",
  38105=>"011001010",
  38106=>"001110010",
  38107=>"011110111",
  38108=>"011010010",
  38109=>"110000001",
  38110=>"011000010",
  38111=>"110000100",
  38112=>"011111111",
  38113=>"010001100",
  38114=>"010101110",
  38115=>"000000001",
  38116=>"110110110",
  38117=>"111111111",
  38118=>"100011110",
  38119=>"100101111",
  38120=>"011111110",
  38121=>"011001000",
  38122=>"001010000",
  38123=>"010001111",
  38124=>"000101000",
  38125=>"010010000",
  38126=>"001011110",
  38127=>"010001101",
  38128=>"110010110",
  38129=>"110111000",
  38130=>"110000000",
  38131=>"001000001",
  38132=>"110101111",
  38133=>"010100000",
  38134=>"010101000",
  38135=>"011101111",
  38136=>"110000010",
  38137=>"110001111",
  38138=>"100101000",
  38139=>"100111100",
  38140=>"101101000",
  38141=>"001000010",
  38142=>"100000000",
  38143=>"001011001",
  38144=>"100001000",
  38145=>"000101001",
  38146=>"010110100",
  38147=>"011011100",
  38148=>"000101010",
  38149=>"111111001",
  38150=>"111111101",
  38151=>"110110111",
  38152=>"101000001",
  38153=>"110111011",
  38154=>"111111000",
  38155=>"110001110",
  38156=>"010001110",
  38157=>"010110100",
  38158=>"001110110",
  38159=>"011010111",
  38160=>"001101111",
  38161=>"111010101",
  38162=>"001111010",
  38163=>"100000110",
  38164=>"100000101",
  38165=>"100100011",
  38166=>"100111101",
  38167=>"010001111",
  38168=>"110100101",
  38169=>"011101100",
  38170=>"010101010",
  38171=>"010111001",
  38172=>"101100001",
  38173=>"111101011",
  38174=>"100101100",
  38175=>"111001111",
  38176=>"001101101",
  38177=>"111100111",
  38178=>"111110010",
  38179=>"101110111",
  38180=>"011000010",
  38181=>"110000011",
  38182=>"010111001",
  38183=>"111100000",
  38184=>"010101110",
  38185=>"010100111",
  38186=>"111011010",
  38187=>"001111100",
  38188=>"001000000",
  38189=>"010110101",
  38190=>"101011100",
  38191=>"001110010",
  38192=>"000100100",
  38193=>"101111000",
  38194=>"111001101",
  38195=>"001000101",
  38196=>"010100000",
  38197=>"011010010",
  38198=>"011010101",
  38199=>"010010111",
  38200=>"111111111",
  38201=>"111011101",
  38202=>"110100100",
  38203=>"111000100",
  38204=>"110101011",
  38205=>"100011011",
  38206=>"100000111",
  38207=>"010001010",
  38208=>"011011001",
  38209=>"011011011",
  38210=>"001010011",
  38211=>"000110010",
  38212=>"000100001",
  38213=>"110101000",
  38214=>"101010101",
  38215=>"110011010",
  38216=>"110010100",
  38217=>"111111111",
  38218=>"111110010",
  38219=>"111101001",
  38220=>"000111001",
  38221=>"111000010",
  38222=>"010111001",
  38223=>"111101110",
  38224=>"111110000",
  38225=>"110111110",
  38226=>"011110000",
  38227=>"000101101",
  38228=>"101011111",
  38229=>"011111101",
  38230=>"110001011",
  38231=>"111111111",
  38232=>"001111111",
  38233=>"100111111",
  38234=>"011011101",
  38235=>"101100110",
  38236=>"001101101",
  38237=>"100001001",
  38238=>"110010011",
  38239=>"101111001",
  38240=>"010000000",
  38241=>"111101111",
  38242=>"101010111",
  38243=>"011101111",
  38244=>"101010000",
  38245=>"111100110",
  38246=>"101011001",
  38247=>"100101010",
  38248=>"100101110",
  38249=>"101100001",
  38250=>"010101011",
  38251=>"111101011",
  38252=>"000011011",
  38253=>"000000101",
  38254=>"011001101",
  38255=>"001110111",
  38256=>"010000111",
  38257=>"010011111",
  38258=>"000010011",
  38259=>"000000000",
  38260=>"011101000",
  38261=>"101110110",
  38262=>"011111111",
  38263=>"000010010",
  38264=>"010111100",
  38265=>"001001101",
  38266=>"111110101",
  38267=>"000000111",
  38268=>"011001000",
  38269=>"000110101",
  38270=>"100110110",
  38271=>"100010000",
  38272=>"011010010",
  38273=>"101101001",
  38274=>"110001111",
  38275=>"111000001",
  38276=>"010001111",
  38277=>"100001100",
  38278=>"101111101",
  38279=>"100101010",
  38280=>"000101101",
  38281=>"010100011",
  38282=>"010010111",
  38283=>"100101111",
  38284=>"001101101",
  38285=>"111100110",
  38286=>"001001111",
  38287=>"010111101",
  38288=>"001011101",
  38289=>"111011111",
  38290=>"111110100",
  38291=>"000000110",
  38292=>"101101000",
  38293=>"100101001",
  38294=>"000100001",
  38295=>"000100100",
  38296=>"111101100",
  38297=>"011001110",
  38298=>"101110110",
  38299=>"010101110",
  38300=>"110001100",
  38301=>"010111100",
  38302=>"110011111",
  38303=>"001010110",
  38304=>"101101001",
  38305=>"011011010",
  38306=>"000000110",
  38307=>"011100111",
  38308=>"101111010",
  38309=>"101101101",
  38310=>"011110000",
  38311=>"000000110",
  38312=>"101011010",
  38313=>"100000000",
  38314=>"011110111",
  38315=>"000000100",
  38316=>"110101000",
  38317=>"000011110",
  38318=>"001010110",
  38319=>"010011000",
  38320=>"100011111",
  38321=>"011000010",
  38322=>"000101000",
  38323=>"011010111",
  38324=>"001010001",
  38325=>"100110100",
  38326=>"111011110",
  38327=>"010011000",
  38328=>"100011111",
  38329=>"100011000",
  38330=>"111000011",
  38331=>"110010111",
  38332=>"000111101",
  38333=>"101001011",
  38334=>"011110110",
  38335=>"100111010",
  38336=>"101111010",
  38337=>"101111111",
  38338=>"100001110",
  38339=>"110011101",
  38340=>"111111111",
  38341=>"010111110",
  38342=>"011101000",
  38343=>"101011010",
  38344=>"011111010",
  38345=>"010001011",
  38346=>"110110100",
  38347=>"100101011",
  38348=>"101000000",
  38349=>"111000000",
  38350=>"111011001",
  38351=>"001001100",
  38352=>"101110110",
  38353=>"001010011",
  38354=>"101110110",
  38355=>"110110000",
  38356=>"010100000",
  38357=>"110010010",
  38358=>"010001100",
  38359=>"010000011",
  38360=>"111111101",
  38361=>"010100111",
  38362=>"011111011",
  38363=>"100010100",
  38364=>"000010110",
  38365=>"001010001",
  38366=>"101110111",
  38367=>"010000101",
  38368=>"111100000",
  38369=>"111111100",
  38370=>"110100110",
  38371=>"000011011",
  38372=>"100101000",
  38373=>"100000010",
  38374=>"110000100",
  38375=>"111101100",
  38376=>"110011111",
  38377=>"111100111",
  38378=>"110101000",
  38379=>"000110011",
  38380=>"111100011",
  38381=>"111111110",
  38382=>"110000100",
  38383=>"000111110",
  38384=>"010111100",
  38385=>"011010111",
  38386=>"011111101",
  38387=>"101110110",
  38388=>"010000101",
  38389=>"011000101",
  38390=>"100111000",
  38391=>"110000110",
  38392=>"001011111",
  38393=>"010101000",
  38394=>"101110011",
  38395=>"001100001",
  38396=>"101100101",
  38397=>"000111111",
  38398=>"111000000",
  38399=>"000101111",
  38400=>"101010100",
  38401=>"011111100",
  38402=>"100000001",
  38403=>"010101111",
  38404=>"111100110",
  38405=>"000101111",
  38406=>"100101100",
  38407=>"111011111",
  38408=>"000011100",
  38409=>"111011000",
  38410=>"000000111",
  38411=>"100111101",
  38412=>"101101010",
  38413=>"110101001",
  38414=>"000001111",
  38415=>"001011010",
  38416=>"101001111",
  38417=>"101101001",
  38418=>"000100010",
  38419=>"110001011",
  38420=>"101101110",
  38421=>"001001110",
  38422=>"001100101",
  38423=>"100101001",
  38424=>"111011000",
  38425=>"110111000",
  38426=>"111110110",
  38427=>"100001101",
  38428=>"101001110",
  38429=>"110010100",
  38430=>"010000110",
  38431=>"001100000",
  38432=>"110110110",
  38433=>"110100000",
  38434=>"011101011",
  38435=>"100100000",
  38436=>"111101101",
  38437=>"100011000",
  38438=>"111000110",
  38439=>"101100100",
  38440=>"101101011",
  38441=>"010001010",
  38442=>"000011100",
  38443=>"101000000",
  38444=>"001101101",
  38445=>"110111100",
  38446=>"010111101",
  38447=>"100001001",
  38448=>"100011111",
  38449=>"111110000",
  38450=>"010001100",
  38451=>"101011100",
  38452=>"101011010",
  38453=>"000101101",
  38454=>"101110011",
  38455=>"101010101",
  38456=>"101110001",
  38457=>"000010011",
  38458=>"011110111",
  38459=>"101100010",
  38460=>"100100101",
  38461=>"100101001",
  38462=>"110111111",
  38463=>"000001001",
  38464=>"100000001",
  38465=>"001011100",
  38466=>"011000101",
  38467=>"010000000",
  38468=>"110011001",
  38469=>"110001001",
  38470=>"010101110",
  38471=>"111000110",
  38472=>"110110101",
  38473=>"001001000",
  38474=>"011110011",
  38475=>"000100001",
  38476=>"110010000",
  38477=>"001110001",
  38478=>"101011111",
  38479=>"110111111",
  38480=>"111000111",
  38481=>"011010101",
  38482=>"111011010",
  38483=>"111111101",
  38484=>"111101001",
  38485=>"110100011",
  38486=>"111011100",
  38487=>"100100010",
  38488=>"010000110",
  38489=>"111010011",
  38490=>"110110100",
  38491=>"111101111",
  38492=>"110010000",
  38493=>"001011111",
  38494=>"110011000",
  38495=>"000000001",
  38496=>"111110100",
  38497=>"011101111",
  38498=>"110101000",
  38499=>"111100100",
  38500=>"100101010",
  38501=>"101101101",
  38502=>"010001011",
  38503=>"001111110",
  38504=>"111111101",
  38505=>"000001010",
  38506=>"100100110",
  38507=>"001101000",
  38508=>"111001110",
  38509=>"000000110",
  38510=>"101010011",
  38511=>"111111110",
  38512=>"010001011",
  38513=>"101101110",
  38514=>"111111111",
  38515=>"011011111",
  38516=>"000011001",
  38517=>"110010101",
  38518=>"100101011",
  38519=>"111101110",
  38520=>"001000010",
  38521=>"001101010",
  38522=>"011111011",
  38523=>"101011110",
  38524=>"001110010",
  38525=>"111111100",
  38526=>"001000100",
  38527=>"101011100",
  38528=>"101000100",
  38529=>"010000010",
  38530=>"111100011",
  38531=>"110110110",
  38532=>"101100111",
  38533=>"101011111",
  38534=>"001000001",
  38535=>"101111010",
  38536=>"101000101",
  38537=>"110011000",
  38538=>"000010110",
  38539=>"001101111",
  38540=>"110111011",
  38541=>"001110110",
  38542=>"000111111",
  38543=>"010111000",
  38544=>"000110111",
  38545=>"000010100",
  38546=>"111001000",
  38547=>"010010000",
  38548=>"001010101",
  38549=>"011110111",
  38550=>"001101101",
  38551=>"001010101",
  38552=>"000011100",
  38553=>"010110101",
  38554=>"101110100",
  38555=>"000001000",
  38556=>"010010110",
  38557=>"101010011",
  38558=>"110111110",
  38559=>"101100010",
  38560=>"101100101",
  38561=>"111100001",
  38562=>"111111110",
  38563=>"010011111",
  38564=>"100101010",
  38565=>"001010110",
  38566=>"101001000",
  38567=>"101011111",
  38568=>"001101000",
  38569=>"101111110",
  38570=>"111110110",
  38571=>"100110000",
  38572=>"010101001",
  38573=>"011111011",
  38574=>"001110111",
  38575=>"010111100",
  38576=>"110110110",
  38577=>"001100110",
  38578=>"111010100",
  38579=>"101100101",
  38580=>"111001010",
  38581=>"011000011",
  38582=>"110001110",
  38583=>"010110111",
  38584=>"110100110",
  38585=>"100110010",
  38586=>"110110011",
  38587=>"010100011",
  38588=>"011111111",
  38589=>"110011110",
  38590=>"010010011",
  38591=>"101010101",
  38592=>"110110011",
  38593=>"100111111",
  38594=>"101111000",
  38595=>"101111001",
  38596=>"000110000",
  38597=>"101010010",
  38598=>"110010110",
  38599=>"010110010",
  38600=>"101111101",
  38601=>"110100001",
  38602=>"101100000",
  38603=>"010100110",
  38604=>"111010101",
  38605=>"111111000",
  38606=>"010011000",
  38607=>"100111010",
  38608=>"111111000",
  38609=>"101111011",
  38610=>"000010011",
  38611=>"010110101",
  38612=>"001001101",
  38613=>"101101111",
  38614=>"100101110",
  38615=>"110101011",
  38616=>"001110001",
  38617=>"110000001",
  38618=>"001010010",
  38619=>"011000010",
  38620=>"010111010",
  38621=>"100100000",
  38622=>"111010011",
  38623=>"010000100",
  38624=>"111000000",
  38625=>"001000100",
  38626=>"001101010",
  38627=>"100111101",
  38628=>"101111011",
  38629=>"101000001",
  38630=>"011010110",
  38631=>"000011010",
  38632=>"111001010",
  38633=>"011011100",
  38634=>"011111101",
  38635=>"001010011",
  38636=>"101000110",
  38637=>"101110110",
  38638=>"000010000",
  38639=>"110111111",
  38640=>"110101101",
  38641=>"111100111",
  38642=>"010111001",
  38643=>"010000001",
  38644=>"111101111",
  38645=>"111101000",
  38646=>"000110000",
  38647=>"000010000",
  38648=>"110110100",
  38649=>"000100110",
  38650=>"110001101",
  38651=>"011111111",
  38652=>"111000010",
  38653=>"100000010",
  38654=>"011110111",
  38655=>"100010000",
  38656=>"000101100",
  38657=>"111111011",
  38658=>"010010100",
  38659=>"110011000",
  38660=>"101010000",
  38661=>"101001111",
  38662=>"111010010",
  38663=>"000000100",
  38664=>"001100101",
  38665=>"101000001",
  38666=>"010000100",
  38667=>"001011101",
  38668=>"100001111",
  38669=>"010101001",
  38670=>"000100011",
  38671=>"011101011",
  38672=>"111010001",
  38673=>"010001010",
  38674=>"101110000",
  38675=>"000011101",
  38676=>"010111011",
  38677=>"111110111",
  38678=>"110001000",
  38679=>"011110011",
  38680=>"111011010",
  38681=>"110110110",
  38682=>"011010101",
  38683=>"111101000",
  38684=>"011110001",
  38685=>"110111101",
  38686=>"100101101",
  38687=>"011011100",
  38688=>"011000000",
  38689=>"010111110",
  38690=>"100001010",
  38691=>"111011111",
  38692=>"111011110",
  38693=>"000100000",
  38694=>"010111111",
  38695=>"110100110",
  38696=>"101010000",
  38697=>"110011111",
  38698=>"010011010",
  38699=>"101001100",
  38700=>"011100100",
  38701=>"111011011",
  38702=>"001111011",
  38703=>"110101011",
  38704=>"010101100",
  38705=>"011000010",
  38706=>"010011011",
  38707=>"101100001",
  38708=>"100100000",
  38709=>"001010010",
  38710=>"001001110",
  38711=>"010001101",
  38712=>"000001010",
  38713=>"110111011",
  38714=>"011011111",
  38715=>"110011100",
  38716=>"001110111",
  38717=>"011110001",
  38718=>"111101001",
  38719=>"111010101",
  38720=>"000000110",
  38721=>"100110001",
  38722=>"101001000",
  38723=>"011010010",
  38724=>"100100011",
  38725=>"000011001",
  38726=>"101001000",
  38727=>"010111110",
  38728=>"011001001",
  38729=>"101000100",
  38730=>"011011000",
  38731=>"001000100",
  38732=>"101100100",
  38733=>"100001111",
  38734=>"001001001",
  38735=>"100001111",
  38736=>"101101000",
  38737=>"111011011",
  38738=>"111111111",
  38739=>"001110010",
  38740=>"011000010",
  38741=>"110111111",
  38742=>"110110010",
  38743=>"010100011",
  38744=>"110110101",
  38745=>"011001011",
  38746=>"111101011",
  38747=>"111010001",
  38748=>"000011010",
  38749=>"111001101",
  38750=>"001011111",
  38751=>"101111101",
  38752=>"111011001",
  38753=>"111110100",
  38754=>"111010111",
  38755=>"010010011",
  38756=>"010011110",
  38757=>"000010011",
  38758=>"011010011",
  38759=>"101010010",
  38760=>"011000001",
  38761=>"010010000",
  38762=>"110100101",
  38763=>"010111000",
  38764=>"001001000",
  38765=>"101110100",
  38766=>"001111111",
  38767=>"101111110",
  38768=>"000101000",
  38769=>"001001010",
  38770=>"010100001",
  38771=>"011000110",
  38772=>"101111001",
  38773=>"101110110",
  38774=>"110100000",
  38775=>"000110010",
  38776=>"101001111",
  38777=>"000010100",
  38778=>"010011110",
  38779=>"011001110",
  38780=>"111110111",
  38781=>"100101011",
  38782=>"101110110",
  38783=>"110111110",
  38784=>"101111011",
  38785=>"110100010",
  38786=>"000001000",
  38787=>"110000111",
  38788=>"110011111",
  38789=>"000010111",
  38790=>"101110101",
  38791=>"010001011",
  38792=>"010100000",
  38793=>"101110110",
  38794=>"010111010",
  38795=>"100001000",
  38796=>"010100110",
  38797=>"101010010",
  38798=>"011010100",
  38799=>"111010000",
  38800=>"110011010",
  38801=>"101101101",
  38802=>"101011111",
  38803=>"100010000",
  38804=>"110010010",
  38805=>"000001010",
  38806=>"110000010",
  38807=>"101101000",
  38808=>"010111111",
  38809=>"010111101",
  38810=>"000111011",
  38811=>"111001011",
  38812=>"110100110",
  38813=>"110110101",
  38814=>"110011001",
  38815=>"110000111",
  38816=>"111110100",
  38817=>"001110100",
  38818=>"110111010",
  38819=>"101001100",
  38820=>"001001110",
  38821=>"010100110",
  38822=>"010110011",
  38823=>"011010110",
  38824=>"010101010",
  38825=>"000000111",
  38826=>"000000110",
  38827=>"110001010",
  38828=>"011101110",
  38829=>"110100101",
  38830=>"010010000",
  38831=>"011011111",
  38832=>"110100000",
  38833=>"110000100",
  38834=>"110001101",
  38835=>"110011100",
  38836=>"100000001",
  38837=>"001101100",
  38838=>"001011100",
  38839=>"100100100",
  38840=>"101010000",
  38841=>"011010110",
  38842=>"110100011",
  38843=>"001100011",
  38844=>"111111010",
  38845=>"110101001",
  38846=>"101010100",
  38847=>"011101110",
  38848=>"111000001",
  38849=>"001010111",
  38850=>"010110110",
  38851=>"000001000",
  38852=>"101101100",
  38853=>"110111001",
  38854=>"111110000",
  38855=>"000011110",
  38856=>"000011100",
  38857=>"111111011",
  38858=>"010011101",
  38859=>"001111001",
  38860=>"001110000",
  38861=>"000000011",
  38862=>"010111010",
  38863=>"111111100",
  38864=>"111110111",
  38865=>"111111010",
  38866=>"111001111",
  38867=>"100001111",
  38868=>"010011011",
  38869=>"111000000",
  38870=>"101000110",
  38871=>"010010000",
  38872=>"110011110",
  38873=>"111111100",
  38874=>"110001011",
  38875=>"000001110",
  38876=>"100000101",
  38877=>"111011011",
  38878=>"100001111",
  38879=>"111000100",
  38880=>"101110111",
  38881=>"011011110",
  38882=>"010001100",
  38883=>"110010110",
  38884=>"000010011",
  38885=>"111011111",
  38886=>"110001111",
  38887=>"011101111",
  38888=>"011010111",
  38889=>"101010111",
  38890=>"011010100",
  38891=>"001101000",
  38892=>"001010101",
  38893=>"111000111",
  38894=>"000111101",
  38895=>"010011100",
  38896=>"011110000",
  38897=>"010011000",
  38898=>"011100000",
  38899=>"100100101",
  38900=>"011111001",
  38901=>"010110010",
  38902=>"010000000",
  38903=>"101100001",
  38904=>"010111011",
  38905=>"011000111",
  38906=>"010011101",
  38907=>"111000001",
  38908=>"111001111",
  38909=>"001010011",
  38910=>"100001011",
  38911=>"011001111",
  38912=>"000011100",
  38913=>"001010000",
  38914=>"010110011",
  38915=>"010110010",
  38916=>"101011111",
  38917=>"101000110",
  38918=>"110100110",
  38919=>"011000000",
  38920=>"111011010",
  38921=>"101111111",
  38922=>"111101110",
  38923=>"110110111",
  38924=>"111100100",
  38925=>"001101000",
  38926=>"101100000",
  38927=>"000010000",
  38928=>"101111100",
  38929=>"100101000",
  38930=>"101001011",
  38931=>"101010110",
  38932=>"011010110",
  38933=>"000101101",
  38934=>"000010110",
  38935=>"100000010",
  38936=>"001110100",
  38937=>"010010100",
  38938=>"010110101",
  38939=>"001111111",
  38940=>"101110100",
  38941=>"000100110",
  38942=>"111111001",
  38943=>"010101010",
  38944=>"101111101",
  38945=>"011001100",
  38946=>"000010010",
  38947=>"001010010",
  38948=>"110101111",
  38949=>"000111000",
  38950=>"010111100",
  38951=>"101100010",
  38952=>"101110100",
  38953=>"000001010",
  38954=>"111000000",
  38955=>"101100111",
  38956=>"111110111",
  38957=>"101100000",
  38958=>"001100110",
  38959=>"100110100",
  38960=>"111001010",
  38961=>"000111000",
  38962=>"111111111",
  38963=>"110011101",
  38964=>"101001110",
  38965=>"110110110",
  38966=>"000111010",
  38967=>"100110010",
  38968=>"110010101",
  38969=>"010110010",
  38970=>"010001010",
  38971=>"010000010",
  38972=>"000111111",
  38973=>"000101111",
  38974=>"010110010",
  38975=>"011100001",
  38976=>"101001100",
  38977=>"011001100",
  38978=>"010010000",
  38979=>"000100111",
  38980=>"001001000",
  38981=>"001110111",
  38982=>"110001100",
  38983=>"100111000",
  38984=>"010100011",
  38985=>"001001101",
  38986=>"011010100",
  38987=>"011001001",
  38988=>"111001100",
  38989=>"101010101",
  38990=>"010011011",
  38991=>"110100010",
  38992=>"001011010",
  38993=>"111010111",
  38994=>"001011111",
  38995=>"110111111",
  38996=>"011111000",
  38997=>"000110110",
  38998=>"101010111",
  38999=>"011000110",
  39000=>"110100001",
  39001=>"011001111",
  39002=>"001011100",
  39003=>"011101000",
  39004=>"000111000",
  39005=>"001000010",
  39006=>"111010001",
  39007=>"001000001",
  39008=>"111100111",
  39009=>"101100011",
  39010=>"101000110",
  39011=>"110101110",
  39012=>"001111111",
  39013=>"100100101",
  39014=>"111010110",
  39015=>"001000010",
  39016=>"001100110",
  39017=>"001001100",
  39018=>"111100100",
  39019=>"010011011",
  39020=>"111110010",
  39021=>"100010110",
  39022=>"110011001",
  39023=>"000111000",
  39024=>"111100011",
  39025=>"101100100",
  39026=>"110101010",
  39027=>"101110100",
  39028=>"111100010",
  39029=>"100100000",
  39030=>"101110011",
  39031=>"011100101",
  39032=>"100111010",
  39033=>"100000100",
  39034=>"000110011",
  39035=>"101001101",
  39036=>"011111101",
  39037=>"000101111",
  39038=>"000100001",
  39039=>"000011100",
  39040=>"000001011",
  39041=>"011101111",
  39042=>"100010010",
  39043=>"001111100",
  39044=>"011010100",
  39045=>"010000101",
  39046=>"000000011",
  39047=>"111100001",
  39048=>"101111101",
  39049=>"010011110",
  39050=>"110110110",
  39051=>"111100100",
  39052=>"101110111",
  39053=>"101001001",
  39054=>"110110111",
  39055=>"001011001",
  39056=>"001001100",
  39057=>"000001110",
  39058=>"111010000",
  39059=>"111110000",
  39060=>"010011101",
  39061=>"101001001",
  39062=>"001100111",
  39063=>"100000101",
  39064=>"100100110",
  39065=>"111010111",
  39066=>"101111101",
  39067=>"011111000",
  39068=>"111100100",
  39069=>"000110000",
  39070=>"000010011",
  39071=>"010000001",
  39072=>"111100011",
  39073=>"000010111",
  39074=>"000000110",
  39075=>"011001001",
  39076=>"001000111",
  39077=>"000011110",
  39078=>"100011110",
  39079=>"100000100",
  39080=>"111111010",
  39081=>"111000011",
  39082=>"001001001",
  39083=>"010011111",
  39084=>"000111110",
  39085=>"001000100",
  39086=>"011011000",
  39087=>"011100011",
  39088=>"100010001",
  39089=>"111001111",
  39090=>"011111000",
  39091=>"000010010",
  39092=>"100010000",
  39093=>"001101101",
  39094=>"011101100",
  39095=>"010000100",
  39096=>"110010001",
  39097=>"101000010",
  39098=>"101100110",
  39099=>"001000111",
  39100=>"011011111",
  39101=>"011111101",
  39102=>"100101110",
  39103=>"111011100",
  39104=>"110100001",
  39105=>"010110101",
  39106=>"011001011",
  39107=>"000101000",
  39108=>"101010100",
  39109=>"101100101",
  39110=>"000110110",
  39111=>"011001111",
  39112=>"111011010",
  39113=>"100010011",
  39114=>"001110010",
  39115=>"000101101",
  39116=>"010011101",
  39117=>"000100110",
  39118=>"101001000",
  39119=>"101000111",
  39120=>"011011010",
  39121=>"001010100",
  39122=>"111111010",
  39123=>"011101100",
  39124=>"000000000",
  39125=>"000101001",
  39126=>"001110010",
  39127=>"000111110",
  39128=>"101110100",
  39129=>"000010100",
  39130=>"110110111",
  39131=>"101111111",
  39132=>"011100000",
  39133=>"110010000",
  39134=>"001011101",
  39135=>"110111100",
  39136=>"000010111",
  39137=>"000100111",
  39138=>"100100101",
  39139=>"111111111",
  39140=>"101011010",
  39141=>"101100110",
  39142=>"111000000",
  39143=>"111100010",
  39144=>"000010001",
  39145=>"000001000",
  39146=>"111110101",
  39147=>"111011111",
  39148=>"010100111",
  39149=>"101110111",
  39150=>"100111011",
  39151=>"000101010",
  39152=>"110000001",
  39153=>"111101111",
  39154=>"011010011",
  39155=>"010011110",
  39156=>"111100000",
  39157=>"110100100",
  39158=>"101011000",
  39159=>"010100000",
  39160=>"000110110",
  39161=>"100110101",
  39162=>"000111111",
  39163=>"001100010",
  39164=>"010111101",
  39165=>"111100100",
  39166=>"111001000",
  39167=>"011010101",
  39168=>"010011100",
  39169=>"100110101",
  39170=>"101110110",
  39171=>"000000001",
  39172=>"010011101",
  39173=>"100010001",
  39174=>"001000100",
  39175=>"100100011",
  39176=>"000000100",
  39177=>"110101101",
  39178=>"010010101",
  39179=>"010001101",
  39180=>"000001110",
  39181=>"111110100",
  39182=>"111100000",
  39183=>"011110000",
  39184=>"000111110",
  39185=>"001000110",
  39186=>"101000100",
  39187=>"100010001",
  39188=>"111000100",
  39189=>"000011000",
  39190=>"010010111",
  39191=>"011011101",
  39192=>"000100010",
  39193=>"000000110",
  39194=>"110111111",
  39195=>"010010111",
  39196=>"101001110",
  39197=>"000001111",
  39198=>"000011011",
  39199=>"100100100",
  39200=>"101110010",
  39201=>"101010011",
  39202=>"011110001",
  39203=>"110101000",
  39204=>"000100100",
  39205=>"110111000",
  39206=>"100010001",
  39207=>"010001001",
  39208=>"011000100",
  39209=>"011111111",
  39210=>"011110011",
  39211=>"111011001",
  39212=>"110101010",
  39213=>"010000000",
  39214=>"000101010",
  39215=>"000110000",
  39216=>"110010100",
  39217=>"010010111",
  39218=>"001101001",
  39219=>"001100000",
  39220=>"010000011",
  39221=>"110110000",
  39222=>"100011111",
  39223=>"110101001",
  39224=>"011011101",
  39225=>"110001000",
  39226=>"000111110",
  39227=>"110100101",
  39228=>"110000111",
  39229=>"111000011",
  39230=>"010000100",
  39231=>"001011010",
  39232=>"011101111",
  39233=>"010100001",
  39234=>"000100100",
  39235=>"000011100",
  39236=>"010100000",
  39237=>"101101101",
  39238=>"000000010",
  39239=>"011010110",
  39240=>"000000010",
  39241=>"101111100",
  39242=>"011011010",
  39243=>"110111101",
  39244=>"101010011",
  39245=>"100001011",
  39246=>"110010001",
  39247=>"011111001",
  39248=>"100101100",
  39249=>"011101001",
  39250=>"011111111",
  39251=>"111001111",
  39252=>"110111011",
  39253=>"010111101",
  39254=>"000100111",
  39255=>"011010000",
  39256=>"001110010",
  39257=>"110100111",
  39258=>"011011100",
  39259=>"001110010",
  39260=>"111100000",
  39261=>"101101011",
  39262=>"101000011",
  39263=>"100111100",
  39264=>"001011100",
  39265=>"110000101",
  39266=>"101110001",
  39267=>"011010001",
  39268=>"100111100",
  39269=>"010011010",
  39270=>"011110100",
  39271=>"111101001",
  39272=>"101101110",
  39273=>"010010010",
  39274=>"111111101",
  39275=>"101000001",
  39276=>"111011001",
  39277=>"100001011",
  39278=>"101100111",
  39279=>"111101111",
  39280=>"110000100",
  39281=>"111000011",
  39282=>"001111010",
  39283=>"010100111",
  39284=>"010111010",
  39285=>"010100100",
  39286=>"000011110",
  39287=>"100011100",
  39288=>"110111101",
  39289=>"010111101",
  39290=>"010111000",
  39291=>"011000001",
  39292=>"000001011",
  39293=>"110101101",
  39294=>"000000111",
  39295=>"000100001",
  39296=>"001101111",
  39297=>"100001101",
  39298=>"101011111",
  39299=>"000011110",
  39300=>"101101110",
  39301=>"001010110",
  39302=>"111010111",
  39303=>"010101010",
  39304=>"000001011",
  39305=>"111001001",
  39306=>"100110011",
  39307=>"111001101",
  39308=>"000001001",
  39309=>"110011101",
  39310=>"110011101",
  39311=>"011111011",
  39312=>"100110111",
  39313=>"100101011",
  39314=>"100110001",
  39315=>"101001111",
  39316=>"010110010",
  39317=>"111001000",
  39318=>"011100101",
  39319=>"111000100",
  39320=>"100101000",
  39321=>"111010111",
  39322=>"000000100",
  39323=>"011001101",
  39324=>"010100001",
  39325=>"001000110",
  39326=>"011111101",
  39327=>"100111100",
  39328=>"111000001",
  39329=>"110000110",
  39330=>"000011100",
  39331=>"111100001",
  39332=>"011011011",
  39333=>"000100001",
  39334=>"110101011",
  39335=>"111100111",
  39336=>"011100100",
  39337=>"101100111",
  39338=>"010000011",
  39339=>"000011111",
  39340=>"000111011",
  39341=>"110000110",
  39342=>"111101100",
  39343=>"111111000",
  39344=>"010110000",
  39345=>"010100011",
  39346=>"010001000",
  39347=>"111110011",
  39348=>"001101111",
  39349=>"001101110",
  39350=>"110111101",
  39351=>"101001000",
  39352=>"001000101",
  39353=>"100111010",
  39354=>"101110111",
  39355=>"111111110",
  39356=>"100000001",
  39357=>"000101001",
  39358=>"110001010",
  39359=>"001111101",
  39360=>"101110100",
  39361=>"010101110",
  39362=>"001110100",
  39363=>"010011010",
  39364=>"010010010",
  39365=>"000010010",
  39366=>"010011001",
  39367=>"000110110",
  39368=>"011100010",
  39369=>"110100100",
  39370=>"111011010",
  39371=>"101111011",
  39372=>"101110100",
  39373=>"111000100",
  39374=>"110101011",
  39375=>"001011111",
  39376=>"110001101",
  39377=>"111101010",
  39378=>"010110110",
  39379=>"001000010",
  39380=>"101000011",
  39381=>"001000001",
  39382=>"110101100",
  39383=>"101000100",
  39384=>"010100101",
  39385=>"111100100",
  39386=>"000001011",
  39387=>"000111111",
  39388=>"001101101",
  39389=>"100011011",
  39390=>"000101011",
  39391=>"111001001",
  39392=>"100100101",
  39393=>"011011111",
  39394=>"001001111",
  39395=>"011100111",
  39396=>"001110000",
  39397=>"011000010",
  39398=>"101100101",
  39399=>"101101001",
  39400=>"011001000",
  39401=>"101101010",
  39402=>"100100011",
  39403=>"000010100",
  39404=>"010001000",
  39405=>"101001011",
  39406=>"001001000",
  39407=>"001011111",
  39408=>"110111011",
  39409=>"001000100",
  39410=>"111110000",
  39411=>"110100100",
  39412=>"000011010",
  39413=>"011110100",
  39414=>"110110001",
  39415=>"000010100",
  39416=>"000001001",
  39417=>"010101111",
  39418=>"001010011",
  39419=>"110010001",
  39420=>"001110001",
  39421=>"111110001",
  39422=>"000100110",
  39423=>"111101011",
  39424=>"100011000",
  39425=>"010101010",
  39426=>"001001101",
  39427=>"101101011",
  39428=>"110001101",
  39429=>"100011001",
  39430=>"100101011",
  39431=>"001111101",
  39432=>"111000111",
  39433=>"111110000",
  39434=>"011110110",
  39435=>"000001000",
  39436=>"101001101",
  39437=>"000111111",
  39438=>"010001101",
  39439=>"110010011",
  39440=>"010011100",
  39441=>"001101111",
  39442=>"010000010",
  39443=>"110000101",
  39444=>"110000001",
  39445=>"111110111",
  39446=>"011100111",
  39447=>"011111011",
  39448=>"101011110",
  39449=>"011001111",
  39450=>"010110101",
  39451=>"111001000",
  39452=>"000101011",
  39453=>"101001100",
  39454=>"101110001",
  39455=>"111101110",
  39456=>"011010101",
  39457=>"010010011",
  39458=>"001001101",
  39459=>"111000010",
  39460=>"000010010",
  39461=>"001110111",
  39462=>"010011100",
  39463=>"001110010",
  39464=>"010100101",
  39465=>"100100111",
  39466=>"111000011",
  39467=>"101110111",
  39468=>"100100000",
  39469=>"001001001",
  39470=>"011001110",
  39471=>"000000101",
  39472=>"001001011",
  39473=>"110101011",
  39474=>"100001000",
  39475=>"110000111",
  39476=>"111010101",
  39477=>"001100001",
  39478=>"111001001",
  39479=>"100111000",
  39480=>"110001010",
  39481=>"010010110",
  39482=>"001100100",
  39483=>"000100010",
  39484=>"010001001",
  39485=>"111001101",
  39486=>"011011111",
  39487=>"110001011",
  39488=>"010100100",
  39489=>"000010011",
  39490=>"100000000",
  39491=>"000000101",
  39492=>"100111000",
  39493=>"011000110",
  39494=>"101010100",
  39495=>"011101111",
  39496=>"001010111",
  39497=>"001000010",
  39498=>"110110001",
  39499=>"101000011",
  39500=>"011010101",
  39501=>"001000000",
  39502=>"100101111",
  39503=>"110101000",
  39504=>"111111110",
  39505=>"100111001",
  39506=>"111101011",
  39507=>"101010111",
  39508=>"100111010",
  39509=>"101101001",
  39510=>"101101111",
  39511=>"100100101",
  39512=>"101111010",
  39513=>"110100001",
  39514=>"010000001",
  39515=>"101110100",
  39516=>"001000100",
  39517=>"000100101",
  39518=>"011110111",
  39519=>"101110001",
  39520=>"111010111",
  39521=>"101000000",
  39522=>"011010011",
  39523=>"000111111",
  39524=>"100101111",
  39525=>"101100110",
  39526=>"111101111",
  39527=>"101110011",
  39528=>"100110011",
  39529=>"100100100",
  39530=>"110011000",
  39531=>"011101010",
  39532=>"001110010",
  39533=>"001001000",
  39534=>"011010111",
  39535=>"111111011",
  39536=>"100001111",
  39537=>"000101111",
  39538=>"110100010",
  39539=>"101110101",
  39540=>"100000101",
  39541=>"011111001",
  39542=>"001001011",
  39543=>"000100001",
  39544=>"111101100",
  39545=>"000000111",
  39546=>"100111110",
  39547=>"110010001",
  39548=>"111101010",
  39549=>"100000100",
  39550=>"111111000",
  39551=>"010100000",
  39552=>"011100111",
  39553=>"000010100",
  39554=>"011000000",
  39555=>"101110101",
  39556=>"100000010",
  39557=>"101111101",
  39558=>"111010010",
  39559=>"100101111",
  39560=>"010000000",
  39561=>"000010011",
  39562=>"000011101",
  39563=>"011011100",
  39564=>"001001011",
  39565=>"111101100",
  39566=>"100100001",
  39567=>"000101000",
  39568=>"101011000",
  39569=>"010101010",
  39570=>"001001011",
  39571=>"010010010",
  39572=>"101101001",
  39573=>"000000101",
  39574=>"111110111",
  39575=>"010111111",
  39576=>"110000100",
  39577=>"001010011",
  39578=>"000100011",
  39579=>"100100100",
  39580=>"101001110",
  39581=>"101001100",
  39582=>"100000001",
  39583=>"110111110",
  39584=>"000110010",
  39585=>"001000100",
  39586=>"001111111",
  39587=>"001001110",
  39588=>"100001110",
  39589=>"010110000",
  39590=>"101000110",
  39591=>"000100111",
  39592=>"101011101",
  39593=>"011011000",
  39594=>"001110010",
  39595=>"001000111",
  39596=>"001000110",
  39597=>"001001001",
  39598=>"000111111",
  39599=>"000010011",
  39600=>"011111000",
  39601=>"111111111",
  39602=>"001001001",
  39603=>"101110000",
  39604=>"001000110",
  39605=>"111000100",
  39606=>"011111000",
  39607=>"010111010",
  39608=>"111101111",
  39609=>"101011100",
  39610=>"100110111",
  39611=>"001000010",
  39612=>"001000001",
  39613=>"100111111",
  39614=>"000101011",
  39615=>"011001110",
  39616=>"011101000",
  39617=>"101011100",
  39618=>"110110101",
  39619=>"110101000",
  39620=>"000001001",
  39621=>"001011101",
  39622=>"101011111",
  39623=>"001001110",
  39624=>"010111100",
  39625=>"101111111",
  39626=>"100101011",
  39627=>"000001101",
  39628=>"100110100",
  39629=>"001111000",
  39630=>"001011110",
  39631=>"000001001",
  39632=>"110100100",
  39633=>"100110011",
  39634=>"100110111",
  39635=>"010010000",
  39636=>"111111001",
  39637=>"001101000",
  39638=>"000010111",
  39639=>"110000111",
  39640=>"001011101",
  39641=>"101010010",
  39642=>"110000000",
  39643=>"101011111",
  39644=>"111101010",
  39645=>"100110111",
  39646=>"101011111",
  39647=>"110100011",
  39648=>"001011011",
  39649=>"100010110",
  39650=>"010101000",
  39651=>"100011110",
  39652=>"000101111",
  39653=>"011101111",
  39654=>"111000000",
  39655=>"010100101",
  39656=>"111001110",
  39657=>"101000101",
  39658=>"111011000",
  39659=>"100000010",
  39660=>"000001001",
  39661=>"011000010",
  39662=>"101101101",
  39663=>"111011101",
  39664=>"101111100",
  39665=>"101010010",
  39666=>"010010110",
  39667=>"101001101",
  39668=>"001101100",
  39669=>"110110101",
  39670=>"010010001",
  39671=>"010100000",
  39672=>"001100000",
  39673=>"000101001",
  39674=>"111011100",
  39675=>"001110010",
  39676=>"101111100",
  39677=>"111100011",
  39678=>"000111000",
  39679=>"101110111",
  39680=>"110101011",
  39681=>"001001010",
  39682=>"100011111",
  39683=>"111101110",
  39684=>"001111010",
  39685=>"000010100",
  39686=>"010010100",
  39687=>"000000000",
  39688=>"011011011",
  39689=>"111011001",
  39690=>"100000001",
  39691=>"001110101",
  39692=>"111000010",
  39693=>"001110100",
  39694=>"001100010",
  39695=>"111111111",
  39696=>"100001101",
  39697=>"001000110",
  39698=>"000011000",
  39699=>"000000101",
  39700=>"000100111",
  39701=>"111101001",
  39702=>"110000000",
  39703=>"111000000",
  39704=>"110010100",
  39705=>"000110111",
  39706=>"100010000",
  39707=>"010100101",
  39708=>"110111011",
  39709=>"100000010",
  39710=>"010110011",
  39711=>"101111000",
  39712=>"110100111",
  39713=>"000011101",
  39714=>"110001010",
  39715=>"101001011",
  39716=>"100010011",
  39717=>"111111100",
  39718=>"001110010",
  39719=>"010001110",
  39720=>"110101101",
  39721=>"111010001",
  39722=>"011001110",
  39723=>"101000011",
  39724=>"001101010",
  39725=>"111101110",
  39726=>"101110001",
  39727=>"110111110",
  39728=>"001111101",
  39729=>"011100100",
  39730=>"010111111",
  39731=>"100110000",
  39732=>"101111111",
  39733=>"110110110",
  39734=>"111000111",
  39735=>"001100011",
  39736=>"100011001",
  39737=>"110101000",
  39738=>"001111111",
  39739=>"101111101",
  39740=>"110100110",
  39741=>"101110101",
  39742=>"101101111",
  39743=>"110011111",
  39744=>"100000001",
  39745=>"000110000",
  39746=>"101010010",
  39747=>"011100001",
  39748=>"111111110",
  39749=>"001101000",
  39750=>"110001100",
  39751=>"001100000",
  39752=>"000100010",
  39753=>"101011110",
  39754=>"110011100",
  39755=>"110011010",
  39756=>"111010000",
  39757=>"110101101",
  39758=>"100111111",
  39759=>"000110011",
  39760=>"110111010",
  39761=>"000001010",
  39762=>"111101011",
  39763=>"001110000",
  39764=>"101110010",
  39765=>"100101000",
  39766=>"101000001",
  39767=>"100100011",
  39768=>"101110011",
  39769=>"111100100",
  39770=>"011001010",
  39771=>"100110111",
  39772=>"110010010",
  39773=>"001001011",
  39774=>"001010011",
  39775=>"001110001",
  39776=>"001100111",
  39777=>"011011011",
  39778=>"001001101",
  39779=>"101110001",
  39780=>"010000100",
  39781=>"010010010",
  39782=>"001100011",
  39783=>"100010100",
  39784=>"100111111",
  39785=>"100101011",
  39786=>"011001110",
  39787=>"101011010",
  39788=>"011000100",
  39789=>"000110101",
  39790=>"010000010",
  39791=>"100001010",
  39792=>"011011010",
  39793=>"101110111",
  39794=>"001111000",
  39795=>"101000110",
  39796=>"001010001",
  39797=>"100110010",
  39798=>"011011010",
  39799=>"111101000",
  39800=>"010110100",
  39801=>"011111100",
  39802=>"100111010",
  39803=>"101100110",
  39804=>"110010111",
  39805=>"001110110",
  39806=>"111101000",
  39807=>"101101011",
  39808=>"001000111",
  39809=>"000010111",
  39810=>"111100000",
  39811=>"100001001",
  39812=>"000001111",
  39813=>"110001100",
  39814=>"000100011",
  39815=>"110100001",
  39816=>"000110100",
  39817=>"101101110",
  39818=>"011111111",
  39819=>"100000000",
  39820=>"001111101",
  39821=>"101000100",
  39822=>"000110001",
  39823=>"100000110",
  39824=>"011111010",
  39825=>"110000000",
  39826=>"110100001",
  39827=>"011001001",
  39828=>"110010111",
  39829=>"001000100",
  39830=>"001111101",
  39831=>"100001000",
  39832=>"111000001",
  39833=>"010011010",
  39834=>"111101100",
  39835=>"000010010",
  39836=>"001000111",
  39837=>"111100011",
  39838=>"000010111",
  39839=>"101011101",
  39840=>"100001101",
  39841=>"011110101",
  39842=>"000101111",
  39843=>"111000110",
  39844=>"000010011",
  39845=>"010111000",
  39846=>"011100011",
  39847=>"100001101",
  39848=>"111100101",
  39849=>"000010000",
  39850=>"110100000",
  39851=>"010101000",
  39852=>"000011101",
  39853=>"110011000",
  39854=>"000100001",
  39855=>"000010010",
  39856=>"100000000",
  39857=>"011011011",
  39858=>"010010001",
  39859=>"111111110",
  39860=>"010011101",
  39861=>"011001010",
  39862=>"101111011",
  39863=>"101011111",
  39864=>"001111001",
  39865=>"101001011",
  39866=>"111110011",
  39867=>"101100000",
  39868=>"111111110",
  39869=>"000011011",
  39870=>"010111100",
  39871=>"100101000",
  39872=>"000110000",
  39873=>"111000000",
  39874=>"011010111",
  39875=>"000100100",
  39876=>"011101010",
  39877=>"100001101",
  39878=>"110000111",
  39879=>"011010011",
  39880=>"001001000",
  39881=>"010110100",
  39882=>"000101101",
  39883=>"111111111",
  39884=>"000000111",
  39885=>"110000000",
  39886=>"111110101",
  39887=>"010101011",
  39888=>"001001000",
  39889=>"010111000",
  39890=>"111000101",
  39891=>"000000101",
  39892=>"111111111",
  39893=>"101110010",
  39894=>"110010010",
  39895=>"101101011",
  39896=>"000010110",
  39897=>"111000010",
  39898=>"100011110",
  39899=>"001110101",
  39900=>"010010010",
  39901=>"101001011",
  39902=>"011000111",
  39903=>"010010000",
  39904=>"111001001",
  39905=>"110110010",
  39906=>"011001001",
  39907=>"111100000",
  39908=>"101000110",
  39909=>"101101111",
  39910=>"000111101",
  39911=>"010101011",
  39912=>"000101010",
  39913=>"010011010",
  39914=>"011011100",
  39915=>"110000100",
  39916=>"001010110",
  39917=>"101100100",
  39918=>"111101001",
  39919=>"010110001",
  39920=>"000011011",
  39921=>"111011011",
  39922=>"101000011",
  39923=>"011001101",
  39924=>"101000100",
  39925=>"011001100",
  39926=>"011001001",
  39927=>"110100010",
  39928=>"001010111",
  39929=>"111111111",
  39930=>"111011000",
  39931=>"111010001",
  39932=>"101010011",
  39933=>"101001000",
  39934=>"011010010",
  39935=>"010010110",
  39936=>"111100010",
  39937=>"001001110",
  39938=>"010010011",
  39939=>"110010001",
  39940=>"001100100",
  39941=>"010110110",
  39942=>"101101100",
  39943=>"000011101",
  39944=>"101001100",
  39945=>"110111101",
  39946=>"000101101",
  39947=>"100010001",
  39948=>"111001010",
  39949=>"000010010",
  39950=>"011101101",
  39951=>"000001101",
  39952=>"011110110",
  39953=>"000000011",
  39954=>"011100000",
  39955=>"100100001",
  39956=>"010111010",
  39957=>"111111111",
  39958=>"111011101",
  39959=>"111100000",
  39960=>"100101111",
  39961=>"111111000",
  39962=>"011110001",
  39963=>"101000010",
  39964=>"010001111",
  39965=>"000100111",
  39966=>"000110100",
  39967=>"110110011",
  39968=>"110100101",
  39969=>"000001000",
  39970=>"111000110",
  39971=>"110100110",
  39972=>"011111000",
  39973=>"000110101",
  39974=>"000101001",
  39975=>"011101101",
  39976=>"111110110",
  39977=>"000111000",
  39978=>"110110111",
  39979=>"001111000",
  39980=>"001100101",
  39981=>"000100000",
  39982=>"011010011",
  39983=>"000111101",
  39984=>"100111101",
  39985=>"111111101",
  39986=>"100010110",
  39987=>"001101000",
  39988=>"010001001",
  39989=>"000110101",
  39990=>"010011110",
  39991=>"110101010",
  39992=>"001001110",
  39993=>"110110101",
  39994=>"100110110",
  39995=>"110101101",
  39996=>"111110010",
  39997=>"110111000",
  39998=>"100000000",
  39999=>"011101000",
  40000=>"010011111",
  40001=>"011100010",
  40002=>"001101010",
  40003=>"101001011",
  40004=>"000111111",
  40005=>"000101100",
  40006=>"010000000",
  40007=>"110010010",
  40008=>"001000111",
  40009=>"100111000",
  40010=>"000100110",
  40011=>"001110111",
  40012=>"111101101",
  40013=>"001000000",
  40014=>"000111000",
  40015=>"010101001",
  40016=>"010100011",
  40017=>"011101110",
  40018=>"010000110",
  40019=>"000000011",
  40020=>"010100010",
  40021=>"100011100",
  40022=>"001110010",
  40023=>"101001111",
  40024=>"101010001",
  40025=>"101110110",
  40026=>"000000010",
  40027=>"100100000",
  40028=>"111011111",
  40029=>"000011000",
  40030=>"001001001",
  40031=>"100000101",
  40032=>"001001110",
  40033=>"101101000",
  40034=>"000001111",
  40035=>"100110001",
  40036=>"001110110",
  40037=>"011000001",
  40038=>"001001001",
  40039=>"010100000",
  40040=>"011111001",
  40041=>"110111010",
  40042=>"010000011",
  40043=>"101101100",
  40044=>"100000111",
  40045=>"101000100",
  40046=>"110100101",
  40047=>"001111001",
  40048=>"001101000",
  40049=>"111010101",
  40050=>"101011001",
  40051=>"101111111",
  40052=>"001001000",
  40053=>"010101100",
  40054=>"101001110",
  40055=>"101110100",
  40056=>"000001000",
  40057=>"011110110",
  40058=>"010010000",
  40059=>"000000111",
  40060=>"101101100",
  40061=>"110011001",
  40062=>"001000110",
  40063=>"011111111",
  40064=>"100001001",
  40065=>"010101110",
  40066=>"101010100",
  40067=>"001100101",
  40068=>"100101101",
  40069=>"010001010",
  40070=>"000000001",
  40071=>"000001010",
  40072=>"000111010",
  40073=>"110100000",
  40074=>"101011111",
  40075=>"100101100",
  40076=>"100000010",
  40077=>"001101111",
  40078=>"101011000",
  40079=>"101000111",
  40080=>"110001101",
  40081=>"100000110",
  40082=>"100011000",
  40083=>"000100111",
  40084=>"000000111",
  40085=>"100101011",
  40086=>"011010101",
  40087=>"000111000",
  40088=>"011110111",
  40089=>"110110010",
  40090=>"011100000",
  40091=>"000010111",
  40092=>"110011101",
  40093=>"101000000",
  40094=>"011011010",
  40095=>"100001111",
  40096=>"110101000",
  40097=>"011001000",
  40098=>"000101101",
  40099=>"001011101",
  40100=>"000110000",
  40101=>"001000110",
  40102=>"011001111",
  40103=>"010110001",
  40104=>"001100010",
  40105=>"110011110",
  40106=>"111010010",
  40107=>"101101101",
  40108=>"111010111",
  40109=>"000011001",
  40110=>"111111000",
  40111=>"000010101",
  40112=>"010101011",
  40113=>"000111010",
  40114=>"101001001",
  40115=>"101101001",
  40116=>"001011000",
  40117=>"000100000",
  40118=>"011100001",
  40119=>"000000101",
  40120=>"000010001",
  40121=>"010110111",
  40122=>"001101101",
  40123=>"010001001",
  40124=>"110110110",
  40125=>"011111010",
  40126=>"000010011",
  40127=>"000111011",
  40128=>"000011011",
  40129=>"100000010",
  40130=>"110011001",
  40131=>"101011100",
  40132=>"101101100",
  40133=>"111001101",
  40134=>"001000001",
  40135=>"100010011",
  40136=>"001000000",
  40137=>"101000000",
  40138=>"111010000",
  40139=>"100010001",
  40140=>"000110100",
  40141=>"111101011",
  40142=>"101001010",
  40143=>"110001001",
  40144=>"110011101",
  40145=>"100101101",
  40146=>"001000101",
  40147=>"000000001",
  40148=>"000001111",
  40149=>"000001111",
  40150=>"011111011",
  40151=>"101100110",
  40152=>"001110001",
  40153=>"101100110",
  40154=>"000110110",
  40155=>"001100001",
  40156=>"111000010",
  40157=>"010111011",
  40158=>"010110000",
  40159=>"111001010",
  40160=>"110101001",
  40161=>"111100110",
  40162=>"101010101",
  40163=>"110100000",
  40164=>"101100101",
  40165=>"011110011",
  40166=>"100010010",
  40167=>"111110111",
  40168=>"001101010",
  40169=>"000011111",
  40170=>"100010110",
  40171=>"000111110",
  40172=>"101001011",
  40173=>"110111010",
  40174=>"111110011",
  40175=>"000011111",
  40176=>"001000101",
  40177=>"000110001",
  40178=>"011010110",
  40179=>"110101010",
  40180=>"000111101",
  40181=>"100101111",
  40182=>"111100011",
  40183=>"010001010",
  40184=>"011111110",
  40185=>"100011111",
  40186=>"001101011",
  40187=>"100000001",
  40188=>"010101111",
  40189=>"111001110",
  40190=>"100000001",
  40191=>"111001110",
  40192=>"111001111",
  40193=>"101011010",
  40194=>"101011101",
  40195=>"000011011",
  40196=>"011011110",
  40197=>"100011110",
  40198=>"010100000",
  40199=>"110101001",
  40200=>"100010110",
  40201=>"010011100",
  40202=>"011111011",
  40203=>"011101001",
  40204=>"111000000",
  40205=>"001111010",
  40206=>"101001000",
  40207=>"010110011",
  40208=>"111100010",
  40209=>"010000011",
  40210=>"100001010",
  40211=>"100010111",
  40212=>"010001010",
  40213=>"101011010",
  40214=>"010110010",
  40215=>"001100101",
  40216=>"110100000",
  40217=>"110111100",
  40218=>"100010100",
  40219=>"001000000",
  40220=>"111101110",
  40221=>"100100111",
  40222=>"001110001",
  40223=>"101111001",
  40224=>"001010000",
  40225=>"001000001",
  40226=>"001111100",
  40227=>"011001111",
  40228=>"110001010",
  40229=>"000100000",
  40230=>"010110000",
  40231=>"010010101",
  40232=>"001001001",
  40233=>"011011111",
  40234=>"111111110",
  40235=>"000111110",
  40236=>"000011111",
  40237=>"100000111",
  40238=>"011110011",
  40239=>"111110010",
  40240=>"011100000",
  40241=>"100000000",
  40242=>"001011010",
  40243=>"111111010",
  40244=>"001001010",
  40245=>"000010000",
  40246=>"110101101",
  40247=>"111101100",
  40248=>"000000110",
  40249=>"001100101",
  40250=>"010000100",
  40251=>"011110110",
  40252=>"110010101",
  40253=>"010000111",
  40254=>"000000010",
  40255=>"101011101",
  40256=>"000000011",
  40257=>"011111010",
  40258=>"001100101",
  40259=>"110110011",
  40260=>"111000101",
  40261=>"101110101",
  40262=>"111100110",
  40263=>"001111001",
  40264=>"101110111",
  40265=>"000101011",
  40266=>"100001100",
  40267=>"100101100",
  40268=>"110111010",
  40269=>"001110111",
  40270=>"111011111",
  40271=>"000101111",
  40272=>"101101101",
  40273=>"111111110",
  40274=>"001010000",
  40275=>"000001101",
  40276=>"111011100",
  40277=>"000110000",
  40278=>"111101010",
  40279=>"110001001",
  40280=>"111000011",
  40281=>"100110000",
  40282=>"001000101",
  40283=>"011111111",
  40284=>"101111010",
  40285=>"001010000",
  40286=>"101110110",
  40287=>"011000100",
  40288=>"001010001",
  40289=>"111010000",
  40290=>"010101100",
  40291=>"001110101",
  40292=>"100101101",
  40293=>"010000110",
  40294=>"101101111",
  40295=>"111100111",
  40296=>"111010100",
  40297=>"111110010",
  40298=>"000011101",
  40299=>"001111001",
  40300=>"110101101",
  40301=>"010001000",
  40302=>"001100100",
  40303=>"010000000",
  40304=>"010100100",
  40305=>"011010011",
  40306=>"011110110",
  40307=>"100000010",
  40308=>"111001011",
  40309=>"011110110",
  40310=>"111010110",
  40311=>"011100001",
  40312=>"101110011",
  40313=>"010010011",
  40314=>"011011001",
  40315=>"000011100",
  40316=>"101001000",
  40317=>"111111110",
  40318=>"011010011",
  40319=>"100001001",
  40320=>"101101111",
  40321=>"110001001",
  40322=>"101000101",
  40323=>"110000110",
  40324=>"110001101",
  40325=>"001010000",
  40326=>"101010001",
  40327=>"000010000",
  40328=>"110000010",
  40329=>"011101101",
  40330=>"111101000",
  40331=>"101010000",
  40332=>"100111000",
  40333=>"011110000",
  40334=>"111000111",
  40335=>"011100101",
  40336=>"100010101",
  40337=>"000001010",
  40338=>"001011000",
  40339=>"000001100",
  40340=>"110010101",
  40341=>"111111101",
  40342=>"001100000",
  40343=>"010010100",
  40344=>"011001100",
  40345=>"000001000",
  40346=>"110010101",
  40347=>"110100101",
  40348=>"011000101",
  40349=>"010011111",
  40350=>"111101101",
  40351=>"101001000",
  40352=>"011011011",
  40353=>"001100101",
  40354=>"001000000",
  40355=>"010000101",
  40356=>"000011110",
  40357=>"010100100",
  40358=>"111001000",
  40359=>"110011011",
  40360=>"011001100",
  40361=>"010011011",
  40362=>"000010110",
  40363=>"010010001",
  40364=>"011001100",
  40365=>"111111101",
  40366=>"011100001",
  40367=>"110011011",
  40368=>"100000100",
  40369=>"110011110",
  40370=>"111110111",
  40371=>"001100110",
  40372=>"010001111",
  40373=>"000100011",
  40374=>"001110101",
  40375=>"100101110",
  40376=>"001000100",
  40377=>"111000011",
  40378=>"101010000",
  40379=>"010000000",
  40380=>"001111000",
  40381=>"011001011",
  40382=>"110101100",
  40383=>"011011000",
  40384=>"001011000",
  40385=>"001100001",
  40386=>"011001110",
  40387=>"011100100",
  40388=>"011111010",
  40389=>"110010010",
  40390=>"111010100",
  40391=>"100001010",
  40392=>"101010100",
  40393=>"100100110",
  40394=>"001111110",
  40395=>"111111111",
  40396=>"001000111",
  40397=>"011100010",
  40398=>"011001001",
  40399=>"001000010",
  40400=>"000011000",
  40401=>"011111000",
  40402=>"000011111",
  40403=>"111010011",
  40404=>"010001011",
  40405=>"101000010",
  40406=>"010010011",
  40407=>"010000100",
  40408=>"000001100",
  40409=>"010100100",
  40410=>"101011111",
  40411=>"001010110",
  40412=>"110100010",
  40413=>"101100111",
  40414=>"001000011",
  40415=>"011101110",
  40416=>"000010000",
  40417=>"010110110",
  40418=>"110111000",
  40419=>"101000011",
  40420=>"110001000",
  40421=>"110011101",
  40422=>"110011011",
  40423=>"001000010",
  40424=>"101010101",
  40425=>"110111100",
  40426=>"010000111",
  40427=>"011110000",
  40428=>"010001011",
  40429=>"110001000",
  40430=>"111111100",
  40431=>"000000000",
  40432=>"101100111",
  40433=>"110100011",
  40434=>"111111110",
  40435=>"110010110",
  40436=>"011101110",
  40437=>"001010011",
  40438=>"001101001",
  40439=>"000011010",
  40440=>"010010100",
  40441=>"000011101",
  40442=>"101000011",
  40443=>"111110110",
  40444=>"000011111",
  40445=>"011101010",
  40446=>"100011101",
  40447=>"111010101",
  40448=>"001101110",
  40449=>"110001010",
  40450=>"100100100",
  40451=>"000001011",
  40452=>"110100101",
  40453=>"000000000",
  40454=>"111100011",
  40455=>"110011110",
  40456=>"100001010",
  40457=>"111001101",
  40458=>"000100010",
  40459=>"011010001",
  40460=>"000101100",
  40461=>"100001000",
  40462=>"111111111",
  40463=>"111010110",
  40464=>"010001110",
  40465=>"001100110",
  40466=>"110101000",
  40467=>"011110011",
  40468=>"011101001",
  40469=>"101010001",
  40470=>"111101110",
  40471=>"100101011",
  40472=>"000000100",
  40473=>"001110100",
  40474=>"110110101",
  40475=>"010111110",
  40476=>"110001110",
  40477=>"101000100",
  40478=>"011100000",
  40479=>"010011110",
  40480=>"001000000",
  40481=>"001000001",
  40482=>"111110000",
  40483=>"010001101",
  40484=>"011100010",
  40485=>"101110100",
  40486=>"001110001",
  40487=>"000011100",
  40488=>"111011000",
  40489=>"111110001",
  40490=>"010110010",
  40491=>"110000011",
  40492=>"111111000",
  40493=>"111111100",
  40494=>"010001111",
  40495=>"111000011",
  40496=>"101011100",
  40497=>"011000101",
  40498=>"010011100",
  40499=>"111100100",
  40500=>"110000110",
  40501=>"111000000",
  40502=>"010011011",
  40503=>"011011111",
  40504=>"010110011",
  40505=>"101011010",
  40506=>"011101110",
  40507=>"110101011",
  40508=>"010111111",
  40509=>"000110000",
  40510=>"111101011",
  40511=>"010000001",
  40512=>"101000101",
  40513=>"110000000",
  40514=>"000010100",
  40515=>"101101000",
  40516=>"111110001",
  40517=>"000111100",
  40518=>"100000111",
  40519=>"111001101",
  40520=>"001000000",
  40521=>"000011001",
  40522=>"101110000",
  40523=>"101010110",
  40524=>"011010010",
  40525=>"100100000",
  40526=>"010100000",
  40527=>"001100110",
  40528=>"011010110",
  40529=>"111001001",
  40530=>"110100101",
  40531=>"000000000",
  40532=>"111110111",
  40533=>"000001101",
  40534=>"110100010",
  40535=>"000110110",
  40536=>"000011011",
  40537=>"100000101",
  40538=>"000110010",
  40539=>"101101101",
  40540=>"000101011",
  40541=>"101010001",
  40542=>"000100001",
  40543=>"001100001",
  40544=>"000000001",
  40545=>"000001010",
  40546=>"111111110",
  40547=>"010000011",
  40548=>"101001000",
  40549=>"000000110",
  40550=>"001001111",
  40551=>"001111100",
  40552=>"101001011",
  40553=>"101011110",
  40554=>"100000000",
  40555=>"000010000",
  40556=>"001110100",
  40557=>"111101110",
  40558=>"101100001",
  40559=>"010010110",
  40560=>"000010111",
  40561=>"000000101",
  40562=>"110111100",
  40563=>"001001101",
  40564=>"100000100",
  40565=>"101001000",
  40566=>"100001111",
  40567=>"101110000",
  40568=>"001011100",
  40569=>"000100000",
  40570=>"111100001",
  40571=>"000101111",
  40572=>"000111100",
  40573=>"111010011",
  40574=>"010010011",
  40575=>"100001000",
  40576=>"010110000",
  40577=>"111010000",
  40578=>"111010011",
  40579=>"001110001",
  40580=>"001010010",
  40581=>"000110011",
  40582=>"101110001",
  40583=>"000100100",
  40584=>"110000110",
  40585=>"001000111",
  40586=>"101100001",
  40587=>"110110110",
  40588=>"000011001",
  40589=>"111010110",
  40590=>"011100011",
  40591=>"011100011",
  40592=>"111101101",
  40593=>"100001111",
  40594=>"001010100",
  40595=>"000001100",
  40596=>"100010000",
  40597=>"100111010",
  40598=>"111010110",
  40599=>"011001111",
  40600=>"110000001",
  40601=>"011000111",
  40602=>"000000000",
  40603=>"110011111",
  40604=>"110111000",
  40605=>"101001010",
  40606=>"100010011",
  40607=>"000100110",
  40608=>"100110011",
  40609=>"001111010",
  40610=>"010100110",
  40611=>"100100000",
  40612=>"111010110",
  40613=>"010101101",
  40614=>"011010111",
  40615=>"111110100",
  40616=>"111111001",
  40617=>"001100000",
  40618=>"110011101",
  40619=>"001011000",
  40620=>"111111001",
  40621=>"110110010",
  40622=>"011001101",
  40623=>"000111111",
  40624=>"111001111",
  40625=>"110100000",
  40626=>"010001011",
  40627=>"110001100",
  40628=>"111100110",
  40629=>"001000001",
  40630=>"011000011",
  40631=>"110111000",
  40632=>"001100001",
  40633=>"110011010",
  40634=>"101010001",
  40635=>"011011011",
  40636=>"010101111",
  40637=>"100001000",
  40638=>"111010000",
  40639=>"100101101",
  40640=>"101011001",
  40641=>"001010010",
  40642=>"101011010",
  40643=>"110100001",
  40644=>"100110000",
  40645=>"110000110",
  40646=>"011010110",
  40647=>"100010110",
  40648=>"010110011",
  40649=>"100111010",
  40650=>"101001011",
  40651=>"101111000",
  40652=>"010110100",
  40653=>"111010010",
  40654=>"101110000",
  40655=>"000100101",
  40656=>"000001000",
  40657=>"010100100",
  40658=>"100011111",
  40659=>"101100110",
  40660=>"111000011",
  40661=>"000001101",
  40662=>"110011000",
  40663=>"010010000",
  40664=>"011000110",
  40665=>"111101011",
  40666=>"111011100",
  40667=>"100110100",
  40668=>"001010011",
  40669=>"010011011",
  40670=>"111100011",
  40671=>"110110111",
  40672=>"011001010",
  40673=>"000100010",
  40674=>"001010000",
  40675=>"001011011",
  40676=>"101101110",
  40677=>"001000011",
  40678=>"111111001",
  40679=>"100111011",
  40680=>"011001000",
  40681=>"111010010",
  40682=>"000101011",
  40683=>"100100001",
  40684=>"001101100",
  40685=>"010010100",
  40686=>"010100001",
  40687=>"000101111",
  40688=>"011110101",
  40689=>"100011000",
  40690=>"110011111",
  40691=>"000000010",
  40692=>"001000111",
  40693=>"100001011",
  40694=>"000101100",
  40695=>"011100010",
  40696=>"011000100",
  40697=>"110010111",
  40698=>"001111100",
  40699=>"001000001",
  40700=>"010101011",
  40701=>"011000110",
  40702=>"101110110",
  40703=>"000011010",
  40704=>"010011101",
  40705=>"001011100",
  40706=>"001001110",
  40707=>"101000010",
  40708=>"100000000",
  40709=>"101001010",
  40710=>"111011111",
  40711=>"010111001",
  40712=>"111101111",
  40713=>"011110111",
  40714=>"110010111",
  40715=>"000000111",
  40716=>"110001111",
  40717=>"000111001",
  40718=>"000010010",
  40719=>"101101111",
  40720=>"101111101",
  40721=>"111100000",
  40722=>"010001101",
  40723=>"100001000",
  40724=>"001110100",
  40725=>"101011111",
  40726=>"111010110",
  40727=>"110111011",
  40728=>"100101110",
  40729=>"001100101",
  40730=>"000000011",
  40731=>"010100100",
  40732=>"010011011",
  40733=>"101110010",
  40734=>"010110010",
  40735=>"101000111",
  40736=>"100111011",
  40737=>"100000110",
  40738=>"101100000",
  40739=>"010000000",
  40740=>"110110110",
  40741=>"011010100",
  40742=>"111100101",
  40743=>"000111110",
  40744=>"001101011",
  40745=>"010000111",
  40746=>"011101001",
  40747=>"100101001",
  40748=>"111111001",
  40749=>"100100001",
  40750=>"001111010",
  40751=>"101000100",
  40752=>"101001111",
  40753=>"100011001",
  40754=>"001001010",
  40755=>"010101010",
  40756=>"001011111",
  40757=>"100000010",
  40758=>"011001110",
  40759=>"111100011",
  40760=>"110101010",
  40761=>"011001001",
  40762=>"011001000",
  40763=>"011000111",
  40764=>"101100000",
  40765=>"001101000",
  40766=>"100110100",
  40767=>"110100010",
  40768=>"100000011",
  40769=>"101000100",
  40770=>"110001010",
  40771=>"100111011",
  40772=>"010111110",
  40773=>"010010011",
  40774=>"101111110",
  40775=>"000001001",
  40776=>"001000101",
  40777=>"111101001",
  40778=>"110100101",
  40779=>"111010100",
  40780=>"010010001",
  40781=>"001101111",
  40782=>"010110100",
  40783=>"110110000",
  40784=>"100011011",
  40785=>"111111010",
  40786=>"000110110",
  40787=>"010010001",
  40788=>"011101001",
  40789=>"000010111",
  40790=>"000000101",
  40791=>"011110111",
  40792=>"011111001",
  40793=>"000101101",
  40794=>"100100111",
  40795=>"000000100",
  40796=>"100101101",
  40797=>"110110100",
  40798=>"100110011",
  40799=>"100100111",
  40800=>"011101101",
  40801=>"000000011",
  40802=>"101110110",
  40803=>"001100101",
  40804=>"000100010",
  40805=>"000110100",
  40806=>"100001101",
  40807=>"001010011",
  40808=>"001111010",
  40809=>"101000100",
  40810=>"111001100",
  40811=>"000010111",
  40812=>"011101111",
  40813=>"101001001",
  40814=>"001111011",
  40815=>"000001100",
  40816=>"100111100",
  40817=>"000100111",
  40818=>"011101100",
  40819=>"101101010",
  40820=>"101010011",
  40821=>"000010111",
  40822=>"000110011",
  40823=>"110011011",
  40824=>"000101011",
  40825=>"100001110",
  40826=>"010110001",
  40827=>"001110011",
  40828=>"110110100",
  40829=>"010111011",
  40830=>"001001111",
  40831=>"010011001",
  40832=>"101000000",
  40833=>"100000101",
  40834=>"100010110",
  40835=>"000100100",
  40836=>"100000011",
  40837=>"010110010",
  40838=>"101010000",
  40839=>"010010010",
  40840=>"101001010",
  40841=>"110111111",
  40842=>"100000000",
  40843=>"001110001",
  40844=>"010100100",
  40845=>"111110101",
  40846=>"100110110",
  40847=>"100101110",
  40848=>"000000011",
  40849=>"010111010",
  40850=>"001000111",
  40851=>"010001110",
  40852=>"111111110",
  40853=>"011000110",
  40854=>"001011011",
  40855=>"010011001",
  40856=>"110010000",
  40857=>"010110011",
  40858=>"000100011",
  40859=>"111000110",
  40860=>"011101110",
  40861=>"001101110",
  40862=>"101101100",
  40863=>"110000111",
  40864=>"000001011",
  40865=>"110101000",
  40866=>"111100000",
  40867=>"100001111",
  40868=>"101111100",
  40869=>"000010111",
  40870=>"010100110",
  40871=>"110001110",
  40872=>"001011000",
  40873=>"000100011",
  40874=>"110110001",
  40875=>"101111101",
  40876=>"010001100",
  40877=>"100101011",
  40878=>"001100111",
  40879=>"000000110",
  40880=>"100101011",
  40881=>"101101101",
  40882=>"110100101",
  40883=>"100001001",
  40884=>"001101110",
  40885=>"100100110",
  40886=>"001100101",
  40887=>"111011110",
  40888=>"101000110",
  40889=>"001100010",
  40890=>"110011100",
  40891=>"111110000",
  40892=>"101101110",
  40893=>"000111100",
  40894=>"111111110",
  40895=>"110101011",
  40896=>"001110110",
  40897=>"000010111",
  40898=>"000001100",
  40899=>"110100010",
  40900=>"011101101",
  40901=>"110100111",
  40902=>"111101111",
  40903=>"001010100",
  40904=>"010110000",
  40905=>"100001010",
  40906=>"001010110",
  40907=>"101010011",
  40908=>"010111111",
  40909=>"110100101",
  40910=>"100001101",
  40911=>"110111011",
  40912=>"011100011",
  40913=>"001010100",
  40914=>"111010010",
  40915=>"000100000",
  40916=>"010101000",
  40917=>"101000110",
  40918=>"101011110",
  40919=>"011001101",
  40920=>"110110110",
  40921=>"010011010",
  40922=>"111011110",
  40923=>"000111111",
  40924=>"000100100",
  40925=>"010011110",
  40926=>"000101101",
  40927=>"010011101",
  40928=>"101110111",
  40929=>"001010001",
  40930=>"111001110",
  40931=>"001001110",
  40932=>"100101000",
  40933=>"111010111",
  40934=>"010111100",
  40935=>"010101000",
  40936=>"100000100",
  40937=>"100111011",
  40938=>"101111110",
  40939=>"010011110",
  40940=>"101011101",
  40941=>"110001101",
  40942=>"011001110",
  40943=>"110110000",
  40944=>"110010001",
  40945=>"110110010",
  40946=>"100011000",
  40947=>"010100011",
  40948=>"101110110",
  40949=>"011111101",
  40950=>"001110111",
  40951=>"001111101",
  40952=>"111001011",
  40953=>"011101110",
  40954=>"011111011",
  40955=>"011100100",
  40956=>"111110100",
  40957=>"001100010",
  40958=>"000000100",
  40959=>"001100011",
  40960=>"110010100",
  40961=>"010101010",
  40962=>"001011111",
  40963=>"001011001",
  40964=>"101001100",
  40965=>"011010111",
  40966=>"011111111",
  40967=>"101000001",
  40968=>"111100011",
  40969=>"111111000",
  40970=>"010001111",
  40971=>"000100100",
  40972=>"110111100",
  40973=>"010110011",
  40974=>"111010100",
  40975=>"101001010",
  40976=>"110011001",
  40977=>"110000011",
  40978=>"010101001",
  40979=>"100110010",
  40980=>"101010110",
  40981=>"110100010",
  40982=>"100101000",
  40983=>"001000111",
  40984=>"111001101",
  40985=>"101011000",
  40986=>"100010001",
  40987=>"010011101",
  40988=>"101011101",
  40989=>"100000001",
  40990=>"111101101",
  40991=>"000010011",
  40992=>"011010010",
  40993=>"101101111",
  40994=>"110010001",
  40995=>"101011011",
  40996=>"000011011",
  40997=>"101110110",
  40998=>"000010111",
  40999=>"111010110",
  41000=>"011011000",
  41001=>"000000101",
  41002=>"001100000",
  41003=>"100111011",
  41004=>"010000111",
  41005=>"010011100",
  41006=>"011101101",
  41007=>"100000111",
  41008=>"010111010",
  41009=>"011011010",
  41010=>"010101010",
  41011=>"101010110",
  41012=>"111001111",
  41013=>"100100001",
  41014=>"111101111",
  41015=>"001001000",
  41016=>"000110011",
  41017=>"010111010",
  41018=>"101110000",
  41019=>"001001001",
  41020=>"100000000",
  41021=>"101100100",
  41022=>"111010111",
  41023=>"001010000",
  41024=>"100100000",
  41025=>"001011100",
  41026=>"001110110",
  41027=>"100000111",
  41028=>"000110010",
  41029=>"110110101",
  41030=>"001011011",
  41031=>"111010001",
  41032=>"011000101",
  41033=>"101101000",
  41034=>"000001011",
  41035=>"001110001",
  41036=>"111110011",
  41037=>"101000110",
  41038=>"110110111",
  41039=>"101111110",
  41040=>"111001100",
  41041=>"110011011",
  41042=>"100100110",
  41043=>"011000001",
  41044=>"110111101",
  41045=>"110001000",
  41046=>"100011101",
  41047=>"110000011",
  41048=>"111100011",
  41049=>"100011010",
  41050=>"110100100",
  41051=>"100100101",
  41052=>"000000000",
  41053=>"001001110",
  41054=>"011110011",
  41055=>"001111101",
  41056=>"010011001",
  41057=>"011000111",
  41058=>"010001111",
  41059=>"110101100",
  41060=>"000100011",
  41061=>"100100001",
  41062=>"000010010",
  41063=>"100010111",
  41064=>"100011111",
  41065=>"011111011",
  41066=>"000111010",
  41067=>"000101110",
  41068=>"011101111",
  41069=>"101001111",
  41070=>"010011110",
  41071=>"000001010",
  41072=>"010100100",
  41073=>"000100000",
  41074=>"101000010",
  41075=>"011010010",
  41076=>"001111010",
  41077=>"111111111",
  41078=>"111111110",
  41079=>"101010111",
  41080=>"100111000",
  41081=>"011010110",
  41082=>"000001000",
  41083=>"011010001",
  41084=>"011011111",
  41085=>"000011101",
  41086=>"011000000",
  41087=>"111110110",
  41088=>"110111011",
  41089=>"100101001",
  41090=>"010001100",
  41091=>"110011011",
  41092=>"110100100",
  41093=>"101100111",
  41094=>"001101011",
  41095=>"100101000",
  41096=>"000111001",
  41097=>"011111100",
  41098=>"001000101",
  41099=>"101111100",
  41100=>"011011110",
  41101=>"100111001",
  41102=>"100010101",
  41103=>"111011101",
  41104=>"010001000",
  41105=>"111010011",
  41106=>"110001001",
  41107=>"101001110",
  41108=>"101010001",
  41109=>"000011001",
  41110=>"000000011",
  41111=>"111111011",
  41112=>"111000100",
  41113=>"010011111",
  41114=>"101111010",
  41115=>"000110100",
  41116=>"110011001",
  41117=>"111111101",
  41118=>"000100010",
  41119=>"000001101",
  41120=>"111010011",
  41121=>"110000110",
  41122=>"000000110",
  41123=>"001001111",
  41124=>"010110110",
  41125=>"100111111",
  41126=>"000111010",
  41127=>"011100001",
  41128=>"111100000",
  41129=>"110010101",
  41130=>"111010010",
  41131=>"010000001",
  41132=>"001101100",
  41133=>"111110010",
  41134=>"010001111",
  41135=>"010111101",
  41136=>"111001100",
  41137=>"000001101",
  41138=>"100100100",
  41139=>"010110101",
  41140=>"111101100",
  41141=>"000000001",
  41142=>"111111010",
  41143=>"000110110",
  41144=>"110100011",
  41145=>"101011010",
  41146=>"010101001",
  41147=>"110001001",
  41148=>"000000000",
  41149=>"111011001",
  41150=>"111001000",
  41151=>"010011000",
  41152=>"110001111",
  41153=>"100000010",
  41154=>"101100000",
  41155=>"110011110",
  41156=>"000000001",
  41157=>"010110011",
  41158=>"000101100",
  41159=>"110001010",
  41160=>"111001100",
  41161=>"011000011",
  41162=>"110011010",
  41163=>"011011001",
  41164=>"110101100",
  41165=>"110110101",
  41166=>"100110011",
  41167=>"110111010",
  41168=>"001001010",
  41169=>"000101010",
  41170=>"101101100",
  41171=>"101100110",
  41172=>"010001101",
  41173=>"001001010",
  41174=>"000000001",
  41175=>"010101101",
  41176=>"011000111",
  41177=>"110111001",
  41178=>"100001111",
  41179=>"110110110",
  41180=>"111001100",
  41181=>"100110101",
  41182=>"011000010",
  41183=>"110001111",
  41184=>"011001111",
  41185=>"001100011",
  41186=>"101100101",
  41187=>"101110101",
  41188=>"010000101",
  41189=>"011001000",
  41190=>"100010001",
  41191=>"100010011",
  41192=>"111110001",
  41193=>"101111100",
  41194=>"100001000",
  41195=>"110000101",
  41196=>"001010101",
  41197=>"111010110",
  41198=>"011111010",
  41199=>"111001000",
  41200=>"011011011",
  41201=>"001111010",
  41202=>"001101011",
  41203=>"101111110",
  41204=>"010011101",
  41205=>"100101111",
  41206=>"000011010",
  41207=>"100001000",
  41208=>"001110010",
  41209=>"110100001",
  41210=>"011001000",
  41211=>"011111111",
  41212=>"100001011",
  41213=>"000001010",
  41214=>"111111001",
  41215=>"110010110",
  41216=>"000010101",
  41217=>"100110010",
  41218=>"101000010",
  41219=>"000110001",
  41220=>"011000001",
  41221=>"101111111",
  41222=>"001001000",
  41223=>"100010011",
  41224=>"001011111",
  41225=>"101101010",
  41226=>"000011111",
  41227=>"010110100",
  41228=>"111110011",
  41229=>"110110000",
  41230=>"101001101",
  41231=>"011011100",
  41232=>"001101111",
  41233=>"000000001",
  41234=>"101001001",
  41235=>"101000110",
  41236=>"110110100",
  41237=>"101101110",
  41238=>"010001100",
  41239=>"100001011",
  41240=>"100000110",
  41241=>"101011110",
  41242=>"111110110",
  41243=>"100111110",
  41244=>"010110110",
  41245=>"000001101",
  41246=>"100000110",
  41247=>"011000010",
  41248=>"101001001",
  41249=>"000000100",
  41250=>"010010000",
  41251=>"001101000",
  41252=>"001101011",
  41253=>"010101101",
  41254=>"011010111",
  41255=>"111000101",
  41256=>"001000001",
  41257=>"001100101",
  41258=>"000111110",
  41259=>"110100011",
  41260=>"000100100",
  41261=>"000100111",
  41262=>"000000100",
  41263=>"011011000",
  41264=>"011111001",
  41265=>"011000011",
  41266=>"111111000",
  41267=>"000110100",
  41268=>"001011010",
  41269=>"000011111",
  41270=>"111000100",
  41271=>"010111101",
  41272=>"101110110",
  41273=>"001101100",
  41274=>"110001011",
  41275=>"000010000",
  41276=>"100010100",
  41277=>"000000101",
  41278=>"110001011",
  41279=>"100110011",
  41280=>"010001001",
  41281=>"001111001",
  41282=>"011111111",
  41283=>"011000100",
  41284=>"001100111",
  41285=>"100000000",
  41286=>"001100111",
  41287=>"000001001",
  41288=>"001010011",
  41289=>"011011000",
  41290=>"010110111",
  41291=>"010011001",
  41292=>"000101011",
  41293=>"000100011",
  41294=>"011000110",
  41295=>"001100100",
  41296=>"111000010",
  41297=>"110011010",
  41298=>"100000100",
  41299=>"101000010",
  41300=>"000010001",
  41301=>"100111100",
  41302=>"111010110",
  41303=>"111010001",
  41304=>"010100010",
  41305=>"100100001",
  41306=>"101100100",
  41307=>"100000100",
  41308=>"000011111",
  41309=>"010000101",
  41310=>"011000111",
  41311=>"000010100",
  41312=>"110110111",
  41313=>"011011101",
  41314=>"011110100",
  41315=>"000100110",
  41316=>"110011001",
  41317=>"111101111",
  41318=>"011000111",
  41319=>"110001011",
  41320=>"101001001",
  41321=>"111001001",
  41322=>"010110110",
  41323=>"000111100",
  41324=>"100010000",
  41325=>"101001110",
  41326=>"001000100",
  41327=>"101111011",
  41328=>"001010100",
  41329=>"010010001",
  41330=>"010000001",
  41331=>"011101101",
  41332=>"011001111",
  41333=>"101101110",
  41334=>"010010110",
  41335=>"110110001",
  41336=>"000111111",
  41337=>"000110010",
  41338=>"001001110",
  41339=>"001101001",
  41340=>"100011100",
  41341=>"001000011",
  41342=>"110011100",
  41343=>"111001111",
  41344=>"001000011",
  41345=>"000011001",
  41346=>"001010100",
  41347=>"111000101",
  41348=>"110000010",
  41349=>"100000000",
  41350=>"111000000",
  41351=>"001001010",
  41352=>"111011100",
  41353=>"011010010",
  41354=>"100011111",
  41355=>"000100001",
  41356=>"001010010",
  41357=>"000000011",
  41358=>"110010110",
  41359=>"101110011",
  41360=>"101000011",
  41361=>"001010001",
  41362=>"100000111",
  41363=>"111111110",
  41364=>"111000001",
  41365=>"010111011",
  41366=>"010011011",
  41367=>"100100000",
  41368=>"111101100",
  41369=>"000110111",
  41370=>"111000110",
  41371=>"101010001",
  41372=>"111000010",
  41373=>"011010011",
  41374=>"010100111",
  41375=>"011101100",
  41376=>"010001010",
  41377=>"010011000",
  41378=>"101000001",
  41379=>"000001000",
  41380=>"011100000",
  41381=>"010010111",
  41382=>"011001000",
  41383=>"010111010",
  41384=>"010010100",
  41385=>"000000110",
  41386=>"100100001",
  41387=>"101011100",
  41388=>"000110111",
  41389=>"110001000",
  41390=>"010000010",
  41391=>"100001110",
  41392=>"010001101",
  41393=>"011001010",
  41394=>"101111000",
  41395=>"110011110",
  41396=>"101100101",
  41397=>"101101101",
  41398=>"101001010",
  41399=>"000110011",
  41400=>"111110000",
  41401=>"000011011",
  41402=>"101011100",
  41403=>"100111000",
  41404=>"111010011",
  41405=>"001010101",
  41406=>"000000000",
  41407=>"001100100",
  41408=>"110010110",
  41409=>"110101100",
  41410=>"010111011",
  41411=>"010001011",
  41412=>"001000001",
  41413=>"011000111",
  41414=>"010011101",
  41415=>"010000001",
  41416=>"101001011",
  41417=>"001100101",
  41418=>"110001110",
  41419=>"011011010",
  41420=>"111101001",
  41421=>"101111111",
  41422=>"000110111",
  41423=>"011011010",
  41424=>"101111001",
  41425=>"101110011",
  41426=>"000000011",
  41427=>"101111011",
  41428=>"001010111",
  41429=>"101001100",
  41430=>"110100001",
  41431=>"011101101",
  41432=>"100101011",
  41433=>"100100101",
  41434=>"111111101",
  41435=>"000010000",
  41436=>"010101100",
  41437=>"001000011",
  41438=>"110100100",
  41439=>"111110001",
  41440=>"101011111",
  41441=>"111110100",
  41442=>"101010111",
  41443=>"111110011",
  41444=>"011101111",
  41445=>"011110011",
  41446=>"001010111",
  41447=>"001001110",
  41448=>"110011010",
  41449=>"001100100",
  41450=>"000010011",
  41451=>"011100110",
  41452=>"000110001",
  41453=>"000100000",
  41454=>"111101011",
  41455=>"110110000",
  41456=>"001101100",
  41457=>"001101111",
  41458=>"011000001",
  41459=>"101010100",
  41460=>"100111110",
  41461=>"001001110",
  41462=>"100101100",
  41463=>"111001100",
  41464=>"100100100",
  41465=>"101001110",
  41466=>"111010101",
  41467=>"101011011",
  41468=>"100110101",
  41469=>"001110000",
  41470=>"100000100",
  41471=>"101000101",
  41472=>"000111100",
  41473=>"110001011",
  41474=>"111110001",
  41475=>"110101100",
  41476=>"011110011",
  41477=>"101011000",
  41478=>"111100011",
  41479=>"111011000",
  41480=>"000000111",
  41481=>"010010101",
  41482=>"011110110",
  41483=>"011100110",
  41484=>"101101111",
  41485=>"111100001",
  41486=>"111001011",
  41487=>"011111110",
  41488=>"001111101",
  41489=>"011011111",
  41490=>"011000011",
  41491=>"101101100",
  41492=>"001101000",
  41493=>"100110000",
  41494=>"100111010",
  41495=>"100010101",
  41496=>"010110011",
  41497=>"011100011",
  41498=>"111110011",
  41499=>"100110110",
  41500=>"111101100",
  41501=>"110111100",
  41502=>"111100000",
  41503=>"010110011",
  41504=>"001001000",
  41505=>"111101101",
  41506=>"100000001",
  41507=>"011111110",
  41508=>"000101100",
  41509=>"110010111",
  41510=>"101111000",
  41511=>"101111000",
  41512=>"101101000",
  41513=>"000000000",
  41514=>"101101100",
  41515=>"101001111",
  41516=>"000001011",
  41517=>"110100000",
  41518=>"000001101",
  41519=>"111111100",
  41520=>"110110101",
  41521=>"111010100",
  41522=>"100010100",
  41523=>"100001011",
  41524=>"001110100",
  41525=>"111001001",
  41526=>"100101001",
  41527=>"000100000",
  41528=>"111010111",
  41529=>"001010110",
  41530=>"110001010",
  41531=>"001101100",
  41532=>"001111100",
  41533=>"100111011",
  41534=>"000000100",
  41535=>"101001011",
  41536=>"110000101",
  41537=>"001100110",
  41538=>"010000111",
  41539=>"110011000",
  41540=>"110111111",
  41541=>"001000011",
  41542=>"110101010",
  41543=>"100100110",
  41544=>"001001000",
  41545=>"111101100",
  41546=>"010100011",
  41547=>"010101001",
  41548=>"011100100",
  41549=>"011000001",
  41550=>"100010000",
  41551=>"110100110",
  41552=>"000000101",
  41553=>"011100010",
  41554=>"001000100",
  41555=>"100000000",
  41556=>"101000010",
  41557=>"111101001",
  41558=>"001000001",
  41559=>"011111000",
  41560=>"001101011",
  41561=>"000010010",
  41562=>"011000010",
  41563=>"000010110",
  41564=>"100000101",
  41565=>"000000001",
  41566=>"001011101",
  41567=>"110001110",
  41568=>"111110001",
  41569=>"101110001",
  41570=>"010011110",
  41571=>"011001010",
  41572=>"110110110",
  41573=>"001111000",
  41574=>"110111101",
  41575=>"000010000",
  41576=>"001010100",
  41577=>"110001001",
  41578=>"101001011",
  41579=>"100101001",
  41580=>"001100001",
  41581=>"110100011",
  41582=>"000111001",
  41583=>"010100100",
  41584=>"100101100",
  41585=>"000110011",
  41586=>"111010000",
  41587=>"111000001",
  41588=>"001110111",
  41589=>"100000010",
  41590=>"111111010",
  41591=>"110000001",
  41592=>"010111100",
  41593=>"100001010",
  41594=>"111111010",
  41595=>"110011010",
  41596=>"100101010",
  41597=>"111011100",
  41598=>"101111011",
  41599=>"111011110",
  41600=>"111111110",
  41601=>"001011111",
  41602=>"110011100",
  41603=>"110101110",
  41604=>"001000000",
  41605=>"001101000",
  41606=>"100000000",
  41607=>"111111000",
  41608=>"011110011",
  41609=>"100010100",
  41610=>"011010100",
  41611=>"111010100",
  41612=>"001101101",
  41613=>"001100010",
  41614=>"111101001",
  41615=>"101110111",
  41616=>"010011010",
  41617=>"111100001",
  41618=>"101000010",
  41619=>"001011111",
  41620=>"010001100",
  41621=>"011101110",
  41622=>"010011001",
  41623=>"111010011",
  41624=>"010100010",
  41625=>"101000010",
  41626=>"100011101",
  41627=>"000100010",
  41628=>"100101100",
  41629=>"000110100",
  41630=>"100010011",
  41631=>"111001011",
  41632=>"010010000",
  41633=>"100111000",
  41634=>"110001100",
  41635=>"010011010",
  41636=>"001011011",
  41637=>"010101110",
  41638=>"000011111",
  41639=>"101111000",
  41640=>"010111010",
  41641=>"000011000",
  41642=>"010001000",
  41643=>"010010011",
  41644=>"101100000",
  41645=>"110000100",
  41646=>"111110000",
  41647=>"110100000",
  41648=>"001101111",
  41649=>"000000011",
  41650=>"000001010",
  41651=>"110001101",
  41652=>"011010100",
  41653=>"101110100",
  41654=>"010100100",
  41655=>"101010110",
  41656=>"001000010",
  41657=>"010101010",
  41658=>"011101010",
  41659=>"100011111",
  41660=>"011000100",
  41661=>"100011101",
  41662=>"001110100",
  41663=>"101001011",
  41664=>"011100000",
  41665=>"010101001",
  41666=>"011101010",
  41667=>"111110001",
  41668=>"000110001",
  41669=>"000110101",
  41670=>"100101111",
  41671=>"000010010",
  41672=>"010101000",
  41673=>"110001101",
  41674=>"011111000",
  41675=>"001111100",
  41676=>"110100101",
  41677=>"011101011",
  41678=>"001111100",
  41679=>"001010000",
  41680=>"111001001",
  41681=>"001011100",
  41682=>"001110101",
  41683=>"110100111",
  41684=>"011110111",
  41685=>"001100010",
  41686=>"100110111",
  41687=>"000000001",
  41688=>"001000000",
  41689=>"110101011",
  41690=>"110101011",
  41691=>"101001110",
  41692=>"010111000",
  41693=>"010100000",
  41694=>"010100000",
  41695=>"000101111",
  41696=>"101101000",
  41697=>"010011000",
  41698=>"010111000",
  41699=>"001010011",
  41700=>"110111000",
  41701=>"011010111",
  41702=>"110110100",
  41703=>"111101100",
  41704=>"010110000",
  41705=>"011101011",
  41706=>"110011100",
  41707=>"111101111",
  41708=>"110010010",
  41709=>"000011110",
  41710=>"111100100",
  41711=>"010100001",
  41712=>"111011101",
  41713=>"010100001",
  41714=>"110000001",
  41715=>"001000100",
  41716=>"010001010",
  41717=>"100010110",
  41718=>"100011111",
  41719=>"010001001",
  41720=>"001000110",
  41721=>"101100001",
  41722=>"000101101",
  41723=>"110111101",
  41724=>"111110110",
  41725=>"111010111",
  41726=>"110101101",
  41727=>"010000101",
  41728=>"010010000",
  41729=>"010101000",
  41730=>"010001010",
  41731=>"001000110",
  41732=>"010000011",
  41733=>"001001000",
  41734=>"101100101",
  41735=>"000000100",
  41736=>"110100110",
  41737=>"001110110",
  41738=>"101011111",
  41739=>"110001001",
  41740=>"111001111",
  41741=>"010001100",
  41742=>"000010001",
  41743=>"101100001",
  41744=>"000101010",
  41745=>"000110010",
  41746=>"000101010",
  41747=>"101000100",
  41748=>"100111001",
  41749=>"110010011",
  41750=>"011101010",
  41751=>"011100101",
  41752=>"100001101",
  41753=>"010101010",
  41754=>"010000111",
  41755=>"111000100",
  41756=>"110011101",
  41757=>"101000000",
  41758=>"000011001",
  41759=>"000010111",
  41760=>"000011011",
  41761=>"010000010",
  41762=>"011011011",
  41763=>"100010111",
  41764=>"001110011",
  41765=>"101100100",
  41766=>"011010001",
  41767=>"111011010",
  41768=>"010100101",
  41769=>"011001010",
  41770=>"100111100",
  41771=>"101111000",
  41772=>"000010011",
  41773=>"000111010",
  41774=>"100010011",
  41775=>"010000000",
  41776=>"101010100",
  41777=>"011001011",
  41778=>"100110010",
  41779=>"100111110",
  41780=>"101110011",
  41781=>"001000101",
  41782=>"101001110",
  41783=>"000100100",
  41784=>"010001101",
  41785=>"000101000",
  41786=>"000101111",
  41787=>"100101001",
  41788=>"100101101",
  41789=>"000110001",
  41790=>"101011000",
  41791=>"010011100",
  41792=>"001111110",
  41793=>"010100111",
  41794=>"000010101",
  41795=>"011110011",
  41796=>"110111000",
  41797=>"111100001",
  41798=>"011000010",
  41799=>"000011110",
  41800=>"001010000",
  41801=>"001100111",
  41802=>"001111111",
  41803=>"001011101",
  41804=>"001111010",
  41805=>"111110001",
  41806=>"111000100",
  41807=>"100010111",
  41808=>"010111100",
  41809=>"101101111",
  41810=>"010001110",
  41811=>"101010100",
  41812=>"101010110",
  41813=>"101110011",
  41814=>"110010100",
  41815=>"000011010",
  41816=>"011011101",
  41817=>"010000111",
  41818=>"111011111",
  41819=>"001101110",
  41820=>"110000101",
  41821=>"110111111",
  41822=>"000100011",
  41823=>"110101011",
  41824=>"000100010",
  41825=>"111010011",
  41826=>"001001100",
  41827=>"100011111",
  41828=>"101100110",
  41829=>"001010000",
  41830=>"010001101",
  41831=>"111111110",
  41832=>"111101111",
  41833=>"011011100",
  41834=>"010111001",
  41835=>"001000100",
  41836=>"111111001",
  41837=>"111101011",
  41838=>"101100010",
  41839=>"000100010",
  41840=>"001100111",
  41841=>"101111110",
  41842=>"111110010",
  41843=>"010000100",
  41844=>"100110000",
  41845=>"001111010",
  41846=>"011001111",
  41847=>"111001101",
  41848=>"111010101",
  41849=>"001011111",
  41850=>"111101011",
  41851=>"001100100",
  41852=>"100001000",
  41853=>"100101010",
  41854=>"110100010",
  41855=>"100010001",
  41856=>"001100010",
  41857=>"001101111",
  41858=>"000100001",
  41859=>"000011010",
  41860=>"011011100",
  41861=>"111000000",
  41862=>"010001001",
  41863=>"010011001",
  41864=>"001011000",
  41865=>"001000001",
  41866=>"101010100",
  41867=>"000000011",
  41868=>"111011101",
  41869=>"100001010",
  41870=>"000011010",
  41871=>"111011111",
  41872=>"101001110",
  41873=>"011010101",
  41874=>"111100001",
  41875=>"101111001",
  41876=>"010011001",
  41877=>"101111011",
  41878=>"001011100",
  41879=>"010010100",
  41880=>"110001010",
  41881=>"111000111",
  41882=>"000111001",
  41883=>"010011110",
  41884=>"011111100",
  41885=>"100000100",
  41886=>"001011000",
  41887=>"010000111",
  41888=>"101100101",
  41889=>"111010101",
  41890=>"010010000",
  41891=>"110101111",
  41892=>"110000000",
  41893=>"000001001",
  41894=>"101101001",
  41895=>"000110100",
  41896=>"011011010",
  41897=>"100010011",
  41898=>"110000100",
  41899=>"100010110",
  41900=>"001010100",
  41901=>"001101101",
  41902=>"100111000",
  41903=>"111101111",
  41904=>"110111101",
  41905=>"000000100",
  41906=>"010000000",
  41907=>"110111111",
  41908=>"011000011",
  41909=>"100101010",
  41910=>"010010100",
  41911=>"010101101",
  41912=>"110000111",
  41913=>"000001110",
  41914=>"101011001",
  41915=>"111000101",
  41916=>"110010101",
  41917=>"011110111",
  41918=>"011110101",
  41919=>"011110000",
  41920=>"001011111",
  41921=>"100000011",
  41922=>"011011001",
  41923=>"110100001",
  41924=>"010110100",
  41925=>"001110110",
  41926=>"111000000",
  41927=>"110010100",
  41928=>"100111100",
  41929=>"000010101",
  41930=>"101011100",
  41931=>"001000101",
  41932=>"010100000",
  41933=>"010011101",
  41934=>"010110111",
  41935=>"111110110",
  41936=>"001111110",
  41937=>"110000011",
  41938=>"011100010",
  41939=>"010000101",
  41940=>"101110100",
  41941=>"111110110",
  41942=>"011110110",
  41943=>"001100110",
  41944=>"100000010",
  41945=>"001000000",
  41946=>"001100000",
  41947=>"011011100",
  41948=>"001001100",
  41949=>"001001011",
  41950=>"100011010",
  41951=>"001010010",
  41952=>"110001111",
  41953=>"011001000",
  41954=>"010111001",
  41955=>"000000000",
  41956=>"001010111",
  41957=>"100011111",
  41958=>"010100001",
  41959=>"010000101",
  41960=>"001100101",
  41961=>"111111110",
  41962=>"111010011",
  41963=>"111011011",
  41964=>"000100110",
  41965=>"111110010",
  41966=>"000111101",
  41967=>"100111101",
  41968=>"100111101",
  41969=>"000010110",
  41970=>"100001111",
  41971=>"010010011",
  41972=>"110010001",
  41973=>"001010100",
  41974=>"100111101",
  41975=>"110100101",
  41976=>"110110100",
  41977=>"101111111",
  41978=>"100011100",
  41979=>"111110100",
  41980=>"010000010",
  41981=>"111101111",
  41982=>"111011100",
  41983=>"000000100",
  41984=>"110111100",
  41985=>"101111010",
  41986=>"011111001",
  41987=>"000000100",
  41988=>"001101001",
  41989=>"111010101",
  41990=>"001010101",
  41991=>"100011011",
  41992=>"010111011",
  41993=>"110111101",
  41994=>"111011010",
  41995=>"000000101",
  41996=>"110001111",
  41997=>"010100111",
  41998=>"011101010",
  41999=>"000100010",
  42000=>"000010010",
  42001=>"001001100",
  42002=>"001000101",
  42003=>"010000000",
  42004=>"011100000",
  42005=>"111111100",
  42006=>"010110110",
  42007=>"111101111",
  42008=>"110101101",
  42009=>"111111000",
  42010=>"010100110",
  42011=>"010011110",
  42012=>"010101111",
  42013=>"101100000",
  42014=>"011001010",
  42015=>"000001100",
  42016=>"000010010",
  42017=>"010010001",
  42018=>"111101110",
  42019=>"101011011",
  42020=>"010110111",
  42021=>"011101101",
  42022=>"001001001",
  42023=>"100011010",
  42024=>"101000001",
  42025=>"001011001",
  42026=>"001000010",
  42027=>"101111000",
  42028=>"111010110",
  42029=>"100110110",
  42030=>"111101001",
  42031=>"001100000",
  42032=>"001010101",
  42033=>"110000001",
  42034=>"111000010",
  42035=>"101101011",
  42036=>"011001110",
  42037=>"111110001",
  42038=>"111001010",
  42039=>"101010000",
  42040=>"011011011",
  42041=>"111111000",
  42042=>"001000000",
  42043=>"101001110",
  42044=>"111101111",
  42045=>"101101101",
  42046=>"011001011",
  42047=>"000100000",
  42048=>"010010111",
  42049=>"110010010",
  42050=>"101010110",
  42051=>"101001010",
  42052=>"111111110",
  42053=>"111100011",
  42054=>"111001110",
  42055=>"101110110",
  42056=>"011100011",
  42057=>"000011100",
  42058=>"001111011",
  42059=>"000100000",
  42060=>"111000100",
  42061=>"100110101",
  42062=>"111001100",
  42063=>"111100111",
  42064=>"000000000",
  42065=>"110000001",
  42066=>"000111111",
  42067=>"111110100",
  42068=>"010010100",
  42069=>"011010001",
  42070=>"101011010",
  42071=>"010001000",
  42072=>"101110110",
  42073=>"011111001",
  42074=>"100000110",
  42075=>"001101000",
  42076=>"111111100",
  42077=>"010110100",
  42078=>"010000011",
  42079=>"001011011",
  42080=>"001000011",
  42081=>"110000010",
  42082=>"000101111",
  42083=>"000100010",
  42084=>"101010011",
  42085=>"011100010",
  42086=>"111111110",
  42087=>"100000111",
  42088=>"001101101",
  42089=>"101000011",
  42090=>"001100101",
  42091=>"101100100",
  42092=>"010110010",
  42093=>"111110001",
  42094=>"000000111",
  42095=>"000101001",
  42096=>"010001011",
  42097=>"010100000",
  42098=>"001010011",
  42099=>"010001011",
  42100=>"010010010",
  42101=>"001011000",
  42102=>"100011011",
  42103=>"001110010",
  42104=>"010100111",
  42105=>"011100110",
  42106=>"101000100",
  42107=>"011001011",
  42108=>"110010001",
  42109=>"111110111",
  42110=>"011011011",
  42111=>"101010101",
  42112=>"101001000",
  42113=>"000101110",
  42114=>"010000010",
  42115=>"000111111",
  42116=>"100010011",
  42117=>"100001110",
  42118=>"010000001",
  42119=>"001010101",
  42120=>"100001111",
  42121=>"001101111",
  42122=>"001001010",
  42123=>"010011010",
  42124=>"111110001",
  42125=>"000110111",
  42126=>"000110011",
  42127=>"011010011",
  42128=>"000101001",
  42129=>"111011110",
  42130=>"000010100",
  42131=>"100100001",
  42132=>"001100000",
  42133=>"000010100",
  42134=>"010110011",
  42135=>"000101110",
  42136=>"011001100",
  42137=>"000000000",
  42138=>"100010110",
  42139=>"011011011",
  42140=>"111111110",
  42141=>"011110011",
  42142=>"100111000",
  42143=>"111100011",
  42144=>"011100001",
  42145=>"001110000",
  42146=>"110000111",
  42147=>"101100110",
  42148=>"101111001",
  42149=>"000111010",
  42150=>"010010001",
  42151=>"000011010",
  42152=>"001110111",
  42153=>"111001110",
  42154=>"110010110",
  42155=>"111101111",
  42156=>"010111101",
  42157=>"001000011",
  42158=>"001110111",
  42159=>"101001101",
  42160=>"000011011",
  42161=>"001010100",
  42162=>"001010101",
  42163=>"010000000",
  42164=>"100000100",
  42165=>"001011111",
  42166=>"001010010",
  42167=>"110100011",
  42168=>"110110011",
  42169=>"111000100",
  42170=>"000010010",
  42171=>"101010010",
  42172=>"110110000",
  42173=>"111101001",
  42174=>"011101010",
  42175=>"110111101",
  42176=>"011101111",
  42177=>"110111000",
  42178=>"100010001",
  42179=>"000011111",
  42180=>"110000000",
  42181=>"000001101",
  42182=>"110101100",
  42183=>"100010101",
  42184=>"011010110",
  42185=>"001001101",
  42186=>"100111111",
  42187=>"111010011",
  42188=>"011100000",
  42189=>"101111100",
  42190=>"000110011",
  42191=>"111100010",
  42192=>"101100011",
  42193=>"011101011",
  42194=>"000011000",
  42195=>"111000000",
  42196=>"010101011",
  42197=>"010101101",
  42198=>"101111110",
  42199=>"001001011",
  42200=>"001001111",
  42201=>"010110110",
  42202=>"000100010",
  42203=>"100100101",
  42204=>"101011010",
  42205=>"101110110",
  42206=>"001000100",
  42207=>"010010001",
  42208=>"000010000",
  42209=>"100100101",
  42210=>"101011001",
  42211=>"011010100",
  42212=>"011110011",
  42213=>"110110011",
  42214=>"100010000",
  42215=>"000001001",
  42216=>"000001000",
  42217=>"101100110",
  42218=>"000000011",
  42219=>"011111110",
  42220=>"101111000",
  42221=>"100100010",
  42222=>"010010100",
  42223=>"100010110",
  42224=>"001111110",
  42225=>"110001001",
  42226=>"000011111",
  42227=>"000111000",
  42228=>"011011111",
  42229=>"111010101",
  42230=>"001000011",
  42231=>"110001010",
  42232=>"001011100",
  42233=>"110100101",
  42234=>"111001110",
  42235=>"111000001",
  42236=>"100001010",
  42237=>"111100000",
  42238=>"100011110",
  42239=>"110101111",
  42240=>"101110000",
  42241=>"001000011",
  42242=>"001100001",
  42243=>"000011111",
  42244=>"001110111",
  42245=>"101011100",
  42246=>"001011111",
  42247=>"111111100",
  42248=>"000011100",
  42249=>"101101000",
  42250=>"000110011",
  42251=>"001001110",
  42252=>"001111000",
  42253=>"001100001",
  42254=>"010010110",
  42255=>"011000010",
  42256=>"011001010",
  42257=>"000101000",
  42258=>"000001000",
  42259=>"001111001",
  42260=>"011001100",
  42261=>"001011110",
  42262=>"101111100",
  42263=>"011100111",
  42264=>"001001010",
  42265=>"010100010",
  42266=>"100010111",
  42267=>"100110101",
  42268=>"001011101",
  42269=>"111100111",
  42270=>"100011100",
  42271=>"000001110",
  42272=>"001001000",
  42273=>"011010001",
  42274=>"010001100",
  42275=>"111000111",
  42276=>"110011111",
  42277=>"001111001",
  42278=>"101011100",
  42279=>"001001011",
  42280=>"001100001",
  42281=>"000001101",
  42282=>"111110110",
  42283=>"001000110",
  42284=>"101000110",
  42285=>"001110110",
  42286=>"000010011",
  42287=>"000101001",
  42288=>"001111111",
  42289=>"010001110",
  42290=>"100011101",
  42291=>"000010001",
  42292=>"011110001",
  42293=>"110001110",
  42294=>"000101110",
  42295=>"000100111",
  42296=>"000001010",
  42297=>"000101100",
  42298=>"011111110",
  42299=>"101110110",
  42300=>"100010001",
  42301=>"001011000",
  42302=>"010110010",
  42303=>"011100101",
  42304=>"010111110",
  42305=>"101000010",
  42306=>"111110100",
  42307=>"001010101",
  42308=>"100001011",
  42309=>"101100100",
  42310=>"011000000",
  42311=>"111010100",
  42312=>"101011111",
  42313=>"001100011",
  42314=>"100111010",
  42315=>"000010100",
  42316=>"101010000",
  42317=>"010000101",
  42318=>"111110010",
  42319=>"010001000",
  42320=>"011101111",
  42321=>"000010111",
  42322=>"111000001",
  42323=>"011110000",
  42324=>"101101101",
  42325=>"100000000",
  42326=>"111010110",
  42327=>"100000111",
  42328=>"100100000",
  42329=>"000000010",
  42330=>"111110100",
  42331=>"000111000",
  42332=>"011111000",
  42333=>"101011110",
  42334=>"000010010",
  42335=>"011100011",
  42336=>"100101101",
  42337=>"100001110",
  42338=>"101100001",
  42339=>"000001100",
  42340=>"001001000",
  42341=>"101000011",
  42342=>"101011111",
  42343=>"100110011",
  42344=>"001000001",
  42345=>"110101100",
  42346=>"001010010",
  42347=>"000010110",
  42348=>"001101001",
  42349=>"000010010",
  42350=>"001000110",
  42351=>"010100111",
  42352=>"000101000",
  42353=>"011101101",
  42354=>"100000010",
  42355=>"011110110",
  42356=>"011001001",
  42357=>"010100100",
  42358=>"110101110",
  42359=>"100011000",
  42360=>"100101010",
  42361=>"011010110",
  42362=>"100101010",
  42363=>"101001001",
  42364=>"001001100",
  42365=>"010001100",
  42366=>"001100000",
  42367=>"011111101",
  42368=>"001100110",
  42369=>"011000001",
  42370=>"111011111",
  42371=>"001011110",
  42372=>"010010100",
  42373=>"110001001",
  42374=>"100010010",
  42375=>"101001101",
  42376=>"111110001",
  42377=>"000101100",
  42378=>"000001100",
  42379=>"111001000",
  42380=>"100111001",
  42381=>"100011110",
  42382=>"110000011",
  42383=>"011010111",
  42384=>"111010111",
  42385=>"111100111",
  42386=>"011000110",
  42387=>"100100011",
  42388=>"101100100",
  42389=>"000001111",
  42390=>"000000100",
  42391=>"011110101",
  42392=>"011101000",
  42393=>"001011011",
  42394=>"010111011",
  42395=>"100001100",
  42396=>"101100011",
  42397=>"011001010",
  42398=>"100100101",
  42399=>"100011101",
  42400=>"010100110",
  42401=>"010111101",
  42402=>"010110011",
  42403=>"010101000",
  42404=>"110011110",
  42405=>"011010010",
  42406=>"001010110",
  42407=>"001110100",
  42408=>"011100001",
  42409=>"100010001",
  42410=>"111111000",
  42411=>"111100101",
  42412=>"100100010",
  42413=>"111010000",
  42414=>"110010101",
  42415=>"011011000",
  42416=>"110101001",
  42417=>"111101111",
  42418=>"010100101",
  42419=>"010000010",
  42420=>"101010001",
  42421=>"101010100",
  42422=>"100101010",
  42423=>"000010010",
  42424=>"111101010",
  42425=>"001101010",
  42426=>"111001011",
  42427=>"000001110",
  42428=>"111011010",
  42429=>"011001110",
  42430=>"101010000",
  42431=>"010011010",
  42432=>"001000001",
  42433=>"000000000",
  42434=>"010100011",
  42435=>"111101011",
  42436=>"110000110",
  42437=>"011101001",
  42438=>"101000011",
  42439=>"111111100",
  42440=>"000001000",
  42441=>"100111001",
  42442=>"111000100",
  42443=>"101101110",
  42444=>"000111011",
  42445=>"110101000",
  42446=>"100011110",
  42447=>"111100111",
  42448=>"101101110",
  42449=>"000010000",
  42450=>"111100110",
  42451=>"110110100",
  42452=>"000010100",
  42453=>"100000111",
  42454=>"111000000",
  42455=>"101001000",
  42456=>"101001001",
  42457=>"111110010",
  42458=>"101011101",
  42459=>"100000110",
  42460=>"100100010",
  42461=>"110110000",
  42462=>"011110111",
  42463=>"010000110",
  42464=>"001111111",
  42465=>"001101000",
  42466=>"111110001",
  42467=>"000100110",
  42468=>"000010001",
  42469=>"111111111",
  42470=>"010100011",
  42471=>"100111100",
  42472=>"001000000",
  42473=>"110100100",
  42474=>"100000101",
  42475=>"011001000",
  42476=>"100100110",
  42477=>"110110011",
  42478=>"110101000",
  42479=>"000111100",
  42480=>"100011111",
  42481=>"010100100",
  42482=>"111100110",
  42483=>"000000000",
  42484=>"010110110",
  42485=>"000000011",
  42486=>"010001111",
  42487=>"011101011",
  42488=>"010111001",
  42489=>"100011000",
  42490=>"111001001",
  42491=>"000101101",
  42492=>"100011000",
  42493=>"001001010",
  42494=>"100001110",
  42495=>"010111000",
  42496=>"000111000",
  42497=>"101100000",
  42498=>"110100011",
  42499=>"101110001",
  42500=>"000000001",
  42501=>"011001000",
  42502=>"101010110",
  42503=>"101101100",
  42504=>"011110110",
  42505=>"101100100",
  42506=>"101101010",
  42507=>"010001010",
  42508=>"010101101",
  42509=>"100010110",
  42510=>"111011001",
  42511=>"101011010",
  42512=>"000100100",
  42513=>"001001101",
  42514=>"011001011",
  42515=>"110100010",
  42516=>"110010101",
  42517=>"011101010",
  42518=>"101111010",
  42519=>"000110000",
  42520=>"010001000",
  42521=>"110110110",
  42522=>"010000010",
  42523=>"100010111",
  42524=>"110111001",
  42525=>"000000011",
  42526=>"101001010",
  42527=>"110100101",
  42528=>"000100010",
  42529=>"100010011",
  42530=>"001000011",
  42531=>"111010000",
  42532=>"110000011",
  42533=>"101011011",
  42534=>"101011011",
  42535=>"101111111",
  42536=>"101111001",
  42537=>"011001110",
  42538=>"101010101",
  42539=>"111110000",
  42540=>"010100001",
  42541=>"001001000",
  42542=>"000000011",
  42543=>"001010011",
  42544=>"011010100",
  42545=>"101100011",
  42546=>"101010101",
  42547=>"011110110",
  42548=>"010101000",
  42549=>"100000000",
  42550=>"001100001",
  42551=>"111101000",
  42552=>"111000110",
  42553=>"011101010",
  42554=>"000111011",
  42555=>"011010011",
  42556=>"000110100",
  42557=>"110101111",
  42558=>"100000001",
  42559=>"111111010",
  42560=>"111000101",
  42561=>"101010001",
  42562=>"001011000",
  42563=>"100101000",
  42564=>"101111111",
  42565=>"101010000",
  42566=>"010001001",
  42567=>"010100001",
  42568=>"001110101",
  42569=>"110111001",
  42570=>"011010011",
  42571=>"100100100",
  42572=>"101010110",
  42573=>"010010010",
  42574=>"101101110",
  42575=>"101011100",
  42576=>"001001010",
  42577=>"111101011",
  42578=>"001001001",
  42579=>"110000001",
  42580=>"100000111",
  42581=>"000100010",
  42582=>"101101101",
  42583=>"001101001",
  42584=>"101011101",
  42585=>"011110000",
  42586=>"001100100",
  42587=>"011010000",
  42588=>"111010001",
  42589=>"010100101",
  42590=>"010101111",
  42591=>"111111100",
  42592=>"110010110",
  42593=>"010110100",
  42594=>"100010111",
  42595=>"000101011",
  42596=>"011010100",
  42597=>"111001111",
  42598=>"110111111",
  42599=>"011100001",
  42600=>"001001000",
  42601=>"100011001",
  42602=>"001111101",
  42603=>"110010001",
  42604=>"001100110",
  42605=>"001001100",
  42606=>"011000011",
  42607=>"100011000",
  42608=>"011001110",
  42609=>"000111010",
  42610=>"101110111",
  42611=>"111111000",
  42612=>"010001101",
  42613=>"111101000",
  42614=>"110010010",
  42615=>"000110101",
  42616=>"111011111",
  42617=>"101111000",
  42618=>"110111100",
  42619=>"110100001",
  42620=>"001011011",
  42621=>"111000011",
  42622=>"111101011",
  42623=>"000000100",
  42624=>"100000110",
  42625=>"110110011",
  42626=>"010111000",
  42627=>"001000010",
  42628=>"001001000",
  42629=>"100100000",
  42630=>"100000101",
  42631=>"101011010",
  42632=>"100100011",
  42633=>"001010000",
  42634=>"111101011",
  42635=>"011010101",
  42636=>"010110110",
  42637=>"001000111",
  42638=>"101000011",
  42639=>"110111010",
  42640=>"110010101",
  42641=>"000111110",
  42642=>"001001001",
  42643=>"110100110",
  42644=>"000100011",
  42645=>"101111110",
  42646=>"010000001",
  42647=>"101111100",
  42648=>"010111100",
  42649=>"001010101",
  42650=>"001100010",
  42651=>"000010111",
  42652=>"111010100",
  42653=>"000001001",
  42654=>"001100000",
  42655=>"011111110",
  42656=>"011101100",
  42657=>"111111011",
  42658=>"101101100",
  42659=>"000000111",
  42660=>"111101010",
  42661=>"101111000",
  42662=>"011111101",
  42663=>"011001100",
  42664=>"111111001",
  42665=>"011101000",
  42666=>"111011100",
  42667=>"101110000",
  42668=>"000010100",
  42669=>"110001011",
  42670=>"110100111",
  42671=>"011000100",
  42672=>"000010110",
  42673=>"110010011",
  42674=>"000001011",
  42675=>"001110001",
  42676=>"011100000",
  42677=>"001010001",
  42678=>"000101100",
  42679=>"101110010",
  42680=>"110100100",
  42681=>"110111110",
  42682=>"100011000",
  42683=>"000001000",
  42684=>"010000001",
  42685=>"001000001",
  42686=>"010010101",
  42687=>"001111010",
  42688=>"011010110",
  42689=>"001010000",
  42690=>"111110111",
  42691=>"011100001",
  42692=>"001100100",
  42693=>"100100101",
  42694=>"111011001",
  42695=>"011110110",
  42696=>"110101000",
  42697=>"110010001",
  42698=>"100000000",
  42699=>"010011010",
  42700=>"010010111",
  42701=>"010110110",
  42702=>"001010001",
  42703=>"010010011",
  42704=>"001001001",
  42705=>"101000111",
  42706=>"010001000",
  42707=>"111000011",
  42708=>"001111100",
  42709=>"010100001",
  42710=>"111111110",
  42711=>"001100101",
  42712=>"001101101",
  42713=>"000110110",
  42714=>"010010011",
  42715=>"011001000",
  42716=>"110110000",
  42717=>"100111001",
  42718=>"110011001",
  42719=>"100101010",
  42720=>"011000101",
  42721=>"001010011",
  42722=>"011011011",
  42723=>"111001011",
  42724=>"000110010",
  42725=>"101001000",
  42726=>"000000010",
  42727=>"110100100",
  42728=>"011000000",
  42729=>"111001100",
  42730=>"101000011",
  42731=>"111111111",
  42732=>"110110000",
  42733=>"010011111",
  42734=>"011010000",
  42735=>"100000101",
  42736=>"100011110",
  42737=>"010000101",
  42738=>"101000010",
  42739=>"011011011",
  42740=>"100000100",
  42741=>"001100100",
  42742=>"000111111",
  42743=>"000110011",
  42744=>"000000000",
  42745=>"010101111",
  42746=>"100100000",
  42747=>"011010101",
  42748=>"100010111",
  42749=>"100010111",
  42750=>"110001000",
  42751=>"010100010",
  42752=>"101011011",
  42753=>"000100010",
  42754=>"110000101",
  42755=>"001010101",
  42756=>"101101000",
  42757=>"011000101",
  42758=>"001010000",
  42759=>"010011101",
  42760=>"000011000",
  42761=>"110110010",
  42762=>"100011110",
  42763=>"011110000",
  42764=>"011111100",
  42765=>"010010011",
  42766=>"000001010",
  42767=>"111110101",
  42768=>"011111110",
  42769=>"100101000",
  42770=>"111001100",
  42771=>"110101010",
  42772=>"000000110",
  42773=>"001111110",
  42774=>"011111101",
  42775=>"010110101",
  42776=>"011001011",
  42777=>"011010001",
  42778=>"101110000",
  42779=>"100000011",
  42780=>"011111010",
  42781=>"001011010",
  42782=>"111000100",
  42783=>"000111001",
  42784=>"111011001",
  42785=>"100010000",
  42786=>"011110011",
  42787=>"101100010",
  42788=>"010111010",
  42789=>"001100000",
  42790=>"000011101",
  42791=>"011110101",
  42792=>"001001100",
  42793=>"111101000",
  42794=>"011100111",
  42795=>"110101100",
  42796=>"010010110",
  42797=>"000000100",
  42798=>"010001100",
  42799=>"110100110",
  42800=>"011000100",
  42801=>"000010111",
  42802=>"100111011",
  42803=>"000110100",
  42804=>"101000111",
  42805=>"101010110",
  42806=>"110010101",
  42807=>"010010010",
  42808=>"101110000",
  42809=>"111111100",
  42810=>"011101010",
  42811=>"001110100",
  42812=>"101001100",
  42813=>"110100000",
  42814=>"101111101",
  42815=>"011011111",
  42816=>"010000101",
  42817=>"110100100",
  42818=>"101000100",
  42819=>"111111110",
  42820=>"111100100",
  42821=>"011111010",
  42822=>"111000011",
  42823=>"101101110",
  42824=>"010000101",
  42825=>"001100001",
  42826=>"000000001",
  42827=>"110011110",
  42828=>"110101100",
  42829=>"111000111",
  42830=>"111100010",
  42831=>"101010010",
  42832=>"101001000",
  42833=>"100010011",
  42834=>"010100000",
  42835=>"111100010",
  42836=>"101011001",
  42837=>"000011001",
  42838=>"000010111",
  42839=>"111011110",
  42840=>"101010010",
  42841=>"101110001",
  42842=>"100111010",
  42843=>"111001001",
  42844=>"110110011",
  42845=>"010001101",
  42846=>"101011000",
  42847=>"101000111",
  42848=>"000001010",
  42849=>"111001100",
  42850=>"000100111",
  42851=>"110111010",
  42852=>"001110101",
  42853=>"111000000",
  42854=>"010111001",
  42855=>"110011001",
  42856=>"111011011",
  42857=>"010101101",
  42858=>"111010110",
  42859=>"011101001",
  42860=>"011010111",
  42861=>"000111100",
  42862=>"010001110",
  42863=>"101010110",
  42864=>"010101011",
  42865=>"111011001",
  42866=>"101101000",
  42867=>"110100000",
  42868=>"010100000",
  42869=>"010101001",
  42870=>"010100010",
  42871=>"000100010",
  42872=>"001001100",
  42873=>"110001001",
  42874=>"101111100",
  42875=>"010110000",
  42876=>"010000000",
  42877=>"111101111",
  42878=>"111101110",
  42879=>"111110110",
  42880=>"001011110",
  42881=>"110010000",
  42882=>"011100011",
  42883=>"010100110",
  42884=>"111111011",
  42885=>"010000110",
  42886=>"000000100",
  42887=>"110101000",
  42888=>"100100010",
  42889=>"000111011",
  42890=>"101111101",
  42891=>"110000111",
  42892=>"110111000",
  42893=>"011001110",
  42894=>"010010000",
  42895=>"111110111",
  42896=>"010101001",
  42897=>"111011100",
  42898=>"111000000",
  42899=>"111011110",
  42900=>"111011001",
  42901=>"111011101",
  42902=>"101110111",
  42903=>"011101010",
  42904=>"010100100",
  42905=>"001000100",
  42906=>"110101000",
  42907=>"111010111",
  42908=>"010000101",
  42909=>"101110010",
  42910=>"010011001",
  42911=>"000000000",
  42912=>"111111000",
  42913=>"011111111",
  42914=>"000010100",
  42915=>"110110110",
  42916=>"110001111",
  42917=>"100001001",
  42918=>"100110110",
  42919=>"001000000",
  42920=>"100011101",
  42921=>"011010000",
  42922=>"001010000",
  42923=>"010001111",
  42924=>"001010110",
  42925=>"000001111",
  42926=>"111010000",
  42927=>"110001110",
  42928=>"000000001",
  42929=>"100001001",
  42930=>"001000011",
  42931=>"010001111",
  42932=>"010010001",
  42933=>"001111111",
  42934=>"010111101",
  42935=>"001010011",
  42936=>"110000001",
  42937=>"111100010",
  42938=>"111110011",
  42939=>"100010100",
  42940=>"111111011",
  42941=>"000100001",
  42942=>"111000011",
  42943=>"100101110",
  42944=>"011100001",
  42945=>"000000001",
  42946=>"000011110",
  42947=>"110110000",
  42948=>"100100110",
  42949=>"011100011",
  42950=>"011101110",
  42951=>"110001110",
  42952=>"100010101",
  42953=>"100100110",
  42954=>"111101101",
  42955=>"101110100",
  42956=>"111111010",
  42957=>"000001110",
  42958=>"100100100",
  42959=>"011011001",
  42960=>"010011110",
  42961=>"111110011",
  42962=>"001010100",
  42963=>"011010000",
  42964=>"111000010",
  42965=>"010101001",
  42966=>"100001100",
  42967=>"110010100",
  42968=>"000101110",
  42969=>"000011010",
  42970=>"111011111",
  42971=>"101011000",
  42972=>"100110000",
  42973=>"110011110",
  42974=>"111010111",
  42975=>"100110100",
  42976=>"000101100",
  42977=>"101010111",
  42978=>"100000111",
  42979=>"111100010",
  42980=>"110100110",
  42981=>"111000010",
  42982=>"100100000",
  42983=>"100101110",
  42984=>"011000010",
  42985=>"000110101",
  42986=>"011011001",
  42987=>"101110101",
  42988=>"100010000",
  42989=>"111010110",
  42990=>"011000000",
  42991=>"110011101",
  42992=>"011000011",
  42993=>"011001001",
  42994=>"001011011",
  42995=>"010111100",
  42996=>"000001110",
  42997=>"010011001",
  42998=>"011011010",
  42999=>"100010011",
  43000=>"010001001",
  43001=>"011011111",
  43002=>"010001010",
  43003=>"100101100",
  43004=>"101110110",
  43005=>"011100010",
  43006=>"000010001",
  43007=>"000101100",
  43008=>"011101101",
  43009=>"001101011",
  43010=>"100111100",
  43011=>"101100111",
  43012=>"100111000",
  43013=>"011000111",
  43014=>"010110000",
  43015=>"001110011",
  43016=>"101110100",
  43017=>"011100101",
  43018=>"010000010",
  43019=>"010010110",
  43020=>"010010010",
  43021=>"111111111",
  43022=>"011100100",
  43023=>"010111110",
  43024=>"001000001",
  43025=>"001000111",
  43026=>"011010000",
  43027=>"001001000",
  43028=>"111111001",
  43029=>"101101010",
  43030=>"100100010",
  43031=>"000001011",
  43032=>"100100011",
  43033=>"010000111",
  43034=>"010000111",
  43035=>"111101111",
  43036=>"101011000",
  43037=>"101001011",
  43038=>"011111001",
  43039=>"000001110",
  43040=>"001100101",
  43041=>"000010011",
  43042=>"110010010",
  43043=>"111010100",
  43044=>"011000111",
  43045=>"100100100",
  43046=>"011000101",
  43047=>"001001111",
  43048=>"110110110",
  43049=>"011010011",
  43050=>"110110101",
  43051=>"111011110",
  43052=>"011010110",
  43053=>"110111101",
  43054=>"101111001",
  43055=>"100001110",
  43056=>"100000111",
  43057=>"000001111",
  43058=>"001111010",
  43059=>"111011101",
  43060=>"110110101",
  43061=>"010010000",
  43062=>"110011110",
  43063=>"000100010",
  43064=>"000001101",
  43065=>"001101101",
  43066=>"000110010",
  43067=>"110010000",
  43068=>"100000001",
  43069=>"101101001",
  43070=>"111010010",
  43071=>"100101100",
  43072=>"000100101",
  43073=>"000000000",
  43074=>"001001111",
  43075=>"110110101",
  43076=>"101111111",
  43077=>"011011000",
  43078=>"100111000",
  43079=>"000100010",
  43080=>"110110010",
  43081=>"010011110",
  43082=>"111001000",
  43083=>"110111011",
  43084=>"010000111",
  43085=>"011101110",
  43086=>"000111111",
  43087=>"110000100",
  43088=>"100101111",
  43089=>"011011011",
  43090=>"010100000",
  43091=>"011011110",
  43092=>"100100011",
  43093=>"011000000",
  43094=>"101011100",
  43095=>"101001000",
  43096=>"111011111",
  43097=>"011001101",
  43098=>"001111001",
  43099=>"010110011",
  43100=>"011010101",
  43101=>"000100000",
  43102=>"011100011",
  43103=>"001101101",
  43104=>"111110101",
  43105=>"001111001",
  43106=>"001010101",
  43107=>"111010010",
  43108=>"100010000",
  43109=>"110111001",
  43110=>"100010000",
  43111=>"111100011",
  43112=>"110101001",
  43113=>"110000110",
  43114=>"000100011",
  43115=>"010010101",
  43116=>"011001011",
  43117=>"011110010",
  43118=>"110100011",
  43119=>"000000111",
  43120=>"111100101",
  43121=>"000100111",
  43122=>"111100000",
  43123=>"001010111",
  43124=>"101110100",
  43125=>"000101011",
  43126=>"101101011",
  43127=>"111110001",
  43128=>"110010000",
  43129=>"010101101",
  43130=>"111111101",
  43131=>"110010110",
  43132=>"001101000",
  43133=>"001100011",
  43134=>"010101111",
  43135=>"001101000",
  43136=>"111110000",
  43137=>"101000111",
  43138=>"111111000",
  43139=>"011000010",
  43140=>"101011000",
  43141=>"011001100",
  43142=>"110000110",
  43143=>"000011000",
  43144=>"001110001",
  43145=>"101111001",
  43146=>"010110110",
  43147=>"010001111",
  43148=>"101000100",
  43149=>"010101010",
  43150=>"101110111",
  43151=>"001111110",
  43152=>"101110000",
  43153=>"110000111",
  43154=>"101010011",
  43155=>"100001000",
  43156=>"100001001",
  43157=>"100101101",
  43158=>"010010010",
  43159=>"001000010",
  43160=>"001010000",
  43161=>"001010110",
  43162=>"110011000",
  43163=>"011101000",
  43164=>"110100010",
  43165=>"111111010",
  43166=>"011000110",
  43167=>"101000011",
  43168=>"101010001",
  43169=>"101111011",
  43170=>"110001111",
  43171=>"001001101",
  43172=>"011000111",
  43173=>"001100111",
  43174=>"000011111",
  43175=>"111000011",
  43176=>"100001010",
  43177=>"010001111",
  43178=>"011001011",
  43179=>"100010101",
  43180=>"100000000",
  43181=>"010011110",
  43182=>"001011001",
  43183=>"011111010",
  43184=>"001011100",
  43185=>"000000000",
  43186=>"110110011",
  43187=>"000011101",
  43188=>"111000111",
  43189=>"101000001",
  43190=>"001000011",
  43191=>"000000010",
  43192=>"000000001",
  43193=>"001000111",
  43194=>"001011010",
  43195=>"111011000",
  43196=>"110001011",
  43197=>"010011001",
  43198=>"100110101",
  43199=>"000000000",
  43200=>"010101001",
  43201=>"011100100",
  43202=>"110000011",
  43203=>"010111111",
  43204=>"100000001",
  43205=>"000101110",
  43206=>"001011010",
  43207=>"111000100",
  43208=>"110111111",
  43209=>"011111011",
  43210=>"111010000",
  43211=>"001110000",
  43212=>"111001110",
  43213=>"000000111",
  43214=>"011111000",
  43215=>"100000000",
  43216=>"011100000",
  43217=>"001100011",
  43218=>"000001111",
  43219=>"110100100",
  43220=>"100001001",
  43221=>"011010100",
  43222=>"010110011",
  43223=>"010111110",
  43224=>"100100000",
  43225=>"011100000",
  43226=>"101100100",
  43227=>"111101011",
  43228=>"100010100",
  43229=>"001011111",
  43230=>"101010011",
  43231=>"001110001",
  43232=>"000000100",
  43233=>"001100010",
  43234=>"110010000",
  43235=>"010111001",
  43236=>"101010100",
  43237=>"001000000",
  43238=>"001000100",
  43239=>"101111111",
  43240=>"011100000",
  43241=>"101110101",
  43242=>"111101111",
  43243=>"111010011",
  43244=>"100110110",
  43245=>"101100001",
  43246=>"011111011",
  43247=>"000001000",
  43248=>"110111001",
  43249=>"111111011",
  43250=>"100110011",
  43251=>"001000100",
  43252=>"100110101",
  43253=>"000100100",
  43254=>"010110111",
  43255=>"010000101",
  43256=>"111100111",
  43257=>"011010000",
  43258=>"101000111",
  43259=>"101000001",
  43260=>"000100000",
  43261=>"010001011",
  43262=>"010111111",
  43263=>"010101101",
  43264=>"111111000",
  43265=>"101110111",
  43266=>"001001101",
  43267=>"000000110",
  43268=>"000001011",
  43269=>"001010110",
  43270=>"011111100",
  43271=>"111000000",
  43272=>"010101110",
  43273=>"110001101",
  43274=>"111111111",
  43275=>"100100000",
  43276=>"111000110",
  43277=>"000101110",
  43278=>"010000001",
  43279=>"111001001",
  43280=>"011110110",
  43281=>"100011011",
  43282=>"110111101",
  43283=>"011010100",
  43284=>"101101010",
  43285=>"100101111",
  43286=>"010110011",
  43287=>"100101101",
  43288=>"000101110",
  43289=>"001111010",
  43290=>"011010001",
  43291=>"001000000",
  43292=>"001000001",
  43293=>"100010001",
  43294=>"011011111",
  43295=>"000001000",
  43296=>"010010100",
  43297=>"100111011",
  43298=>"111111010",
  43299=>"111001101",
  43300=>"111110011",
  43301=>"011110101",
  43302=>"101001010",
  43303=>"101001011",
  43304=>"001001001",
  43305=>"111110101",
  43306=>"100010110",
  43307=>"000100000",
  43308=>"000100111",
  43309=>"011110101",
  43310=>"000000010",
  43311=>"111010110",
  43312=>"111010000",
  43313=>"010010011",
  43314=>"111110100",
  43315=>"100101111",
  43316=>"000100111",
  43317=>"001101110",
  43318=>"000010011",
  43319=>"001111000",
  43320=>"110010110",
  43321=>"101101001",
  43322=>"110011110",
  43323=>"111100101",
  43324=>"000010111",
  43325=>"000011001",
  43326=>"001110010",
  43327=>"010010000",
  43328=>"110000000",
  43329=>"100000010",
  43330=>"000011110",
  43331=>"110000001",
  43332=>"101111110",
  43333=>"010110101",
  43334=>"000101000",
  43335=>"011101111",
  43336=>"000110101",
  43337=>"001110100",
  43338=>"001010111",
  43339=>"110101010",
  43340=>"011011010",
  43341=>"000011011",
  43342=>"110011111",
  43343=>"101111111",
  43344=>"010001000",
  43345=>"111000110",
  43346=>"001011010",
  43347=>"101011100",
  43348=>"000101111",
  43349=>"000011001",
  43350=>"100011000",
  43351=>"111110000",
  43352=>"100100000",
  43353=>"010010110",
  43354=>"001110010",
  43355=>"010000100",
  43356=>"110101111",
  43357=>"010101100",
  43358=>"101111010",
  43359=>"001111001",
  43360=>"110010111",
  43361=>"011010011",
  43362=>"110001001",
  43363=>"001011001",
  43364=>"010010100",
  43365=>"101100001",
  43366=>"111010010",
  43367=>"000110011",
  43368=>"000100010",
  43369=>"101110100",
  43370=>"000110100",
  43371=>"101100110",
  43372=>"000000010",
  43373=>"110111100",
  43374=>"001000011",
  43375=>"011011001",
  43376=>"011001111",
  43377=>"000110011",
  43378=>"110010010",
  43379=>"100011000",
  43380=>"111011110",
  43381=>"011111000",
  43382=>"010001110",
  43383=>"110111001",
  43384=>"110000010",
  43385=>"111000111",
  43386=>"101111100",
  43387=>"000000111",
  43388=>"110110010",
  43389=>"000110010",
  43390=>"100101001",
  43391=>"111110111",
  43392=>"110000000",
  43393=>"001000110",
  43394=>"101111001",
  43395=>"010011000",
  43396=>"010001011",
  43397=>"010100010",
  43398=>"011101001",
  43399=>"011010010",
  43400=>"010001100",
  43401=>"011111011",
  43402=>"000101011",
  43403=>"101001011",
  43404=>"010010110",
  43405=>"101101110",
  43406=>"011000111",
  43407=>"001001110",
  43408=>"100100111",
  43409=>"100001001",
  43410=>"001010001",
  43411=>"110011011",
  43412=>"101100000",
  43413=>"000001000",
  43414=>"111111110",
  43415=>"111101011",
  43416=>"000100000",
  43417=>"011100010",
  43418=>"010011100",
  43419=>"111101110",
  43420=>"100011010",
  43421=>"010011001",
  43422=>"011011001",
  43423=>"101000111",
  43424=>"011011000",
  43425=>"111101001",
  43426=>"010011111",
  43427=>"100000000",
  43428=>"111100001",
  43429=>"010000100",
  43430=>"000001111",
  43431=>"010111111",
  43432=>"011111011",
  43433=>"101010010",
  43434=>"000100010",
  43435=>"100001001",
  43436=>"010101000",
  43437=>"000100010",
  43438=>"000110010",
  43439=>"000100010",
  43440=>"101110100",
  43441=>"110000001",
  43442=>"000101101",
  43443=>"111000011",
  43444=>"110111000",
  43445=>"100011110",
  43446=>"001100000",
  43447=>"010100101",
  43448=>"000010101",
  43449=>"101101011",
  43450=>"111101111",
  43451=>"111110100",
  43452=>"100110001",
  43453=>"111111101",
  43454=>"010011100",
  43455=>"000010111",
  43456=>"110111001",
  43457=>"111001001",
  43458=>"101101011",
  43459=>"010010110",
  43460=>"010010000",
  43461=>"101001000",
  43462=>"001011101",
  43463=>"010110111",
  43464=>"010011000",
  43465=>"001111010",
  43466=>"011100001",
  43467=>"010011101",
  43468=>"111110001",
  43469=>"001110000",
  43470=>"101110110",
  43471=>"100011011",
  43472=>"001110101",
  43473=>"001100101",
  43474=>"011001111",
  43475=>"111111111",
  43476=>"110000100",
  43477=>"000100000",
  43478=>"011100100",
  43479=>"110110111",
  43480=>"110110000",
  43481=>"011110111",
  43482=>"000010111",
  43483=>"011111011",
  43484=>"001011100",
  43485=>"000111110",
  43486=>"110101000",
  43487=>"001101000",
  43488=>"001100001",
  43489=>"101101111",
  43490=>"010000000",
  43491=>"010101101",
  43492=>"100110011",
  43493=>"110110100",
  43494=>"001110100",
  43495=>"011001011",
  43496=>"111000001",
  43497=>"011010111",
  43498=>"000110010",
  43499=>"101011000",
  43500=>"010100100",
  43501=>"101000110",
  43502=>"111010100",
  43503=>"000111110",
  43504=>"001010010",
  43505=>"110110010",
  43506=>"000010101",
  43507=>"110001000",
  43508=>"010101110",
  43509=>"010011010",
  43510=>"010000110",
  43511=>"001110110",
  43512=>"001001010",
  43513=>"111011011",
  43514=>"011000110",
  43515=>"011000011",
  43516=>"010110010",
  43517=>"000010010",
  43518=>"000010100",
  43519=>"110100101",
  43520=>"101001110",
  43521=>"100001011",
  43522=>"001101111",
  43523=>"101101000",
  43524=>"010000110",
  43525=>"101110111",
  43526=>"011100000",
  43527=>"111011000",
  43528=>"101100110",
  43529=>"001010010",
  43530=>"101000100",
  43531=>"000111011",
  43532=>"001100011",
  43533=>"100001101",
  43534=>"011000111",
  43535=>"001010011",
  43536=>"000011111",
  43537=>"011011010",
  43538=>"001010011",
  43539=>"011101101",
  43540=>"011001001",
  43541=>"100001110",
  43542=>"100101000",
  43543=>"010100001",
  43544=>"001100001",
  43545=>"101001010",
  43546=>"000000110",
  43547=>"111001000",
  43548=>"010100111",
  43549=>"000001111",
  43550=>"011001000",
  43551=>"010011000",
  43552=>"101011110",
  43553=>"011110000",
  43554=>"000000011",
  43555=>"100001100",
  43556=>"101110000",
  43557=>"010101111",
  43558=>"000010011",
  43559=>"010110010",
  43560=>"001010100",
  43561=>"110000000",
  43562=>"100001011",
  43563=>"011001100",
  43564=>"101011100",
  43565=>"000000110",
  43566=>"100010000",
  43567=>"101100001",
  43568=>"101100111",
  43569=>"110001110",
  43570=>"001000010",
  43571=>"011001000",
  43572=>"100001111",
  43573=>"000110111",
  43574=>"100010110",
  43575=>"100011101",
  43576=>"000011110",
  43577=>"000100001",
  43578=>"101110001",
  43579=>"100010111",
  43580=>"101101100",
  43581=>"010110110",
  43582=>"100000110",
  43583=>"011101000",
  43584=>"011111110",
  43585=>"101000011",
  43586=>"011110011",
  43587=>"001011001",
  43588=>"101000000",
  43589=>"100111101",
  43590=>"011010101",
  43591=>"100000110",
  43592=>"001011111",
  43593=>"000111011",
  43594=>"000001010",
  43595=>"110110000",
  43596=>"101010001",
  43597=>"010011100",
  43598=>"011100100",
  43599=>"101001000",
  43600=>"000110010",
  43601=>"100110100",
  43602=>"010011111",
  43603=>"001100000",
  43604=>"000100001",
  43605=>"011011101",
  43606=>"001110111",
  43607=>"011110100",
  43608=>"100101111",
  43609=>"110010100",
  43610=>"110010000",
  43611=>"111111111",
  43612=>"100110110",
  43613=>"011000010",
  43614=>"000010110",
  43615=>"111001011",
  43616=>"101100001",
  43617=>"111000011",
  43618=>"111000111",
  43619=>"100010111",
  43620=>"101111011",
  43621=>"100111110",
  43622=>"111000111",
  43623=>"000001011",
  43624=>"100000110",
  43625=>"000100111",
  43626=>"100110010",
  43627=>"110100010",
  43628=>"100001101",
  43629=>"111111111",
  43630=>"011110111",
  43631=>"111000110",
  43632=>"100000110",
  43633=>"111111111",
  43634=>"000101000",
  43635=>"010100000",
  43636=>"101110101",
  43637=>"110011111",
  43638=>"100011011",
  43639=>"010101100",
  43640=>"000110000",
  43641=>"110110110",
  43642=>"011001100",
  43643=>"011001111",
  43644=>"001001100",
  43645=>"001111001",
  43646=>"011011101",
  43647=>"111001001",
  43648=>"000001010",
  43649=>"100100010",
  43650=>"010110110",
  43651=>"001001100",
  43652=>"011010010",
  43653=>"000100100",
  43654=>"100011111",
  43655=>"110010101",
  43656=>"000100111",
  43657=>"011110111",
  43658=>"111011000",
  43659=>"000001100",
  43660=>"000100000",
  43661=>"101100001",
  43662=>"011000111",
  43663=>"101111111",
  43664=>"001110110",
  43665=>"111100110",
  43666=>"111100011",
  43667=>"011111110",
  43668=>"001001101",
  43669=>"110011010",
  43670=>"001001111",
  43671=>"111010010",
  43672=>"010110001",
  43673=>"000000000",
  43674=>"101000110",
  43675=>"010111011",
  43676=>"010101010",
  43677=>"111101111",
  43678=>"110111100",
  43679=>"100000100",
  43680=>"001111000",
  43681=>"101011110",
  43682=>"011111010",
  43683=>"011101111",
  43684=>"000110000",
  43685=>"010001001",
  43686=>"000100010",
  43687=>"000111000",
  43688=>"010100110",
  43689=>"111011010",
  43690=>"010001001",
  43691=>"000111011",
  43692=>"101110110",
  43693=>"010110100",
  43694=>"000011001",
  43695=>"000010010",
  43696=>"100001000",
  43697=>"011110011",
  43698=>"101010111",
  43699=>"001101001",
  43700=>"110000011",
  43701=>"010011100",
  43702=>"111111101",
  43703=>"110000110",
  43704=>"001111010",
  43705=>"100101001",
  43706=>"010111010",
  43707=>"010010011",
  43708=>"110101001",
  43709=>"100110011",
  43710=>"011001001",
  43711=>"010001000",
  43712=>"100001100",
  43713=>"101101011",
  43714=>"000101110",
  43715=>"111110000",
  43716=>"110011000",
  43717=>"101101100",
  43718=>"010110011",
  43719=>"111111001",
  43720=>"001010101",
  43721=>"111001000",
  43722=>"110100001",
  43723=>"010110001",
  43724=>"000000101",
  43725=>"000100111",
  43726=>"100100110",
  43727=>"100110000",
  43728=>"011100110",
  43729=>"001101100",
  43730=>"100101011",
  43731=>"111101111",
  43732=>"110110111",
  43733=>"111001001",
  43734=>"011101001",
  43735=>"000100100",
  43736=>"000001000",
  43737=>"110111110",
  43738=>"110001100",
  43739=>"100111011",
  43740=>"010101111",
  43741=>"110000000",
  43742=>"000111111",
  43743=>"010010001",
  43744=>"010010010",
  43745=>"101111010",
  43746=>"011101100",
  43747=>"010111000",
  43748=>"110101000",
  43749=>"101011101",
  43750=>"001101000",
  43751=>"110000110",
  43752=>"111111110",
  43753=>"011100011",
  43754=>"111011001",
  43755=>"101011000",
  43756=>"110001011",
  43757=>"011011110",
  43758=>"101000101",
  43759=>"010000100",
  43760=>"011011110",
  43761=>"010100110",
  43762=>"101110001",
  43763=>"000011000",
  43764=>"101010001",
  43765=>"111010011",
  43766=>"100011110",
  43767=>"111110111",
  43768=>"101111001",
  43769=>"010001111",
  43770=>"001101111",
  43771=>"001101010",
  43772=>"011100000",
  43773=>"010001100",
  43774=>"011001011",
  43775=>"101111011",
  43776=>"101010011",
  43777=>"001011011",
  43778=>"100101110",
  43779=>"000110100",
  43780=>"011110100",
  43781=>"000001100",
  43782=>"010110010",
  43783=>"110111010",
  43784=>"101010010",
  43785=>"000000010",
  43786=>"000011100",
  43787=>"010000000",
  43788=>"011111111",
  43789=>"001010101",
  43790=>"010101100",
  43791=>"010000010",
  43792=>"110101111",
  43793=>"100110110",
  43794=>"001111011",
  43795=>"001101011",
  43796=>"111111001",
  43797=>"110001011",
  43798=>"011101111",
  43799=>"011000100",
  43800=>"110010101",
  43801=>"100001001",
  43802=>"111111101",
  43803=>"000110001",
  43804=>"110000011",
  43805=>"011011111",
  43806=>"001101000",
  43807=>"011000011",
  43808=>"100110111",
  43809=>"000110011",
  43810=>"010001100",
  43811=>"100010011",
  43812=>"000010000",
  43813=>"010000000",
  43814=>"010101000",
  43815=>"111100000",
  43816=>"011100101",
  43817=>"101111001",
  43818=>"100010010",
  43819=>"011100110",
  43820=>"111000000",
  43821=>"111001000",
  43822=>"111010101",
  43823=>"101011100",
  43824=>"111101110",
  43825=>"010101101",
  43826=>"110110010",
  43827=>"010001101",
  43828=>"010111000",
  43829=>"100100111",
  43830=>"011010001",
  43831=>"100110011",
  43832=>"011011101",
  43833=>"100000001",
  43834=>"000000001",
  43835=>"101100000",
  43836=>"110101101",
  43837=>"111100101",
  43838=>"101100010",
  43839=>"101100011",
  43840=>"100100010",
  43841=>"110110100",
  43842=>"000001011",
  43843=>"100111000",
  43844=>"010001010",
  43845=>"001110010",
  43846=>"110010101",
  43847=>"100000011",
  43848=>"111010100",
  43849=>"100000010",
  43850=>"011011010",
  43851=>"111111110",
  43852=>"010010010",
  43853=>"100111010",
  43854=>"000001101",
  43855=>"000100001",
  43856=>"011101110",
  43857=>"100111000",
  43858=>"110000010",
  43859=>"000001011",
  43860=>"101000101",
  43861=>"011001111",
  43862=>"011100101",
  43863=>"101100111",
  43864=>"110101110",
  43865=>"110110010",
  43866=>"101100111",
  43867=>"011110000",
  43868=>"001111101",
  43869=>"100000100",
  43870=>"000000001",
  43871=>"000000001",
  43872=>"111110100",
  43873=>"000011000",
  43874=>"000100101",
  43875=>"111101010",
  43876=>"000010010",
  43877=>"010010001",
  43878=>"011110111",
  43879=>"011000010",
  43880=>"011100110",
  43881=>"101111110",
  43882=>"001111111",
  43883=>"100100010",
  43884=>"001101110",
  43885=>"000000000",
  43886=>"010010011",
  43887=>"110101100",
  43888=>"010011100",
  43889=>"010100100",
  43890=>"101001101",
  43891=>"101101111",
  43892=>"000001011",
  43893=>"111100111",
  43894=>"111101101",
  43895=>"111010001",
  43896=>"101010011",
  43897=>"101001100",
  43898=>"011001110",
  43899=>"001010000",
  43900=>"000000001",
  43901=>"111001110",
  43902=>"001011111",
  43903=>"110101111",
  43904=>"101101001",
  43905=>"010101100",
  43906=>"100110101",
  43907=>"110011101",
  43908=>"111001000",
  43909=>"000001011",
  43910=>"011101001",
  43911=>"000111101",
  43912=>"110110010",
  43913=>"011110110",
  43914=>"000101101",
  43915=>"011000000",
  43916=>"110101101",
  43917=>"111110111",
  43918=>"000100100",
  43919=>"111010100",
  43920=>"100110100",
  43921=>"110001100",
  43922=>"011010111",
  43923=>"100110010",
  43924=>"001001000",
  43925=>"010110110",
  43926=>"100000110",
  43927=>"101111111",
  43928=>"001010110",
  43929=>"000001011",
  43930=>"111101010",
  43931=>"111101001",
  43932=>"000001101",
  43933=>"011111101",
  43934=>"010010100",
  43935=>"001111000",
  43936=>"100100101",
  43937=>"011111000",
  43938=>"001001011",
  43939=>"010010000",
  43940=>"100001111",
  43941=>"101110010",
  43942=>"110101100",
  43943=>"100010010",
  43944=>"011010011",
  43945=>"001100101",
  43946=>"110010001",
  43947=>"011100000",
  43948=>"000001110",
  43949=>"110010001",
  43950=>"110100010",
  43951=>"101110010",
  43952=>"011111110",
  43953=>"000011011",
  43954=>"111011111",
  43955=>"001100001",
  43956=>"110001110",
  43957=>"011011110",
  43958=>"111110111",
  43959=>"001011011",
  43960=>"110011110",
  43961=>"110110000",
  43962=>"100110010",
  43963=>"000001100",
  43964=>"000100011",
  43965=>"100001010",
  43966=>"001000110",
  43967=>"000010011",
  43968=>"010111111",
  43969=>"010001010",
  43970=>"110110100",
  43971=>"111001011",
  43972=>"110000111",
  43973=>"010100010",
  43974=>"100111110",
  43975=>"110011101",
  43976=>"000011001",
  43977=>"110010011",
  43978=>"001010010",
  43979=>"100101001",
  43980=>"010110111",
  43981=>"101000000",
  43982=>"010110110",
  43983=>"001001011",
  43984=>"010001100",
  43985=>"110000011",
  43986=>"011001010",
  43987=>"001111011",
  43988=>"100100010",
  43989=>"110100011",
  43990=>"110001111",
  43991=>"000111010",
  43992=>"011001111",
  43993=>"000110110",
  43994=>"000001010",
  43995=>"111010001",
  43996=>"001001010",
  43997=>"110001001",
  43998=>"001111011",
  43999=>"000000011",
  44000=>"101001111",
  44001=>"000000111",
  44002=>"111010011",
  44003=>"010010110",
  44004=>"011001000",
  44005=>"110100001",
  44006=>"000110111",
  44007=>"011000010",
  44008=>"001000011",
  44009=>"100001100",
  44010=>"010010111",
  44011=>"000010001",
  44012=>"010111010",
  44013=>"100111000",
  44014=>"010111000",
  44015=>"111011110",
  44016=>"001001100",
  44017=>"111001110",
  44018=>"101110111",
  44019=>"000001010",
  44020=>"010111011",
  44021=>"111001100",
  44022=>"011010010",
  44023=>"101001100",
  44024=>"100101100",
  44025=>"111010010",
  44026=>"011101110",
  44027=>"111100100",
  44028=>"101111001",
  44029=>"101001001",
  44030=>"110000110",
  44031=>"101101101",
  44032=>"011000101",
  44033=>"011011110",
  44034=>"100011110",
  44035=>"110111110",
  44036=>"001000011",
  44037=>"100010000",
  44038=>"100111001",
  44039=>"110110010",
  44040=>"111110010",
  44041=>"110010110",
  44042=>"011011000",
  44043=>"101000101",
  44044=>"010001110",
  44045=>"001111010",
  44046=>"110110011",
  44047=>"111001111",
  44048=>"101001110",
  44049=>"111111011",
  44050=>"111010011",
  44051=>"001011010",
  44052=>"111011000",
  44053=>"101011010",
  44054=>"011100101",
  44055=>"101101110",
  44056=>"110101000",
  44057=>"100111110",
  44058=>"111101001",
  44059=>"000011100",
  44060=>"000000100",
  44061=>"011100111",
  44062=>"001010011",
  44063=>"111011001",
  44064=>"110101100",
  44065=>"111101100",
  44066=>"100001111",
  44067=>"011110000",
  44068=>"010010000",
  44069=>"110101110",
  44070=>"101011111",
  44071=>"010001001",
  44072=>"010101010",
  44073=>"110011011",
  44074=>"001001110",
  44075=>"111101110",
  44076=>"010011001",
  44077=>"100011100",
  44078=>"110110101",
  44079=>"100100101",
  44080=>"101001111",
  44081=>"101111100",
  44082=>"000011110",
  44083=>"000111001",
  44084=>"001110101",
  44085=>"101100011",
  44086=>"001000010",
  44087=>"100100111",
  44088=>"100110111",
  44089=>"111000000",
  44090=>"110110111",
  44091=>"011000011",
  44092=>"111101011",
  44093=>"000111101",
  44094=>"101101000",
  44095=>"100010011",
  44096=>"111001110",
  44097=>"101101000",
  44098=>"011001011",
  44099=>"101101011",
  44100=>"111011100",
  44101=>"111110111",
  44102=>"101110111",
  44103=>"110011001",
  44104=>"110011110",
  44105=>"001000010",
  44106=>"101101100",
  44107=>"001011010",
  44108=>"101110100",
  44109=>"100110100",
  44110=>"010101110",
  44111=>"011111010",
  44112=>"110111000",
  44113=>"000011000",
  44114=>"111001011",
  44115=>"100111101",
  44116=>"101110011",
  44117=>"101101101",
  44118=>"101111000",
  44119=>"001100101",
  44120=>"011100100",
  44121=>"010000100",
  44122=>"100111100",
  44123=>"100110100",
  44124=>"101111011",
  44125=>"101100001",
  44126=>"010111000",
  44127=>"001110111",
  44128=>"010101000",
  44129=>"000010001",
  44130=>"110110110",
  44131=>"101000100",
  44132=>"010100100",
  44133=>"001110010",
  44134=>"111100111",
  44135=>"001011011",
  44136=>"101100101",
  44137=>"101010110",
  44138=>"001100010",
  44139=>"111000011",
  44140=>"001000100",
  44141=>"101111100",
  44142=>"111100011",
  44143=>"101000101",
  44144=>"010010101",
  44145=>"001100011",
  44146=>"111010110",
  44147=>"000011010",
  44148=>"011100110",
  44149=>"100011111",
  44150=>"011111010",
  44151=>"111100101",
  44152=>"110011100",
  44153=>"010001110",
  44154=>"111111001",
  44155=>"001111101",
  44156=>"011001001",
  44157=>"010101010",
  44158=>"111011101",
  44159=>"101000100",
  44160=>"001010111",
  44161=>"010100101",
  44162=>"000010001",
  44163=>"110111011",
  44164=>"100011111",
  44165=>"101111101",
  44166=>"001001010",
  44167=>"101110100",
  44168=>"001010110",
  44169=>"110111010",
  44170=>"101001111",
  44171=>"000010110",
  44172=>"000000100",
  44173=>"100100110",
  44174=>"100100100",
  44175=>"101001110",
  44176=>"000001000",
  44177=>"010111100",
  44178=>"010110111",
  44179=>"000011000",
  44180=>"000010000",
  44181=>"001011100",
  44182=>"010110000",
  44183=>"010000000",
  44184=>"101011111",
  44185=>"000110000",
  44186=>"010001000",
  44187=>"101111100",
  44188=>"011000111",
  44189=>"111101001",
  44190=>"110110110",
  44191=>"100000000",
  44192=>"101010010",
  44193=>"111111101",
  44194=>"000010101",
  44195=>"100000000",
  44196=>"110010011",
  44197=>"011101010",
  44198=>"000000000",
  44199=>"001110001",
  44200=>"111011101",
  44201=>"000011111",
  44202=>"100000110",
  44203=>"000000000",
  44204=>"100101110",
  44205=>"010101101",
  44206=>"110011010",
  44207=>"101101010",
  44208=>"000000101",
  44209=>"110010010",
  44210=>"101111011",
  44211=>"000000110",
  44212=>"010001101",
  44213=>"001010100",
  44214=>"110011101",
  44215=>"001100101",
  44216=>"001001100",
  44217=>"000010110",
  44218=>"010000100",
  44219=>"001110101",
  44220=>"001100111",
  44221=>"111000101",
  44222=>"000110011",
  44223=>"100010011",
  44224=>"000100110",
  44225=>"001100011",
  44226=>"101111011",
  44227=>"111010111",
  44228=>"000010001",
  44229=>"111101011",
  44230=>"010101111",
  44231=>"110010100",
  44232=>"001010001",
  44233=>"010110111",
  44234=>"100000011",
  44235=>"100111010",
  44236=>"101000100",
  44237=>"100110000",
  44238=>"011100110",
  44239=>"111110110",
  44240=>"101001001",
  44241=>"100101101",
  44242=>"000000110",
  44243=>"100001100",
  44244=>"100010111",
  44245=>"011111010",
  44246=>"001100010",
  44247=>"111100000",
  44248=>"000101110",
  44249=>"001000010",
  44250=>"111110110",
  44251=>"111001010",
  44252=>"110100110",
  44253=>"110010011",
  44254=>"000100111",
  44255=>"111100000",
  44256=>"111111110",
  44257=>"001010101",
  44258=>"011010111",
  44259=>"011011000",
  44260=>"111011100",
  44261=>"010010010",
  44262=>"111010000",
  44263=>"100010010",
  44264=>"110111000",
  44265=>"110100001",
  44266=>"110110001",
  44267=>"101101101",
  44268=>"110101010",
  44269=>"101110101",
  44270=>"111101010",
  44271=>"000111111",
  44272=>"101111000",
  44273=>"000111011",
  44274=>"011000001",
  44275=>"101001111",
  44276=>"010010110",
  44277=>"111101101",
  44278=>"110001010",
  44279=>"011100110",
  44280=>"010001100",
  44281=>"110101010",
  44282=>"010001110",
  44283=>"011100100",
  44284=>"110010010",
  44285=>"000100110",
  44286=>"001111101",
  44287=>"010001101",
  44288=>"111110001",
  44289=>"011011101",
  44290=>"111000101",
  44291=>"011101000",
  44292=>"101001100",
  44293=>"100010000",
  44294=>"111000010",
  44295=>"111001100",
  44296=>"111111101",
  44297=>"000010100",
  44298=>"000010011",
  44299=>"010001110",
  44300=>"010111101",
  44301=>"101000011",
  44302=>"001100101",
  44303=>"000111001",
  44304=>"101101001",
  44305=>"001001001",
  44306=>"000011110",
  44307=>"101011100",
  44308=>"110100011",
  44309=>"000001001",
  44310=>"010000010",
  44311=>"101101011",
  44312=>"101111110",
  44313=>"010110101",
  44314=>"000000001",
  44315=>"101111000",
  44316=>"001001111",
  44317=>"100010101",
  44318=>"111010100",
  44319=>"111011111",
  44320=>"101100110",
  44321=>"001110111",
  44322=>"111100001",
  44323=>"111001111",
  44324=>"010010100",
  44325=>"100011010",
  44326=>"001000111",
  44327=>"100110001",
  44328=>"110010010",
  44329=>"110000000",
  44330=>"100111110",
  44331=>"110110111",
  44332=>"010010110",
  44333=>"000010000",
  44334=>"000001101",
  44335=>"110001111",
  44336=>"101101111",
  44337=>"100111011",
  44338=>"101000000",
  44339=>"100010101",
  44340=>"100011010",
  44341=>"101100101",
  44342=>"011101110",
  44343=>"010101010",
  44344=>"101100110",
  44345=>"000000101",
  44346=>"111100101",
  44347=>"101111110",
  44348=>"001111110",
  44349=>"110110011",
  44350=>"111101001",
  44351=>"011001011",
  44352=>"011100110",
  44353=>"111000000",
  44354=>"010110100",
  44355=>"101000110",
  44356=>"110010101",
  44357=>"000001101",
  44358=>"110001000",
  44359=>"100000001",
  44360=>"101001111",
  44361=>"000001010",
  44362=>"111001100",
  44363=>"110000111",
  44364=>"100101111",
  44365=>"110010100",
  44366=>"111110011",
  44367=>"111001001",
  44368=>"110110011",
  44369=>"000111010",
  44370=>"010000001",
  44371=>"011111000",
  44372=>"110100110",
  44373=>"010101010",
  44374=>"000100100",
  44375=>"000100111",
  44376=>"010000001",
  44377=>"000010110",
  44378=>"000011010",
  44379=>"110001100",
  44380=>"110001001",
  44381=>"100010110",
  44382=>"101011011",
  44383=>"100010000",
  44384=>"010110001",
  44385=>"001001001",
  44386=>"000111101",
  44387=>"100011100",
  44388=>"011001100",
  44389=>"110000011",
  44390=>"111101100",
  44391=>"001000101",
  44392=>"100101011",
  44393=>"000011000",
  44394=>"111011111",
  44395=>"000100000",
  44396=>"100000111",
  44397=>"110110011",
  44398=>"110001110",
  44399=>"010110000",
  44400=>"011001000",
  44401=>"110010100",
  44402=>"101111111",
  44403=>"111001100",
  44404=>"101010101",
  44405=>"110101100",
  44406=>"111110001",
  44407=>"101011101",
  44408=>"011011010",
  44409=>"100000111",
  44410=>"011111101",
  44411=>"100010011",
  44412=>"011010010",
  44413=>"110011101",
  44414=>"101110011",
  44415=>"100100001",
  44416=>"010010100",
  44417=>"101001100",
  44418=>"110111101",
  44419=>"101110100",
  44420=>"110000111",
  44421=>"110100001",
  44422=>"111110001",
  44423=>"111111110",
  44424=>"011101001",
  44425=>"001101110",
  44426=>"000011010",
  44427=>"110111110",
  44428=>"110111111",
  44429=>"001011001",
  44430=>"101101100",
  44431=>"101001001",
  44432=>"110101110",
  44433=>"000101000",
  44434=>"100001101",
  44435=>"100000100",
  44436=>"010111100",
  44437=>"110101000",
  44438=>"100111111",
  44439=>"000001010",
  44440=>"010101101",
  44441=>"000111000",
  44442=>"001001011",
  44443=>"000001001",
  44444=>"100011000",
  44445=>"000110111",
  44446=>"010101100",
  44447=>"111111100",
  44448=>"000011110",
  44449=>"001011111",
  44450=>"110000101",
  44451=>"000000110",
  44452=>"001100110",
  44453=>"000010110",
  44454=>"000000111",
  44455=>"001110110",
  44456=>"101010000",
  44457=>"100011101",
  44458=>"101101110",
  44459=>"110110010",
  44460=>"001110111",
  44461=>"000110000",
  44462=>"110011010",
  44463=>"111101101",
  44464=>"111111110",
  44465=>"000101000",
  44466=>"110010111",
  44467=>"111010110",
  44468=>"011110100",
  44469=>"111000101",
  44470=>"100010100",
  44471=>"011110111",
  44472=>"010111010",
  44473=>"001011110",
  44474=>"111100110",
  44475=>"111100001",
  44476=>"000010100",
  44477=>"101011110",
  44478=>"001111110",
  44479=>"110111101",
  44480=>"001011011",
  44481=>"010011001",
  44482=>"110110010",
  44483=>"010110111",
  44484=>"101010111",
  44485=>"000010110",
  44486=>"100110111",
  44487=>"011111011",
  44488=>"100100100",
  44489=>"010000101",
  44490=>"010001011",
  44491=>"011100110",
  44492=>"000001110",
  44493=>"100110100",
  44494=>"000101111",
  44495=>"110111100",
  44496=>"111010011",
  44497=>"100110111",
  44498=>"001010111",
  44499=>"100101001",
  44500=>"111101111",
  44501=>"000100110",
  44502=>"101100110",
  44503=>"101110000",
  44504=>"010110011",
  44505=>"100100111",
  44506=>"100001110",
  44507=>"000100000",
  44508=>"011100100",
  44509=>"011100011",
  44510=>"011101010",
  44511=>"111000000",
  44512=>"000000001",
  44513=>"111010000",
  44514=>"010000000",
  44515=>"000111000",
  44516=>"110011110",
  44517=>"001100010",
  44518=>"010101010",
  44519=>"111100001",
  44520=>"001111000",
  44521=>"001010100",
  44522=>"010000100",
  44523=>"011010101",
  44524=>"101100011",
  44525=>"101000000",
  44526=>"111011100",
  44527=>"010100100",
  44528=>"111110011",
  44529=>"010110110",
  44530=>"000010011",
  44531=>"001001000",
  44532=>"110011110",
  44533=>"000100100",
  44534=>"011110101",
  44535=>"111100101",
  44536=>"100111110",
  44537=>"011011000",
  44538=>"000111001",
  44539=>"010000110",
  44540=>"111010100",
  44541=>"000001100",
  44542=>"001011001",
  44543=>"000111001",
  44544=>"001000011",
  44545=>"111111010",
  44546=>"000100010",
  44547=>"011101110",
  44548=>"110001111",
  44549=>"011001101",
  44550=>"000100010",
  44551=>"001010000",
  44552=>"001111000",
  44553=>"100011111",
  44554=>"011100000",
  44555=>"110101110",
  44556=>"110001110",
  44557=>"110001010",
  44558=>"000000110",
  44559=>"110111101",
  44560=>"010100110",
  44561=>"111101011",
  44562=>"001111101",
  44563=>"100001110",
  44564=>"101101111",
  44565=>"110001011",
  44566=>"010110100",
  44567=>"110011101",
  44568=>"001010000",
  44569=>"100010110",
  44570=>"100010111",
  44571=>"110100000",
  44572=>"101001100",
  44573=>"001011100",
  44574=>"100000110",
  44575=>"001101110",
  44576=>"111111001",
  44577=>"110010101",
  44578=>"100100111",
  44579=>"110001110",
  44580=>"000000011",
  44581=>"110010111",
  44582=>"110111111",
  44583=>"001010010",
  44584=>"010001000",
  44585=>"010111010",
  44586=>"100100100",
  44587=>"111001000",
  44588=>"111101101",
  44589=>"101000010",
  44590=>"111100101",
  44591=>"110101001",
  44592=>"101000000",
  44593=>"010101100",
  44594=>"001000001",
  44595=>"111110101",
  44596=>"001110011",
  44597=>"110000111",
  44598=>"110011000",
  44599=>"110101111",
  44600=>"011110001",
  44601=>"010001010",
  44602=>"111101000",
  44603=>"111001001",
  44604=>"101001100",
  44605=>"011101000",
  44606=>"011001001",
  44607=>"011001110",
  44608=>"101110101",
  44609=>"110111111",
  44610=>"011100100",
  44611=>"100011000",
  44612=>"010001100",
  44613=>"110011111",
  44614=>"001101101",
  44615=>"101111000",
  44616=>"100011000",
  44617=>"000000000",
  44618=>"001101000",
  44619=>"000101110",
  44620=>"110001001",
  44621=>"100100010",
  44622=>"101011100",
  44623=>"001111010",
  44624=>"110001000",
  44625=>"100010111",
  44626=>"111110111",
  44627=>"001101011",
  44628=>"110011011",
  44629=>"010011101",
  44630=>"011011101",
  44631=>"011111111",
  44632=>"010100101",
  44633=>"001001101",
  44634=>"100111110",
  44635=>"001110100",
  44636=>"110001011",
  44637=>"001100111",
  44638=>"100111000",
  44639=>"010111100",
  44640=>"011110100",
  44641=>"000100010",
  44642=>"111100000",
  44643=>"111000000",
  44644=>"001100110",
  44645=>"011101000",
  44646=>"100000110",
  44647=>"011001010",
  44648=>"011011000",
  44649=>"110001000",
  44650=>"101011101",
  44651=>"000000010",
  44652=>"111111011",
  44653=>"000011011",
  44654=>"101100010",
  44655=>"100010001",
  44656=>"111111111",
  44657=>"010011001",
  44658=>"001000101",
  44659=>"110101011",
  44660=>"011101011",
  44661=>"110110110",
  44662=>"101100110",
  44663=>"011100111",
  44664=>"101001011",
  44665=>"100000110",
  44666=>"110010111",
  44667=>"100000010",
  44668=>"100011100",
  44669=>"010011111",
  44670=>"110001010",
  44671=>"111111001",
  44672=>"101101010",
  44673=>"100101000",
  44674=>"111101101",
  44675=>"010010011",
  44676=>"100001011",
  44677=>"110110111",
  44678=>"100011100",
  44679=>"100001101",
  44680=>"011001100",
  44681=>"100010110",
  44682=>"101000000",
  44683=>"100111010",
  44684=>"011001010",
  44685=>"010001011",
  44686=>"011011010",
  44687=>"101001110",
  44688=>"001101111",
  44689=>"101100000",
  44690=>"001101000",
  44691=>"100111100",
  44692=>"000010111",
  44693=>"011000111",
  44694=>"111011000",
  44695=>"101011011",
  44696=>"110010010",
  44697=>"000101100",
  44698=>"101000111",
  44699=>"011000001",
  44700=>"011100100",
  44701=>"101010011",
  44702=>"010000000",
  44703=>"011001010",
  44704=>"010001010",
  44705=>"010000110",
  44706=>"010000000",
  44707=>"000011100",
  44708=>"110111110",
  44709=>"111111101",
  44710=>"110011011",
  44711=>"101000000",
  44712=>"000000000",
  44713=>"000101001",
  44714=>"000111101",
  44715=>"001000010",
  44716=>"101100010",
  44717=>"000000000",
  44718=>"111101101",
  44719=>"111011111",
  44720=>"111001100",
  44721=>"110010110",
  44722=>"011000100",
  44723=>"110000100",
  44724=>"010011010",
  44725=>"100111001",
  44726=>"110101101",
  44727=>"100101111",
  44728=>"110100000",
  44729=>"111110001",
  44730=>"100000000",
  44731=>"001101101",
  44732=>"101111110",
  44733=>"110001111",
  44734=>"100111100",
  44735=>"100110100",
  44736=>"111001000",
  44737=>"110010101",
  44738=>"010010110",
  44739=>"100000001",
  44740=>"001101100",
  44741=>"000000000",
  44742=>"101111000",
  44743=>"100010000",
  44744=>"011110011",
  44745=>"000000000",
  44746=>"000010001",
  44747=>"100001101",
  44748=>"100101111",
  44749=>"001000000",
  44750=>"000010101",
  44751=>"111010111",
  44752=>"111011001",
  44753=>"001110010",
  44754=>"010100100",
  44755=>"111011101",
  44756=>"001011001",
  44757=>"001100000",
  44758=>"010001001",
  44759=>"000110101",
  44760=>"100011100",
  44761=>"110010100",
  44762=>"111010110",
  44763=>"110100001",
  44764=>"110110110",
  44765=>"000010000",
  44766=>"010110101",
  44767=>"001011111",
  44768=>"000100001",
  44769=>"000001111",
  44770=>"111110111",
  44771=>"010101011",
  44772=>"000011111",
  44773=>"011101110",
  44774=>"101101000",
  44775=>"111111101",
  44776=>"111000101",
  44777=>"010111100",
  44778=>"001000000",
  44779=>"001110011",
  44780=>"001111000",
  44781=>"001010010",
  44782=>"101000101",
  44783=>"000101101",
  44784=>"000110001",
  44785=>"110000111",
  44786=>"100001100",
  44787=>"111000100",
  44788=>"111010011",
  44789=>"010111001",
  44790=>"001011100",
  44791=>"000000101",
  44792=>"111111010",
  44793=>"100000010",
  44794=>"111111000",
  44795=>"011110100",
  44796=>"110100011",
  44797=>"001100001",
  44798=>"000001001",
  44799=>"100011110",
  44800=>"000000101",
  44801=>"101101110",
  44802=>"111011111",
  44803=>"000111010",
  44804=>"100001110",
  44805=>"110010001",
  44806=>"111100101",
  44807=>"001011111",
  44808=>"111001010",
  44809=>"010110000",
  44810=>"111101010",
  44811=>"101010001",
  44812=>"100100001",
  44813=>"010010000",
  44814=>"011100000",
  44815=>"000000010",
  44816=>"100010011",
  44817=>"110010110",
  44818=>"000011111",
  44819=>"001111001",
  44820=>"010011011",
  44821=>"110011101",
  44822=>"010001001",
  44823=>"100000111",
  44824=>"101101001",
  44825=>"111011101",
  44826=>"111110011",
  44827=>"010011101",
  44828=>"001100110",
  44829=>"000101101",
  44830=>"001111110",
  44831=>"010000111",
  44832=>"100011110",
  44833=>"001001110",
  44834=>"110101111",
  44835=>"011110011",
  44836=>"001010110",
  44837=>"000101110",
  44838=>"110110000",
  44839=>"110011000",
  44840=>"001111001",
  44841=>"011000001",
  44842=>"110100011",
  44843=>"111111111",
  44844=>"000111100",
  44845=>"000111010",
  44846=>"111001001",
  44847=>"010100011",
  44848=>"110111010",
  44849=>"001000011",
  44850=>"001111000",
  44851=>"000001001",
  44852=>"101101100",
  44853=>"001000000",
  44854=>"101010010",
  44855=>"001011110",
  44856=>"011111000",
  44857=>"100100101",
  44858=>"110100100",
  44859=>"011100110",
  44860=>"100100101",
  44861=>"100001101",
  44862=>"010001010",
  44863=>"000011001",
  44864=>"001100010",
  44865=>"111110010",
  44866=>"110000100",
  44867=>"011000100",
  44868=>"000001000",
  44869=>"001101101",
  44870=>"010001001",
  44871=>"001101110",
  44872=>"010010000",
  44873=>"101001111",
  44874=>"010000010",
  44875=>"011010000",
  44876=>"110110001",
  44877=>"110101110",
  44878=>"011010001",
  44879=>"001011110",
  44880=>"101011011",
  44881=>"010110110",
  44882=>"110111111",
  44883=>"000000000",
  44884=>"110001011",
  44885=>"010010101",
  44886=>"000011001",
  44887=>"101011001",
  44888=>"000110000",
  44889=>"011010000",
  44890=>"101011010",
  44891=>"000101111",
  44892=>"000011110",
  44893=>"101001010",
  44894=>"110010111",
  44895=>"110011110",
  44896=>"110001011",
  44897=>"110000011",
  44898=>"111100101",
  44899=>"111100010",
  44900=>"110110111",
  44901=>"101101001",
  44902=>"101011110",
  44903=>"110011101",
  44904=>"010111001",
  44905=>"100110101",
  44906=>"100010001",
  44907=>"010111101",
  44908=>"110110111",
  44909=>"110110110",
  44910=>"011010011",
  44911=>"100101111",
  44912=>"100000111",
  44913=>"010010110",
  44914=>"111110100",
  44915=>"100010001",
  44916=>"001001111",
  44917=>"101100011",
  44918=>"000110100",
  44919=>"000011010",
  44920=>"000000111",
  44921=>"110111111",
  44922=>"011000000",
  44923=>"011110111",
  44924=>"101011001",
  44925=>"001100010",
  44926=>"010010001",
  44927=>"111011111",
  44928=>"110100001",
  44929=>"111001110",
  44930=>"101011000",
  44931=>"000110010",
  44932=>"010101001",
  44933=>"100110000",
  44934=>"000111111",
  44935=>"110111110",
  44936=>"011101001",
  44937=>"001100010",
  44938=>"011110010",
  44939=>"110010111",
  44940=>"011100110",
  44941=>"101000111",
  44942=>"111110000",
  44943=>"101011011",
  44944=>"101101101",
  44945=>"111001000",
  44946=>"001111000",
  44947=>"101110110",
  44948=>"111001001",
  44949=>"000111110",
  44950=>"001001010",
  44951=>"111101010",
  44952=>"100100111",
  44953=>"001101111",
  44954=>"111111001",
  44955=>"011011100",
  44956=>"110100110",
  44957=>"010000001",
  44958=>"001011010",
  44959=>"000100110",
  44960=>"000011000",
  44961=>"011101111",
  44962=>"010000101",
  44963=>"110000110",
  44964=>"110101011",
  44965=>"111111001",
  44966=>"110110001",
  44967=>"111111111",
  44968=>"101101001",
  44969=>"001011111",
  44970=>"101011100",
  44971=>"010100011",
  44972=>"011101101",
  44973=>"010011110",
  44974=>"100010001",
  44975=>"010110110",
  44976=>"111011110",
  44977=>"010100011",
  44978=>"000101001",
  44979=>"010000010",
  44980=>"000010111",
  44981=>"111111100",
  44982=>"110110111",
  44983=>"100101000",
  44984=>"000010111",
  44985=>"010001111",
  44986=>"110001101",
  44987=>"110100000",
  44988=>"011000101",
  44989=>"000010101",
  44990=>"100111111",
  44991=>"010001100",
  44992=>"000100010",
  44993=>"111110111",
  44994=>"110110110",
  44995=>"110100111",
  44996=>"001100110",
  44997=>"111000110",
  44998=>"100010100",
  44999=>"100100101",
  45000=>"010000110",
  45001=>"111100011",
  45002=>"000000001",
  45003=>"011111011",
  45004=>"011000000",
  45005=>"001000110",
  45006=>"010110101",
  45007=>"001001110",
  45008=>"100010011",
  45009=>"000101001",
  45010=>"001110101",
  45011=>"000001000",
  45012=>"000001001",
  45013=>"101100000",
  45014=>"001010101",
  45015=>"101101110",
  45016=>"010011001",
  45017=>"010001000",
  45018=>"001111101",
  45019=>"101011000",
  45020=>"111110000",
  45021=>"101001101",
  45022=>"010010010",
  45023=>"001001101",
  45024=>"000010111",
  45025=>"100010001",
  45026=>"101011000",
  45027=>"100100101",
  45028=>"000101100",
  45029=>"110011001",
  45030=>"001000000",
  45031=>"110110111",
  45032=>"001101000",
  45033=>"011011000",
  45034=>"010101101",
  45035=>"001110000",
  45036=>"001110110",
  45037=>"110101110",
  45038=>"000010001",
  45039=>"010111010",
  45040=>"100110100",
  45041=>"110110001",
  45042=>"100000000",
  45043=>"000110110",
  45044=>"000110111",
  45045=>"000010011",
  45046=>"011000010",
  45047=>"011011100",
  45048=>"110111101",
  45049=>"001111111",
  45050=>"111100011",
  45051=>"010100001",
  45052=>"100010010",
  45053=>"101101000",
  45054=>"010010001",
  45055=>"000000001",
  45056=>"110111001",
  45057=>"001110111",
  45058=>"010000001",
  45059=>"111101011",
  45060=>"101010101",
  45061=>"010100100",
  45062=>"011110101",
  45063=>"010001000",
  45064=>"100100001",
  45065=>"101101100",
  45066=>"011100000",
  45067=>"111110010",
  45068=>"001111101",
  45069=>"000101100",
  45070=>"101110001",
  45071=>"000110010",
  45072=>"011001010",
  45073=>"100000110",
  45074=>"111100001",
  45075=>"011010110",
  45076=>"010111011",
  45077=>"011101001",
  45078=>"010011101",
  45079=>"000010011",
  45080=>"111101100",
  45081=>"100100000",
  45082=>"100000010",
  45083=>"100100011",
  45084=>"101111000",
  45085=>"101111010",
  45086=>"001111111",
  45087=>"101011111",
  45088=>"100100010",
  45089=>"010000011",
  45090=>"011001111",
  45091=>"110001011",
  45092=>"101011001",
  45093=>"111010011",
  45094=>"110000000",
  45095=>"110111010",
  45096=>"100111010",
  45097=>"010011001",
  45098=>"111010000",
  45099=>"100001010",
  45100=>"011001010",
  45101=>"110001100",
  45102=>"010011111",
  45103=>"000000111",
  45104=>"101000011",
  45105=>"010011110",
  45106=>"011110010",
  45107=>"011000011",
  45108=>"100111110",
  45109=>"100011000",
  45110=>"011000001",
  45111=>"011010001",
  45112=>"000111101",
  45113=>"100001110",
  45114=>"010001101",
  45115=>"011111011",
  45116=>"011100110",
  45117=>"110111010",
  45118=>"100011111",
  45119=>"110011000",
  45120=>"000011011",
  45121=>"000110110",
  45122=>"010000011",
  45123=>"010001010",
  45124=>"101111000",
  45125=>"010001100",
  45126=>"100110000",
  45127=>"100111100",
  45128=>"000110100",
  45129=>"110010000",
  45130=>"111101001",
  45131=>"001101000",
  45132=>"001111100",
  45133=>"110011110",
  45134=>"110000000",
  45135=>"100111010",
  45136=>"100001001",
  45137=>"001011110",
  45138=>"110111010",
  45139=>"111011110",
  45140=>"000000011",
  45141=>"101011011",
  45142=>"100011111",
  45143=>"100111000",
  45144=>"001001001",
  45145=>"100001101",
  45146=>"101011110",
  45147=>"010101001",
  45148=>"101100010",
  45149=>"011101000",
  45150=>"100010100",
  45151=>"001010001",
  45152=>"010111011",
  45153=>"010111010",
  45154=>"011001001",
  45155=>"001111000",
  45156=>"011011010",
  45157=>"100011010",
  45158=>"001001001",
  45159=>"001101110",
  45160=>"001110100",
  45161=>"101011010",
  45162=>"010011010",
  45163=>"111011011",
  45164=>"000100110",
  45165=>"100110001",
  45166=>"100101111",
  45167=>"000011111",
  45168=>"001010001",
  45169=>"010001001",
  45170=>"011001111",
  45171=>"110110101",
  45172=>"101110011",
  45173=>"101101010",
  45174=>"001110010",
  45175=>"000001100",
  45176=>"000111110",
  45177=>"011001001",
  45178=>"100001000",
  45179=>"000001001",
  45180=>"000000110",
  45181=>"101001101",
  45182=>"010000001",
  45183=>"111111000",
  45184=>"101000110",
  45185=>"100010011",
  45186=>"110110000",
  45187=>"110101001",
  45188=>"100101001",
  45189=>"110101000",
  45190=>"011101111",
  45191=>"100000101",
  45192=>"001101100",
  45193=>"101010000",
  45194=>"100011010",
  45195=>"111010010",
  45196=>"111000101",
  45197=>"110000111",
  45198=>"101001100",
  45199=>"100001000",
  45200=>"001001010",
  45201=>"000000100",
  45202=>"111100110",
  45203=>"001101011",
  45204=>"000001011",
  45205=>"101011111",
  45206=>"110111100",
  45207=>"110000101",
  45208=>"010100110",
  45209=>"000100110",
  45210=>"101101011",
  45211=>"000001000",
  45212=>"111010011",
  45213=>"110011110",
  45214=>"110001000",
  45215=>"010101000",
  45216=>"011010111",
  45217=>"011001111",
  45218=>"100110100",
  45219=>"111001110",
  45220=>"011000101",
  45221=>"000010100",
  45222=>"101010011",
  45223=>"000110010",
  45224=>"111010111",
  45225=>"100111000",
  45226=>"001111000",
  45227=>"110001111",
  45228=>"010110010",
  45229=>"100101000",
  45230=>"111101000",
  45231=>"111111111",
  45232=>"101110010",
  45233=>"100000100",
  45234=>"101100111",
  45235=>"000100100",
  45236=>"111101010",
  45237=>"110001100",
  45238=>"011101000",
  45239=>"111001000",
  45240=>"111100001",
  45241=>"001011010",
  45242=>"010101000",
  45243=>"000000010",
  45244=>"001010000",
  45245=>"011010111",
  45246=>"000110111",
  45247=>"011101111",
  45248=>"111110101",
  45249=>"111100111",
  45250=>"010010001",
  45251=>"010111111",
  45252=>"001001011",
  45253=>"001010000",
  45254=>"111111110",
  45255=>"101011011",
  45256=>"111010001",
  45257=>"111011100",
  45258=>"111101010",
  45259=>"011010100",
  45260=>"100001000",
  45261=>"100110001",
  45262=>"000010001",
  45263=>"111000110",
  45264=>"101111010",
  45265=>"100000010",
  45266=>"010101110",
  45267=>"100100000",
  45268=>"111101101",
  45269=>"000010011",
  45270=>"100010011",
  45271=>"010011001",
  45272=>"101100001",
  45273=>"000000110",
  45274=>"010100011",
  45275=>"111111000",
  45276=>"101010011",
  45277=>"100100000",
  45278=>"000001111",
  45279=>"101001010",
  45280=>"111000000",
  45281=>"101000011",
  45282=>"011101000",
  45283=>"000011010",
  45284=>"001100111",
  45285=>"000010111",
  45286=>"100000001",
  45287=>"011100000",
  45288=>"001100111",
  45289=>"100010001",
  45290=>"100100001",
  45291=>"001100101",
  45292=>"010100010",
  45293=>"100011100",
  45294=>"010100101",
  45295=>"101001010",
  45296=>"101111001",
  45297=>"100100001",
  45298=>"000010000",
  45299=>"100111110",
  45300=>"011000101",
  45301=>"000110101",
  45302=>"001100101",
  45303=>"111100000",
  45304=>"100011001",
  45305=>"011010000",
  45306=>"000011101",
  45307=>"111001110",
  45308=>"111000110",
  45309=>"110001011",
  45310=>"010000010",
  45311=>"000110111",
  45312=>"010010010",
  45313=>"110101000",
  45314=>"010101010",
  45315=>"000011011",
  45316=>"000101110",
  45317=>"110001000",
  45318=>"001100000",
  45319=>"110010010",
  45320=>"000000000",
  45321=>"011110110",
  45322=>"101000110",
  45323=>"111101101",
  45324=>"110101111",
  45325=>"100000101",
  45326=>"110110110",
  45327=>"011000001",
  45328=>"111101111",
  45329=>"000101011",
  45330=>"010000000",
  45331=>"100101110",
  45332=>"011111111",
  45333=>"101011111",
  45334=>"101000000",
  45335=>"101001100",
  45336=>"100110110",
  45337=>"011111111",
  45338=>"011010011",
  45339=>"110010001",
  45340=>"101000010",
  45341=>"111100010",
  45342=>"110110111",
  45343=>"000101111",
  45344=>"011000110",
  45345=>"000101010",
  45346=>"010011111",
  45347=>"000001100",
  45348=>"000011011",
  45349=>"011001101",
  45350=>"000011100",
  45351=>"110110010",
  45352=>"111000011",
  45353=>"111011100",
  45354=>"111111001",
  45355=>"010000011",
  45356=>"100101010",
  45357=>"111110011",
  45358=>"011000001",
  45359=>"000101001",
  45360=>"110001001",
  45361=>"000110000",
  45362=>"011110010",
  45363=>"000011011",
  45364=>"100010110",
  45365=>"101000101",
  45366=>"011011101",
  45367=>"001100001",
  45368=>"111010111",
  45369=>"101111101",
  45370=>"111000000",
  45371=>"111011010",
  45372=>"001100000",
  45373=>"001110101",
  45374=>"110001110",
  45375=>"000001000",
  45376=>"011111010",
  45377=>"101100110",
  45378=>"101010101",
  45379=>"001000100",
  45380=>"000101010",
  45381=>"010101010",
  45382=>"000100101",
  45383=>"010110010",
  45384=>"110001010",
  45385=>"111101001",
  45386=>"001000000",
  45387=>"101000011",
  45388=>"110100001",
  45389=>"001011100",
  45390=>"100100000",
  45391=>"001111011",
  45392=>"100001000",
  45393=>"101011010",
  45394=>"100000100",
  45395=>"000010100",
  45396=>"000100100",
  45397=>"001010011",
  45398=>"111001011",
  45399=>"011011010",
  45400=>"000000000",
  45401=>"100010101",
  45402=>"000011111",
  45403=>"111100111",
  45404=>"111101101",
  45405=>"101011111",
  45406=>"110100001",
  45407=>"101010001",
  45408=>"100001110",
  45409=>"001001110",
  45410=>"011010001",
  45411=>"000110011",
  45412=>"111101011",
  45413=>"100000110",
  45414=>"110101000",
  45415=>"100001110",
  45416=>"101101001",
  45417=>"100110010",
  45418=>"110111000",
  45419=>"100100001",
  45420=>"001101001",
  45421=>"000100101",
  45422=>"101001111",
  45423=>"100011011",
  45424=>"010001100",
  45425=>"100101111",
  45426=>"101101111",
  45427=>"010000011",
  45428=>"011111011",
  45429=>"101100010",
  45430=>"100001100",
  45431=>"100010110",
  45432=>"010111011",
  45433=>"010011001",
  45434=>"000011101",
  45435=>"000011110",
  45436=>"100111011",
  45437=>"110110100",
  45438=>"110011110",
  45439=>"110100111",
  45440=>"110110000",
  45441=>"000101000",
  45442=>"110101111",
  45443=>"101111000",
  45444=>"011000010",
  45445=>"001111111",
  45446=>"110111000",
  45447=>"101110111",
  45448=>"010010100",
  45449=>"001110101",
  45450=>"001110011",
  45451=>"010110000",
  45452=>"111001111",
  45453=>"011001011",
  45454=>"001110100",
  45455=>"010010110",
  45456=>"111011001",
  45457=>"000101100",
  45458=>"101000011",
  45459=>"100100110",
  45460=>"100000101",
  45461=>"011110000",
  45462=>"111010100",
  45463=>"001011000",
  45464=>"100110100",
  45465=>"100000100",
  45466=>"001111111",
  45467=>"000001101",
  45468=>"110011111",
  45469=>"100111000",
  45470=>"010110111",
  45471=>"001100001",
  45472=>"100100010",
  45473=>"101000000",
  45474=>"111100000",
  45475=>"100101011",
  45476=>"011100011",
  45477=>"111000100",
  45478=>"101001011",
  45479=>"011010010",
  45480=>"001101100",
  45481=>"100111001",
  45482=>"010000110",
  45483=>"111101000",
  45484=>"010010100",
  45485=>"000111110",
  45486=>"011001000",
  45487=>"001110111",
  45488=>"001000101",
  45489=>"110100100",
  45490=>"101111100",
  45491=>"111100001",
  45492=>"111001100",
  45493=>"000001000",
  45494=>"100000111",
  45495=>"101111100",
  45496=>"110100101",
  45497=>"000100000",
  45498=>"100001010",
  45499=>"110010010",
  45500=>"111110111",
  45501=>"011110001",
  45502=>"000101101",
  45503=>"010101001",
  45504=>"100100100",
  45505=>"000010100",
  45506=>"000101000",
  45507=>"100011111",
  45508=>"010011000",
  45509=>"100101000",
  45510=>"000000010",
  45511=>"001010110",
  45512=>"000010111",
  45513=>"000001100",
  45514=>"001001100",
  45515=>"010010000",
  45516=>"011001110",
  45517=>"100100101",
  45518=>"101111100",
  45519=>"001010010",
  45520=>"001001110",
  45521=>"011100111",
  45522=>"011111001",
  45523=>"001000010",
  45524=>"010011110",
  45525=>"101101010",
  45526=>"101010001",
  45527=>"101110110",
  45528=>"111010010",
  45529=>"110011000",
  45530=>"011001001",
  45531=>"100100001",
  45532=>"100010101",
  45533=>"010000110",
  45534=>"111001111",
  45535=>"100000100",
  45536=>"110100010",
  45537=>"001111001",
  45538=>"111111100",
  45539=>"001101001",
  45540=>"101100100",
  45541=>"000000110",
  45542=>"110100110",
  45543=>"010111100",
  45544=>"100100101",
  45545=>"001010110",
  45546=>"101001100",
  45547=>"110101101",
  45548=>"001101011",
  45549=>"101010001",
  45550=>"101100011",
  45551=>"110110010",
  45552=>"000110010",
  45553=>"010110111",
  45554=>"101110110",
  45555=>"010110111",
  45556=>"101011111",
  45557=>"010110110",
  45558=>"001111101",
  45559=>"110101010",
  45560=>"101000000",
  45561=>"111000111",
  45562=>"100101001",
  45563=>"110001101",
  45564=>"110010000",
  45565=>"010000101",
  45566=>"001000001",
  45567=>"010011000",
  45568=>"000000110",
  45569=>"000101100",
  45570=>"011111011",
  45571=>"011001000",
  45572=>"010001011",
  45573=>"011010011",
  45574=>"110110001",
  45575=>"111010001",
  45576=>"011110111",
  45577=>"000100011",
  45578=>"110110001",
  45579=>"101010011",
  45580=>"001010110",
  45581=>"111111001",
  45582=>"010010100",
  45583=>"001000001",
  45584=>"010010010",
  45585=>"010010011",
  45586=>"111101100",
  45587=>"100100110",
  45588=>"111100000",
  45589=>"000001011",
  45590=>"100101001",
  45591=>"111111011",
  45592=>"101110110",
  45593=>"000001100",
  45594=>"000010101",
  45595=>"010000010",
  45596=>"000110000",
  45597=>"100001010",
  45598=>"111101011",
  45599=>"110101111",
  45600=>"001010101",
  45601=>"000100110",
  45602=>"011000001",
  45603=>"001101111",
  45604=>"111100111",
  45605=>"110000101",
  45606=>"010110111",
  45607=>"011111111",
  45608=>"100000000",
  45609=>"101010000",
  45610=>"111100111",
  45611=>"001100101",
  45612=>"110000011",
  45613=>"000110110",
  45614=>"000011111",
  45615=>"000101010",
  45616=>"011001101",
  45617=>"111000101",
  45618=>"000001000",
  45619=>"011000011",
  45620=>"001011101",
  45621=>"110100110",
  45622=>"010111000",
  45623=>"000001000",
  45624=>"111111110",
  45625=>"111001010",
  45626=>"000011101",
  45627=>"000100010",
  45628=>"010001101",
  45629=>"111101011",
  45630=>"101100100",
  45631=>"111011010",
  45632=>"111110000",
  45633=>"010110101",
  45634=>"100001001",
  45635=>"111100010",
  45636=>"100001101",
  45637=>"110000111",
  45638=>"111000101",
  45639=>"010111101",
  45640=>"111010100",
  45641=>"101111111",
  45642=>"110100101",
  45643=>"100010001",
  45644=>"110110000",
  45645=>"110111100",
  45646=>"000110000",
  45647=>"001001011",
  45648=>"101110111",
  45649=>"110010010",
  45650=>"110011110",
  45651=>"000000110",
  45652=>"010001001",
  45653=>"110100000",
  45654=>"001000010",
  45655=>"110001000",
  45656=>"010110011",
  45657=>"001011010",
  45658=>"000110111",
  45659=>"101101010",
  45660=>"100100100",
  45661=>"111010111",
  45662=>"111000000",
  45663=>"010010011",
  45664=>"001010010",
  45665=>"001000010",
  45666=>"011011100",
  45667=>"001111111",
  45668=>"110111001",
  45669=>"101011111",
  45670=>"011000110",
  45671=>"100011101",
  45672=>"001001100",
  45673=>"010110100",
  45674=>"101011100",
  45675=>"101010110",
  45676=>"010100000",
  45677=>"000011011",
  45678=>"001001000",
  45679=>"100010010",
  45680=>"110101010",
  45681=>"111011010",
  45682=>"011010111",
  45683=>"101110111",
  45684=>"010110010",
  45685=>"001000000",
  45686=>"101011110",
  45687=>"001001010",
  45688=>"100100110",
  45689=>"101011100",
  45690=>"000110110",
  45691=>"000010111",
  45692=>"100001100",
  45693=>"101111100",
  45694=>"011100110",
  45695=>"001100011",
  45696=>"001101010",
  45697=>"000000001",
  45698=>"000001000",
  45699=>"000001100",
  45700=>"111010111",
  45701=>"101001100",
  45702=>"110100111",
  45703=>"000001000",
  45704=>"010110101",
  45705=>"000000001",
  45706=>"110111000",
  45707=>"110010110",
  45708=>"000001111",
  45709=>"001100000",
  45710=>"101110000",
  45711=>"111101110",
  45712=>"010010011",
  45713=>"111011111",
  45714=>"000010110",
  45715=>"101001111",
  45716=>"100100100",
  45717=>"001011011",
  45718=>"010000011",
  45719=>"100001000",
  45720=>"100101100",
  45721=>"101011100",
  45722=>"011100100",
  45723=>"101101011",
  45724=>"100111100",
  45725=>"011110110",
  45726=>"100101111",
  45727=>"001011111",
  45728=>"001111111",
  45729=>"101110011",
  45730=>"000111101",
  45731=>"110001011",
  45732=>"110000001",
  45733=>"110011110",
  45734=>"000010100",
  45735=>"100001100",
  45736=>"010000100",
  45737=>"011100011",
  45738=>"010010000",
  45739=>"110011001",
  45740=>"000000001",
  45741=>"000000011",
  45742=>"001001010",
  45743=>"101100011",
  45744=>"001100000",
  45745=>"001000101",
  45746=>"101100001",
  45747=>"101011000",
  45748=>"110101101",
  45749=>"100010101",
  45750=>"001001111",
  45751=>"000111011",
  45752=>"100100011",
  45753=>"110011110",
  45754=>"100000110",
  45755=>"011010011",
  45756=>"110101001",
  45757=>"001010000",
  45758=>"110101010",
  45759=>"000101000",
  45760=>"010111010",
  45761=>"010100100",
  45762=>"101001011",
  45763=>"000001100",
  45764=>"001001110",
  45765=>"111111111",
  45766=>"001111011",
  45767=>"000110101",
  45768=>"101000101",
  45769=>"111010011",
  45770=>"111110101",
  45771=>"000100001",
  45772=>"100110001",
  45773=>"101000110",
  45774=>"111110110",
  45775=>"011000000",
  45776=>"010001111",
  45777=>"001001101",
  45778=>"010000001",
  45779=>"111101001",
  45780=>"100100010",
  45781=>"001111001",
  45782=>"010001101",
  45783=>"000000001",
  45784=>"000000101",
  45785=>"110000100",
  45786=>"001000011",
  45787=>"111000111",
  45788=>"100101001",
  45789=>"010000000",
  45790=>"001010101",
  45791=>"010111101",
  45792=>"101101001",
  45793=>"110001001",
  45794=>"101001010",
  45795=>"010011101",
  45796=>"110100111",
  45797=>"111001001",
  45798=>"101111010",
  45799=>"010011000",
  45800=>"101001011",
  45801=>"110100100",
  45802=>"011011100",
  45803=>"011100110",
  45804=>"011011011",
  45805=>"100111111",
  45806=>"101011100",
  45807=>"101010110",
  45808=>"001110011",
  45809=>"110101011",
  45810=>"100100101",
  45811=>"001101001",
  45812=>"001100011",
  45813=>"110011010",
  45814=>"111111110",
  45815=>"010001000",
  45816=>"000110100",
  45817=>"111100100",
  45818=>"111110001",
  45819=>"101011000",
  45820=>"010010011",
  45821=>"100100100",
  45822=>"000111100",
  45823=>"000110011",
  45824=>"001110110",
  45825=>"100101101",
  45826=>"001111000",
  45827=>"010001100",
  45828=>"011011100",
  45829=>"001011101",
  45830=>"101011100",
  45831=>"000000111",
  45832=>"100111110",
  45833=>"111000100",
  45834=>"100100000",
  45835=>"001011011",
  45836=>"111000100",
  45837=>"101110010",
  45838=>"011001001",
  45839=>"011111011",
  45840=>"000101101",
  45841=>"101001111",
  45842=>"101001000",
  45843=>"110001101",
  45844=>"001101100",
  45845=>"001011000",
  45846=>"111100001",
  45847=>"111001000",
  45848=>"001011011",
  45849=>"000001011",
  45850=>"010101100",
  45851=>"000000111",
  45852=>"001110100",
  45853=>"110111101",
  45854=>"111101000",
  45855=>"100101110",
  45856=>"011100101",
  45857=>"111111111",
  45858=>"100111011",
  45859=>"101011000",
  45860=>"000100111",
  45861=>"111011101",
  45862=>"001001110",
  45863=>"101110000",
  45864=>"100001100",
  45865=>"101001001",
  45866=>"100011100",
  45867=>"011100110",
  45868=>"000011011",
  45869=>"111000001",
  45870=>"100001110",
  45871=>"100100000",
  45872=>"100100101",
  45873=>"101000100",
  45874=>"000111011",
  45875=>"001100010",
  45876=>"101000011",
  45877=>"000100110",
  45878=>"111010100",
  45879=>"010011001",
  45880=>"000011000",
  45881=>"000010010",
  45882=>"011010100",
  45883=>"000001001",
  45884=>"100101111",
  45885=>"100010100",
  45886=>"110101001",
  45887=>"100110111",
  45888=>"101000111",
  45889=>"011011011",
  45890=>"000010101",
  45891=>"100110100",
  45892=>"110001101",
  45893=>"010000111",
  45894=>"101100011",
  45895=>"011101000",
  45896=>"100010101",
  45897=>"110111001",
  45898=>"011000000",
  45899=>"001011001",
  45900=>"101011100",
  45901=>"111000001",
  45902=>"001100010",
  45903=>"000000000",
  45904=>"100000010",
  45905=>"100001000",
  45906=>"010000100",
  45907=>"111111000",
  45908=>"000000000",
  45909=>"010100100",
  45910=>"010101111",
  45911=>"011000100",
  45912=>"001000100",
  45913=>"011100101",
  45914=>"110010111",
  45915=>"011001100",
  45916=>"001010101",
  45917=>"111111111",
  45918=>"011110010",
  45919=>"111110001",
  45920=>"110010001",
  45921=>"011110010",
  45922=>"100111111",
  45923=>"111101110",
  45924=>"100100000",
  45925=>"011001101",
  45926=>"010101100",
  45927=>"000000111",
  45928=>"100011100",
  45929=>"110011110",
  45930=>"111111100",
  45931=>"010110111",
  45932=>"101100110",
  45933=>"101011110",
  45934=>"100010101",
  45935=>"100101001",
  45936=>"010111111",
  45937=>"100011000",
  45938=>"111100011",
  45939=>"101100000",
  45940=>"111010011",
  45941=>"111011010",
  45942=>"110110011",
  45943=>"101111101",
  45944=>"111111011",
  45945=>"000000100",
  45946=>"101000001",
  45947=>"100110010",
  45948=>"010100010",
  45949=>"001010111",
  45950=>"000110100",
  45951=>"111111111",
  45952=>"001111111",
  45953=>"110110110",
  45954=>"101100100",
  45955=>"001000101",
  45956=>"111000110",
  45957=>"010101100",
  45958=>"000000011",
  45959=>"111000011",
  45960=>"011100111",
  45961=>"100010101",
  45962=>"001111100",
  45963=>"001011011",
  45964=>"110101100",
  45965=>"111110011",
  45966=>"110010000",
  45967=>"011100000",
  45968=>"011111001",
  45969=>"001010000",
  45970=>"000110110",
  45971=>"110001010",
  45972=>"011011110",
  45973=>"111110011",
  45974=>"001101011",
  45975=>"110101101",
  45976=>"111110000",
  45977=>"011000111",
  45978=>"000101111",
  45979=>"110100101",
  45980=>"000111010",
  45981=>"101010000",
  45982=>"000011000",
  45983=>"100111100",
  45984=>"111000100",
  45985=>"011111101",
  45986=>"001101110",
  45987=>"111111010",
  45988=>"110110001",
  45989=>"010001101",
  45990=>"111001111",
  45991=>"110110111",
  45992=>"011001000",
  45993=>"100100001",
  45994=>"000110011",
  45995=>"010100100",
  45996=>"101001010",
  45997=>"100111101",
  45998=>"100111001",
  45999=>"000011011",
  46000=>"011010101",
  46001=>"010111010",
  46002=>"011010001",
  46003=>"111110101",
  46004=>"000001001",
  46005=>"010111111",
  46006=>"100001011",
  46007=>"111111000",
  46008=>"011110001",
  46009=>"011101011",
  46010=>"101001001",
  46011=>"001100000",
  46012=>"001001000",
  46013=>"010001010",
  46014=>"101111100",
  46015=>"110001100",
  46016=>"000110110",
  46017=>"000000111",
  46018=>"000111110",
  46019=>"111101010",
  46020=>"010101111",
  46021=>"011001010",
  46022=>"011000110",
  46023=>"000100000",
  46024=>"110001000",
  46025=>"001110101",
  46026=>"011101100",
  46027=>"100010000",
  46028=>"010001011",
  46029=>"110111111",
  46030=>"011010110",
  46031=>"101001000",
  46032=>"010111101",
  46033=>"111111101",
  46034=>"100010111",
  46035=>"000000111",
  46036=>"010011000",
  46037=>"111011011",
  46038=>"011111001",
  46039=>"000100111",
  46040=>"110010011",
  46041=>"111110011",
  46042=>"111101110",
  46043=>"111110011",
  46044=>"011110110",
  46045=>"111111111",
  46046=>"100110011",
  46047=>"011010010",
  46048=>"001101011",
  46049=>"110010100",
  46050=>"011101111",
  46051=>"001111000",
  46052=>"100001000",
  46053=>"101101111",
  46054=>"010111011",
  46055=>"011110001",
  46056=>"010000000",
  46057=>"000101011",
  46058=>"110100110",
  46059=>"110001001",
  46060=>"101101100",
  46061=>"000010010",
  46062=>"000000110",
  46063=>"100000111",
  46064=>"100111001",
  46065=>"101111101",
  46066=>"100101001",
  46067=>"011010000",
  46068=>"110110110",
  46069=>"110110011",
  46070=>"001101100",
  46071=>"111100010",
  46072=>"101101010",
  46073=>"011001000",
  46074=>"010101011",
  46075=>"111101001",
  46076=>"001011101",
  46077=>"001110000",
  46078=>"111000001",
  46079=>"111110001",
  46080=>"000110000",
  46081=>"010000101",
  46082=>"000000111",
  46083=>"100100101",
  46084=>"010011101",
  46085=>"011000000",
  46086=>"000000111",
  46087=>"111101111",
  46088=>"111010001",
  46089=>"001110000",
  46090=>"010001011",
  46091=>"001111001",
  46092=>"100000000",
  46093=>"100110000",
  46094=>"010010000",
  46095=>"010101110",
  46096=>"100111011",
  46097=>"011110110",
  46098=>"001111010",
  46099=>"100110011",
  46100=>"100000000",
  46101=>"111000111",
  46102=>"110110101",
  46103=>"000001100",
  46104=>"100000100",
  46105=>"100111001",
  46106=>"101100101",
  46107=>"101101000",
  46108=>"111110000",
  46109=>"111010000",
  46110=>"101011011",
  46111=>"100111111",
  46112=>"010010101",
  46113=>"100111011",
  46114=>"010011010",
  46115=>"010100001",
  46116=>"000001000",
  46117=>"010010111",
  46118=>"110110110",
  46119=>"011101001",
  46120=>"110010001",
  46121=>"101111001",
  46122=>"000100000",
  46123=>"011101000",
  46124=>"111010101",
  46125=>"010100011",
  46126=>"000101100",
  46127=>"000110100",
  46128=>"100110110",
  46129=>"010000110",
  46130=>"110111001",
  46131=>"100010101",
  46132=>"001000001",
  46133=>"001110001",
  46134=>"000111110",
  46135=>"000011101",
  46136=>"000010111",
  46137=>"011000010",
  46138=>"111001100",
  46139=>"001110010",
  46140=>"011001000",
  46141=>"011010100",
  46142=>"111111010",
  46143=>"000001001",
  46144=>"110100000",
  46145=>"100101100",
  46146=>"010101111",
  46147=>"110011101",
  46148=>"100110110",
  46149=>"111000010",
  46150=>"100100011",
  46151=>"100100100",
  46152=>"100001001",
  46153=>"101000001",
  46154=>"001010011",
  46155=>"110000011",
  46156=>"011011010",
  46157=>"100110010",
  46158=>"100011110",
  46159=>"001001000",
  46160=>"000001101",
  46161=>"011000100",
  46162=>"001101111",
  46163=>"010111000",
  46164=>"110011100",
  46165=>"101011100",
  46166=>"111111110",
  46167=>"111110010",
  46168=>"001101011",
  46169=>"001010000",
  46170=>"011111110",
  46171=>"100000111",
  46172=>"100101010",
  46173=>"000100000",
  46174=>"111101110",
  46175=>"010000111",
  46176=>"000111000",
  46177=>"011000001",
  46178=>"000101110",
  46179=>"010110000",
  46180=>"000101110",
  46181=>"001111000",
  46182=>"110000000",
  46183=>"110111101",
  46184=>"001001110",
  46185=>"110110011",
  46186=>"001111010",
  46187=>"111111001",
  46188=>"111111000",
  46189=>"111010101",
  46190=>"101010100",
  46191=>"010110000",
  46192=>"111100101",
  46193=>"100111000",
  46194=>"110110110",
  46195=>"101010010",
  46196=>"011110100",
  46197=>"000101110",
  46198=>"110011011",
  46199=>"100111100",
  46200=>"101100000",
  46201=>"100100001",
  46202=>"000111010",
  46203=>"100000110",
  46204=>"010111001",
  46205=>"000101010",
  46206=>"010010000",
  46207=>"000000000",
  46208=>"100111111",
  46209=>"111001001",
  46210=>"101101010",
  46211=>"010011100",
  46212=>"111111011",
  46213=>"010100101",
  46214=>"001001010",
  46215=>"001010000",
  46216=>"110011110",
  46217=>"000100111",
  46218=>"000100110",
  46219=>"001110101",
  46220=>"100001100",
  46221=>"111100100",
  46222=>"100100100",
  46223=>"100100000",
  46224=>"011011110",
  46225=>"010111110",
  46226=>"010011110",
  46227=>"110011010",
  46228=>"110010111",
  46229=>"000110101",
  46230=>"110110000",
  46231=>"100000100",
  46232=>"111100101",
  46233=>"110101101",
  46234=>"100001000",
  46235=>"101011111",
  46236=>"000001000",
  46237=>"100001111",
  46238=>"100110010",
  46239=>"111011100",
  46240=>"100101000",
  46241=>"101011111",
  46242=>"111101011",
  46243=>"111110100",
  46244=>"001101001",
  46245=>"001101100",
  46246=>"001111100",
  46247=>"110111001",
  46248=>"000101101",
  46249=>"010001100",
  46250=>"000011111",
  46251=>"001010001",
  46252=>"001011000",
  46253=>"111111110",
  46254=>"111101111",
  46255=>"010111110",
  46256=>"100110001",
  46257=>"011101101",
  46258=>"100101011",
  46259=>"001001110",
  46260=>"001101111",
  46261=>"000100100",
  46262=>"110111001",
  46263=>"011100000",
  46264=>"110101100",
  46265=>"001110111",
  46266=>"011011101",
  46267=>"011101001",
  46268=>"111000111",
  46269=>"000010011",
  46270=>"110100111",
  46271=>"011010011",
  46272=>"000011100",
  46273=>"100010010",
  46274=>"000001010",
  46275=>"110011100",
  46276=>"110011001",
  46277=>"000100111",
  46278=>"110000110",
  46279=>"110111010",
  46280=>"100111111",
  46281=>"011110000",
  46282=>"101111111",
  46283=>"110011110",
  46284=>"001000100",
  46285=>"010000111",
  46286=>"010100010",
  46287=>"101101100",
  46288=>"111101101",
  46289=>"001011010",
  46290=>"001001000",
  46291=>"000110000",
  46292=>"101110111",
  46293=>"000110011",
  46294=>"001000100",
  46295=>"001000000",
  46296=>"110100000",
  46297=>"010110101",
  46298=>"010010000",
  46299=>"100010000",
  46300=>"101010010",
  46301=>"100100110",
  46302=>"001010111",
  46303=>"100101101",
  46304=>"110011101",
  46305=>"000001010",
  46306=>"000000111",
  46307=>"001101000",
  46308=>"101001110",
  46309=>"100000110",
  46310=>"100001011",
  46311=>"110010101",
  46312=>"110010011",
  46313=>"101011101",
  46314=>"001000110",
  46315=>"010110011",
  46316=>"110010110",
  46317=>"011100010",
  46318=>"100001100",
  46319=>"111001101",
  46320=>"101000101",
  46321=>"110101111",
  46322=>"100111110",
  46323=>"001001110",
  46324=>"011110100",
  46325=>"010100011",
  46326=>"011010011",
  46327=>"110001101",
  46328=>"111010000",
  46329=>"010001010",
  46330=>"010110011",
  46331=>"001110000",
  46332=>"101011101",
  46333=>"001100101",
  46334=>"011111111",
  46335=>"001010101",
  46336=>"111000111",
  46337=>"011011110",
  46338=>"010010000",
  46339=>"100001010",
  46340=>"011111111",
  46341=>"011111000",
  46342=>"001111011",
  46343=>"000000001",
  46344=>"111100100",
  46345=>"100111010",
  46346=>"110000101",
  46347=>"101101110",
  46348=>"100111010",
  46349=>"110001011",
  46350=>"110111011",
  46351=>"011000101",
  46352=>"010110111",
  46353=>"101101111",
  46354=>"000010001",
  46355=>"010000011",
  46356=>"001010110",
  46357=>"101010101",
  46358=>"001011011",
  46359=>"000111111",
  46360=>"100011000",
  46361=>"000101101",
  46362=>"011001000",
  46363=>"010100000",
  46364=>"100010111",
  46365=>"001111010",
  46366=>"000100001",
  46367=>"111110101",
  46368=>"010101100",
  46369=>"111111010",
  46370=>"010101110",
  46371=>"010101001",
  46372=>"110101001",
  46373=>"010000101",
  46374=>"010010110",
  46375=>"010000001",
  46376=>"100011111",
  46377=>"001101010",
  46378=>"010101101",
  46379=>"011110111",
  46380=>"111100111",
  46381=>"010110000",
  46382=>"100001100",
  46383=>"101111001",
  46384=>"001010110",
  46385=>"011110001",
  46386=>"111111110",
  46387=>"111000101",
  46388=>"010000001",
  46389=>"001111010",
  46390=>"111001011",
  46391=>"000110000",
  46392=>"111001111",
  46393=>"001110100",
  46394=>"001000000",
  46395=>"111000010",
  46396=>"101110001",
  46397=>"010100111",
  46398=>"010011010",
  46399=>"011010011",
  46400=>"000010000",
  46401=>"000010001",
  46402=>"011001000",
  46403=>"110010011",
  46404=>"000110011",
  46405=>"001001101",
  46406=>"000111100",
  46407=>"100110000",
  46408=>"011000100",
  46409=>"101101101",
  46410=>"011110111",
  46411=>"000000000",
  46412=>"001001011",
  46413=>"100111001",
  46414=>"001001010",
  46415=>"001100000",
  46416=>"100111110",
  46417=>"111101000",
  46418=>"110000011",
  46419=>"011111011",
  46420=>"000001011",
  46421=>"111010110",
  46422=>"001001100",
  46423=>"010101111",
  46424=>"110110111",
  46425=>"001011010",
  46426=>"101010001",
  46427=>"001110011",
  46428=>"001010011",
  46429=>"111011001",
  46430=>"100100000",
  46431=>"000010001",
  46432=>"100000100",
  46433=>"110001000",
  46434=>"111100110",
  46435=>"100000110",
  46436=>"001001100",
  46437=>"111100010",
  46438=>"010100111",
  46439=>"010111101",
  46440=>"101111011",
  46441=>"000000100",
  46442=>"100101110",
  46443=>"011000010",
  46444=>"100010111",
  46445=>"100100010",
  46446=>"000001000",
  46447=>"010100000",
  46448=>"111001100",
  46449=>"101001101",
  46450=>"101101111",
  46451=>"001011101",
  46452=>"000010001",
  46453=>"110100101",
  46454=>"010111010",
  46455=>"011011001",
  46456=>"100111100",
  46457=>"001100110",
  46458=>"000011101",
  46459=>"110110100",
  46460=>"101100010",
  46461=>"110111011",
  46462=>"110110011",
  46463=>"000110111",
  46464=>"000111110",
  46465=>"011010110",
  46466=>"010111010",
  46467=>"100010111",
  46468=>"000010100",
  46469=>"011011110",
  46470=>"000111100",
  46471=>"111101010",
  46472=>"000010100",
  46473=>"111000011",
  46474=>"110011000",
  46475=>"101100001",
  46476=>"001111011",
  46477=>"101101110",
  46478=>"111100001",
  46479=>"111000011",
  46480=>"001000100",
  46481=>"010000100",
  46482=>"010000000",
  46483=>"001010010",
  46484=>"010100001",
  46485=>"000100111",
  46486=>"001010001",
  46487=>"101110001",
  46488=>"111100110",
  46489=>"100010101",
  46490=>"010100000",
  46491=>"011100100",
  46492=>"010010010",
  46493=>"011011110",
  46494=>"010001101",
  46495=>"000000011",
  46496=>"111000100",
  46497=>"010011100",
  46498=>"100101101",
  46499=>"110110111",
  46500=>"011100100",
  46501=>"100100011",
  46502=>"100001000",
  46503=>"000111111",
  46504=>"100011111",
  46505=>"110001111",
  46506=>"011000000",
  46507=>"110110010",
  46508=>"101100011",
  46509=>"100111110",
  46510=>"000100010",
  46511=>"010010001",
  46512=>"110011001",
  46513=>"011011010",
  46514=>"111101110",
  46515=>"010011111",
  46516=>"101110010",
  46517=>"010010000",
  46518=>"100010001",
  46519=>"011100110",
  46520=>"110000011",
  46521=>"000100110",
  46522=>"100100000",
  46523=>"010100000",
  46524=>"111000010",
  46525=>"110111000",
  46526=>"000111110",
  46527=>"100001000",
  46528=>"000001100",
  46529=>"000011010",
  46530=>"010110111",
  46531=>"100011010",
  46532=>"100001000",
  46533=>"010101100",
  46534=>"001100001",
  46535=>"011011100",
  46536=>"110010001",
  46537=>"010111111",
  46538=>"110110001",
  46539=>"010101101",
  46540=>"010001000",
  46541=>"110010010",
  46542=>"100010000",
  46543=>"001110001",
  46544=>"011111011",
  46545=>"010001110",
  46546=>"101101000",
  46547=>"110000011",
  46548=>"100010111",
  46549=>"000001100",
  46550=>"011110000",
  46551=>"100010101",
  46552=>"111010111",
  46553=>"001111000",
  46554=>"110100010",
  46555=>"100000011",
  46556=>"111011100",
  46557=>"111110111",
  46558=>"100011110",
  46559=>"010001100",
  46560=>"111111101",
  46561=>"001101001",
  46562=>"111000011",
  46563=>"100001101",
  46564=>"111111010",
  46565=>"010001110",
  46566=>"001100000",
  46567=>"101010000",
  46568=>"010011100",
  46569=>"000000100",
  46570=>"011101011",
  46571=>"111011001",
  46572=>"111011000",
  46573=>"000101010",
  46574=>"001011000",
  46575=>"011100110",
  46576=>"110101011",
  46577=>"101001111",
  46578=>"011010101",
  46579=>"000110010",
  46580=>"110110010",
  46581=>"000001001",
  46582=>"110000110",
  46583=>"110011000",
  46584=>"010101001",
  46585=>"010101110",
  46586=>"011111110",
  46587=>"101000100",
  46588=>"111100110",
  46589=>"010111010",
  46590=>"011101001",
  46591=>"010110110",
  46592=>"111001010",
  46593=>"100111101",
  46594=>"101011011",
  46595=>"101110001",
  46596=>"001001010",
  46597=>"010001111",
  46598=>"000111110",
  46599=>"100000111",
  46600=>"101100001",
  46601=>"011100010",
  46602=>"001101010",
  46603=>"111010111",
  46604=>"001000100",
  46605=>"100111010",
  46606=>"010000011",
  46607=>"010110001",
  46608=>"011111110",
  46609=>"001111111",
  46610=>"111101111",
  46611=>"011100010",
  46612=>"011001010",
  46613=>"110101001",
  46614=>"011101000",
  46615=>"111011111",
  46616=>"111000001",
  46617=>"001001110",
  46618=>"110001001",
  46619=>"000110111",
  46620=>"000100100",
  46621=>"110101011",
  46622=>"011011011",
  46623=>"011011011",
  46624=>"011100101",
  46625=>"100010011",
  46626=>"001110110",
  46627=>"001100001",
  46628=>"001111010",
  46629=>"001001101",
  46630=>"010111011",
  46631=>"111100101",
  46632=>"000011111",
  46633=>"110000110",
  46634=>"001000011",
  46635=>"000101010",
  46636=>"010000000",
  46637=>"110100000",
  46638=>"110100001",
  46639=>"000100001",
  46640=>"011101111",
  46641=>"111000000",
  46642=>"110101010",
  46643=>"001111001",
  46644=>"011110001",
  46645=>"110000100",
  46646=>"000100101",
  46647=>"010010011",
  46648=>"110010111",
  46649=>"110010011",
  46650=>"001010001",
  46651=>"000000010",
  46652=>"101100100",
  46653=>"000111011",
  46654=>"111000100",
  46655=>"001000011",
  46656=>"110110100",
  46657=>"001101001",
  46658=>"110110000",
  46659=>"000010001",
  46660=>"101110111",
  46661=>"110100101",
  46662=>"000100100",
  46663=>"011110010",
  46664=>"010001110",
  46665=>"110111111",
  46666=>"000000001",
  46667=>"000000100",
  46668=>"110101111",
  46669=>"000000011",
  46670=>"111100011",
  46671=>"011100010",
  46672=>"101100110",
  46673=>"000110110",
  46674=>"010100110",
  46675=>"110010100",
  46676=>"101001001",
  46677=>"101001101",
  46678=>"101111011",
  46679=>"111100011",
  46680=>"001011110",
  46681=>"011101011",
  46682=>"100010001",
  46683=>"010100100",
  46684=>"100001111",
  46685=>"011011111",
  46686=>"111011011",
  46687=>"110000000",
  46688=>"000000101",
  46689=>"110000011",
  46690=>"111010111",
  46691=>"100010110",
  46692=>"010110001",
  46693=>"001011101",
  46694=>"011011101",
  46695=>"101101010",
  46696=>"100111111",
  46697=>"101011110",
  46698=>"011001110",
  46699=>"010000001",
  46700=>"110001100",
  46701=>"000111101",
  46702=>"110111100",
  46703=>"010100000",
  46704=>"100010010",
  46705=>"000100000",
  46706=>"100001001",
  46707=>"000101101",
  46708=>"000011011",
  46709=>"111110111",
  46710=>"101001101",
  46711=>"110101101",
  46712=>"010000000",
  46713=>"011100011",
  46714=>"001110011",
  46715=>"101011110",
  46716=>"000011000",
  46717=>"001100001",
  46718=>"110101010",
  46719=>"000011010",
  46720=>"010001110",
  46721=>"001100000",
  46722=>"110001101",
  46723=>"001010100",
  46724=>"000100100",
  46725=>"101001001",
  46726=>"111101111",
  46727=>"111111110",
  46728=>"100110100",
  46729=>"010100111",
  46730=>"000100000",
  46731=>"011000001",
  46732=>"011100010",
  46733=>"111011000",
  46734=>"111010011",
  46735=>"000000010",
  46736=>"000110011",
  46737=>"001010100",
  46738=>"000000011",
  46739=>"111001000",
  46740=>"000000110",
  46741=>"010101100",
  46742=>"010110010",
  46743=>"001111111",
  46744=>"010001111",
  46745=>"110100101",
  46746=>"111001110",
  46747=>"000000000",
  46748=>"110000110",
  46749=>"111010000",
  46750=>"010111011",
  46751=>"010100010",
  46752=>"010101010",
  46753=>"100000001",
  46754=>"000011110",
  46755=>"100011000",
  46756=>"100010101",
  46757=>"110111001",
  46758=>"010010110",
  46759=>"101111101",
  46760=>"011010011",
  46761=>"010101101",
  46762=>"011101101",
  46763=>"100001001",
  46764=>"110100101",
  46765=>"001001000",
  46766=>"111101111",
  46767=>"100010100",
  46768=>"110000011",
  46769=>"010110010",
  46770=>"110100010",
  46771=>"001000111",
  46772=>"001011011",
  46773=>"011110011",
  46774=>"110011100",
  46775=>"001001100",
  46776=>"101111011",
  46777=>"000100100",
  46778=>"111111001",
  46779=>"101010000",
  46780=>"011101011",
  46781=>"010001000",
  46782=>"011111110",
  46783=>"000000010",
  46784=>"100110111",
  46785=>"001010111",
  46786=>"101111100",
  46787=>"110010101",
  46788=>"100011011",
  46789=>"010011000",
  46790=>"000001011",
  46791=>"100011100",
  46792=>"000100010",
  46793=>"000101000",
  46794=>"100101000",
  46795=>"110001000",
  46796=>"000100000",
  46797=>"100101001",
  46798=>"000010101",
  46799=>"011101100",
  46800=>"101101000",
  46801=>"001011001",
  46802=>"101011011",
  46803=>"101101011",
  46804=>"001100000",
  46805=>"110000010",
  46806=>"001011110",
  46807=>"100110101",
  46808=>"000001110",
  46809=>"110111010",
  46810=>"011000001",
  46811=>"111100010",
  46812=>"101111100",
  46813=>"001001001",
  46814=>"000000100",
  46815=>"101000101",
  46816=>"001010011",
  46817=>"000011011",
  46818=>"010111111",
  46819=>"111011000",
  46820=>"100011001",
  46821=>"111100110",
  46822=>"000010110",
  46823=>"000110110",
  46824=>"010111001",
  46825=>"111111111",
  46826=>"000110010",
  46827=>"111101010",
  46828=>"111100000",
  46829=>"101110011",
  46830=>"111000001",
  46831=>"100100000",
  46832=>"100101110",
  46833=>"101100011",
  46834=>"100101010",
  46835=>"111101101",
  46836=>"111111100",
  46837=>"110110010",
  46838=>"111001000",
  46839=>"100000011",
  46840=>"100000001",
  46841=>"100101101",
  46842=>"110100010",
  46843=>"101010101",
  46844=>"110111011",
  46845=>"100101010",
  46846=>"000010000",
  46847=>"100001000",
  46848=>"100101111",
  46849=>"111000010",
  46850=>"001010101",
  46851=>"011111011",
  46852=>"101101101",
  46853=>"100010000",
  46854=>"111101001",
  46855=>"000000111",
  46856=>"001000110",
  46857=>"010110010",
  46858=>"001011111",
  46859=>"111000011",
  46860=>"100110000",
  46861=>"100010011",
  46862=>"110110110",
  46863=>"101110011",
  46864=>"101011000",
  46865=>"000001101",
  46866=>"011011011",
  46867=>"010010111",
  46868=>"000010111",
  46869=>"101000111",
  46870=>"000010000",
  46871=>"110110100",
  46872=>"010000010",
  46873=>"111101001",
  46874=>"001111111",
  46875=>"001001000",
  46876=>"011001101",
  46877=>"100010000",
  46878=>"011010100",
  46879=>"011101000",
  46880=>"111001111",
  46881=>"100000111",
  46882=>"111010000",
  46883=>"000100011",
  46884=>"001100101",
  46885=>"111110001",
  46886=>"010110100",
  46887=>"010010010",
  46888=>"000110011",
  46889=>"111101110",
  46890=>"110101100",
  46891=>"101101001",
  46892=>"010100111",
  46893=>"000100110",
  46894=>"101111110",
  46895=>"011010110",
  46896=>"011100010",
  46897=>"111100000",
  46898=>"101001100",
  46899=>"101000000",
  46900=>"010101111",
  46901=>"101111100",
  46902=>"001000000",
  46903=>"101111100",
  46904=>"110000000",
  46905=>"001000010",
  46906=>"100010000",
  46907=>"101010111",
  46908=>"000100011",
  46909=>"111000010",
  46910=>"101111001",
  46911=>"000100111",
  46912=>"101110010",
  46913=>"100011000",
  46914=>"001111010",
  46915=>"100100000",
  46916=>"100010100",
  46917=>"011101111",
  46918=>"101111111",
  46919=>"011011001",
  46920=>"101111111",
  46921=>"001101111",
  46922=>"010010101",
  46923=>"111100111",
  46924=>"001000100",
  46925=>"100011011",
  46926=>"011001001",
  46927=>"011101100",
  46928=>"101010001",
  46929=>"111010001",
  46930=>"110010010",
  46931=>"101001101",
  46932=>"111100000",
  46933=>"110001111",
  46934=>"010111111",
  46935=>"011111101",
  46936=>"000111111",
  46937=>"111010000",
  46938=>"010011110",
  46939=>"101111101",
  46940=>"000001100",
  46941=>"111000100",
  46942=>"111110000",
  46943=>"110001001",
  46944=>"000110100",
  46945=>"110000011",
  46946=>"011000111",
  46947=>"000110101",
  46948=>"000001000",
  46949=>"001001110",
  46950=>"100011110",
  46951=>"100111101",
  46952=>"100000001",
  46953=>"001110100",
  46954=>"111101111",
  46955=>"001011000",
  46956=>"111111001",
  46957=>"001010001",
  46958=>"011111010",
  46959=>"100111100",
  46960=>"011101111",
  46961=>"001101001",
  46962=>"110110000",
  46963=>"010100010",
  46964=>"001000000",
  46965=>"011010110",
  46966=>"011011101",
  46967=>"111110111",
  46968=>"000110010",
  46969=>"011111101",
  46970=>"010001100",
  46971=>"000101010",
  46972=>"100101000",
  46973=>"101110100",
  46974=>"110001110",
  46975=>"000000001",
  46976=>"110110010",
  46977=>"110100000",
  46978=>"010011111",
  46979=>"001110000",
  46980=>"011100101",
  46981=>"101101100",
  46982=>"000100000",
  46983=>"110100010",
  46984=>"101011010",
  46985=>"101110111",
  46986=>"100011111",
  46987=>"000101101",
  46988=>"110111100",
  46989=>"111110111",
  46990=>"011011101",
  46991=>"110101111",
  46992=>"111101100",
  46993=>"110101011",
  46994=>"011001110",
  46995=>"111101011",
  46996=>"111011010",
  46997=>"110011000",
  46998=>"010001010",
  46999=>"101100100",
  47000=>"001100110",
  47001=>"001110111",
  47002=>"011011101",
  47003=>"010011110",
  47004=>"001110111",
  47005=>"000110011",
  47006=>"011110010",
  47007=>"111100101",
  47008=>"010110100",
  47009=>"011101000",
  47010=>"100111110",
  47011=>"100000101",
  47012=>"001001011",
  47013=>"101110111",
  47014=>"111000011",
  47015=>"000001000",
  47016=>"111010010",
  47017=>"110000101",
  47018=>"111100011",
  47019=>"001011001",
  47020=>"001110110",
  47021=>"010011100",
  47022=>"110101100",
  47023=>"011101111",
  47024=>"000010011",
  47025=>"100110000",
  47026=>"010100010",
  47027=>"111000101",
  47028=>"010111000",
  47029=>"001010111",
  47030=>"011010001",
  47031=>"111000111",
  47032=>"001100010",
  47033=>"011010100",
  47034=>"100100110",
  47035=>"000100111",
  47036=>"011011011",
  47037=>"101100111",
  47038=>"010001111",
  47039=>"101111100",
  47040=>"001010010",
  47041=>"010111000",
  47042=>"111101000",
  47043=>"110100010",
  47044=>"000111001",
  47045=>"011000111",
  47046=>"000110100",
  47047=>"110111111",
  47048=>"111011011",
  47049=>"010011010",
  47050=>"000100110",
  47051=>"111010011",
  47052=>"111000110",
  47053=>"011110010",
  47054=>"010100011",
  47055=>"111111010",
  47056=>"110110110",
  47057=>"111000011",
  47058=>"001010101",
  47059=>"101100010",
  47060=>"101110111",
  47061=>"100000111",
  47062=>"010001001",
  47063=>"110000010",
  47064=>"110000110",
  47065=>"101111100",
  47066=>"100101100",
  47067=>"100000000",
  47068=>"110101101",
  47069=>"101111100",
  47070=>"000111011",
  47071=>"000111110",
  47072=>"111101110",
  47073=>"000000100",
  47074=>"001000010",
  47075=>"011001101",
  47076=>"010001000",
  47077=>"001010010",
  47078=>"010010000",
  47079=>"110101001",
  47080=>"000100110",
  47081=>"011101001",
  47082=>"010011100",
  47083=>"011101001",
  47084=>"110101111",
  47085=>"110011001",
  47086=>"000011000",
  47087=>"110101101",
  47088=>"111100010",
  47089=>"001111101",
  47090=>"100111111",
  47091=>"101001010",
  47092=>"110010010",
  47093=>"000100110",
  47094=>"001010000",
  47095=>"100000010",
  47096=>"111110110",
  47097=>"011100000",
  47098=>"100100000",
  47099=>"010001111",
  47100=>"110001111",
  47101=>"010001100",
  47102=>"100000110",
  47103=>"000100001",
  47104=>"100000100",
  47105=>"101111000",
  47106=>"011110010",
  47107=>"011110000",
  47108=>"001111001",
  47109=>"100011000",
  47110=>"011111100",
  47111=>"101011101",
  47112=>"010011010",
  47113=>"111101111",
  47114=>"111000101",
  47115=>"110011010",
  47116=>"101101001",
  47117=>"100000100",
  47118=>"011001010",
  47119=>"111001101",
  47120=>"110111111",
  47121=>"110010001",
  47122=>"100000101",
  47123=>"100001110",
  47124=>"000100010",
  47125=>"010010011",
  47126=>"110101111",
  47127=>"000100001",
  47128=>"000010111",
  47129=>"101111111",
  47130=>"100010001",
  47131=>"111110111",
  47132=>"111100001",
  47133=>"000010011",
  47134=>"100101111",
  47135=>"111110101",
  47136=>"010110001",
  47137=>"101100010",
  47138=>"100001000",
  47139=>"000001001",
  47140=>"101100111",
  47141=>"111010001",
  47142=>"110101011",
  47143=>"000011010",
  47144=>"001111011",
  47145=>"100110110",
  47146=>"000110111",
  47147=>"010000000",
  47148=>"000100010",
  47149=>"111100001",
  47150=>"011001000",
  47151=>"100111000",
  47152=>"111111001",
  47153=>"000010100",
  47154=>"011000111",
  47155=>"000000011",
  47156=>"010100001",
  47157=>"010000000",
  47158=>"101111100",
  47159=>"110010100",
  47160=>"111111101",
  47161=>"000010101",
  47162=>"111000001",
  47163=>"000011001",
  47164=>"100010111",
  47165=>"100001000",
  47166=>"111001000",
  47167=>"011101010",
  47168=>"001101110",
  47169=>"001000011",
  47170=>"101000100",
  47171=>"010000010",
  47172=>"001011000",
  47173=>"101101100",
  47174=>"101110101",
  47175=>"101011001",
  47176=>"111110001",
  47177=>"111111001",
  47178=>"110100001",
  47179=>"100001010",
  47180=>"101100011",
  47181=>"011111111",
  47182=>"010000000",
  47183=>"000100110",
  47184=>"011001010",
  47185=>"011000100",
  47186=>"010101110",
  47187=>"111111111",
  47188=>"011100111",
  47189=>"110101100",
  47190=>"111101000",
  47191=>"011101000",
  47192=>"010101111",
  47193=>"101010001",
  47194=>"110010000",
  47195=>"110000010",
  47196=>"011010011",
  47197=>"101100101",
  47198=>"100000100",
  47199=>"110010101",
  47200=>"111011000",
  47201=>"100101011",
  47202=>"000111101",
  47203=>"000001110",
  47204=>"001001111",
  47205=>"010000110",
  47206=>"100110110",
  47207=>"111010100",
  47208=>"100111100",
  47209=>"001011000",
  47210=>"110101001",
  47211=>"100011010",
  47212=>"101001011",
  47213=>"111000001",
  47214=>"101000001",
  47215=>"101001011",
  47216=>"100010101",
  47217=>"000011001",
  47218=>"001101001",
  47219=>"100111010",
  47220=>"111100000",
  47221=>"100101001",
  47222=>"100101100",
  47223=>"111010000",
  47224=>"111011111",
  47225=>"110011101",
  47226=>"110110010",
  47227=>"000111111",
  47228=>"000010001",
  47229=>"101110000",
  47230=>"000101100",
  47231=>"110010010",
  47232=>"001011011",
  47233=>"111010111",
  47234=>"111000001",
  47235=>"111011101",
  47236=>"001101001",
  47237=>"100011010",
  47238=>"111110010",
  47239=>"000000100",
  47240=>"011011000",
  47241=>"100110001",
  47242=>"010010111",
  47243=>"111000100",
  47244=>"000111000",
  47245=>"001110100",
  47246=>"100001010",
  47247=>"000111110",
  47248=>"000111000",
  47249=>"001110111",
  47250=>"111100101",
  47251=>"000101001",
  47252=>"111101110",
  47253=>"111001010",
  47254=>"000111011",
  47255=>"110001111",
  47256=>"111110100",
  47257=>"000111111",
  47258=>"010010011",
  47259=>"011110000",
  47260=>"101110010",
  47261=>"011111101",
  47262=>"000110110",
  47263=>"001110011",
  47264=>"100101101",
  47265=>"110010110",
  47266=>"101100101",
  47267=>"001111010",
  47268=>"000111110",
  47269=>"000100101",
  47270=>"100110110",
  47271=>"101100101",
  47272=>"001110111",
  47273=>"010010001",
  47274=>"110000000",
  47275=>"010001111",
  47276=>"110111100",
  47277=>"100001110",
  47278=>"010001100",
  47279=>"111010110",
  47280=>"100111100",
  47281=>"011011001",
  47282=>"001011001",
  47283=>"100111010",
  47284=>"000000000",
  47285=>"110001010",
  47286=>"011001101",
  47287=>"000000110",
  47288=>"011010100",
  47289=>"000101100",
  47290=>"110011000",
  47291=>"001101010",
  47292=>"110001001",
  47293=>"000000010",
  47294=>"011010000",
  47295=>"001111010",
  47296=>"100000100",
  47297=>"011000100",
  47298=>"001111010",
  47299=>"010010111",
  47300=>"011011111",
  47301=>"101001101",
  47302=>"000000010",
  47303=>"101111111",
  47304=>"011011010",
  47305=>"010000010",
  47306=>"100100100",
  47307=>"000111010",
  47308=>"000010001",
  47309=>"100100110",
  47310=>"000010100",
  47311=>"110111010",
  47312=>"011110011",
  47313=>"010101111",
  47314=>"001100000",
  47315=>"101001101",
  47316=>"000111100",
  47317=>"100001101",
  47318=>"001010000",
  47319=>"010110000",
  47320=>"001011010",
  47321=>"110100000",
  47322=>"000110111",
  47323=>"011011111",
  47324=>"111010000",
  47325=>"011101101",
  47326=>"001100010",
  47327=>"011000010",
  47328=>"100000001",
  47329=>"110010101",
  47330=>"101110010",
  47331=>"111010110",
  47332=>"101110000",
  47333=>"000000110",
  47334=>"101101001",
  47335=>"010001111",
  47336=>"011101010",
  47337=>"000010000",
  47338=>"001100011",
  47339=>"101000001",
  47340=>"100010100",
  47341=>"111011110",
  47342=>"111100011",
  47343=>"010100111",
  47344=>"010000010",
  47345=>"001000010",
  47346=>"001101101",
  47347=>"000000010",
  47348=>"111100000",
  47349=>"000100100",
  47350=>"001101010",
  47351=>"000100001",
  47352=>"101010001",
  47353=>"101001000",
  47354=>"111011010",
  47355=>"101001101",
  47356=>"010100111",
  47357=>"111111110",
  47358=>"110111011",
  47359=>"110110011",
  47360=>"001100111",
  47361=>"011101101",
  47362=>"010001101",
  47363=>"100001101",
  47364=>"001011101",
  47365=>"100011110",
  47366=>"110000101",
  47367=>"001000011",
  47368=>"110110101",
  47369=>"101010110",
  47370=>"101011000",
  47371=>"101011000",
  47372=>"100110100",
  47373=>"111010100",
  47374=>"010000001",
  47375=>"010010111",
  47376=>"100010001",
  47377=>"010001110",
  47378=>"111111100",
  47379=>"011011010",
  47380=>"000000110",
  47381=>"001111001",
  47382=>"001100010",
  47383=>"101011110",
  47384=>"111010101",
  47385=>"100001010",
  47386=>"111111100",
  47387=>"000110110",
  47388=>"110101111",
  47389=>"111001001",
  47390=>"010100001",
  47391=>"000010011",
  47392=>"110110010",
  47393=>"111000011",
  47394=>"111001111",
  47395=>"110101001",
  47396=>"000110011",
  47397=>"101010011",
  47398=>"010110000",
  47399=>"001001101",
  47400=>"011101001",
  47401=>"101010101",
  47402=>"111010001",
  47403=>"111110000",
  47404=>"010111110",
  47405=>"100000000",
  47406=>"110001011",
  47407=>"100000111",
  47408=>"000011101",
  47409=>"010001111",
  47410=>"111000111",
  47411=>"111111110",
  47412=>"010000000",
  47413=>"001011101",
  47414=>"001100010",
  47415=>"110001101",
  47416=>"100010110",
  47417=>"011011110",
  47418=>"111100110",
  47419=>"010000010",
  47420=>"110100100",
  47421=>"101101111",
  47422=>"000100011",
  47423=>"111100011",
  47424=>"111110110",
  47425=>"100101011",
  47426=>"010001000",
  47427=>"000001111",
  47428=>"000000001",
  47429=>"011111101",
  47430=>"100001111",
  47431=>"111110010",
  47432=>"111000011",
  47433=>"010010011",
  47434=>"001110011",
  47435=>"010000110",
  47436=>"110100101",
  47437=>"111110011",
  47438=>"011001111",
  47439=>"110111100",
  47440=>"111010010",
  47441=>"110101000",
  47442=>"001001010",
  47443=>"100110001",
  47444=>"111101011",
  47445=>"011000110",
  47446=>"110001111",
  47447=>"001100000",
  47448=>"010111100",
  47449=>"100011001",
  47450=>"001110100",
  47451=>"001110101",
  47452=>"101011001",
  47453=>"011010110",
  47454=>"000010010",
  47455=>"111000000",
  47456=>"111110111",
  47457=>"010011001",
  47458=>"001010111",
  47459=>"111111010",
  47460=>"101000111",
  47461=>"011100011",
  47462=>"110111110",
  47463=>"110100011",
  47464=>"001111001",
  47465=>"100011111",
  47466=>"010110111",
  47467=>"010000110",
  47468=>"000011100",
  47469=>"110011110",
  47470=>"001111110",
  47471=>"011111111",
  47472=>"001100100",
  47473=>"001100011",
  47474=>"011100001",
  47475=>"001010111",
  47476=>"000011110",
  47477=>"000001111",
  47478=>"111111110",
  47479=>"010011101",
  47480=>"000000000",
  47481=>"010011111",
  47482=>"001001001",
  47483=>"111011101",
  47484=>"010111001",
  47485=>"001110110",
  47486=>"111010100",
  47487=>"000000010",
  47488=>"111011111",
  47489=>"011101000",
  47490=>"101110110",
  47491=>"000010110",
  47492=>"011010001",
  47493=>"010110001",
  47494=>"101101001",
  47495=>"000010111",
  47496=>"000000011",
  47497=>"101110000",
  47498=>"111011011",
  47499=>"010001110",
  47500=>"001100011",
  47501=>"111011010",
  47502=>"000111100",
  47503=>"001001011",
  47504=>"110000100",
  47505=>"110011111",
  47506=>"010001011",
  47507=>"011010011",
  47508=>"011100011",
  47509=>"101101010",
  47510=>"100011000",
  47511=>"101000001",
  47512=>"011110011",
  47513=>"101100000",
  47514=>"001011011",
  47515=>"110100010",
  47516=>"100110000",
  47517=>"110000000",
  47518=>"111011100",
  47519=>"110010000",
  47520=>"100100100",
  47521=>"101000000",
  47522=>"010010111",
  47523=>"001000001",
  47524=>"100100111",
  47525=>"010011101",
  47526=>"011110110",
  47527=>"001000100",
  47528=>"001011001",
  47529=>"000100010",
  47530=>"001000000",
  47531=>"001010001",
  47532=>"111111010",
  47533=>"100001010",
  47534=>"111001100",
  47535=>"001101100",
  47536=>"110100111",
  47537=>"010100110",
  47538=>"000110000",
  47539=>"101000101",
  47540=>"111011100",
  47541=>"010111100",
  47542=>"111010100",
  47543=>"100100101",
  47544=>"000011101",
  47545=>"110000110",
  47546=>"110100001",
  47547=>"100001110",
  47548=>"110010101",
  47549=>"010001000",
  47550=>"111101000",
  47551=>"110010101",
  47552=>"101000000",
  47553=>"101000100",
  47554=>"100100001",
  47555=>"011001001",
  47556=>"000101100",
  47557=>"001101111",
  47558=>"100001000",
  47559=>"100001111",
  47560=>"100011111",
  47561=>"111111101",
  47562=>"100010110",
  47563=>"101100110",
  47564=>"001000000",
  47565=>"110110110",
  47566=>"000100010",
  47567=>"111101111",
  47568=>"001101110",
  47569=>"110101111",
  47570=>"000101110",
  47571=>"010100110",
  47572=>"100001010",
  47573=>"101000000",
  47574=>"010110110",
  47575=>"111000000",
  47576=>"111000101",
  47577=>"010001101",
  47578=>"110110111",
  47579=>"010111010",
  47580=>"111101101",
  47581=>"011001111",
  47582=>"100000110",
  47583=>"101100010",
  47584=>"001011110",
  47585=>"111000111",
  47586=>"000001110",
  47587=>"001000101",
  47588=>"110101011",
  47589=>"001100010",
  47590=>"000101011",
  47591=>"111101010",
  47592=>"101111001",
  47593=>"101010000",
  47594=>"100100100",
  47595=>"001001101",
  47596=>"111110001",
  47597=>"010000110",
  47598=>"100011011",
  47599=>"110001011",
  47600=>"000110111",
  47601=>"000101011",
  47602=>"010001011",
  47603=>"110100111",
  47604=>"000100010",
  47605=>"001000100",
  47606=>"111100010",
  47607=>"010011011",
  47608=>"101000010",
  47609=>"101110000",
  47610=>"010001000",
  47611=>"110111011",
  47612=>"110100100",
  47613=>"111010000",
  47614=>"101110100",
  47615=>"011000001",
  47616=>"110111011",
  47617=>"111010100",
  47618=>"010010011",
  47619=>"111101000",
  47620=>"111101111",
  47621=>"001111001",
  47622=>"111011010",
  47623=>"110110100",
  47624=>"110000010",
  47625=>"001011101",
  47626=>"100011110",
  47627=>"011010000",
  47628=>"010100111",
  47629=>"011100011",
  47630=>"100101000",
  47631=>"001001010",
  47632=>"001011001",
  47633=>"011011100",
  47634=>"111010111",
  47635=>"100101100",
  47636=>"010011111",
  47637=>"111111010",
  47638=>"100111110",
  47639=>"101100000",
  47640=>"100100111",
  47641=>"011111000",
  47642=>"101010110",
  47643=>"011110000",
  47644=>"011011000",
  47645=>"110010100",
  47646=>"011001000",
  47647=>"000100110",
  47648=>"010010101",
  47649=>"101101010",
  47650=>"011000110",
  47651=>"011101111",
  47652=>"101111110",
  47653=>"111110001",
  47654=>"101100101",
  47655=>"110011000",
  47656=>"010000100",
  47657=>"011011100",
  47658=>"000111001",
  47659=>"000000010",
  47660=>"000110011",
  47661=>"011010011",
  47662=>"010100111",
  47663=>"010001100",
  47664=>"100111111",
  47665=>"110100110",
  47666=>"010100000",
  47667=>"011111011",
  47668=>"001111100",
  47669=>"101001000",
  47670=>"001011111",
  47671=>"110110001",
  47672=>"000100010",
  47673=>"101110110",
  47674=>"101011000",
  47675=>"101011101",
  47676=>"010010110",
  47677=>"010011101",
  47678=>"110000101",
  47679=>"010001111",
  47680=>"011011111",
  47681=>"111111011",
  47682=>"010010001",
  47683=>"001011010",
  47684=>"110000111",
  47685=>"110001110",
  47686=>"101110100",
  47687=>"000011110",
  47688=>"011101110",
  47689=>"111111001",
  47690=>"111001001",
  47691=>"111011111",
  47692=>"111101001",
  47693=>"000110011",
  47694=>"011010111",
  47695=>"011010101",
  47696=>"111011111",
  47697=>"000110100",
  47698=>"110101101",
  47699=>"110011111",
  47700=>"111010111",
  47701=>"001001101",
  47702=>"001101001",
  47703=>"000010101",
  47704=>"111100101",
  47705=>"101000010",
  47706=>"011100010",
  47707=>"000000000",
  47708=>"001011100",
  47709=>"011111110",
  47710=>"101110101",
  47711=>"100000110",
  47712=>"010100110",
  47713=>"001000000",
  47714=>"110010110",
  47715=>"111001001",
  47716=>"010001110",
  47717=>"101110001",
  47718=>"111111111",
  47719=>"001011100",
  47720=>"010010110",
  47721=>"010101100",
  47722=>"010001011",
  47723=>"111111001",
  47724=>"100000001",
  47725=>"011101000",
  47726=>"111000111",
  47727=>"101001000",
  47728=>"100010100",
  47729=>"101100101",
  47730=>"111101101",
  47731=>"111100001",
  47732=>"000111111",
  47733=>"011001000",
  47734=>"101111111",
  47735=>"111110100",
  47736=>"111000000",
  47737=>"001001000",
  47738=>"011000000",
  47739=>"010000011",
  47740=>"110111001",
  47741=>"110110101",
  47742=>"111111111",
  47743=>"011100100",
  47744=>"100011111",
  47745=>"101010011",
  47746=>"111101011",
  47747=>"110100001",
  47748=>"110100000",
  47749=>"000001101",
  47750=>"001000011",
  47751=>"110010010",
  47752=>"111010011",
  47753=>"110111000",
  47754=>"011101111",
  47755=>"110011010",
  47756=>"111010011",
  47757=>"001000101",
  47758=>"010011001",
  47759=>"111111001",
  47760=>"000101100",
  47761=>"000111101",
  47762=>"011000101",
  47763=>"011100100",
  47764=>"100101010",
  47765=>"001110000",
  47766=>"101100100",
  47767=>"100111011",
  47768=>"010011001",
  47769=>"011100100",
  47770=>"001011110",
  47771=>"001000110",
  47772=>"110000101",
  47773=>"000100010",
  47774=>"101110100",
  47775=>"111101011",
  47776=>"000010111",
  47777=>"100101000",
  47778=>"101111111",
  47779=>"001010001",
  47780=>"110011110",
  47781=>"101111001",
  47782=>"001010101",
  47783=>"110110111",
  47784=>"000110110",
  47785=>"001000100",
  47786=>"100101010",
  47787=>"110011000",
  47788=>"101110010",
  47789=>"111011100",
  47790=>"011011111",
  47791=>"000010001",
  47792=>"001100101",
  47793=>"111101001",
  47794=>"001100110",
  47795=>"001010110",
  47796=>"011001001",
  47797=>"000001101",
  47798=>"001010111",
  47799=>"011000001",
  47800=>"101111101",
  47801=>"111100000",
  47802=>"001001011",
  47803=>"101010100",
  47804=>"100010000",
  47805=>"111101110",
  47806=>"111000111",
  47807=>"100011100",
  47808=>"000001010",
  47809=>"001110001",
  47810=>"110101111",
  47811=>"001010110",
  47812=>"111111001",
  47813=>"110011000",
  47814=>"110000101",
  47815=>"001110011",
  47816=>"010111001",
  47817=>"111001011",
  47818=>"110100011",
  47819=>"000000000",
  47820=>"110001110",
  47821=>"110000010",
  47822=>"110100100",
  47823=>"001111110",
  47824=>"010100010",
  47825=>"000000010",
  47826=>"000100100",
  47827=>"000011010",
  47828=>"110001001",
  47829=>"011000110",
  47830=>"011001111",
  47831=>"100100000",
  47832=>"101101010",
  47833=>"010010011",
  47834=>"011101001",
  47835=>"001100011",
  47836=>"001001100",
  47837=>"101001000",
  47838=>"010100111",
  47839=>"011111110",
  47840=>"000100111",
  47841=>"000101001",
  47842=>"111110110",
  47843=>"100110100",
  47844=>"010111101",
  47845=>"101011001",
  47846=>"000111111",
  47847=>"101011000",
  47848=>"110000010",
  47849=>"101101010",
  47850=>"001100110",
  47851=>"110010000",
  47852=>"101001101",
  47853=>"000101100",
  47854=>"101011010",
  47855=>"111101111",
  47856=>"100111110",
  47857=>"000101100",
  47858=>"000011010",
  47859=>"000011101",
  47860=>"100110111",
  47861=>"011100010",
  47862=>"001111101",
  47863=>"010000000",
  47864=>"111011011",
  47865=>"010011001",
  47866=>"101111111",
  47867=>"001010100",
  47868=>"000110010",
  47869=>"011111111",
  47870=>"111011000",
  47871=>"011101100",
  47872=>"010011001",
  47873=>"110011111",
  47874=>"001111000",
  47875=>"111100101",
  47876=>"110101010",
  47877=>"100110101",
  47878=>"111101000",
  47879=>"001001110",
  47880=>"110011000",
  47881=>"011100001",
  47882=>"101011111",
  47883=>"111110011",
  47884=>"010010011",
  47885=>"001011111",
  47886=>"111100001",
  47887=>"111110101",
  47888=>"001101011",
  47889=>"011110100",
  47890=>"000001011",
  47891=>"111011000",
  47892=>"011101010",
  47893=>"000111010",
  47894=>"101110001",
  47895=>"111100100",
  47896=>"000001001",
  47897=>"001001111",
  47898=>"001010111",
  47899=>"101010001",
  47900=>"000001111",
  47901=>"110000001",
  47902=>"111110011",
  47903=>"000111010",
  47904=>"000100010",
  47905=>"111000010",
  47906=>"010010000",
  47907=>"111001111",
  47908=>"101100001",
  47909=>"000111010",
  47910=>"000101101",
  47911=>"010010101",
  47912=>"011100100",
  47913=>"101000101",
  47914=>"101111000",
  47915=>"110110011",
  47916=>"011010010",
  47917=>"011010011",
  47918=>"001001111",
  47919=>"010100010",
  47920=>"010011110",
  47921=>"101100111",
  47922=>"000110001",
  47923=>"110000000",
  47924=>"101001100",
  47925=>"011010110",
  47926=>"100010100",
  47927=>"001000001",
  47928=>"001011000",
  47929=>"100110100",
  47930=>"010000101",
  47931=>"100110111",
  47932=>"001111100",
  47933=>"001001110",
  47934=>"111100101",
  47935=>"111110000",
  47936=>"100111111",
  47937=>"001000011",
  47938=>"001101011",
  47939=>"000110011",
  47940=>"101100111",
  47941=>"100110110",
  47942=>"010010010",
  47943=>"111110111",
  47944=>"000101110",
  47945=>"010101101",
  47946=>"010100100",
  47947=>"100001001",
  47948=>"111001011",
  47949=>"001101010",
  47950=>"001001110",
  47951=>"110011011",
  47952=>"100001001",
  47953=>"000000010",
  47954=>"111101110",
  47955=>"001100000",
  47956=>"110101110",
  47957=>"010101011",
  47958=>"011100100",
  47959=>"111011101",
  47960=>"111110000",
  47961=>"110100111",
  47962=>"100101000",
  47963=>"000111010",
  47964=>"010010100",
  47965=>"010100010",
  47966=>"101000001",
  47967=>"101010000",
  47968=>"101010111",
  47969=>"110011010",
  47970=>"101000100",
  47971=>"011111010",
  47972=>"001010001",
  47973=>"001011111",
  47974=>"011001111",
  47975=>"100100100",
  47976=>"001001101",
  47977=>"000001110",
  47978=>"000000000",
  47979=>"010100001",
  47980=>"100011110",
  47981=>"000101101",
  47982=>"010110101",
  47983=>"011110011",
  47984=>"111000000",
  47985=>"001000010",
  47986=>"011101101",
  47987=>"100111011",
  47988=>"001101000",
  47989=>"000110000",
  47990=>"010111111",
  47991=>"000010111",
  47992=>"011000011",
  47993=>"000110100",
  47994=>"111101011",
  47995=>"110101101",
  47996=>"111110111",
  47997=>"001001110",
  47998=>"100011000",
  47999=>"000101011",
  48000=>"000011111",
  48001=>"111001001",
  48002=>"011010000",
  48003=>"000001010",
  48004=>"011000110",
  48005=>"111001000",
  48006=>"110100101",
  48007=>"000001000",
  48008=>"101001101",
  48009=>"010111100",
  48010=>"100000111",
  48011=>"111001111",
  48012=>"001010010",
  48013=>"011001001",
  48014=>"001011100",
  48015=>"101000111",
  48016=>"001001101",
  48017=>"100101011",
  48018=>"100111001",
  48019=>"101101000",
  48020=>"100101010",
  48021=>"011000110",
  48022=>"101111011",
  48023=>"010001001",
  48024=>"100100101",
  48025=>"000000100",
  48026=>"001010100",
  48027=>"001100100",
  48028=>"011110000",
  48029=>"000011001",
  48030=>"011110110",
  48031=>"100100000",
  48032=>"001111001",
  48033=>"001101101",
  48034=>"001000101",
  48035=>"001000101",
  48036=>"100110100",
  48037=>"111111000",
  48038=>"110000001",
  48039=>"000001110",
  48040=>"100011000",
  48041=>"011000010",
  48042=>"011000001",
  48043=>"000100101",
  48044=>"110000011",
  48045=>"100000000",
  48046=>"011110000",
  48047=>"000000000",
  48048=>"111010010",
  48049=>"111000010",
  48050=>"011000100",
  48051=>"101001000",
  48052=>"011111010",
  48053=>"101001111",
  48054=>"100001111",
  48055=>"011001011",
  48056=>"011001111",
  48057=>"100101100",
  48058=>"001001101",
  48059=>"101010011",
  48060=>"111111000",
  48061=>"111101111",
  48062=>"000101000",
  48063=>"001001111",
  48064=>"110110101",
  48065=>"001100100",
  48066=>"001101101",
  48067=>"100100000",
  48068=>"101001000",
  48069=>"111101111",
  48070=>"100001101",
  48071=>"010100001",
  48072=>"010010011",
  48073=>"100111111",
  48074=>"010001011",
  48075=>"011110001",
  48076=>"000101010",
  48077=>"100010000",
  48078=>"010011111",
  48079=>"110100010",
  48080=>"110111111",
  48081=>"111010010",
  48082=>"101101111",
  48083=>"010110110",
  48084=>"110011010",
  48085=>"100100101",
  48086=>"100000001",
  48087=>"001110001",
  48088=>"001000001",
  48089=>"100100011",
  48090=>"010100100",
  48091=>"000011100",
  48092=>"001010011",
  48093=>"010101101",
  48094=>"011011111",
  48095=>"010101011",
  48096=>"101001101",
  48097=>"001001011",
  48098=>"111110101",
  48099=>"110011101",
  48100=>"010100111",
  48101=>"111100111",
  48102=>"100001110",
  48103=>"000100000",
  48104=>"000001101",
  48105=>"101010001",
  48106=>"000000101",
  48107=>"100010000",
  48108=>"110110010",
  48109=>"111011001",
  48110=>"111011010",
  48111=>"011010001",
  48112=>"111100001",
  48113=>"100011110",
  48114=>"101100100",
  48115=>"011000011",
  48116=>"011110110",
  48117=>"010100000",
  48118=>"111101001",
  48119=>"000111100",
  48120=>"010001001",
  48121=>"111001111",
  48122=>"001011100",
  48123=>"001100100",
  48124=>"010101101",
  48125=>"100001000",
  48126=>"101011100",
  48127=>"111001011",
  48128=>"101110000",
  48129=>"101101100",
  48130=>"100110111",
  48131=>"001110101",
  48132=>"101000000",
  48133=>"011000001",
  48134=>"101000101",
  48135=>"100001000",
  48136=>"000000001",
  48137=>"000010000",
  48138=>"011011001",
  48139=>"010110011",
  48140=>"110000000",
  48141=>"000110010",
  48142=>"001010110",
  48143=>"100100111",
  48144=>"000111010",
  48145=>"001001001",
  48146=>"100111010",
  48147=>"110100110",
  48148=>"011001000",
  48149=>"000010010",
  48150=>"110111111",
  48151=>"001110001",
  48152=>"011100000",
  48153=>"001111010",
  48154=>"011000111",
  48155=>"000011011",
  48156=>"011000000",
  48157=>"101001101",
  48158=>"001000010",
  48159=>"111100110",
  48160=>"111011110",
  48161=>"100110011",
  48162=>"010110000",
  48163=>"100001100",
  48164=>"101110101",
  48165=>"011110010",
  48166=>"011000011",
  48167=>"011100110",
  48168=>"010011000",
  48169=>"111111110",
  48170=>"000011011",
  48171=>"101000101",
  48172=>"010000000",
  48173=>"011001101",
  48174=>"001010110",
  48175=>"101111111",
  48176=>"100111100",
  48177=>"111001000",
  48178=>"010111011",
  48179=>"111011110",
  48180=>"100110010",
  48181=>"011001110",
  48182=>"111111000",
  48183=>"011000101",
  48184=>"101001000",
  48185=>"101011000",
  48186=>"000100111",
  48187=>"111110111",
  48188=>"001011001",
  48189=>"111110101",
  48190=>"001110001",
  48191=>"100010010",
  48192=>"001000101",
  48193=>"011100100",
  48194=>"111111000",
  48195=>"011101001",
  48196=>"000000000",
  48197=>"110110111",
  48198=>"011100010",
  48199=>"010001101",
  48200=>"010000000",
  48201=>"001010011",
  48202=>"110011111",
  48203=>"001001111",
  48204=>"111101001",
  48205=>"100000000",
  48206=>"010101100",
  48207=>"011000001",
  48208=>"110111101",
  48209=>"110111101",
  48210=>"110000110",
  48211=>"001001100",
  48212=>"101101111",
  48213=>"000000100",
  48214=>"000010110",
  48215=>"001100010",
  48216=>"101000110",
  48217=>"110010111",
  48218=>"111010010",
  48219=>"010110100",
  48220=>"100111000",
  48221=>"110001001",
  48222=>"000110110",
  48223=>"000101101",
  48224=>"111001101",
  48225=>"111011111",
  48226=>"010011111",
  48227=>"100000010",
  48228=>"101010110",
  48229=>"110011111",
  48230=>"110001100",
  48231=>"011011011",
  48232=>"110101100",
  48233=>"100000000",
  48234=>"011010101",
  48235=>"000100110",
  48236=>"001001001",
  48237=>"010110010",
  48238=>"100111001",
  48239=>"001110010",
  48240=>"001011000",
  48241=>"000000100",
  48242=>"001101011",
  48243=>"111011110",
  48244=>"001100100",
  48245=>"000011000",
  48246=>"111111111",
  48247=>"000101011",
  48248=>"010111000",
  48249=>"001001010",
  48250=>"101100000",
  48251=>"100101001",
  48252=>"111010101",
  48253=>"110001000",
  48254=>"000100011",
  48255=>"100000000",
  48256=>"000001010",
  48257=>"000111111",
  48258=>"010000111",
  48259=>"100111111",
  48260=>"100000100",
  48261=>"100111110",
  48262=>"100011000",
  48263=>"001000110",
  48264=>"111111110",
  48265=>"000101001",
  48266=>"110000001",
  48267=>"110000011",
  48268=>"010001000",
  48269=>"001111101",
  48270=>"011100111",
  48271=>"100100111",
  48272=>"000011100",
  48273=>"000100101",
  48274=>"010100010",
  48275=>"001111010",
  48276=>"111001000",
  48277=>"010100011",
  48278=>"000101100",
  48279=>"000101001",
  48280=>"100101011",
  48281=>"000101000",
  48282=>"010001010",
  48283=>"011001001",
  48284=>"101011110",
  48285=>"000100000",
  48286=>"000000111",
  48287=>"000000000",
  48288=>"010111001",
  48289=>"011011010",
  48290=>"111001010",
  48291=>"110000011",
  48292=>"010101110",
  48293=>"000000000",
  48294=>"011000100",
  48295=>"000100100",
  48296=>"011000010",
  48297=>"110101010",
  48298=>"000000100",
  48299=>"101011010",
  48300=>"101011011",
  48301=>"010011011",
  48302=>"100000010",
  48303=>"010000100",
  48304=>"011000101",
  48305=>"111001101",
  48306=>"110010000",
  48307=>"011101011",
  48308=>"010001110",
  48309=>"001110100",
  48310=>"100000000",
  48311=>"011011111",
  48312=>"000110000",
  48313=>"100000111",
  48314=>"000011011",
  48315=>"101010000",
  48316=>"111101011",
  48317=>"010011000",
  48318=>"000100111",
  48319=>"000001010",
  48320=>"110101111",
  48321=>"000101100",
  48322=>"101100111",
  48323=>"010110111",
  48324=>"111000111",
  48325=>"000000001",
  48326=>"100010001",
  48327=>"101100000",
  48328=>"100101110",
  48329=>"000111111",
  48330=>"100101111",
  48331=>"110111111",
  48332=>"101101111",
  48333=>"000001011",
  48334=>"100111110",
  48335=>"000000110",
  48336=>"001010110",
  48337=>"000010100",
  48338=>"001010110",
  48339=>"110001010",
  48340=>"000100110",
  48341=>"011000001",
  48342=>"011101110",
  48343=>"001111000",
  48344=>"000010000",
  48345=>"000110101",
  48346=>"000011110",
  48347=>"011000010",
  48348=>"010111011",
  48349=>"000011101",
  48350=>"000110010",
  48351=>"101111110",
  48352=>"011010101",
  48353=>"011110000",
  48354=>"001111100",
  48355=>"101001111",
  48356=>"011110111",
  48357=>"110101101",
  48358=>"110010011",
  48359=>"101010110",
  48360=>"001001011",
  48361=>"111011000",
  48362=>"101100000",
  48363=>"101110110",
  48364=>"011011000",
  48365=>"110001111",
  48366=>"000101000",
  48367=>"011101000",
  48368=>"011100001",
  48369=>"000111011",
  48370=>"100101110",
  48371=>"000110001",
  48372=>"110010110",
  48373=>"011001000",
  48374=>"000111001",
  48375=>"010101111",
  48376=>"001010001",
  48377=>"010100010",
  48378=>"111011111",
  48379=>"000011000",
  48380=>"011001001",
  48381=>"001100010",
  48382=>"001010000",
  48383=>"111011011",
  48384=>"010010101",
  48385=>"111011001",
  48386=>"110101110",
  48387=>"010001001",
  48388=>"100101011",
  48389=>"000001000",
  48390=>"011011101",
  48391=>"111011001",
  48392=>"011011010",
  48393=>"000001010",
  48394=>"111110001",
  48395=>"000001100",
  48396=>"110111010",
  48397=>"100001000",
  48398=>"100111100",
  48399=>"001000001",
  48400=>"101100111",
  48401=>"011111000",
  48402=>"101000100",
  48403=>"100011111",
  48404=>"000000100",
  48405=>"110000111",
  48406=>"011101101",
  48407=>"101111111",
  48408=>"000000001",
  48409=>"101000010",
  48410=>"110000011",
  48411=>"100101101",
  48412=>"010000010",
  48413=>"110110100",
  48414=>"000001111",
  48415=>"100001000",
  48416=>"100010111",
  48417=>"111011000",
  48418=>"111011100",
  48419=>"000101101",
  48420=>"100111111",
  48421=>"011000010",
  48422=>"100111111",
  48423=>"100100110",
  48424=>"110111000",
  48425=>"110000010",
  48426=>"001011111",
  48427=>"101110100",
  48428=>"111010101",
  48429=>"010011000",
  48430=>"111001001",
  48431=>"100100011",
  48432=>"101110000",
  48433=>"100010001",
  48434=>"011100000",
  48435=>"001100111",
  48436=>"011111011",
  48437=>"000101000",
  48438=>"000001001",
  48439=>"001001110",
  48440=>"111100110",
  48441=>"100100011",
  48442=>"101111010",
  48443=>"111111101",
  48444=>"110100001",
  48445=>"111100011",
  48446=>"000110111",
  48447=>"011001000",
  48448=>"111100110",
  48449=>"111101001",
  48450=>"110100000",
  48451=>"110111000",
  48452=>"001100111",
  48453=>"000100010",
  48454=>"000010001",
  48455=>"010010111",
  48456=>"110010110",
  48457=>"100011000",
  48458=>"111110010",
  48459=>"010010000",
  48460=>"111011011",
  48461=>"111000001",
  48462=>"001010110",
  48463=>"010000101",
  48464=>"100001010",
  48465=>"110000011",
  48466=>"000010110",
  48467=>"111001110",
  48468=>"100011100",
  48469=>"101100011",
  48470=>"000101111",
  48471=>"110011011",
  48472=>"001010011",
  48473=>"010111001",
  48474=>"001000100",
  48475=>"111110100",
  48476=>"101011110",
  48477=>"111110001",
  48478=>"101110011",
  48479=>"001000001",
  48480=>"000111101",
  48481=>"000010100",
  48482=>"010100111",
  48483=>"001101000",
  48484=>"011111101",
  48485=>"101000001",
  48486=>"100001101",
  48487=>"101001101",
  48488=>"010011111",
  48489=>"001110000",
  48490=>"110110101",
  48491=>"111010110",
  48492=>"111101001",
  48493=>"101011011",
  48494=>"100000010",
  48495=>"111001011",
  48496=>"101101001",
  48497=>"000100011",
  48498=>"011000111",
  48499=>"010111001",
  48500=>"111000010",
  48501=>"000011010",
  48502=>"001101010",
  48503=>"010110110",
  48504=>"101010111",
  48505=>"010101000",
  48506=>"000000101",
  48507=>"100110101",
  48508=>"011000110",
  48509=>"001111110",
  48510=>"110000101",
  48511=>"001101111",
  48512=>"111101110",
  48513=>"100111010",
  48514=>"100010111",
  48515=>"100010100",
  48516=>"001110101",
  48517=>"001001110",
  48518=>"101111111",
  48519=>"100100101",
  48520=>"110101001",
  48521=>"000001010",
  48522=>"000001010",
  48523=>"110010010",
  48524=>"001001001",
  48525=>"011011001",
  48526=>"011111111",
  48527=>"011111010",
  48528=>"001000111",
  48529=>"101100110",
  48530=>"011100001",
  48531=>"011100000",
  48532=>"001000111",
  48533=>"000000000",
  48534=>"100110110",
  48535=>"011000001",
  48536=>"110000011",
  48537=>"011000110",
  48538=>"001000001",
  48539=>"111001000",
  48540=>"111111001",
  48541=>"001111100",
  48542=>"001100100",
  48543=>"111111101",
  48544=>"000111110",
  48545=>"110100001",
  48546=>"001110010",
  48547=>"010111011",
  48548=>"000111100",
  48549=>"001111011",
  48550=>"011001010",
  48551=>"010110001",
  48552=>"000001001",
  48553=>"011110110",
  48554=>"000100101",
  48555=>"000001110",
  48556=>"010111111",
  48557=>"100100011",
  48558=>"111110101",
  48559=>"010010011",
  48560=>"001110010",
  48561=>"110101111",
  48562=>"001010000",
  48563=>"100111010",
  48564=>"110001000",
  48565=>"001101100",
  48566=>"011111101",
  48567=>"011001000",
  48568=>"010111001",
  48569=>"110010011",
  48570=>"000001000",
  48571=>"011010101",
  48572=>"000000111",
  48573=>"101100011",
  48574=>"001010110",
  48575=>"110111000",
  48576=>"011011110",
  48577=>"001100101",
  48578=>"001101100",
  48579=>"111111001",
  48580=>"100101111",
  48581=>"011011010",
  48582=>"110011100",
  48583=>"100000101",
  48584=>"111100101",
  48585=>"101101111",
  48586=>"000111000",
  48587=>"000110111",
  48588=>"011110110",
  48589=>"101111111",
  48590=>"100100000",
  48591=>"111010011",
  48592=>"000101011",
  48593=>"010111010",
  48594=>"010100111",
  48595=>"010001010",
  48596=>"001101100",
  48597=>"000010011",
  48598=>"000011000",
  48599=>"011010010",
  48600=>"101100011",
  48601=>"000101000",
  48602=>"011000000",
  48603=>"011001000",
  48604=>"010010111",
  48605=>"111011101",
  48606=>"000101011",
  48607=>"110100000",
  48608=>"010001101",
  48609=>"000010000",
  48610=>"100110110",
  48611=>"111110101",
  48612=>"111000100",
  48613=>"101000011",
  48614=>"010001110",
  48615=>"011101111",
  48616=>"000011111",
  48617=>"101000010",
  48618=>"100011101",
  48619=>"000101100",
  48620=>"010000101",
  48621=>"111010011",
  48622=>"110110000",
  48623=>"101100011",
  48624=>"101101000",
  48625=>"010100001",
  48626=>"001000110",
  48627=>"110011001",
  48628=>"111000000",
  48629=>"101101110",
  48630=>"101001110",
  48631=>"011110111",
  48632=>"011001100",
  48633=>"010011000",
  48634=>"111011010",
  48635=>"100010110",
  48636=>"101101110",
  48637=>"010100111",
  48638=>"010101000",
  48639=>"100100011",
  48640=>"100001010",
  48641=>"000010110",
  48642=>"101011011",
  48643=>"101011110",
  48644=>"001010010",
  48645=>"110110011",
  48646=>"110101001",
  48647=>"111111110",
  48648=>"000010011",
  48649=>"010010101",
  48650=>"000111001",
  48651=>"010110000",
  48652=>"010111000",
  48653=>"110010010",
  48654=>"100000111",
  48655=>"011000011",
  48656=>"000111011",
  48657=>"111111001",
  48658=>"111011101",
  48659=>"011001010",
  48660=>"000110001",
  48661=>"010001100",
  48662=>"111001101",
  48663=>"101001000",
  48664=>"001011111",
  48665=>"000100101",
  48666=>"001010110",
  48667=>"101010001",
  48668=>"101010000",
  48669=>"111001000",
  48670=>"110110111",
  48671=>"011110000",
  48672=>"001010101",
  48673=>"011011000",
  48674=>"111100101",
  48675=>"101010101",
  48676=>"110001011",
  48677=>"110111101",
  48678=>"110110000",
  48679=>"100101011",
  48680=>"010110100",
  48681=>"011010000",
  48682=>"001000010",
  48683=>"010010110",
  48684=>"110100010",
  48685=>"001001001",
  48686=>"011111111",
  48687=>"010011111",
  48688=>"000000010",
  48689=>"011010101",
  48690=>"110111101",
  48691=>"110000101",
  48692=>"000000011",
  48693=>"000111010",
  48694=>"000100011",
  48695=>"101010100",
  48696=>"111110111",
  48697=>"110111001",
  48698=>"000011100",
  48699=>"000111001",
  48700=>"010101001",
  48701=>"100111010",
  48702=>"111000110",
  48703=>"011100111",
  48704=>"111110101",
  48705=>"111011110",
  48706=>"000000000",
  48707=>"100110011",
  48708=>"000011111",
  48709=>"110011010",
  48710=>"000000010",
  48711=>"011000101",
  48712=>"001010000",
  48713=>"100001011",
  48714=>"100011111",
  48715=>"001011101",
  48716=>"111110111",
  48717=>"011100100",
  48718=>"101110010",
  48719=>"110111000",
  48720=>"111000011",
  48721=>"100101110",
  48722=>"011111100",
  48723=>"011111011",
  48724=>"111111000",
  48725=>"101001010",
  48726=>"101111100",
  48727=>"000100001",
  48728=>"000011001",
  48729=>"100111110",
  48730=>"000010001",
  48731=>"000100010",
  48732=>"110101000",
  48733=>"101110010",
  48734=>"101111111",
  48735=>"111011000",
  48736=>"110101100",
  48737=>"010111010",
  48738=>"001100000",
  48739=>"001000111",
  48740=>"010101011",
  48741=>"111011100",
  48742=>"000001111",
  48743=>"101011111",
  48744=>"110011111",
  48745=>"100100011",
  48746=>"010111100",
  48747=>"011001010",
  48748=>"111010110",
  48749=>"010010110",
  48750=>"111101110",
  48751=>"011111110",
  48752=>"011001001",
  48753=>"000000100",
  48754=>"011101010",
  48755=>"001010011",
  48756=>"111000011",
  48757=>"001111100",
  48758=>"011011001",
  48759=>"100010001",
  48760=>"100011000",
  48761=>"001011100",
  48762=>"111010101",
  48763=>"011100011",
  48764=>"110010110",
  48765=>"011101011",
  48766=>"110111100",
  48767=>"001001101",
  48768=>"011100110",
  48769=>"110010101",
  48770=>"000101110",
  48771=>"010010000",
  48772=>"101101011",
  48773=>"001011110",
  48774=>"000011111",
  48775=>"000001001",
  48776=>"101011000",
  48777=>"011000111",
  48778=>"111111010",
  48779=>"110111000",
  48780=>"100000100",
  48781=>"100101010",
  48782=>"010010100",
  48783=>"010000111",
  48784=>"111010010",
  48785=>"111111101",
  48786=>"010000011",
  48787=>"100100001",
  48788=>"000001001",
  48789=>"001001101",
  48790=>"110011101",
  48791=>"101111101",
  48792=>"100111101",
  48793=>"000111000",
  48794=>"100110011",
  48795=>"010011101",
  48796=>"001010011",
  48797=>"110010100",
  48798=>"111100111",
  48799=>"001110000",
  48800=>"000000100",
  48801=>"111101010",
  48802=>"111100111",
  48803=>"011001111",
  48804=>"001010001",
  48805=>"101101111",
  48806=>"111100100",
  48807=>"001101010",
  48808=>"110110010",
  48809=>"110100000",
  48810=>"110100111",
  48811=>"000100010",
  48812=>"010011000",
  48813=>"010000100",
  48814=>"111100101",
  48815=>"000010101",
  48816=>"000001100",
  48817=>"100001010",
  48818=>"010111100",
  48819=>"010001000",
  48820=>"001000000",
  48821=>"000010101",
  48822=>"000110010",
  48823=>"011011101",
  48824=>"100010000",
  48825=>"000001100",
  48826=>"100001111",
  48827=>"101110111",
  48828=>"000010111",
  48829=>"101000001",
  48830=>"000011000",
  48831=>"011000001",
  48832=>"000111010",
  48833=>"101011111",
  48834=>"111101101",
  48835=>"110110110",
  48836=>"100000111",
  48837=>"111011011",
  48838=>"110111101",
  48839=>"010110111",
  48840=>"100100001",
  48841=>"011000001",
  48842=>"001001010",
  48843=>"100001000",
  48844=>"010001100",
  48845=>"010100000",
  48846=>"010111111",
  48847=>"100100010",
  48848=>"010011000",
  48849=>"010111100",
  48850=>"000010010",
  48851=>"110011010",
  48852=>"000000111",
  48853=>"000100010",
  48854=>"001101100",
  48855=>"110100001",
  48856=>"000110110",
  48857=>"011000110",
  48858=>"111000100",
  48859=>"011110010",
  48860=>"001101111",
  48861=>"011100000",
  48862=>"000101101",
  48863=>"100111110",
  48864=>"110010000",
  48865=>"001010010",
  48866=>"000101001",
  48867=>"100010000",
  48868=>"101100111",
  48869=>"100011110",
  48870=>"000000101",
  48871=>"010000000",
  48872=>"010011100",
  48873=>"111100101",
  48874=>"011010001",
  48875=>"001111110",
  48876=>"000100010",
  48877=>"111010110",
  48878=>"001000110",
  48879=>"110001101",
  48880=>"000000010",
  48881=>"000100000",
  48882=>"000010010",
  48883=>"111111001",
  48884=>"000101001",
  48885=>"110100000",
  48886=>"010111111",
  48887=>"111001010",
  48888=>"101110111",
  48889=>"000011001",
  48890=>"110001101",
  48891=>"001101001",
  48892=>"111111110",
  48893=>"101110100",
  48894=>"000011100",
  48895=>"110000000",
  48896=>"000000100",
  48897=>"100011100",
  48898=>"011110011",
  48899=>"000000010",
  48900=>"111110110",
  48901=>"100110001",
  48902=>"100100111",
  48903=>"101010001",
  48904=>"000110111",
  48905=>"100001010",
  48906=>"110010111",
  48907=>"011100111",
  48908=>"010011111",
  48909=>"001000011",
  48910=>"111010001",
  48911=>"101110011",
  48912=>"111111010",
  48913=>"101000010",
  48914=>"100101011",
  48915=>"110111000",
  48916=>"010001111",
  48917=>"011101010",
  48918=>"101001100",
  48919=>"100011111",
  48920=>"011000100",
  48921=>"100100111",
  48922=>"011010010",
  48923=>"101010110",
  48924=>"110011110",
  48925=>"100001010",
  48926=>"111011100",
  48927=>"011110110",
  48928=>"000101110",
  48929=>"101000001",
  48930=>"000100001",
  48931=>"011000000",
  48932=>"000011011",
  48933=>"110110100",
  48934=>"010000010",
  48935=>"010101000",
  48936=>"111101111",
  48937=>"100011100",
  48938=>"010101001",
  48939=>"100000100",
  48940=>"111011111",
  48941=>"110011001",
  48942=>"001000000",
  48943=>"000100010",
  48944=>"010111010",
  48945=>"001010110",
  48946=>"000111000",
  48947=>"001111111",
  48948=>"010111110",
  48949=>"011110111",
  48950=>"011100111",
  48951=>"000010001",
  48952=>"101100110",
  48953=>"101100111",
  48954=>"110101001",
  48955=>"000110111",
  48956=>"000111011",
  48957=>"111100000",
  48958=>"001111011",
  48959=>"001100110",
  48960=>"000001111",
  48961=>"001110001",
  48962=>"110111011",
  48963=>"001111000",
  48964=>"110110011",
  48965=>"010010101",
  48966=>"011001011",
  48967=>"011010000",
  48968=>"111010101",
  48969=>"010000100",
  48970=>"001100110",
  48971=>"011111001",
  48972=>"000001100",
  48973=>"110000100",
  48974=>"110110101",
  48975=>"001011001",
  48976=>"110011110",
  48977=>"110110111",
  48978=>"010101100",
  48979=>"010000110",
  48980=>"010110111",
  48981=>"111111010",
  48982=>"101111010",
  48983=>"001110011",
  48984=>"001101100",
  48985=>"000110111",
  48986=>"111100100",
  48987=>"111111100",
  48988=>"010100100",
  48989=>"011001100",
  48990=>"011010111",
  48991=>"101111110",
  48992=>"011010011",
  48993=>"010111101",
  48994=>"110000000",
  48995=>"000111001",
  48996=>"010000111",
  48997=>"101111000",
  48998=>"010110100",
  48999=>"100010100",
  49000=>"110101001",
  49001=>"001111010",
  49002=>"111000110",
  49003=>"111011101",
  49004=>"010111100",
  49005=>"000001100",
  49006=>"000111000",
  49007=>"110010000",
  49008=>"010101100",
  49009=>"101100110",
  49010=>"101110100",
  49011=>"010111101",
  49012=>"111101000",
  49013=>"010000100",
  49014=>"010000010",
  49015=>"010100100",
  49016=>"100010011",
  49017=>"101101111",
  49018=>"001001000",
  49019=>"100100000",
  49020=>"001000011",
  49021=>"111110101",
  49022=>"000111111",
  49023=>"001000011",
  49024=>"111110010",
  49025=>"100101011",
  49026=>"011011001",
  49027=>"101101011",
  49028=>"100110111",
  49029=>"110000011",
  49030=>"110111001",
  49031=>"001110101",
  49032=>"100110010",
  49033=>"000001000",
  49034=>"111101100",
  49035=>"010001100",
  49036=>"100011011",
  49037=>"011110001",
  49038=>"010011011",
  49039=>"111110111",
  49040=>"111110001",
  49041=>"110000001",
  49042=>"000110111",
  49043=>"001000010",
  49044=>"111100110",
  49045=>"101100000",
  49046=>"100100001",
  49047=>"110010101",
  49048=>"110000000",
  49049=>"111001100",
  49050=>"111000110",
  49051=>"100001110",
  49052=>"111111011",
  49053=>"001111101",
  49054=>"100111101",
  49055=>"110001101",
  49056=>"010000010",
  49057=>"101001000",
  49058=>"001110011",
  49059=>"010100010",
  49060=>"010111101",
  49061=>"111011011",
  49062=>"101100011",
  49063=>"011100100",
  49064=>"000000010",
  49065=>"101101000",
  49066=>"111111110",
  49067=>"010001001",
  49068=>"001101100",
  49069=>"000010101",
  49070=>"111110110",
  49071=>"001010000",
  49072=>"101001111",
  49073=>"110101010",
  49074=>"110000000",
  49075=>"110000111",
  49076=>"101100001",
  49077=>"111011110",
  49078=>"101000000",
  49079=>"100000011",
  49080=>"010111101",
  49081=>"010100011",
  49082=>"100001011",
  49083=>"110010011",
  49084=>"001000111",
  49085=>"001010010",
  49086=>"110000010",
  49087=>"100011000",
  49088=>"100100000",
  49089=>"111111000",
  49090=>"110010101",
  49091=>"001000010",
  49092=>"101111011",
  49093=>"001100100",
  49094=>"000010011",
  49095=>"011101101",
  49096=>"000111111",
  49097=>"101101110",
  49098=>"000010100",
  49099=>"101000101",
  49100=>"010101000",
  49101=>"001010101",
  49102=>"110010001",
  49103=>"011001110",
  49104=>"111111101",
  49105=>"111101000",
  49106=>"110110000",
  49107=>"011011100",
  49108=>"101000101",
  49109=>"011001000",
  49110=>"010110100",
  49111=>"010001110",
  49112=>"100101011",
  49113=>"000110010",
  49114=>"100100010",
  49115=>"010000000",
  49116=>"000110000",
  49117=>"000001110",
  49118=>"001101110",
  49119=>"110000000",
  49120=>"110101011",
  49121=>"001011000",
  49122=>"110010001",
  49123=>"100000000",
  49124=>"001101110",
  49125=>"110000101",
  49126=>"110100111",
  49127=>"111000000",
  49128=>"110100000",
  49129=>"011000011",
  49130=>"110110111",
  49131=>"100000101",
  49132=>"000011100",
  49133=>"011111010",
  49134=>"100011000",
  49135=>"111010110",
  49136=>"100110110",
  49137=>"001101011",
  49138=>"100011111",
  49139=>"100100011",
  49140=>"100110110",
  49141=>"010010010",
  49142=>"111110110",
  49143=>"101010101",
  49144=>"000001000",
  49145=>"110110001",
  49146=>"010010000",
  49147=>"001001000",
  49148=>"011101010",
  49149=>"001001111",
  49150=>"001001001",
  49151=>"011000001",
  49152=>"000011110",
  49153=>"001100010",
  49154=>"001001111",
  49155=>"001100010",
  49156=>"110100101",
  49157=>"111000110",
  49158=>"110010001",
  49159=>"101110111",
  49160=>"000001000",
  49161=>"000001100",
  49162=>"010100001",
  49163=>"100101110",
  49164=>"010111101",
  49165=>"000100010",
  49166=>"111100111",
  49167=>"110111011",
  49168=>"010100010",
  49169=>"110010001",
  49170=>"001110111",
  49171=>"111110111",
  49172=>"000110111",
  49173=>"110000010",
  49174=>"011010100",
  49175=>"001101110",
  49176=>"110100100",
  49177=>"000110011",
  49178=>"111111101",
  49179=>"001110101",
  49180=>"000011001",
  49181=>"111011000",
  49182=>"111101011",
  49183=>"110011101",
  49184=>"100010001",
  49185=>"100000001",
  49186=>"010000110",
  49187=>"011001101",
  49188=>"000001110",
  49189=>"010101100",
  49190=>"110010101",
  49191=>"101001000",
  49192=>"001001101",
  49193=>"100000101",
  49194=>"101011100",
  49195=>"111100110",
  49196=>"100001100",
  49197=>"000011101",
  49198=>"100000010",
  49199=>"011000111",
  49200=>"111110010",
  49201=>"010011010",
  49202=>"011010001",
  49203=>"101110101",
  49204=>"011100101",
  49205=>"001111001",
  49206=>"000100011",
  49207=>"010110001",
  49208=>"111100001",
  49209=>"000111101",
  49210=>"001010010",
  49211=>"101110011",
  49212=>"001000001",
  49213=>"000001101",
  49214=>"101011001",
  49215=>"000010111",
  49216=>"000000011",
  49217=>"000000000",
  49218=>"010001000",
  49219=>"101001110",
  49220=>"101110111",
  49221=>"110011000",
  49222=>"000011010",
  49223=>"011111000",
  49224=>"101101101",
  49225=>"011111001",
  49226=>"100111101",
  49227=>"000000011",
  49228=>"111100010",
  49229=>"111111110",
  49230=>"100001110",
  49231=>"101001011",
  49232=>"110110001",
  49233=>"000011110",
  49234=>"011010000",
  49235=>"111001100",
  49236=>"111110010",
  49237=>"101000110",
  49238=>"110001111",
  49239=>"100001000",
  49240=>"011011110",
  49241=>"010001001",
  49242=>"010011010",
  49243=>"111100111",
  49244=>"101100101",
  49245=>"111100000",
  49246=>"000100000",
  49247=>"111101110",
  49248=>"011001001",
  49249=>"010001000",
  49250=>"110101101",
  49251=>"100100101",
  49252=>"001000100",
  49253=>"111100101",
  49254=>"010101101",
  49255=>"000010001",
  49256=>"001111001",
  49257=>"011111010",
  49258=>"101111101",
  49259=>"000010011",
  49260=>"101100100",
  49261=>"000101010",
  49262=>"011101101",
  49263=>"000000001",
  49264=>"011000000",
  49265=>"010011011",
  49266=>"010010101",
  49267=>"011111100",
  49268=>"110000010",
  49269=>"111111011",
  49270=>"110011011",
  49271=>"000100010",
  49272=>"001000000",
  49273=>"110100101",
  49274=>"111011000",
  49275=>"000011010",
  49276=>"001101111",
  49277=>"010010011",
  49278=>"101100011",
  49279=>"001100110",
  49280=>"100101101",
  49281=>"111111111",
  49282=>"100111101",
  49283=>"001011000",
  49284=>"001101010",
  49285=>"000100001",
  49286=>"001001111",
  49287=>"011100110",
  49288=>"001100101",
  49289=>"001010100",
  49290=>"001011011",
  49291=>"011011111",
  49292=>"110111110",
  49293=>"101011100",
  49294=>"100010001",
  49295=>"111110101",
  49296=>"110101111",
  49297=>"001110001",
  49298=>"001000111",
  49299=>"010101010",
  49300=>"011110110",
  49301=>"010101011",
  49302=>"100100100",
  49303=>"100010110",
  49304=>"000001001",
  49305=>"010101000",
  49306=>"000010011",
  49307=>"010011010",
  49308=>"100111100",
  49309=>"000110000",
  49310=>"110000001",
  49311=>"011001110",
  49312=>"100001011",
  49313=>"000010110",
  49314=>"001000011",
  49315=>"000001101",
  49316=>"111011100",
  49317=>"010101011",
  49318=>"111111100",
  49319=>"100010111",
  49320=>"110001001",
  49321=>"111110110",
  49322=>"001001101",
  49323=>"000010010",
  49324=>"101100011",
  49325=>"111111011",
  49326=>"011111010",
  49327=>"011110010",
  49328=>"000000101",
  49329=>"010110111",
  49330=>"011111110",
  49331=>"110110101",
  49332=>"000111001",
  49333=>"010011101",
  49334=>"111111101",
  49335=>"000100101",
  49336=>"101010010",
  49337=>"011001110",
  49338=>"010001011",
  49339=>"011100101",
  49340=>"110010110",
  49341=>"001011100",
  49342=>"001011010",
  49343=>"001000000",
  49344=>"100101110",
  49345=>"000011111",
  49346=>"000111010",
  49347=>"100111010",
  49348=>"101010001",
  49349=>"000101010",
  49350=>"101100000",
  49351=>"011011011",
  49352=>"010000000",
  49353=>"100000001",
  49354=>"011110011",
  49355=>"001100110",
  49356=>"110010001",
  49357=>"101010101",
  49358=>"111111000",
  49359=>"000011011",
  49360=>"001110010",
  49361=>"110000010",
  49362=>"110000000",
  49363=>"010100111",
  49364=>"001010101",
  49365=>"000000000",
  49366=>"111001011",
  49367=>"111011011",
  49368=>"100100001",
  49369=>"110010000",
  49370=>"010011111",
  49371=>"101100100",
  49372=>"011100011",
  49373=>"001001000",
  49374=>"000100001",
  49375=>"111100101",
  49376=>"000110100",
  49377=>"101111111",
  49378=>"111101001",
  49379=>"111011100",
  49380=>"101011010",
  49381=>"100000010",
  49382=>"000010001",
  49383=>"111001011",
  49384=>"001011001",
  49385=>"101001011",
  49386=>"011110101",
  49387=>"111001100",
  49388=>"101100001",
  49389=>"010110010",
  49390=>"100001100",
  49391=>"101010000",
  49392=>"111010101",
  49393=>"101010000",
  49394=>"101011100",
  49395=>"101010111",
  49396=>"100100100",
  49397=>"110011101",
  49398=>"101101010",
  49399=>"100000110",
  49400=>"101000111",
  49401=>"010001000",
  49402=>"011101110",
  49403=>"101000100",
  49404=>"000111000",
  49405=>"000100011",
  49406=>"010011010",
  49407=>"111110001",
  49408=>"011011100",
  49409=>"100001100",
  49410=>"111110011",
  49411=>"000000111",
  49412=>"100000011",
  49413=>"000001011",
  49414=>"101101011",
  49415=>"011010011",
  49416=>"101001001",
  49417=>"101101100",
  49418=>"101000001",
  49419=>"011110011",
  49420=>"011010111",
  49421=>"111001111",
  49422=>"100100000",
  49423=>"111110111",
  49424=>"111111110",
  49425=>"000010110",
  49426=>"101110001",
  49427=>"010000001",
  49428=>"100010000",
  49429=>"001100011",
  49430=>"011110000",
  49431=>"100001010",
  49432=>"110110110",
  49433=>"010101111",
  49434=>"101000100",
  49435=>"011001100",
  49436=>"010110110",
  49437=>"000101111",
  49438=>"100001010",
  49439=>"100101101",
  49440=>"010000101",
  49441=>"010111110",
  49442=>"011000101",
  49443=>"111101011",
  49444=>"110011100",
  49445=>"100011100",
  49446=>"001111100",
  49447=>"011010000",
  49448=>"000011010",
  49449=>"011001011",
  49450=>"110110111",
  49451=>"001101111",
  49452=>"101000010",
  49453=>"010111110",
  49454=>"100000010",
  49455=>"011101010",
  49456=>"110010011",
  49457=>"100001011",
  49458=>"101000001",
  49459=>"000000101",
  49460=>"100001101",
  49461=>"001011000",
  49462=>"100111011",
  49463=>"001000110",
  49464=>"011000100",
  49465=>"111000111",
  49466=>"001010010",
  49467=>"101010101",
  49468=>"000010101",
  49469=>"011101001",
  49470=>"010001001",
  49471=>"100000010",
  49472=>"010011100",
  49473=>"110110110",
  49474=>"111110110",
  49475=>"100110000",
  49476=>"000010110",
  49477=>"111011001",
  49478=>"001100001",
  49479=>"001010011",
  49480=>"101111100",
  49481=>"011011011",
  49482=>"010010101",
  49483=>"100000000",
  49484=>"111111001",
  49485=>"001011010",
  49486=>"111100110",
  49487=>"110110000",
  49488=>"000111101",
  49489=>"011100111",
  49490=>"010000101",
  49491=>"011010111",
  49492=>"010111110",
  49493=>"100111110",
  49494=>"010011001",
  49495=>"111011111",
  49496=>"111101110",
  49497=>"110110110",
  49498=>"110000110",
  49499=>"001000101",
  49500=>"111000110",
  49501=>"110100010",
  49502=>"001011000",
  49503=>"100100100",
  49504=>"100011010",
  49505=>"010100110",
  49506=>"111011000",
  49507=>"100000010",
  49508=>"000010000",
  49509=>"100011011",
  49510=>"001001100",
  49511=>"000110001",
  49512=>"010110100",
  49513=>"100001001",
  49514=>"101001000",
  49515=>"101111101",
  49516=>"001011110",
  49517=>"001111000",
  49518=>"001110001",
  49519=>"000000100",
  49520=>"110010100",
  49521=>"010110010",
  49522=>"001001100",
  49523=>"000010010",
  49524=>"111100010",
  49525=>"101100110",
  49526=>"000111001",
  49527=>"011000100",
  49528=>"011001000",
  49529=>"110001100",
  49530=>"000110000",
  49531=>"001100011",
  49532=>"011110011",
  49533=>"111010111",
  49534=>"101011110",
  49535=>"011101000",
  49536=>"000101101",
  49537=>"111000010",
  49538=>"001011010",
  49539=>"110110011",
  49540=>"001001010",
  49541=>"011100010",
  49542=>"100011000",
  49543=>"010000100",
  49544=>"000010011",
  49545=>"011110110",
  49546=>"100111110",
  49547=>"010100110",
  49548=>"101011100",
  49549=>"100111110",
  49550=>"010111100",
  49551=>"000010111",
  49552=>"010111100",
  49553=>"011000111",
  49554=>"010010010",
  49555=>"111011100",
  49556=>"000000000",
  49557=>"111110101",
  49558=>"011100010",
  49559=>"100010101",
  49560=>"011001100",
  49561=>"100101110",
  49562=>"101100000",
  49563=>"101111110",
  49564=>"100010100",
  49565=>"011111111",
  49566=>"000110000",
  49567=>"011000101",
  49568=>"101111000",
  49569=>"111001011",
  49570=>"100101110",
  49571=>"101100011",
  49572=>"111101110",
  49573=>"101110100",
  49574=>"011101000",
  49575=>"111001000",
  49576=>"011011101",
  49577=>"101111110",
  49578=>"111001000",
  49579=>"000010011",
  49580=>"010011111",
  49581=>"111100000",
  49582=>"110101110",
  49583=>"111100011",
  49584=>"101010111",
  49585=>"000111101",
  49586=>"000100101",
  49587=>"110101111",
  49588=>"100101010",
  49589=>"111100010",
  49590=>"111111100",
  49591=>"010111011",
  49592=>"101000000",
  49593=>"111101010",
  49594=>"111110111",
  49595=>"010011000",
  49596=>"011001110",
  49597=>"101011000",
  49598=>"110001111",
  49599=>"011100100",
  49600=>"000101100",
  49601=>"010100110",
  49602=>"101011011",
  49603=>"110001100",
  49604=>"010100101",
  49605=>"101011001",
  49606=>"101110000",
  49607=>"010000000",
  49608=>"111001111",
  49609=>"110010000",
  49610=>"000000000",
  49611=>"000110100",
  49612=>"010111001",
  49613=>"001011100",
  49614=>"101001111",
  49615=>"101011000",
  49616=>"011111100",
  49617=>"000011010",
  49618=>"000111000",
  49619=>"101111111",
  49620=>"001111001",
  49621=>"111111001",
  49622=>"000101010",
  49623=>"101010000",
  49624=>"001111011",
  49625=>"101000110",
  49626=>"110111111",
  49627=>"001000011",
  49628=>"101011011",
  49629=>"011100100",
  49630=>"010000011",
  49631=>"001001110",
  49632=>"010001111",
  49633=>"001111110",
  49634=>"011100100",
  49635=>"110010100",
  49636=>"110000110",
  49637=>"010100000",
  49638=>"000000010",
  49639=>"000000100",
  49640=>"000101010",
  49641=>"100111011",
  49642=>"011000010",
  49643=>"001111100",
  49644=>"000100111",
  49645=>"011000000",
  49646=>"110101011",
  49647=>"011101100",
  49648=>"101101011",
  49649=>"100001001",
  49650=>"111001111",
  49651=>"100100111",
  49652=>"010000011",
  49653=>"001111101",
  49654=>"011011001",
  49655=>"011101100",
  49656=>"000101110",
  49657=>"011011110",
  49658=>"111100011",
  49659=>"110101110",
  49660=>"110101100",
  49661=>"000010110",
  49662=>"000110110",
  49663=>"000011011",
  49664=>"000000000",
  49665=>"000100110",
  49666=>"010000000",
  49667=>"110010101",
  49668=>"110100111",
  49669=>"110010011",
  49670=>"100001011",
  49671=>"011101011",
  49672=>"111010110",
  49673=>"010110110",
  49674=>"100000000",
  49675=>"110001110",
  49676=>"010010111",
  49677=>"001000111",
  49678=>"111110101",
  49679=>"100011011",
  49680=>"100001000",
  49681=>"001101011",
  49682=>"011010011",
  49683=>"000111001",
  49684=>"100001101",
  49685=>"111000001",
  49686=>"001011101",
  49687=>"101101110",
  49688=>"000101001",
  49689=>"110101011",
  49690=>"011100011",
  49691=>"010010110",
  49692=>"100111110",
  49693=>"000101111",
  49694=>"101000000",
  49695=>"101001111",
  49696=>"000110111",
  49697=>"000011001",
  49698=>"011111010",
  49699=>"100011111",
  49700=>"110000100",
  49701=>"000011100",
  49702=>"000110100",
  49703=>"111010010",
  49704=>"111000101",
  49705=>"111001011",
  49706=>"011101100",
  49707=>"010110000",
  49708=>"011010011",
  49709=>"001010001",
  49710=>"100000100",
  49711=>"110000110",
  49712=>"010000101",
  49713=>"010100011",
  49714=>"101100000",
  49715=>"101111110",
  49716=>"011110011",
  49717=>"010010001",
  49718=>"010110100",
  49719=>"001100100",
  49720=>"111001000",
  49721=>"111100100",
  49722=>"011000001",
  49723=>"010001010",
  49724=>"101000011",
  49725=>"100010111",
  49726=>"000101010",
  49727=>"100110000",
  49728=>"100011111",
  49729=>"011010011",
  49730=>"001101101",
  49731=>"110001111",
  49732=>"011100001",
  49733=>"111111110",
  49734=>"101010001",
  49735=>"100010000",
  49736=>"011001101",
  49737=>"010100000",
  49738=>"010011000",
  49739=>"100100100",
  49740=>"010000101",
  49741=>"110110011",
  49742=>"111111111",
  49743=>"000100000",
  49744=>"110011111",
  49745=>"111000000",
  49746=>"101110111",
  49747=>"101010110",
  49748=>"101110101",
  49749=>"100110101",
  49750=>"111101111",
  49751=>"000001110",
  49752=>"000000010",
  49753=>"101101001",
  49754=>"100011001",
  49755=>"101101001",
  49756=>"010001001",
  49757=>"011000011",
  49758=>"001011100",
  49759=>"111110000",
  49760=>"111111110",
  49761=>"101101100",
  49762=>"101110001",
  49763=>"110000100",
  49764=>"110100101",
  49765=>"110100011",
  49766=>"000001100",
  49767=>"101110101",
  49768=>"001110101",
  49769=>"011011011",
  49770=>"001101001",
  49771=>"011101101",
  49772=>"100001001",
  49773=>"110011001",
  49774=>"011111010",
  49775=>"000000010",
  49776=>"011111001",
  49777=>"101110100",
  49778=>"011011000",
  49779=>"101011010",
  49780=>"110011010",
  49781=>"101100110",
  49782=>"110101001",
  49783=>"110000000",
  49784=>"111000011",
  49785=>"111111001",
  49786=>"011110001",
  49787=>"111011011",
  49788=>"001000110",
  49789=>"001000101",
  49790=>"110011011",
  49791=>"100100000",
  49792=>"000011011",
  49793=>"010011010",
  49794=>"001101100",
  49795=>"011110001",
  49796=>"001100011",
  49797=>"111110000",
  49798=>"101011010",
  49799=>"011101110",
  49800=>"111110100",
  49801=>"101010011",
  49802=>"101000100",
  49803=>"000000000",
  49804=>"000011000",
  49805=>"011000001",
  49806=>"111010000",
  49807=>"101101001",
  49808=>"100001101",
  49809=>"010011111",
  49810=>"100110111",
  49811=>"101000001",
  49812=>"000110111",
  49813=>"110011111",
  49814=>"000111110",
  49815=>"100101100",
  49816=>"100000111",
  49817=>"000010101",
  49818=>"011110100",
  49819=>"000111011",
  49820=>"000011010",
  49821=>"011000110",
  49822=>"111110110",
  49823=>"011001001",
  49824=>"000001100",
  49825=>"000001011",
  49826=>"100011101",
  49827=>"100000111",
  49828=>"000110101",
  49829=>"110011110",
  49830=>"010001001",
  49831=>"110101111",
  49832=>"111010100",
  49833=>"011101011",
  49834=>"101101110",
  49835=>"000000011",
  49836=>"101100111",
  49837=>"011100100",
  49838=>"110111100",
  49839=>"111101010",
  49840=>"100110111",
  49841=>"000100111",
  49842=>"111100000",
  49843=>"010111100",
  49844=>"011000000",
  49845=>"010100100",
  49846=>"011100111",
  49847=>"111101101",
  49848=>"000110111",
  49849=>"001111101",
  49850=>"111011011",
  49851=>"001000011",
  49852=>"010111111",
  49853=>"000011000",
  49854=>"110111100",
  49855=>"101111001",
  49856=>"111101111",
  49857=>"011111001",
  49858=>"101101110",
  49859=>"010010000",
  49860=>"100000001",
  49861=>"011110001",
  49862=>"011111000",
  49863=>"001111001",
  49864=>"000111110",
  49865=>"010100011",
  49866=>"111001001",
  49867=>"000101100",
  49868=>"011101110",
  49869=>"001101101",
  49870=>"110110101",
  49871=>"101111101",
  49872=>"001001000",
  49873=>"110111001",
  49874=>"001101100",
  49875=>"111101101",
  49876=>"110110001",
  49877=>"010110011",
  49878=>"010111010",
  49879=>"101110001",
  49880=>"010111001",
  49881=>"011011010",
  49882=>"111111001",
  49883=>"100011100",
  49884=>"100010011",
  49885=>"010111010",
  49886=>"101010001",
  49887=>"011000110",
  49888=>"101110010",
  49889=>"011000011",
  49890=>"010101101",
  49891=>"000000000",
  49892=>"101011110",
  49893=>"001111111",
  49894=>"110010101",
  49895=>"001000001",
  49896=>"101101000",
  49897=>"010110010",
  49898=>"111011000",
  49899=>"111001001",
  49900=>"011001010",
  49901=>"000010111",
  49902=>"110001110",
  49903=>"010110100",
  49904=>"010100001",
  49905=>"000000001",
  49906=>"010010010",
  49907=>"011011011",
  49908=>"000000000",
  49909=>"111111010",
  49910=>"000101011",
  49911=>"000111101",
  49912=>"011110001",
  49913=>"111001110",
  49914=>"100010000",
  49915=>"101100000",
  49916=>"011100111",
  49917=>"000001010",
  49918=>"111010101",
  49919=>"111111010",
  49920=>"011101010",
  49921=>"010110101",
  49922=>"110001100",
  49923=>"100110010",
  49924=>"011011010",
  49925=>"001001011",
  49926=>"100001100",
  49927=>"110101111",
  49928=>"100001001",
  49929=>"110011010",
  49930=>"010101100",
  49931=>"100110000",
  49932=>"111111010",
  49933=>"011011111",
  49934=>"111011001",
  49935=>"000011100",
  49936=>"110101111",
  49937=>"000110101",
  49938=>"001011111",
  49939=>"110100111",
  49940=>"110010100",
  49941=>"000011101",
  49942=>"110000100",
  49943=>"000101000",
  49944=>"000100110",
  49945=>"000100011",
  49946=>"000111001",
  49947=>"010110110",
  49948=>"101100000",
  49949=>"001000001",
  49950=>"000101111",
  49951=>"111111100",
  49952=>"110000011",
  49953=>"101100010",
  49954=>"110100000",
  49955=>"110101010",
  49956=>"001101110",
  49957=>"110010001",
  49958=>"000001010",
  49959=>"000001000",
  49960=>"011011010",
  49961=>"001100000",
  49962=>"010100000",
  49963=>"011011000",
  49964=>"101001010",
  49965=>"001011101",
  49966=>"100101111",
  49967=>"011010100",
  49968=>"101111111",
  49969=>"001110011",
  49970=>"101100011",
  49971=>"111100011",
  49972=>"101001001",
  49973=>"101000110",
  49974=>"101110100",
  49975=>"100010100",
  49976=>"101000011",
  49977=>"100100111",
  49978=>"000100100",
  49979=>"110011001",
  49980=>"001101111",
  49981=>"111010000",
  49982=>"000010001",
  49983=>"011010000",
  49984=>"100111011",
  49985=>"001000010",
  49986=>"111110111",
  49987=>"001101011",
  49988=>"001101110",
  49989=>"110111011",
  49990=>"001001101",
  49991=>"101001001",
  49992=>"101110011",
  49993=>"110000100",
  49994=>"111111000",
  49995=>"000100000",
  49996=>"000000000",
  49997=>"101101011",
  49998=>"010001110",
  49999=>"000001011",
  50000=>"000111011",
  50001=>"000000010",
  50002=>"000000001",
  50003=>"111011100",
  50004=>"000011110",
  50005=>"001000010",
  50006=>"100001101",
  50007=>"001110000",
  50008=>"100100010",
  50009=>"110011111",
  50010=>"010111111",
  50011=>"000100100",
  50012=>"111001000",
  50013=>"110100000",
  50014=>"110110100",
  50015=>"110010010",
  50016=>"111011001",
  50017=>"111111001",
  50018=>"011001010",
  50019=>"000011001",
  50020=>"100011100",
  50021=>"000100001",
  50022=>"101001011",
  50023=>"001110110",
  50024=>"110001000",
  50025=>"011010010",
  50026=>"110110111",
  50027=>"001101001",
  50028=>"111000011",
  50029=>"111100101",
  50030=>"000011110",
  50031=>"101000010",
  50032=>"111100011",
  50033=>"011010100",
  50034=>"001110000",
  50035=>"000100110",
  50036=>"010011000",
  50037=>"001001110",
  50038=>"000001101",
  50039=>"011000110",
  50040=>"010111101",
  50041=>"001101110",
  50042=>"111010010",
  50043=>"110111110",
  50044=>"100111100",
  50045=>"001110011",
  50046=>"111000010",
  50047=>"110011100",
  50048=>"111101111",
  50049=>"001110010",
  50050=>"000110111",
  50051=>"010101000",
  50052=>"011010110",
  50053=>"010010101",
  50054=>"110100100",
  50055=>"100110100",
  50056=>"101000000",
  50057=>"001000111",
  50058=>"001100011",
  50059=>"000000011",
  50060=>"110000100",
  50061=>"010101101",
  50062=>"001100001",
  50063=>"100010000",
  50064=>"110110110",
  50065=>"001011101",
  50066=>"000110000",
  50067=>"010011000",
  50068=>"100100110",
  50069=>"010100100",
  50070=>"111110011",
  50071=>"001111110",
  50072=>"111110111",
  50073=>"000010111",
  50074=>"110011000",
  50075=>"001100111",
  50076=>"100100011",
  50077=>"100011101",
  50078=>"011001010",
  50079=>"001000111",
  50080=>"100100100",
  50081=>"101001011",
  50082=>"010011001",
  50083=>"010001000",
  50084=>"110001101",
  50085=>"000100011",
  50086=>"100110011",
  50087=>"000011111",
  50088=>"000010111",
  50089=>"100100010",
  50090=>"001011011",
  50091=>"011111001",
  50092=>"001000100",
  50093=>"000010100",
  50094=>"100001111",
  50095=>"111100001",
  50096=>"010110001",
  50097=>"110111000",
  50098=>"111110100",
  50099=>"001001001",
  50100=>"000000010",
  50101=>"100110110",
  50102=>"011010010",
  50103=>"110001000",
  50104=>"110110010",
  50105=>"001000111",
  50106=>"001010100",
  50107=>"111101000",
  50108=>"000000011",
  50109=>"011001111",
  50110=>"000011010",
  50111=>"110010011",
  50112=>"111101001",
  50113=>"100101110",
  50114=>"111110111",
  50115=>"000110100",
  50116=>"000001001",
  50117=>"000000100",
  50118=>"110110010",
  50119=>"011100000",
  50120=>"001010111",
  50121=>"011001000",
  50122=>"100011100",
  50123=>"110111110",
  50124=>"101001010",
  50125=>"011111110",
  50126=>"101100010",
  50127=>"110101000",
  50128=>"101111100",
  50129=>"000101101",
  50130=>"001010010",
  50131=>"001000111",
  50132=>"101111011",
  50133=>"000010110",
  50134=>"000011111",
  50135=>"011000001",
  50136=>"000011010",
  50137=>"100011110",
  50138=>"111111011",
  50139=>"001100001",
  50140=>"111100111",
  50141=>"011100110",
  50142=>"000101101",
  50143=>"010001100",
  50144=>"101111111",
  50145=>"011001000",
  50146=>"001100001",
  50147=>"100110111",
  50148=>"010000110",
  50149=>"010100000",
  50150=>"101001101",
  50151=>"111000001",
  50152=>"000110010",
  50153=>"110111101",
  50154=>"011101010",
  50155=>"101000101",
  50156=>"001110111",
  50157=>"101000101",
  50158=>"110100110",
  50159=>"110111110",
  50160=>"010100101",
  50161=>"001010110",
  50162=>"110011010",
  50163=>"110011011",
  50164=>"111000100",
  50165=>"010010110",
  50166=>"000101111",
  50167=>"011001011",
  50168=>"000111100",
  50169=>"000111101",
  50170=>"000000011",
  50171=>"111001010",
  50172=>"001110001",
  50173=>"100001011",
  50174=>"110010011",
  50175=>"010110001",
  50176=>"000000001",
  50177=>"011101000",
  50178=>"010111000",
  50179=>"010001101",
  50180=>"010011110",
  50181=>"111000011",
  50182=>"101000000",
  50183=>"001000000",
  50184=>"001011111",
  50185=>"001101100",
  50186=>"111011101",
  50187=>"000010011",
  50188=>"111010000",
  50189=>"100000100",
  50190=>"000000011",
  50191=>"010010100",
  50192=>"101001101",
  50193=>"100100101",
  50194=>"001001110",
  50195=>"000001001",
  50196=>"100010111",
  50197=>"001010100",
  50198=>"110101010",
  50199=>"111101001",
  50200=>"010000101",
  50201=>"000111100",
  50202=>"011000101",
  50203=>"101111111",
  50204=>"010111010",
  50205=>"001011111",
  50206=>"110000000",
  50207=>"001001000",
  50208=>"100000001",
  50209=>"111110101",
  50210=>"011011000",
  50211=>"100000010",
  50212=>"101110011",
  50213=>"000011001",
  50214=>"001010010",
  50215=>"101111010",
  50216=>"001000010",
  50217=>"000110010",
  50218=>"000010111",
  50219=>"011011010",
  50220=>"000000110",
  50221=>"000111110",
  50222=>"011010100",
  50223=>"110010000",
  50224=>"110000010",
  50225=>"110111111",
  50226=>"011001000",
  50227=>"110110110",
  50228=>"111100101",
  50229=>"010001100",
  50230=>"110111110",
  50231=>"001000001",
  50232=>"111101011",
  50233=>"000011001",
  50234=>"000001011",
  50235=>"011011000",
  50236=>"001010100",
  50237=>"010111001",
  50238=>"000010000",
  50239=>"000011111",
  50240=>"000011001",
  50241=>"011010111",
  50242=>"000011110",
  50243=>"000001010",
  50244=>"101000100",
  50245=>"000101010",
  50246=>"111010101",
  50247=>"010101100",
  50248=>"000010011",
  50249=>"010000011",
  50250=>"000001000",
  50251=>"111110001",
  50252=>"110111010",
  50253=>"010101011",
  50254=>"011011001",
  50255=>"011000010",
  50256=>"011101100",
  50257=>"101000100",
  50258=>"011010011",
  50259=>"101101101",
  50260=>"011011101",
  50261=>"111111001",
  50262=>"000111001",
  50263=>"101011111",
  50264=>"111100010",
  50265=>"110100011",
  50266=>"100111010",
  50267=>"010100000",
  50268=>"100100110",
  50269=>"110100111",
  50270=>"101000100",
  50271=>"110000100",
  50272=>"111011011",
  50273=>"111101000",
  50274=>"100110101",
  50275=>"011111001",
  50276=>"100101010",
  50277=>"010010110",
  50278=>"001111100",
  50279=>"010100100",
  50280=>"111111000",
  50281=>"111011110",
  50282=>"100001100",
  50283=>"100001111",
  50284=>"001110110",
  50285=>"000000111",
  50286=>"000101001",
  50287=>"000100000",
  50288=>"111000000",
  50289=>"101110011",
  50290=>"011011000",
  50291=>"110110100",
  50292=>"111000001",
  50293=>"101010011",
  50294=>"000010011",
  50295=>"011110010",
  50296=>"010010110",
  50297=>"001000010",
  50298=>"011001110",
  50299=>"000111011",
  50300=>"010100100",
  50301=>"110100100",
  50302=>"001101110",
  50303=>"110000100",
  50304=>"010100100",
  50305=>"000011001",
  50306=>"100010100",
  50307=>"111010101",
  50308=>"100000010",
  50309=>"010110000",
  50310=>"010011000",
  50311=>"111010101",
  50312=>"011011100",
  50313=>"100100100",
  50314=>"100010001",
  50315=>"110011110",
  50316=>"101010111",
  50317=>"111101010",
  50318=>"001010000",
  50319=>"101010100",
  50320=>"010111010",
  50321=>"010101000",
  50322=>"001100001",
  50323=>"101101100",
  50324=>"110010000",
  50325=>"110011001",
  50326=>"000011110",
  50327=>"010001000",
  50328=>"010010001",
  50329=>"101101110",
  50330=>"000001100",
  50331=>"111111010",
  50332=>"100001011",
  50333=>"100110010",
  50334=>"100011100",
  50335=>"101111011",
  50336=>"011010110",
  50337=>"010111110",
  50338=>"111100011",
  50339=>"110100010",
  50340=>"111110101",
  50341=>"101000110",
  50342=>"011111001",
  50343=>"010100011",
  50344=>"011010010",
  50345=>"011111100",
  50346=>"001111101",
  50347=>"111001000",
  50348=>"011110011",
  50349=>"010000001",
  50350=>"000011001",
  50351=>"100111101",
  50352=>"010110100",
  50353=>"000011001",
  50354=>"000100000",
  50355=>"110100111",
  50356=>"110100000",
  50357=>"001110110",
  50358=>"010110000",
  50359=>"001001001",
  50360=>"101000000",
  50361=>"001111001",
  50362=>"000100011",
  50363=>"111010000",
  50364=>"111100111",
  50365=>"001010101",
  50366=>"110101011",
  50367=>"010111001",
  50368=>"011000001",
  50369=>"011110101",
  50370=>"001001000",
  50371=>"001111011",
  50372=>"000001110",
  50373=>"111001000",
  50374=>"110010110",
  50375=>"010100100",
  50376=>"100011101",
  50377=>"000001000",
  50378=>"111011110",
  50379=>"111011111",
  50380=>"100010010",
  50381=>"101101111",
  50382=>"000001100",
  50383=>"100110111",
  50384=>"001100100",
  50385=>"011100100",
  50386=>"000001000",
  50387=>"110010010",
  50388=>"001101111",
  50389=>"100101100",
  50390=>"000100110",
  50391=>"001010010",
  50392=>"100101101",
  50393=>"110000001",
  50394=>"010000011",
  50395=>"010111101",
  50396=>"100101100",
  50397=>"010000000",
  50398=>"110001011",
  50399=>"111100110",
  50400=>"000100000",
  50401=>"111100100",
  50402=>"110000001",
  50403=>"011110011",
  50404=>"111100010",
  50405=>"111010111",
  50406=>"101011100",
  50407=>"101111001",
  50408=>"111010101",
  50409=>"011100011",
  50410=>"000010000",
  50411=>"100000000",
  50412=>"111110111",
  50413=>"110001101",
  50414=>"000000111",
  50415=>"000111010",
  50416=>"011101011",
  50417=>"010001000",
  50418=>"110110010",
  50419=>"111010000",
  50420=>"011011001",
  50421=>"000010110",
  50422=>"011010101",
  50423=>"000000001",
  50424=>"010000110",
  50425=>"101111010",
  50426=>"111110001",
  50427=>"000010010",
  50428=>"110101100",
  50429=>"001100000",
  50430=>"110001000",
  50431=>"010101100",
  50432=>"000011001",
  50433=>"011111011",
  50434=>"101011111",
  50435=>"100110001",
  50436=>"100111000",
  50437=>"100100110",
  50438=>"011010001",
  50439=>"100001010",
  50440=>"001100111",
  50441=>"001000100",
  50442=>"001001000",
  50443=>"101010000",
  50444=>"101001010",
  50445=>"000111111",
  50446=>"110111100",
  50447=>"110100111",
  50448=>"110101001",
  50449=>"110100110",
  50450=>"000111010",
  50451=>"111101110",
  50452=>"110010100",
  50453=>"101110000",
  50454=>"001010101",
  50455=>"100100010",
  50456=>"000001000",
  50457=>"110111010",
  50458=>"111000100",
  50459=>"101110011",
  50460=>"100011000",
  50461=>"011101010",
  50462=>"000111110",
  50463=>"001100100",
  50464=>"000110101",
  50465=>"000010100",
  50466=>"001000010",
  50467=>"110101011",
  50468=>"001110111",
  50469=>"000010001",
  50470=>"000000100",
  50471=>"111011011",
  50472=>"001000010",
  50473=>"100001010",
  50474=>"010010111",
  50475=>"101000101",
  50476=>"010000111",
  50477=>"001111011",
  50478=>"001011100",
  50479=>"100000111",
  50480=>"001001000",
  50481=>"111010010",
  50482=>"010001111",
  50483=>"110101010",
  50484=>"000000011",
  50485=>"001000100",
  50486=>"010110000",
  50487=>"111000110",
  50488=>"010000011",
  50489=>"001001000",
  50490=>"110110110",
  50491=>"011101110",
  50492=>"010101101",
  50493=>"100011010",
  50494=>"100101000",
  50495=>"001011101",
  50496=>"000010001",
  50497=>"111001110",
  50498=>"100101010",
  50499=>"100011011",
  50500=>"011011101",
  50501=>"111001110",
  50502=>"001011101",
  50503=>"000010001",
  50504=>"111111011",
  50505=>"011001100",
  50506=>"100111111",
  50507=>"111101100",
  50508=>"000001111",
  50509=>"010111001",
  50510=>"011110111",
  50511=>"001110111",
  50512=>"100010111",
  50513=>"001011101",
  50514=>"001001011",
  50515=>"010001111",
  50516=>"101101110",
  50517=>"111010010",
  50518=>"101111110",
  50519=>"001000111",
  50520=>"000100111",
  50521=>"011111100",
  50522=>"101010110",
  50523=>"000001101",
  50524=>"100100111",
  50525=>"011111111",
  50526=>"110101000",
  50527=>"110110110",
  50528=>"001111110",
  50529=>"110011111",
  50530=>"000110101",
  50531=>"100001101",
  50532=>"110100101",
  50533=>"100100100",
  50534=>"111100010",
  50535=>"010100100",
  50536=>"001101011",
  50537=>"100010000",
  50538=>"001000101",
  50539=>"011000000",
  50540=>"011111010",
  50541=>"110001110",
  50542=>"010000011",
  50543=>"001001000",
  50544=>"010000000",
  50545=>"001010011",
  50546=>"111000011",
  50547=>"111110001",
  50548=>"001010101",
  50549=>"111101101",
  50550=>"100000110",
  50551=>"010111011",
  50552=>"101100001",
  50553=>"110111000",
  50554=>"000101111",
  50555=>"100010100",
  50556=>"010110100",
  50557=>"100110001",
  50558=>"010101011",
  50559=>"101111110",
  50560=>"111101000",
  50561=>"001001100",
  50562=>"001111110",
  50563=>"001110111",
  50564=>"011101001",
  50565=>"011000011",
  50566=>"000111101",
  50567=>"111000111",
  50568=>"000000010",
  50569=>"111000101",
  50570=>"001101101",
  50571=>"001010000",
  50572=>"010000010",
  50573=>"011100010",
  50574=>"001010100",
  50575=>"111011101",
  50576=>"101001101",
  50577=>"111010110",
  50578=>"110010010",
  50579=>"100110111",
  50580=>"011000100",
  50581=>"000011010",
  50582=>"110111100",
  50583=>"010101111",
  50584=>"000000100",
  50585=>"000100011",
  50586=>"000101000",
  50587=>"101101111",
  50588=>"110001010",
  50589=>"101111010",
  50590=>"111110011",
  50591=>"101001100",
  50592=>"101110111",
  50593=>"000010001",
  50594=>"000101011",
  50595=>"011010000",
  50596=>"011101001",
  50597=>"110010111",
  50598=>"001000011",
  50599=>"010000000",
  50600=>"011100110",
  50601=>"010000001",
  50602=>"110010100",
  50603=>"000101000",
  50604=>"001111101",
  50605=>"110001110",
  50606=>"101011110",
  50607=>"010001010",
  50608=>"101000110",
  50609=>"001000001",
  50610=>"100010000",
  50611=>"010101011",
  50612=>"101101111",
  50613=>"111110010",
  50614=>"001101001",
  50615=>"101111010",
  50616=>"011011010",
  50617=>"110000001",
  50618=>"101100010",
  50619=>"000001010",
  50620=>"110001000",
  50621=>"111010010",
  50622=>"010001000",
  50623=>"001100111",
  50624=>"010100011",
  50625=>"010100100",
  50626=>"111111000",
  50627=>"111101110",
  50628=>"001111001",
  50629=>"000011110",
  50630=>"110011111",
  50631=>"101110111",
  50632=>"010010000",
  50633=>"111111111",
  50634=>"111100001",
  50635=>"110101100",
  50636=>"101111100",
  50637=>"110100111",
  50638=>"001000000",
  50639=>"101010111",
  50640=>"010111110",
  50641=>"110010111",
  50642=>"000011101",
  50643=>"110110000",
  50644=>"100011001",
  50645=>"101101001",
  50646=>"111001101",
  50647=>"000000000",
  50648=>"000101110",
  50649=>"101011001",
  50650=>"101100110",
  50651=>"110011111",
  50652=>"101011010",
  50653=>"001010000",
  50654=>"011011110",
  50655=>"100000001",
  50656=>"101011011",
  50657=>"010110101",
  50658=>"011101111",
  50659=>"010100110",
  50660=>"101101101",
  50661=>"011111001",
  50662=>"001100101",
  50663=>"000011001",
  50664=>"101000000",
  50665=>"001010110",
  50666=>"111110100",
  50667=>"001001000",
  50668=>"000111101",
  50669=>"110011001",
  50670=>"000001010",
  50671=>"010001101",
  50672=>"011000101",
  50673=>"010010001",
  50674=>"100001011",
  50675=>"011101001",
  50676=>"100100110",
  50677=>"001101101",
  50678=>"000001000",
  50679=>"110110011",
  50680=>"011000000",
  50681=>"011000111",
  50682=>"110111011",
  50683=>"110101011",
  50684=>"111010001",
  50685=>"000111111",
  50686=>"100001111",
  50687=>"111010110",
  50688=>"010101110",
  50689=>"111010000",
  50690=>"010011110",
  50691=>"000010000",
  50692=>"111100111",
  50693=>"100000010",
  50694=>"010101011",
  50695=>"110001101",
  50696=>"011011000",
  50697=>"011110010",
  50698=>"100001100",
  50699=>"000000100",
  50700=>"100111111",
  50701=>"011111010",
  50702=>"111011101",
  50703=>"100011011",
  50704=>"010011110",
  50705=>"010010010",
  50706=>"000000001",
  50707=>"110101001",
  50708=>"010001011",
  50709=>"010011000",
  50710=>"000100000",
  50711=>"001100011",
  50712=>"011101000",
  50713=>"101101000",
  50714=>"010110011",
  50715=>"101000011",
  50716=>"010110010",
  50717=>"011110100",
  50718=>"011110010",
  50719=>"110110101",
  50720=>"111000111",
  50721=>"000001000",
  50722=>"010010101",
  50723=>"110010010",
  50724=>"111000111",
  50725=>"011110000",
  50726=>"100111011",
  50727=>"011101111",
  50728=>"101001001",
  50729=>"110110100",
  50730=>"101011001",
  50731=>"110001010",
  50732=>"100010011",
  50733=>"110100100",
  50734=>"100011110",
  50735=>"010110010",
  50736=>"000001000",
  50737=>"110100111",
  50738=>"111001110",
  50739=>"010101111",
  50740=>"011001000",
  50741=>"100101110",
  50742=>"001111100",
  50743=>"100110011",
  50744=>"011001010",
  50745=>"111110001",
  50746=>"100000111",
  50747=>"101111011",
  50748=>"000011001",
  50749=>"000000000",
  50750=>"100110100",
  50751=>"010101000",
  50752=>"001100010",
  50753=>"001101011",
  50754=>"010111011",
  50755=>"100001001",
  50756=>"100011111",
  50757=>"111101110",
  50758=>"110110001",
  50759=>"000110010",
  50760=>"110111000",
  50761=>"101011011",
  50762=>"100100111",
  50763=>"011110101",
  50764=>"010000010",
  50765=>"000100010",
  50766=>"001001111",
  50767=>"101110101",
  50768=>"011010010",
  50769=>"010010001",
  50770=>"011110101",
  50771=>"000001111",
  50772=>"010000001",
  50773=>"110101101",
  50774=>"110101100",
  50775=>"101100110",
  50776=>"101101001",
  50777=>"010111000",
  50778=>"100101010",
  50779=>"111011010",
  50780=>"010010001",
  50781=>"010011101",
  50782=>"010010000",
  50783=>"011010000",
  50784=>"101000011",
  50785=>"011101000",
  50786=>"111011100",
  50787=>"010001100",
  50788=>"110011010",
  50789=>"101001010",
  50790=>"101000110",
  50791=>"000100101",
  50792=>"111110001",
  50793=>"110000101",
  50794=>"111100010",
  50795=>"010010101",
  50796=>"011110100",
  50797=>"111011010",
  50798=>"101111010",
  50799=>"111011000",
  50800=>"100000100",
  50801=>"010110101",
  50802=>"000111101",
  50803=>"011000100",
  50804=>"001111100",
  50805=>"110111111",
  50806=>"101000011",
  50807=>"001011000",
  50808=>"101110100",
  50809=>"001001010",
  50810=>"001010000",
  50811=>"000100010",
  50812=>"111100000",
  50813=>"000010001",
  50814=>"000101110",
  50815=>"001111101",
  50816=>"110110100",
  50817=>"001011011",
  50818=>"011001010",
  50819=>"101010110",
  50820=>"110111010",
  50821=>"100101011",
  50822=>"011110001",
  50823=>"001110010",
  50824=>"110110111",
  50825=>"001011000",
  50826=>"111010001",
  50827=>"000110100",
  50828=>"000010000",
  50829=>"111111011",
  50830=>"000110010",
  50831=>"110111100",
  50832=>"001000000",
  50833=>"000011001",
  50834=>"110101001",
  50835=>"101010100",
  50836=>"101010000",
  50837=>"010101110",
  50838=>"000001000",
  50839=>"000101000",
  50840=>"000110100",
  50841=>"110100011",
  50842=>"110010100",
  50843=>"010111000",
  50844=>"001111110",
  50845=>"111011000",
  50846=>"011101010",
  50847=>"001011001",
  50848=>"101110110",
  50849=>"010110110",
  50850=>"010011010",
  50851=>"011101000",
  50852=>"101001001",
  50853=>"010101101",
  50854=>"010111110",
  50855=>"101101101",
  50856=>"010111101",
  50857=>"010001011",
  50858=>"110001101",
  50859=>"001010000",
  50860=>"010100001",
  50861=>"010010110",
  50862=>"000000001",
  50863=>"011011101",
  50864=>"000101001",
  50865=>"101101010",
  50866=>"011100110",
  50867=>"111011110",
  50868=>"111000110",
  50869=>"110011110",
  50870=>"011101010",
  50871=>"000100110",
  50872=>"111001001",
  50873=>"001010000",
  50874=>"110011011",
  50875=>"000001000",
  50876=>"010111000",
  50877=>"000001001",
  50878=>"110110101",
  50879=>"110110011",
  50880=>"100011010",
  50881=>"111110101",
  50882=>"010110001",
  50883=>"001001010",
  50884=>"010011001",
  50885=>"111111110",
  50886=>"011110110",
  50887=>"000101101",
  50888=>"110000000",
  50889=>"100001001",
  50890=>"011101110",
  50891=>"110010101",
  50892=>"001101001",
  50893=>"111101011",
  50894=>"011001001",
  50895=>"101011001",
  50896=>"000110100",
  50897=>"101101011",
  50898=>"000111000",
  50899=>"011011001",
  50900=>"100111111",
  50901=>"011001110",
  50902=>"101000101",
  50903=>"000010010",
  50904=>"000000011",
  50905=>"111001100",
  50906=>"001111010",
  50907=>"011101111",
  50908=>"000010110",
  50909=>"110100001",
  50910=>"101010001",
  50911=>"111101101",
  50912=>"011011101",
  50913=>"001011100",
  50914=>"101011001",
  50915=>"101001111",
  50916=>"100010100",
  50917=>"100100110",
  50918=>"010110010",
  50919=>"110100110",
  50920=>"000010101",
  50921=>"000000011",
  50922=>"001001001",
  50923=>"010100110",
  50924=>"010110001",
  50925=>"101001000",
  50926=>"110110100",
  50927=>"100101111",
  50928=>"011100110",
  50929=>"010101111",
  50930=>"110000101",
  50931=>"000000100",
  50932=>"110000100",
  50933=>"110010001",
  50934=>"110001100",
  50935=>"111111101",
  50936=>"011101001",
  50937=>"111000111",
  50938=>"010010100",
  50939=>"000000010",
  50940=>"100110000",
  50941=>"111100101",
  50942=>"100000001",
  50943=>"001101010",
  50944=>"111011011",
  50945=>"110110110",
  50946=>"000110001",
  50947=>"011100100",
  50948=>"010100110",
  50949=>"000101100",
  50950=>"011001101",
  50951=>"010011100",
  50952=>"000111000",
  50953=>"111011001",
  50954=>"110101100",
  50955=>"101010011",
  50956=>"010011001",
  50957=>"111101101",
  50958=>"100011100",
  50959=>"010011000",
  50960=>"000001000",
  50961=>"000110010",
  50962=>"111010011",
  50963=>"000011101",
  50964=>"110100001",
  50965=>"101000110",
  50966=>"010110000",
  50967=>"101111110",
  50968=>"111110010",
  50969=>"110010011",
  50970=>"110001100",
  50971=>"100010111",
  50972=>"101011010",
  50973=>"000011101",
  50974=>"011101001",
  50975=>"111001001",
  50976=>"110000000",
  50977=>"000101000",
  50978=>"000010100",
  50979=>"111011011",
  50980=>"111111000",
  50981=>"110101111",
  50982=>"010111100",
  50983=>"110111001",
  50984=>"000100011",
  50985=>"100100101",
  50986=>"100011000",
  50987=>"011110100",
  50988=>"100001110",
  50989=>"010111010",
  50990=>"110010010",
  50991=>"000011100",
  50992=>"000001000",
  50993=>"100001011",
  50994=>"100110101",
  50995=>"010010110",
  50996=>"001101101",
  50997=>"101110011",
  50998=>"100111100",
  50999=>"110001011",
  51000=>"111100000",
  51001=>"111010111",
  51002=>"001000000",
  51003=>"110111010",
  51004=>"000001011",
  51005=>"000100110",
  51006=>"111100000",
  51007=>"101011110",
  51008=>"010100011",
  51009=>"100000101",
  51010=>"001100101",
  51011=>"000110110",
  51012=>"000111011",
  51013=>"011100110",
  51014=>"110111111",
  51015=>"000010100",
  51016=>"001111111",
  51017=>"111111011",
  51018=>"110101111",
  51019=>"011000011",
  51020=>"010000101",
  51021=>"111011111",
  51022=>"010111101",
  51023=>"101011111",
  51024=>"000111100",
  51025=>"011100010",
  51026=>"101101110",
  51027=>"000000000",
  51028=>"010000010",
  51029=>"100011111",
  51030=>"010111100",
  51031=>"010010000",
  51032=>"000100000",
  51033=>"111101011",
  51034=>"101100010",
  51035=>"010011011",
  51036=>"111110011",
  51037=>"110100011",
  51038=>"100110011",
  51039=>"000000010",
  51040=>"101000011",
  51041=>"100111111",
  51042=>"001101100",
  51043=>"110110100",
  51044=>"010000001",
  51045=>"001000100",
  51046=>"000110110",
  51047=>"001110111",
  51048=>"111101100",
  51049=>"110000101",
  51050=>"000101010",
  51051=>"111110101",
  51052=>"101111100",
  51053=>"110100011",
  51054=>"110100100",
  51055=>"010110100",
  51056=>"010010100",
  51057=>"011101011",
  51058=>"101001111",
  51059=>"100110001",
  51060=>"010000001",
  51061=>"100010000",
  51062=>"110101100",
  51063=>"100100000",
  51064=>"011011001",
  51065=>"100001011",
  51066=>"011000100",
  51067=>"011100001",
  51068=>"000000000",
  51069=>"100100110",
  51070=>"110111111",
  51071=>"010001000",
  51072=>"001001010",
  51073=>"001000000",
  51074=>"010110101",
  51075=>"000011010",
  51076=>"000001101",
  51077=>"111001110",
  51078=>"000111000",
  51079=>"100110111",
  51080=>"110011011",
  51081=>"100001100",
  51082=>"101100001",
  51083=>"011000011",
  51084=>"100110001",
  51085=>"011110001",
  51086=>"010001100",
  51087=>"001101101",
  51088=>"101011100",
  51089=>"111000001",
  51090=>"100000000",
  51091=>"011010101",
  51092=>"111011101",
  51093=>"110001010",
  51094=>"000010110",
  51095=>"010100110",
  51096=>"000100000",
  51097=>"000110010",
  51098=>"010010010",
  51099=>"010100001",
  51100=>"001110010",
  51101=>"110000001",
  51102=>"101101001",
  51103=>"100010010",
  51104=>"010101101",
  51105=>"110111110",
  51106=>"000010010",
  51107=>"101000001",
  51108=>"001110010",
  51109=>"100010000",
  51110=>"111111110",
  51111=>"111011010",
  51112=>"000101101",
  51113=>"000010011",
  51114=>"000110000",
  51115=>"100010100",
  51116=>"001000110",
  51117=>"111000010",
  51118=>"110011000",
  51119=>"011010111",
  51120=>"110000010",
  51121=>"000000101",
  51122=>"010100001",
  51123=>"101000101",
  51124=>"100000001",
  51125=>"110111111",
  51126=>"110110010",
  51127=>"100010101",
  51128=>"110101111",
  51129=>"011011001",
  51130=>"011101101",
  51131=>"011111000",
  51132=>"110101010",
  51133=>"100101010",
  51134=>"010110111",
  51135=>"010010110",
  51136=>"000100011",
  51137=>"000000000",
  51138=>"101111100",
  51139=>"110000010",
  51140=>"011001100",
  51141=>"111100101",
  51142=>"010101110",
  51143=>"001111011",
  51144=>"101001000",
  51145=>"010001010",
  51146=>"010000011",
  51147=>"011101110",
  51148=>"000100010",
  51149=>"010100100",
  51150=>"111110001",
  51151=>"001011110",
  51152=>"010011101",
  51153=>"100110111",
  51154=>"110101101",
  51155=>"100000010",
  51156=>"001001111",
  51157=>"100000100",
  51158=>"101011110",
  51159=>"001000000",
  51160=>"110000111",
  51161=>"100100011",
  51162=>"001111000",
  51163=>"100000111",
  51164=>"010101101",
  51165=>"010110101",
  51166=>"110111001",
  51167=>"111010110",
  51168=>"011010000",
  51169=>"000010110",
  51170=>"010001111",
  51171=>"100010101",
  51172=>"001011000",
  51173=>"111111011",
  51174=>"000101011",
  51175=>"010010110",
  51176=>"101000000",
  51177=>"111110011",
  51178=>"110111001",
  51179=>"001100101",
  51180=>"010101011",
  51181=>"011111110",
  51182=>"111000100",
  51183=>"010101111",
  51184=>"111010000",
  51185=>"101011101",
  51186=>"101101011",
  51187=>"110100010",
  51188=>"111011111",
  51189=>"001001101",
  51190=>"101001100",
  51191=>"111011110",
  51192=>"000011110",
  51193=>"110101110",
  51194=>"010001000",
  51195=>"011111111",
  51196=>"101100011",
  51197=>"010011010",
  51198=>"100000101",
  51199=>"010011111",
  51200=>"011110101",
  51201=>"101101000",
  51202=>"100010111",
  51203=>"010000010",
  51204=>"001001000",
  51205=>"011111101",
  51206=>"010000000",
  51207=>"000110001",
  51208=>"011011001",
  51209=>"000100000",
  51210=>"101001011",
  51211=>"111010100",
  51212=>"100100001",
  51213=>"010010111",
  51214=>"001011000",
  51215=>"111101101",
  51216=>"111111001",
  51217=>"011001101",
  51218=>"110101001",
  51219=>"010111110",
  51220=>"010000101",
  51221=>"011011011",
  51222=>"100101110",
  51223=>"000111011",
  51224=>"001011000",
  51225=>"100100111",
  51226=>"100011101",
  51227=>"011101101",
  51228=>"100010000",
  51229=>"000100010",
  51230=>"011100011",
  51231=>"111001001",
  51232=>"100010010",
  51233=>"101101101",
  51234=>"111010000",
  51235=>"111100100",
  51236=>"111101100",
  51237=>"000001111",
  51238=>"011110001",
  51239=>"011011001",
  51240=>"100111000",
  51241=>"100000001",
  51242=>"100010000",
  51243=>"100100110",
  51244=>"101111100",
  51245=>"010101010",
  51246=>"110010010",
  51247=>"100001110",
  51248=>"111011111",
  51249=>"110110011",
  51250=>"100001101",
  51251=>"011011010",
  51252=>"110000111",
  51253=>"000010110",
  51254=>"110110100",
  51255=>"010101101",
  51256=>"011101111",
  51257=>"011110000",
  51258=>"001100111",
  51259=>"110001010",
  51260=>"010111101",
  51261=>"101101111",
  51262=>"110000000",
  51263=>"011010010",
  51264=>"010111111",
  51265=>"011110100",
  51266=>"100100111",
  51267=>"100010101",
  51268=>"000010010",
  51269=>"000100011",
  51270=>"011010001",
  51271=>"101101110",
  51272=>"011000000",
  51273=>"100101000",
  51274=>"111010001",
  51275=>"100010010",
  51276=>"001010011",
  51277=>"010100010",
  51278=>"101011000",
  51279=>"100101110",
  51280=>"001001010",
  51281=>"000110010",
  51282=>"000110111",
  51283=>"011101110",
  51284=>"001110011",
  51285=>"011101001",
  51286=>"001010111",
  51287=>"101101001",
  51288=>"100010000",
  51289=>"010111100",
  51290=>"001110111",
  51291=>"101010101",
  51292=>"010111111",
  51293=>"001101101",
  51294=>"111011001",
  51295=>"001000010",
  51296=>"011001011",
  51297=>"000001101",
  51298=>"101110100",
  51299=>"110010100",
  51300=>"001000000",
  51301=>"111000010",
  51302=>"010101100",
  51303=>"000011000",
  51304=>"000111010",
  51305=>"000001111",
  51306=>"010010110",
  51307=>"110001010",
  51308=>"110001001",
  51309=>"110111001",
  51310=>"001110000",
  51311=>"100001101",
  51312=>"000100011",
  51313=>"000111000",
  51314=>"111001001",
  51315=>"010011011",
  51316=>"010011000",
  51317=>"011111111",
  51318=>"001001101",
  51319=>"110011101",
  51320=>"111000000",
  51321=>"011001110",
  51322=>"111111111",
  51323=>"010000101",
  51324=>"010101010",
  51325=>"010000101",
  51326=>"011101010",
  51327=>"011111111",
  51328=>"110101110",
  51329=>"110110110",
  51330=>"000001001",
  51331=>"110010010",
  51332=>"010111000",
  51333=>"000110111",
  51334=>"001101111",
  51335=>"100000101",
  51336=>"001100010",
  51337=>"000000001",
  51338=>"110011000",
  51339=>"000001101",
  51340=>"000011100",
  51341=>"100000100",
  51342=>"011000101",
  51343=>"000010000",
  51344=>"011001001",
  51345=>"000101011",
  51346=>"100110111",
  51347=>"010111110",
  51348=>"101111101",
  51349=>"001010011",
  51350=>"001000100",
  51351=>"000000101",
  51352=>"011010110",
  51353=>"011011101",
  51354=>"011111111",
  51355=>"010101000",
  51356=>"000110010",
  51357=>"111111101",
  51358=>"100000110",
  51359=>"001101100",
  51360=>"101101000",
  51361=>"100100011",
  51362=>"000110110",
  51363=>"010001011",
  51364=>"001101110",
  51365=>"011000000",
  51366=>"011100011",
  51367=>"100101001",
  51368=>"000000011",
  51369=>"011000001",
  51370=>"010110101",
  51371=>"000000110",
  51372=>"110001111",
  51373=>"001000101",
  51374=>"010001010",
  51375=>"001101110",
  51376=>"111101000",
  51377=>"111001000",
  51378=>"111111111",
  51379=>"101110010",
  51380=>"001101001",
  51381=>"010011101",
  51382=>"000010100",
  51383=>"011000110",
  51384=>"001000001",
  51385=>"110001011",
  51386=>"110110110",
  51387=>"111111111",
  51388=>"101111001",
  51389=>"010000100",
  51390=>"101101100",
  51391=>"111011001",
  51392=>"010100111",
  51393=>"001010001",
  51394=>"011111011",
  51395=>"011001010",
  51396=>"111000011",
  51397=>"010010101",
  51398=>"110101101",
  51399=>"101001011",
  51400=>"011110010",
  51401=>"011100010",
  51402=>"011110110",
  51403=>"110011111",
  51404=>"010001101",
  51405=>"011110011",
  51406=>"001110100",
  51407=>"110010000",
  51408=>"101100100",
  51409=>"001010000",
  51410=>"101110110",
  51411=>"001101010",
  51412=>"010111001",
  51413=>"101110111",
  51414=>"101001100",
  51415=>"101011000",
  51416=>"000100000",
  51417=>"101000011",
  51418=>"011011011",
  51419=>"101000110",
  51420=>"100001110",
  51421=>"110100100",
  51422=>"110010110",
  51423=>"000001100",
  51424=>"101101111",
  51425=>"100100101",
  51426=>"001100011",
  51427=>"101100100",
  51428=>"110001110",
  51429=>"011011010",
  51430=>"011100101",
  51431=>"100011100",
  51432=>"001101000",
  51433=>"100011000",
  51434=>"000001000",
  51435=>"111001011",
  51436=>"110110100",
  51437=>"101111001",
  51438=>"010110000",
  51439=>"100100111",
  51440=>"010001100",
  51441=>"000010000",
  51442=>"010111111",
  51443=>"101100011",
  51444=>"100001100",
  51445=>"010001011",
  51446=>"110110111",
  51447=>"000000000",
  51448=>"000101111",
  51449=>"111010001",
  51450=>"000111110",
  51451=>"101001010",
  51452=>"000010111",
  51453=>"110101110",
  51454=>"111111010",
  51455=>"110111011",
  51456=>"010010100",
  51457=>"010010000",
  51458=>"011000011",
  51459=>"111000001",
  51460=>"111101100",
  51461=>"000010001",
  51462=>"100100011",
  51463=>"101111110",
  51464=>"111100110",
  51465=>"000001111",
  51466=>"000111101",
  51467=>"110100100",
  51468=>"010000111",
  51469=>"100101010",
  51470=>"110110101",
  51471=>"110011000",
  51472=>"110001100",
  51473=>"101100011",
  51474=>"110010001",
  51475=>"010001111",
  51476=>"001101111",
  51477=>"001011010",
  51478=>"000001000",
  51479=>"100111101",
  51480=>"001111011",
  51481=>"010101101",
  51482=>"111001000",
  51483=>"011010011",
  51484=>"010110011",
  51485=>"101100001",
  51486=>"110001011",
  51487=>"111001011",
  51488=>"010011000",
  51489=>"011010001",
  51490=>"010000010",
  51491=>"111001001",
  51492=>"000010101",
  51493=>"011110101",
  51494=>"101000000",
  51495=>"011100111",
  51496=>"101100110",
  51497=>"011111010",
  51498=>"100000111",
  51499=>"111110101",
  51500=>"010100011",
  51501=>"001001101",
  51502=>"011110101",
  51503=>"111011111",
  51504=>"111100000",
  51505=>"000010101",
  51506=>"010110110",
  51507=>"111100001",
  51508=>"100111000",
  51509=>"110101101",
  51510=>"011010001",
  51511=>"011000001",
  51512=>"010000010",
  51513=>"110000011",
  51514=>"111001101",
  51515=>"100110101",
  51516=>"101010000",
  51517=>"010001001",
  51518=>"101110110",
  51519=>"110111111",
  51520=>"011101100",
  51521=>"000111010",
  51522=>"100101111",
  51523=>"011101101",
  51524=>"110101001",
  51525=>"111000011",
  51526=>"110000100",
  51527=>"101011111",
  51528=>"010101100",
  51529=>"100101000",
  51530=>"000011101",
  51531=>"110111100",
  51532=>"101100010",
  51533=>"001010101",
  51534=>"111001101",
  51535=>"000110010",
  51536=>"000100010",
  51537=>"000000000",
  51538=>"110001100",
  51539=>"100000011",
  51540=>"110110010",
  51541=>"001110011",
  51542=>"001000001",
  51543=>"001101101",
  51544=>"001111011",
  51545=>"010100110",
  51546=>"011100001",
  51547=>"010101011",
  51548=>"000000000",
  51549=>"101001011",
  51550=>"001101001",
  51551=>"011100101",
  51552=>"101000100",
  51553=>"000010110",
  51554=>"000010000",
  51555=>"101001001",
  51556=>"000111001",
  51557=>"010001110",
  51558=>"111000100",
  51559=>"111110100",
  51560=>"110010100",
  51561=>"110010100",
  51562=>"011110100",
  51563=>"101110100",
  51564=>"001000101",
  51565=>"111111110",
  51566=>"000010100",
  51567=>"001011100",
  51568=>"010100101",
  51569=>"001101101",
  51570=>"000101010",
  51571=>"010010100",
  51572=>"101001000",
  51573=>"011101011",
  51574=>"100000111",
  51575=>"100011110",
  51576=>"110100010",
  51577=>"110110010",
  51578=>"011000001",
  51579=>"101011011",
  51580=>"000111110",
  51581=>"100011110",
  51582=>"000001100",
  51583=>"000100100",
  51584=>"111001101",
  51585=>"000101111",
  51586=>"001101101",
  51587=>"010010000",
  51588=>"111001111",
  51589=>"001111001",
  51590=>"000100000",
  51591=>"010100000",
  51592=>"111010010",
  51593=>"000001101",
  51594=>"010001000",
  51595=>"010100110",
  51596=>"011001110",
  51597=>"111110010",
  51598=>"101000101",
  51599=>"001000011",
  51600=>"011100010",
  51601=>"000101010",
  51602=>"011100001",
  51603=>"011100110",
  51604=>"000110101",
  51605=>"011010011",
  51606=>"100100100",
  51607=>"110000011",
  51608=>"001100110",
  51609=>"011101100",
  51610=>"111001011",
  51611=>"010100110",
  51612=>"000000100",
  51613=>"101110011",
  51614=>"100001001",
  51615=>"111010100",
  51616=>"100100010",
  51617=>"000010001",
  51618=>"000001101",
  51619=>"010001111",
  51620=>"001011111",
  51621=>"101100100",
  51622=>"111110000",
  51623=>"010010101",
  51624=>"111011001",
  51625=>"000101110",
  51626=>"100101001",
  51627=>"001011100",
  51628=>"111110100",
  51629=>"110110010",
  51630=>"010100000",
  51631=>"001110001",
  51632=>"101101110",
  51633=>"100000000",
  51634=>"010001010",
  51635=>"001101100",
  51636=>"100100101",
  51637=>"011011101",
  51638=>"101101000",
  51639=>"001101111",
  51640=>"101001011",
  51641=>"111000110",
  51642=>"001100010",
  51643=>"100001010",
  51644=>"110101011",
  51645=>"111101110",
  51646=>"100110111",
  51647=>"001100110",
  51648=>"001110111",
  51649=>"000100110",
  51650=>"000010001",
  51651=>"110011110",
  51652=>"100111101",
  51653=>"011001000",
  51654=>"111010111",
  51655=>"011111110",
  51656=>"010110101",
  51657=>"111001101",
  51658=>"100000000",
  51659=>"110100000",
  51660=>"010101100",
  51661=>"101101111",
  51662=>"111011101",
  51663=>"110011110",
  51664=>"000011101",
  51665=>"111001000",
  51666=>"110111111",
  51667=>"100111010",
  51668=>"111111001",
  51669=>"101000000",
  51670=>"011010001",
  51671=>"111111100",
  51672=>"100001011",
  51673=>"101101101",
  51674=>"011100011",
  51675=>"111100010",
  51676=>"100010011",
  51677=>"101000001",
  51678=>"010101000",
  51679=>"000100111",
  51680=>"110011100",
  51681=>"000111101",
  51682=>"011100111",
  51683=>"110011101",
  51684=>"111101100",
  51685=>"100011101",
  51686=>"111111110",
  51687=>"110100110",
  51688=>"110101101",
  51689=>"101101010",
  51690=>"011101100",
  51691=>"111000100",
  51692=>"100010000",
  51693=>"001110101",
  51694=>"000100011",
  51695=>"001010000",
  51696=>"100101010",
  51697=>"001010000",
  51698=>"111000010",
  51699=>"011001101",
  51700=>"011110110",
  51701=>"100010010",
  51702=>"001111000",
  51703=>"010001111",
  51704=>"111101001",
  51705=>"111101110",
  51706=>"101100011",
  51707=>"001100001",
  51708=>"000011111",
  51709=>"101110000",
  51710=>"101010010",
  51711=>"000101110",
  51712=>"100110011",
  51713=>"000110111",
  51714=>"110010011",
  51715=>"010001000",
  51716=>"111101001",
  51717=>"010111011",
  51718=>"101111101",
  51719=>"010110000",
  51720=>"001010010",
  51721=>"000011100",
  51722=>"000111000",
  51723=>"010000100",
  51724=>"011111111",
  51725=>"010000000",
  51726=>"101111101",
  51727=>"110001110",
  51728=>"100110110",
  51729=>"000011111",
  51730=>"001001001",
  51731=>"100001111",
  51732=>"101000111",
  51733=>"001010100",
  51734=>"000100011",
  51735=>"000001010",
  51736=>"101011101",
  51737=>"011000100",
  51738=>"101000100",
  51739=>"011000100",
  51740=>"110110011",
  51741=>"011010011",
  51742=>"000101110",
  51743=>"000011100",
  51744=>"000110100",
  51745=>"001010010",
  51746=>"000000010",
  51747=>"001000001",
  51748=>"011011000",
  51749=>"001100100",
  51750=>"010001000",
  51751=>"000001001",
  51752=>"111100111",
  51753=>"010100111",
  51754=>"110000001",
  51755=>"011100110",
  51756=>"010110100",
  51757=>"101011110",
  51758=>"001100000",
  51759=>"110111110",
  51760=>"101001011",
  51761=>"001001100",
  51762=>"110001011",
  51763=>"110011001",
  51764=>"000100010",
  51765=>"111010011",
  51766=>"001111001",
  51767=>"100101000",
  51768=>"110000011",
  51769=>"101001100",
  51770=>"011100000",
  51771=>"001110100",
  51772=>"000010001",
  51773=>"100001000",
  51774=>"001100110",
  51775=>"100010100",
  51776=>"011101010",
  51777=>"000100101",
  51778=>"110101111",
  51779=>"001100101",
  51780=>"011001100",
  51781=>"000001010",
  51782=>"100111110",
  51783=>"001100111",
  51784=>"111100100",
  51785=>"111010001",
  51786=>"110010111",
  51787=>"101001001",
  51788=>"011010110",
  51789=>"010111000",
  51790=>"111110001",
  51791=>"101000000",
  51792=>"111111111",
  51793=>"011011000",
  51794=>"111001110",
  51795=>"000110111",
  51796=>"100001010",
  51797=>"101000100",
  51798=>"000011101",
  51799=>"101111100",
  51800=>"100011111",
  51801=>"111110100",
  51802=>"111011111",
  51803=>"111101111",
  51804=>"001000001",
  51805=>"000011011",
  51806=>"100111000",
  51807=>"011101100",
  51808=>"101111100",
  51809=>"111000000",
  51810=>"000010101",
  51811=>"011010000",
  51812=>"001110011",
  51813=>"111110001",
  51814=>"010100111",
  51815=>"000100110",
  51816=>"111011100",
  51817=>"000110110",
  51818=>"100010110",
  51819=>"100110101",
  51820=>"101000111",
  51821=>"110001011",
  51822=>"000010100",
  51823=>"100000100",
  51824=>"100101101",
  51825=>"001010000",
  51826=>"000010111",
  51827=>"110010000",
  51828=>"100110100",
  51829=>"100011110",
  51830=>"001100101",
  51831=>"100001110",
  51832=>"101100000",
  51833=>"110011011",
  51834=>"001000110",
  51835=>"001110010",
  51836=>"111111110",
  51837=>"000011001",
  51838=>"011011111",
  51839=>"000100110",
  51840=>"011100110",
  51841=>"010000010",
  51842=>"011101100",
  51843=>"011111000",
  51844=>"111111111",
  51845=>"000000111",
  51846=>"111100101",
  51847=>"001110000",
  51848=>"010110011",
  51849=>"010000000",
  51850=>"101110111",
  51851=>"011011010",
  51852=>"110001100",
  51853=>"011111110",
  51854=>"001000110",
  51855=>"101000001",
  51856=>"111001111",
  51857=>"000111101",
  51858=>"101011111",
  51859=>"000110100",
  51860=>"001010011",
  51861=>"100110010",
  51862=>"110110110",
  51863=>"100011001",
  51864=>"010000010",
  51865=>"100111110",
  51866=>"010010010",
  51867=>"011100111",
  51868=>"010000000",
  51869=>"100110111",
  51870=>"110010111",
  51871=>"001111011",
  51872=>"110010101",
  51873=>"110000110",
  51874=>"011111101",
  51875=>"000000110",
  51876=>"000111000",
  51877=>"100111110",
  51878=>"011100010",
  51879=>"110110010",
  51880=>"101010011",
  51881=>"011111011",
  51882=>"011110101",
  51883=>"001101111",
  51884=>"100101110",
  51885=>"101110000",
  51886=>"000011100",
  51887=>"011110100",
  51888=>"111110101",
  51889=>"000010110",
  51890=>"100110111",
  51891=>"110000101",
  51892=>"110001000",
  51893=>"101010010",
  51894=>"111000100",
  51895=>"100110100",
  51896=>"011110011",
  51897=>"101110001",
  51898=>"010110000",
  51899=>"000111101",
  51900=>"110100111",
  51901=>"101001100",
  51902=>"001001100",
  51903=>"010010110",
  51904=>"100100111",
  51905=>"110111101",
  51906=>"101011101",
  51907=>"010110111",
  51908=>"100111111",
  51909=>"001011111",
  51910=>"100000111",
  51911=>"010111100",
  51912=>"010100100",
  51913=>"100111101",
  51914=>"110101110",
  51915=>"101010011",
  51916=>"111101011",
  51917=>"100000110",
  51918=>"011000100",
  51919=>"011000011",
  51920=>"101111110",
  51921=>"100101100",
  51922=>"010011001",
  51923=>"001001001",
  51924=>"011110110",
  51925=>"110100011",
  51926=>"110111110",
  51927=>"100010010",
  51928=>"000001110",
  51929=>"011011111",
  51930=>"010001111",
  51931=>"111101000",
  51932=>"001101100",
  51933=>"011001001",
  51934=>"000101001",
  51935=>"010000000",
  51936=>"100110100",
  51937=>"001011011",
  51938=>"000001111",
  51939=>"011011010",
  51940=>"110001111",
  51941=>"110100101",
  51942=>"001001100",
  51943=>"111110010",
  51944=>"010100010",
  51945=>"111111000",
  51946=>"010000101",
  51947=>"111111100",
  51948=>"100011011",
  51949=>"001001010",
  51950=>"110111011",
  51951=>"100001000",
  51952=>"111011010",
  51953=>"100111001",
  51954=>"000101101",
  51955=>"001000011",
  51956=>"111011001",
  51957=>"011100111",
  51958=>"011111111",
  51959=>"011110010",
  51960=>"011110100",
  51961=>"110001110",
  51962=>"001101101",
  51963=>"010001110",
  51964=>"011000010",
  51965=>"100000001",
  51966=>"111111001",
  51967=>"001000111",
  51968=>"010111000",
  51969=>"000000010",
  51970=>"010101111",
  51971=>"110010110",
  51972=>"000100011",
  51973=>"000000100",
  51974=>"011110110",
  51975=>"010100111",
  51976=>"011111100",
  51977=>"110100111",
  51978=>"111010000",
  51979=>"010011111",
  51980=>"100100010",
  51981=>"011011110",
  51982=>"001111111",
  51983=>"000011011",
  51984=>"011111010",
  51985=>"110110001",
  51986=>"110000000",
  51987=>"011100111",
  51988=>"001111101",
  51989=>"101001011",
  51990=>"100101101",
  51991=>"110101110",
  51992=>"011100111",
  51993=>"000001000",
  51994=>"010110010",
  51995=>"011100001",
  51996=>"011100000",
  51997=>"010011101",
  51998=>"100010010",
  51999=>"111010100",
  52000=>"110000000",
  52001=>"000101001",
  52002=>"000101110",
  52003=>"111001111",
  52004=>"100000000",
  52005=>"100000110",
  52006=>"111010011",
  52007=>"101011100",
  52008=>"110000111",
  52009=>"011000101",
  52010=>"011001111",
  52011=>"101100101",
  52012=>"011110000",
  52013=>"010000000",
  52014=>"100010000",
  52015=>"101101011",
  52016=>"000010001",
  52017=>"100100110",
  52018=>"001100010",
  52019=>"110011000",
  52020=>"010001110",
  52021=>"111000010",
  52022=>"011111101",
  52023=>"000111100",
  52024=>"000001001",
  52025=>"001000000",
  52026=>"000011000",
  52027=>"011001010",
  52028=>"011000111",
  52029=>"001111111",
  52030=>"101001100",
  52031=>"111011101",
  52032=>"111100111",
  52033=>"111011111",
  52034=>"110101101",
  52035=>"000000010",
  52036=>"000001100",
  52037=>"000011111",
  52038=>"100000100",
  52039=>"010001101",
  52040=>"011100111",
  52041=>"001011111",
  52042=>"001101011",
  52043=>"100111101",
  52044=>"100100110",
  52045=>"001000010",
  52046=>"010111000",
  52047=>"101111000",
  52048=>"100101011",
  52049=>"001100001",
  52050=>"100000110",
  52051=>"111101001",
  52052=>"000000001",
  52053=>"001000101",
  52054=>"111101000",
  52055=>"010101011",
  52056=>"111101111",
  52057=>"101011111",
  52058=>"100101110",
  52059=>"000011100",
  52060=>"101001011",
  52061=>"010000000",
  52062=>"000001111",
  52063=>"100111100",
  52064=>"011010011",
  52065=>"100110001",
  52066=>"110100000",
  52067=>"010000011",
  52068=>"101010011",
  52069=>"110000001",
  52070=>"111101000",
  52071=>"010000000",
  52072=>"010001000",
  52073=>"110000100",
  52074=>"110011011",
  52075=>"001110010",
  52076=>"101010101",
  52077=>"101010101",
  52078=>"001111000",
  52079=>"100001101",
  52080=>"101101011",
  52081=>"011000001",
  52082=>"110011110",
  52083=>"100001001",
  52084=>"000000010",
  52085=>"010010011",
  52086=>"101110101",
  52087=>"011010011",
  52088=>"001100000",
  52089=>"011001101",
  52090=>"110101001",
  52091=>"011110101",
  52092=>"100011011",
  52093=>"100100100",
  52094=>"100011111",
  52095=>"100101100",
  52096=>"010011000",
  52097=>"000011110",
  52098=>"001101110",
  52099=>"101100110",
  52100=>"011001001",
  52101=>"101001101",
  52102=>"111110001",
  52103=>"010100111",
  52104=>"110000101",
  52105=>"000010111",
  52106=>"100001000",
  52107=>"100111011",
  52108=>"110110011",
  52109=>"111111100",
  52110=>"110111011",
  52111=>"101010110",
  52112=>"100101001",
  52113=>"010000101",
  52114=>"101011001",
  52115=>"010011100",
  52116=>"010000000",
  52117=>"101000010",
  52118=>"011101110",
  52119=>"111101101",
  52120=>"000000010",
  52121=>"010000011",
  52122=>"101110110",
  52123=>"110001001",
  52124=>"101000000",
  52125=>"100011111",
  52126=>"100101110",
  52127=>"100101010",
  52128=>"100000000",
  52129=>"001111011",
  52130=>"111001010",
  52131=>"001010100",
  52132=>"001111101",
  52133=>"111100000",
  52134=>"110100100",
  52135=>"111001101",
  52136=>"111111001",
  52137=>"001101001",
  52138=>"110010110",
  52139=>"110100111",
  52140=>"101001000",
  52141=>"100101110",
  52142=>"110111000",
  52143=>"000100001",
  52144=>"011110100",
  52145=>"110011110",
  52146=>"110101001",
  52147=>"010101100",
  52148=>"110001010",
  52149=>"000010111",
  52150=>"111001000",
  52151=>"010000011",
  52152=>"001101011",
  52153=>"000100010",
  52154=>"001001010",
  52155=>"011110010",
  52156=>"001101000",
  52157=>"110011111",
  52158=>"110111111",
  52159=>"101101111",
  52160=>"110111110",
  52161=>"001111111",
  52162=>"000011111",
  52163=>"000010101",
  52164=>"000000000",
  52165=>"010100010",
  52166=>"111000011",
  52167=>"111111111",
  52168=>"000100101",
  52169=>"000010010",
  52170=>"000010001",
  52171=>"011000001",
  52172=>"011101000",
  52173=>"110110000",
  52174=>"110010001",
  52175=>"001111011",
  52176=>"010011011",
  52177=>"111001101",
  52178=>"001010011",
  52179=>"010110101",
  52180=>"010000010",
  52181=>"111010010",
  52182=>"011011000",
  52183=>"111101101",
  52184=>"000000111",
  52185=>"010010110",
  52186=>"001111101",
  52187=>"000000111",
  52188=>"100110111",
  52189=>"100110101",
  52190=>"110010101",
  52191=>"110001000",
  52192=>"111010011",
  52193=>"110001101",
  52194=>"011010001",
  52195=>"011001000",
  52196=>"011100100",
  52197=>"111000100",
  52198=>"000101111",
  52199=>"010010001",
  52200=>"101010110",
  52201=>"010010111",
  52202=>"000010110",
  52203=>"101110111",
  52204=>"011101010",
  52205=>"001010000",
  52206=>"101111101",
  52207=>"101110000",
  52208=>"011110010",
  52209=>"100001000",
  52210=>"110100011",
  52211=>"100000011",
  52212=>"000111000",
  52213=>"000001010",
  52214=>"101100000",
  52215=>"010001111",
  52216=>"101101111",
  52217=>"111110100",
  52218=>"110000100",
  52219=>"111010110",
  52220=>"010000110",
  52221=>"111000110",
  52222=>"110100100",
  52223=>"110001000",
  52224=>"101100000",
  52225=>"011010100",
  52226=>"000101101",
  52227=>"100101101",
  52228=>"000100010",
  52229=>"110110101",
  52230=>"001001111",
  52231=>"111111000",
  52232=>"110011011",
  52233=>"110001001",
  52234=>"101010001",
  52235=>"010100101",
  52236=>"111000010",
  52237=>"000111111",
  52238=>"111101010",
  52239=>"100100111",
  52240=>"000100100",
  52241=>"011011111",
  52242=>"111110111",
  52243=>"100001100",
  52244=>"010100101",
  52245=>"010110101",
  52246=>"111101011",
  52247=>"001010000",
  52248=>"001001100",
  52249=>"110111000",
  52250=>"011110110",
  52251=>"001111111",
  52252=>"111101001",
  52253=>"011010011",
  52254=>"100111100",
  52255=>"101100101",
  52256=>"111010100",
  52257=>"000000110",
  52258=>"001011110",
  52259=>"111000100",
  52260=>"000011011",
  52261=>"001001001",
  52262=>"000011110",
  52263=>"011001001",
  52264=>"001101010",
  52265=>"000100001",
  52266=>"011011011",
  52267=>"001100001",
  52268=>"011001100",
  52269=>"011110101",
  52270=>"001000001",
  52271=>"000001110",
  52272=>"111011111",
  52273=>"000010111",
  52274=>"011100110",
  52275=>"110111010",
  52276=>"001001000",
  52277=>"000000001",
  52278=>"011110111",
  52279=>"000001101",
  52280=>"110001000",
  52281=>"100000110",
  52282=>"101001100",
  52283=>"000010010",
  52284=>"000111001",
  52285=>"001001000",
  52286=>"101000101",
  52287=>"000101011",
  52288=>"101111011",
  52289=>"000000000",
  52290=>"011000000",
  52291=>"000110000",
  52292=>"111111101",
  52293=>"011011100",
  52294=>"010011000",
  52295=>"010011100",
  52296=>"001011010",
  52297=>"110011101",
  52298=>"000111101",
  52299=>"011100100",
  52300=>"000000101",
  52301=>"111010010",
  52302=>"100000110",
  52303=>"010011101",
  52304=>"111100110",
  52305=>"100011110",
  52306=>"111010111",
  52307=>"101001010",
  52308=>"111010011",
  52309=>"111011111",
  52310=>"010001111",
  52311=>"011110001",
  52312=>"111100011",
  52313=>"001110011",
  52314=>"110000101",
  52315=>"101100000",
  52316=>"010011111",
  52317=>"010101000",
  52318=>"110101101",
  52319=>"010110011",
  52320=>"110010010",
  52321=>"000010011",
  52322=>"010001011",
  52323=>"011000010",
  52324=>"101101011",
  52325=>"000100000",
  52326=>"001111101",
  52327=>"110001000",
  52328=>"111001000",
  52329=>"100110100",
  52330=>"100111100",
  52331=>"000010011",
  52332=>"100011010",
  52333=>"101111110",
  52334=>"101101100",
  52335=>"110011011",
  52336=>"011001111",
  52337=>"010001100",
  52338=>"000101011",
  52339=>"100001101",
  52340=>"001010111",
  52341=>"100110011",
  52342=>"110010100",
  52343=>"111001100",
  52344=>"101010111",
  52345=>"110110000",
  52346=>"001100100",
  52347=>"011100001",
  52348=>"111011100",
  52349=>"000101110",
  52350=>"110101010",
  52351=>"100110001",
  52352=>"000011001",
  52353=>"101110111",
  52354=>"000101011",
  52355=>"101100111",
  52356=>"100111100",
  52357=>"000010010",
  52358=>"000111101",
  52359=>"000101000",
  52360=>"011101101",
  52361=>"110010011",
  52362=>"010110011",
  52363=>"011111010",
  52364=>"100000110",
  52365=>"100101001",
  52366=>"101100101",
  52367=>"100100110",
  52368=>"010000000",
  52369=>"101110111",
  52370=>"101111000",
  52371=>"000101110",
  52372=>"110110100",
  52373=>"000000110",
  52374=>"000001000",
  52375=>"011010111",
  52376=>"100001001",
  52377=>"100111011",
  52378=>"010101001",
  52379=>"101100010",
  52380=>"000011111",
  52381=>"000110000",
  52382=>"001110110",
  52383=>"110000110",
  52384=>"011100111",
  52385=>"001001001",
  52386=>"110010010",
  52387=>"101001111",
  52388=>"011100011",
  52389=>"101011111",
  52390=>"100100101",
  52391=>"000101101",
  52392=>"100000010",
  52393=>"001010011",
  52394=>"101110110",
  52395=>"101001010",
  52396=>"101100110",
  52397=>"001101101",
  52398=>"100010000",
  52399=>"010110111",
  52400=>"100110101",
  52401=>"110111000",
  52402=>"111101110",
  52403=>"000101001",
  52404=>"110100000",
  52405=>"110000100",
  52406=>"000111101",
  52407=>"101101000",
  52408=>"001010011",
  52409=>"010000111",
  52410=>"100000011",
  52411=>"011001011",
  52412=>"110000110",
  52413=>"110111101",
  52414=>"001111110",
  52415=>"001111001",
  52416=>"100000001",
  52417=>"010101010",
  52418=>"000111111",
  52419=>"001010101",
  52420=>"011111011",
  52421=>"001111001",
  52422=>"010110100",
  52423=>"010110111",
  52424=>"010011110",
  52425=>"011010111",
  52426=>"010011011",
  52427=>"001110010",
  52428=>"101011100",
  52429=>"100110101",
  52430=>"101001100",
  52431=>"000000010",
  52432=>"000001000",
  52433=>"001010101",
  52434=>"001100110",
  52435=>"011000000",
  52436=>"010100110",
  52437=>"000111101",
  52438=>"001100001",
  52439=>"111111100",
  52440=>"001100101",
  52441=>"110110000",
  52442=>"011110101",
  52443=>"100100011",
  52444=>"111111101",
  52445=>"101010110",
  52446=>"101100010",
  52447=>"100100111",
  52448=>"111110001",
  52449=>"100001101",
  52450=>"001100010",
  52451=>"001011000",
  52452=>"011111010",
  52453=>"010110101",
  52454=>"100111100",
  52455=>"000100010",
  52456=>"110011011",
  52457=>"111010110",
  52458=>"000101110",
  52459=>"111111111",
  52460=>"101011011",
  52461=>"001010100",
  52462=>"001011000",
  52463=>"101111110",
  52464=>"110101110",
  52465=>"100010010",
  52466=>"101011001",
  52467=>"100100000",
  52468=>"111111000",
  52469=>"100001111",
  52470=>"110010101",
  52471=>"101000011",
  52472=>"100010011",
  52473=>"011010001",
  52474=>"110011001",
  52475=>"101001101",
  52476=>"111001100",
  52477=>"011001111",
  52478=>"100000011",
  52479=>"110101011",
  52480=>"110011000",
  52481=>"011110101",
  52482=>"010001011",
  52483=>"010010000",
  52484=>"000010111",
  52485=>"100000110",
  52486=>"010110001",
  52487=>"000100000",
  52488=>"111110101",
  52489=>"100001000",
  52490=>"011000010",
  52491=>"101011001",
  52492=>"010010010",
  52493=>"011100000",
  52494=>"100000100",
  52495=>"100010011",
  52496=>"101111111",
  52497=>"110001010",
  52498=>"110001111",
  52499=>"111111111",
  52500=>"010001010",
  52501=>"100011011",
  52502=>"000100000",
  52503=>"011110100",
  52504=>"101101111",
  52505=>"011000000",
  52506=>"110110011",
  52507=>"101001001",
  52508=>"100110000",
  52509=>"011011011",
  52510=>"011100110",
  52511=>"010101000",
  52512=>"011110010",
  52513=>"011010101",
  52514=>"100101001",
  52515=>"101010010",
  52516=>"101110110",
  52517=>"101111011",
  52518=>"001110000",
  52519=>"110000111",
  52520=>"000000101",
  52521=>"111011111",
  52522=>"000111010",
  52523=>"111101010",
  52524=>"001010010",
  52525=>"100011100",
  52526=>"011110001",
  52527=>"010001100",
  52528=>"010011000",
  52529=>"100101001",
  52530=>"010111011",
  52531=>"100011001",
  52532=>"001101110",
  52533=>"000001100",
  52534=>"010011101",
  52535=>"101011001",
  52536=>"110011111",
  52537=>"110011001",
  52538=>"011100111",
  52539=>"111011100",
  52540=>"110011110",
  52541=>"100000101",
  52542=>"000100001",
  52543=>"001111111",
  52544=>"110000100",
  52545=>"100100000",
  52546=>"110111000",
  52547=>"011001011",
  52548=>"100000011",
  52549=>"011111011",
  52550=>"101000111",
  52551=>"001001001",
  52552=>"101011011",
  52553=>"110000010",
  52554=>"000011100",
  52555=>"001011000",
  52556=>"111011001",
  52557=>"000101111",
  52558=>"101110100",
  52559=>"001110111",
  52560=>"001001100",
  52561=>"101110011",
  52562=>"000111100",
  52563=>"000101111",
  52564=>"100001110",
  52565=>"010000011",
  52566=>"110000010",
  52567=>"100101000",
  52568=>"000101100",
  52569=>"010010010",
  52570=>"100001001",
  52571=>"000110110",
  52572=>"110010011",
  52573=>"001110101",
  52574=>"101010100",
  52575=>"001110100",
  52576=>"110101000",
  52577=>"101010001",
  52578=>"100100110",
  52579=>"000111100",
  52580=>"000100010",
  52581=>"010101101",
  52582=>"001010101",
  52583=>"101101010",
  52584=>"011110011",
  52585=>"100011010",
  52586=>"000100010",
  52587=>"000000101",
  52588=>"000001000",
  52589=>"110011001",
  52590=>"100010110",
  52591=>"010011011",
  52592=>"000000000",
  52593=>"010111011",
  52594=>"111000000",
  52595=>"110011011",
  52596=>"110000001",
  52597=>"000000100",
  52598=>"011010011",
  52599=>"001100001",
  52600=>"011100001",
  52601=>"010101101",
  52602=>"111111010",
  52603=>"000101101",
  52604=>"110000000",
  52605=>"010100000",
  52606=>"010000001",
  52607=>"010001001",
  52608=>"111110001",
  52609=>"111101011",
  52610=>"101000010",
  52611=>"110101100",
  52612=>"101101101",
  52613=>"000110011",
  52614=>"100100111",
  52615=>"001100111",
  52616=>"011010010",
  52617=>"110100100",
  52618=>"111010110",
  52619=>"000001001",
  52620=>"110101100",
  52621=>"010011111",
  52622=>"000011001",
  52623=>"010100011",
  52624=>"101101000",
  52625=>"101000110",
  52626=>"001000111",
  52627=>"111010011",
  52628=>"110111100",
  52629=>"000110000",
  52630=>"101001111",
  52631=>"010100101",
  52632=>"010100100",
  52633=>"000000000",
  52634=>"001100101",
  52635=>"000010011",
  52636=>"011010100",
  52637=>"101010100",
  52638=>"001100000",
  52639=>"110011100",
  52640=>"011000011",
  52641=>"010111101",
  52642=>"111101100",
  52643=>"100000000",
  52644=>"110111100",
  52645=>"011110000",
  52646=>"000001001",
  52647=>"010011000",
  52648=>"111010111",
  52649=>"011110000",
  52650=>"011001100",
  52651=>"000101011",
  52652=>"110100100",
  52653=>"100100100",
  52654=>"000010100",
  52655=>"000011011",
  52656=>"001100000",
  52657=>"001101000",
  52658=>"001110111",
  52659=>"001000001",
  52660=>"100010110",
  52661=>"111001011",
  52662=>"010011101",
  52663=>"011100111",
  52664=>"111010010",
  52665=>"000000111",
  52666=>"000000101",
  52667=>"100111000",
  52668=>"101000010",
  52669=>"010001001",
  52670=>"101000111",
  52671=>"101110111",
  52672=>"110010011",
  52673=>"011101110",
  52674=>"101100001",
  52675=>"111010000",
  52676=>"000110011",
  52677=>"000100000",
  52678=>"010000010",
  52679=>"000111000",
  52680=>"111100010",
  52681=>"000100000",
  52682=>"000000001",
  52683=>"010101011",
  52684=>"000101001",
  52685=>"000000111",
  52686=>"111011001",
  52687=>"101100110",
  52688=>"011001111",
  52689=>"110011000",
  52690=>"011000010",
  52691=>"011001001",
  52692=>"111100010",
  52693=>"000101111",
  52694=>"011010000",
  52695=>"011010000",
  52696=>"111011000",
  52697=>"101100010",
  52698=>"100101110",
  52699=>"001101000",
  52700=>"111101000",
  52701=>"100011110",
  52702=>"001111100",
  52703=>"010100001",
  52704=>"011111111",
  52705=>"110011110",
  52706=>"110111000",
  52707=>"111101110",
  52708=>"001010101",
  52709=>"101111011",
  52710=>"100010010",
  52711=>"001111000",
  52712=>"110100000",
  52713=>"100001000",
  52714=>"001010011",
  52715=>"011011110",
  52716=>"000110010",
  52717=>"001000000",
  52718=>"010011001",
  52719=>"111001100",
  52720=>"110010101",
  52721=>"010011000",
  52722=>"001101001",
  52723=>"010010100",
  52724=>"011000010",
  52725=>"010110010",
  52726=>"101111001",
  52727=>"001101011",
  52728=>"010001011",
  52729=>"000000011",
  52730=>"001001001",
  52731=>"101101110",
  52732=>"001001101",
  52733=>"011110001",
  52734=>"111100111",
  52735=>"110100001",
  52736=>"101100110",
  52737=>"000101110",
  52738=>"110000001",
  52739=>"011001010",
  52740=>"000001101",
  52741=>"100100110",
  52742=>"110110001",
  52743=>"100100101",
  52744=>"101010100",
  52745=>"000011111",
  52746=>"111100100",
  52747=>"011001110",
  52748=>"111111111",
  52749=>"001100101",
  52750=>"000110000",
  52751=>"000111010",
  52752=>"001011101",
  52753=>"110001000",
  52754=>"011101010",
  52755=>"011010110",
  52756=>"100010001",
  52757=>"001101111",
  52758=>"001001001",
  52759=>"100110010",
  52760=>"011100110",
  52761=>"110100001",
  52762=>"011000001",
  52763=>"001000001",
  52764=>"010010000",
  52765=>"001010010",
  52766=>"001010110",
  52767=>"110100001",
  52768=>"011001111",
  52769=>"011111111",
  52770=>"011011111",
  52771=>"100000000",
  52772=>"100000111",
  52773=>"011000000",
  52774=>"010011101",
  52775=>"100000101",
  52776=>"101111100",
  52777=>"010110101",
  52778=>"101000110",
  52779=>"010001001",
  52780=>"101100111",
  52781=>"000101000",
  52782=>"110111000",
  52783=>"000000010",
  52784=>"010011011",
  52785=>"001001001",
  52786=>"001010000",
  52787=>"010100001",
  52788=>"100101011",
  52789=>"011001101",
  52790=>"010111111",
  52791=>"110110010",
  52792=>"111101001",
  52793=>"100101111",
  52794=>"011111101",
  52795=>"100001011",
  52796=>"100110111",
  52797=>"110100000",
  52798=>"011100000",
  52799=>"100100100",
  52800=>"011000001",
  52801=>"110111000",
  52802=>"100111000",
  52803=>"000100100",
  52804=>"011111010",
  52805=>"101111010",
  52806=>"010001110",
  52807=>"100100001",
  52808=>"000001101",
  52809=>"110010110",
  52810=>"110111001",
  52811=>"010000111",
  52812=>"100001101",
  52813=>"000011111",
  52814=>"010010010",
  52815=>"010100011",
  52816=>"010110000",
  52817=>"000100001",
  52818=>"011101100",
  52819=>"010011011",
  52820=>"011101110",
  52821=>"011010011",
  52822=>"000000000",
  52823=>"111101111",
  52824=>"100110110",
  52825=>"000111101",
  52826=>"000111101",
  52827=>"110000101",
  52828=>"011000001",
  52829=>"000000101",
  52830=>"110001110",
  52831=>"010000110",
  52832=>"100000011",
  52833=>"101101000",
  52834=>"111101001",
  52835=>"000001101",
  52836=>"000011011",
  52837=>"110110110",
  52838=>"110001111",
  52839=>"010010100",
  52840=>"001111010",
  52841=>"011000000",
  52842=>"111110111",
  52843=>"000000000",
  52844=>"010100011",
  52845=>"001111011",
  52846=>"001001010",
  52847=>"010000101",
  52848=>"111111011",
  52849=>"111100010",
  52850=>"010001100",
  52851=>"001000111",
  52852=>"111010011",
  52853=>"000000000",
  52854=>"001110100",
  52855=>"011101011",
  52856=>"110011111",
  52857=>"110011001",
  52858=>"011011100",
  52859=>"111001101",
  52860=>"000010101",
  52861=>"100000111",
  52862=>"100111110",
  52863=>"001001111",
  52864=>"101110110",
  52865=>"110101111",
  52866=>"100100111",
  52867=>"100110101",
  52868=>"001110011",
  52869=>"010101000",
  52870=>"000110100",
  52871=>"101111001",
  52872=>"010011010",
  52873=>"111001100",
  52874=>"000100011",
  52875=>"000010010",
  52876=>"100111101",
  52877=>"100011000",
  52878=>"110110010",
  52879=>"010110100",
  52880=>"000011000",
  52881=>"001010010",
  52882=>"100011001",
  52883=>"101111101",
  52884=>"000010000",
  52885=>"101011011",
  52886=>"011101000",
  52887=>"001001010",
  52888=>"010111010",
  52889=>"011101100",
  52890=>"011001100",
  52891=>"011001100",
  52892=>"110010110",
  52893=>"100011010",
  52894=>"000010010",
  52895=>"001100100",
  52896=>"100010001",
  52897=>"000100111",
  52898=>"010001110",
  52899=>"010100110",
  52900=>"000000111",
  52901=>"110111001",
  52902=>"000000001",
  52903=>"000101110",
  52904=>"010001011",
  52905=>"000100001",
  52906=>"001111001",
  52907=>"100110100",
  52908=>"110111011",
  52909=>"111000101",
  52910=>"000000101",
  52911=>"001111001",
  52912=>"001110000",
  52913=>"100110101",
  52914=>"101010001",
  52915=>"010011011",
  52916=>"001001011",
  52917=>"100110101",
  52918=>"110111010",
  52919=>"010101101",
  52920=>"100001001",
  52921=>"100000011",
  52922=>"001100110",
  52923=>"001110001",
  52924=>"000100010",
  52925=>"010001011",
  52926=>"001100000",
  52927=>"110111001",
  52928=>"111100011",
  52929=>"111100100",
  52930=>"111000000",
  52931=>"001011111",
  52932=>"000011000",
  52933=>"000111010",
  52934=>"100011000",
  52935=>"100010110",
  52936=>"111101111",
  52937=>"000101001",
  52938=>"000000010",
  52939=>"111100110",
  52940=>"000010011",
  52941=>"111110111",
  52942=>"000011011",
  52943=>"001111111",
  52944=>"001110001",
  52945=>"010100110",
  52946=>"111100011",
  52947=>"000011000",
  52948=>"101110110",
  52949=>"011011001",
  52950=>"010001000",
  52951=>"011010100",
  52952=>"000010001",
  52953=>"110010110",
  52954=>"100010111",
  52955=>"100010111",
  52956=>"101110000",
  52957=>"000111011",
  52958=>"111100101",
  52959=>"001101111",
  52960=>"101100101",
  52961=>"001010011",
  52962=>"011010100",
  52963=>"100000000",
  52964=>"011101011",
  52965=>"010101100",
  52966=>"111000000",
  52967=>"110010101",
  52968=>"010000110",
  52969=>"111010011",
  52970=>"000010111",
  52971=>"010101001",
  52972=>"001100010",
  52973=>"111011111",
  52974=>"110111111",
  52975=>"110110110",
  52976=>"111111001",
  52977=>"100001000",
  52978=>"001011101",
  52979=>"010100101",
  52980=>"000111011",
  52981=>"100000011",
  52982=>"100010001",
  52983=>"110110110",
  52984=>"010000011",
  52985=>"010001110",
  52986=>"100011001",
  52987=>"001001000",
  52988=>"011101011",
  52989=>"100100010",
  52990=>"001110010",
  52991=>"000110010",
  52992=>"100101000",
  52993=>"011110010",
  52994=>"110000011",
  52995=>"010111000",
  52996=>"100110110",
  52997=>"001111111",
  52998=>"100111110",
  52999=>"111111001",
  53000=>"000011001",
  53001=>"110011100",
  53002=>"000011100",
  53003=>"111010001",
  53004=>"010001101",
  53005=>"101101011",
  53006=>"101010001",
  53007=>"111010010",
  53008=>"010000001",
  53009=>"000100100",
  53010=>"000011101",
  53011=>"001010110",
  53012=>"011101011",
  53013=>"110111011",
  53014=>"111100001",
  53015=>"000100000",
  53016=>"001001011",
  53017=>"011110110",
  53018=>"100011110",
  53019=>"101011011",
  53020=>"011001101",
  53021=>"110110100",
  53022=>"110110111",
  53023=>"000010011",
  53024=>"100000101",
  53025=>"111001000",
  53026=>"111111001",
  53027=>"101011010",
  53028=>"100100000",
  53029=>"011110000",
  53030=>"010101010",
  53031=>"101101100",
  53032=>"001001001",
  53033=>"101111110",
  53034=>"001110100",
  53035=>"001101110",
  53036=>"100011010",
  53037=>"000001000",
  53038=>"011000010",
  53039=>"110000001",
  53040=>"101011110",
  53041=>"011110101",
  53042=>"101001001",
  53043=>"101100001",
  53044=>"000010110",
  53045=>"001010100",
  53046=>"100011100",
  53047=>"000011100",
  53048=>"011110100",
  53049=>"010100010",
  53050=>"111111000",
  53051=>"010000001",
  53052=>"010100101",
  53053=>"010000000",
  53054=>"100000001",
  53055=>"011000000",
  53056=>"010010100",
  53057=>"110010110",
  53058=>"101011010",
  53059=>"100111011",
  53060=>"010100111",
  53061=>"101011101",
  53062=>"001110111",
  53063=>"001001101",
  53064=>"000010100",
  53065=>"111011101",
  53066=>"110111101",
  53067=>"010000101",
  53068=>"010000111",
  53069=>"111011100",
  53070=>"110110100",
  53071=>"111111100",
  53072=>"101100000",
  53073=>"010010000",
  53074=>"110010111",
  53075=>"000000011",
  53076=>"001001101",
  53077=>"000111100",
  53078=>"100001101",
  53079=>"100010010",
  53080=>"101000110",
  53081=>"110101010",
  53082=>"110101000",
  53083=>"010000000",
  53084=>"010011101",
  53085=>"011011001",
  53086=>"100010001",
  53087=>"101001000",
  53088=>"101100101",
  53089=>"001000000",
  53090=>"000100111",
  53091=>"010110100",
  53092=>"010101100",
  53093=>"101110011",
  53094=>"110110100",
  53095=>"101101010",
  53096=>"100011000",
  53097=>"001100011",
  53098=>"001010010",
  53099=>"101000100",
  53100=>"010101001",
  53101=>"000011011",
  53102=>"000011000",
  53103=>"001101001",
  53104=>"101000110",
  53105=>"011100000",
  53106=>"110100011",
  53107=>"110111110",
  53108=>"000011111",
  53109=>"101001110",
  53110=>"111101100",
  53111=>"001000000",
  53112=>"100100100",
  53113=>"110110111",
  53114=>"000110101",
  53115=>"010000110",
  53116=>"000100001",
  53117=>"011111000",
  53118=>"111011111",
  53119=>"100101101",
  53120=>"100100101",
  53121=>"101000011",
  53122=>"111111101",
  53123=>"111111100",
  53124=>"100010000",
  53125=>"101011100",
  53126=>"000110010",
  53127=>"000100110",
  53128=>"100010110",
  53129=>"011001101",
  53130=>"011101110",
  53131=>"001101011",
  53132=>"000110001",
  53133=>"001011101",
  53134=>"110111110",
  53135=>"110001101",
  53136=>"010101000",
  53137=>"100010110",
  53138=>"000001110",
  53139=>"000000010",
  53140=>"101011101",
  53141=>"110011011",
  53142=>"000111001",
  53143=>"000001101",
  53144=>"011010010",
  53145=>"001000110",
  53146=>"110010001",
  53147=>"001111010",
  53148=>"110011011",
  53149=>"000110110",
  53150=>"000000000",
  53151=>"101000001",
  53152=>"111101111",
  53153=>"011001000",
  53154=>"101010001",
  53155=>"011010100",
  53156=>"110010101",
  53157=>"111110110",
  53158=>"100111100",
  53159=>"110011010",
  53160=>"110101100",
  53161=>"111100000",
  53162=>"110000101",
  53163=>"110001001",
  53164=>"010101100",
  53165=>"100101001",
  53166=>"011111000",
  53167=>"100101010",
  53168=>"100100111",
  53169=>"100001101",
  53170=>"101001111",
  53171=>"010110011",
  53172=>"111101011",
  53173=>"110110010",
  53174=>"000110011",
  53175=>"111011001",
  53176=>"111110101",
  53177=>"111111001",
  53178=>"000101111",
  53179=>"011001100",
  53180=>"011010010",
  53181=>"010111011",
  53182=>"110110011",
  53183=>"011111111",
  53184=>"100110010",
  53185=>"010001001",
  53186=>"110000010",
  53187=>"010100000",
  53188=>"110110010",
  53189=>"100001011",
  53190=>"101111111",
  53191=>"111010111",
  53192=>"001000000",
  53193=>"000000011",
  53194=>"000000001",
  53195=>"000001010",
  53196=>"001111010",
  53197=>"110000101",
  53198=>"000110100",
  53199=>"101010101",
  53200=>"010110101",
  53201=>"001000000",
  53202=>"101111100",
  53203=>"111001110",
  53204=>"011010010",
  53205=>"101100010",
  53206=>"100000000",
  53207=>"110101110",
  53208=>"100111101",
  53209=>"010010101",
  53210=>"001110101",
  53211=>"100000110",
  53212=>"001001110",
  53213=>"111001111",
  53214=>"011111101",
  53215=>"110110001",
  53216=>"101011101",
  53217=>"000100011",
  53218=>"111101110",
  53219=>"001110101",
  53220=>"000000110",
  53221=>"000010000",
  53222=>"000100000",
  53223=>"000010000",
  53224=>"011101101",
  53225=>"111010011",
  53226=>"001001101",
  53227=>"000111011",
  53228=>"100001000",
  53229=>"010101001",
  53230=>"100000100",
  53231=>"111000011",
  53232=>"010101001",
  53233=>"110101010",
  53234=>"010001100",
  53235=>"011001111",
  53236=>"111011100",
  53237=>"001000101",
  53238=>"101001011",
  53239=>"101111100",
  53240=>"000000000",
  53241=>"110010000",
  53242=>"001010110",
  53243=>"000010001",
  53244=>"111011001",
  53245=>"111001000",
  53246=>"010001001",
  53247=>"111011000",
  53248=>"100110010",
  53249=>"110000100",
  53250=>"001101010",
  53251=>"110010100",
  53252=>"000100000",
  53253=>"000000110",
  53254=>"100111001",
  53255=>"111001011",
  53256=>"000010011",
  53257=>"011101101",
  53258=>"010000100",
  53259=>"100100010",
  53260=>"111101001",
  53261=>"000010000",
  53262=>"011111101",
  53263=>"001010001",
  53264=>"111100001",
  53265=>"011001010",
  53266=>"010001101",
  53267=>"000000011",
  53268=>"011010000",
  53269=>"110000100",
  53270=>"101010110",
  53271=>"000101101",
  53272=>"010100010",
  53273=>"101101000",
  53274=>"101100111",
  53275=>"111110010",
  53276=>"011100100",
  53277=>"111001001",
  53278=>"001000010",
  53279=>"111101000",
  53280=>"100011000",
  53281=>"101101010",
  53282=>"110000111",
  53283=>"100101100",
  53284=>"101101000",
  53285=>"111001100",
  53286=>"100111101",
  53287=>"000111011",
  53288=>"110111011",
  53289=>"000000000",
  53290=>"101110101",
  53291=>"101010000",
  53292=>"000011000",
  53293=>"100000010",
  53294=>"010010100",
  53295=>"000000001",
  53296=>"010001110",
  53297=>"010101100",
  53298=>"011011101",
  53299=>"111111110",
  53300=>"111111101",
  53301=>"101011101",
  53302=>"010110101",
  53303=>"011100101",
  53304=>"000010001",
  53305=>"110001100",
  53306=>"101111010",
  53307=>"011011101",
  53308=>"100110111",
  53309=>"001001000",
  53310=>"000001101",
  53311=>"011100011",
  53312=>"000111100",
  53313=>"000110000",
  53314=>"011100111",
  53315=>"111010101",
  53316=>"100100000",
  53317=>"011110010",
  53318=>"110001111",
  53319=>"110100101",
  53320=>"000101001",
  53321=>"101010101",
  53322=>"010000000",
  53323=>"111001111",
  53324=>"000001111",
  53325=>"110000001",
  53326=>"011101001",
  53327=>"101110110",
  53328=>"011111001",
  53329=>"000011010",
  53330=>"111001000",
  53331=>"000000001",
  53332=>"110000101",
  53333=>"000001011",
  53334=>"011111111",
  53335=>"101100111",
  53336=>"011000010",
  53337=>"001000100",
  53338=>"100101100",
  53339=>"111000000",
  53340=>"000100010",
  53341=>"111100001",
  53342=>"100100100",
  53343=>"010101111",
  53344=>"011011000",
  53345=>"101101101",
  53346=>"100101010",
  53347=>"011111010",
  53348=>"101001100",
  53349=>"100101001",
  53350=>"000010111",
  53351=>"111111011",
  53352=>"001000110",
  53353=>"010111010",
  53354=>"010000111",
  53355=>"110000001",
  53356=>"001000100",
  53357=>"010011111",
  53358=>"101001111",
  53359=>"010100011",
  53360=>"110110110",
  53361=>"011011110",
  53362=>"011110101",
  53363=>"001010001",
  53364=>"111000111",
  53365=>"101101001",
  53366=>"111111001",
  53367=>"010000100",
  53368=>"001111000",
  53369=>"000100011",
  53370=>"010001010",
  53371=>"000111010",
  53372=>"001000001",
  53373=>"110100000",
  53374=>"101010110",
  53375=>"101000001",
  53376=>"000011010",
  53377=>"110011111",
  53378=>"011101100",
  53379=>"111101101",
  53380=>"110101100",
  53381=>"000011110",
  53382=>"101100000",
  53383=>"111010001",
  53384=>"000011011",
  53385=>"011010000",
  53386=>"110100111",
  53387=>"100101011",
  53388=>"000001011",
  53389=>"100010101",
  53390=>"110111011",
  53391=>"000100100",
  53392=>"101111110",
  53393=>"101001100",
  53394=>"110011110",
  53395=>"001101011",
  53396=>"111010101",
  53397=>"000111011",
  53398=>"111011000",
  53399=>"110011100",
  53400=>"011101100",
  53401=>"110101000",
  53402=>"100110110",
  53403=>"110010111",
  53404=>"111110000",
  53405=>"001111100",
  53406=>"100110011",
  53407=>"011110001",
  53408=>"100000010",
  53409=>"010101100",
  53410=>"100100000",
  53411=>"001001001",
  53412=>"011011100",
  53413=>"000110011",
  53414=>"100111000",
  53415=>"100000000",
  53416=>"001011001",
  53417=>"111101011",
  53418=>"111110110",
  53419=>"000000000",
  53420=>"111010110",
  53421=>"110101101",
  53422=>"111011011",
  53423=>"000110111",
  53424=>"011000001",
  53425=>"110000011",
  53426=>"111101100",
  53427=>"101100001",
  53428=>"011101111",
  53429=>"011111101",
  53430=>"000110010",
  53431=>"011001110",
  53432=>"110010110",
  53433=>"010010111",
  53434=>"011101000",
  53435=>"110101000",
  53436=>"001001101",
  53437=>"010100000",
  53438=>"011000001",
  53439=>"000110111",
  53440=>"100010100",
  53441=>"001111100",
  53442=>"111101101",
  53443=>"010001000",
  53444=>"110001101",
  53445=>"100110110",
  53446=>"111110011",
  53447=>"101011010",
  53448=>"011011010",
  53449=>"011111001",
  53450=>"000101101",
  53451=>"110101001",
  53452=>"100110011",
  53453=>"011010000",
  53454=>"001110111",
  53455=>"011010110",
  53456=>"011001101",
  53457=>"010010100",
  53458=>"001000000",
  53459=>"010100000",
  53460=>"000101111",
  53461=>"010011011",
  53462=>"111100011",
  53463=>"101100000",
  53464=>"110100100",
  53465=>"011110100",
  53466=>"010101100",
  53467=>"000000010",
  53468=>"000111011",
  53469=>"000101000",
  53470=>"101001000",
  53471=>"110100010",
  53472=>"110101000",
  53473=>"101101101",
  53474=>"010100101",
  53475=>"000010100",
  53476=>"010001101",
  53477=>"111000111",
  53478=>"110110100",
  53479=>"011001100",
  53480=>"101000011",
  53481=>"101000110",
  53482=>"000000010",
  53483=>"010100011",
  53484=>"101011011",
  53485=>"100001011",
  53486=>"101001011",
  53487=>"111111000",
  53488=>"100111111",
  53489=>"001001000",
  53490=>"110111001",
  53491=>"011111111",
  53492=>"001010000",
  53493=>"000000001",
  53494=>"111110001",
  53495=>"000011100",
  53496=>"001100000",
  53497=>"111000100",
  53498=>"111100101",
  53499=>"000101001",
  53500=>"110100100",
  53501=>"011111111",
  53502=>"111111101",
  53503=>"011110010",
  53504=>"000111101",
  53505=>"011100000",
  53506=>"101000100",
  53507=>"111110011",
  53508=>"101110101",
  53509=>"100010100",
  53510=>"010001001",
  53511=>"001100111",
  53512=>"111101100",
  53513=>"111111000",
  53514=>"011001110",
  53515=>"010010110",
  53516=>"001110001",
  53517=>"110111111",
  53518=>"001110100",
  53519=>"110101001",
  53520=>"101010110",
  53521=>"101010010",
  53522=>"111101011",
  53523=>"101011000",
  53524=>"000010000",
  53525=>"101010100",
  53526=>"000101111",
  53527=>"111000001",
  53528=>"011100011",
  53529=>"100001010",
  53530=>"110000100",
  53531=>"000110101",
  53532=>"101101001",
  53533=>"001001001",
  53534=>"100001100",
  53535=>"101000001",
  53536=>"100101110",
  53537=>"011000001",
  53538=>"100010001",
  53539=>"100100000",
  53540=>"010001100",
  53541=>"010110000",
  53542=>"000010011",
  53543=>"001000011",
  53544=>"110001010",
  53545=>"101011000",
  53546=>"111111101",
  53547=>"000000010",
  53548=>"110010100",
  53549=>"110000011",
  53550=>"001100101",
  53551=>"010111111",
  53552=>"011001110",
  53553=>"111111100",
  53554=>"001111100",
  53555=>"100011000",
  53556=>"100100111",
  53557=>"000111111",
  53558=>"000000100",
  53559=>"100001000",
  53560=>"001010100",
  53561=>"111011001",
  53562=>"100000100",
  53563=>"001010101",
  53564=>"010011111",
  53565=>"101101001",
  53566=>"000111101",
  53567=>"101001100",
  53568=>"001010110",
  53569=>"111111101",
  53570=>"111101000",
  53571=>"001011001",
  53572=>"110100100",
  53573=>"001100111",
  53574=>"100000001",
  53575=>"011101100",
  53576=>"111111011",
  53577=>"110010011",
  53578=>"001001001",
  53579=>"000111111",
  53580=>"011101010",
  53581=>"111100111",
  53582=>"010010000",
  53583=>"101100001",
  53584=>"000010001",
  53585=>"110010111",
  53586=>"000110011",
  53587=>"101001111",
  53588=>"000101011",
  53589=>"101111111",
  53590=>"010101100",
  53591=>"111011010",
  53592=>"010101010",
  53593=>"011101001",
  53594=>"000100100",
  53595=>"101011100",
  53596=>"011110111",
  53597=>"111101111",
  53598=>"111100101",
  53599=>"100001101",
  53600=>"111000100",
  53601=>"010001100",
  53602=>"000111100",
  53603=>"111111000",
  53604=>"010100101",
  53605=>"101100001",
  53606=>"001011100",
  53607=>"100110000",
  53608=>"001010011",
  53609=>"011000001",
  53610=>"101100111",
  53611=>"011001101",
  53612=>"110000010",
  53613=>"011001010",
  53614=>"111011001",
  53615=>"101100111",
  53616=>"010000011",
  53617=>"011001111",
  53618=>"111011001",
  53619=>"100000010",
  53620=>"100111010",
  53621=>"011110011",
  53622=>"001111010",
  53623=>"011111100",
  53624=>"111110110",
  53625=>"110100001",
  53626=>"100100001",
  53627=>"000011011",
  53628=>"100100010",
  53629=>"110000111",
  53630=>"000000010",
  53631=>"101110111",
  53632=>"101011011",
  53633=>"111110101",
  53634=>"001001011",
  53635=>"111101100",
  53636=>"011001001",
  53637=>"001101110",
  53638=>"001110010",
  53639=>"111101110",
  53640=>"010111011",
  53641=>"001001010",
  53642=>"000010110",
  53643=>"100101100",
  53644=>"110100101",
  53645=>"000101001",
  53646=>"000101100",
  53647=>"110010000",
  53648=>"111110010",
  53649=>"011101010",
  53650=>"111100001",
  53651=>"111000100",
  53652=>"001111001",
  53653=>"001001101",
  53654=>"100100000",
  53655=>"000111100",
  53656=>"011010001",
  53657=>"011010001",
  53658=>"110001001",
  53659=>"000000010",
  53660=>"110000111",
  53661=>"010110011",
  53662=>"010010000",
  53663=>"110101110",
  53664=>"101100001",
  53665=>"111101101",
  53666=>"101111100",
  53667=>"110111110",
  53668=>"100101000",
  53669=>"100000011",
  53670=>"111001111",
  53671=>"000000110",
  53672=>"100111101",
  53673=>"101101101",
  53674=>"101000111",
  53675=>"110100111",
  53676=>"110100001",
  53677=>"100110111",
  53678=>"101100110",
  53679=>"011011001",
  53680=>"100100100",
  53681=>"010011111",
  53682=>"100101100",
  53683=>"011010000",
  53684=>"011001100",
  53685=>"011110001",
  53686=>"010010001",
  53687=>"010101000",
  53688=>"100000101",
  53689=>"001100000",
  53690=>"100101111",
  53691=>"100100000",
  53692=>"101010101",
  53693=>"011001001",
  53694=>"011100000",
  53695=>"001100111",
  53696=>"011010111",
  53697=>"001000001",
  53698=>"000110001",
  53699=>"001010111",
  53700=>"111101111",
  53701=>"010010001",
  53702=>"000010111",
  53703=>"101100000",
  53704=>"111000000",
  53705=>"100010111",
  53706=>"110101100",
  53707=>"000000001",
  53708=>"111000111",
  53709=>"001000101",
  53710=>"010111011",
  53711=>"110000010",
  53712=>"101011111",
  53713=>"010110011",
  53714=>"001100001",
  53715=>"011101000",
  53716=>"100101100",
  53717=>"111100011",
  53718=>"000011100",
  53719=>"000001110",
  53720=>"010000000",
  53721=>"110101000",
  53722=>"111101010",
  53723=>"101000010",
  53724=>"111110110",
  53725=>"011100000",
  53726=>"110010110",
  53727=>"100110001",
  53728=>"100111000",
  53729=>"101000000",
  53730=>"001110011",
  53731=>"101011011",
  53732=>"001000101",
  53733=>"001011011",
  53734=>"000000110",
  53735=>"100010010",
  53736=>"111100110",
  53737=>"111101011",
  53738=>"100101000",
  53739=>"000110111",
  53740=>"010001000",
  53741=>"001100000",
  53742=>"100000000",
  53743=>"111101111",
  53744=>"100100000",
  53745=>"001111010",
  53746=>"101110111",
  53747=>"100110110",
  53748=>"001101101",
  53749=>"101111110",
  53750=>"111011011",
  53751=>"001110111",
  53752=>"001011111",
  53753=>"100000100",
  53754=>"111100001",
  53755=>"010000100",
  53756=>"111110111",
  53757=>"000000110",
  53758=>"111110110",
  53759=>"010010011",
  53760=>"010011000",
  53761=>"000110010",
  53762=>"100101000",
  53763=>"000111001",
  53764=>"101011011",
  53765=>"000111100",
  53766=>"001110111",
  53767=>"011000011",
  53768=>"010100001",
  53769=>"000001110",
  53770=>"111110100",
  53771=>"101000100",
  53772=>"011111000",
  53773=>"110011001",
  53774=>"000000011",
  53775=>"001101000",
  53776=>"001100010",
  53777=>"011101110",
  53778=>"101010000",
  53779=>"110011100",
  53780=>"001011100",
  53781=>"000101010",
  53782=>"111111111",
  53783=>"101100011",
  53784=>"110011001",
  53785=>"110001000",
  53786=>"011001100",
  53787=>"000111001",
  53788=>"001111010",
  53789=>"100100101",
  53790=>"001010010",
  53791=>"110000010",
  53792=>"000100101",
  53793=>"010001100",
  53794=>"001000001",
  53795=>"101110000",
  53796=>"000101100",
  53797=>"001111100",
  53798=>"010100101",
  53799=>"100010010",
  53800=>"010001110",
  53801=>"111110110",
  53802=>"001001000",
  53803=>"100011011",
  53804=>"011100010",
  53805=>"011111110",
  53806=>"010101111",
  53807=>"100111101",
  53808=>"001010100",
  53809=>"101101000",
  53810=>"000110011",
  53811=>"100101111",
  53812=>"101111001",
  53813=>"010110010",
  53814=>"111100000",
  53815=>"001100001",
  53816=>"010111001",
  53817=>"010000101",
  53818=>"101010011",
  53819=>"001000001",
  53820=>"001100001",
  53821=>"001000111",
  53822=>"000101001",
  53823=>"111110110",
  53824=>"001011011",
  53825=>"011010101",
  53826=>"000000010",
  53827=>"110110010",
  53828=>"010111001",
  53829=>"110101010",
  53830=>"100101100",
  53831=>"001101101",
  53832=>"011111011",
  53833=>"111001000",
  53834=>"000001010",
  53835=>"100010101",
  53836=>"000000101",
  53837=>"101000010",
  53838=>"110110011",
  53839=>"000011111",
  53840=>"111101000",
  53841=>"100000011",
  53842=>"010101010",
  53843=>"101000111",
  53844=>"001011110",
  53845=>"000100011",
  53846=>"110100110",
  53847=>"100010010",
  53848=>"011010100",
  53849=>"111001000",
  53850=>"110001001",
  53851=>"001001010",
  53852=>"101100101",
  53853=>"100110001",
  53854=>"110110000",
  53855=>"011000110",
  53856=>"010100100",
  53857=>"100111100",
  53858=>"001000000",
  53859=>"100000000",
  53860=>"111101001",
  53861=>"000100010",
  53862=>"001110001",
  53863=>"000100011",
  53864=>"001001010",
  53865=>"010100110",
  53866=>"111001011",
  53867=>"001100000",
  53868=>"110100100",
  53869=>"110110000",
  53870=>"000000000",
  53871=>"010100010",
  53872=>"010000001",
  53873=>"100000011",
  53874=>"011000101",
  53875=>"101100011",
  53876=>"001000101",
  53877=>"100010000",
  53878=>"111001000",
  53879=>"000100111",
  53880=>"101000101",
  53881=>"101010001",
  53882=>"110011011",
  53883=>"100001011",
  53884=>"100001011",
  53885=>"111110100",
  53886=>"001101010",
  53887=>"100011101",
  53888=>"001110000",
  53889=>"110001110",
  53890=>"000111100",
  53891=>"000001101",
  53892=>"110011110",
  53893=>"000110010",
  53894=>"101111101",
  53895=>"000011010",
  53896=>"001011010",
  53897=>"001100001",
  53898=>"110110101",
  53899=>"101101110",
  53900=>"011000001",
  53901=>"001000000",
  53902=>"000010111",
  53903=>"010100100",
  53904=>"110001110",
  53905=>"010001000",
  53906=>"010011001",
  53907=>"011110111",
  53908=>"111110101",
  53909=>"101110111",
  53910=>"110101010",
  53911=>"011111001",
  53912=>"101011101",
  53913=>"000000001",
  53914=>"000010011",
  53915=>"100110000",
  53916=>"001110010",
  53917=>"010111101",
  53918=>"100100010",
  53919=>"000101110",
  53920=>"011101001",
  53921=>"011111110",
  53922=>"100110010",
  53923=>"000010000",
  53924=>"111010101",
  53925=>"101111111",
  53926=>"010011000",
  53927=>"101011101",
  53928=>"010010111",
  53929=>"000110110",
  53930=>"001000001",
  53931=>"010110101",
  53932=>"010011111",
  53933=>"100101011",
  53934=>"011011001",
  53935=>"111100011",
  53936=>"000100101",
  53937=>"111111111",
  53938=>"111000101",
  53939=>"111111001",
  53940=>"000011000",
  53941=>"110001101",
  53942=>"110001010",
  53943=>"010000001",
  53944=>"000000001",
  53945=>"010011101",
  53946=>"101101000",
  53947=>"000011000",
  53948=>"110001110",
  53949=>"000100101",
  53950=>"000001111",
  53951=>"111011011",
  53952=>"101111011",
  53953=>"101000110",
  53954=>"010101000",
  53955=>"010011011",
  53956=>"111101110",
  53957=>"100011000",
  53958=>"001011100",
  53959=>"000101110",
  53960=>"000100010",
  53961=>"011010000",
  53962=>"000111101",
  53963=>"111000101",
  53964=>"000000110",
  53965=>"100000101",
  53966=>"000001100",
  53967=>"010101011",
  53968=>"001001000",
  53969=>"010011011",
  53970=>"010110110",
  53971=>"000111001",
  53972=>"000011001",
  53973=>"111101010",
  53974=>"110000010",
  53975=>"101100111",
  53976=>"110001000",
  53977=>"111001000",
  53978=>"011010000",
  53979=>"000011000",
  53980=>"011010110",
  53981=>"001111000",
  53982=>"111010001",
  53983=>"101000110",
  53984=>"000110110",
  53985=>"001000000",
  53986=>"000001001",
  53987=>"000000010",
  53988=>"001000010",
  53989=>"001111101",
  53990=>"001011000",
  53991=>"101010011",
  53992=>"010100011",
  53993=>"110011000",
  53994=>"001000001",
  53995=>"101011111",
  53996=>"000110100",
  53997=>"000110101",
  53998=>"011001100",
  53999=>"010000001",
  54000=>"000101111",
  54001=>"110001100",
  54002=>"101111000",
  54003=>"000011101",
  54004=>"101110100",
  54005=>"111111011",
  54006=>"111111000",
  54007=>"100101110",
  54008=>"110010110",
  54009=>"101001001",
  54010=>"001101110",
  54011=>"001000100",
  54012=>"001001001",
  54013=>"111010100",
  54014=>"001011001",
  54015=>"101111011",
  54016=>"010100101",
  54017=>"100000010",
  54018=>"100011100",
  54019=>"110111100",
  54020=>"101001100",
  54021=>"010000000",
  54022=>"101111110",
  54023=>"101101000",
  54024=>"001000100",
  54025=>"011001110",
  54026=>"010000011",
  54027=>"110011101",
  54028=>"100100000",
  54029=>"100010001",
  54030=>"001100100",
  54031=>"011101101",
  54032=>"110011010",
  54033=>"101001011",
  54034=>"011000110",
  54035=>"010011111",
  54036=>"100011101",
  54037=>"001111111",
  54038=>"011000110",
  54039=>"100000000",
  54040=>"001000000",
  54041=>"100000010",
  54042=>"111000101",
  54043=>"110000110",
  54044=>"111110101",
  54045=>"011000010",
  54046=>"000000111",
  54047=>"100101010",
  54048=>"111010101",
  54049=>"101111010",
  54050=>"101110111",
  54051=>"101010010",
  54052=>"111001100",
  54053=>"100100000",
  54054=>"110110000",
  54055=>"100011111",
  54056=>"011100000",
  54057=>"111011100",
  54058=>"010000001",
  54059=>"111100001",
  54060=>"000000111",
  54061=>"000101110",
  54062=>"000000111",
  54063=>"100110011",
  54064=>"011011001",
  54065=>"101000101",
  54066=>"000000100",
  54067=>"100111011",
  54068=>"101100000",
  54069=>"110000001",
  54070=>"110101100",
  54071=>"101111111",
  54072=>"110000000",
  54073=>"000000101",
  54074=>"111000000",
  54075=>"011110001",
  54076=>"001101011",
  54077=>"000100101",
  54078=>"100100000",
  54079=>"100010010",
  54080=>"111101101",
  54081=>"101010010",
  54082=>"001101100",
  54083=>"100000011",
  54084=>"011001111",
  54085=>"101011111",
  54086=>"110011111",
  54087=>"001111001",
  54088=>"000011100",
  54089=>"100111101",
  54090=>"111111001",
  54091=>"110100000",
  54092=>"101001011",
  54093=>"011100110",
  54094=>"000010000",
  54095=>"111000100",
  54096=>"101000100",
  54097=>"010000100",
  54098=>"010110100",
  54099=>"001111110",
  54100=>"010110101",
  54101=>"100001111",
  54102=>"101100011",
  54103=>"111100111",
  54104=>"101001001",
  54105=>"001000010",
  54106=>"000111111",
  54107=>"000111101",
  54108=>"010000000",
  54109=>"011010111",
  54110=>"001010111",
  54111=>"000110010",
  54112=>"001100100",
  54113=>"111100100",
  54114=>"111011111",
  54115=>"110000111",
  54116=>"001100010",
  54117=>"101111000",
  54118=>"110011000",
  54119=>"111000110",
  54120=>"010100011",
  54121=>"110010011",
  54122=>"111101000",
  54123=>"010111011",
  54124=>"010001010",
  54125=>"100111100",
  54126=>"110100111",
  54127=>"100010001",
  54128=>"001100010",
  54129=>"101011011",
  54130=>"010011110",
  54131=>"001100100",
  54132=>"001000101",
  54133=>"110111111",
  54134=>"000100001",
  54135=>"001000010",
  54136=>"001100000",
  54137=>"011101010",
  54138=>"000101110",
  54139=>"001000001",
  54140=>"011111001",
  54141=>"101001100",
  54142=>"000000101",
  54143=>"010110010",
  54144=>"100000101",
  54145=>"010100100",
  54146=>"001001011",
  54147=>"011100011",
  54148=>"010000111",
  54149=>"101010010",
  54150=>"100011011",
  54151=>"001100000",
  54152=>"000111100",
  54153=>"000100010",
  54154=>"010000000",
  54155=>"111011111",
  54156=>"000110010",
  54157=>"000101010",
  54158=>"010001111",
  54159=>"010100010",
  54160=>"110100111",
  54161=>"100110011",
  54162=>"100110111",
  54163=>"010111010",
  54164=>"000000001",
  54165=>"101000010",
  54166=>"000110010",
  54167=>"011000000",
  54168=>"010010111",
  54169=>"000010111",
  54170=>"110110110",
  54171=>"011111010",
  54172=>"110011111",
  54173=>"100111101",
  54174=>"111000101",
  54175=>"000111010",
  54176=>"101111101",
  54177=>"100101100",
  54178=>"100110111",
  54179=>"110001111",
  54180=>"110110000",
  54181=>"101000010",
  54182=>"111001010",
  54183=>"110100100",
  54184=>"010100111",
  54185=>"001011000",
  54186=>"001000101",
  54187=>"101101000",
  54188=>"100100010",
  54189=>"100101110",
  54190=>"111101001",
  54191=>"000101100",
  54192=>"000000001",
  54193=>"000111111",
  54194=>"011000000",
  54195=>"100000001",
  54196=>"100001011",
  54197=>"011001101",
  54198=>"011001100",
  54199=>"011001110",
  54200=>"100100100",
  54201=>"100111010",
  54202=>"101010100",
  54203=>"101111010",
  54204=>"011011100",
  54205=>"000010110",
  54206=>"011000000",
  54207=>"100101000",
  54208=>"000001111",
  54209=>"110010011",
  54210=>"100111100",
  54211=>"101111000",
  54212=>"110001111",
  54213=>"101011000",
  54214=>"111110011",
  54215=>"010001110",
  54216=>"110000100",
  54217=>"001001100",
  54218=>"011001010",
  54219=>"101001000",
  54220=>"010101110",
  54221=>"001011011",
  54222=>"111110110",
  54223=>"001000100",
  54224=>"101110110",
  54225=>"011000000",
  54226=>"000110000",
  54227=>"111010110",
  54228=>"001001001",
  54229=>"110010000",
  54230=>"010101101",
  54231=>"111110101",
  54232=>"111110111",
  54233=>"111101110",
  54234=>"111110110",
  54235=>"000000011",
  54236=>"000100100",
  54237=>"000111000",
  54238=>"100001100",
  54239=>"110110010",
  54240=>"011101111",
  54241=>"011000001",
  54242=>"000000000",
  54243=>"101010100",
  54244=>"010110110",
  54245=>"111010100",
  54246=>"010001111",
  54247=>"000111000",
  54248=>"001010000",
  54249=>"011011111",
  54250=>"010101000",
  54251=>"100000111",
  54252=>"010011100",
  54253=>"000011101",
  54254=>"011010110",
  54255=>"010101101",
  54256=>"001101111",
  54257=>"000010001",
  54258=>"011001111",
  54259=>"111011010",
  54260=>"000111101",
  54261=>"100100110",
  54262=>"110011101",
  54263=>"101101011",
  54264=>"111001100",
  54265=>"001100101",
  54266=>"101111010",
  54267=>"010111010",
  54268=>"110110111",
  54269=>"000000010",
  54270=>"001001000",
  54271=>"010001111",
  54272=>"001010010",
  54273=>"100100111",
  54274=>"011111101",
  54275=>"111011001",
  54276=>"100101011",
  54277=>"110000010",
  54278=>"111100010",
  54279=>"010101001",
  54280=>"101000110",
  54281=>"110101000",
  54282=>"101100010",
  54283=>"111000110",
  54284=>"101010011",
  54285=>"011010010",
  54286=>"010100011",
  54287=>"001001011",
  54288=>"101100010",
  54289=>"101001000",
  54290=>"101110111",
  54291=>"011101110",
  54292=>"111111100",
  54293=>"000001001",
  54294=>"111110111",
  54295=>"000000101",
  54296=>"111110101",
  54297=>"011110000",
  54298=>"111100010",
  54299=>"011000010",
  54300=>"111110100",
  54301=>"000000011",
  54302=>"111010100",
  54303=>"010011011",
  54304=>"101001111",
  54305=>"011010110",
  54306=>"111011000",
  54307=>"000001011",
  54308=>"111000001",
  54309=>"011100000",
  54310=>"110111001",
  54311=>"111001101",
  54312=>"010001110",
  54313=>"001011001",
  54314=>"101111101",
  54315=>"110110101",
  54316=>"101011110",
  54317=>"101000000",
  54318=>"001010101",
  54319=>"110000011",
  54320=>"111101010",
  54321=>"001001000",
  54322=>"001011000",
  54323=>"101100010",
  54324=>"111001110",
  54325=>"000000010",
  54326=>"001000010",
  54327=>"110110010",
  54328=>"000011110",
  54329=>"101010010",
  54330=>"001110001",
  54331=>"011110000",
  54332=>"111110011",
  54333=>"111101111",
  54334=>"101000001",
  54335=>"101001010",
  54336=>"000111001",
  54337=>"111101010",
  54338=>"100101101",
  54339=>"101010000",
  54340=>"000110000",
  54341=>"111101001",
  54342=>"011011000",
  54343=>"010010110",
  54344=>"001000010",
  54345=>"111111111",
  54346=>"011110000",
  54347=>"100011111",
  54348=>"001110001",
  54349=>"000000110",
  54350=>"001001000",
  54351=>"001100000",
  54352=>"111011111",
  54353=>"000101000",
  54354=>"100000101",
  54355=>"011000100",
  54356=>"001000110",
  54357=>"000110010",
  54358=>"011001110",
  54359=>"100110100",
  54360=>"101111100",
  54361=>"111010101",
  54362=>"000000100",
  54363=>"001111000",
  54364=>"011010000",
  54365=>"100000000",
  54366=>"110001100",
  54367=>"011111110",
  54368=>"010111000",
  54369=>"110000010",
  54370=>"001101101",
  54371=>"000100001",
  54372=>"100010111",
  54373=>"111101111",
  54374=>"101010110",
  54375=>"111111011",
  54376=>"000011111",
  54377=>"111011100",
  54378=>"001011011",
  54379=>"111001101",
  54380=>"101011010",
  54381=>"110000010",
  54382=>"011111011",
  54383=>"010000101",
  54384=>"011110001",
  54385=>"000100101",
  54386=>"011110011",
  54387=>"110000001",
  54388=>"000110001",
  54389=>"101101100",
  54390=>"000111110",
  54391=>"101111100",
  54392=>"111111100",
  54393=>"111001011",
  54394=>"000100011",
  54395=>"100001010",
  54396=>"111001111",
  54397=>"111001011",
  54398=>"111010011",
  54399=>"111111100",
  54400=>"001011101",
  54401=>"110010001",
  54402=>"101111111",
  54403=>"001011101",
  54404=>"001111000",
  54405=>"011000111",
  54406=>"110010110",
  54407=>"000001110",
  54408=>"100011111",
  54409=>"111100100",
  54410=>"011001001",
  54411=>"000011110",
  54412=>"010110111",
  54413=>"101101111",
  54414=>"110000100",
  54415=>"001011010",
  54416=>"100101000",
  54417=>"110100001",
  54418=>"101010110",
  54419=>"101011101",
  54420=>"011101000",
  54421=>"001010000",
  54422=>"110110010",
  54423=>"011010011",
  54424=>"000011001",
  54425=>"101111111",
  54426=>"100000100",
  54427=>"001110100",
  54428=>"000000010",
  54429=>"111001000",
  54430=>"111111100",
  54431=>"011000100",
  54432=>"010001001",
  54433=>"010101100",
  54434=>"011100000",
  54435=>"101000000",
  54436=>"011011100",
  54437=>"010110010",
  54438=>"101011011",
  54439=>"101101001",
  54440=>"010111101",
  54441=>"110000110",
  54442=>"000001111",
  54443=>"100000100",
  54444=>"111110001",
  54445=>"001111000",
  54446=>"101101111",
  54447=>"011111100",
  54448=>"011111111",
  54449=>"111111111",
  54450=>"110101010",
  54451=>"000000000",
  54452=>"101011101",
  54453=>"011111111",
  54454=>"100001100",
  54455=>"111111100",
  54456=>"111000000",
  54457=>"101000000",
  54458=>"000000100",
  54459=>"000110100",
  54460=>"011011000",
  54461=>"011100111",
  54462=>"000000000",
  54463=>"010110000",
  54464=>"111010100",
  54465=>"011101100",
  54466=>"011000011",
  54467=>"101000101",
  54468=>"100101101",
  54469=>"010011011",
  54470=>"101000100",
  54471=>"111101110",
  54472=>"110101111",
  54473=>"101010100",
  54474=>"010010000",
  54475=>"100111001",
  54476=>"001100011",
  54477=>"110111011",
  54478=>"111110111",
  54479=>"110010001",
  54480=>"100010011",
  54481=>"001111001",
  54482=>"000011101",
  54483=>"000110011",
  54484=>"000010101",
  54485=>"110000010",
  54486=>"011011011",
  54487=>"010000000",
  54488=>"100110100",
  54489=>"000110110",
  54490=>"101000011",
  54491=>"000000100",
  54492=>"000000000",
  54493=>"110101010",
  54494=>"100001001",
  54495=>"010110101",
  54496=>"011001001",
  54497=>"010010001",
  54498=>"000001011",
  54499=>"010000101",
  54500=>"000010101",
  54501=>"110010001",
  54502=>"001000011",
  54503=>"000011000",
  54504=>"110000100",
  54505=>"110000000",
  54506=>"111100010",
  54507=>"100000111",
  54508=>"100100110",
  54509=>"010010001",
  54510=>"111101100",
  54511=>"011100000",
  54512=>"000000111",
  54513=>"110111011",
  54514=>"110100111",
  54515=>"011111100",
  54516=>"010110000",
  54517=>"111110100",
  54518=>"100001001",
  54519=>"011000010",
  54520=>"101010011",
  54521=>"101111111",
  54522=>"110010000",
  54523=>"110111001",
  54524=>"111101111",
  54525=>"111010100",
  54526=>"101011110",
  54527=>"001010100",
  54528=>"100101001",
  54529=>"111010101",
  54530=>"111101101",
  54531=>"110011101",
  54532=>"100010101",
  54533=>"100110110",
  54534=>"010010101",
  54535=>"010000000",
  54536=>"101101111",
  54537=>"101111110",
  54538=>"111110110",
  54539=>"001011001",
  54540=>"101110001",
  54541=>"101100010",
  54542=>"111000111",
  54543=>"111110010",
  54544=>"001010010",
  54545=>"100110010",
  54546=>"010000010",
  54547=>"000010000",
  54548=>"001000011",
  54549=>"101010000",
  54550=>"001111001",
  54551=>"111100100",
  54552=>"100000000",
  54553=>"010010111",
  54554=>"010001001",
  54555=>"100011000",
  54556=>"000001101",
  54557=>"011001011",
  54558=>"100111010",
  54559=>"101100000",
  54560=>"010010010",
  54561=>"100100010",
  54562=>"110110011",
  54563=>"101101001",
  54564=>"011111111",
  54565=>"111001001",
  54566=>"001101011",
  54567=>"101101011",
  54568=>"000010011",
  54569=>"011111101",
  54570=>"100001011",
  54571=>"101100001",
  54572=>"100101001",
  54573=>"101111011",
  54574=>"111111111",
  54575=>"111011100",
  54576=>"111101010",
  54577=>"000010011",
  54578=>"101110101",
  54579=>"101110001",
  54580=>"011001010",
  54581=>"110000000",
  54582=>"001011011",
  54583=>"101001010",
  54584=>"000001010",
  54585=>"101110100",
  54586=>"011110100",
  54587=>"100101001",
  54588=>"111010011",
  54589=>"000001001",
  54590=>"010110011",
  54591=>"010111101",
  54592=>"100110111",
  54593=>"111101100",
  54594=>"110111111",
  54595=>"101001111",
  54596=>"010010000",
  54597=>"101100111",
  54598=>"000100100",
  54599=>"110000001",
  54600=>"111111111",
  54601=>"100000001",
  54602=>"000000100",
  54603=>"110101100",
  54604=>"010100100",
  54605=>"001100000",
  54606=>"010111100",
  54607=>"100101100",
  54608=>"010011011",
  54609=>"010001110",
  54610=>"000100111",
  54611=>"111100000",
  54612=>"010010000",
  54613=>"111000100",
  54614=>"110110110",
  54615=>"010101100",
  54616=>"101100101",
  54617=>"010010110",
  54618=>"010110110",
  54619=>"000100000",
  54620=>"101001001",
  54621=>"100011001",
  54622=>"111001110",
  54623=>"110001100",
  54624=>"110000110",
  54625=>"101110011",
  54626=>"100101000",
  54627=>"000010000",
  54628=>"000000010",
  54629=>"110011110",
  54630=>"110110010",
  54631=>"101110000",
  54632=>"001111010",
  54633=>"100100001",
  54634=>"111001001",
  54635=>"101110011",
  54636=>"111111010",
  54637=>"101000110",
  54638=>"101000000",
  54639=>"101011010",
  54640=>"110110000",
  54641=>"111001101",
  54642=>"100110100",
  54643=>"001111011",
  54644=>"111110111",
  54645=>"001100000",
  54646=>"110100101",
  54647=>"100010101",
  54648=>"100000001",
  54649=>"101100101",
  54650=>"110111111",
  54651=>"101001100",
  54652=>"000101111",
  54653=>"010011000",
  54654=>"101111001",
  54655=>"011010111",
  54656=>"100101010",
  54657=>"010001001",
  54658=>"110111101",
  54659=>"001111000",
  54660=>"110101010",
  54661=>"110111110",
  54662=>"101011010",
  54663=>"001111111",
  54664=>"010010000",
  54665=>"000111000",
  54666=>"110010101",
  54667=>"111111010",
  54668=>"101100100",
  54669=>"011010011",
  54670=>"111001010",
  54671=>"101100100",
  54672=>"011000000",
  54673=>"000100111",
  54674=>"010100100",
  54675=>"000000110",
  54676=>"111001110",
  54677=>"001010101",
  54678=>"000000111",
  54679=>"101010111",
  54680=>"000101001",
  54681=>"010100001",
  54682=>"111010111",
  54683=>"000110001",
  54684=>"000100000",
  54685=>"000110111",
  54686=>"101001111",
  54687=>"000010010",
  54688=>"010010010",
  54689=>"111010101",
  54690=>"110101101",
  54691=>"100000000",
  54692=>"010011011",
  54693=>"000000101",
  54694=>"010011010",
  54695=>"111111110",
  54696=>"001111000",
  54697=>"000110110",
  54698=>"100111111",
  54699=>"000000100",
  54700=>"011011010",
  54701=>"110100001",
  54702=>"110000001",
  54703=>"001010100",
  54704=>"110000001",
  54705=>"001001000",
  54706=>"111111001",
  54707=>"011010011",
  54708=>"100110010",
  54709=>"001110110",
  54710=>"111010000",
  54711=>"101100101",
  54712=>"000110010",
  54713=>"100000101",
  54714=>"011010011",
  54715=>"001110010",
  54716=>"100101111",
  54717=>"000000001",
  54718=>"100001001",
  54719=>"000101101",
  54720=>"001001110",
  54721=>"000001110",
  54722=>"111010101",
  54723=>"001110110",
  54724=>"101110000",
  54725=>"000110001",
  54726=>"100110101",
  54727=>"101011010",
  54728=>"110010100",
  54729=>"101111110",
  54730=>"101011001",
  54731=>"111111111",
  54732=>"111111000",
  54733=>"011000010",
  54734=>"110111000",
  54735=>"000001110",
  54736=>"100100110",
  54737=>"010000001",
  54738=>"011111111",
  54739=>"110011110",
  54740=>"100001001",
  54741=>"001000001",
  54742=>"110010111",
  54743=>"101110110",
  54744=>"001010100",
  54745=>"010000010",
  54746=>"010100110",
  54747=>"111000011",
  54748=>"001101110",
  54749=>"110001001",
  54750=>"101100000",
  54751=>"001010100",
  54752=>"000110100",
  54753=>"011011111",
  54754=>"010111000",
  54755=>"110001010",
  54756=>"000110011",
  54757=>"000110000",
  54758=>"101000000",
  54759=>"101010000",
  54760=>"100111111",
  54761=>"111000100",
  54762=>"011010011",
  54763=>"101000001",
  54764=>"110111011",
  54765=>"101100001",
  54766=>"101111010",
  54767=>"110011000",
  54768=>"111111001",
  54769=>"011001001",
  54770=>"100010011",
  54771=>"010111100",
  54772=>"101110000",
  54773=>"000000000",
  54774=>"011011000",
  54775=>"111100001",
  54776=>"110101101",
  54777=>"100111011",
  54778=>"001101010",
  54779=>"000010010",
  54780=>"111100111",
  54781=>"001101111",
  54782=>"101111111",
  54783=>"111010100",
  54784=>"001111110",
  54785=>"110010011",
  54786=>"110101100",
  54787=>"100101101",
  54788=>"100010001",
  54789=>"111000000",
  54790=>"000101001",
  54791=>"011011111",
  54792=>"011100100",
  54793=>"111110100",
  54794=>"100010011",
  54795=>"000000000",
  54796=>"001111100",
  54797=>"010100000",
  54798=>"001010100",
  54799=>"110100000",
  54800=>"111110011",
  54801=>"000111111",
  54802=>"011000111",
  54803=>"010010111",
  54804=>"000001000",
  54805=>"010010000",
  54806=>"111011001",
  54807=>"001001011",
  54808=>"001000110",
  54809=>"110110010",
  54810=>"110111101",
  54811=>"011101111",
  54812=>"011110011",
  54813=>"100100100",
  54814=>"011010010",
  54815=>"101101010",
  54816=>"110000010",
  54817=>"011001011",
  54818=>"111001000",
  54819=>"110011000",
  54820=>"110001010",
  54821=>"001011110",
  54822=>"110000011",
  54823=>"000000010",
  54824=>"010001000",
  54825=>"000011001",
  54826=>"100001101",
  54827=>"000110000",
  54828=>"111001001",
  54829=>"011100011",
  54830=>"001111111",
  54831=>"111011101",
  54832=>"100111010",
  54833=>"101101001",
  54834=>"010100111",
  54835=>"001010000",
  54836=>"000000101",
  54837=>"111100000",
  54838=>"001010111",
  54839=>"000110000",
  54840=>"101111011",
  54841=>"001010000",
  54842=>"111001101",
  54843=>"000000111",
  54844=>"110001000",
  54845=>"000111001",
  54846=>"011100100",
  54847=>"000000010",
  54848=>"111010001",
  54849=>"111111111",
  54850=>"100001101",
  54851=>"111011101",
  54852=>"010101101",
  54853=>"010010100",
  54854=>"001001110",
  54855=>"000100100",
  54856=>"111100010",
  54857=>"100110111",
  54858=>"100101100",
  54859=>"101000011",
  54860=>"111011100",
  54861=>"000011000",
  54862=>"001001111",
  54863=>"100100001",
  54864=>"010111000",
  54865=>"000000110",
  54866=>"001000011",
  54867=>"000000000",
  54868=>"010011110",
  54869=>"000011010",
  54870=>"100100011",
  54871=>"100101011",
  54872=>"100001111",
  54873=>"101101011",
  54874=>"010011111",
  54875=>"011010111",
  54876=>"000000101",
  54877=>"101001010",
  54878=>"101100001",
  54879=>"111011010",
  54880=>"110001110",
  54881=>"100001001",
  54882=>"111110000",
  54883=>"000001101",
  54884=>"101011001",
  54885=>"001000010",
  54886=>"110110100",
  54887=>"100001110",
  54888=>"111100111",
  54889=>"010110100",
  54890=>"000101010",
  54891=>"011111010",
  54892=>"001000000",
  54893=>"110001101",
  54894=>"011110001",
  54895=>"100011110",
  54896=>"001000100",
  54897=>"000000101",
  54898=>"001100001",
  54899=>"001000011",
  54900=>"100111000",
  54901=>"000101000",
  54902=>"111111101",
  54903=>"111101011",
  54904=>"100100000",
  54905=>"010010100",
  54906=>"001000000",
  54907=>"010000000",
  54908=>"010100000",
  54909=>"101111101",
  54910=>"101011010",
  54911=>"010100010",
  54912=>"000111011",
  54913=>"101110111",
  54914=>"000001001",
  54915=>"100011000",
  54916=>"100001111",
  54917=>"000101110",
  54918=>"100001001",
  54919=>"110100111",
  54920=>"000001110",
  54921=>"010101011",
  54922=>"110101000",
  54923=>"011101000",
  54924=>"010000111",
  54925=>"100011010",
  54926=>"001000001",
  54927=>"000011100",
  54928=>"100010000",
  54929=>"011110000",
  54930=>"101100101",
  54931=>"100000000",
  54932=>"000100011",
  54933=>"100111111",
  54934=>"000001001",
  54935=>"100110100",
  54936=>"001010110",
  54937=>"001010010",
  54938=>"000011110",
  54939=>"100010000",
  54940=>"000010000",
  54941=>"100110010",
  54942=>"111010011",
  54943=>"110011100",
  54944=>"111110111",
  54945=>"011011010",
  54946=>"001001101",
  54947=>"011111110",
  54948=>"111010000",
  54949=>"111110000",
  54950=>"111101110",
  54951=>"001010101",
  54952=>"101110100",
  54953=>"000100010",
  54954=>"110100000",
  54955=>"100010000",
  54956=>"110001000",
  54957=>"110010110",
  54958=>"001011110",
  54959=>"111111011",
  54960=>"001001110",
  54961=>"000010001",
  54962=>"000111000",
  54963=>"000100111",
  54964=>"010011000",
  54965=>"011001001",
  54966=>"010100001",
  54967=>"011001001",
  54968=>"011111000",
  54969=>"000010000",
  54970=>"111101100",
  54971=>"011010000",
  54972=>"010001101",
  54973=>"100011011",
  54974=>"101011011",
  54975=>"000101111",
  54976=>"010110000",
  54977=>"110111110",
  54978=>"110100101",
  54979=>"101001000",
  54980=>"011111110",
  54981=>"111010001",
  54982=>"011100111",
  54983=>"111010111",
  54984=>"000000011",
  54985=>"110101000",
  54986=>"010001101",
  54987=>"001010100",
  54988=>"101101111",
  54989=>"000110100",
  54990=>"111010000",
  54991=>"111111000",
  54992=>"001110101",
  54993=>"001011101",
  54994=>"001111010",
  54995=>"100000000",
  54996=>"000010010",
  54997=>"010111001",
  54998=>"111001111",
  54999=>"011001001",
  55000=>"100010110",
  55001=>"011010101",
  55002=>"111110110",
  55003=>"101001101",
  55004=>"100100000",
  55005=>"101101101",
  55006=>"000011101",
  55007=>"001111111",
  55008=>"101100001",
  55009=>"110100010",
  55010=>"011001010",
  55011=>"111011010",
  55012=>"010000000",
  55013=>"001011010",
  55014=>"011111010",
  55015=>"001010110",
  55016=>"001110101",
  55017=>"111110011",
  55018=>"111011100",
  55019=>"000100000",
  55020=>"011100001",
  55021=>"110010110",
  55022=>"011100111",
  55023=>"110000010",
  55024=>"101011001",
  55025=>"100111110",
  55026=>"111011101",
  55027=>"101011000",
  55028=>"111110011",
  55029=>"011001111",
  55030=>"101000100",
  55031=>"100111100",
  55032=>"100001011",
  55033=>"101110101",
  55034=>"000000110",
  55035=>"000101010",
  55036=>"111011001",
  55037=>"100010001",
  55038=>"000111110",
  55039=>"010001010",
  55040=>"010101011",
  55041=>"010101000",
  55042=>"011010001",
  55043=>"000000000",
  55044=>"110110110",
  55045=>"001000100",
  55046=>"001110001",
  55047=>"000101111",
  55048=>"011100001",
  55049=>"111111101",
  55050=>"001001011",
  55051=>"011010110",
  55052=>"001100000",
  55053=>"001101111",
  55054=>"101111011",
  55055=>"100001001",
  55056=>"010101001",
  55057=>"010110100",
  55058=>"000101010",
  55059=>"010100100",
  55060=>"111000011",
  55061=>"110111010",
  55062=>"010000101",
  55063=>"111011111",
  55064=>"000010000",
  55065=>"100000010",
  55066=>"000100100",
  55067=>"011011101",
  55068=>"001011000",
  55069=>"000110111",
  55070=>"001000001",
  55071=>"100010110",
  55072=>"100011010",
  55073=>"110110001",
  55074=>"101001101",
  55075=>"110000000",
  55076=>"000011011",
  55077=>"101101111",
  55078=>"110100100",
  55079=>"000100010",
  55080=>"011010110",
  55081=>"001000000",
  55082=>"110001100",
  55083=>"110111110",
  55084=>"111000110",
  55085=>"111111110",
  55086=>"110101001",
  55087=>"011011111",
  55088=>"000001110",
  55089=>"101110010",
  55090=>"001011110",
  55091=>"000011100",
  55092=>"100101111",
  55093=>"000101011",
  55094=>"110000001",
  55095=>"100011001",
  55096=>"101001100",
  55097=>"001000100",
  55098=>"101000011",
  55099=>"110010101",
  55100=>"111000000",
  55101=>"011010011",
  55102=>"000010000",
  55103=>"100111010",
  55104=>"010000111",
  55105=>"111100100",
  55106=>"110101110",
  55107=>"100010011",
  55108=>"010000000",
  55109=>"000111110",
  55110=>"011010111",
  55111=>"010100010",
  55112=>"011001111",
  55113=>"000010011",
  55114=>"110110111",
  55115=>"100100001",
  55116=>"000111011",
  55117=>"000011000",
  55118=>"010001000",
  55119=>"111001100",
  55120=>"011010001",
  55121=>"001111111",
  55122=>"111111000",
  55123=>"110011110",
  55124=>"101100000",
  55125=>"001111111",
  55126=>"011011110",
  55127=>"001110100",
  55128=>"111101111",
  55129=>"110000011",
  55130=>"111001011",
  55131=>"000101000",
  55132=>"001110001",
  55133=>"001000100",
  55134=>"010011011",
  55135=>"010001101",
  55136=>"101010011",
  55137=>"011011110",
  55138=>"100000010",
  55139=>"111111100",
  55140=>"000111001",
  55141=>"001011100",
  55142=>"101011111",
  55143=>"001101101",
  55144=>"101001001",
  55145=>"000001000",
  55146=>"111101000",
  55147=>"010111000",
  55148=>"010011001",
  55149=>"000000010",
  55150=>"011000000",
  55151=>"011100100",
  55152=>"010011100",
  55153=>"111011111",
  55154=>"100011100",
  55155=>"111101010",
  55156=>"110010111",
  55157=>"000000001",
  55158=>"001111011",
  55159=>"100111111",
  55160=>"101101110",
  55161=>"010101100",
  55162=>"011000100",
  55163=>"011000010",
  55164=>"011011111",
  55165=>"010101000",
  55166=>"000111100",
  55167=>"100111001",
  55168=>"111010010",
  55169=>"010011111",
  55170=>"101100010",
  55171=>"010001111",
  55172=>"000000110",
  55173=>"111100100",
  55174=>"000001100",
  55175=>"101011110",
  55176=>"110101010",
  55177=>"000111111",
  55178=>"111001001",
  55179=>"011111101",
  55180=>"011000010",
  55181=>"011110111",
  55182=>"001000111",
  55183=>"011001101",
  55184=>"011000100",
  55185=>"000101111",
  55186=>"101011011",
  55187=>"111110110",
  55188=>"010100100",
  55189=>"011010001",
  55190=>"011111100",
  55191=>"000000100",
  55192=>"110000010",
  55193=>"111111011",
  55194=>"101001000",
  55195=>"010110010",
  55196=>"001100000",
  55197=>"100100000",
  55198=>"000011100",
  55199=>"010110011",
  55200=>"101011001",
  55201=>"000011001",
  55202=>"001111110",
  55203=>"000000100",
  55204=>"001110000",
  55205=>"111101010",
  55206=>"110000101",
  55207=>"100000111",
  55208=>"010110010",
  55209=>"100011010",
  55210=>"110100101",
  55211=>"000010110",
  55212=>"001001100",
  55213=>"000110111",
  55214=>"010111011",
  55215=>"101000010",
  55216=>"111000110",
  55217=>"001111111",
  55218=>"110101100",
  55219=>"100011001",
  55220=>"100101111",
  55221=>"110100011",
  55222=>"011010100",
  55223=>"010110010",
  55224=>"000101001",
  55225=>"111010001",
  55226=>"010010010",
  55227=>"111010010",
  55228=>"011101110",
  55229=>"010100111",
  55230=>"010110110",
  55231=>"000000100",
  55232=>"000001110",
  55233=>"110010111",
  55234=>"010111110",
  55235=>"000101100",
  55236=>"110101111",
  55237=>"010100001",
  55238=>"010011100",
  55239=>"100101100",
  55240=>"100000010",
  55241=>"100001111",
  55242=>"110110111",
  55243=>"111001110",
  55244=>"101110100",
  55245=>"011010100",
  55246=>"000001000",
  55247=>"001011011",
  55248=>"011001000",
  55249=>"111100110",
  55250=>"111110010",
  55251=>"011100100",
  55252=>"111001100",
  55253=>"001010010",
  55254=>"110000110",
  55255=>"111100111",
  55256=>"000001111",
  55257=>"000100100",
  55258=>"100101010",
  55259=>"101000011",
  55260=>"110101110",
  55261=>"001101101",
  55262=>"111111111",
  55263=>"110010110",
  55264=>"101010100",
  55265=>"110110001",
  55266=>"011111110",
  55267=>"110111110",
  55268=>"100010100",
  55269=>"010010101",
  55270=>"011000000",
  55271=>"001001001",
  55272=>"110100010",
  55273=>"000000011",
  55274=>"110000110",
  55275=>"000010001",
  55276=>"000111010",
  55277=>"001000001",
  55278=>"011001000",
  55279=>"101100011",
  55280=>"111101101",
  55281=>"010001110",
  55282=>"101011010",
  55283=>"000000101",
  55284=>"111101111",
  55285=>"100000110",
  55286=>"110000000",
  55287=>"000010111",
  55288=>"001000101",
  55289=>"110100111",
  55290=>"001111111",
  55291=>"101110100",
  55292=>"111111100",
  55293=>"101100000",
  55294=>"011110000",
  55295=>"010111100",
  55296=>"101111111",
  55297=>"001101000",
  55298=>"111111110",
  55299=>"101111101",
  55300=>"010100110",
  55301=>"111001101",
  55302=>"010011100",
  55303=>"100000000",
  55304=>"010011110",
  55305=>"100100011",
  55306=>"100010100",
  55307=>"011101000",
  55308=>"001010110",
  55309=>"111001000",
  55310=>"001100011",
  55311=>"110110000",
  55312=>"001100000",
  55313=>"101010100",
  55314=>"001111101",
  55315=>"001010010",
  55316=>"001111111",
  55317=>"111110101",
  55318=>"000110110",
  55319=>"111000001",
  55320=>"011110011",
  55321=>"100011010",
  55322=>"111001011",
  55323=>"011011000",
  55324=>"100011000",
  55325=>"010011110",
  55326=>"110110000",
  55327=>"001101101",
  55328=>"011100000",
  55329=>"001111101",
  55330=>"110010100",
  55331=>"101011011",
  55332=>"111110101",
  55333=>"010101011",
  55334=>"100001110",
  55335=>"111111001",
  55336=>"011010010",
  55337=>"101110110",
  55338=>"010110111",
  55339=>"101111111",
  55340=>"010011001",
  55341=>"001110001",
  55342=>"011101100",
  55343=>"011101101",
  55344=>"000010011",
  55345=>"110110010",
  55346=>"001000010",
  55347=>"011000001",
  55348=>"111000100",
  55349=>"111011001",
  55350=>"001100101",
  55351=>"011001101",
  55352=>"101111111",
  55353=>"000010011",
  55354=>"010011011",
  55355=>"110110111",
  55356=>"000100010",
  55357=>"111001000",
  55358=>"110011010",
  55359=>"001001100",
  55360=>"100100110",
  55361=>"100010010",
  55362=>"100111111",
  55363=>"101110010",
  55364=>"001001000",
  55365=>"000110011",
  55366=>"101011001",
  55367=>"011011011",
  55368=>"010100110",
  55369=>"111000101",
  55370=>"100111100",
  55371=>"010011010",
  55372=>"111101001",
  55373=>"000010000",
  55374=>"110000001",
  55375=>"011100010",
  55376=>"101111010",
  55377=>"011010111",
  55378=>"110001000",
  55379=>"001100000",
  55380=>"100111110",
  55381=>"000000010",
  55382=>"011100111",
  55383=>"101110000",
  55384=>"000011110",
  55385=>"101111101",
  55386=>"010101111",
  55387=>"110001100",
  55388=>"001010010",
  55389=>"000000101",
  55390=>"011011110",
  55391=>"100100101",
  55392=>"001000101",
  55393=>"100110001",
  55394=>"111110010",
  55395=>"000010011",
  55396=>"000000000",
  55397=>"100001100",
  55398=>"011101110",
  55399=>"110110111",
  55400=>"001010010",
  55401=>"001100011",
  55402=>"100011001",
  55403=>"101100101",
  55404=>"110011110",
  55405=>"001000000",
  55406=>"000011001",
  55407=>"010101111",
  55408=>"001011011",
  55409=>"101110010",
  55410=>"110010000",
  55411=>"001010110",
  55412=>"101100001",
  55413=>"100111000",
  55414=>"111100010",
  55415=>"100101111",
  55416=>"111011001",
  55417=>"001101101",
  55418=>"110101111",
  55419=>"101111010",
  55420=>"000000111",
  55421=>"101010000",
  55422=>"000000100",
  55423=>"111111111",
  55424=>"111111110",
  55425=>"001000110",
  55426=>"010100110",
  55427=>"001011010",
  55428=>"101001110",
  55429=>"001111011",
  55430=>"011011001",
  55431=>"110100001",
  55432=>"000000010",
  55433=>"010001101",
  55434=>"000001100",
  55435=>"001111000",
  55436=>"111011101",
  55437=>"000100011",
  55438=>"101100000",
  55439=>"001010101",
  55440=>"101011110",
  55441=>"011010011",
  55442=>"011110000",
  55443=>"100011100",
  55444=>"100111111",
  55445=>"111101101",
  55446=>"001111111",
  55447=>"110001010",
  55448=>"000100111",
  55449=>"100011000",
  55450=>"001011001",
  55451=>"011010110",
  55452=>"000010001",
  55453=>"100110010",
  55454=>"001000110",
  55455=>"011110110",
  55456=>"011100001",
  55457=>"101101111",
  55458=>"000000001",
  55459=>"101100001",
  55460=>"000100110",
  55461=>"000011110",
  55462=>"110101001",
  55463=>"000001001",
  55464=>"101000011",
  55465=>"110110000",
  55466=>"100011110",
  55467=>"000011000",
  55468=>"000001110",
  55469=>"101011000",
  55470=>"000101011",
  55471=>"110000001",
  55472=>"001010010",
  55473=>"001000010",
  55474=>"011110011",
  55475=>"000000011",
  55476=>"111011110",
  55477=>"101001111",
  55478=>"011101101",
  55479=>"010111010",
  55480=>"101110111",
  55481=>"110011111",
  55482=>"010111110",
  55483=>"010111011",
  55484=>"001011001",
  55485=>"010010001",
  55486=>"010100011",
  55487=>"001111011",
  55488=>"001110010",
  55489=>"000010100",
  55490=>"100100001",
  55491=>"001001100",
  55492=>"000010000",
  55493=>"110110000",
  55494=>"011010110",
  55495=>"010001111",
  55496=>"000011011",
  55497=>"011101111",
  55498=>"111100101",
  55499=>"110010000",
  55500=>"001101100",
  55501=>"111001110",
  55502=>"010100110",
  55503=>"000011000",
  55504=>"101110111",
  55505=>"010010000",
  55506=>"100101010",
  55507=>"011110000",
  55508=>"011010000",
  55509=>"111101000",
  55510=>"010111100",
  55511=>"101111111",
  55512=>"001000100",
  55513=>"110001010",
  55514=>"010000011",
  55515=>"000101000",
  55516=>"011001111",
  55517=>"010100011",
  55518=>"100111000",
  55519=>"011010011",
  55520=>"000110010",
  55521=>"010100010",
  55522=>"001000001",
  55523=>"001010010",
  55524=>"111100101",
  55525=>"011110000",
  55526=>"001010000",
  55527=>"101111010",
  55528=>"111100100",
  55529=>"110111101",
  55530=>"011000000",
  55531=>"011000111",
  55532=>"011001101",
  55533=>"000001110",
  55534=>"000001110",
  55535=>"100000100",
  55536=>"101101110",
  55537=>"001001100",
  55538=>"101101100",
  55539=>"011001000",
  55540=>"011000010",
  55541=>"010001101",
  55542=>"100001110",
  55543=>"000100001",
  55544=>"101010001",
  55545=>"100010110",
  55546=>"010100000",
  55547=>"111000100",
  55548=>"010000010",
  55549=>"010100010",
  55550=>"001101111",
  55551=>"001010111",
  55552=>"011100000",
  55553=>"000101101",
  55554=>"000010111",
  55555=>"101111111",
  55556=>"111011010",
  55557=>"010101100",
  55558=>"000001111",
  55559=>"000111101",
  55560=>"000010000",
  55561=>"000010000",
  55562=>"000111110",
  55563=>"100000111",
  55564=>"010011100",
  55565=>"011111010",
  55566=>"110001110",
  55567=>"011111000",
  55568=>"101000000",
  55569=>"101101010",
  55570=>"111011011",
  55571=>"111011100",
  55572=>"101011100",
  55573=>"010110111",
  55574=>"011110010",
  55575=>"010001111",
  55576=>"111100001",
  55577=>"110110110",
  55578=>"011101000",
  55579=>"101110110",
  55580=>"001111001",
  55581=>"000001000",
  55582=>"001000010",
  55583=>"111011000",
  55584=>"111001010",
  55585=>"000101010",
  55586=>"011010010",
  55587=>"011110001",
  55588=>"011000010",
  55589=>"000000111",
  55590=>"101101010",
  55591=>"110001110",
  55592=>"111010100",
  55593=>"110101111",
  55594=>"010110110",
  55595=>"100101101",
  55596=>"111011110",
  55597=>"000111011",
  55598=>"110111001",
  55599=>"000110100",
  55600=>"101000000",
  55601=>"010100101",
  55602=>"101000101",
  55603=>"100110101",
  55604=>"101000111",
  55605=>"100101101",
  55606=>"111011011",
  55607=>"101001110",
  55608=>"000001000",
  55609=>"100101111",
  55610=>"100111101",
  55611=>"000000111",
  55612=>"010010011",
  55613=>"010100010",
  55614=>"101111100",
  55615=>"101000000",
  55616=>"111010101",
  55617=>"101101011",
  55618=>"000000101",
  55619=>"011010001",
  55620=>"100011111",
  55621=>"110101100",
  55622=>"011000110",
  55623=>"010011110",
  55624=>"010110000",
  55625=>"000000110",
  55626=>"011011111",
  55627=>"001100100",
  55628=>"010111000",
  55629=>"010111100",
  55630=>"110110101",
  55631=>"100101011",
  55632=>"110000010",
  55633=>"100001011",
  55634=>"101011010",
  55635=>"001111001",
  55636=>"101101001",
  55637=>"111011000",
  55638=>"110100110",
  55639=>"100010111",
  55640=>"011001110",
  55641=>"000010110",
  55642=>"000110110",
  55643=>"111110001",
  55644=>"011111001",
  55645=>"010101111",
  55646=>"011100010",
  55647=>"100111000",
  55648=>"000000000",
  55649=>"000110000",
  55650=>"011010001",
  55651=>"000010101",
  55652=>"110011110",
  55653=>"111001101",
  55654=>"010011001",
  55655=>"110010110",
  55656=>"010111111",
  55657=>"110011111",
  55658=>"001011000",
  55659=>"101010011",
  55660=>"100011110",
  55661=>"110010010",
  55662=>"100000001",
  55663=>"010111100",
  55664=>"100111100",
  55665=>"001010101",
  55666=>"010010010",
  55667=>"011001101",
  55668=>"111111111",
  55669=>"001000010",
  55670=>"100100111",
  55671=>"001001110",
  55672=>"001010011",
  55673=>"101001010",
  55674=>"001111010",
  55675=>"010101100",
  55676=>"110101101",
  55677=>"001110010",
  55678=>"010101010",
  55679=>"100001001",
  55680=>"110100000",
  55681=>"000000000",
  55682=>"011000101",
  55683=>"111011110",
  55684=>"100001110",
  55685=>"011110101",
  55686=>"111000001",
  55687=>"111011010",
  55688=>"000100001",
  55689=>"011111011",
  55690=>"110111011",
  55691=>"010011000",
  55692=>"101110111",
  55693=>"101110000",
  55694=>"000110010",
  55695=>"000010100",
  55696=>"001001101",
  55697=>"101001000",
  55698=>"101101101",
  55699=>"000000000",
  55700=>"001101100",
  55701=>"000010001",
  55702=>"100101010",
  55703=>"001101111",
  55704=>"101110001",
  55705=>"100100011",
  55706=>"011101000",
  55707=>"111100100",
  55708=>"110110000",
  55709=>"110010001",
  55710=>"100100111",
  55711=>"111100101",
  55712=>"010111101",
  55713=>"101001111",
  55714=>"011100101",
  55715=>"000000010",
  55716=>"011111001",
  55717=>"001000000",
  55718=>"101111110",
  55719=>"101101000",
  55720=>"110110100",
  55721=>"101010110",
  55722=>"000100010",
  55723=>"001011101",
  55724=>"001110101",
  55725=>"101000000",
  55726=>"110000011",
  55727=>"110011010",
  55728=>"000101110",
  55729=>"101011101",
  55730=>"000000110",
  55731=>"001000001",
  55732=>"011111001",
  55733=>"010001110",
  55734=>"100110101",
  55735=>"000000110",
  55736=>"000001000",
  55737=>"000111110",
  55738=>"100011110",
  55739=>"010010101",
  55740=>"110110100",
  55741=>"111011110",
  55742=>"010101111",
  55743=>"111000100",
  55744=>"110100100",
  55745=>"000111100",
  55746=>"011111100",
  55747=>"000001100",
  55748=>"101110111",
  55749=>"101111111",
  55750=>"000000111",
  55751=>"001000000",
  55752=>"101000111",
  55753=>"000111100",
  55754=>"011110100",
  55755=>"111110110",
  55756=>"100011110",
  55757=>"010000001",
  55758=>"011010100",
  55759=>"010001010",
  55760=>"010111101",
  55761=>"101111010",
  55762=>"111011000",
  55763=>"100111101",
  55764=>"101100011",
  55765=>"100000001",
  55766=>"101000010",
  55767=>"010110101",
  55768=>"000111000",
  55769=>"000001001",
  55770=>"001001100",
  55771=>"000001101",
  55772=>"111100100",
  55773=>"100111100",
  55774=>"110100000",
  55775=>"001110110",
  55776=>"100101110",
  55777=>"000100110",
  55778=>"111110000",
  55779=>"111000100",
  55780=>"100011101",
  55781=>"101010001",
  55782=>"011000011",
  55783=>"011001101",
  55784=>"101111100",
  55785=>"101101010",
  55786=>"001000011",
  55787=>"001111000",
  55788=>"010011010",
  55789=>"010001001",
  55790=>"110110000",
  55791=>"011110011",
  55792=>"010110001",
  55793=>"010111101",
  55794=>"000111011",
  55795=>"100010010",
  55796=>"010000001",
  55797=>"001100111",
  55798=>"110011111",
  55799=>"111101001",
  55800=>"011010110",
  55801=>"000110101",
  55802=>"110100111",
  55803=>"111100110",
  55804=>"101010101",
  55805=>"110111011",
  55806=>"011011101",
  55807=>"000001001",
  55808=>"010110001",
  55809=>"111100011",
  55810=>"011010001",
  55811=>"111110000",
  55812=>"010010101",
  55813=>"011110110",
  55814=>"111101110",
  55815=>"101101110",
  55816=>"100101001",
  55817=>"000000001",
  55818=>"001111011",
  55819=>"001001010",
  55820=>"000110001",
  55821=>"100000010",
  55822=>"100101000",
  55823=>"111000011",
  55824=>"100110001",
  55825=>"100001110",
  55826=>"011011011",
  55827=>"101101111",
  55828=>"000111000",
  55829=>"111001011",
  55830=>"001001110",
  55831=>"101101001",
  55832=>"001001111",
  55833=>"111110010",
  55834=>"011000001",
  55835=>"001101110",
  55836=>"010010111",
  55837=>"101010011",
  55838=>"000001110",
  55839=>"101110011",
  55840=>"101101001",
  55841=>"000010010",
  55842=>"000001110",
  55843=>"010101001",
  55844=>"010101000",
  55845=>"111011101",
  55846=>"010100011",
  55847=>"000011101",
  55848=>"110010010",
  55849=>"110000100",
  55850=>"001010001",
  55851=>"010011110",
  55852=>"110110101",
  55853=>"101010010",
  55854=>"000101110",
  55855=>"100111011",
  55856=>"001100000",
  55857=>"000010001",
  55858=>"001011110",
  55859=>"001000001",
  55860=>"000101101",
  55861=>"011000001",
  55862=>"001101110",
  55863=>"010101011",
  55864=>"010100100",
  55865=>"111111010",
  55866=>"100000100",
  55867=>"000000000",
  55868=>"111100100",
  55869=>"001000100",
  55870=>"100101110",
  55871=>"010110111",
  55872=>"001110101",
  55873=>"100001100",
  55874=>"011000000",
  55875=>"011000011",
  55876=>"000000001",
  55877=>"110111100",
  55878=>"110000000",
  55879=>"010001111",
  55880=>"010001000",
  55881=>"001100101",
  55882=>"000110111",
  55883=>"100010010",
  55884=>"010101101",
  55885=>"000101000",
  55886=>"000111000",
  55887=>"110100000",
  55888=>"111001101",
  55889=>"111010011",
  55890=>"000100000",
  55891=>"000000011",
  55892=>"011100011",
  55893=>"011000110",
  55894=>"101000111",
  55895=>"110010101",
  55896=>"111111110",
  55897=>"110010011",
  55898=>"000100010",
  55899=>"010011111",
  55900=>"001100000",
  55901=>"000010001",
  55902=>"110100000",
  55903=>"111110000",
  55904=>"101010000",
  55905=>"010010000",
  55906=>"001100011",
  55907=>"001110010",
  55908=>"110001010",
  55909=>"011110110",
  55910=>"001111111",
  55911=>"001001010",
  55912=>"000000000",
  55913=>"000110111",
  55914=>"101000010",
  55915=>"100010011",
  55916=>"100000011",
  55917=>"100111110",
  55918=>"101010101",
  55919=>"111111001",
  55920=>"001111000",
  55921=>"010100010",
  55922=>"101000110",
  55923=>"000101100",
  55924=>"100100111",
  55925=>"111010110",
  55926=>"101101000",
  55927=>"110111111",
  55928=>"001001100",
  55929=>"101000000",
  55930=>"101010100",
  55931=>"001000010",
  55932=>"110111110",
  55933=>"110000010",
  55934=>"001011001",
  55935=>"000010111",
  55936=>"010000111",
  55937=>"011000011",
  55938=>"011100010",
  55939=>"011100111",
  55940=>"011011000",
  55941=>"111111001",
  55942=>"110111011",
  55943=>"101110110",
  55944=>"111100011",
  55945=>"101110110",
  55946=>"111111011",
  55947=>"001001010",
  55948=>"011110100",
  55949=>"101010100",
  55950=>"000110101",
  55951=>"100100101",
  55952=>"111011111",
  55953=>"001110110",
  55954=>"011100101",
  55955=>"110111010",
  55956=>"010010111",
  55957=>"000110100",
  55958=>"101100111",
  55959=>"011100000",
  55960=>"100011111",
  55961=>"010110000",
  55962=>"101111010",
  55963=>"111001001",
  55964=>"101111011",
  55965=>"100110111",
  55966=>"100001110",
  55967=>"111011011",
  55968=>"100000001",
  55969=>"001101101",
  55970=>"000010010",
  55971=>"010110110",
  55972=>"101101001",
  55973=>"000010111",
  55974=>"101010000",
  55975=>"100000101",
  55976=>"010011001",
  55977=>"111010111",
  55978=>"100100111",
  55979=>"001001000",
  55980=>"100100111",
  55981=>"111101000",
  55982=>"101101001",
  55983=>"110001100",
  55984=>"110011101",
  55985=>"110010000",
  55986=>"110001010",
  55987=>"001101110",
  55988=>"010001011",
  55989=>"011000010",
  55990=>"100000001",
  55991=>"110101000",
  55992=>"011111110",
  55993=>"001000110",
  55994=>"011100001",
  55995=>"100010001",
  55996=>"100001000",
  55997=>"011111000",
  55998=>"110010010",
  55999=>"101101000",
  56000=>"100110001",
  56001=>"010000111",
  56002=>"101000000",
  56003=>"010101110",
  56004=>"100001010",
  56005=>"110010000",
  56006=>"011101111",
  56007=>"000001110",
  56008=>"000010110",
  56009=>"001011101",
  56010=>"000011101",
  56011=>"110011100",
  56012=>"011010011",
  56013=>"010000001",
  56014=>"001101001",
  56015=>"111101100",
  56016=>"010100001",
  56017=>"000010011",
  56018=>"111111111",
  56019=>"001010100",
  56020=>"010111010",
  56021=>"111011010",
  56022=>"001000111",
  56023=>"100001101",
  56024=>"000010100",
  56025=>"111110101",
  56026=>"010111111",
  56027=>"010000000",
  56028=>"101110110",
  56029=>"100001100",
  56030=>"101111011",
  56031=>"000110011",
  56032=>"100000010",
  56033=>"000100000",
  56034=>"001011010",
  56035=>"100101000",
  56036=>"110101111",
  56037=>"000001011",
  56038=>"110001100",
  56039=>"000111011",
  56040=>"100000101",
  56041=>"111101010",
  56042=>"010100100",
  56043=>"100111001",
  56044=>"100111000",
  56045=>"101110001",
  56046=>"000110101",
  56047=>"110110101",
  56048=>"011000000",
  56049=>"100110100",
  56050=>"001100011",
  56051=>"110111011",
  56052=>"111101001",
  56053=>"100001101",
  56054=>"011000010",
  56055=>"111010001",
  56056=>"010101111",
  56057=>"100011011",
  56058=>"111101100",
  56059=>"100110101",
  56060=>"000110101",
  56061=>"100011100",
  56062=>"010001100",
  56063=>"011101110",
  56064=>"010100010",
  56065=>"011011000",
  56066=>"010100010",
  56067=>"000000100",
  56068=>"000001110",
  56069=>"000110110",
  56070=>"010010000",
  56071=>"010101001",
  56072=>"100011100",
  56073=>"000101101",
  56074=>"010000110",
  56075=>"010001110",
  56076=>"101111001",
  56077=>"010101011",
  56078=>"001101000",
  56079=>"000111010",
  56080=>"010010010",
  56081=>"000001001",
  56082=>"110101110",
  56083=>"000100101",
  56084=>"011101000",
  56085=>"001101011",
  56086=>"110011001",
  56087=>"000100000",
  56088=>"011111000",
  56089=>"010101010",
  56090=>"101101010",
  56091=>"101111111",
  56092=>"000000101",
  56093=>"001110010",
  56094=>"111001100",
  56095=>"111011000",
  56096=>"100000000",
  56097=>"001011100",
  56098=>"000010110",
  56099=>"101111100",
  56100=>"100110110",
  56101=>"100101000",
  56102=>"111100110",
  56103=>"010001100",
  56104=>"111010011",
  56105=>"101111110",
  56106=>"101000011",
  56107=>"001001000",
  56108=>"011101101",
  56109=>"000001000",
  56110=>"101000110",
  56111=>"111001000",
  56112=>"011111011",
  56113=>"101110111",
  56114=>"111000110",
  56115=>"110110001",
  56116=>"011101100",
  56117=>"100101000",
  56118=>"001110010",
  56119=>"011111111",
  56120=>"100110011",
  56121=>"011011010",
  56122=>"111100001",
  56123=>"110100100",
  56124=>"111111011",
  56125=>"110010100",
  56126=>"010000010",
  56127=>"001000110",
  56128=>"010110011",
  56129=>"010001010",
  56130=>"000111110",
  56131=>"111111100",
  56132=>"000011010",
  56133=>"000010011",
  56134=>"111111110",
  56135=>"010101000",
  56136=>"010111110",
  56137=>"000011010",
  56138=>"010000110",
  56139=>"100101011",
  56140=>"101011101",
  56141=>"010100010",
  56142=>"011101100",
  56143=>"101111000",
  56144=>"111001101",
  56145=>"101110100",
  56146=>"100000000",
  56147=>"011101011",
  56148=>"011010111",
  56149=>"110010110",
  56150=>"001111001",
  56151=>"101000010",
  56152=>"001010111",
  56153=>"111011001",
  56154=>"110110001",
  56155=>"110010001",
  56156=>"011000011",
  56157=>"110010111",
  56158=>"110010010",
  56159=>"010000100",
  56160=>"010110001",
  56161=>"010001111",
  56162=>"100010000",
  56163=>"000000001",
  56164=>"101111011",
  56165=>"010111101",
  56166=>"001011010",
  56167=>"000010101",
  56168=>"010110001",
  56169=>"000111101",
  56170=>"101101011",
  56171=>"000111011",
  56172=>"010000010",
  56173=>"010110010",
  56174=>"111000000",
  56175=>"001000000",
  56176=>"110110110",
  56177=>"001011001",
  56178=>"011110110",
  56179=>"101010101",
  56180=>"001011100",
  56181=>"001010010",
  56182=>"000100000",
  56183=>"001100010",
  56184=>"101000010",
  56185=>"010100101",
  56186=>"000010001",
  56187=>"011001010",
  56188=>"111101111",
  56189=>"011000000",
  56190=>"100011000",
  56191=>"101111110",
  56192=>"000111111",
  56193=>"100110000",
  56194=>"000001000",
  56195=>"111110010",
  56196=>"101111001",
  56197=>"011010101",
  56198=>"001101101",
  56199=>"100110111",
  56200=>"010100100",
  56201=>"000100110",
  56202=>"000010011",
  56203=>"010101100",
  56204=>"000000101",
  56205=>"000000110",
  56206=>"001111100",
  56207=>"100100011",
  56208=>"100000111",
  56209=>"011100111",
  56210=>"010000000",
  56211=>"110101110",
  56212=>"111101111",
  56213=>"111111111",
  56214=>"011101110",
  56215=>"100101100",
  56216=>"011010111",
  56217=>"010011101",
  56218=>"000101100",
  56219=>"110100101",
  56220=>"101000101",
  56221=>"010000111",
  56222=>"001000101",
  56223=>"001111110",
  56224=>"100110100",
  56225=>"110101001",
  56226=>"101100001",
  56227=>"001000110",
  56228=>"100000100",
  56229=>"111001111",
  56230=>"111110101",
  56231=>"110010000",
  56232=>"111101110",
  56233=>"101101001",
  56234=>"111011110",
  56235=>"100001100",
  56236=>"111001010",
  56237=>"100111111",
  56238=>"000010000",
  56239=>"000001000",
  56240=>"100101000",
  56241=>"111100111",
  56242=>"010100110",
  56243=>"110001001",
  56244=>"101101111",
  56245=>"111000001",
  56246=>"010001101",
  56247=>"010011100",
  56248=>"101010000",
  56249=>"100001001",
  56250=>"100100001",
  56251=>"100100110",
  56252=>"010100100",
  56253=>"101101100",
  56254=>"000100001",
  56255=>"011011101",
  56256=>"010111010",
  56257=>"100001100",
  56258=>"011110000",
  56259=>"011111101",
  56260=>"100101100",
  56261=>"111101111",
  56262=>"111111110",
  56263=>"010001011",
  56264=>"011011110",
  56265=>"100010110",
  56266=>"010001100",
  56267=>"110111000",
  56268=>"010000101",
  56269=>"000000011",
  56270=>"111101100",
  56271=>"111000011",
  56272=>"010011111",
  56273=>"000101100",
  56274=>"011110000",
  56275=>"011011101",
  56276=>"011111101",
  56277=>"000110001",
  56278=>"000001001",
  56279=>"011010110",
  56280=>"100010101",
  56281=>"010111011",
  56282=>"000110110",
  56283=>"011010010",
  56284=>"111101101",
  56285=>"100110000",
  56286=>"001001000",
  56287=>"011001110",
  56288=>"110011010",
  56289=>"110100100",
  56290=>"111011100",
  56291=>"000111111",
  56292=>"000000100",
  56293=>"000110000",
  56294=>"010110111",
  56295=>"101010101",
  56296=>"110101110",
  56297=>"100100000",
  56298=>"011001001",
  56299=>"011111111",
  56300=>"001001110",
  56301=>"000001010",
  56302=>"010101100",
  56303=>"011000000",
  56304=>"010110100",
  56305=>"100001110",
  56306=>"011010010",
  56307=>"000111100",
  56308=>"100101101",
  56309=>"101101001",
  56310=>"111001010",
  56311=>"100011001",
  56312=>"110110010",
  56313=>"010111000",
  56314=>"001000101",
  56315=>"110111100",
  56316=>"001001000",
  56317=>"011110000",
  56318=>"000010000",
  56319=>"110011101",
  56320=>"100010011",
  56321=>"001000001",
  56322=>"001001101",
  56323=>"100111100",
  56324=>"101111011",
  56325=>"010000110",
  56326=>"110011010",
  56327=>"111001110",
  56328=>"000011010",
  56329=>"000111000",
  56330=>"100001100",
  56331=>"101111110",
  56332=>"110011000",
  56333=>"011000111",
  56334=>"110100100",
  56335=>"110100101",
  56336=>"010111100",
  56337=>"000010011",
  56338=>"010101000",
  56339=>"000100001",
  56340=>"110000000",
  56341=>"110111111",
  56342=>"111100001",
  56343=>"001011110",
  56344=>"001100110",
  56345=>"100101110",
  56346=>"110000000",
  56347=>"110110000",
  56348=>"100011011",
  56349=>"000010100",
  56350=>"001000100",
  56351=>"011101110",
  56352=>"000011011",
  56353=>"010111000",
  56354=>"110011111",
  56355=>"010101001",
  56356=>"000110110",
  56357=>"000100101",
  56358=>"111000000",
  56359=>"100111111",
  56360=>"000000100",
  56361=>"111100011",
  56362=>"001111111",
  56363=>"110010001",
  56364=>"101011010",
  56365=>"101011101",
  56366=>"101011111",
  56367=>"111111001",
  56368=>"001011001",
  56369=>"101111000",
  56370=>"010110100",
  56371=>"110111000",
  56372=>"000100000",
  56373=>"111001110",
  56374=>"000001111",
  56375=>"001001001",
  56376=>"111100000",
  56377=>"100111010",
  56378=>"011110011",
  56379=>"001100010",
  56380=>"100000011",
  56381=>"001000010",
  56382=>"001100101",
  56383=>"110011011",
  56384=>"101001011",
  56385=>"111100101",
  56386=>"010001001",
  56387=>"010101110",
  56388=>"100000000",
  56389=>"010010000",
  56390=>"011111011",
  56391=>"101000000",
  56392=>"010110110",
  56393=>"110010100",
  56394=>"111000000",
  56395=>"001011100",
  56396=>"010010111",
  56397=>"010001101",
  56398=>"010110101",
  56399=>"101101011",
  56400=>"011110010",
  56401=>"001010010",
  56402=>"000110101",
  56403=>"100001000",
  56404=>"001110100",
  56405=>"101101000",
  56406=>"101001011",
  56407=>"011001111",
  56408=>"011000001",
  56409=>"001100000",
  56410=>"111010000",
  56411=>"000101100",
  56412=>"011110000",
  56413=>"111101101",
  56414=>"111001000",
  56415=>"111110000",
  56416=>"000111101",
  56417=>"110000000",
  56418=>"111001110",
  56419=>"011001101",
  56420=>"011000000",
  56421=>"111010100",
  56422=>"000000110",
  56423=>"000100011",
  56424=>"101011100",
  56425=>"111101110",
  56426=>"111001000",
  56427=>"110000010",
  56428=>"100100000",
  56429=>"101001100",
  56430=>"100001000",
  56431=>"000111001",
  56432=>"010100110",
  56433=>"110101100",
  56434=>"100100010",
  56435=>"111000011",
  56436=>"100001011",
  56437=>"010001101",
  56438=>"000100010",
  56439=>"100000101",
  56440=>"110100110",
  56441=>"000111001",
  56442=>"010101111",
  56443=>"011001101",
  56444=>"110011110",
  56445=>"011000110",
  56446=>"000111100",
  56447=>"010110011",
  56448=>"101001001",
  56449=>"101100100",
  56450=>"100001000",
  56451=>"011010010",
  56452=>"111110101",
  56453=>"011001010",
  56454=>"001010001",
  56455=>"101111100",
  56456=>"100000000",
  56457=>"111010101",
  56458=>"011000101",
  56459=>"010110000",
  56460=>"100101000",
  56461=>"000001011",
  56462=>"001011011",
  56463=>"010000011",
  56464=>"100010011",
  56465=>"011011011",
  56466=>"011110100",
  56467=>"100000011",
  56468=>"101110011",
  56469=>"011010110",
  56470=>"111000001",
  56471=>"110000011",
  56472=>"100000100",
  56473=>"011111011",
  56474=>"111100100",
  56475=>"010100010",
  56476=>"111101100",
  56477=>"110111111",
  56478=>"111111010",
  56479=>"100111110",
  56480=>"000100110",
  56481=>"111001100",
  56482=>"000111111",
  56483=>"100110111",
  56484=>"000000000",
  56485=>"100000100",
  56486=>"100011001",
  56487=>"100000110",
  56488=>"101011000",
  56489=>"101111011",
  56490=>"000110101",
  56491=>"100010101",
  56492=>"101001110",
  56493=>"000000000",
  56494=>"101011111",
  56495=>"011100000",
  56496=>"000100110",
  56497=>"000011100",
  56498=>"111000011",
  56499=>"000010101",
  56500=>"000000110",
  56501=>"010111110",
  56502=>"001100111",
  56503=>"010101010",
  56504=>"001011000",
  56505=>"111010000",
  56506=>"110000100",
  56507=>"001100111",
  56508=>"101110010",
  56509=>"111101011",
  56510=>"111101111",
  56511=>"001111100",
  56512=>"010000001",
  56513=>"001000111",
  56514=>"010001011",
  56515=>"010001111",
  56516=>"100110000",
  56517=>"111100010",
  56518=>"010110000",
  56519=>"101100110",
  56520=>"010100001",
  56521=>"000100000",
  56522=>"011111111",
  56523=>"000100100",
  56524=>"100010100",
  56525=>"110111000",
  56526=>"101001000",
  56527=>"111011101",
  56528=>"010111101",
  56529=>"111110110",
  56530=>"010101110",
  56531=>"010111001",
  56532=>"100011000",
  56533=>"010101110",
  56534=>"100111101",
  56535=>"111001011",
  56536=>"001011101",
  56537=>"001111110",
  56538=>"110000100",
  56539=>"111111001",
  56540=>"111100011",
  56541=>"111000100",
  56542=>"101011101",
  56543=>"101001111",
  56544=>"101001101",
  56545=>"101110001",
  56546=>"000111111",
  56547=>"001000010",
  56548=>"110011000",
  56549=>"011011010",
  56550=>"100111100",
  56551=>"100010111",
  56552=>"001100000",
  56553=>"011000100",
  56554=>"101101001",
  56555=>"000111101",
  56556=>"000111101",
  56557=>"101010110",
  56558=>"010001101",
  56559=>"110001011",
  56560=>"000100101",
  56561=>"111001001",
  56562=>"001101111",
  56563=>"101110000",
  56564=>"110110011",
  56565=>"000000100",
  56566=>"010010101",
  56567=>"111101010",
  56568=>"110010010",
  56569=>"000110011",
  56570=>"111000000",
  56571=>"100000000",
  56572=>"011100101",
  56573=>"101110000",
  56574=>"101101001",
  56575=>"010110000",
  56576=>"000011100",
  56577=>"001011111",
  56578=>"110111011",
  56579=>"000010111",
  56580=>"111110001",
  56581=>"000000110",
  56582=>"111111100",
  56583=>"001011000",
  56584=>"011100000",
  56585=>"101111101",
  56586=>"011011001",
  56587=>"111011010",
  56588=>"000111010",
  56589=>"111000010",
  56590=>"101010001",
  56591=>"011001111",
  56592=>"000000000",
  56593=>"110100110",
  56594=>"110110010",
  56595=>"000110100",
  56596=>"001110110",
  56597=>"101111000",
  56598=>"010111100",
  56599=>"001011001",
  56600=>"011001001",
  56601=>"110100111",
  56602=>"010101010",
  56603=>"110010111",
  56604=>"001000110",
  56605=>"100100001",
  56606=>"001010011",
  56607=>"011000100",
  56608=>"001001100",
  56609=>"100011011",
  56610=>"100111110",
  56611=>"111010110",
  56612=>"110110010",
  56613=>"100011100",
  56614=>"110101010",
  56615=>"001110011",
  56616=>"110110000",
  56617=>"101010011",
  56618=>"100011111",
  56619=>"110010101",
  56620=>"010100001",
  56621=>"111111111",
  56622=>"010101110",
  56623=>"001100110",
  56624=>"111100111",
  56625=>"101000001",
  56626=>"100101001",
  56627=>"000101010",
  56628=>"111000011",
  56629=>"101000111",
  56630=>"001101111",
  56631=>"101111111",
  56632=>"111111011",
  56633=>"101001000",
  56634=>"111110111",
  56635=>"001011100",
  56636=>"110110011",
  56637=>"011010011",
  56638=>"110000000",
  56639=>"111111100",
  56640=>"011101101",
  56641=>"010100010",
  56642=>"111010101",
  56643=>"000000000",
  56644=>"100110010",
  56645=>"000111010",
  56646=>"010011001",
  56647=>"001001000",
  56648=>"000110000",
  56649=>"111011111",
  56650=>"101010000",
  56651=>"000111110",
  56652=>"111010010",
  56653=>"110001010",
  56654=>"101100011",
  56655=>"111111110",
  56656=>"010001010",
  56657=>"101011110",
  56658=>"011000100",
  56659=>"011110101",
  56660=>"101001000",
  56661=>"010001000",
  56662=>"100010110",
  56663=>"000011101",
  56664=>"110001000",
  56665=>"001000000",
  56666=>"100111010",
  56667=>"110101000",
  56668=>"101011110",
  56669=>"001011110",
  56670=>"001111011",
  56671=>"111110011",
  56672=>"010011101",
  56673=>"100100100",
  56674=>"101000110",
  56675=>"011000000",
  56676=>"101011110",
  56677=>"100010100",
  56678=>"011100000",
  56679=>"100100000",
  56680=>"111011011",
  56681=>"011001000",
  56682=>"010000110",
  56683=>"001001111",
  56684=>"100010000",
  56685=>"011011011",
  56686=>"111010110",
  56687=>"111101010",
  56688=>"110110111",
  56689=>"001010110",
  56690=>"010011011",
  56691=>"110100000",
  56692=>"000000110",
  56693=>"011010100",
  56694=>"111011111",
  56695=>"010000001",
  56696=>"100000111",
  56697=>"011101010",
  56698=>"011110001",
  56699=>"011111010",
  56700=>"011001010",
  56701=>"111100110",
  56702=>"010100001",
  56703=>"101110110",
  56704=>"110110110",
  56705=>"100000000",
  56706=>"000001000",
  56707=>"000111010",
  56708=>"001001000",
  56709=>"010100111",
  56710=>"000110110",
  56711=>"110110101",
  56712=>"000010101",
  56713=>"001110110",
  56714=>"000111011",
  56715=>"100011010",
  56716=>"111110111",
  56717=>"011001001",
  56718=>"100010001",
  56719=>"001011011",
  56720=>"000010010",
  56721=>"001011100",
  56722=>"111011100",
  56723=>"111110001",
  56724=>"000000001",
  56725=>"110101001",
  56726=>"101111010",
  56727=>"100001110",
  56728=>"000011001",
  56729=>"011100000",
  56730=>"111001110",
  56731=>"001110111",
  56732=>"010111111",
  56733=>"101101101",
  56734=>"110101100",
  56735=>"100111111",
  56736=>"101111110",
  56737=>"011101001",
  56738=>"010011100",
  56739=>"111011101",
  56740=>"000110111",
  56741=>"011110001",
  56742=>"110110100",
  56743=>"011001110",
  56744=>"111000110",
  56745=>"110111111",
  56746=>"101111110",
  56747=>"111111111",
  56748=>"000010000",
  56749=>"001010011",
  56750=>"101110101",
  56751=>"010111001",
  56752=>"111101001",
  56753=>"111111111",
  56754=>"000000000",
  56755=>"000100010",
  56756=>"000001110",
  56757=>"110000101",
  56758=>"010101000",
  56759=>"110001011",
  56760=>"111010011",
  56761=>"110100101",
  56762=>"101011001",
  56763=>"001101110",
  56764=>"111101011",
  56765=>"011110000",
  56766=>"110001101",
  56767=>"010111010",
  56768=>"100111101",
  56769=>"001000101",
  56770=>"000110111",
  56771=>"100100100",
  56772=>"011011000",
  56773=>"110011110",
  56774=>"110111101",
  56775=>"011111001",
  56776=>"000001111",
  56777=>"111100111",
  56778=>"001010000",
  56779=>"111100111",
  56780=>"110001000",
  56781=>"111010110",
  56782=>"000110011",
  56783=>"100110010",
  56784=>"010000011",
  56785=>"010100010",
  56786=>"001000000",
  56787=>"111111000",
  56788=>"000010100",
  56789=>"111001001",
  56790=>"010000000",
  56791=>"111101101",
  56792=>"000101000",
  56793=>"111100101",
  56794=>"101000001",
  56795=>"000011001",
  56796=>"000001100",
  56797=>"001100101",
  56798=>"000001010",
  56799=>"001100011",
  56800=>"111010110",
  56801=>"001001100",
  56802=>"111010010",
  56803=>"010101110",
  56804=>"001100001",
  56805=>"000100000",
  56806=>"111000000",
  56807=>"111000011",
  56808=>"010100011",
  56809=>"010000100",
  56810=>"010000010",
  56811=>"000010011",
  56812=>"111010010",
  56813=>"011000000",
  56814=>"001010110",
  56815=>"101001011",
  56816=>"010010100",
  56817=>"011011001",
  56818=>"101010000",
  56819=>"100011011",
  56820=>"110111000",
  56821=>"001000000",
  56822=>"010111111",
  56823=>"100111111",
  56824=>"101000101",
  56825=>"000010011",
  56826=>"000101111",
  56827=>"111100100",
  56828=>"101100010",
  56829=>"111000110",
  56830=>"000000100",
  56831=>"110011101",
  56832=>"110000110",
  56833=>"000011101",
  56834=>"010011110",
  56835=>"111011011",
  56836=>"111011001",
  56837=>"101001000",
  56838=>"000101010",
  56839=>"000101001",
  56840=>"011001110",
  56841=>"001101110",
  56842=>"101000100",
  56843=>"110010011",
  56844=>"010001111",
  56845=>"010110001",
  56846=>"101110000",
  56847=>"100000110",
  56848=>"100010011",
  56849=>"111001001",
  56850=>"101110000",
  56851=>"011000001",
  56852=>"110010001",
  56853=>"000000010",
  56854=>"000010011",
  56855=>"011000010",
  56856=>"100111010",
  56857=>"111011000",
  56858=>"001111011",
  56859=>"110000000",
  56860=>"111011011",
  56861=>"111000011",
  56862=>"010010111",
  56863=>"001001010",
  56864=>"011101111",
  56865=>"010000101",
  56866=>"001001111",
  56867=>"100100001",
  56868=>"100111110",
  56869=>"100100101",
  56870=>"111101110",
  56871=>"011101100",
  56872=>"100101000",
  56873=>"111000110",
  56874=>"111111001",
  56875=>"100011011",
  56876=>"111011101",
  56877=>"100101101",
  56878=>"001000101",
  56879=>"011111110",
  56880=>"010100011",
  56881=>"000111011",
  56882=>"000000001",
  56883=>"101100001",
  56884=>"001000010",
  56885=>"001111011",
  56886=>"011100000",
  56887=>"001010000",
  56888=>"010111010",
  56889=>"110110111",
  56890=>"100010110",
  56891=>"111001110",
  56892=>"011111101",
  56893=>"110000000",
  56894=>"101001111",
  56895=>"000111101",
  56896=>"110001000",
  56897=>"010011110",
  56898=>"001110101",
  56899=>"101110101",
  56900=>"000000111",
  56901=>"111101010",
  56902=>"111010000",
  56903=>"100111000",
  56904=>"000011100",
  56905=>"011101111",
  56906=>"010010100",
  56907=>"000010000",
  56908=>"010000001",
  56909=>"010111100",
  56910=>"010000101",
  56911=>"010001111",
  56912=>"100001001",
  56913=>"000001011",
  56914=>"000010010",
  56915=>"100100110",
  56916=>"100000111",
  56917=>"001001100",
  56918=>"111111100",
  56919=>"001000110",
  56920=>"000011101",
  56921=>"110101010",
  56922=>"110011001",
  56923=>"001101001",
  56924=>"101110100",
  56925=>"110111011",
  56926=>"000100001",
  56927=>"000001101",
  56928=>"010000000",
  56929=>"100000100",
  56930=>"011100011",
  56931=>"011010101",
  56932=>"010000111",
  56933=>"001001001",
  56934=>"111010111",
  56935=>"011111101",
  56936=>"000101100",
  56937=>"101110010",
  56938=>"010111111",
  56939=>"001011010",
  56940=>"110001011",
  56941=>"110100101",
  56942=>"110001101",
  56943=>"110010010",
  56944=>"000100010",
  56945=>"010110011",
  56946=>"111010110",
  56947=>"111010000",
  56948=>"100111111",
  56949=>"111000001",
  56950=>"101111000",
  56951=>"000101110",
  56952=>"100001101",
  56953=>"100110100",
  56954=>"011101111",
  56955=>"111000000",
  56956=>"101100011",
  56957=>"110001110",
  56958=>"100110111",
  56959=>"100010010",
  56960=>"010101010",
  56961=>"001001111",
  56962=>"001101101",
  56963=>"110110001",
  56964=>"110001111",
  56965=>"100101010",
  56966=>"011000101",
  56967=>"101001101",
  56968=>"010010100",
  56969=>"111110011",
  56970=>"010000111",
  56971=>"001111110",
  56972=>"011000010",
  56973=>"110001101",
  56974=>"111111010",
  56975=>"011110000",
  56976=>"100001011",
  56977=>"100101011",
  56978=>"001110101",
  56979=>"111000000",
  56980=>"011010011",
  56981=>"010011100",
  56982=>"100100101",
  56983=>"010010011",
  56984=>"100000100",
  56985=>"000011010",
  56986=>"110010111",
  56987=>"101111001",
  56988=>"110110010",
  56989=>"101011000",
  56990=>"001000110",
  56991=>"100011100",
  56992=>"100100100",
  56993=>"010001000",
  56994=>"000110111",
  56995=>"101000010",
  56996=>"101110111",
  56997=>"111110101",
  56998=>"001110100",
  56999=>"111101100",
  57000=>"000111111",
  57001=>"111111001",
  57002=>"101101001",
  57003=>"111110110",
  57004=>"101100000",
  57005=>"011011101",
  57006=>"110001010",
  57007=>"000001010",
  57008=>"100101100",
  57009=>"011111100",
  57010=>"011010101",
  57011=>"100101010",
  57012=>"011110110",
  57013=>"101100100",
  57014=>"001100010",
  57015=>"100111011",
  57016=>"111011100",
  57017=>"001000110",
  57018=>"110011000",
  57019=>"001101100",
  57020=>"001001000",
  57021=>"000100100",
  57022=>"010010000",
  57023=>"101011110",
  57024=>"001100010",
  57025=>"001111111",
  57026=>"000111100",
  57027=>"000000000",
  57028=>"000101111",
  57029=>"111111111",
  57030=>"001110101",
  57031=>"110011110",
  57032=>"001111111",
  57033=>"010100010",
  57034=>"100001000",
  57035=>"001000011",
  57036=>"100000000",
  57037=>"101110010",
  57038=>"000100110",
  57039=>"100010101",
  57040=>"110101100",
  57041=>"000000101",
  57042=>"010001011",
  57043=>"101110011",
  57044=>"000110100",
  57045=>"110000000",
  57046=>"111111111",
  57047=>"010001010",
  57048=>"100100010",
  57049=>"101111011",
  57050=>"000110011",
  57051=>"010110010",
  57052=>"010011001",
  57053=>"110111011",
  57054=>"111001110",
  57055=>"101001100",
  57056=>"011111101",
  57057=>"000110010",
  57058=>"110011011",
  57059=>"110111011",
  57060=>"001110011",
  57061=>"101101101",
  57062=>"101000000",
  57063=>"000001111",
  57064=>"010100100",
  57065=>"101111100",
  57066=>"110001001",
  57067=>"000100110",
  57068=>"000100000",
  57069=>"000010010",
  57070=>"100100000",
  57071=>"100100001",
  57072=>"001101110",
  57073=>"100000011",
  57074=>"101100111",
  57075=>"001111100",
  57076=>"000100100",
  57077=>"011111111",
  57078=>"101000101",
  57079=>"110011011",
  57080=>"011011011",
  57081=>"000000011",
  57082=>"001100000",
  57083=>"100011101",
  57084=>"110111111",
  57085=>"010001101",
  57086=>"100011010",
  57087=>"000000001",
  57088=>"101100000",
  57089=>"011101001",
  57090=>"110011100",
  57091=>"000100001",
  57092=>"000100001",
  57093=>"011000111",
  57094=>"111110011",
  57095=>"101000101",
  57096=>"010110101",
  57097=>"000110110",
  57098=>"011110100",
  57099=>"111101000",
  57100=>"010100000",
  57101=>"000100001",
  57102=>"011111011",
  57103=>"011001111",
  57104=>"001001100",
  57105=>"110000000",
  57106=>"101111111",
  57107=>"011111000",
  57108=>"000000100",
  57109=>"111000100",
  57110=>"110111001",
  57111=>"010000100",
  57112=>"000101000",
  57113=>"000011010",
  57114=>"011010001",
  57115=>"010101010",
  57116=>"101011011",
  57117=>"010001001",
  57118=>"111111011",
  57119=>"011011111",
  57120=>"000100010",
  57121=>"011111110",
  57122=>"110110001",
  57123=>"011111111",
  57124=>"110011110",
  57125=>"001101101",
  57126=>"111100110",
  57127=>"000000110",
  57128=>"001100100",
  57129=>"111011101",
  57130=>"000100100",
  57131=>"000011110",
  57132=>"000010011",
  57133=>"010100111",
  57134=>"100101111",
  57135=>"010110010",
  57136=>"110011010",
  57137=>"001100010",
  57138=>"011101101",
  57139=>"000000011",
  57140=>"001011011",
  57141=>"111111111",
  57142=>"000110011",
  57143=>"001001010",
  57144=>"111001010",
  57145=>"111110110",
  57146=>"010100101",
  57147=>"001111001",
  57148=>"101011111",
  57149=>"100000100",
  57150=>"110001010",
  57151=>"110100010",
  57152=>"010101100",
  57153=>"001011000",
  57154=>"001001101",
  57155=>"000101101",
  57156=>"111000001",
  57157=>"011010001",
  57158=>"111111100",
  57159=>"110000000",
  57160=>"111110000",
  57161=>"000101111",
  57162=>"101110011",
  57163=>"100101011",
  57164=>"111111011",
  57165=>"000110010",
  57166=>"111000000",
  57167=>"110001001",
  57168=>"110000100",
  57169=>"011000001",
  57170=>"010100011",
  57171=>"000111000",
  57172=>"101101100",
  57173=>"001011000",
  57174=>"110010011",
  57175=>"110111100",
  57176=>"000111111",
  57177=>"000110101",
  57178=>"111101010",
  57179=>"111010111",
  57180=>"010101111",
  57181=>"000000010",
  57182=>"110111111",
  57183=>"111110110",
  57184=>"001101011",
  57185=>"011101100",
  57186=>"101011001",
  57187=>"100101000",
  57188=>"000010111",
  57189=>"110100000",
  57190=>"011101000",
  57191=>"010101100",
  57192=>"101111111",
  57193=>"111101011",
  57194=>"111101011",
  57195=>"101100111",
  57196=>"110000000",
  57197=>"010110111",
  57198=>"010001111",
  57199=>"100110001",
  57200=>"000100001",
  57201=>"100000001",
  57202=>"110111111",
  57203=>"011001000",
  57204=>"100010100",
  57205=>"000010000",
  57206=>"101101000",
  57207=>"100000101",
  57208=>"100110111",
  57209=>"000000010",
  57210=>"111010101",
  57211=>"111100100",
  57212=>"011000000",
  57213=>"101101001",
  57214=>"011000011",
  57215=>"111101101",
  57216=>"101010010",
  57217=>"111000000",
  57218=>"000100110",
  57219=>"011100100",
  57220=>"100001000",
  57221=>"000111011",
  57222=>"111110100",
  57223=>"001111101",
  57224=>"100111101",
  57225=>"111101001",
  57226=>"010010100",
  57227=>"110000110",
  57228=>"010110010",
  57229=>"001101101",
  57230=>"001001100",
  57231=>"111001110",
  57232=>"000110001",
  57233=>"000000110",
  57234=>"111001001",
  57235=>"111100011",
  57236=>"111001101",
  57237=>"100110000",
  57238=>"011011111",
  57239=>"000011110",
  57240=>"011111010",
  57241=>"010111011",
  57242=>"011111001",
  57243=>"010001101",
  57244=>"100111101",
  57245=>"111100110",
  57246=>"100001000",
  57247=>"000011000",
  57248=>"001111001",
  57249=>"101111100",
  57250=>"110101000",
  57251=>"111000101",
  57252=>"110111000",
  57253=>"001011110",
  57254=>"010010110",
  57255=>"010001010",
  57256=>"110001000",
  57257=>"000010111",
  57258=>"011010110",
  57259=>"101001011",
  57260=>"110100100",
  57261=>"111111000",
  57262=>"000011011",
  57263=>"001100110",
  57264=>"001000010",
  57265=>"111001110",
  57266=>"100101000",
  57267=>"001000110",
  57268=>"011011100",
  57269=>"100111001",
  57270=>"100110111",
  57271=>"100010000",
  57272=>"000010110",
  57273=>"011011011",
  57274=>"011000110",
  57275=>"001000101",
  57276=>"001011110",
  57277=>"110000000",
  57278=>"111001111",
  57279=>"110100101",
  57280=>"000000110",
  57281=>"111011001",
  57282=>"101001011",
  57283=>"111111011",
  57284=>"000111010",
  57285=>"101110100",
  57286=>"011010100",
  57287=>"001000000",
  57288=>"101100111",
  57289=>"100111100",
  57290=>"000010010",
  57291=>"000001001",
  57292=>"011010000",
  57293=>"100001000",
  57294=>"111110100",
  57295=>"000001010",
  57296=>"111010110",
  57297=>"101110010",
  57298=>"010101111",
  57299=>"001011110",
  57300=>"010101001",
  57301=>"100010100",
  57302=>"010000100",
  57303=>"000101001",
  57304=>"000111010",
  57305=>"000110111",
  57306=>"110001100",
  57307=>"000010000",
  57308=>"100111001",
  57309=>"010110110",
  57310=>"010011000",
  57311=>"101110111",
  57312=>"111110001",
  57313=>"100100010",
  57314=>"101001110",
  57315=>"101000110",
  57316=>"011101000",
  57317=>"100010110",
  57318=>"010100100",
  57319=>"000001101",
  57320=>"011100111",
  57321=>"001101111",
  57322=>"000010111",
  57323=>"100111000",
  57324=>"100111111",
  57325=>"001100011",
  57326=>"111011001",
  57327=>"011100111",
  57328=>"100101111",
  57329=>"111111010",
  57330=>"100011001",
  57331=>"101101111",
  57332=>"001011100",
  57333=>"010110111",
  57334=>"100110001",
  57335=>"110100111",
  57336=>"000111100",
  57337=>"010000010",
  57338=>"110010100",
  57339=>"001100000",
  57340=>"101001001",
  57341=>"111011010",
  57342=>"100000011",
  57343=>"101111101",
  57344=>"010010011",
  57345=>"111111101",
  57346=>"100010110",
  57347=>"001010101",
  57348=>"000100111",
  57349=>"000010100",
  57350=>"011101111",
  57351=>"111011000",
  57352=>"101000010",
  57353=>"110000010",
  57354=>"010101000",
  57355=>"010001011",
  57356=>"000110100",
  57357=>"001011011",
  57358=>"010101001",
  57359=>"000010010",
  57360=>"110111010",
  57361=>"110110110",
  57362=>"010101001",
  57363=>"010001111",
  57364=>"111111111",
  57365=>"001010110",
  57366=>"111001111",
  57367=>"011001000",
  57368=>"001000111",
  57369=>"001110101",
  57370=>"011110111",
  57371=>"010000001",
  57372=>"000000110",
  57373=>"001111010",
  57374=>"101001100",
  57375=>"111100111",
  57376=>"000001101",
  57377=>"110000000",
  57378=>"111011101",
  57379=>"100011111",
  57380=>"110011010",
  57381=>"110011011",
  57382=>"111110100",
  57383=>"011111011",
  57384=>"100001000",
  57385=>"000100111",
  57386=>"001001010",
  57387=>"110110011",
  57388=>"101111011",
  57389=>"011111111",
  57390=>"011011001",
  57391=>"101011010",
  57392=>"001110101",
  57393=>"101010000",
  57394=>"000101010",
  57395=>"011000000",
  57396=>"101011101",
  57397=>"111110010",
  57398=>"100010101",
  57399=>"001111001",
  57400=>"011000100",
  57401=>"011100111",
  57402=>"101010000",
  57403=>"010101000",
  57404=>"001001111",
  57405=>"111000111",
  57406=>"001001010",
  57407=>"011101110",
  57408=>"001000111",
  57409=>"100111010",
  57410=>"001111000",
  57411=>"001011111",
  57412=>"010110111",
  57413=>"011010001",
  57414=>"010000100",
  57415=>"100000001",
  57416=>"100000001",
  57417=>"010010111",
  57418=>"011101110",
  57419=>"101100011",
  57420=>"001000010",
  57421=>"111000110",
  57422=>"111010001",
  57423=>"000110111",
  57424=>"101111101",
  57425=>"011010010",
  57426=>"111010111",
  57427=>"001111111",
  57428=>"011010100",
  57429=>"111011001",
  57430=>"001001000",
  57431=>"110100000",
  57432=>"000111101",
  57433=>"001001000",
  57434=>"110010000",
  57435=>"001111111",
  57436=>"101111010",
  57437=>"000000010",
  57438=>"001100100",
  57439=>"011001010",
  57440=>"011001000",
  57441=>"110101011",
  57442=>"011111100",
  57443=>"011111111",
  57444=>"010011101",
  57445=>"001101110",
  57446=>"000010000",
  57447=>"011111000",
  57448=>"101000000",
  57449=>"110110001",
  57450=>"100101101",
  57451=>"000110000",
  57452=>"110000011",
  57453=>"100110111",
  57454=>"111011001",
  57455=>"110000110",
  57456=>"110101011",
  57457=>"100011000",
  57458=>"011101100",
  57459=>"011111011",
  57460=>"111001111",
  57461=>"011111111",
  57462=>"001011101",
  57463=>"001000111",
  57464=>"000000001",
  57465=>"100000001",
  57466=>"100101100",
  57467=>"000000010",
  57468=>"011011101",
  57469=>"101100000",
  57470=>"010000001",
  57471=>"011100011",
  57472=>"100100010",
  57473=>"001000110",
  57474=>"011101011",
  57475=>"010000011",
  57476=>"100000010",
  57477=>"011111101",
  57478=>"010010000",
  57479=>"000101010",
  57480=>"110101101",
  57481=>"100001100",
  57482=>"111000000",
  57483=>"000001000",
  57484=>"001111000",
  57485=>"111000111",
  57486=>"100000011",
  57487=>"001001001",
  57488=>"100100001",
  57489=>"101101101",
  57490=>"000110101",
  57491=>"101000110",
  57492=>"000001010",
  57493=>"101000001",
  57494=>"010000110",
  57495=>"110110010",
  57496=>"110101000",
  57497=>"100010111",
  57498=>"000010100",
  57499=>"111010000",
  57500=>"011001011",
  57501=>"111011111",
  57502=>"110100010",
  57503=>"100000111",
  57504=>"101011101",
  57505=>"011100001",
  57506=>"010001100",
  57507=>"001111011",
  57508=>"011100001",
  57509=>"011111100",
  57510=>"111111110",
  57511=>"110010000",
  57512=>"100001110",
  57513=>"111110010",
  57514=>"101011010",
  57515=>"000101011",
  57516=>"111001110",
  57517=>"011111010",
  57518=>"100110011",
  57519=>"110110110",
  57520=>"001101011",
  57521=>"001111001",
  57522=>"010000101",
  57523=>"110001010",
  57524=>"100010001",
  57525=>"100010001",
  57526=>"011011111",
  57527=>"011111101",
  57528=>"111100000",
  57529=>"001110110",
  57530=>"000000101",
  57531=>"111010001",
  57532=>"101000101",
  57533=>"001011010",
  57534=>"111101000",
  57535=>"000100101",
  57536=>"010101110",
  57537=>"001110010",
  57538=>"111111010",
  57539=>"100010010",
  57540=>"101100001",
  57541=>"110010000",
  57542=>"001100001",
  57543=>"010111101",
  57544=>"100111000",
  57545=>"001110000",
  57546=>"001110111",
  57547=>"010010010",
  57548=>"010101010",
  57549=>"101010110",
  57550=>"101111101",
  57551=>"100110001",
  57552=>"011001001",
  57553=>"010011000",
  57554=>"011111100",
  57555=>"011111011",
  57556=>"010001011",
  57557=>"101001101",
  57558=>"100000100",
  57559=>"000010010",
  57560=>"000100101",
  57561=>"101010010",
  57562=>"000001101",
  57563=>"010110001",
  57564=>"110100100",
  57565=>"111111001",
  57566=>"111110101",
  57567=>"110001010",
  57568=>"001000010",
  57569=>"100000001",
  57570=>"101001110",
  57571=>"110101011",
  57572=>"101111001",
  57573=>"000110000",
  57574=>"011101111",
  57575=>"001101111",
  57576=>"001010000",
  57577=>"000101101",
  57578=>"101001101",
  57579=>"111000011",
  57580=>"000110111",
  57581=>"110100000",
  57582=>"001011001",
  57583=>"001100011",
  57584=>"111011000",
  57585=>"011111010",
  57586=>"100101001",
  57587=>"101111000",
  57588=>"100010100",
  57589=>"000010100",
  57590=>"010110101",
  57591=>"010110111",
  57592=>"101001010",
  57593=>"000100100",
  57594=>"100011000",
  57595=>"010100111",
  57596=>"010001101",
  57597=>"110110001",
  57598=>"001100101",
  57599=>"001110111",
  57600=>"001000110",
  57601=>"110010001",
  57602=>"011000110",
  57603=>"011101001",
  57604=>"110101111",
  57605=>"011001101",
  57606=>"000000010",
  57607=>"101011111",
  57608=>"001100000",
  57609=>"101001100",
  57610=>"111000111",
  57611=>"000001101",
  57612=>"011111010",
  57613=>"011011011",
  57614=>"011001000",
  57615=>"101100011",
  57616=>"001100011",
  57617=>"011000100",
  57618=>"101001101",
  57619=>"101111000",
  57620=>"001001011",
  57621=>"001100001",
  57622=>"001000100",
  57623=>"110100001",
  57624=>"011110111",
  57625=>"000111111",
  57626=>"001000111",
  57627=>"001010010",
  57628=>"000010010",
  57629=>"101100110",
  57630=>"001110010",
  57631=>"101001000",
  57632=>"101100111",
  57633=>"000111100",
  57634=>"001000010",
  57635=>"111011101",
  57636=>"010101111",
  57637=>"111010010",
  57638=>"011101000",
  57639=>"001110011",
  57640=>"010011110",
  57641=>"000001000",
  57642=>"001101000",
  57643=>"011111001",
  57644=>"101001010",
  57645=>"000001000",
  57646=>"101000001",
  57647=>"000100100",
  57648=>"000100011",
  57649=>"000000101",
  57650=>"011010010",
  57651=>"100111110",
  57652=>"011010000",
  57653=>"010010011",
  57654=>"000011101",
  57655=>"000000010",
  57656=>"010100000",
  57657=>"010010101",
  57658=>"000000000",
  57659=>"110100110",
  57660=>"001011111",
  57661=>"111001000",
  57662=>"111101000",
  57663=>"000110110",
  57664=>"001000001",
  57665=>"001011010",
  57666=>"000011110",
  57667=>"110100110",
  57668=>"000000011",
  57669=>"110111011",
  57670=>"100100100",
  57671=>"001110110",
  57672=>"010100000",
  57673=>"000010011",
  57674=>"111100101",
  57675=>"010010011",
  57676=>"100111111",
  57677=>"000111110",
  57678=>"000100010",
  57679=>"101010101",
  57680=>"001101000",
  57681=>"000001101",
  57682=>"101111101",
  57683=>"101100000",
  57684=>"011010000",
  57685=>"111001111",
  57686=>"000110111",
  57687=>"101011101",
  57688=>"011100111",
  57689=>"001001001",
  57690=>"111001000",
  57691=>"100000111",
  57692=>"000000001",
  57693=>"011000100",
  57694=>"001111001",
  57695=>"111000011",
  57696=>"100101010",
  57697=>"110101101",
  57698=>"111101101",
  57699=>"000100011",
  57700=>"001000111",
  57701=>"001010100",
  57702=>"001000111",
  57703=>"001100001",
  57704=>"101000100",
  57705=>"001010000",
  57706=>"000000100",
  57707=>"101011010",
  57708=>"011011001",
  57709=>"111111010",
  57710=>"101001010",
  57711=>"010101011",
  57712=>"011100101",
  57713=>"111100001",
  57714=>"010110101",
  57715=>"000010001",
  57716=>"001110110",
  57717=>"101001111",
  57718=>"101000001",
  57719=>"110010010",
  57720=>"110000000",
  57721=>"101011000",
  57722=>"010111001",
  57723=>"111010010",
  57724=>"101101111",
  57725=>"010100101",
  57726=>"100110000",
  57727=>"100111111",
  57728=>"000000101",
  57729=>"100100010",
  57730=>"000111010",
  57731=>"111100111",
  57732=>"011010000",
  57733=>"011111100",
  57734=>"000101110",
  57735=>"000011010",
  57736=>"001001000",
  57737=>"011100110",
  57738=>"101100010",
  57739=>"100010001",
  57740=>"111001101",
  57741=>"110010010",
  57742=>"111011000",
  57743=>"101100101",
  57744=>"000001101",
  57745=>"100001100",
  57746=>"111000100",
  57747=>"011001011",
  57748=>"000001111",
  57749=>"110101000",
  57750=>"000100000",
  57751=>"000000101",
  57752=>"000010010",
  57753=>"011111110",
  57754=>"001100111",
  57755=>"000100000",
  57756=>"011110000",
  57757=>"000100111",
  57758=>"010010010",
  57759=>"000111001",
  57760=>"110100000",
  57761=>"000100001",
  57762=>"111010101",
  57763=>"000010010",
  57764=>"011101000",
  57765=>"011001011",
  57766=>"000000000",
  57767=>"110010100",
  57768=>"111100000",
  57769=>"011111101",
  57770=>"000011110",
  57771=>"010000100",
  57772=>"101000000",
  57773=>"000000100",
  57774=>"110111000",
  57775=>"100100000",
  57776=>"110001111",
  57777=>"010101101",
  57778=>"100001011",
  57779=>"110101010",
  57780=>"111101111",
  57781=>"111110010",
  57782=>"111010000",
  57783=>"011011011",
  57784=>"101100010",
  57785=>"011000010",
  57786=>"000100001",
  57787=>"010011111",
  57788=>"111100101",
  57789=>"011100101",
  57790=>"110000101",
  57791=>"111010011",
  57792=>"100000001",
  57793=>"011000101",
  57794=>"101010001",
  57795=>"101011000",
  57796=>"110101010",
  57797=>"100011100",
  57798=>"101111001",
  57799=>"001000001",
  57800=>"000100001",
  57801=>"000110010",
  57802=>"101000000",
  57803=>"110101110",
  57804=>"110100100",
  57805=>"010110001",
  57806=>"101101000",
  57807=>"111010000",
  57808=>"000110111",
  57809=>"000111110",
  57810=>"111011110",
  57811=>"001110101",
  57812=>"000101111",
  57813=>"000110011",
  57814=>"011110001",
  57815=>"000000001",
  57816=>"001101001",
  57817=>"011010000",
  57818=>"011000001",
  57819=>"010100001",
  57820=>"100011100",
  57821=>"000000100",
  57822=>"101011101",
  57823=>"111110111",
  57824=>"001101100",
  57825=>"101010001",
  57826=>"110100010",
  57827=>"100110001",
  57828=>"000110001",
  57829=>"100001001",
  57830=>"001010000",
  57831=>"010000000",
  57832=>"111101111",
  57833=>"001011110",
  57834=>"011001100",
  57835=>"010011100",
  57836=>"011111000",
  57837=>"100010010",
  57838=>"101010110",
  57839=>"110100110",
  57840=>"110100011",
  57841=>"010111010",
  57842=>"110111111",
  57843=>"101110010",
  57844=>"011001111",
  57845=>"001110000",
  57846=>"000010110",
  57847=>"100110110",
  57848=>"101011110",
  57849=>"101001001",
  57850=>"110001000",
  57851=>"101110101",
  57852=>"011111111",
  57853=>"110011110",
  57854=>"010111110",
  57855=>"100110111",
  57856=>"001011011",
  57857=>"100110001",
  57858=>"111001100",
  57859=>"100110110",
  57860=>"111010111",
  57861=>"111010111",
  57862=>"001100101",
  57863=>"011011000",
  57864=>"010100111",
  57865=>"000101111",
  57866=>"101011001",
  57867=>"111000000",
  57868=>"010111011",
  57869=>"110011001",
  57870=>"000110010",
  57871=>"110001111",
  57872=>"000110001",
  57873=>"111101111",
  57874=>"101001001",
  57875=>"001101011",
  57876=>"000010110",
  57877=>"101000010",
  57878=>"111101101",
  57879=>"101111111",
  57880=>"100101110",
  57881=>"111011111",
  57882=>"101010011",
  57883=>"110001111",
  57884=>"010001011",
  57885=>"110000001",
  57886=>"011100001",
  57887=>"111000111",
  57888=>"000101101",
  57889=>"100111101",
  57890=>"100110100",
  57891=>"001110110",
  57892=>"111110101",
  57893=>"011010000",
  57894=>"010011001",
  57895=>"001100011",
  57896=>"011001100",
  57897=>"000010000",
  57898=>"001110000",
  57899=>"110001001",
  57900=>"101000111",
  57901=>"011110111",
  57902=>"101010000",
  57903=>"000101100",
  57904=>"001100100",
  57905=>"010001001",
  57906=>"011111011",
  57907=>"000000000",
  57908=>"101000000",
  57909=>"011111010",
  57910=>"110111000",
  57911=>"101101011",
  57912=>"101001000",
  57913=>"000101010",
  57914=>"100111010",
  57915=>"111110011",
  57916=>"111001001",
  57917=>"100001001",
  57918=>"000000000",
  57919=>"011001110",
  57920=>"000001101",
  57921=>"101000110",
  57922=>"001010011",
  57923=>"001111001",
  57924=>"000110111",
  57925=>"000011001",
  57926=>"000011101",
  57927=>"010010010",
  57928=>"001000110",
  57929=>"110001100",
  57930=>"001010010",
  57931=>"000110100",
  57932=>"010011010",
  57933=>"010001010",
  57934=>"110010110",
  57935=>"010110111",
  57936=>"100100010",
  57937=>"111111011",
  57938=>"110111111",
  57939=>"100010111",
  57940=>"101011010",
  57941=>"011100110",
  57942=>"100010000",
  57943=>"010110001",
  57944=>"001111001",
  57945=>"101111001",
  57946=>"101011011",
  57947=>"111000001",
  57948=>"110100000",
  57949=>"111011110",
  57950=>"111101110",
  57951=>"110111100",
  57952=>"111111110",
  57953=>"011000011",
  57954=>"000010101",
  57955=>"101111110",
  57956=>"100100111",
  57957=>"000010010",
  57958=>"111000001",
  57959=>"010111011",
  57960=>"001011111",
  57961=>"001100001",
  57962=>"000011010",
  57963=>"110011100",
  57964=>"100101111",
  57965=>"100000110",
  57966=>"001010100",
  57967=>"101010101",
  57968=>"010000000",
  57969=>"101001101",
  57970=>"110101100",
  57971=>"111100010",
  57972=>"111111011",
  57973=>"111010001",
  57974=>"101000111",
  57975=>"110000101",
  57976=>"101110110",
  57977=>"100101001",
  57978=>"110000000",
  57979=>"100100001",
  57980=>"111110011",
  57981=>"111011000",
  57982=>"011011001",
  57983=>"001001011",
  57984=>"010100111",
  57985=>"000010111",
  57986=>"111101110",
  57987=>"100011010",
  57988=>"011010111",
  57989=>"110000000",
  57990=>"011000010",
  57991=>"001111101",
  57992=>"010000011",
  57993=>"010111000",
  57994=>"000010100",
  57995=>"100011110",
  57996=>"111011011",
  57997=>"011000010",
  57998=>"100101000",
  57999=>"110100110",
  58000=>"100110111",
  58001=>"010010010",
  58002=>"011101000",
  58003=>"111101110",
  58004=>"101001110",
  58005=>"101000000",
  58006=>"101100110",
  58007=>"100101110",
  58008=>"100011100",
  58009=>"110000111",
  58010=>"010101101",
  58011=>"111011111",
  58012=>"001000000",
  58013=>"100001011",
  58014=>"010000100",
  58015=>"011100110",
  58016=>"100000001",
  58017=>"001101000",
  58018=>"110100101",
  58019=>"100011101",
  58020=>"010110101",
  58021=>"011001110",
  58022=>"000100110",
  58023=>"001001111",
  58024=>"101010000",
  58025=>"110100010",
  58026=>"000100001",
  58027=>"011100101",
  58028=>"001001000",
  58029=>"001010100",
  58030=>"111010110",
  58031=>"001010010",
  58032=>"100001110",
  58033=>"001110011",
  58034=>"010000001",
  58035=>"001101001",
  58036=>"011000011",
  58037=>"011101011",
  58038=>"111100000",
  58039=>"111010001",
  58040=>"000000101",
  58041=>"000010001",
  58042=>"001011111",
  58043=>"001101011",
  58044=>"011100011",
  58045=>"000101111",
  58046=>"110110010",
  58047=>"011111111",
  58048=>"110101000",
  58049=>"111001101",
  58050=>"010011011",
  58051=>"100101001",
  58052=>"101011000",
  58053=>"011010000",
  58054=>"011100100",
  58055=>"101100100",
  58056=>"101101011",
  58057=>"101111001",
  58058=>"010011100",
  58059=>"011000010",
  58060=>"101010101",
  58061=>"001001100",
  58062=>"000101010",
  58063=>"011101111",
  58064=>"011101001",
  58065=>"001001010",
  58066=>"111111110",
  58067=>"101011000",
  58068=>"111011000",
  58069=>"010000001",
  58070=>"110000111",
  58071=>"010001011",
  58072=>"000110111",
  58073=>"010011011",
  58074=>"000011000",
  58075=>"011110100",
  58076=>"100111111",
  58077=>"000001010",
  58078=>"101100110",
  58079=>"110011001",
  58080=>"010100111",
  58081=>"101001101",
  58082=>"011110110",
  58083=>"011110001",
  58084=>"000011001",
  58085=>"101111010",
  58086=>"111011111",
  58087=>"111110100",
  58088=>"000001011",
  58089=>"101110110",
  58090=>"110000110",
  58091=>"111011001",
  58092=>"101001010",
  58093=>"100101100",
  58094=>"001100000",
  58095=>"111101011",
  58096=>"011101110",
  58097=>"111110001",
  58098=>"111011101",
  58099=>"110011101",
  58100=>"101011111",
  58101=>"100001100",
  58102=>"101111011",
  58103=>"110011110",
  58104=>"100010101",
  58105=>"001001001",
  58106=>"000000001",
  58107=>"101111001",
  58108=>"001100000",
  58109=>"001110010",
  58110=>"010011101",
  58111=>"001010001",
  58112=>"101000100",
  58113=>"010100101",
  58114=>"100101111",
  58115=>"000000101",
  58116=>"100101111",
  58117=>"000000001",
  58118=>"111000000",
  58119=>"110000001",
  58120=>"110101110",
  58121=>"000011111",
  58122=>"101010011",
  58123=>"111011100",
  58124=>"000010000",
  58125=>"110010101",
  58126=>"000000011",
  58127=>"110011010",
  58128=>"110010110",
  58129=>"100011110",
  58130=>"101110001",
  58131=>"100000101",
  58132=>"010001110",
  58133=>"100100100",
  58134=>"000000000",
  58135=>"101000111",
  58136=>"001001101",
  58137=>"011010100",
  58138=>"001101000",
  58139=>"111011011",
  58140=>"011111111",
  58141=>"001000000",
  58142=>"011011010",
  58143=>"110101010",
  58144=>"011001111",
  58145=>"110000111",
  58146=>"010110000",
  58147=>"110001010",
  58148=>"001011001",
  58149=>"010011000",
  58150=>"101001010",
  58151=>"010000100",
  58152=>"110100000",
  58153=>"111010111",
  58154=>"110110110",
  58155=>"011010000",
  58156=>"001011110",
  58157=>"001101101",
  58158=>"100000110",
  58159=>"000110010",
  58160=>"110001011",
  58161=>"101101100",
  58162=>"001000101",
  58163=>"111011000",
  58164=>"111111001",
  58165=>"000100011",
  58166=>"001000100",
  58167=>"011110100",
  58168=>"110010100",
  58169=>"010001011",
  58170=>"110010101",
  58171=>"111000110",
  58172=>"101000111",
  58173=>"111101111",
  58174=>"100010001",
  58175=>"000101011",
  58176=>"111001100",
  58177=>"001000111",
  58178=>"011110000",
  58179=>"111100010",
  58180=>"001010011",
  58181=>"000010101",
  58182=>"111000010",
  58183=>"111101111",
  58184=>"011100011",
  58185=>"100100101",
  58186=>"111011111",
  58187=>"110100001",
  58188=>"100100111",
  58189=>"001011100",
  58190=>"010000100",
  58191=>"010101111",
  58192=>"011101111",
  58193=>"001000100",
  58194=>"000011000",
  58195=>"000101101",
  58196=>"011101110",
  58197=>"010011100",
  58198=>"110110110",
  58199=>"101101001",
  58200=>"010010111",
  58201=>"001111110",
  58202=>"101001010",
  58203=>"110011101",
  58204=>"001011001",
  58205=>"110011111",
  58206=>"101111101",
  58207=>"011000100",
  58208=>"101101100",
  58209=>"101110010",
  58210=>"100011000",
  58211=>"110011101",
  58212=>"100100100",
  58213=>"011000010",
  58214=>"100110011",
  58215=>"101001000",
  58216=>"111110101",
  58217=>"100111111",
  58218=>"111100110",
  58219=>"100001011",
  58220=>"001000110",
  58221=>"110110000",
  58222=>"100101101",
  58223=>"001010110",
  58224=>"010110111",
  58225=>"100011001",
  58226=>"010001111",
  58227=>"100111001",
  58228=>"000110000",
  58229=>"011101001",
  58230=>"111011111",
  58231=>"111010011",
  58232=>"101101101",
  58233=>"001101110",
  58234=>"011001110",
  58235=>"111000010",
  58236=>"010000000",
  58237=>"000101001",
  58238=>"010110001",
  58239=>"001111001",
  58240=>"010110110",
  58241=>"001101010",
  58242=>"000001111",
  58243=>"001011001",
  58244=>"010110010",
  58245=>"101011001",
  58246=>"000010011",
  58247=>"000011001",
  58248=>"111110111",
  58249=>"100001110",
  58250=>"100100010",
  58251=>"100100001",
  58252=>"111011100",
  58253=>"011000100",
  58254=>"000001101",
  58255=>"100110001",
  58256=>"001000011",
  58257=>"110111010",
  58258=>"111111101",
  58259=>"010110101",
  58260=>"000011110",
  58261=>"110001100",
  58262=>"010000100",
  58263=>"010100100",
  58264=>"111101101",
  58265=>"011011100",
  58266=>"000000111",
  58267=>"010100101",
  58268=>"001111101",
  58269=>"111100111",
  58270=>"010001110",
  58271=>"100001000",
  58272=>"000110110",
  58273=>"111011001",
  58274=>"010111101",
  58275=>"011000001",
  58276=>"101100001",
  58277=>"001101010",
  58278=>"100101110",
  58279=>"000011010",
  58280=>"001011010",
  58281=>"011111100",
  58282=>"111110001",
  58283=>"101010010",
  58284=>"101011100",
  58285=>"101101110",
  58286=>"110111110",
  58287=>"110010110",
  58288=>"011100000",
  58289=>"100110011",
  58290=>"101101100",
  58291=>"010110001",
  58292=>"001101100",
  58293=>"001011111",
  58294=>"110100011",
  58295=>"011111100",
  58296=>"000111101",
  58297=>"100110110",
  58298=>"101011100",
  58299=>"010101111",
  58300=>"110001110",
  58301=>"000100001",
  58302=>"010101110",
  58303=>"011000100",
  58304=>"001110110",
  58305=>"001011111",
  58306=>"011000011",
  58307=>"000010001",
  58308=>"000110011",
  58309=>"101111000",
  58310=>"101000011",
  58311=>"000011100",
  58312=>"110100000",
  58313=>"010000111",
  58314=>"001101010",
  58315=>"010110000",
  58316=>"111110101",
  58317=>"011010111",
  58318=>"111100010",
  58319=>"010101000",
  58320=>"101000111",
  58321=>"010011010",
  58322=>"111110111",
  58323=>"010100000",
  58324=>"100001101",
  58325=>"010101011",
  58326=>"100110111",
  58327=>"101100100",
  58328=>"001111001",
  58329=>"000101001",
  58330=>"011111101",
  58331=>"100011110",
  58332=>"010011100",
  58333=>"110110111",
  58334=>"110110101",
  58335=>"101111111",
  58336=>"010001101",
  58337=>"110001000",
  58338=>"101001110",
  58339=>"000011100",
  58340=>"110010111",
  58341=>"001010110",
  58342=>"010101100",
  58343=>"110101000",
  58344=>"101100101",
  58345=>"101010111",
  58346=>"001101010",
  58347=>"101011000",
  58348=>"001001000",
  58349=>"110011011",
  58350=>"111011110",
  58351=>"111001111",
  58352=>"110001010",
  58353=>"000001000",
  58354=>"001001000",
  58355=>"111111111",
  58356=>"001111011",
  58357=>"101000110",
  58358=>"000100011",
  58359=>"000011010",
  58360=>"101001110",
  58361=>"100111101",
  58362=>"101010101",
  58363=>"100111011",
  58364=>"000110100",
  58365=>"101101111",
  58366=>"000011101",
  58367=>"010111010",
  58368=>"100101011",
  58369=>"100001001",
  58370=>"100001001",
  58371=>"110111001",
  58372=>"101100001",
  58373=>"001000010",
  58374=>"110001001",
  58375=>"011010000",
  58376=>"011110111",
  58377=>"101001000",
  58378=>"000011100",
  58379=>"111011110",
  58380=>"100100010",
  58381=>"001110110",
  58382=>"010111000",
  58383=>"110001000",
  58384=>"110110101",
  58385=>"010001000",
  58386=>"100100100",
  58387=>"000100101",
  58388=>"010000101",
  58389=>"110010000",
  58390=>"111000110",
  58391=>"000000101",
  58392=>"010101000",
  58393=>"000100000",
  58394=>"110010101",
  58395=>"110110111",
  58396=>"011100000",
  58397=>"111001001",
  58398=>"011010000",
  58399=>"110000110",
  58400=>"011100100",
  58401=>"101110110",
  58402=>"010100111",
  58403=>"101010111",
  58404=>"010111011",
  58405=>"111011000",
  58406=>"101010111",
  58407=>"000010011",
  58408=>"111101011",
  58409=>"001101000",
  58410=>"100000110",
  58411=>"100100111",
  58412=>"111010000",
  58413=>"001100011",
  58414=>"000100000",
  58415=>"111101000",
  58416=>"001000001",
  58417=>"100110011",
  58418=>"101001111",
  58419=>"101000101",
  58420=>"100010010",
  58421=>"011011111",
  58422=>"011111111",
  58423=>"011001011",
  58424=>"010001010",
  58425=>"000001101",
  58426=>"001001001",
  58427=>"011101100",
  58428=>"111010001",
  58429=>"011001000",
  58430=>"001111111",
  58431=>"011001111",
  58432=>"001111111",
  58433=>"101010101",
  58434=>"110111001",
  58435=>"101100001",
  58436=>"001011011",
  58437=>"010001001",
  58438=>"001001110",
  58439=>"001000110",
  58440=>"111101110",
  58441=>"110000001",
  58442=>"001000101",
  58443=>"011111001",
  58444=>"000001010",
  58445=>"100100001",
  58446=>"101001111",
  58447=>"001101100",
  58448=>"111101001",
  58449=>"000110000",
  58450=>"010101111",
  58451=>"010101010",
  58452=>"100101111",
  58453=>"001101011",
  58454=>"101010111",
  58455=>"101001001",
  58456=>"010110111",
  58457=>"011010111",
  58458=>"100101000",
  58459=>"111110111",
  58460=>"011111010",
  58461=>"001001000",
  58462=>"000111100",
  58463=>"011011110",
  58464=>"010001100",
  58465=>"100111100",
  58466=>"000000000",
  58467=>"001001011",
  58468=>"011000101",
  58469=>"101110100",
  58470=>"101101001",
  58471=>"011110001",
  58472=>"011100111",
  58473=>"011101010",
  58474=>"111011100",
  58475=>"000110100",
  58476=>"100100000",
  58477=>"101000011",
  58478=>"110111011",
  58479=>"010101100",
  58480=>"101001111",
  58481=>"011100001",
  58482=>"010100111",
  58483=>"100000010",
  58484=>"001011110",
  58485=>"110110000",
  58486=>"111001010",
  58487=>"101111110",
  58488=>"001111001",
  58489=>"010101110",
  58490=>"000000001",
  58491=>"101000101",
  58492=>"111110111",
  58493=>"111011000",
  58494=>"101101100",
  58495=>"101010101",
  58496=>"011100000",
  58497=>"010101011",
  58498=>"100000011",
  58499=>"011010001",
  58500=>"101111111",
  58501=>"011101011",
  58502=>"000111110",
  58503=>"101001110",
  58504=>"001100101",
  58505=>"001011000",
  58506=>"010101111",
  58507=>"010110010",
  58508=>"101101000",
  58509=>"011100111",
  58510=>"000111001",
  58511=>"111001100",
  58512=>"000010000",
  58513=>"001011111",
  58514=>"010001110",
  58515=>"011000011",
  58516=>"100101111",
  58517=>"100110111",
  58518=>"000111000",
  58519=>"011011101",
  58520=>"100011000",
  58521=>"111011010",
  58522=>"011100100",
  58523=>"010000110",
  58524=>"111000000",
  58525=>"111101100",
  58526=>"100001100",
  58527=>"000000100",
  58528=>"001010010",
  58529=>"000000010",
  58530=>"011011100",
  58531=>"100001011",
  58532=>"111001010",
  58533=>"001101111",
  58534=>"100000010",
  58535=>"001010101",
  58536=>"010011011",
  58537=>"011010111",
  58538=>"100101111",
  58539=>"100001011",
  58540=>"101101110",
  58541=>"110000111",
  58542=>"100110011",
  58543=>"011001111",
  58544=>"001011000",
  58545=>"100000101",
  58546=>"101110111",
  58547=>"011000100",
  58548=>"110000001",
  58549=>"100011001",
  58550=>"101101001",
  58551=>"100110010",
  58552=>"001101101",
  58553=>"101101101",
  58554=>"011101001",
  58555=>"001111010",
  58556=>"001110010",
  58557=>"111010010",
  58558=>"101111000",
  58559=>"000010100",
  58560=>"111001010",
  58561=>"010010001",
  58562=>"111000000",
  58563=>"001000111",
  58564=>"011100010",
  58565=>"001011000",
  58566=>"111110000",
  58567=>"110100010",
  58568=>"010000000",
  58569=>"011110011",
  58570=>"010100100",
  58571=>"011011000",
  58572=>"000101011",
  58573=>"010101010",
  58574=>"011111111",
  58575=>"001000101",
  58576=>"011011000",
  58577=>"110011101",
  58578=>"100100101",
  58579=>"010010010",
  58580=>"101101101",
  58581=>"111101111",
  58582=>"111011010",
  58583=>"011110010",
  58584=>"111111111",
  58585=>"100111101",
  58586=>"101111010",
  58587=>"101101100",
  58588=>"101001110",
  58589=>"101010101",
  58590=>"011101000",
  58591=>"010011101",
  58592=>"010100000",
  58593=>"000001110",
  58594=>"110110011",
  58595=>"001100011",
  58596=>"111100000",
  58597=>"001001000",
  58598=>"110111111",
  58599=>"110110110",
  58600=>"010111101",
  58601=>"010101110",
  58602=>"001101111",
  58603=>"101011011",
  58604=>"101111101",
  58605=>"111011011",
  58606=>"111001101",
  58607=>"110010000",
  58608=>"000011111",
  58609=>"100010110",
  58610=>"111001110",
  58611=>"001001111",
  58612=>"101011100",
  58613=>"100011000",
  58614=>"000101010",
  58615=>"101101111",
  58616=>"011111011",
  58617=>"101001110",
  58618=>"001001100",
  58619=>"100001101",
  58620=>"110111111",
  58621=>"101101010",
  58622=>"011101111",
  58623=>"101110001",
  58624=>"101100011",
  58625=>"110011110",
  58626=>"000101000",
  58627=>"111110100",
  58628=>"110001000",
  58629=>"011001110",
  58630=>"001010111",
  58631=>"101000000",
  58632=>"111011001",
  58633=>"001111101",
  58634=>"110011110",
  58635=>"101011010",
  58636=>"011010000",
  58637=>"010010110",
  58638=>"110110111",
  58639=>"011101101",
  58640=>"110010001",
  58641=>"111110101",
  58642=>"110100000",
  58643=>"010001000",
  58644=>"011001110",
  58645=>"100100001",
  58646=>"011000000",
  58647=>"001111011",
  58648=>"001100011",
  58649=>"010010110",
  58650=>"111101111",
  58651=>"110000000",
  58652=>"001101101",
  58653=>"111001111",
  58654=>"001110100",
  58655=>"101100010",
  58656=>"010000000",
  58657=>"000001111",
  58658=>"111101001",
  58659=>"101000111",
  58660=>"101111100",
  58661=>"011100001",
  58662=>"111000000",
  58663=>"111011010",
  58664=>"100100101",
  58665=>"010111100",
  58666=>"011111111",
  58667=>"111111111",
  58668=>"100000000",
  58669=>"000101000",
  58670=>"110101100",
  58671=>"101111000",
  58672=>"000000111",
  58673=>"111000000",
  58674=>"111011101",
  58675=>"011010101",
  58676=>"000100011",
  58677=>"000000100",
  58678=>"101011011",
  58679=>"001011111",
  58680=>"011000001",
  58681=>"011001011",
  58682=>"100101110",
  58683=>"001010000",
  58684=>"110011000",
  58685=>"001101010",
  58686=>"000101001",
  58687=>"111001010",
  58688=>"001001010",
  58689=>"000101010",
  58690=>"010100101",
  58691=>"001001001",
  58692=>"101101110",
  58693=>"101001100",
  58694=>"110000001",
  58695=>"100111101",
  58696=>"111101101",
  58697=>"000101100",
  58698=>"001100001",
  58699=>"111110000",
  58700=>"011001011",
  58701=>"011110110",
  58702=>"111111000",
  58703=>"111100111",
  58704=>"010001111",
  58705=>"010101011",
  58706=>"111100001",
  58707=>"101101001",
  58708=>"000101111",
  58709=>"101111001",
  58710=>"010111110",
  58711=>"110100111",
  58712=>"111111011",
  58713=>"110111111",
  58714=>"000010000",
  58715=>"110111000",
  58716=>"000101011",
  58717=>"000011111",
  58718=>"111000010",
  58719=>"100011001",
  58720=>"010001001",
  58721=>"010111001",
  58722=>"100001000",
  58723=>"111101001",
  58724=>"110110101",
  58725=>"011010110",
  58726=>"001101011",
  58727=>"000001000",
  58728=>"101000000",
  58729=>"101111101",
  58730=>"010001001",
  58731=>"110010111",
  58732=>"000010010",
  58733=>"111111001",
  58734=>"100110011",
  58735=>"011110101",
  58736=>"011011000",
  58737=>"000000001",
  58738=>"101110010",
  58739=>"111100110",
  58740=>"111110110",
  58741=>"001001111",
  58742=>"000010100",
  58743=>"000011100",
  58744=>"100000110",
  58745=>"100010110",
  58746=>"111011001",
  58747=>"101100101",
  58748=>"001111101",
  58749=>"001100000",
  58750=>"101111111",
  58751=>"110110110",
  58752=>"100000110",
  58753=>"001011101",
  58754=>"001010000",
  58755=>"011110001",
  58756=>"111001101",
  58757=>"100111000",
  58758=>"101110110",
  58759=>"110111010",
  58760=>"001000101",
  58761=>"100010110",
  58762=>"100001010",
  58763=>"001100111",
  58764=>"100101100",
  58765=>"010010011",
  58766=>"100101111",
  58767=>"011001001",
  58768=>"101011001",
  58769=>"110001100",
  58770=>"111100000",
  58771=>"110010001",
  58772=>"110000111",
  58773=>"001001001",
  58774=>"100111100",
  58775=>"100110101",
  58776=>"010101101",
  58777=>"011000000",
  58778=>"010110000",
  58779=>"001101101",
  58780=>"001111110",
  58781=>"001001100",
  58782=>"011100111",
  58783=>"111100111",
  58784=>"101110101",
  58785=>"000100100",
  58786=>"001011011",
  58787=>"111111111",
  58788=>"111000000",
  58789=>"111111110",
  58790=>"100100110",
  58791=>"011101110",
  58792=>"100101000",
  58793=>"100000000",
  58794=>"100011000",
  58795=>"000000001",
  58796=>"100011000",
  58797=>"001100100",
  58798=>"111010100",
  58799=>"011101011",
  58800=>"001010100",
  58801=>"000100100",
  58802=>"111000111",
  58803=>"001111111",
  58804=>"000111001",
  58805=>"000110000",
  58806=>"100110100",
  58807=>"010001001",
  58808=>"011011011",
  58809=>"101010001",
  58810=>"001011011",
  58811=>"011101001",
  58812=>"000100110",
  58813=>"111110011",
  58814=>"110010010",
  58815=>"110010111",
  58816=>"110001101",
  58817=>"101111111",
  58818=>"011111100",
  58819=>"111010011",
  58820=>"000111101",
  58821=>"110011111",
  58822=>"001010100",
  58823=>"100010011",
  58824=>"111100010",
  58825=>"100001110",
  58826=>"001010110",
  58827=>"111111011",
  58828=>"000000101",
  58829=>"110001100",
  58830=>"111100111",
  58831=>"010111111",
  58832=>"011101001",
  58833=>"111111010",
  58834=>"011110110",
  58835=>"010101111",
  58836=>"100100101",
  58837=>"111110010",
  58838=>"101111101",
  58839=>"001001110",
  58840=>"111110000",
  58841=>"000100110",
  58842=>"011000100",
  58843=>"001110001",
  58844=>"111100110",
  58845=>"100010110",
  58846=>"011100000",
  58847=>"101011001",
  58848=>"001110010",
  58849=>"010011010",
  58850=>"110101001",
  58851=>"101111110",
  58852=>"100001010",
  58853=>"001011101",
  58854=>"101000010",
  58855=>"011011011",
  58856=>"111010111",
  58857=>"100000100",
  58858=>"101100110",
  58859=>"001110100",
  58860=>"101101110",
  58861=>"111100111",
  58862=>"011011011",
  58863=>"001101011",
  58864=>"111101011",
  58865=>"000111001",
  58866=>"100011011",
  58867=>"001011100",
  58868=>"011111010",
  58869=>"000100011",
  58870=>"111001101",
  58871=>"111110111",
  58872=>"101100101",
  58873=>"011001111",
  58874=>"100100000",
  58875=>"001010001",
  58876=>"101110111",
  58877=>"010011100",
  58878=>"110100110",
  58879=>"001111111",
  58880=>"101001010",
  58881=>"011011001",
  58882=>"101100010",
  58883=>"101011100",
  58884=>"110101100",
  58885=>"100001001",
  58886=>"111111010",
  58887=>"111101101",
  58888=>"011000010",
  58889=>"110000001",
  58890=>"101100111",
  58891=>"111101011",
  58892=>"011111110",
  58893=>"001001001",
  58894=>"101001100",
  58895=>"100100001",
  58896=>"000110001",
  58897=>"001010101",
  58898=>"011101011",
  58899=>"000100010",
  58900=>"101110000",
  58901=>"110101100",
  58902=>"100001101",
  58903=>"001111001",
  58904=>"011111111",
  58905=>"000110100",
  58906=>"011001011",
  58907=>"010100101",
  58908=>"011111110",
  58909=>"010000000",
  58910=>"001101011",
  58911=>"010001110",
  58912=>"011000011",
  58913=>"111100011",
  58914=>"001101000",
  58915=>"011111001",
  58916=>"001101011",
  58917=>"101011010",
  58918=>"101000110",
  58919=>"110001010",
  58920=>"111000001",
  58921=>"001001110",
  58922=>"010001010",
  58923=>"110101111",
  58924=>"110101001",
  58925=>"000101110",
  58926=>"101011001",
  58927=>"111111111",
  58928=>"001001000",
  58929=>"001001000",
  58930=>"101100011",
  58931=>"000110111",
  58932=>"101110110",
  58933=>"010010100",
  58934=>"110011100",
  58935=>"011001000",
  58936=>"011011001",
  58937=>"101010001",
  58938=>"100000111",
  58939=>"111011000",
  58940=>"101100110",
  58941=>"111111111",
  58942=>"010001011",
  58943=>"111110100",
  58944=>"001000100",
  58945=>"101011010",
  58946=>"001100100",
  58947=>"100001111",
  58948=>"010001000",
  58949=>"100110011",
  58950=>"101111100",
  58951=>"111000101",
  58952=>"001110110",
  58953=>"011110100",
  58954=>"100110000",
  58955=>"110001011",
  58956=>"111001111",
  58957=>"100101100",
  58958=>"111100000",
  58959=>"001011111",
  58960=>"011111001",
  58961=>"110001001",
  58962=>"100110110",
  58963=>"001101111",
  58964=>"010010000",
  58965=>"000101100",
  58966=>"010001011",
  58967=>"011011010",
  58968=>"101000010",
  58969=>"111101101",
  58970=>"111000101",
  58971=>"010110100",
  58972=>"100000010",
  58973=>"100001100",
  58974=>"000100110",
  58975=>"110001011",
  58976=>"001010110",
  58977=>"111100011",
  58978=>"011000101",
  58979=>"111110001",
  58980=>"100000110",
  58981=>"100011111",
  58982=>"111110000",
  58983=>"000000100",
  58984=>"101011010",
  58985=>"100101000",
  58986=>"001011110",
  58987=>"100001100",
  58988=>"000111000",
  58989=>"000111100",
  58990=>"111100001",
  58991=>"011110001",
  58992=>"100001011",
  58993=>"000000100",
  58994=>"011110100",
  58995=>"110110101",
  58996=>"000101010",
  58997=>"100100100",
  58998=>"100101010",
  58999=>"001100001",
  59000=>"100111110",
  59001=>"000101100",
  59002=>"101000001",
  59003=>"001000111",
  59004=>"111100011",
  59005=>"110111110",
  59006=>"110001110",
  59007=>"000000101",
  59008=>"001000000",
  59009=>"011011000",
  59010=>"001001000",
  59011=>"010000111",
  59012=>"000001011",
  59013=>"101101001",
  59014=>"001001010",
  59015=>"001011110",
  59016=>"011000111",
  59017=>"001111110",
  59018=>"101100010",
  59019=>"001000000",
  59020=>"110011010",
  59021=>"111000000",
  59022=>"000000011",
  59023=>"000011001",
  59024=>"100100111",
  59025=>"000010000",
  59026=>"101101001",
  59027=>"101111011",
  59028=>"000110101",
  59029=>"110100010",
  59030=>"111011111",
  59031=>"001111101",
  59032=>"011111101",
  59033=>"010100011",
  59034=>"100101100",
  59035=>"010100111",
  59036=>"010101001",
  59037=>"110010011",
  59038=>"110000110",
  59039=>"111101110",
  59040=>"001100000",
  59041=>"011110010",
  59042=>"000100010",
  59043=>"000110100",
  59044=>"011010100",
  59045=>"001110011",
  59046=>"001110110",
  59047=>"101000100",
  59048=>"001111010",
  59049=>"101110101",
  59050=>"110100001",
  59051=>"110100000",
  59052=>"100001001",
  59053=>"011110010",
  59054=>"000001101",
  59055=>"010111011",
  59056=>"001101101",
  59057=>"111111110",
  59058=>"010001011",
  59059=>"101001001",
  59060=>"010101011",
  59061=>"011001001",
  59062=>"011101010",
  59063=>"001000001",
  59064=>"101010110",
  59065=>"100001000",
  59066=>"110001101",
  59067=>"111000001",
  59068=>"101111000",
  59069=>"001000000",
  59070=>"001100000",
  59071=>"101010001",
  59072=>"101110000",
  59073=>"111011100",
  59074=>"110001011",
  59075=>"000111111",
  59076=>"001000001",
  59077=>"000100000",
  59078=>"010110000",
  59079=>"100011111",
  59080=>"000100000",
  59081=>"001100011",
  59082=>"100011000",
  59083=>"000100101",
  59084=>"001001011",
  59085=>"111101001",
  59086=>"010010000",
  59087=>"100000010",
  59088=>"101110101",
  59089=>"100100110",
  59090=>"101001110",
  59091=>"010010011",
  59092=>"000100111",
  59093=>"111111101",
  59094=>"011100110",
  59095=>"000110001",
  59096=>"001010011",
  59097=>"001011101",
  59098=>"011100110",
  59099=>"001011111",
  59100=>"011110110",
  59101=>"100101111",
  59102=>"101011110",
  59103=>"010110010",
  59104=>"011000001",
  59105=>"110110011",
  59106=>"101011101",
  59107=>"000000001",
  59108=>"101001110",
  59109=>"000001110",
  59110=>"011100111",
  59111=>"011000010",
  59112=>"101110001",
  59113=>"111110101",
  59114=>"001101100",
  59115=>"110011100",
  59116=>"000111111",
  59117=>"000000100",
  59118=>"100111001",
  59119=>"110010010",
  59120=>"110011000",
  59121=>"110000000",
  59122=>"011100101",
  59123=>"101110101",
  59124=>"110100101",
  59125=>"001100100",
  59126=>"011010101",
  59127=>"001111001",
  59128=>"101000011",
  59129=>"011011110",
  59130=>"010100111",
  59131=>"000010101",
  59132=>"010100001",
  59133=>"101100101",
  59134=>"011001000",
  59135=>"101101111",
  59136=>"101010111",
  59137=>"011111001",
  59138=>"110010001",
  59139=>"100100110",
  59140=>"001100000",
  59141=>"111110100",
  59142=>"010110001",
  59143=>"101000001",
  59144=>"100001101",
  59145=>"011000010",
  59146=>"100010001",
  59147=>"001101101",
  59148=>"101001000",
  59149=>"101100111",
  59150=>"010010111",
  59151=>"101001000",
  59152=>"001011011",
  59153=>"000001001",
  59154=>"110001101",
  59155=>"010011001",
  59156=>"100111000",
  59157=>"101100001",
  59158=>"111110110",
  59159=>"101000111",
  59160=>"001111001",
  59161=>"110000001",
  59162=>"101011111",
  59163=>"111111101",
  59164=>"101101011",
  59165=>"010100111",
  59166=>"101110101",
  59167=>"011010110",
  59168=>"011110111",
  59169=>"011111110",
  59170=>"100100110",
  59171=>"100110000",
  59172=>"110011100",
  59173=>"000100011",
  59174=>"011000101",
  59175=>"010101000",
  59176=>"011011001",
  59177=>"111001011",
  59178=>"001011100",
  59179=>"101101000",
  59180=>"101111010",
  59181=>"101100110",
  59182=>"001001001",
  59183=>"110110100",
  59184=>"000101011",
  59185=>"010110001",
  59186=>"001010011",
  59187=>"101110110",
  59188=>"000101001",
  59189=>"001101111",
  59190=>"110111110",
  59191=>"111111100",
  59192=>"000111110",
  59193=>"101001000",
  59194=>"011100001",
  59195=>"110101101",
  59196=>"110100110",
  59197=>"001101101",
  59198=>"101011111",
  59199=>"001001111",
  59200=>"010110011",
  59201=>"001110001",
  59202=>"111011001",
  59203=>"001111100",
  59204=>"001011000",
  59205=>"010010010",
  59206=>"100001000",
  59207=>"100101000",
  59208=>"011111100",
  59209=>"011001000",
  59210=>"110011001",
  59211=>"100011001",
  59212=>"101101111",
  59213=>"100100110",
  59214=>"111010010",
  59215=>"011100100",
  59216=>"100111110",
  59217=>"110101101",
  59218=>"100010001",
  59219=>"100100100",
  59220=>"111111100",
  59221=>"110010111",
  59222=>"111010101",
  59223=>"110000010",
  59224=>"011000100",
  59225=>"100110011",
  59226=>"010011111",
  59227=>"000100100",
  59228=>"111011001",
  59229=>"100110100",
  59230=>"001011100",
  59231=>"111100110",
  59232=>"001011111",
  59233=>"000100000",
  59234=>"101101000",
  59235=>"111000000",
  59236=>"111111101",
  59237=>"010000100",
  59238=>"101100111",
  59239=>"111000101",
  59240=>"111011010",
  59241=>"110001111",
  59242=>"100001101",
  59243=>"011100110",
  59244=>"001101101",
  59245=>"001000000",
  59246=>"100110110",
  59247=>"000011001",
  59248=>"001010110",
  59249=>"101010011",
  59250=>"000010000",
  59251=>"001110111",
  59252=>"101111111",
  59253=>"110110000",
  59254=>"110010010",
  59255=>"011111110",
  59256=>"001111011",
  59257=>"011000110",
  59258=>"011011110",
  59259=>"010110001",
  59260=>"111111111",
  59261=>"000000001",
  59262=>"100100101",
  59263=>"010110110",
  59264=>"101011111",
  59265=>"110100000",
  59266=>"100101101",
  59267=>"111110110",
  59268=>"101001110",
  59269=>"000001000",
  59270=>"000010000",
  59271=>"000010000",
  59272=>"110011011",
  59273=>"001110111",
  59274=>"110000111",
  59275=>"011011000",
  59276=>"110010010",
  59277=>"001001010",
  59278=>"001001101",
  59279=>"100111111",
  59280=>"001000000",
  59281=>"110100111",
  59282=>"101111100",
  59283=>"010110101",
  59284=>"001010011",
  59285=>"100010100",
  59286=>"001100000",
  59287=>"010010010",
  59288=>"110001000",
  59289=>"111111001",
  59290=>"011100111",
  59291=>"011101110",
  59292=>"111101111",
  59293=>"001001100",
  59294=>"100000111",
  59295=>"011101101",
  59296=>"100011011",
  59297=>"100100010",
  59298=>"011101101",
  59299=>"111001101",
  59300=>"101111100",
  59301=>"100011011",
  59302=>"001000010",
  59303=>"100000111",
  59304=>"011001100",
  59305=>"100001000",
  59306=>"111010010",
  59307=>"110111100",
  59308=>"101000001",
  59309=>"111100111",
  59310=>"100011000",
  59311=>"101000100",
  59312=>"001000101",
  59313=>"000100100",
  59314=>"101001101",
  59315=>"110001110",
  59316=>"111111111",
  59317=>"000000000",
  59318=>"110110010",
  59319=>"011011001",
  59320=>"101110110",
  59321=>"010010111",
  59322=>"101001011",
  59323=>"101111100",
  59324=>"100100011",
  59325=>"101001001",
  59326=>"100011110",
  59327=>"101100000",
  59328=>"000011111",
  59329=>"111111101",
  59330=>"100011111",
  59331=>"111110101",
  59332=>"101111000",
  59333=>"000001000",
  59334=>"010101111",
  59335=>"100100101",
  59336=>"100111111",
  59337=>"101100101",
  59338=>"110111100",
  59339=>"010101010",
  59340=>"110010101",
  59341=>"110110001",
  59342=>"100101110",
  59343=>"001110011",
  59344=>"000101000",
  59345=>"000010110",
  59346=>"010000000",
  59347=>"001000111",
  59348=>"001001101",
  59349=>"000001111",
  59350=>"011011000",
  59351=>"110110111",
  59352=>"101100000",
  59353=>"000111111",
  59354=>"101010011",
  59355=>"011010011",
  59356=>"100100100",
  59357=>"111111010",
  59358=>"111001001",
  59359=>"001011011",
  59360=>"111101110",
  59361=>"010000011",
  59362=>"010111001",
  59363=>"100101000",
  59364=>"101101111",
  59365=>"111101111",
  59366=>"001000110",
  59367=>"101101011",
  59368=>"101001011",
  59369=>"100100010",
  59370=>"100001110",
  59371=>"101101101",
  59372=>"110100110",
  59373=>"000101100",
  59374=>"001010100",
  59375=>"100011101",
  59376=>"110101100",
  59377=>"001001010",
  59378=>"001001110",
  59379=>"100010100",
  59380=>"111101010",
  59381=>"110001111",
  59382=>"110110010",
  59383=>"001110000",
  59384=>"100110100",
  59385=>"100011000",
  59386=>"110010011",
  59387=>"001001001",
  59388=>"101011000",
  59389=>"010111111",
  59390=>"110110011",
  59391=>"011100000",
  59392=>"111010001",
  59393=>"111101101",
  59394=>"100001001",
  59395=>"101111010",
  59396=>"010010101",
  59397=>"001000001",
  59398=>"010010001",
  59399=>"000110110",
  59400=>"111101011",
  59401=>"000000011",
  59402=>"011101011",
  59403=>"110110101",
  59404=>"010011010",
  59405=>"001100000",
  59406=>"010101101",
  59407=>"001110010",
  59408=>"100010100",
  59409=>"011000110",
  59410=>"111010111",
  59411=>"011101110",
  59412=>"001100111",
  59413=>"110001100",
  59414=>"100101000",
  59415=>"000101001",
  59416=>"111000000",
  59417=>"000100101",
  59418=>"111000000",
  59419=>"111110011",
  59420=>"001110111",
  59421=>"001101101",
  59422=>"100011101",
  59423=>"111000010",
  59424=>"000011011",
  59425=>"100100110",
  59426=>"001000000",
  59427=>"001110011",
  59428=>"010011000",
  59429=>"101100111",
  59430=>"111000010",
  59431=>"111101101",
  59432=>"001110111",
  59433=>"000000000",
  59434=>"010000010",
  59435=>"011111111",
  59436=>"101001111",
  59437=>"000110101",
  59438=>"011001110",
  59439=>"011101000",
  59440=>"101100111",
  59441=>"011101111",
  59442=>"011010111",
  59443=>"100110100",
  59444=>"101100000",
  59445=>"011010001",
  59446=>"010110000",
  59447=>"000100010",
  59448=>"111110010",
  59449=>"010010010",
  59450=>"111101010",
  59451=>"100000000",
  59452=>"100011111",
  59453=>"100101011",
  59454=>"001101100",
  59455=>"010111011",
  59456=>"010010000",
  59457=>"110000011",
  59458=>"010011110",
  59459=>"110010011",
  59460=>"100111000",
  59461=>"110101110",
  59462=>"110000001",
  59463=>"000001010",
  59464=>"011011000",
  59465=>"000101111",
  59466=>"110101011",
  59467=>"111001101",
  59468=>"110001001",
  59469=>"000001011",
  59470=>"100010000",
  59471=>"001101111",
  59472=>"100001101",
  59473=>"001011001",
  59474=>"100100101",
  59475=>"000111001",
  59476=>"101100011",
  59477=>"000011110",
  59478=>"111111000",
  59479=>"111000011",
  59480=>"000001011",
  59481=>"110011110",
  59482=>"001110010",
  59483=>"100100101",
  59484=>"010100011",
  59485=>"100011110",
  59486=>"010100101",
  59487=>"010101001",
  59488=>"010111011",
  59489=>"110000111",
  59490=>"011111000",
  59491=>"111110010",
  59492=>"011101011",
  59493=>"100100001",
  59494=>"010111111",
  59495=>"110101110",
  59496=>"000001011",
  59497=>"001111001",
  59498=>"011111101",
  59499=>"101000110",
  59500=>"100011010",
  59501=>"100000011",
  59502=>"010101011",
  59503=>"110100111",
  59504=>"011000011",
  59505=>"111010011",
  59506=>"001110001",
  59507=>"010010110",
  59508=>"110000110",
  59509=>"001100101",
  59510=>"100010101",
  59511=>"101010011",
  59512=>"010000001",
  59513=>"010001111",
  59514=>"101101001",
  59515=>"110101111",
  59516=>"010001000",
  59517=>"111011000",
  59518=>"101110110",
  59519=>"001110111",
  59520=>"001111000",
  59521=>"000101111",
  59522=>"000000111",
  59523=>"111101100",
  59524=>"001011101",
  59525=>"000001010",
  59526=>"001011101",
  59527=>"111100110",
  59528=>"101110110",
  59529=>"100101100",
  59530=>"001011011",
  59531=>"100011101",
  59532=>"000110111",
  59533=>"000110010",
  59534=>"000111111",
  59535=>"011110011",
  59536=>"101000101",
  59537=>"011110011",
  59538=>"101000100",
  59539=>"001110111",
  59540=>"100111100",
  59541=>"110110011",
  59542=>"111011011",
  59543=>"000000000",
  59544=>"011101101",
  59545=>"111000110",
  59546=>"001010010",
  59547=>"000000010",
  59548=>"101100000",
  59549=>"010100000",
  59550=>"000111100",
  59551=>"100010100",
  59552=>"101011101",
  59553=>"110001111",
  59554=>"111011000",
  59555=>"000101011",
  59556=>"100110000",
  59557=>"011111111",
  59558=>"011111001",
  59559=>"000000010",
  59560=>"100100010",
  59561=>"001111110",
  59562=>"010001101",
  59563=>"011001100",
  59564=>"110100100",
  59565=>"111110101",
  59566=>"000001111",
  59567=>"101100010",
  59568=>"010100000",
  59569=>"100010011",
  59570=>"110111001",
  59571=>"101010001",
  59572=>"111011111",
  59573=>"010110010",
  59574=>"101010000",
  59575=>"111101010",
  59576=>"010111000",
  59577=>"010100110",
  59578=>"101010100",
  59579=>"111110110",
  59580=>"011110011",
  59581=>"111111001",
  59582=>"011101100",
  59583=>"110111011",
  59584=>"110110101",
  59585=>"111001110",
  59586=>"000111111",
  59587=>"111011001",
  59588=>"001111111",
  59589=>"111100001",
  59590=>"010100111",
  59591=>"011110111",
  59592=>"010000000",
  59593=>"100000001",
  59594=>"010001011",
  59595=>"000110010",
  59596=>"000101011",
  59597=>"100111111",
  59598=>"111010111",
  59599=>"000101000",
  59600=>"110110011",
  59601=>"011100101",
  59602=>"110000001",
  59603=>"100000001",
  59604=>"101000100",
  59605=>"011100011",
  59606=>"010011110",
  59607=>"000101110",
  59608=>"010010001",
  59609=>"010100000",
  59610=>"101000001",
  59611=>"010010100",
  59612=>"111110000",
  59613=>"000111111",
  59614=>"101001101",
  59615=>"010011111",
  59616=>"000011111",
  59617=>"000010000",
  59618=>"101101101",
  59619=>"100000001",
  59620=>"000111001",
  59621=>"001001010",
  59622=>"110011011",
  59623=>"100111011",
  59624=>"110011001",
  59625=>"100111000",
  59626=>"101100011",
  59627=>"101010101",
  59628=>"101010010",
  59629=>"100101111",
  59630=>"011111001",
  59631=>"011011011",
  59632=>"001011000",
  59633=>"001011001",
  59634=>"011101100",
  59635=>"001010001",
  59636=>"111001100",
  59637=>"111110001",
  59638=>"111100101",
  59639=>"101111000",
  59640=>"011000111",
  59641=>"010111010",
  59642=>"001000001",
  59643=>"100101010",
  59644=>"101111100",
  59645=>"110000111",
  59646=>"011111101",
  59647=>"000100001",
  59648=>"110110110",
  59649=>"101010000",
  59650=>"110110001",
  59651=>"101101001",
  59652=>"010101100",
  59653=>"010010010",
  59654=>"111011101",
  59655=>"100011000",
  59656=>"011000000",
  59657=>"100110011",
  59658=>"010001011",
  59659=>"110000110",
  59660=>"010110111",
  59661=>"111101001",
  59662=>"001100101",
  59663=>"101101100",
  59664=>"111111011",
  59665=>"111101011",
  59666=>"100000011",
  59667=>"111011101",
  59668=>"111000100",
  59669=>"100101001",
  59670=>"011000000",
  59671=>"110101000",
  59672=>"101000001",
  59673=>"001000111",
  59674=>"010011000",
  59675=>"110101001",
  59676=>"111011000",
  59677=>"110001100",
  59678=>"111110010",
  59679=>"101010000",
  59680=>"101110000",
  59681=>"111011000",
  59682=>"001011001",
  59683=>"011111011",
  59684=>"111011111",
  59685=>"111100111",
  59686=>"110111011",
  59687=>"010100111",
  59688=>"101111110",
  59689=>"101101100",
  59690=>"110010011",
  59691=>"000000000",
  59692=>"010011111",
  59693=>"111111010",
  59694=>"110000111",
  59695=>"011111100",
  59696=>"011101101",
  59697=>"001111101",
  59698=>"011100110",
  59699=>"000110011",
  59700=>"101010110",
  59701=>"000010111",
  59702=>"011110101",
  59703=>"001010001",
  59704=>"000110001",
  59705=>"111000111",
  59706=>"100000000",
  59707=>"011000111",
  59708=>"101101001",
  59709=>"111100100",
  59710=>"000110010",
  59711=>"001001000",
  59712=>"011011100",
  59713=>"110000111",
  59714=>"111100100",
  59715=>"010010111",
  59716=>"011011011",
  59717=>"100100001",
  59718=>"000110100",
  59719=>"110001010",
  59720=>"000101110",
  59721=>"000100001",
  59722=>"111101010",
  59723=>"100011101",
  59724=>"010010111",
  59725=>"000011111",
  59726=>"110011001",
  59727=>"010011000",
  59728=>"110101101",
  59729=>"110110011",
  59730=>"001010000",
  59731=>"011111001",
  59732=>"110001101",
  59733=>"010010010",
  59734=>"001101000",
  59735=>"011100010",
  59736=>"100010111",
  59737=>"011001000",
  59738=>"110010101",
  59739=>"110000110",
  59740=>"011010111",
  59741=>"111111010",
  59742=>"111011110",
  59743=>"111000001",
  59744=>"101110110",
  59745=>"000110110",
  59746=>"000000010",
  59747=>"011111101",
  59748=>"110110010",
  59749=>"001101010",
  59750=>"000100010",
  59751=>"110011001",
  59752=>"101110111",
  59753=>"110110011",
  59754=>"001011110",
  59755=>"010001000",
  59756=>"011101101",
  59757=>"110110000",
  59758=>"101111000",
  59759=>"100000001",
  59760=>"110010000",
  59761=>"111101000",
  59762=>"000100001",
  59763=>"111101100",
  59764=>"010100000",
  59765=>"000001111",
  59766=>"100101010",
  59767=>"110000110",
  59768=>"101100000",
  59769=>"100101011",
  59770=>"010011011",
  59771=>"101110111",
  59772=>"100001011",
  59773=>"010010111",
  59774=>"111110110",
  59775=>"101110110",
  59776=>"010110110",
  59777=>"110100000",
  59778=>"111111101",
  59779=>"010000111",
  59780=>"110110101",
  59781=>"001011010",
  59782=>"010110000",
  59783=>"010011100",
  59784=>"000100110",
  59785=>"010101111",
  59786=>"011101101",
  59787=>"010000110",
  59788=>"111101011",
  59789=>"011111000",
  59790=>"111111111",
  59791=>"111100101",
  59792=>"100101111",
  59793=>"001101000",
  59794=>"000111010",
  59795=>"110010010",
  59796=>"100011000",
  59797=>"110100010",
  59798=>"100000001",
  59799=>"000011010",
  59800=>"101000100",
  59801=>"000011111",
  59802=>"010011110",
  59803=>"000010001",
  59804=>"100101011",
  59805=>"100100101",
  59806=>"101101110",
  59807=>"110100100",
  59808=>"001001101",
  59809=>"010000001",
  59810=>"011110101",
  59811=>"011100001",
  59812=>"111100001",
  59813=>"001001100",
  59814=>"001000010",
  59815=>"111011111",
  59816=>"011000001",
  59817=>"000100010",
  59818=>"110001011",
  59819=>"100010000",
  59820=>"000010000",
  59821=>"000100100",
  59822=>"110000010",
  59823=>"000001010",
  59824=>"100110110",
  59825=>"011101100",
  59826=>"010010111",
  59827=>"000100110",
  59828=>"110011010",
  59829=>"101110101",
  59830=>"011101011",
  59831=>"000100110",
  59832=>"111110010",
  59833=>"110110100",
  59834=>"000111111",
  59835=>"110100101",
  59836=>"011000001",
  59837=>"011110011",
  59838=>"111100001",
  59839=>"100111110",
  59840=>"101010110",
  59841=>"001000111",
  59842=>"000110111",
  59843=>"110001100",
  59844=>"010000010",
  59845=>"000000000",
  59846=>"101011010",
  59847=>"000001010",
  59848=>"110100011",
  59849=>"001111110",
  59850=>"000011000",
  59851=>"110010111",
  59852=>"100111110",
  59853=>"000111001",
  59854=>"011111111",
  59855=>"010111011",
  59856=>"100001100",
  59857=>"111010001",
  59858=>"010111111",
  59859=>"010000001",
  59860=>"110011111",
  59861=>"010111101",
  59862=>"000001100",
  59863=>"111010011",
  59864=>"110110111",
  59865=>"100010101",
  59866=>"001101010",
  59867=>"010000001",
  59868=>"101011001",
  59869=>"111000011",
  59870=>"110000111",
  59871=>"100110000",
  59872=>"000001001",
  59873=>"001100000",
  59874=>"110000000",
  59875=>"100101010",
  59876=>"011001101",
  59877=>"110110111",
  59878=>"001100100",
  59879=>"101001100",
  59880=>"001000011",
  59881=>"111110100",
  59882=>"100001101",
  59883=>"110001101",
  59884=>"111110111",
  59885=>"111000000",
  59886=>"000100000",
  59887=>"110000001",
  59888=>"101100101",
  59889=>"111110010",
  59890=>"101100011",
  59891=>"011011001",
  59892=>"010100100",
  59893=>"000010111",
  59894=>"000000111",
  59895=>"010100010",
  59896=>"010011111",
  59897=>"100011110",
  59898=>"101000101",
  59899=>"011111100",
  59900=>"111100011",
  59901=>"100100111",
  59902=>"010110100",
  59903=>"000100111",
  59904=>"010101100",
  59905=>"000000000",
  59906=>"110001111",
  59907=>"110000001",
  59908=>"101101010",
  59909=>"010111100",
  59910=>"010001010",
  59911=>"100110001",
  59912=>"010001000",
  59913=>"100010001",
  59914=>"010001000",
  59915=>"111010010",
  59916=>"000011010",
  59917=>"111010001",
  59918=>"101001110",
  59919=>"011100111",
  59920=>"011100000",
  59921=>"101000001",
  59922=>"111100110",
  59923=>"111101001",
  59924=>"010101011",
  59925=>"111000001",
  59926=>"000100100",
  59927=>"010111000",
  59928=>"101101010",
  59929=>"111000111",
  59930=>"101110011",
  59931=>"000010101",
  59932=>"010100010",
  59933=>"010111111",
  59934=>"100110110",
  59935=>"011101011",
  59936=>"001010000",
  59937=>"011010100",
  59938=>"000111000",
  59939=>"100111100",
  59940=>"111111100",
  59941=>"101100101",
  59942=>"110001000",
  59943=>"110011000",
  59944=>"011111100",
  59945=>"111001110",
  59946=>"001111001",
  59947=>"111011010",
  59948=>"101010101",
  59949=>"000000100",
  59950=>"101110100",
  59951=>"001000011",
  59952=>"100111111",
  59953=>"011001101",
  59954=>"010001011",
  59955=>"011001111",
  59956=>"011100100",
  59957=>"101100111",
  59958=>"010000011",
  59959=>"100110111",
  59960=>"000100111",
  59961=>"000110100",
  59962=>"110010101",
  59963=>"010100000",
  59964=>"111110000",
  59965=>"001100101",
  59966=>"000101100",
  59967=>"000101111",
  59968=>"100000000",
  59969=>"011001010",
  59970=>"010011000",
  59971=>"011011000",
  59972=>"101010111",
  59973=>"111010100",
  59974=>"011101001",
  59975=>"111100101",
  59976=>"011011111",
  59977=>"101110011",
  59978=>"101000010",
  59979=>"010010010",
  59980=>"101000001",
  59981=>"100100111",
  59982=>"111000001",
  59983=>"100101010",
  59984=>"110101000",
  59985=>"011011110",
  59986=>"000010111",
  59987=>"010111100",
  59988=>"100111100",
  59989=>"110111010",
  59990=>"000100010",
  59991=>"010011001",
  59992=>"111111001",
  59993=>"111110110",
  59994=>"011001100",
  59995=>"010100110",
  59996=>"000111100",
  59997=>"100000010",
  59998=>"101110010",
  59999=>"100101010",
  60000=>"110010111",
  60001=>"110011000",
  60002=>"011110010",
  60003=>"111000010",
  60004=>"101000111",
  60005=>"011001000",
  60006=>"000101100",
  60007=>"111000101",
  60008=>"011100110",
  60009=>"001110110",
  60010=>"000110111",
  60011=>"111011001",
  60012=>"111001101",
  60013=>"100011100",
  60014=>"111101111",
  60015=>"001001010",
  60016=>"000100001",
  60017=>"000011010",
  60018=>"000111101",
  60019=>"000111101",
  60020=>"000010000",
  60021=>"010110000",
  60022=>"010001111",
  60023=>"011100010",
  60024=>"001110110",
  60025=>"001011100",
  60026=>"100010111",
  60027=>"010001011",
  60028=>"001101111",
  60029=>"111000001",
  60030=>"100101001",
  60031=>"111101000",
  60032=>"000111011",
  60033=>"000110010",
  60034=>"110011001",
  60035=>"111011001",
  60036=>"000111011",
  60037=>"000100111",
  60038=>"010110111",
  60039=>"000000101",
  60040=>"100000001",
  60041=>"011010011",
  60042=>"111001000",
  60043=>"000011010",
  60044=>"000101001",
  60045=>"001010111",
  60046=>"111101011",
  60047=>"011011111",
  60048=>"011000101",
  60049=>"001111010",
  60050=>"000001100",
  60051=>"011001101",
  60052=>"001101111",
  60053=>"000011011",
  60054=>"101011111",
  60055=>"001111110",
  60056=>"100101011",
  60057=>"101000101",
  60058=>"101110101",
  60059=>"101111011",
  60060=>"110001111",
  60061=>"000000111",
  60062=>"000010000",
  60063=>"101100101",
  60064=>"000000000",
  60065=>"001010011",
  60066=>"110110011",
  60067=>"000010011",
  60068=>"000111100",
  60069=>"101111100",
  60070=>"000111100",
  60071=>"000001010",
  60072=>"010010001",
  60073=>"100001001",
  60074=>"001000010",
  60075=>"000001110",
  60076=>"011011011",
  60077=>"100100001",
  60078=>"110101110",
  60079=>"001111110",
  60080=>"011111100",
  60081=>"011111001",
  60082=>"001011110",
  60083=>"111110011",
  60084=>"011000110",
  60085=>"101101011",
  60086=>"100000000",
  60087=>"111001001",
  60088=>"001111000",
  60089=>"001000000",
  60090=>"111111100",
  60091=>"001011101",
  60092=>"111011110",
  60093=>"001011000",
  60094=>"010001100",
  60095=>"010110010",
  60096=>"010010000",
  60097=>"110100100",
  60098=>"001001100",
  60099=>"110000011",
  60100=>"110100010",
  60101=>"011111000",
  60102=>"010010110",
  60103=>"100110000",
  60104=>"000001001",
  60105=>"011011101",
  60106=>"000111110",
  60107=>"101011101",
  60108=>"011010000",
  60109=>"100000110",
  60110=>"011111000",
  60111=>"011101110",
  60112=>"001111001",
  60113=>"111001101",
  60114=>"001111110",
  60115=>"001111011",
  60116=>"111101110",
  60117=>"101011101",
  60118=>"010110100",
  60119=>"111000001",
  60120=>"010110010",
  60121=>"111100110",
  60122=>"000110000",
  60123=>"011101000",
  60124=>"011110000",
  60125=>"000011101",
  60126=>"101011111",
  60127=>"010100101",
  60128=>"000100111",
  60129=>"000001100",
  60130=>"111100001",
  60131=>"011100000",
  60132=>"000011011",
  60133=>"110001011",
  60134=>"010000010",
  60135=>"001101100",
  60136=>"011000001",
  60137=>"111000110",
  60138=>"010110001",
  60139=>"001010011",
  60140=>"010001000",
  60141=>"111101110",
  60142=>"001100101",
  60143=>"111101101",
  60144=>"111101101",
  60145=>"000101111",
  60146=>"100100100",
  60147=>"111001101",
  60148=>"101001101",
  60149=>"001110011",
  60150=>"111101000",
  60151=>"000011011",
  60152=>"011011101",
  60153=>"111010100",
  60154=>"010101011",
  60155=>"100000001",
  60156=>"000011101",
  60157=>"100010101",
  60158=>"011001011",
  60159=>"110100100",
  60160=>"010010010",
  60161=>"101110011",
  60162=>"101101101",
  60163=>"100101111",
  60164=>"110011000",
  60165=>"100101001",
  60166=>"110110111",
  60167=>"111010101",
  60168=>"001110001",
  60169=>"001001010",
  60170=>"110101011",
  60171=>"001011110",
  60172=>"111000100",
  60173=>"000101011",
  60174=>"110101000",
  60175=>"101001011",
  60176=>"001010011",
  60177=>"011011011",
  60178=>"010000010",
  60179=>"111111101",
  60180=>"011101001",
  60181=>"010110011",
  60182=>"010011000",
  60183=>"001000100",
  60184=>"011010001",
  60185=>"001101000",
  60186=>"110010110",
  60187=>"010100101",
  60188=>"110111111",
  60189=>"010110110",
  60190=>"111001101",
  60191=>"010111001",
  60192=>"101111000",
  60193=>"001001001",
  60194=>"101101100",
  60195=>"001001110",
  60196=>"000011001",
  60197=>"101000000",
  60198=>"001000010",
  60199=>"100001110",
  60200=>"110111000",
  60201=>"111011010",
  60202=>"011101011",
  60203=>"100100011",
  60204=>"010011011",
  60205=>"000001000",
  60206=>"101111010",
  60207=>"001000010",
  60208=>"110100110",
  60209=>"101011111",
  60210=>"111101100",
  60211=>"001000101",
  60212=>"101111011",
  60213=>"010000100",
  60214=>"101101110",
  60215=>"000010000",
  60216=>"010101010",
  60217=>"001101000",
  60218=>"011101001",
  60219=>"110111110",
  60220=>"111010010",
  60221=>"110000110",
  60222=>"010100101",
  60223=>"100110000",
  60224=>"000100100",
  60225=>"110000111",
  60226=>"110010000",
  60227=>"010000100",
  60228=>"100000000",
  60229=>"110110101",
  60230=>"011000001",
  60231=>"111101011",
  60232=>"110110011",
  60233=>"000000011",
  60234=>"101010011",
  60235=>"000010001",
  60236=>"110011110",
  60237=>"101111001",
  60238=>"010011000",
  60239=>"001000101",
  60240=>"111101001",
  60241=>"010001100",
  60242=>"011110010",
  60243=>"010000110",
  60244=>"111100111",
  60245=>"001011100",
  60246=>"010110000",
  60247=>"000111011",
  60248=>"000111110",
  60249=>"110111000",
  60250=>"011101111",
  60251=>"110110111",
  60252=>"000011111",
  60253=>"000101101",
  60254=>"011111101",
  60255=>"010000101",
  60256=>"111001110",
  60257=>"000010111",
  60258=>"011111000",
  60259=>"010010100",
  60260=>"100111110",
  60261=>"110001001",
  60262=>"001010110",
  60263=>"111001011",
  60264=>"001110100",
  60265=>"111011001",
  60266=>"110111010",
  60267=>"001000110",
  60268=>"001100000",
  60269=>"010001101",
  60270=>"110100111",
  60271=>"000000110",
  60272=>"101011010",
  60273=>"001100001",
  60274=>"111011001",
  60275=>"111010011",
  60276=>"101110100",
  60277=>"111100000",
  60278=>"000000000",
  60279=>"000010011",
  60280=>"000101001",
  60281=>"000011101",
  60282=>"010000011",
  60283=>"000001101",
  60284=>"011001011",
  60285=>"011011011",
  60286=>"101001010",
  60287=>"101100110",
  60288=>"110001100",
  60289=>"000000001",
  60290=>"100101110",
  60291=>"101011001",
  60292=>"100111001",
  60293=>"101000011",
  60294=>"100000100",
  60295=>"100010111",
  60296=>"001100110",
  60297=>"010110010",
  60298=>"011000001",
  60299=>"111011010",
  60300=>"110001001",
  60301=>"111100010",
  60302=>"010011001",
  60303=>"011001111",
  60304=>"111001111",
  60305=>"001010001",
  60306=>"001011110",
  60307=>"001010011",
  60308=>"011110011",
  60309=>"111100101",
  60310=>"000011001",
  60311=>"111110111",
  60312=>"111011001",
  60313=>"011100111",
  60314=>"111011100",
  60315=>"110100011",
  60316=>"110110010",
  60317=>"001111111",
  60318=>"010011100",
  60319=>"001000110",
  60320=>"011000001",
  60321=>"011000010",
  60322=>"100011110",
  60323=>"001011101",
  60324=>"101111000",
  60325=>"111100000",
  60326=>"010110010",
  60327=>"011010001",
  60328=>"111010100",
  60329=>"000010000",
  60330=>"110110111",
  60331=>"110010001",
  60332=>"111000100",
  60333=>"000001101",
  60334=>"111111111",
  60335=>"100010010",
  60336=>"111100000",
  60337=>"101111000",
  60338=>"100010100",
  60339=>"000000010",
  60340=>"011011111",
  60341=>"011001111",
  60342=>"001000111",
  60343=>"100111011",
  60344=>"011101111",
  60345=>"000000111",
  60346=>"001110011",
  60347=>"101100100",
  60348=>"110000000",
  60349=>"101100100",
  60350=>"000001110",
  60351=>"010001000",
  60352=>"000011010",
  60353=>"000000000",
  60354=>"100111011",
  60355=>"000011101",
  60356=>"100011001",
  60357=>"100100101",
  60358=>"100001100",
  60359=>"111111010",
  60360=>"111011011",
  60361=>"100000111",
  60362=>"000110001",
  60363=>"011000010",
  60364=>"101100101",
  60365=>"000110000",
  60366=>"011011000",
  60367=>"010110101",
  60368=>"011100111",
  60369=>"000100000",
  60370=>"001010011",
  60371=>"101001000",
  60372=>"010000011",
  60373=>"110111101",
  60374=>"111101110",
  60375=>"000110010",
  60376=>"101001111",
  60377=>"001011111",
  60378=>"101101000",
  60379=>"000111100",
  60380=>"111110000",
  60381=>"100111110",
  60382=>"011101010",
  60383=>"011010000",
  60384=>"100100100",
  60385=>"001101001",
  60386=>"110010111",
  60387=>"101100000",
  60388=>"001101000",
  60389=>"111101000",
  60390=>"000110111",
  60391=>"011001110",
  60392=>"001100010",
  60393=>"001101101",
  60394=>"100010010",
  60395=>"111000010",
  60396=>"100110100",
  60397=>"111101010",
  60398=>"010011010",
  60399=>"000110111",
  60400=>"110011000",
  60401=>"101001110",
  60402=>"110111100",
  60403=>"001110001",
  60404=>"101101110",
  60405=>"011100110",
  60406=>"110110110",
  60407=>"111101000",
  60408=>"001111000",
  60409=>"011011110",
  60410=>"100111000",
  60411=>"011100011",
  60412=>"110001110",
  60413=>"111010010",
  60414=>"011101111",
  60415=>"010010011",
  60416=>"111000010",
  60417=>"011001111",
  60418=>"010001110",
  60419=>"010110000",
  60420=>"110111101",
  60421=>"001110011",
  60422=>"100101100",
  60423=>"111001111",
  60424=>"101010101",
  60425=>"011101000",
  60426=>"101100111",
  60427=>"100101110",
  60428=>"111111010",
  60429=>"010010000",
  60430=>"101111010",
  60431=>"100000110",
  60432=>"000001100",
  60433=>"100100010",
  60434=>"000010000",
  60435=>"001101110",
  60436=>"100001101",
  60437=>"111100111",
  60438=>"010000001",
  60439=>"001000101",
  60440=>"101001001",
  60441=>"001000011",
  60442=>"101000110",
  60443=>"111001010",
  60444=>"111100111",
  60445=>"101010011",
  60446=>"001101001",
  60447=>"000100000",
  60448=>"110000100",
  60449=>"110011111",
  60450=>"110001100",
  60451=>"011101110",
  60452=>"100111101",
  60453=>"110011000",
  60454=>"110110111",
  60455=>"001000110",
  60456=>"010001010",
  60457=>"001101101",
  60458=>"010101001",
  60459=>"001011010",
  60460=>"101110011",
  60461=>"111001111",
  60462=>"000010111",
  60463=>"100100010",
  60464=>"010111100",
  60465=>"110000101",
  60466=>"111100001",
  60467=>"101001000",
  60468=>"111010011",
  60469=>"111111110",
  60470=>"110010101",
  60471=>"011111010",
  60472=>"010100001",
  60473=>"010011010",
  60474=>"111001010",
  60475=>"011011100",
  60476=>"011010011",
  60477=>"001111111",
  60478=>"010000011",
  60479=>"101001101",
  60480=>"011011100",
  60481=>"000010110",
  60482=>"111110000",
  60483=>"011000101",
  60484=>"101010110",
  60485=>"101000000",
  60486=>"010010011",
  60487=>"010011011",
  60488=>"100001001",
  60489=>"110010010",
  60490=>"110001000",
  60491=>"110011001",
  60492=>"010011111",
  60493=>"000010101",
  60494=>"001100000",
  60495=>"111000110",
  60496=>"100000110",
  60497=>"000101000",
  60498=>"100100111",
  60499=>"010101111",
  60500=>"110111001",
  60501=>"000001101",
  60502=>"011110110",
  60503=>"001011001",
  60504=>"010111001",
  60505=>"111111001",
  60506=>"000100000",
  60507=>"010111011",
  60508=>"111101100",
  60509=>"110000001",
  60510=>"101111011",
  60511=>"010110010",
  60512=>"011000001",
  60513=>"011100100",
  60514=>"101000010",
  60515=>"001010010",
  60516=>"101010001",
  60517=>"111101011",
  60518=>"011000010",
  60519=>"000110010",
  60520=>"100011101",
  60521=>"100010000",
  60522=>"000010011",
  60523=>"101001101",
  60524=>"101111010",
  60525=>"011100000",
  60526=>"010000110",
  60527=>"101011110",
  60528=>"110000100",
  60529=>"001001010",
  60530=>"101000111",
  60531=>"111101001",
  60532=>"001101110",
  60533=>"001100101",
  60534=>"111100000",
  60535=>"101110000",
  60536=>"010100100",
  60537=>"111111000",
  60538=>"000101010",
  60539=>"000110001",
  60540=>"111010111",
  60541=>"010000111",
  60542=>"001010111",
  60543=>"010110111",
  60544=>"100110100",
  60545=>"000001000",
  60546=>"100110101",
  60547=>"011110000",
  60548=>"111001110",
  60549=>"001111010",
  60550=>"101111000",
  60551=>"111011101",
  60552=>"111101011",
  60553=>"000010000",
  60554=>"110000100",
  60555=>"100001001",
  60556=>"111110001",
  60557=>"100101000",
  60558=>"101011101",
  60559=>"111010011",
  60560=>"011011101",
  60561=>"001101111",
  60562=>"001110101",
  60563=>"111111001",
  60564=>"111000100",
  60565=>"111000000",
  60566=>"000011001",
  60567=>"001001101",
  60568=>"101111101",
  60569=>"000010000",
  60570=>"001110111",
  60571=>"111101001",
  60572=>"101001101",
  60573=>"011100111",
  60574=>"101000001",
  60575=>"001100010",
  60576=>"011110011",
  60577=>"101001100",
  60578=>"010111101",
  60579=>"110010111",
  60580=>"001011110",
  60581=>"100100101",
  60582=>"100001001",
  60583=>"000000100",
  60584=>"101100010",
  60585=>"011010011",
  60586=>"101001110",
  60587=>"011010110",
  60588=>"001010011",
  60589=>"011110100",
  60590=>"010010000",
  60591=>"011000111",
  60592=>"001011100",
  60593=>"100110100",
  60594=>"100100101",
  60595=>"000110100",
  60596=>"001010101",
  60597=>"101001010",
  60598=>"010111010",
  60599=>"101100111",
  60600=>"110000000",
  60601=>"110101001",
  60602=>"000001000",
  60603=>"100011001",
  60604=>"000010111",
  60605=>"011000111",
  60606=>"101011001",
  60607=>"100111000",
  60608=>"001111011",
  60609=>"111011111",
  60610=>"111110100",
  60611=>"100110100",
  60612=>"111101000",
  60613=>"110001001",
  60614=>"011010110",
  60615=>"001000010",
  60616=>"110011000",
  60617=>"000100111",
  60618=>"011000100",
  60619=>"010110011",
  60620=>"101100001",
  60621=>"101101011",
  60622=>"000000001",
  60623=>"001001000",
  60624=>"010100010",
  60625=>"010111001",
  60626=>"000001100",
  60627=>"101110110",
  60628=>"101001000",
  60629=>"100100000",
  60630=>"000011100",
  60631=>"101001010",
  60632=>"100010101",
  60633=>"010110000",
  60634=>"110011010",
  60635=>"110000110",
  60636=>"001001110",
  60637=>"010000011",
  60638=>"011111110",
  60639=>"011010010",
  60640=>"000000001",
  60641=>"110100010",
  60642=>"111110101",
  60643=>"100001001",
  60644=>"100000110",
  60645=>"100011111",
  60646=>"001100000",
  60647=>"001011011",
  60648=>"101011001",
  60649=>"001001100",
  60650=>"100000011",
  60651=>"111110111",
  60652=>"101001101",
  60653=>"100000010",
  60654=>"111111110",
  60655=>"000010101",
  60656=>"111001000",
  60657=>"111111100",
  60658=>"011101001",
  60659=>"101110111",
  60660=>"011110000",
  60661=>"110101010",
  60662=>"000111101",
  60663=>"001010001",
  60664=>"110110110",
  60665=>"111100000",
  60666=>"101001111",
  60667=>"000111011",
  60668=>"110100110",
  60669=>"111111010",
  60670=>"010111110",
  60671=>"111000100",
  60672=>"110100001",
  60673=>"101111000",
  60674=>"100110101",
  60675=>"000110010",
  60676=>"111110111",
  60677=>"011101100",
  60678=>"010010000",
  60679=>"011010100",
  60680=>"111011011",
  60681=>"010111111",
  60682=>"110100101",
  60683=>"001011000",
  60684=>"000011101",
  60685=>"010011011",
  60686=>"000110010",
  60687=>"011110101",
  60688=>"110000101",
  60689=>"010010011",
  60690=>"001111100",
  60691=>"101110100",
  60692=>"100110110",
  60693=>"000001110",
  60694=>"011100000",
  60695=>"000100001",
  60696=>"101111110",
  60697=>"110001110",
  60698=>"101001011",
  60699=>"001110110",
  60700=>"000001000",
  60701=>"001001000",
  60702=>"100110101",
  60703=>"011011001",
  60704=>"000000010",
  60705=>"010011001",
  60706=>"100101011",
  60707=>"111110100",
  60708=>"001010010",
  60709=>"001101110",
  60710=>"111000100",
  60711=>"001110111",
  60712=>"000001101",
  60713=>"101010111",
  60714=>"010011100",
  60715=>"100010111",
  60716=>"110010111",
  60717=>"101000101",
  60718=>"010010101",
  60719=>"001010000",
  60720=>"010011101",
  60721=>"111101111",
  60722=>"001100000",
  60723=>"000010000",
  60724=>"010100100",
  60725=>"011101110",
  60726=>"000000110",
  60727=>"000001110",
  60728=>"101001000",
  60729=>"100101000",
  60730=>"101101111",
  60731=>"101101000",
  60732=>"011111010",
  60733=>"101111111",
  60734=>"100011111",
  60735=>"101001100",
  60736=>"100100100",
  60737=>"011011110",
  60738=>"110011010",
  60739=>"010100101",
  60740=>"011001000",
  60741=>"100010101",
  60742=>"000000001",
  60743=>"001011100",
  60744=>"100001010",
  60745=>"001000001",
  60746=>"001100110",
  60747=>"111100001",
  60748=>"011101100",
  60749=>"111100101",
  60750=>"110001100",
  60751=>"111011111",
  60752=>"100101110",
  60753=>"010100011",
  60754=>"001100110",
  60755=>"101100101",
  60756=>"110100110",
  60757=>"101110000",
  60758=>"111110100",
  60759=>"000100010",
  60760=>"010001000",
  60761=>"101111110",
  60762=>"011010100",
  60763=>"000111111",
  60764=>"001111111",
  60765=>"011010000",
  60766=>"111001010",
  60767=>"001110000",
  60768=>"100001001",
  60769=>"001001101",
  60770=>"111111110",
  60771=>"101110001",
  60772=>"101110111",
  60773=>"001000110",
  60774=>"011100010",
  60775=>"100001011",
  60776=>"000110000",
  60777=>"000000100",
  60778=>"010010111",
  60779=>"110101111",
  60780=>"001111100",
  60781=>"001001111",
  60782=>"000100000",
  60783=>"000100110",
  60784=>"111001101",
  60785=>"110101011",
  60786=>"001100011",
  60787=>"101100101",
  60788=>"001111001",
  60789=>"000011111",
  60790=>"011100000",
  60791=>"110010010",
  60792=>"000111001",
  60793=>"010111100",
  60794=>"100000010",
  60795=>"110110011",
  60796=>"000001000",
  60797=>"011110111",
  60798=>"000100100",
  60799=>"101111000",
  60800=>"100000001",
  60801=>"111110000",
  60802=>"010011010",
  60803=>"010010010",
  60804=>"000111011",
  60805=>"011111100",
  60806=>"101000011",
  60807=>"001011001",
  60808=>"110001111",
  60809=>"010101000",
  60810=>"110101001",
  60811=>"010101010",
  60812=>"101110111",
  60813=>"010101001",
  60814=>"110111110",
  60815=>"001100110",
  60816=>"111011110",
  60817=>"010001011",
  60818=>"101101001",
  60819=>"110001111",
  60820=>"000001101",
  60821=>"100000001",
  60822=>"110111111",
  60823=>"110001111",
  60824=>"000001010",
  60825=>"011001000",
  60826=>"000000010",
  60827=>"001110011",
  60828=>"000000000",
  60829=>"111000000",
  60830=>"101000001",
  60831=>"000000111",
  60832=>"100101000",
  60833=>"011111111",
  60834=>"111110011",
  60835=>"001111000",
  60836=>"001000100",
  60837=>"000000011",
  60838=>"100110110",
  60839=>"011011011",
  60840=>"111001011",
  60841=>"001100011",
  60842=>"000011011",
  60843=>"010010011",
  60844=>"011001011",
  60845=>"001110010",
  60846=>"101000100",
  60847=>"011101011",
  60848=>"010001100",
  60849=>"000010001",
  60850=>"110111000",
  60851=>"101001001",
  60852=>"011001111",
  60853=>"001011001",
  60854=>"111111100",
  60855=>"011011011",
  60856=>"011111111",
  60857=>"111011010",
  60858=>"101010110",
  60859=>"110011010",
  60860=>"110101010",
  60861=>"000101101",
  60862=>"001011001",
  60863=>"001100111",
  60864=>"111011000",
  60865=>"000000110",
  60866=>"101010100",
  60867=>"110101010",
  60868=>"101001000",
  60869=>"001110001",
  60870=>"110010000",
  60871=>"110101001",
  60872=>"110100000",
  60873=>"111100100",
  60874=>"111000110",
  60875=>"001000010",
  60876=>"100100110",
  60877=>"101110001",
  60878=>"110010100",
  60879=>"001011111",
  60880=>"100001010",
  60881=>"010011011",
  60882=>"011110100",
  60883=>"001000110",
  60884=>"111111000",
  60885=>"001010010",
  60886=>"000010000",
  60887=>"001010010",
  60888=>"111101101",
  60889=>"000010000",
  60890=>"101011110",
  60891=>"001111010",
  60892=>"000101001",
  60893=>"011100000",
  60894=>"011011010",
  60895=>"001000100",
  60896=>"011010110",
  60897=>"110110000",
  60898=>"101011100",
  60899=>"111000100",
  60900=>"001011001",
  60901=>"011001000",
  60902=>"001100001",
  60903=>"101001101",
  60904=>"100000011",
  60905=>"100000110",
  60906=>"000111000",
  60907=>"110110101",
  60908=>"000100101",
  60909=>"001000110",
  60910=>"000100111",
  60911=>"001100000",
  60912=>"000100101",
  60913=>"001001011",
  60914=>"110010011",
  60915=>"001001001",
  60916=>"110000001",
  60917=>"110001100",
  60918=>"110000100",
  60919=>"110010001",
  60920=>"101111001",
  60921=>"111100111",
  60922=>"100010101",
  60923=>"000010010",
  60924=>"110011101",
  60925=>"010111110",
  60926=>"010011000",
  60927=>"110100001",
  60928=>"000001000",
  60929=>"000100001",
  60930=>"100110010",
  60931=>"001000000",
  60932=>"111011111",
  60933=>"111100000",
  60934=>"000001001",
  60935=>"110010100",
  60936=>"011010011",
  60937=>"010010101",
  60938=>"010100010",
  60939=>"000011011",
  60940=>"000001010",
  60941=>"011111011",
  60942=>"011001001",
  60943=>"011011010",
  60944=>"011100110",
  60945=>"110101110",
  60946=>"001000000",
  60947=>"010001010",
  60948=>"100001000",
  60949=>"011010111",
  60950=>"010010000",
  60951=>"010101111",
  60952=>"110010000",
  60953=>"001111011",
  60954=>"111010001",
  60955=>"100100101",
  60956=>"001001000",
  60957=>"110011110",
  60958=>"011111001",
  60959=>"001000001",
  60960=>"001010011",
  60961=>"110110011",
  60962=>"001101100",
  60963=>"110011101",
  60964=>"010101101",
  60965=>"111111110",
  60966=>"111111010",
  60967=>"111010111",
  60968=>"001000101",
  60969=>"111100101",
  60970=>"001010010",
  60971=>"001110111",
  60972=>"011100001",
  60973=>"111101011",
  60974=>"110111110",
  60975=>"000110111",
  60976=>"001011101",
  60977=>"110101001",
  60978=>"110000101",
  60979=>"111001001",
  60980=>"111010101",
  60981=>"011001100",
  60982=>"110101011",
  60983=>"111011011",
  60984=>"101000000",
  60985=>"001101010",
  60986=>"000011000",
  60987=>"010111101",
  60988=>"100011001",
  60989=>"111011000",
  60990=>"001101001",
  60991=>"010010001",
  60992=>"100000100",
  60993=>"000111100",
  60994=>"111010010",
  60995=>"010111101",
  60996=>"100111010",
  60997=>"111101001",
  60998=>"001101000",
  60999=>"111010111",
  61000=>"010001011",
  61001=>"110111010",
  61002=>"100011100",
  61003=>"100001100",
  61004=>"101010100",
  61005=>"101100101",
  61006=>"101000000",
  61007=>"000010000",
  61008=>"111100110",
  61009=>"100011001",
  61010=>"100101111",
  61011=>"011000001",
  61012=>"000010000",
  61013=>"011100001",
  61014=>"110000000",
  61015=>"011111111",
  61016=>"011111010",
  61017=>"100110100",
  61018=>"101000010",
  61019=>"111101111",
  61020=>"010010010",
  61021=>"111011101",
  61022=>"100100100",
  61023=>"011011101",
  61024=>"011111011",
  61025=>"110011101",
  61026=>"100111111",
  61027=>"011010000",
  61028=>"001100010",
  61029=>"111011011",
  61030=>"100011110",
  61031=>"010011010",
  61032=>"110111010",
  61033=>"011110101",
  61034=>"010110110",
  61035=>"010000100",
  61036=>"100001000",
  61037=>"010000000",
  61038=>"101110001",
  61039=>"001101111",
  61040=>"110011010",
  61041=>"110011000",
  61042=>"111011100",
  61043=>"001111010",
  61044=>"100000001",
  61045=>"111011000",
  61046=>"010111010",
  61047=>"010011111",
  61048=>"010011111",
  61049=>"001110110",
  61050=>"010101111",
  61051=>"000100110",
  61052=>"011100000",
  61053=>"111101111",
  61054=>"110100011",
  61055=>"111100101",
  61056=>"011110001",
  61057=>"100101111",
  61058=>"011011001",
  61059=>"010001100",
  61060=>"110011001",
  61061=>"001101010",
  61062=>"010000100",
  61063=>"011010000",
  61064=>"110111111",
  61065=>"000010101",
  61066=>"010100110",
  61067=>"010011011",
  61068=>"100111000",
  61069=>"111100110",
  61070=>"100101010",
  61071=>"011010101",
  61072=>"111001101",
  61073=>"100011010",
  61074=>"011101010",
  61075=>"111010010",
  61076=>"100101011",
  61077=>"111011101",
  61078=>"011101110",
  61079=>"111010101",
  61080=>"000010101",
  61081=>"110001000",
  61082=>"110011111",
  61083=>"011111001",
  61084=>"011101011",
  61085=>"110010011",
  61086=>"011110010",
  61087=>"010010110",
  61088=>"110111111",
  61089=>"100101011",
  61090=>"000000101",
  61091=>"101010000",
  61092=>"100010001",
  61093=>"000111101",
  61094=>"011111100",
  61095=>"010010100",
  61096=>"011110010",
  61097=>"000100000",
  61098=>"101100111",
  61099=>"100011111",
  61100=>"000001100",
  61101=>"100000111",
  61102=>"100100101",
  61103=>"000001011",
  61104=>"000100011",
  61105=>"000011101",
  61106=>"101110011",
  61107=>"111100110",
  61108=>"010001011",
  61109=>"010100111",
  61110=>"110101001",
  61111=>"011001000",
  61112=>"010111101",
  61113=>"100000111",
  61114=>"010000000",
  61115=>"011010101",
  61116=>"000011101",
  61117=>"010000010",
  61118=>"001110111",
  61119=>"110110000",
  61120=>"110010110",
  61121=>"101100111",
  61122=>"101100100",
  61123=>"000010001",
  61124=>"011110010",
  61125=>"000101010",
  61126=>"110110110",
  61127=>"100110101",
  61128=>"101001100",
  61129=>"000010101",
  61130=>"101101000",
  61131=>"111010010",
  61132=>"110101011",
  61133=>"001111110",
  61134=>"000010100",
  61135=>"110001111",
  61136=>"110101011",
  61137=>"111001101",
  61138=>"101010001",
  61139=>"111111001",
  61140=>"001100000",
  61141=>"111111111",
  61142=>"100100011",
  61143=>"000100010",
  61144=>"001100110",
  61145=>"101101010",
  61146=>"001000010",
  61147=>"100100011",
  61148=>"001001001",
  61149=>"000011101",
  61150=>"110000001",
  61151=>"110010111",
  61152=>"101000101",
  61153=>"100001101",
  61154=>"010101111",
  61155=>"000001011",
  61156=>"000000000",
  61157=>"101101010",
  61158=>"100100000",
  61159=>"110110110",
  61160=>"001111111",
  61161=>"011111100",
  61162=>"001000110",
  61163=>"111011101",
  61164=>"101010000",
  61165=>"011110101",
  61166=>"100100100",
  61167=>"101001110",
  61168=>"000101001",
  61169=>"010100000",
  61170=>"110101010",
  61171=>"111111010",
  61172=>"110101010",
  61173=>"101010111",
  61174=>"111110001",
  61175=>"000000110",
  61176=>"000100001",
  61177=>"010001100",
  61178=>"110110000",
  61179=>"011000011",
  61180=>"111100100",
  61181=>"101111100",
  61182=>"000010000",
  61183=>"000100111",
  61184=>"011001011",
  61185=>"110010100",
  61186=>"110001101",
  61187=>"111110101",
  61188=>"110010000",
  61189=>"111010000",
  61190=>"011000100",
  61191=>"011000110",
  61192=>"010011111",
  61193=>"101011111",
  61194=>"011110001",
  61195=>"010110101",
  61196=>"011011100",
  61197=>"010011100",
  61198=>"001011001",
  61199=>"111001101",
  61200=>"101110110",
  61201=>"101010111",
  61202=>"101011101",
  61203=>"110000100",
  61204=>"001110000",
  61205=>"010000000",
  61206=>"101011100",
  61207=>"000001001",
  61208=>"111001001",
  61209=>"100101111",
  61210=>"001101110",
  61211=>"110110010",
  61212=>"100111101",
  61213=>"110110101",
  61214=>"001101000",
  61215=>"011011111",
  61216=>"000010010",
  61217=>"111100010",
  61218=>"101011110",
  61219=>"110101100",
  61220=>"011100110",
  61221=>"100000101",
  61222=>"001100111",
  61223=>"010001001",
  61224=>"011100110",
  61225=>"101011011",
  61226=>"111000100",
  61227=>"110101100",
  61228=>"101000110",
  61229=>"110111010",
  61230=>"000000000",
  61231=>"011111101",
  61232=>"010010001",
  61233=>"001001100",
  61234=>"010100001",
  61235=>"010111001",
  61236=>"011111000",
  61237=>"001001011",
  61238=>"101101000",
  61239=>"111011100",
  61240=>"111111001",
  61241=>"001101110",
  61242=>"111011000",
  61243=>"111010100",
  61244=>"110010010",
  61245=>"010101110",
  61246=>"001011010",
  61247=>"111110000",
  61248=>"010100101",
  61249=>"010100010",
  61250=>"110101000",
  61251=>"001110000",
  61252=>"001100011",
  61253=>"000110100",
  61254=>"110001100",
  61255=>"001111000",
  61256=>"110100011",
  61257=>"010011110",
  61258=>"111000011",
  61259=>"000001011",
  61260=>"011110000",
  61261=>"000011010",
  61262=>"010110100",
  61263=>"000011111",
  61264=>"001010001",
  61265=>"000010110",
  61266=>"010100101",
  61267=>"101000010",
  61268=>"010111000",
  61269=>"100101000",
  61270=>"100111101",
  61271=>"100001101",
  61272=>"100110100",
  61273=>"010110010",
  61274=>"110000111",
  61275=>"111011101",
  61276=>"010111101",
  61277=>"000010001",
  61278=>"011111111",
  61279=>"011010001",
  61280=>"101100111",
  61281=>"000001110",
  61282=>"100111011",
  61283=>"000010001",
  61284=>"100010000",
  61285=>"010100111",
  61286=>"111010101",
  61287=>"100010011",
  61288=>"101111011",
  61289=>"111000001",
  61290=>"011000011",
  61291=>"101110110",
  61292=>"111110110",
  61293=>"111000001",
  61294=>"101011100",
  61295=>"110111100",
  61296=>"100010100",
  61297=>"000010110",
  61298=>"000000010",
  61299=>"010010000",
  61300=>"000110010",
  61301=>"110001000",
  61302=>"110110001",
  61303=>"011001101",
  61304=>"001100100",
  61305=>"111111010",
  61306=>"000001010",
  61307=>"101111100",
  61308=>"001111100",
  61309=>"000111111",
  61310=>"111001111",
  61311=>"111111110",
  61312=>"001110001",
  61313=>"100100011",
  61314=>"001110110",
  61315=>"110111110",
  61316=>"110010101",
  61317=>"010111100",
  61318=>"010101001",
  61319=>"110000011",
  61320=>"100111110",
  61321=>"001111101",
  61322=>"011111001",
  61323=>"011010001",
  61324=>"110100001",
  61325=>"110101100",
  61326=>"000011110",
  61327=>"111101101",
  61328=>"000000010",
  61329=>"001011111",
  61330=>"110001100",
  61331=>"110001100",
  61332=>"011110000",
  61333=>"011011110",
  61334=>"010100010",
  61335=>"011010001",
  61336=>"010110101",
  61337=>"011000000",
  61338=>"101100011",
  61339=>"010010001",
  61340=>"010100101",
  61341=>"010011111",
  61342=>"010100000",
  61343=>"111111111",
  61344=>"101101000",
  61345=>"101001101",
  61346=>"011101111",
  61347=>"000110101",
  61348=>"101000010",
  61349=>"110100010",
  61350=>"110011010",
  61351=>"111000001",
  61352=>"011101001",
  61353=>"111001000",
  61354=>"110111011",
  61355=>"100011100",
  61356=>"111000000",
  61357=>"111001010",
  61358=>"110100001",
  61359=>"010111100",
  61360=>"111000111",
  61361=>"011111101",
  61362=>"110111100",
  61363=>"110011110",
  61364=>"100110011",
  61365=>"100111000",
  61366=>"101110111",
  61367=>"000001101",
  61368=>"101000000",
  61369=>"001001101",
  61370=>"010111000",
  61371=>"011111000",
  61372=>"111111000",
  61373=>"110011111",
  61374=>"110000101",
  61375=>"100010111",
  61376=>"000001111",
  61377=>"100100100",
  61378=>"011011111",
  61379=>"000011001",
  61380=>"000111011",
  61381=>"100010111",
  61382=>"011000111",
  61383=>"000100001",
  61384=>"110101000",
  61385=>"010110000",
  61386=>"110010111",
  61387=>"100010111",
  61388=>"110111111",
  61389=>"101001110",
  61390=>"000110000",
  61391=>"000101011",
  61392=>"110100110",
  61393=>"101010000",
  61394=>"101100111",
  61395=>"100111010",
  61396=>"101010010",
  61397=>"101001110",
  61398=>"010110000",
  61399=>"011001001",
  61400=>"001000100",
  61401=>"100001001",
  61402=>"001101111",
  61403=>"010000100",
  61404=>"101101000",
  61405=>"110100111",
  61406=>"110100101",
  61407=>"101000100",
  61408=>"001110000",
  61409=>"010011001",
  61410=>"000100100",
  61411=>"100010100",
  61412=>"001001000",
  61413=>"110000001",
  61414=>"001100101",
  61415=>"001110010",
  61416=>"001111110",
  61417=>"001111100",
  61418=>"110101000",
  61419=>"010011001",
  61420=>"011011010",
  61421=>"000000010",
  61422=>"011111000",
  61423=>"111110110",
  61424=>"101100000",
  61425=>"001110111",
  61426=>"010011000",
  61427=>"010000000",
  61428=>"000011111",
  61429=>"010011010",
  61430=>"000011000",
  61431=>"000011001",
  61432=>"101100101",
  61433=>"111111000",
  61434=>"000001010",
  61435=>"111111001",
  61436=>"110010000",
  61437=>"010011101",
  61438=>"111010000",
  61439=>"110110001",
  61440=>"111101110",
  61441=>"011000111",
  61442=>"010010011",
  61443=>"011000001",
  61444=>"110001100",
  61445=>"100110111",
  61446=>"111100101",
  61447=>"101011101",
  61448=>"100101111",
  61449=>"110101011",
  61450=>"000010101",
  61451=>"010000110",
  61452=>"111110101",
  61453=>"000001101",
  61454=>"001111011",
  61455=>"101101101",
  61456=>"011111001",
  61457=>"100101111",
  61458=>"001000001",
  61459=>"111000010",
  61460=>"100001110",
  61461=>"101000100",
  61462=>"010110000",
  61463=>"100100100",
  61464=>"110111100",
  61465=>"101101011",
  61466=>"011011001",
  61467=>"000110011",
  61468=>"101001111",
  61469=>"101001100",
  61470=>"100110110",
  61471=>"110000000",
  61472=>"010010110",
  61473=>"010011111",
  61474=>"100100111",
  61475=>"100110101",
  61476=>"010101110",
  61477=>"000011110",
  61478=>"010001101",
  61479=>"001101111",
  61480=>"000001101",
  61481=>"000100000",
  61482=>"101000101",
  61483=>"010011111",
  61484=>"100010101",
  61485=>"000110110",
  61486=>"100011000",
  61487=>"000011011",
  61488=>"110011000",
  61489=>"001100010",
  61490=>"000111010",
  61491=>"100010100",
  61492=>"011000000",
  61493=>"000011000",
  61494=>"110010100",
  61495=>"010011100",
  61496=>"100010000",
  61497=>"101010001",
  61498=>"111111101",
  61499=>"101100101",
  61500=>"011101010",
  61501=>"000100110",
  61502=>"110000000",
  61503=>"001011000",
  61504=>"000000010",
  61505=>"000101000",
  61506=>"001101100",
  61507=>"011010101",
  61508=>"000001101",
  61509=>"010111011",
  61510=>"000111010",
  61511=>"010111011",
  61512=>"100110011",
  61513=>"010010001",
  61514=>"001000101",
  61515=>"100000101",
  61516=>"100110100",
  61517=>"011010111",
  61518=>"001011110",
  61519=>"100110110",
  61520=>"000111000",
  61521=>"011000001",
  61522=>"110011001",
  61523=>"100101110",
  61524=>"101111111",
  61525=>"110110001",
  61526=>"100000111",
  61527=>"001001001",
  61528=>"111011101",
  61529=>"010001011",
  61530=>"101000001",
  61531=>"101110100",
  61532=>"001100011",
  61533=>"000010000",
  61534=>"100000001",
  61535=>"111110011",
  61536=>"000110010",
  61537=>"111111010",
  61538=>"010011100",
  61539=>"010100000",
  61540=>"001001100",
  61541=>"100000101",
  61542=>"100111010",
  61543=>"100000001",
  61544=>"010111000",
  61545=>"100011101",
  61546=>"111101110",
  61547=>"000010111",
  61548=>"000111100",
  61549=>"011000110",
  61550=>"011101101",
  61551=>"001001000",
  61552=>"101100011",
  61553=>"100110100",
  61554=>"101111110",
  61555=>"111111010",
  61556=>"001000110",
  61557=>"010111110",
  61558=>"001011111",
  61559=>"100111101",
  61560=>"111100010",
  61561=>"001001001",
  61562=>"100011101",
  61563=>"010010111",
  61564=>"000001110",
  61565=>"100010101",
  61566=>"010101000",
  61567=>"110000100",
  61568=>"000000110",
  61569=>"111100000",
  61570=>"100000111",
  61571=>"100001110",
  61572=>"100001000",
  61573=>"000001010",
  61574=>"100000000",
  61575=>"011010001",
  61576=>"000001111",
  61577=>"111000110",
  61578=>"001011011",
  61579=>"101101110",
  61580=>"111111010",
  61581=>"001111111",
  61582=>"100111101",
  61583=>"101110101",
  61584=>"001011110",
  61585=>"101000111",
  61586=>"000100000",
  61587=>"110110011",
  61588=>"110001011",
  61589=>"000110011",
  61590=>"101010110",
  61591=>"011000110",
  61592=>"111010010",
  61593=>"111001000",
  61594=>"101110101",
  61595=>"000010000",
  61596=>"101111101",
  61597=>"100101101",
  61598=>"100110111",
  61599=>"111111111",
  61600=>"001110001",
  61601=>"011110101",
  61602=>"010010101",
  61603=>"100011100",
  61604=>"100101000",
  61605=>"011001110",
  61606=>"100111111",
  61607=>"111000000",
  61608=>"000110101",
  61609=>"001000000",
  61610=>"000111000",
  61611=>"000111011",
  61612=>"011110101",
  61613=>"100000010",
  61614=>"100011000",
  61615=>"000110010",
  61616=>"100100101",
  61617=>"100000010",
  61618=>"100001000",
  61619=>"000001111",
  61620=>"000100001",
  61621=>"100100011",
  61622=>"101110110",
  61623=>"011010000",
  61624=>"111100011",
  61625=>"100001000",
  61626=>"111000010",
  61627=>"010110100",
  61628=>"111000101",
  61629=>"011000001",
  61630=>"111100110",
  61631=>"101000011",
  61632=>"010001011",
  61633=>"100101001",
  61634=>"001000101",
  61635=>"011000000",
  61636=>"010111101",
  61637=>"100111101",
  61638=>"000101010",
  61639=>"101101000",
  61640=>"100111111",
  61641=>"001001100",
  61642=>"101100100",
  61643=>"010010100",
  61644=>"110001100",
  61645=>"111101101",
  61646=>"011010000",
  61647=>"111110111",
  61648=>"011101110",
  61649=>"110000110",
  61650=>"010101011",
  61651=>"011111011",
  61652=>"011000110",
  61653=>"110010111",
  61654=>"101100011",
  61655=>"101101010",
  61656=>"110001111",
  61657=>"001111101",
  61658=>"110111001",
  61659=>"011110111",
  61660=>"111011111",
  61661=>"000101000",
  61662=>"101110101",
  61663=>"001000010",
  61664=>"100111110",
  61665=>"010111000",
  61666=>"101110111",
  61667=>"010110100",
  61668=>"001000000",
  61669=>"001101001",
  61670=>"111101111",
  61671=>"101101110",
  61672=>"000110101",
  61673=>"101111001",
  61674=>"110101110",
  61675=>"110111000",
  61676=>"001111100",
  61677=>"111000100",
  61678=>"000001010",
  61679=>"011001101",
  61680=>"000010010",
  61681=>"000000000",
  61682=>"100001110",
  61683=>"101001111",
  61684=>"101001001",
  61685=>"100000001",
  61686=>"000001110",
  61687=>"100101011",
  61688=>"011010010",
  61689=>"001100010",
  61690=>"010111110",
  61691=>"010110101",
  61692=>"111011111",
  61693=>"010010000",
  61694=>"110101101",
  61695=>"110100110",
  61696=>"001100011",
  61697=>"000100100",
  61698=>"110110011",
  61699=>"001000001",
  61700=>"000001110",
  61701=>"110010001",
  61702=>"101000001",
  61703=>"111000110",
  61704=>"111110101",
  61705=>"100101101",
  61706=>"000011111",
  61707=>"001001101",
  61708=>"011010010",
  61709=>"101110010",
  61710=>"101110000",
  61711=>"010010010",
  61712=>"011111000",
  61713=>"110101100",
  61714=>"111110100",
  61715=>"001011010",
  61716=>"101000001",
  61717=>"011000100",
  61718=>"000001110",
  61719=>"010010000",
  61720=>"110010001",
  61721=>"100001100",
  61722=>"000110100",
  61723=>"010000011",
  61724=>"100011001",
  61725=>"000111111",
  61726=>"111110100",
  61727=>"110100010",
  61728=>"000000110",
  61729=>"101010100",
  61730=>"111101100",
  61731=>"011000110",
  61732=>"010000010",
  61733=>"001100101",
  61734=>"010001000",
  61735=>"100000000",
  61736=>"111000111",
  61737=>"001011101",
  61738=>"011101000",
  61739=>"011000000",
  61740=>"001010111",
  61741=>"001100101",
  61742=>"000001001",
  61743=>"100100111",
  61744=>"001001001",
  61745=>"100011110",
  61746=>"001011110",
  61747=>"111100101",
  61748=>"000010110",
  61749=>"000000111",
  61750=>"111010110",
  61751=>"101111101",
  61752=>"000010001",
  61753=>"101101110",
  61754=>"001100110",
  61755=>"110101111",
  61756=>"100111010",
  61757=>"101101110",
  61758=>"100111101",
  61759=>"011001001",
  61760=>"000011110",
  61761=>"100111110",
  61762=>"110101101",
  61763=>"010011111",
  61764=>"000000010",
  61765=>"111011010",
  61766=>"000001111",
  61767=>"101110110",
  61768=>"010010010",
  61769=>"001001010",
  61770=>"011101110",
  61771=>"111110001",
  61772=>"000001001",
  61773=>"000010010",
  61774=>"000001111",
  61775=>"001010111",
  61776=>"000001101",
  61777=>"011000110",
  61778=>"101010011",
  61779=>"101011000",
  61780=>"101101011",
  61781=>"001010000",
  61782=>"001010011",
  61783=>"011111000",
  61784=>"011000110",
  61785=>"110000000",
  61786=>"001100010",
  61787=>"000100000",
  61788=>"000000100",
  61789=>"000000100",
  61790=>"010001111",
  61791=>"100110010",
  61792=>"000101100",
  61793=>"001010101",
  61794=>"111101100",
  61795=>"001110010",
  61796=>"111110101",
  61797=>"101111010",
  61798=>"010101111",
  61799=>"100011011",
  61800=>"011001010",
  61801=>"000001001",
  61802=>"001100001",
  61803=>"100010000",
  61804=>"100010011",
  61805=>"011110110",
  61806=>"011110100",
  61807=>"101100001",
  61808=>"000100101",
  61809=>"101000100",
  61810=>"010001001",
  61811=>"001111010",
  61812=>"001101000",
  61813=>"101000010",
  61814=>"010111111",
  61815=>"000010001",
  61816=>"101000001",
  61817=>"110100010",
  61818=>"110100100",
  61819=>"110111010",
  61820=>"110010100",
  61821=>"000000110",
  61822=>"000000011",
  61823=>"000000000",
  61824=>"100011101",
  61825=>"110110110",
  61826=>"100111111",
  61827=>"100111100",
  61828=>"010100101",
  61829=>"011110011",
  61830=>"110000000",
  61831=>"110100011",
  61832=>"011001100",
  61833=>"000010110",
  61834=>"110010110",
  61835=>"010000001",
  61836=>"111001111",
  61837=>"011001001",
  61838=>"011101011",
  61839=>"101010101",
  61840=>"100011000",
  61841=>"100110010",
  61842=>"100111111",
  61843=>"011101111",
  61844=>"011010100",
  61845=>"000110001",
  61846=>"111101111",
  61847=>"110000011",
  61848=>"111001011",
  61849=>"101110101",
  61850=>"011100111",
  61851=>"111101001",
  61852=>"111100110",
  61853=>"110101000",
  61854=>"110000000",
  61855=>"011100110",
  61856=>"101101101",
  61857=>"110100001",
  61858=>"101000100",
  61859=>"011000000",
  61860=>"010001000",
  61861=>"000011100",
  61862=>"010100011",
  61863=>"001100111",
  61864=>"010101011",
  61865=>"001001101",
  61866=>"101111001",
  61867=>"100110010",
  61868=>"000000011",
  61869=>"100111011",
  61870=>"101011111",
  61871=>"100000001",
  61872=>"101001011",
  61873=>"110001110",
  61874=>"001001000",
  61875=>"101110100",
  61876=>"010010110",
  61877=>"010000000",
  61878=>"011110001",
  61879=>"101111111",
  61880=>"111010001",
  61881=>"110001111",
  61882=>"101101000",
  61883=>"000001011",
  61884=>"101001000",
  61885=>"100000100",
  61886=>"101100011",
  61887=>"101110110",
  61888=>"110011001",
  61889=>"100000001",
  61890=>"100101110",
  61891=>"101111001",
  61892=>"010010000",
  61893=>"011000000",
  61894=>"000100100",
  61895=>"001110010",
  61896=>"011001010",
  61897=>"001110000",
  61898=>"101011100",
  61899=>"111011000",
  61900=>"101010000",
  61901=>"001111101",
  61902=>"010000010",
  61903=>"010011000",
  61904=>"101111001",
  61905=>"101101110",
  61906=>"011001011",
  61907=>"011110101",
  61908=>"000010011",
  61909=>"000111111",
  61910=>"010010001",
  61911=>"000000110",
  61912=>"011010111",
  61913=>"111100010",
  61914=>"010000110",
  61915=>"101001000",
  61916=>"010011100",
  61917=>"100000111",
  61918=>"100100111",
  61919=>"111001100",
  61920=>"101100000",
  61921=>"111010100",
  61922=>"001011111",
  61923=>"000111011",
  61924=>"111111111",
  61925=>"010001100",
  61926=>"001000001",
  61927=>"010010010",
  61928=>"000000110",
  61929=>"010100100",
  61930=>"110100000",
  61931=>"001111110",
  61932=>"000001111",
  61933=>"000000001",
  61934=>"111100010",
  61935=>"011110111",
  61936=>"100111000",
  61937=>"101100111",
  61938=>"111001101",
  61939=>"100100000",
  61940=>"011101010",
  61941=>"001101111",
  61942=>"100101111",
  61943=>"011010111",
  61944=>"100101110",
  61945=>"000101011",
  61946=>"100100010",
  61947=>"011101001",
  61948=>"011001110",
  61949=>"111110001",
  61950=>"100001110",
  61951=>"000000100",
  61952=>"110111001",
  61953=>"110111111",
  61954=>"101111011",
  61955=>"010101101",
  61956=>"111111101",
  61957=>"100101001",
  61958=>"110111000",
  61959=>"010110000",
  61960=>"010010101",
  61961=>"100100010",
  61962=>"110110011",
  61963=>"101101000",
  61964=>"001111101",
  61965=>"111111111",
  61966=>"000000000",
  61967=>"110011110",
  61968=>"011010010",
  61969=>"110000100",
  61970=>"011011010",
  61971=>"100011100",
  61972=>"000011101",
  61973=>"000011011",
  61974=>"110011011",
  61975=>"011101101",
  61976=>"000000111",
  61977=>"111000110",
  61978=>"010101100",
  61979=>"101001110",
  61980=>"101101000",
  61981=>"011001101",
  61982=>"100010101",
  61983=>"110110100",
  61984=>"001001111",
  61985=>"110110110",
  61986=>"000000101",
  61987=>"110100110",
  61988=>"001011110",
  61989=>"100011011",
  61990=>"001001000",
  61991=>"110100110",
  61992=>"100010010",
  61993=>"101110000",
  61994=>"001001011",
  61995=>"000000000",
  61996=>"011010000",
  61997=>"100011110",
  61998=>"000010010",
  61999=>"001000000",
  62000=>"100101101",
  62001=>"000011010",
  62002=>"110100011",
  62003=>"111100100",
  62004=>"110001100",
  62005=>"011101110",
  62006=>"100110101",
  62007=>"001100010",
  62008=>"100111100",
  62009=>"111111101",
  62010=>"010100100",
  62011=>"011110001",
  62012=>"111000110",
  62013=>"110010110",
  62014=>"011011001",
  62015=>"000001100",
  62016=>"010101011",
  62017=>"000111110",
  62018=>"011001001",
  62019=>"000011110",
  62020=>"101010111",
  62021=>"111011111",
  62022=>"001100001",
  62023=>"110111011",
  62024=>"010100100",
  62025=>"000110100",
  62026=>"111100100",
  62027=>"011110011",
  62028=>"000001000",
  62029=>"100110100",
  62030=>"001110000",
  62031=>"011000111",
  62032=>"010100100",
  62033=>"100000110",
  62034=>"010000011",
  62035=>"000011000",
  62036=>"100110001",
  62037=>"110101000",
  62038=>"111101100",
  62039=>"110000010",
  62040=>"000010110",
  62041=>"001010000",
  62042=>"100100000",
  62043=>"000000001",
  62044=>"101111000",
  62045=>"101110010",
  62046=>"001110110",
  62047=>"100111110",
  62048=>"000011000",
  62049=>"000111000",
  62050=>"100100000",
  62051=>"000000101",
  62052=>"000011111",
  62053=>"011000100",
  62054=>"000011111",
  62055=>"100111010",
  62056=>"001011010",
  62057=>"111111010",
  62058=>"111101011",
  62059=>"111110101",
  62060=>"111000111",
  62061=>"010011110",
  62062=>"111001001",
  62063=>"001010110",
  62064=>"111111000",
  62065=>"111101101",
  62066=>"100111110",
  62067=>"000101010",
  62068=>"111111110",
  62069=>"010000001",
  62070=>"101111111",
  62071=>"110100001",
  62072=>"101000010",
  62073=>"000110111",
  62074=>"000101110",
  62075=>"000100001",
  62076=>"010010010",
  62077=>"001000011",
  62078=>"110111011",
  62079=>"011001011",
  62080=>"101100100",
  62081=>"110001101",
  62082=>"001101001",
  62083=>"001001000",
  62084=>"111100011",
  62085=>"001110000",
  62086=>"101110101",
  62087=>"000010101",
  62088=>"111010011",
  62089=>"000010010",
  62090=>"000100010",
  62091=>"011011100",
  62092=>"000000010",
  62093=>"111000011",
  62094=>"000110111",
  62095=>"111111110",
  62096=>"101111111",
  62097=>"101010111",
  62098=>"100010011",
  62099=>"010000000",
  62100=>"000000100",
  62101=>"010001011",
  62102=>"001100011",
  62103=>"110100000",
  62104=>"011000010",
  62105=>"000100001",
  62106=>"010000000",
  62107=>"110000110",
  62108=>"000001101",
  62109=>"110011000",
  62110=>"101110111",
  62111=>"000010001",
  62112=>"011000000",
  62113=>"010001000",
  62114=>"000110111",
  62115=>"100011010",
  62116=>"100000110",
  62117=>"101111010",
  62118=>"001010000",
  62119=>"010000100",
  62120=>"100001101",
  62121=>"110110110",
  62122=>"001100111",
  62123=>"101100001",
  62124=>"110010010",
  62125=>"011011100",
  62126=>"101010010",
  62127=>"000010010",
  62128=>"100101111",
  62129=>"110100111",
  62130=>"111001010",
  62131=>"110111010",
  62132=>"110001001",
  62133=>"001000101",
  62134=>"111010100",
  62135=>"001100111",
  62136=>"000000110",
  62137=>"011010111",
  62138=>"000001011",
  62139=>"011011000",
  62140=>"010101000",
  62141=>"001001110",
  62142=>"001000100",
  62143=>"100110011",
  62144=>"100001110",
  62145=>"001101000",
  62146=>"100011110",
  62147=>"110110111",
  62148=>"000110111",
  62149=>"010010100",
  62150=>"011011010",
  62151=>"111110001",
  62152=>"110011001",
  62153=>"111010111",
  62154=>"111101100",
  62155=>"101110101",
  62156=>"111111010",
  62157=>"111001001",
  62158=>"110000111",
  62159=>"101101110",
  62160=>"010000011",
  62161=>"001010001",
  62162=>"011111111",
  62163=>"001100010",
  62164=>"000100001",
  62165=>"100110011",
  62166=>"010110011",
  62167=>"010110100",
  62168=>"111111001",
  62169=>"011110100",
  62170=>"000111111",
  62171=>"101000101",
  62172=>"100101101",
  62173=>"101011111",
  62174=>"011111000",
  62175=>"010111110",
  62176=>"100100110",
  62177=>"011001100",
  62178=>"000110110",
  62179=>"100100111",
  62180=>"010110100",
  62181=>"011101111",
  62182=>"001110101",
  62183=>"100111101",
  62184=>"010000010",
  62185=>"110011010",
  62186=>"000100000",
  62187=>"010010000",
  62188=>"000101101",
  62189=>"101111001",
  62190=>"010011011",
  62191=>"111010100",
  62192=>"001011101",
  62193=>"001111100",
  62194=>"100100100",
  62195=>"111011001",
  62196=>"111110110",
  62197=>"101101111",
  62198=>"100001001",
  62199=>"111101100",
  62200=>"101101000",
  62201=>"010011011",
  62202=>"010110111",
  62203=>"100001110",
  62204=>"100110111",
  62205=>"101001111",
  62206=>"000100110",
  62207=>"001011001",
  62208=>"010100100",
  62209=>"111011010",
  62210=>"110000000",
  62211=>"000110110",
  62212=>"001111010",
  62213=>"101111001",
  62214=>"110000011",
  62215=>"010101101",
  62216=>"000000100",
  62217=>"111100111",
  62218=>"010000101",
  62219=>"011000001",
  62220=>"111000000",
  62221=>"111101001",
  62222=>"111101000",
  62223=>"111011011",
  62224=>"110110000",
  62225=>"100100111",
  62226=>"000110111",
  62227=>"000010001",
  62228=>"011100000",
  62229=>"110010111",
  62230=>"101101110",
  62231=>"001000001",
  62232=>"101001011",
  62233=>"101100101",
  62234=>"001001110",
  62235=>"000100111",
  62236=>"101000011",
  62237=>"000011111",
  62238=>"111110111",
  62239=>"101101001",
  62240=>"001100010",
  62241=>"110001011",
  62242=>"000100000",
  62243=>"110111111",
  62244=>"101011001",
  62245=>"001000100",
  62246=>"100100010",
  62247=>"111110010",
  62248=>"110110101",
  62249=>"111110110",
  62250=>"110011100",
  62251=>"000001001",
  62252=>"111101001",
  62253=>"010110111",
  62254=>"001110110",
  62255=>"001100011",
  62256=>"101001111",
  62257=>"100110001",
  62258=>"111000110",
  62259=>"010010001",
  62260=>"000001010",
  62261=>"101101100",
  62262=>"111011101",
  62263=>"110000110",
  62264=>"100110000",
  62265=>"101101101",
  62266=>"011000000",
  62267=>"001111101",
  62268=>"011011001",
  62269=>"110000000",
  62270=>"001011001",
  62271=>"111001110",
  62272=>"111111100",
  62273=>"000001001",
  62274=>"001011011",
  62275=>"111001110",
  62276=>"111111001",
  62277=>"011100101",
  62278=>"101000101",
  62279=>"001110010",
  62280=>"011100011",
  62281=>"111100010",
  62282=>"100010000",
  62283=>"101001001",
  62284=>"001110101",
  62285=>"001100011",
  62286=>"011010000",
  62287=>"100111011",
  62288=>"101100100",
  62289=>"000101101",
  62290=>"100001111",
  62291=>"000100101",
  62292=>"100100100",
  62293=>"110011111",
  62294=>"000010010",
  62295=>"011011000",
  62296=>"111000010",
  62297=>"001110011",
  62298=>"100111110",
  62299=>"000011111",
  62300=>"100111101",
  62301=>"110100001",
  62302=>"110100110",
  62303=>"100010111",
  62304=>"010111100",
  62305=>"100000010",
  62306=>"101000001",
  62307=>"111111100",
  62308=>"111110010",
  62309=>"110110110",
  62310=>"001000011",
  62311=>"110011100",
  62312=>"100000100",
  62313=>"100001011",
  62314=>"001001000",
  62315=>"001101001",
  62316=>"010110011",
  62317=>"001001011",
  62318=>"101000000",
  62319=>"011011010",
  62320=>"100101110",
  62321=>"011110111",
  62322=>"100001101",
  62323=>"110111111",
  62324=>"001111000",
  62325=>"111101100",
  62326=>"011101001",
  62327=>"000010100",
  62328=>"011100110",
  62329=>"011110110",
  62330=>"101001000",
  62331=>"101010111",
  62332=>"111011101",
  62333=>"111011100",
  62334=>"101100111",
  62335=>"100001001",
  62336=>"001101001",
  62337=>"101010000",
  62338=>"001000000",
  62339=>"000001000",
  62340=>"010100101",
  62341=>"110011111",
  62342=>"101011010",
  62343=>"010101110",
  62344=>"000001001",
  62345=>"011011000",
  62346=>"010101010",
  62347=>"011010100",
  62348=>"000010100",
  62349=>"000111101",
  62350=>"100110111",
  62351=>"100011100",
  62352=>"000001100",
  62353=>"000010111",
  62354=>"000100000",
  62355=>"010100001",
  62356=>"000010000",
  62357=>"011100100",
  62358=>"101111011",
  62359=>"110000101",
  62360=>"001011011",
  62361=>"000010011",
  62362=>"010100010",
  62363=>"001110111",
  62364=>"100001000",
  62365=>"010011110",
  62366=>"011010011",
  62367=>"001001110",
  62368=>"010100000",
  62369=>"000001011",
  62370=>"011000101",
  62371=>"100110010",
  62372=>"110001001",
  62373=>"100110110",
  62374=>"001110111",
  62375=>"001001100",
  62376=>"001100111",
  62377=>"001101101",
  62378=>"101101011",
  62379=>"001111100",
  62380=>"111100111",
  62381=>"011001110",
  62382=>"000001000",
  62383=>"010010000",
  62384=>"111011011",
  62385=>"011000110",
  62386=>"000010100",
  62387=>"000111000",
  62388=>"101101000",
  62389=>"110000110",
  62390=>"000111001",
  62391=>"111111101",
  62392=>"110100110",
  62393=>"101010011",
  62394=>"010111011",
  62395=>"000011001",
  62396=>"010011011",
  62397=>"001000010",
  62398=>"111100101",
  62399=>"111110100",
  62400=>"111010111",
  62401=>"110001110",
  62402=>"111110000",
  62403=>"000011000",
  62404=>"110011110",
  62405=>"100101001",
  62406=>"000110000",
  62407=>"110001100",
  62408=>"101010101",
  62409=>"000101110",
  62410=>"100101001",
  62411=>"000000011",
  62412=>"101110000",
  62413=>"100110010",
  62414=>"100101011",
  62415=>"010000000",
  62416=>"011111111",
  62417=>"111011100",
  62418=>"111111100",
  62419=>"100100010",
  62420=>"000000011",
  62421=>"110001101",
  62422=>"000011111",
  62423=>"001010001",
  62424=>"000010101",
  62425=>"010000000",
  62426=>"110100100",
  62427=>"011010000",
  62428=>"110110001",
  62429=>"101011110",
  62430=>"111100111",
  62431=>"010011000",
  62432=>"100100101",
  62433=>"000010011",
  62434=>"000100001",
  62435=>"100000111",
  62436=>"000010000",
  62437=>"101001100",
  62438=>"100001001",
  62439=>"010101000",
  62440=>"111101110",
  62441=>"111111001",
  62442=>"000111000",
  62443=>"101001100",
  62444=>"011000100",
  62445=>"011010001",
  62446=>"010101001",
  62447=>"110101110",
  62448=>"011010111",
  62449=>"010101110",
  62450=>"111110110",
  62451=>"110111101",
  62452=>"000100000",
  62453=>"011001111",
  62454=>"100010110",
  62455=>"010101001",
  62456=>"011101100",
  62457=>"111010100",
  62458=>"010001010",
  62459=>"011101101",
  62460=>"101100001",
  62461=>"100110010",
  62462=>"101101100",
  62463=>"101010110",
  62464=>"101100100",
  62465=>"100011010",
  62466=>"111001010",
  62467=>"000010001",
  62468=>"000101000",
  62469=>"100101001",
  62470=>"111001110",
  62471=>"001111010",
  62472=>"110000000",
  62473=>"001000001",
  62474=>"000001010",
  62475=>"000011000",
  62476=>"111101101",
  62477=>"010101010",
  62478=>"011111111",
  62479=>"101110001",
  62480=>"010000100",
  62481=>"011010000",
  62482=>"001011010",
  62483=>"001101001",
  62484=>"011000011",
  62485=>"110100000",
  62486=>"000110011",
  62487=>"110100010",
  62488=>"110100110",
  62489=>"111100111",
  62490=>"010010000",
  62491=>"111000111",
  62492=>"110100000",
  62493=>"000100011",
  62494=>"001010010",
  62495=>"000100000",
  62496=>"001111100",
  62497=>"010001010",
  62498=>"010100101",
  62499=>"001101010",
  62500=>"110101111",
  62501=>"011110100",
  62502=>"000100010",
  62503=>"001001001",
  62504=>"100111111",
  62505=>"000010110",
  62506=>"000111011",
  62507=>"111111111",
  62508=>"100101111",
  62509=>"100011100",
  62510=>"000000101",
  62511=>"001111110",
  62512=>"101000000",
  62513=>"010001100",
  62514=>"100110000",
  62515=>"001011101",
  62516=>"010010000",
  62517=>"011000011",
  62518=>"101101001",
  62519=>"001100000",
  62520=>"000100000",
  62521=>"110000010",
  62522=>"010010010",
  62523=>"111000011",
  62524=>"000100101",
  62525=>"100000000",
  62526=>"100000000",
  62527=>"010011100",
  62528=>"010010101",
  62529=>"000100010",
  62530=>"001011011",
  62531=>"010010111",
  62532=>"010000101",
  62533=>"001101110",
  62534=>"000011001",
  62535=>"010001001",
  62536=>"100001010",
  62537=>"011011010",
  62538=>"000000100",
  62539=>"101001110",
  62540=>"010001000",
  62541=>"111011101",
  62542=>"101001001",
  62543=>"101101111",
  62544=>"001000000",
  62545=>"101101101",
  62546=>"110010111",
  62547=>"000101101",
  62548=>"000000110",
  62549=>"111101110",
  62550=>"100010000",
  62551=>"101101010",
  62552=>"010101110",
  62553=>"011011000",
  62554=>"001000111",
  62555=>"000000001",
  62556=>"010000011",
  62557=>"110101001",
  62558=>"101001010",
  62559=>"101011101",
  62560=>"001000000",
  62561=>"010000011",
  62562=>"000111000",
  62563=>"001001010",
  62564=>"000100101",
  62565=>"010100010",
  62566=>"010100101",
  62567=>"000000101",
  62568=>"000100001",
  62569=>"111111110",
  62570=>"010101000",
  62571=>"100011011",
  62572=>"110101101",
  62573=>"011101111",
  62574=>"100111010",
  62575=>"001101000",
  62576=>"110000010",
  62577=>"110110011",
  62578=>"111010011",
  62579=>"101101001",
  62580=>"011010100",
  62581=>"100101111",
  62582=>"000101101",
  62583=>"000111101",
  62584=>"111010100",
  62585=>"011110011",
  62586=>"101000101",
  62587=>"011110111",
  62588=>"000101100",
  62589=>"000110010",
  62590=>"001010110",
  62591=>"010011100",
  62592=>"100000011",
  62593=>"101010011",
  62594=>"110000111",
  62595=>"001001011",
  62596=>"101001010",
  62597=>"010011100",
  62598=>"111100001",
  62599=>"011001011",
  62600=>"110001011",
  62601=>"000011000",
  62602=>"110000110",
  62603=>"010000000",
  62604=>"010011000",
  62605=>"000000110",
  62606=>"100111111",
  62607=>"111100100",
  62608=>"101110010",
  62609=>"101100111",
  62610=>"110110101",
  62611=>"101010111",
  62612=>"110101111",
  62613=>"100000101",
  62614=>"011110111",
  62615=>"010100001",
  62616=>"110011101",
  62617=>"100001000",
  62618=>"010011001",
  62619=>"111111101",
  62620=>"111011000",
  62621=>"010100100",
  62622=>"000010001",
  62623=>"000111001",
  62624=>"010000010",
  62625=>"100010110",
  62626=>"001001011",
  62627=>"000111010",
  62628=>"001100000",
  62629=>"010110010",
  62630=>"010100110",
  62631=>"101100000",
  62632=>"011000111",
  62633=>"101001001",
  62634=>"101011111",
  62635=>"100111101",
  62636=>"111011000",
  62637=>"000101000",
  62638=>"000111111",
  62639=>"101111011",
  62640=>"111010000",
  62641=>"000000000",
  62642=>"010100010",
  62643=>"011110100",
  62644=>"010010100",
  62645=>"110000010",
  62646=>"110100100",
  62647=>"011110101",
  62648=>"100011111",
  62649=>"101100111",
  62650=>"000100000",
  62651=>"111011010",
  62652=>"101101110",
  62653=>"011101100",
  62654=>"111010010",
  62655=>"110111110",
  62656=>"000010010",
  62657=>"101001100",
  62658=>"100101101",
  62659=>"011110100",
  62660=>"111010111",
  62661=>"011111111",
  62662=>"110001011",
  62663=>"001110101",
  62664=>"100110001",
  62665=>"110110000",
  62666=>"101010000",
  62667=>"110111100",
  62668=>"001110110",
  62669=>"111101111",
  62670=>"011001010",
  62671=>"111101010",
  62672=>"000001111",
  62673=>"010010100",
  62674=>"010110101",
  62675=>"100011011",
  62676=>"101101001",
  62677=>"011111110",
  62678=>"010111000",
  62679=>"110111000",
  62680=>"100000010",
  62681=>"010110111",
  62682=>"010011100",
  62683=>"111101110",
  62684=>"100101011",
  62685=>"011100110",
  62686=>"011101010",
  62687=>"100000000",
  62688=>"010011000",
  62689=>"101001001",
  62690=>"101100110",
  62691=>"010110110",
  62692=>"111011100",
  62693=>"001011010",
  62694=>"001111101",
  62695=>"001110001",
  62696=>"011101001",
  62697=>"001110001",
  62698=>"111110110",
  62699=>"000011001",
  62700=>"110110100",
  62701=>"110111001",
  62702=>"000101110",
  62703=>"010111111",
  62704=>"101001011",
  62705=>"101110010",
  62706=>"100101111",
  62707=>"000000000",
  62708=>"010110111",
  62709=>"111000010",
  62710=>"011110101",
  62711=>"100001000",
  62712=>"111000000",
  62713=>"010100110",
  62714=>"111111111",
  62715=>"001010001",
  62716=>"010100011",
  62717=>"110111101",
  62718=>"011111001",
  62719=>"101111001",
  62720=>"001111000",
  62721=>"010111001",
  62722=>"010001000",
  62723=>"100111110",
  62724=>"110011011",
  62725=>"101110010",
  62726=>"010001100",
  62727=>"010010011",
  62728=>"010111110",
  62729=>"101001100",
  62730=>"001000110",
  62731=>"001001000",
  62732=>"101101100",
  62733=>"011001000",
  62734=>"000001001",
  62735=>"010111011",
  62736=>"001111101",
  62737=>"000000111",
  62738=>"110011010",
  62739=>"100001010",
  62740=>"010100100",
  62741=>"010100101",
  62742=>"110010100",
  62743=>"001011110",
  62744=>"000010001",
  62745=>"011100010",
  62746=>"100101000",
  62747=>"001001101",
  62748=>"100011011",
  62749=>"110111100",
  62750=>"101101010",
  62751=>"110111000",
  62752=>"101111100",
  62753=>"101111100",
  62754=>"110011111",
  62755=>"011111101",
  62756=>"101110111",
  62757=>"010101110",
  62758=>"000010100",
  62759=>"100010010",
  62760=>"001110000",
  62761=>"111010010",
  62762=>"010010110",
  62763=>"110000100",
  62764=>"011100111",
  62765=>"111011101",
  62766=>"110010010",
  62767=>"110011001",
  62768=>"010011001",
  62769=>"010000111",
  62770=>"001110011",
  62771=>"001011000",
  62772=>"000111000",
  62773=>"011110000",
  62774=>"111000000",
  62775=>"111000000",
  62776=>"000101100",
  62777=>"100101100",
  62778=>"000011100",
  62779=>"011000101",
  62780=>"010111111",
  62781=>"101110010",
  62782=>"110001111",
  62783=>"001011101",
  62784=>"000111100",
  62785=>"010000000",
  62786=>"111001010",
  62787=>"100010000",
  62788=>"001101101",
  62789=>"111001100",
  62790=>"000110101",
  62791=>"010111001",
  62792=>"010010100",
  62793=>"110100010",
  62794=>"001010010",
  62795=>"100100000",
  62796=>"010100101",
  62797=>"100111011",
  62798=>"100100010",
  62799=>"010100111",
  62800=>"011100101",
  62801=>"111101101",
  62802=>"001110001",
  62803=>"000001001",
  62804=>"101111111",
  62805=>"101110111",
  62806=>"111100011",
  62807=>"111111001",
  62808=>"000101110",
  62809=>"011000111",
  62810=>"101010000",
  62811=>"100101001",
  62812=>"111010101",
  62813=>"001001011",
  62814=>"010110001",
  62815=>"011001000",
  62816=>"111001000",
  62817=>"101101100",
  62818=>"001000100",
  62819=>"010111111",
  62820=>"111100111",
  62821=>"001111010",
  62822=>"111001101",
  62823=>"011011110",
  62824=>"000111000",
  62825=>"010011010",
  62826=>"110000001",
  62827=>"000100011",
  62828=>"100000011",
  62829=>"011000011",
  62830=>"011010010",
  62831=>"101100100",
  62832=>"100110011",
  62833=>"101100000",
  62834=>"111101100",
  62835=>"110011010",
  62836=>"000000111",
  62837=>"000011111",
  62838=>"010010110",
  62839=>"010000000",
  62840=>"110010001",
  62841=>"010100111",
  62842=>"010100100",
  62843=>"011100000",
  62844=>"100111000",
  62845=>"101000100",
  62846=>"101000111",
  62847=>"111100000",
  62848=>"001011110",
  62849=>"100110101",
  62850=>"101000101",
  62851=>"101101011",
  62852=>"101001101",
  62853=>"101101000",
  62854=>"000101110",
  62855=>"000100100",
  62856=>"010000000",
  62857=>"101000011",
  62858=>"001010010",
  62859=>"010100011",
  62860=>"001100000",
  62861=>"110010100",
  62862=>"010111010",
  62863=>"110010000",
  62864=>"011010010",
  62865=>"101110010",
  62866=>"110000000",
  62867=>"000110010",
  62868=>"000010110",
  62869=>"011010101",
  62870=>"111011111",
  62871=>"110011000",
  62872=>"100100001",
  62873=>"100100010",
  62874=>"110001001",
  62875=>"010000111",
  62876=>"101100110",
  62877=>"110101111",
  62878=>"100100110",
  62879=>"010000010",
  62880=>"110101010",
  62881=>"011010001",
  62882=>"011100110",
  62883=>"000010010",
  62884=>"000010001",
  62885=>"110000110",
  62886=>"101010010",
  62887=>"000000010",
  62888=>"111101111",
  62889=>"000101101",
  62890=>"100010001",
  62891=>"010110001",
  62892=>"011111101",
  62893=>"111011101",
  62894=>"001001111",
  62895=>"001100001",
  62896=>"110001001",
  62897=>"101000000",
  62898=>"000001100",
  62899=>"111000010",
  62900=>"001111100",
  62901=>"111000010",
  62902=>"000010011",
  62903=>"101001001",
  62904=>"100000011",
  62905=>"000000000",
  62906=>"000010001",
  62907=>"101000101",
  62908=>"110100110",
  62909=>"011101111",
  62910=>"111001111",
  62911=>"110011001",
  62912=>"111001011",
  62913=>"000101110",
  62914=>"000001010",
  62915=>"001000100",
  62916=>"000100001",
  62917=>"110011001",
  62918=>"011110010",
  62919=>"100010000",
  62920=>"110110100",
  62921=>"111110010",
  62922=>"010111000",
  62923=>"000110000",
  62924=>"100110000",
  62925=>"111011101",
  62926=>"001100001",
  62927=>"100100100",
  62928=>"010111111",
  62929=>"001000101",
  62930=>"000010001",
  62931=>"101111000",
  62932=>"111101000",
  62933=>"100111111",
  62934=>"100001011",
  62935=>"101101011",
  62936=>"000000010",
  62937=>"011000010",
  62938=>"110100110",
  62939=>"001100000",
  62940=>"110111110",
  62941=>"101111101",
  62942=>"111011111",
  62943=>"101011011",
  62944=>"000011001",
  62945=>"010011111",
  62946=>"111011111",
  62947=>"110000111",
  62948=>"100001101",
  62949=>"011101111",
  62950=>"011001010",
  62951=>"111111011",
  62952=>"101011010",
  62953=>"101100101",
  62954=>"011010000",
  62955=>"100010100",
  62956=>"001011100",
  62957=>"110000001",
  62958=>"000010000",
  62959=>"110110011",
  62960=>"011001100",
  62961=>"000111000",
  62962=>"101101000",
  62963=>"111000011",
  62964=>"101000010",
  62965=>"100011010",
  62966=>"111001101",
  62967=>"100101011",
  62968=>"111001111",
  62969=>"010100011",
  62970=>"101101101",
  62971=>"110001010",
  62972=>"010101010",
  62973=>"011010000",
  62974=>"101010001",
  62975=>"001001001",
  62976=>"110100111",
  62977=>"011101001",
  62978=>"111111010",
  62979=>"110001000",
  62980=>"101111000",
  62981=>"010100110",
  62982=>"111111010",
  62983=>"000010100",
  62984=>"001010010",
  62985=>"011111110",
  62986=>"001000010",
  62987=>"111010101",
  62988=>"011001111",
  62989=>"011011011",
  62990=>"111101111",
  62991=>"111111011",
  62992=>"010011110",
  62993=>"010010001",
  62994=>"111010100",
  62995=>"010101001",
  62996=>"010110111",
  62997=>"100110001",
  62998=>"100001001",
  62999=>"010101010",
  63000=>"001001101",
  63001=>"001001010",
  63002=>"001000011",
  63003=>"010101000",
  63004=>"100000011",
  63005=>"000000111",
  63006=>"001100011",
  63007=>"010110001",
  63008=>"100001110",
  63009=>"010001011",
  63010=>"100010011",
  63011=>"000010101",
  63012=>"101010111",
  63013=>"110101011",
  63014=>"011001001",
  63015=>"001010011",
  63016=>"011100010",
  63017=>"111001000",
  63018=>"011100101",
  63019=>"101100001",
  63020=>"000000000",
  63021=>"010111100",
  63022=>"100100011",
  63023=>"010001000",
  63024=>"100011000",
  63025=>"000010111",
  63026=>"010010000",
  63027=>"111010010",
  63028=>"000101111",
  63029=>"010111111",
  63030=>"100100111",
  63031=>"011000000",
  63032=>"000101101",
  63033=>"111010010",
  63034=>"001101101",
  63035=>"100001011",
  63036=>"010001101",
  63037=>"100110010",
  63038=>"011101010",
  63039=>"010101101",
  63040=>"110001000",
  63041=>"100001010",
  63042=>"000010001",
  63043=>"010001111",
  63044=>"010100011",
  63045=>"011000100",
  63046=>"011101101",
  63047=>"100000111",
  63048=>"010100001",
  63049=>"011001101",
  63050=>"101000110",
  63051=>"001111011",
  63052=>"110000110",
  63053=>"100011001",
  63054=>"000001001",
  63055=>"000011111",
  63056=>"110101111",
  63057=>"000011100",
  63058=>"100000010",
  63059=>"000111010",
  63060=>"101010100",
  63061=>"111100101",
  63062=>"010010010",
  63063=>"000100100",
  63064=>"001001111",
  63065=>"000011001",
  63066=>"010101000",
  63067=>"011010100",
  63068=>"000011010",
  63069=>"101001111",
  63070=>"110101011",
  63071=>"110100111",
  63072=>"101011001",
  63073=>"110100101",
  63074=>"110100110",
  63075=>"100101011",
  63076=>"111011110",
  63077=>"010101000",
  63078=>"010111001",
  63079=>"100000010",
  63080=>"100110001",
  63081=>"111101110",
  63082=>"011010011",
  63083=>"000111110",
  63084=>"100100010",
  63085=>"100001101",
  63086=>"111011000",
  63087=>"010010101",
  63088=>"000001001",
  63089=>"000011101",
  63090=>"010110011",
  63091=>"110011001",
  63092=>"110100100",
  63093=>"101000101",
  63094=>"001011011",
  63095=>"101001011",
  63096=>"111000110",
  63097=>"110001001",
  63098=>"110000111",
  63099=>"000000110",
  63100=>"000010000",
  63101=>"001101101",
  63102=>"001110101",
  63103=>"110010000",
  63104=>"010111101",
  63105=>"100110010",
  63106=>"010110111",
  63107=>"010000001",
  63108=>"000110010",
  63109=>"001001000",
  63110=>"101101100",
  63111=>"000111001",
  63112=>"110110011",
  63113=>"010000000",
  63114=>"000101010",
  63115=>"111110010",
  63116=>"010000000",
  63117=>"010100011",
  63118=>"111010101",
  63119=>"101011000",
  63120=>"111100011",
  63121=>"010011010",
  63122=>"011010010",
  63123=>"001000000",
  63124=>"000110100",
  63125=>"110011010",
  63126=>"100100110",
  63127=>"111011111",
  63128=>"011001000",
  63129=>"000110111",
  63130=>"110011111",
  63131=>"111010000",
  63132=>"011011101",
  63133=>"011110011",
  63134=>"111101011",
  63135=>"010011111",
  63136=>"111011111",
  63137=>"010111000",
  63138=>"011100110",
  63139=>"010001011",
  63140=>"000010101",
  63141=>"111000101",
  63142=>"000010101",
  63143=>"000101010",
  63144=>"011110001",
  63145=>"001100011",
  63146=>"011110001",
  63147=>"101000100",
  63148=>"100001001",
  63149=>"000011011",
  63150=>"111011111",
  63151=>"110110001",
  63152=>"011110011",
  63153=>"110101110",
  63154=>"110101111",
  63155=>"011010110",
  63156=>"010110101",
  63157=>"110111110",
  63158=>"111010010",
  63159=>"110111110",
  63160=>"100000110",
  63161=>"011110010",
  63162=>"100010110",
  63163=>"001100010",
  63164=>"000010011",
  63165=>"110110000",
  63166=>"011110010",
  63167=>"010101101",
  63168=>"110100001",
  63169=>"110011101",
  63170=>"100010110",
  63171=>"011101111",
  63172=>"100110110",
  63173=>"110010010",
  63174=>"100100111",
  63175=>"111101101",
  63176=>"011000011",
  63177=>"011001000",
  63178=>"010111101",
  63179=>"101000100",
  63180=>"100101011",
  63181=>"101001000",
  63182=>"010001000",
  63183=>"001101011",
  63184=>"000000011",
  63185=>"001000110",
  63186=>"010100000",
  63187=>"001011100",
  63188=>"011111000",
  63189=>"000110010",
  63190=>"001111101",
  63191=>"011101111",
  63192=>"000100000",
  63193=>"101010111",
  63194=>"000100100",
  63195=>"111100100",
  63196=>"111111111",
  63197=>"110000000",
  63198=>"100010001",
  63199=>"011111010",
  63200=>"001000110",
  63201=>"110110000",
  63202=>"001111110",
  63203=>"011000100",
  63204=>"011000101",
  63205=>"101000111",
  63206=>"000000010",
  63207=>"011000100",
  63208=>"000001001",
  63209=>"011010000",
  63210=>"100110110",
  63211=>"111111011",
  63212=>"000101001",
  63213=>"001010110",
  63214=>"000111001",
  63215=>"001100101",
  63216=>"110010001",
  63217=>"001101110",
  63218=>"100000100",
  63219=>"001111101",
  63220=>"101100001",
  63221=>"000101010",
  63222=>"000110000",
  63223=>"111001000",
  63224=>"010111001",
  63225=>"001010101",
  63226=>"101000010",
  63227=>"000000000",
  63228=>"110001000",
  63229=>"010010110",
  63230=>"000000000",
  63231=>"110111001",
  63232=>"010101101",
  63233=>"001111101",
  63234=>"010110101",
  63235=>"111100111",
  63236=>"001011100",
  63237=>"011000101",
  63238=>"111110110",
  63239=>"100010111",
  63240=>"000011110",
  63241=>"100110111",
  63242=>"011110100",
  63243=>"001010011",
  63244=>"011000100",
  63245=>"110100000",
  63246=>"100101100",
  63247=>"010111100",
  63248=>"111100001",
  63249=>"000001000",
  63250=>"110010110",
  63251=>"010101000",
  63252=>"000001100",
  63253=>"110110011",
  63254=>"100110000",
  63255=>"110101001",
  63256=>"000111110",
  63257=>"100111010",
  63258=>"010011111",
  63259=>"010101110",
  63260=>"001010100",
  63261=>"101011010",
  63262=>"010101011",
  63263=>"000011000",
  63264=>"000110101",
  63265=>"001000111",
  63266=>"010000100",
  63267=>"000101011",
  63268=>"001001111",
  63269=>"010101001",
  63270=>"100100010",
  63271=>"001101100",
  63272=>"000101111",
  63273=>"111000001",
  63274=>"011111111",
  63275=>"001010000",
  63276=>"100110101",
  63277=>"110110100",
  63278=>"001111010",
  63279=>"011111010",
  63280=>"001000010",
  63281=>"110101100",
  63282=>"111101010",
  63283=>"110000000",
  63284=>"110110100",
  63285=>"000100000",
  63286=>"100001110",
  63287=>"100111101",
  63288=>"100011101",
  63289=>"111100111",
  63290=>"101111000",
  63291=>"111100011",
  63292=>"100010001",
  63293=>"100000111",
  63294=>"001001010",
  63295=>"001010001",
  63296=>"111001100",
  63297=>"011100010",
  63298=>"011000011",
  63299=>"111001101",
  63300=>"100101101",
  63301=>"100111100",
  63302=>"101101110",
  63303=>"111001111",
  63304=>"010001000",
  63305=>"110110111",
  63306=>"001010100",
  63307=>"000001000",
  63308=>"000010110",
  63309=>"001001110",
  63310=>"101011100",
  63311=>"010111000",
  63312=>"110110110",
  63313=>"000101101",
  63314=>"000111111",
  63315=>"111000110",
  63316=>"111101101",
  63317=>"010000100",
  63318=>"100000011",
  63319=>"000100111",
  63320=>"111011101",
  63321=>"010001111",
  63322=>"011101001",
  63323=>"001000111",
  63324=>"011110101",
  63325=>"111100011",
  63326=>"101110111",
  63327=>"100001001",
  63328=>"001011101",
  63329=>"001000000",
  63330=>"000110000",
  63331=>"010101101",
  63332=>"010001000",
  63333=>"000100011",
  63334=>"101101011",
  63335=>"011111100",
  63336=>"000101100",
  63337=>"100000100",
  63338=>"000001001",
  63339=>"001010101",
  63340=>"111100011",
  63341=>"001111110",
  63342=>"100000110",
  63343=>"011101100",
  63344=>"100110000",
  63345=>"001010100",
  63346=>"101100000",
  63347=>"000001000",
  63348=>"010101100",
  63349=>"101011111",
  63350=>"110101111",
  63351=>"010000100",
  63352=>"111011010",
  63353=>"010000010",
  63354=>"111010000",
  63355=>"001101110",
  63356=>"100001010",
  63357=>"000111101",
  63358=>"011101001",
  63359=>"010010011",
  63360=>"001111100",
  63361=>"100001010",
  63362=>"010100101",
  63363=>"011101000",
  63364=>"001111101",
  63365=>"100111100",
  63366=>"111110010",
  63367=>"000101011",
  63368=>"111101111",
  63369=>"111111101",
  63370=>"100111010",
  63371=>"100101011",
  63372=>"001000001",
  63373=>"111111011",
  63374=>"010010011",
  63375=>"001000100",
  63376=>"000111100",
  63377=>"001111000",
  63378=>"100000101",
  63379=>"001100000",
  63380=>"110001001",
  63381=>"110011000",
  63382=>"010010011",
  63383=>"001001100",
  63384=>"101100111",
  63385=>"101111101",
  63386=>"000011001",
  63387=>"110011101",
  63388=>"111001010",
  63389=>"010100001",
  63390=>"101101100",
  63391=>"001100001",
  63392=>"100000000",
  63393=>"110111101",
  63394=>"001111001",
  63395=>"100101000",
  63396=>"000001111",
  63397=>"001011000",
  63398=>"010111000",
  63399=>"000000100",
  63400=>"110000101",
  63401=>"000011000",
  63402=>"001011110",
  63403=>"001101111",
  63404=>"001010001",
  63405=>"000101011",
  63406=>"000001000",
  63407=>"101110011",
  63408=>"110111100",
  63409=>"111011100",
  63410=>"000100011",
  63411=>"100111111",
  63412=>"010001101",
  63413=>"000011101",
  63414=>"011101101",
  63415=>"110011101",
  63416=>"101011111",
  63417=>"100011000",
  63418=>"110001111",
  63419=>"000110011",
  63420=>"001100011",
  63421=>"110111100",
  63422=>"111000000",
  63423=>"110011010",
  63424=>"110110000",
  63425=>"010000010",
  63426=>"111000101",
  63427=>"101001100",
  63428=>"001010101",
  63429=>"001110001",
  63430=>"010010001",
  63431=>"101000110",
  63432=>"011111101",
  63433=>"011111000",
  63434=>"000000000",
  63435=>"110011110",
  63436=>"111011011",
  63437=>"111110110",
  63438=>"010110110",
  63439=>"001010100",
  63440=>"101000011",
  63441=>"010111000",
  63442=>"110111101",
  63443=>"001000100",
  63444=>"001001101",
  63445=>"111001010",
  63446=>"101110000",
  63447=>"010100011",
  63448=>"001110000",
  63449=>"010011100",
  63450=>"000011100",
  63451=>"010000111",
  63452=>"010100101",
  63453=>"100000100",
  63454=>"000111111",
  63455=>"110010100",
  63456=>"001011000",
  63457=>"001100100",
  63458=>"111101111",
  63459=>"000110010",
  63460=>"101001001",
  63461=>"111100110",
  63462=>"010101101",
  63463=>"010100111",
  63464=>"101011110",
  63465=>"100010100",
  63466=>"000110000",
  63467=>"100110000",
  63468=>"111110110",
  63469=>"110000101",
  63470=>"100110000",
  63471=>"100110110",
  63472=>"110010011",
  63473=>"111101111",
  63474=>"010110110",
  63475=>"000111001",
  63476=>"001010111",
  63477=>"100101111",
  63478=>"010011000",
  63479=>"011010101",
  63480=>"010101010",
  63481=>"000010100",
  63482=>"011100000",
  63483=>"010011010",
  63484=>"110101111",
  63485=>"100011110",
  63486=>"110100010",
  63487=>"011001000",
  63488=>"010010111",
  63489=>"110111101",
  63490=>"010010000",
  63491=>"101101010",
  63492=>"110000111",
  63493=>"110011110",
  63494=>"110011111",
  63495=>"011100110",
  63496=>"000111111",
  63497=>"111100110",
  63498=>"001010011",
  63499=>"000101101",
  63500=>"100000100",
  63501=>"001011101",
  63502=>"000011100",
  63503=>"010111011",
  63504=>"001001010",
  63505=>"000111010",
  63506=>"101111010",
  63507=>"011010000",
  63508=>"100011111",
  63509=>"110011000",
  63510=>"111100100",
  63511=>"111000011",
  63512=>"011100001",
  63513=>"110001100",
  63514=>"100111000",
  63515=>"101011001",
  63516=>"000011110",
  63517=>"111101001",
  63518=>"111001010",
  63519=>"110001111",
  63520=>"001110000",
  63521=>"011111011",
  63522=>"010110000",
  63523=>"111000101",
  63524=>"010011111",
  63525=>"100000101",
  63526=>"100011000",
  63527=>"011010010",
  63528=>"011111000",
  63529=>"010010110",
  63530=>"100100101",
  63531=>"110100110",
  63532=>"100101011",
  63533=>"111111111",
  63534=>"010001101",
  63535=>"101111010",
  63536=>"010111011",
  63537=>"100011010",
  63538=>"000000100",
  63539=>"001110000",
  63540=>"101000110",
  63541=>"000000101",
  63542=>"011100011",
  63543=>"100001011",
  63544=>"100010001",
  63545=>"001001000",
  63546=>"011000011",
  63547=>"100000100",
  63548=>"100010101",
  63549=>"101110111",
  63550=>"111001011",
  63551=>"000010110",
  63552=>"010101101",
  63553=>"000000101",
  63554=>"100110100",
  63555=>"101001000",
  63556=>"110101001",
  63557=>"010010110",
  63558=>"101001001",
  63559=>"111101000",
  63560=>"000010011",
  63561=>"101000100",
  63562=>"111010001",
  63563=>"011000101",
  63564=>"111110001",
  63565=>"000111000",
  63566=>"111000010",
  63567=>"001001011",
  63568=>"001000001",
  63569=>"000101110",
  63570=>"111001010",
  63571=>"011101100",
  63572=>"111101110",
  63573=>"111101111",
  63574=>"001001000",
  63575=>"000110010",
  63576=>"010001100",
  63577=>"111010010",
  63578=>"000111001",
  63579=>"010011010",
  63580=>"011001111",
  63581=>"101101110",
  63582=>"101010110",
  63583=>"010111100",
  63584=>"001000000",
  63585=>"100010001",
  63586=>"010000000",
  63587=>"010010000",
  63588=>"001100101",
  63589=>"110111001",
  63590=>"010111101",
  63591=>"001110111",
  63592=>"111110100",
  63593=>"000011001",
  63594=>"101100000",
  63595=>"100010001",
  63596=>"011100001",
  63597=>"101100100",
  63598=>"111000110",
  63599=>"110100010",
  63600=>"010111100",
  63601=>"100000011",
  63602=>"010010010",
  63603=>"000101011",
  63604=>"000000110",
  63605=>"110010111",
  63606=>"111100111",
  63607=>"100101110",
  63608=>"010111001",
  63609=>"111100100",
  63610=>"100100011",
  63611=>"010000001",
  63612=>"001110110",
  63613=>"100111000",
  63614=>"011011100",
  63615=>"110111010",
  63616=>"100100000",
  63617=>"101111110",
  63618=>"101110111",
  63619=>"011000000",
  63620=>"010111111",
  63621=>"100000110",
  63622=>"111110101",
  63623=>"100111001",
  63624=>"010111101",
  63625=>"001111011",
  63626=>"000001101",
  63627=>"100010001",
  63628=>"101101001",
  63629=>"101110100",
  63630=>"101010101",
  63631=>"110011000",
  63632=>"010010110",
  63633=>"000000110",
  63634=>"101111001",
  63635=>"101110110",
  63636=>"000011100",
  63637=>"001100001",
  63638=>"001010001",
  63639=>"101110010",
  63640=>"010011001",
  63641=>"011010001",
  63642=>"010001110",
  63643=>"000001111",
  63644=>"110100101",
  63645=>"100011101",
  63646=>"011001000",
  63647=>"000110000",
  63648=>"000100001",
  63649=>"111101101",
  63650=>"000110001",
  63651=>"101101111",
  63652=>"111011011",
  63653=>"000011010",
  63654=>"011000000",
  63655=>"101111000",
  63656=>"011000100",
  63657=>"001111110",
  63658=>"001001101",
  63659=>"010101100",
  63660=>"110000100",
  63661=>"010110000",
  63662=>"001111101",
  63663=>"110110011",
  63664=>"001100110",
  63665=>"011111010",
  63666=>"101100000",
  63667=>"001010101",
  63668=>"000001010",
  63669=>"100000011",
  63670=>"001010001",
  63671=>"110000111",
  63672=>"011011010",
  63673=>"101000011",
  63674=>"011001011",
  63675=>"111101110",
  63676=>"010001010",
  63677=>"101100101",
  63678=>"111010011",
  63679=>"100011000",
  63680=>"110100100",
  63681=>"011001110",
  63682=>"010110110",
  63683=>"100100101",
  63684=>"011111001",
  63685=>"010000111",
  63686=>"111111001",
  63687=>"000011101",
  63688=>"001001101",
  63689=>"011011100",
  63690=>"111100101",
  63691=>"001010111",
  63692=>"011010100",
  63693=>"011000111",
  63694=>"001010011",
  63695=>"100110001",
  63696=>"111111100",
  63697=>"101000001",
  63698=>"111011100",
  63699=>"010110110",
  63700=>"000001011",
  63701=>"010001011",
  63702=>"111001011",
  63703=>"100111001",
  63704=>"100110111",
  63705=>"101011010",
  63706=>"000111111",
  63707=>"111010001",
  63708=>"101111000",
  63709=>"010110000",
  63710=>"001110101",
  63711=>"110011100",
  63712=>"000011100",
  63713=>"011011110",
  63714=>"110100111",
  63715=>"110110011",
  63716=>"010010111",
  63717=>"000101010",
  63718=>"010001010",
  63719=>"010011100",
  63720=>"100011001",
  63721=>"011111101",
  63722=>"000100111",
  63723=>"101111111",
  63724=>"100101001",
  63725=>"101100110",
  63726=>"010110011",
  63727=>"101001001",
  63728=>"011101101",
  63729=>"100010000",
  63730=>"100111011",
  63731=>"000001101",
  63732=>"010110000",
  63733=>"000100010",
  63734=>"010100000",
  63735=>"000100000",
  63736=>"100011011",
  63737=>"101011011",
  63738=>"011110011",
  63739=>"010000110",
  63740=>"001011110",
  63741=>"001110010",
  63742=>"101001000",
  63743=>"111101001",
  63744=>"001111001",
  63745=>"110110101",
  63746=>"101111110",
  63747=>"011001010",
  63748=>"011100100",
  63749=>"100111100",
  63750=>"111001111",
  63751=>"010111000",
  63752=>"100110010",
  63753=>"111100001",
  63754=>"000111010",
  63755=>"100011110",
  63756=>"001010011",
  63757=>"100000100",
  63758=>"101000010",
  63759=>"100110011",
  63760=>"100111000",
  63761=>"111101100",
  63762=>"110001000",
  63763=>"010110000",
  63764=>"001010111",
  63765=>"100101000",
  63766=>"100001000",
  63767=>"111110001",
  63768=>"110001111",
  63769=>"111110001",
  63770=>"000101001",
  63771=>"001001100",
  63772=>"111011010",
  63773=>"110011001",
  63774=>"001111100",
  63775=>"110101111",
  63776=>"111001000",
  63777=>"110111111",
  63778=>"111101111",
  63779=>"001100101",
  63780=>"100101001",
  63781=>"010101011",
  63782=>"001010110",
  63783=>"010101100",
  63784=>"000000011",
  63785=>"111111110",
  63786=>"110111001",
  63787=>"001010110",
  63788=>"110111110",
  63789=>"000101100",
  63790=>"100010000",
  63791=>"011111110",
  63792=>"110001101",
  63793=>"001011000",
  63794=>"101111001",
  63795=>"100011101",
  63796=>"011011001",
  63797=>"101111111",
  63798=>"111011001",
  63799=>"011100110",
  63800=>"111010100",
  63801=>"011011100",
  63802=>"010010111",
  63803=>"010110111",
  63804=>"111100100",
  63805=>"011000000",
  63806=>"000001100",
  63807=>"011111111",
  63808=>"001011101",
  63809=>"000010001",
  63810=>"000001010",
  63811=>"101100101",
  63812=>"001001111",
  63813=>"101100110",
  63814=>"100100100",
  63815=>"111010001",
  63816=>"110111100",
  63817=>"100110110",
  63818=>"010101111",
  63819=>"111010010",
  63820=>"100110110",
  63821=>"010110101",
  63822=>"101010111",
  63823=>"000000110",
  63824=>"011101010",
  63825=>"011100001",
  63826=>"100111100",
  63827=>"010111110",
  63828=>"110011010",
  63829=>"001011100",
  63830=>"101100110",
  63831=>"101110000",
  63832=>"000000111",
  63833=>"100000111",
  63834=>"111000100",
  63835=>"011111100",
  63836=>"100111101",
  63837=>"011100011",
  63838=>"101000110",
  63839=>"100001010",
  63840=>"011010101",
  63841=>"011111010",
  63842=>"100001000",
  63843=>"011111010",
  63844=>"010011000",
  63845=>"011110111",
  63846=>"101100110",
  63847=>"110001011",
  63848=>"011111100",
  63849=>"000110000",
  63850=>"100001000",
  63851=>"001111100",
  63852=>"101001011",
  63853=>"100000000",
  63854=>"010011010",
  63855=>"111001111",
  63856=>"010011011",
  63857=>"010001101",
  63858=>"000010100",
  63859=>"110001111",
  63860=>"110000000",
  63861=>"100001111",
  63862=>"001011010",
  63863=>"001011011",
  63864=>"110111101",
  63865=>"000101110",
  63866=>"000001000",
  63867=>"101110110",
  63868=>"100000000",
  63869=>"111000001",
  63870=>"010101010",
  63871=>"110000001",
  63872=>"111111111",
  63873=>"000101000",
  63874=>"111011011",
  63875=>"000111111",
  63876=>"010011100",
  63877=>"010110011",
  63878=>"111010111",
  63879=>"111010101",
  63880=>"010000111",
  63881=>"010010101",
  63882=>"111100000",
  63883=>"000000110",
  63884=>"010111011",
  63885=>"000000110",
  63886=>"001011000",
  63887=>"101101100",
  63888=>"111000001",
  63889=>"001101011",
  63890=>"001111100",
  63891=>"011110011",
  63892=>"101000001",
  63893=>"011101110",
  63894=>"001111010",
  63895=>"100010100",
  63896=>"000101000",
  63897=>"101011000",
  63898=>"010001011",
  63899=>"111010111",
  63900=>"110011010",
  63901=>"010100011",
  63902=>"110001001",
  63903=>"110100111",
  63904=>"010100111",
  63905=>"010100010",
  63906=>"011101011",
  63907=>"001101001",
  63908=>"000100011",
  63909=>"000100100",
  63910=>"000000000",
  63911=>"100110000",
  63912=>"110000101",
  63913=>"111100001",
  63914=>"100101100",
  63915=>"011100111",
  63916=>"010000101",
  63917=>"011100101",
  63918=>"001100010",
  63919=>"111101000",
  63920=>"101001011",
  63921=>"100010100",
  63922=>"100000010",
  63923=>"000010000",
  63924=>"100011110",
  63925=>"110011010",
  63926=>"001100111",
  63927=>"110100010",
  63928=>"100001000",
  63929=>"010000010",
  63930=>"001010011",
  63931=>"111100110",
  63932=>"111110100",
  63933=>"000001011",
  63934=>"100111110",
  63935=>"111100000",
  63936=>"010110100",
  63937=>"101000001",
  63938=>"011001101",
  63939=>"011011001",
  63940=>"010001010",
  63941=>"000001100",
  63942=>"001000010",
  63943=>"001100101",
  63944=>"010010100",
  63945=>"100000110",
  63946=>"101000001",
  63947=>"100011101",
  63948=>"001110111",
  63949=>"010011011",
  63950=>"010000010",
  63951=>"010111100",
  63952=>"110001111",
  63953=>"010110011",
  63954=>"010011110",
  63955=>"010010110",
  63956=>"011111010",
  63957=>"011000000",
  63958=>"101101011",
  63959=>"001111101",
  63960=>"111100001",
  63961=>"111001110",
  63962=>"001001101",
  63963=>"011101011",
  63964=>"100101001",
  63965=>"101111100",
  63966=>"110010010",
  63967=>"110111111",
  63968=>"000000010",
  63969=>"100000001",
  63970=>"010100001",
  63971=>"111110110",
  63972=>"011010100",
  63973=>"101110111",
  63974=>"011011100",
  63975=>"100110000",
  63976=>"100100010",
  63977=>"010010000",
  63978=>"000001100",
  63979=>"111001000",
  63980=>"110001101",
  63981=>"101100000",
  63982=>"010010011",
  63983=>"010011011",
  63984=>"011000001",
  63985=>"111110000",
  63986=>"111011000",
  63987=>"010111101",
  63988=>"111111001",
  63989=>"100001001",
  63990=>"111011101",
  63991=>"011110101",
  63992=>"110011011",
  63993=>"010011000",
  63994=>"111001000",
  63995=>"111011110",
  63996=>"000110101",
  63997=>"101000011",
  63998=>"111001010",
  63999=>"100111001",
  64000=>"001100100",
  64001=>"001100001",
  64002=>"110101000",
  64003=>"101000000",
  64004=>"011110100",
  64005=>"000000000",
  64006=>"001011000",
  64007=>"000110100",
  64008=>"110110010",
  64009=>"011101011",
  64010=>"011011101",
  64011=>"101110000",
  64012=>"111101011",
  64013=>"100000011",
  64014=>"000000001",
  64015=>"110100110",
  64016=>"010010110",
  64017=>"110110111",
  64018=>"111001101",
  64019=>"111100101",
  64020=>"011011001",
  64021=>"111111001",
  64022=>"110011111",
  64023=>"010110101",
  64024=>"010110101",
  64025=>"011111110",
  64026=>"001000100",
  64027=>"111100110",
  64028=>"101110001",
  64029=>"110000101",
  64030=>"011111101",
  64031=>"001010101",
  64032=>"110101001",
  64033=>"110110001",
  64034=>"101101011",
  64035=>"000001000",
  64036=>"101111101",
  64037=>"111001000",
  64038=>"111010110",
  64039=>"011111010",
  64040=>"000011000",
  64041=>"111101101",
  64042=>"111010100",
  64043=>"011011101",
  64044=>"100000100",
  64045=>"100010111",
  64046=>"000111010",
  64047=>"011010100",
  64048=>"111111001",
  64049=>"000011000",
  64050=>"110011101",
  64051=>"101011011",
  64052=>"101001100",
  64053=>"111100000",
  64054=>"000100000",
  64055=>"000100111",
  64056=>"100000100",
  64057=>"101100010",
  64058=>"111010110",
  64059=>"110001110",
  64060=>"000000001",
  64061=>"010011111",
  64062=>"000110000",
  64063=>"011000000",
  64064=>"101000011",
  64065=>"000000001",
  64066=>"011010011",
  64067=>"100010111",
  64068=>"101100010",
  64069=>"111010001",
  64070=>"111001011",
  64071=>"100101001",
  64072=>"101111001",
  64073=>"000011110",
  64074=>"110001101",
  64075=>"000010010",
  64076=>"110000001",
  64077=>"001100111",
  64078=>"111001011",
  64079=>"111110000",
  64080=>"111011010",
  64081=>"111110101",
  64082=>"110110011",
  64083=>"011110001",
  64084=>"000010110",
  64085=>"101010000",
  64086=>"001010001",
  64087=>"000000010",
  64088=>"111000110",
  64089=>"001011101",
  64090=>"101110111",
  64091=>"011011010",
  64092=>"011100111",
  64093=>"100010110",
  64094=>"011111000",
  64095=>"010110100",
  64096=>"011011111",
  64097=>"010010111",
  64098=>"000110100",
  64099=>"110000111",
  64100=>"000000111",
  64101=>"111110101",
  64102=>"101001001",
  64103=>"111001100",
  64104=>"010000010",
  64105=>"001100100",
  64106=>"111000100",
  64107=>"111101111",
  64108=>"001100000",
  64109=>"101111011",
  64110=>"000101110",
  64111=>"010000010",
  64112=>"101011000",
  64113=>"110101101",
  64114=>"111010010",
  64115=>"110010010",
  64116=>"111011001",
  64117=>"011100000",
  64118=>"110011010",
  64119=>"110010111",
  64120=>"101001110",
  64121=>"000010111",
  64122=>"001110010",
  64123=>"011101100",
  64124=>"010010111",
  64125=>"011001101",
  64126=>"001010001",
  64127=>"111001011",
  64128=>"001001000",
  64129=>"000101100",
  64130=>"111111111",
  64131=>"100011111",
  64132=>"001001100",
  64133=>"111101110",
  64134=>"011000010",
  64135=>"101001000",
  64136=>"001010110",
  64137=>"100011111",
  64138=>"000111101",
  64139=>"110010110",
  64140=>"111010011",
  64141=>"001001101",
  64142=>"010010010",
  64143=>"010101011",
  64144=>"010011100",
  64145=>"100110110",
  64146=>"010001010",
  64147=>"000111011",
  64148=>"011010001",
  64149=>"101100011",
  64150=>"111101000",
  64151=>"000010001",
  64152=>"000010111",
  64153=>"010010100",
  64154=>"011100101",
  64155=>"100110110",
  64156=>"011111110",
  64157=>"001011100",
  64158=>"001111100",
  64159=>"000101101",
  64160=>"001001011",
  64161=>"001010001",
  64162=>"000101000",
  64163=>"100110100",
  64164=>"101110011",
  64165=>"000001101",
  64166=>"100101010",
  64167=>"000010001",
  64168=>"110100001",
  64169=>"100000011",
  64170=>"000010111",
  64171=>"101010101",
  64172=>"100001001",
  64173=>"111001100",
  64174=>"110110010",
  64175=>"100111111",
  64176=>"001101001",
  64177=>"000100111",
  64178=>"001001110",
  64179=>"010010110",
  64180=>"101100100",
  64181=>"111100010",
  64182=>"101010011",
  64183=>"111001110",
  64184=>"010010001",
  64185=>"000001010",
  64186=>"010000100",
  64187=>"100001110",
  64188=>"011100000",
  64189=>"010111000",
  64190=>"001010100",
  64191=>"011101001",
  64192=>"000111110",
  64193=>"010111001",
  64194=>"101111101",
  64195=>"111010010",
  64196=>"101010110",
  64197=>"001111010",
  64198=>"110011000",
  64199=>"000000110",
  64200=>"000100101",
  64201=>"001100000",
  64202=>"100011001",
  64203=>"100010001",
  64204=>"111100000",
  64205=>"101000011",
  64206=>"101111100",
  64207=>"010000001",
  64208=>"011100010",
  64209=>"011011101",
  64210=>"101001110",
  64211=>"010000110",
  64212=>"110101100",
  64213=>"001001100",
  64214=>"001001001",
  64215=>"000100100",
  64216=>"111001100",
  64217=>"000010001",
  64218=>"110010110",
  64219=>"010000000",
  64220=>"010101100",
  64221=>"000011001",
  64222=>"000100010",
  64223=>"111101011",
  64224=>"001110010",
  64225=>"011101001",
  64226=>"011100011",
  64227=>"000110101",
  64228=>"011010101",
  64229=>"110011110",
  64230=>"000100101",
  64231=>"100101000",
  64232=>"001011011",
  64233=>"110110101",
  64234=>"010000000",
  64235=>"001111111",
  64236=>"001110101",
  64237=>"110101100",
  64238=>"110001100",
  64239=>"101010100",
  64240=>"010010001",
  64241=>"100001100",
  64242=>"010001011",
  64243=>"011101001",
  64244=>"100101111",
  64245=>"101101010",
  64246=>"100001001",
  64247=>"010000111",
  64248=>"110101010",
  64249=>"101110111",
  64250=>"101000111",
  64251=>"001000111",
  64252=>"011011001",
  64253=>"000110111",
  64254=>"001011111",
  64255=>"000100011",
  64256=>"100101100",
  64257=>"000000100",
  64258=>"001000101",
  64259=>"100100011",
  64260=>"110010011",
  64261=>"000110101",
  64262=>"000010100",
  64263=>"010000100",
  64264=>"001110000",
  64265=>"011100111",
  64266=>"100011100",
  64267=>"111101111",
  64268=>"000101101",
  64269=>"011101001",
  64270=>"001011111",
  64271=>"111111101",
  64272=>"000001110",
  64273=>"010011010",
  64274=>"100001110",
  64275=>"001001010",
  64276=>"001110000",
  64277=>"001000000",
  64278=>"100110101",
  64279=>"010101000",
  64280=>"111100100",
  64281=>"111001000",
  64282=>"011010010",
  64283=>"111000001",
  64284=>"000100001",
  64285=>"111000000",
  64286=>"011101110",
  64287=>"001111101",
  64288=>"000101011",
  64289=>"111001011",
  64290=>"111010101",
  64291=>"101100101",
  64292=>"111011001",
  64293=>"001000101",
  64294=>"000100111",
  64295=>"011110000",
  64296=>"110110111",
  64297=>"110110101",
  64298=>"001101000",
  64299=>"111101100",
  64300=>"010110001",
  64301=>"000001011",
  64302=>"100010011",
  64303=>"110111011",
  64304=>"001100000",
  64305=>"000001000",
  64306=>"100101111",
  64307=>"111011110",
  64308=>"000011111",
  64309=>"010111001",
  64310=>"111111011",
  64311=>"111011111",
  64312=>"010001001",
  64313=>"000000110",
  64314=>"001100111",
  64315=>"101011011",
  64316=>"000111001",
  64317=>"101101100",
  64318=>"001111111",
  64319=>"110111101",
  64320=>"000001101",
  64321=>"100100000",
  64322=>"111100000",
  64323=>"111100000",
  64324=>"111111010",
  64325=>"000000001",
  64326=>"011111001",
  64327=>"011111100",
  64328=>"100110001",
  64329=>"101011100",
  64330=>"001011100",
  64331=>"100000011",
  64332=>"011100101",
  64333=>"101110110",
  64334=>"111110111",
  64335=>"000010111",
  64336=>"001100100",
  64337=>"010101101",
  64338=>"110001000",
  64339=>"101000010",
  64340=>"111011110",
  64341=>"000010000",
  64342=>"010011011",
  64343=>"101011101",
  64344=>"010000100",
  64345=>"110110001",
  64346=>"001111101",
  64347=>"011000000",
  64348=>"111100000",
  64349=>"010011101",
  64350=>"111001111",
  64351=>"010100111",
  64352=>"001001000",
  64353=>"001110011",
  64354=>"001111011",
  64355=>"001101100",
  64356=>"011011011",
  64357=>"100000001",
  64358=>"110111101",
  64359=>"110101101",
  64360=>"010001010",
  64361=>"011000101",
  64362=>"010111000",
  64363=>"101110110",
  64364=>"000111100",
  64365=>"111100100",
  64366=>"101101011",
  64367=>"001110101",
  64368=>"101011111",
  64369=>"001011111",
  64370=>"111100011",
  64371=>"010001001",
  64372=>"100101100",
  64373=>"001101111",
  64374=>"101100011",
  64375=>"011110111",
  64376=>"001100110",
  64377=>"000001010",
  64378=>"101001100",
  64379=>"010101101",
  64380=>"001111101",
  64381=>"001010000",
  64382=>"100010001",
  64383=>"000010101",
  64384=>"001101011",
  64385=>"100110001",
  64386=>"010011010",
  64387=>"111001110",
  64388=>"110110101",
  64389=>"000011010",
  64390=>"101110110",
  64391=>"011011000",
  64392=>"100010010",
  64393=>"000110011",
  64394=>"001010101",
  64395=>"010101110",
  64396=>"001000011",
  64397=>"101000101",
  64398=>"010011010",
  64399=>"001001010",
  64400=>"010001011",
  64401=>"110011011",
  64402=>"000000011",
  64403=>"010100101",
  64404=>"000111011",
  64405=>"100011110",
  64406=>"101101111",
  64407=>"011110011",
  64408=>"111010101",
  64409=>"010011010",
  64410=>"100001000",
  64411=>"100100111",
  64412=>"101111000",
  64413=>"001100111",
  64414=>"001000101",
  64415=>"110000000",
  64416=>"010111000",
  64417=>"110000011",
  64418=>"101101010",
  64419=>"110111001",
  64420=>"101000001",
  64421=>"100101010",
  64422=>"111100000",
  64423=>"100001000",
  64424=>"100001111",
  64425=>"101101110",
  64426=>"000011101",
  64427=>"111100010",
  64428=>"010000001",
  64429=>"000001111",
  64430=>"001110100",
  64431=>"110011010",
  64432=>"010100011",
  64433=>"100010110",
  64434=>"111010010",
  64435=>"001011101",
  64436=>"010101000",
  64437=>"101101111",
  64438=>"110101101",
  64439=>"110011110",
  64440=>"011000000",
  64441=>"010100010",
  64442=>"111111101",
  64443=>"010011100",
  64444=>"010011001",
  64445=>"111110000",
  64446=>"110001000",
  64447=>"001001111",
  64448=>"110101111",
  64449=>"000000110",
  64450=>"011110100",
  64451=>"011101110",
  64452=>"110101010",
  64453=>"101010100",
  64454=>"001100001",
  64455=>"110000101",
  64456=>"000000001",
  64457=>"000000111",
  64458=>"111111110",
  64459=>"000111001",
  64460=>"001010100",
  64461=>"011110100",
  64462=>"001000100",
  64463=>"010101100",
  64464=>"111011110",
  64465=>"001010001",
  64466=>"111110110",
  64467=>"111011111",
  64468=>"010111000",
  64469=>"100000010",
  64470=>"111001000",
  64471=>"110001111",
  64472=>"001110000",
  64473=>"001100111",
  64474=>"111111111",
  64475=>"011111010",
  64476=>"011110100",
  64477=>"011100111",
  64478=>"001010100",
  64479=>"011101110",
  64480=>"101100100",
  64481=>"000011000",
  64482=>"011100101",
  64483=>"110011111",
  64484=>"101000000",
  64485=>"010100111",
  64486=>"011101000",
  64487=>"111010000",
  64488=>"001000111",
  64489=>"111010011",
  64490=>"010110000",
  64491=>"010101110",
  64492=>"001001111",
  64493=>"010100011",
  64494=>"100111101",
  64495=>"100111111",
  64496=>"100100000",
  64497=>"011100011",
  64498=>"110010110",
  64499=>"010100001",
  64500=>"100101101",
  64501=>"101001100",
  64502=>"000011110",
  64503=>"010101001",
  64504=>"110101111",
  64505=>"010111110",
  64506=>"101101001",
  64507=>"100100101",
  64508=>"011000110",
  64509=>"011111011",
  64510=>"110100010",
  64511=>"111100101",
  64512=>"110000100",
  64513=>"111100101",
  64514=>"011010000",
  64515=>"010111001",
  64516=>"001110011",
  64517=>"000001101",
  64518=>"101001101",
  64519=>"011001111",
  64520=>"010001000",
  64521=>"000000001",
  64522=>"000001001",
  64523=>"100111110",
  64524=>"111110000",
  64525=>"101011011",
  64526=>"100000001",
  64527=>"111100000",
  64528=>"101111100",
  64529=>"000000000",
  64530=>"111100001",
  64531=>"110101000",
  64532=>"010101101",
  64533=>"011011010",
  64534=>"100110111",
  64535=>"011000110",
  64536=>"111011000",
  64537=>"100010001",
  64538=>"100110101",
  64539=>"110001011",
  64540=>"111001001",
  64541=>"110001100",
  64542=>"110010111",
  64543=>"100011101",
  64544=>"110001110",
  64545=>"111111010",
  64546=>"000000000",
  64547=>"101110101",
  64548=>"101010010",
  64549=>"000111111",
  64550=>"011110001",
  64551=>"000001101",
  64552=>"110011100",
  64553=>"000001001",
  64554=>"000010001",
  64555=>"010111001",
  64556=>"101000001",
  64557=>"001100111",
  64558=>"011011010",
  64559=>"010100110",
  64560=>"110110011",
  64561=>"010000101",
  64562=>"111010001",
  64563=>"010110100",
  64564=>"000001001",
  64565=>"000011110",
  64566=>"001111011",
  64567=>"101111011",
  64568=>"100110000",
  64569=>"110000000",
  64570=>"100001000",
  64571=>"000000010",
  64572=>"000000110",
  64573=>"010011101",
  64574=>"011101000",
  64575=>"101110100",
  64576=>"001010100",
  64577=>"000010100",
  64578=>"100100111",
  64579=>"111010100",
  64580=>"011001000",
  64581=>"001001111",
  64582=>"111110110",
  64583=>"000000001",
  64584=>"110000100",
  64585=>"100110010",
  64586=>"100000001",
  64587=>"101010001",
  64588=>"110010000",
  64589=>"111000011",
  64590=>"101011001",
  64591=>"111001110",
  64592=>"101110111",
  64593=>"111011010",
  64594=>"101100101",
  64595=>"100011100",
  64596=>"011011110",
  64597=>"000110110",
  64598=>"011000101",
  64599=>"000110011",
  64600=>"011101101",
  64601=>"000101101",
  64602=>"010011100",
  64603=>"110011100",
  64604=>"000100001",
  64605=>"010111011",
  64606=>"100111101",
  64607=>"110000101",
  64608=>"111010010",
  64609=>"011110001",
  64610=>"111101110",
  64611=>"101011001",
  64612=>"010111110",
  64613=>"111010001",
  64614=>"010011101",
  64615=>"101010000",
  64616=>"011111101",
  64617=>"011100010",
  64618=>"010100111",
  64619=>"000000001",
  64620=>"110000110",
  64621=>"001000111",
  64622=>"000110111",
  64623=>"011111001",
  64624=>"001101100",
  64625=>"011110111",
  64626=>"011111110",
  64627=>"110101110",
  64628=>"010011000",
  64629=>"101100111",
  64630=>"111110100",
  64631=>"010001110",
  64632=>"101111111",
  64633=>"101100010",
  64634=>"010010001",
  64635=>"011101010",
  64636=>"101000100",
  64637=>"000010111",
  64638=>"000111000",
  64639=>"101010001",
  64640=>"111100010",
  64641=>"001001011",
  64642=>"001000110",
  64643=>"000110100",
  64644=>"001011110",
  64645=>"111010100",
  64646=>"000000001",
  64647=>"011100001",
  64648=>"001001000",
  64649=>"001001011",
  64650=>"010100110",
  64651=>"000001110",
  64652=>"010100001",
  64653=>"110111110",
  64654=>"110111000",
  64655=>"111101010",
  64656=>"001010000",
  64657=>"000010001",
  64658=>"110111110",
  64659=>"001110011",
  64660=>"110001000",
  64661=>"010111010",
  64662=>"010111010",
  64663=>"001011111",
  64664=>"000111101",
  64665=>"110001011",
  64666=>"100100110",
  64667=>"000010000",
  64668=>"001011100",
  64669=>"100011110",
  64670=>"001000001",
  64671=>"000011101",
  64672=>"101110000",
  64673=>"001001100",
  64674=>"000101000",
  64675=>"101110100",
  64676=>"111111011",
  64677=>"011110110",
  64678=>"000000110",
  64679=>"100111011",
  64680=>"110110110",
  64681=>"100100000",
  64682=>"010011111",
  64683=>"110001101",
  64684=>"111001000",
  64685=>"100011101",
  64686=>"110011011",
  64687=>"000101000",
  64688=>"010010101",
  64689=>"010000001",
  64690=>"111111111",
  64691=>"100100111",
  64692=>"000101000",
  64693=>"111111101",
  64694=>"000000111",
  64695=>"011010010",
  64696=>"000001000",
  64697=>"011101111",
  64698=>"001001001",
  64699=>"000010100",
  64700=>"111010100",
  64701=>"001000011",
  64702=>"011100100",
  64703=>"000101000",
  64704=>"111011000",
  64705=>"010011001",
  64706=>"000101100",
  64707=>"110100011",
  64708=>"010011010",
  64709=>"000011100",
  64710=>"100101000",
  64711=>"010010000",
  64712=>"011001110",
  64713=>"001011101",
  64714=>"101010000",
  64715=>"011111001",
  64716=>"110000111",
  64717=>"100011011",
  64718=>"111101011",
  64719=>"011101101",
  64720=>"001000011",
  64721=>"111010001",
  64722=>"101000101",
  64723=>"100001001",
  64724=>"110100011",
  64725=>"011000111",
  64726=>"111100101",
  64727=>"000000111",
  64728=>"110000001",
  64729=>"001001010",
  64730=>"010011101",
  64731=>"100011000",
  64732=>"111111001",
  64733=>"101100100",
  64734=>"000110110",
  64735=>"100101011",
  64736=>"001110110",
  64737=>"110110110",
  64738=>"000011111",
  64739=>"101101101",
  64740=>"110001110",
  64741=>"111100110",
  64742=>"001000110",
  64743=>"010001010",
  64744=>"100011011",
  64745=>"100111111",
  64746=>"101111010",
  64747=>"001001011",
  64748=>"010101000",
  64749=>"111100100",
  64750=>"000000111",
  64751=>"110011110",
  64752=>"110111110",
  64753=>"001100101",
  64754=>"100001011",
  64755=>"000100010",
  64756=>"111011110",
  64757=>"001101111",
  64758=>"111000110",
  64759=>"010010000",
  64760=>"001000111",
  64761=>"111100000",
  64762=>"000101101",
  64763=>"011010010",
  64764=>"110001101",
  64765=>"001001010",
  64766=>"010010001",
  64767=>"011101110",
  64768=>"010110001",
  64769=>"111110011",
  64770=>"000101110",
  64771=>"001111100",
  64772=>"111100010",
  64773=>"110110111",
  64774=>"010100111",
  64775=>"001101010",
  64776=>"001011000",
  64777=>"000110100",
  64778=>"010010011",
  64779=>"101101101",
  64780=>"000110011",
  64781=>"110011011",
  64782=>"011011101",
  64783=>"101110101",
  64784=>"011010111",
  64785=>"011000100",
  64786=>"101111110",
  64787=>"100110001",
  64788=>"000111000",
  64789=>"111011101",
  64790=>"000001111",
  64791=>"111010000",
  64792=>"010010010",
  64793=>"001110000",
  64794=>"011000000",
  64795=>"001110000",
  64796=>"000101000",
  64797=>"011100011",
  64798=>"101110001",
  64799=>"111011010",
  64800=>"001110000",
  64801=>"010101000",
  64802=>"011101101",
  64803=>"100100011",
  64804=>"001000111",
  64805=>"011110110",
  64806=>"000001110",
  64807=>"110100011",
  64808=>"000000010",
  64809=>"001011100",
  64810=>"110100010",
  64811=>"101011101",
  64812=>"001000000",
  64813=>"101010111",
  64814=>"111001101",
  64815=>"111100111",
  64816=>"000101000",
  64817=>"100110000",
  64818=>"011011000",
  64819=>"011000001",
  64820=>"111010100",
  64821=>"110001001",
  64822=>"011011111",
  64823=>"000101111",
  64824=>"000011100",
  64825=>"101010010",
  64826=>"111110100",
  64827=>"111101111",
  64828=>"100111100",
  64829=>"101100001",
  64830=>"101100111",
  64831=>"100110110",
  64832=>"101110000",
  64833=>"001010110",
  64834=>"001100100",
  64835=>"011100000",
  64836=>"000111110",
  64837=>"110001010",
  64838=>"010100101",
  64839=>"101101011",
  64840=>"110000010",
  64841=>"010001110",
  64842=>"100101011",
  64843=>"001101000",
  64844=>"011111101",
  64845=>"011010101",
  64846=>"000011111",
  64847=>"011011001",
  64848=>"111101111",
  64849=>"001110011",
  64850=>"110100111",
  64851=>"000110101",
  64852=>"001101111",
  64853=>"001011001",
  64854=>"010000111",
  64855=>"010110111",
  64856=>"011011010",
  64857=>"101001110",
  64858=>"111110110",
  64859=>"100111011",
  64860=>"111011000",
  64861=>"010011001",
  64862=>"111110001",
  64863=>"000100000",
  64864=>"010010101",
  64865=>"100110011",
  64866=>"010010000",
  64867=>"011001100",
  64868=>"010011100",
  64869=>"101110110",
  64870=>"011011001",
  64871=>"100010111",
  64872=>"101010110",
  64873=>"000101011",
  64874=>"001000000",
  64875=>"100111011",
  64876=>"110111110",
  64877=>"111000000",
  64878=>"011111110",
  64879=>"001010000",
  64880=>"000001011",
  64881=>"000100111",
  64882=>"100000001",
  64883=>"110111110",
  64884=>"001011000",
  64885=>"101110000",
  64886=>"001010110",
  64887=>"010010001",
  64888=>"101101101",
  64889=>"001010010",
  64890=>"101111110",
  64891=>"010010111",
  64892=>"101111011",
  64893=>"000011000",
  64894=>"101011010",
  64895=>"001001100",
  64896=>"110010100",
  64897=>"011101101",
  64898=>"000011110",
  64899=>"111000000",
  64900=>"001010101",
  64901=>"100100100",
  64902=>"111001111",
  64903=>"001001010",
  64904=>"000000011",
  64905=>"110101100",
  64906=>"001110111",
  64907=>"010000001",
  64908=>"110100111",
  64909=>"100111100",
  64910=>"000011000",
  64911=>"101100011",
  64912=>"011000100",
  64913=>"010001000",
  64914=>"111101111",
  64915=>"010100100",
  64916=>"101001111",
  64917=>"000000000",
  64918=>"110001000",
  64919=>"011101000",
  64920=>"101000101",
  64921=>"000110110",
  64922=>"010110001",
  64923=>"011000010",
  64924=>"010010100",
  64925=>"100011101",
  64926=>"010111111",
  64927=>"101000101",
  64928=>"000101110",
  64929=>"001011010",
  64930=>"100100001",
  64931=>"000001100",
  64932=>"010101011",
  64933=>"001000110",
  64934=>"001101000",
  64935=>"010110101",
  64936=>"111011101",
  64937=>"111011010",
  64938=>"000110101",
  64939=>"100000010",
  64940=>"011110100",
  64941=>"001110001",
  64942=>"011011000",
  64943=>"010110011",
  64944=>"101110111",
  64945=>"101011000",
  64946=>"101011000",
  64947=>"010001000",
  64948=>"100010000",
  64949=>"100001000",
  64950=>"011100101",
  64951=>"011101101",
  64952=>"010000101",
  64953=>"011111111",
  64954=>"101010000",
  64955=>"101101111",
  64956=>"001100000",
  64957=>"101010001",
  64958=>"000101111",
  64959=>"111010011",
  64960=>"100101110",
  64961=>"010001101",
  64962=>"001010100",
  64963=>"001110010",
  64964=>"000011000",
  64965=>"110101001",
  64966=>"101001000",
  64967=>"000111111",
  64968=>"111011001",
  64969=>"000110001",
  64970=>"011111111",
  64971=>"011111110",
  64972=>"100000010",
  64973=>"100001101",
  64974=>"100110011",
  64975=>"011101101",
  64976=>"111100011",
  64977=>"111100110",
  64978=>"000011111",
  64979=>"110011011",
  64980=>"000011101",
  64981=>"011010011",
  64982=>"101110100",
  64983=>"000000010",
  64984=>"101100101",
  64985=>"110111001",
  64986=>"011101000",
  64987=>"111000101",
  64988=>"100000111",
  64989=>"010000101",
  64990=>"110100111",
  64991=>"101010100",
  64992=>"111101100",
  64993=>"011000001",
  64994=>"011011001",
  64995=>"011010000",
  64996=>"101010111",
  64997=>"101011010",
  64998=>"011101100",
  64999=>"101001000",
  65000=>"000000010",
  65001=>"001101001",
  65002=>"010011000",
  65003=>"001111010",
  65004=>"101101110",
  65005=>"000010101",
  65006=>"110010010",
  65007=>"010000111",
  65008=>"101110001",
  65009=>"011000010",
  65010=>"110110100",
  65011=>"000110010",
  65012=>"111001011",
  65013=>"100010010",
  65014=>"010010010",
  65015=>"101011111",
  65016=>"010100000",
  65017=>"000101011",
  65018=>"000111000",
  65019=>"110101010",
  65020=>"000111001",
  65021=>"100100010",
  65022=>"101000010",
  65023=>"000011110",
  65024=>"011010100",
  65025=>"011001001",
  65026=>"111001111",
  65027=>"011100011",
  65028=>"000101110",
  65029=>"011000011",
  65030=>"011100011",
  65031=>"001011111",
  65032=>"001111000",
  65033=>"110111011",
  65034=>"110101100",
  65035=>"011000110",
  65036=>"111110100",
  65037=>"111001111",
  65038=>"011100100",
  65039=>"011000101",
  65040=>"111100111",
  65041=>"010100100",
  65042=>"100000111",
  65043=>"101101000",
  65044=>"011001110",
  65045=>"100101011",
  65046=>"100001000",
  65047=>"100110110",
  65048=>"111100101",
  65049=>"010001111",
  65050=>"111100011",
  65051=>"001010000",
  65052=>"010000100",
  65053=>"101110110",
  65054=>"000101111",
  65055=>"100010101",
  65056=>"111001101",
  65057=>"011101100",
  65058=>"000100100",
  65059=>"100001001",
  65060=>"110111111",
  65061=>"000110110",
  65062=>"111111001",
  65063=>"101101011",
  65064=>"100010100",
  65065=>"101001101",
  65066=>"101011111",
  65067=>"111010100",
  65068=>"000101001",
  65069=>"101100010",
  65070=>"101101011",
  65071=>"111101011",
  65072=>"110110111",
  65073=>"111110101",
  65074=>"110000110",
  65075=>"100100111",
  65076=>"010110011",
  65077=>"001101001",
  65078=>"001111111",
  65079=>"101111000",
  65080=>"001100110",
  65081=>"001101101",
  65082=>"110111101",
  65083=>"000010101",
  65084=>"011010111",
  65085=>"111001010",
  65086=>"100101100",
  65087=>"101011111",
  65088=>"111000000",
  65089=>"100010001",
  65090=>"000101111",
  65091=>"010101000",
  65092=>"010111111",
  65093=>"000000101",
  65094=>"100010000",
  65095=>"001010101",
  65096=>"011011001",
  65097=>"101010111",
  65098=>"110001110",
  65099=>"001111001",
  65100=>"101010000",
  65101=>"110110110",
  65102=>"110111101",
  65103=>"011111101",
  65104=>"011111100",
  65105=>"100001000",
  65106=>"110000100",
  65107=>"010000010",
  65108=>"111000110",
  65109=>"000010101",
  65110=>"111101001",
  65111=>"111011100",
  65112=>"110111110",
  65113=>"000100101",
  65114=>"110111010",
  65115=>"000011101",
  65116=>"000001100",
  65117=>"000111101",
  65118=>"111111001",
  65119=>"010000001",
  65120=>"110110011",
  65121=>"001100100",
  65122=>"101011101",
  65123=>"100101101",
  65124=>"110111100",
  65125=>"001110001",
  65126=>"110010101",
  65127=>"100001110",
  65128=>"100111100",
  65129=>"000000011",
  65130=>"010111000",
  65131=>"101010010",
  65132=>"000011100",
  65133=>"111111010",
  65134=>"011011011",
  65135=>"101101011",
  65136=>"100101100",
  65137=>"111011101",
  65138=>"110101001",
  65139=>"100101101",
  65140=>"100111101",
  65141=>"011010001",
  65142=>"101100000",
  65143=>"100111100",
  65144=>"000110100",
  65145=>"100001010",
  65146=>"000110001",
  65147=>"000010110",
  65148=>"001101110",
  65149=>"100110000",
  65150=>"011011000",
  65151=>"001100010",
  65152=>"010010110",
  65153=>"010010101",
  65154=>"011011010",
  65155=>"110000111",
  65156=>"100111011",
  65157=>"000011101",
  65158=>"111000111",
  65159=>"101111000",
  65160=>"010101000",
  65161=>"000100101",
  65162=>"110110110",
  65163=>"111111110",
  65164=>"010011111",
  65165=>"000100011",
  65166=>"010011001",
  65167=>"010000111",
  65168=>"011110111",
  65169=>"111101011",
  65170=>"011101000",
  65171=>"011001111",
  65172=>"010110110",
  65173=>"011111111",
  65174=>"011111011",
  65175=>"011001101",
  65176=>"110010010",
  65177=>"100011000",
  65178=>"011011001",
  65179=>"001100000",
  65180=>"100100110",
  65181=>"101011100",
  65182=>"011111100",
  65183=>"011100100",
  65184=>"000111101",
  65185=>"000000000",
  65186=>"001001111",
  65187=>"010000000",
  65188=>"100101101",
  65189=>"010111011",
  65190=>"101001010",
  65191=>"100111110",
  65192=>"101110111",
  65193=>"010100010",
  65194=>"000000101",
  65195=>"000101000",
  65196=>"000101000",
  65197=>"000101000",
  65198=>"010000011",
  65199=>"011010011",
  65200=>"110110101",
  65201=>"111111000",
  65202=>"011101101",
  65203=>"111100011",
  65204=>"110001001",
  65205=>"101100101",
  65206=>"100011111",
  65207=>"110100111",
  65208=>"101001000",
  65209=>"101001001",
  65210=>"010110001",
  65211=>"100011100",
  65212=>"100011000",
  65213=>"111111100",
  65214=>"011100000",
  65215=>"000101011",
  65216=>"111111110",
  65217=>"010010010",
  65218=>"111110000",
  65219=>"100001110",
  65220=>"100000110",
  65221=>"101111111",
  65222=>"111010010",
  65223=>"010010100",
  65224=>"010000110",
  65225=>"001010010",
  65226=>"000001011",
  65227=>"011011010",
  65228=>"011101011",
  65229=>"110100101",
  65230=>"100101100",
  65231=>"100111111",
  65232=>"111010110",
  65233=>"011111011",
  65234=>"101000000",
  65235=>"110110000",
  65236=>"010001011",
  65237=>"100011001",
  65238=>"101101000",
  65239=>"100010000",
  65240=>"000010110",
  65241=>"110101011",
  65242=>"101000001",
  65243=>"011000001",
  65244=>"110111111",
  65245=>"000001001",
  65246=>"010010000",
  65247=>"010001010",
  65248=>"110100001",
  65249=>"101100111",
  65250=>"010011000",
  65251=>"000001111",
  65252=>"100000101",
  65253=>"001100100",
  65254=>"100111111",
  65255=>"000001110",
  65256=>"110111011",
  65257=>"110000011",
  65258=>"110101110",
  65259=>"001101010",
  65260=>"111101101",
  65261=>"111011111",
  65262=>"110101101",
  65263=>"001100010",
  65264=>"010111010",
  65265=>"110101000",
  65266=>"100111110",
  65267=>"000101000",
  65268=>"110010000",
  65269=>"001100111",
  65270=>"000011100",
  65271=>"110100011",
  65272=>"011101110",
  65273=>"111100001",
  65274=>"010001101",
  65275=>"100011101",
  65276=>"111110101",
  65277=>"100100110",
  65278=>"001011100",
  65279=>"010110011",
  65280=>"110101010",
  65281=>"110110000",
  65282=>"101101010",
  65283=>"100101100",
  65284=>"010001011",
  65285=>"101001100",
  65286=>"000100011",
  65287=>"110011001",
  65288=>"111010000",
  65289=>"000011000",
  65290=>"011000000",
  65291=>"100000011",
  65292=>"011101000",
  65293=>"111101111",
  65294=>"010011000",
  65295=>"110010010",
  65296=>"011100111",
  65297=>"010011101",
  65298=>"111100010",
  65299=>"001000000",
  65300=>"101000010",
  65301=>"000111010",
  65302=>"000000011",
  65303=>"011100101",
  65304=>"000110110",
  65305=>"100000011",
  65306=>"111001011",
  65307=>"001010101",
  65308=>"001001110",
  65309=>"110011010",
  65310=>"010010010",
  65311=>"001100010",
  65312=>"000001000",
  65313=>"001101101",
  65314=>"010000111",
  65315=>"100011011",
  65316=>"000010001",
  65317=>"100101101",
  65318=>"011100001",
  65319=>"111111111",
  65320=>"001001010",
  65321=>"100000010",
  65322=>"001000110",
  65323=>"111010000",
  65324=>"001011110",
  65325=>"100011011",
  65326=>"000001001",
  65327=>"111100001",
  65328=>"011011110",
  65329=>"111000010",
  65330=>"110001011",
  65331=>"000010001",
  65332=>"011001010",
  65333=>"100010010",
  65334=>"100111111",
  65335=>"100110111",
  65336=>"000010000",
  65337=>"101010100",
  65338=>"111101000",
  65339=>"001100011",
  65340=>"001110000",
  65341=>"000011110",
  65342=>"011001000",
  65343=>"111011011",
  65344=>"010000001",
  65345=>"010000111",
  65346=>"101101011",
  65347=>"011111100",
  65348=>"111110101",
  65349=>"011101011",
  65350=>"101000000",
  65351=>"010110011",
  65352=>"001011100",
  65353=>"000000101",
  65354=>"001001110",
  65355=>"110101010",
  65356=>"000011001",
  65357=>"100000110",
  65358=>"000100111",
  65359=>"100111001",
  65360=>"110100101",
  65361=>"100111001",
  65362=>"001110011",
  65363=>"011011001",
  65364=>"100000001",
  65365=>"100111010",
  65366=>"010010001",
  65367=>"100101111",
  65368=>"010100000",
  65369=>"111000010",
  65370=>"010011001",
  65371=>"110100100",
  65372=>"101101001",
  65373=>"000010011",
  65374=>"011111011",
  65375=>"111010010",
  65376=>"110101110",
  65377=>"111000000",
  65378=>"001001001",
  65379=>"000101110",
  65380=>"000110101",
  65381=>"111010010",
  65382=>"110001011",
  65383=>"010001110",
  65384=>"001000001",
  65385=>"111101010",
  65386=>"111010101",
  65387=>"010111001",
  65388=>"010001001",
  65389=>"111100110",
  65390=>"011000100",
  65391=>"011000000",
  65392=>"101101000",
  65393=>"110001100",
  65394=>"011000101",
  65395=>"111111001",
  65396=>"101001000",
  65397=>"100000110",
  65398=>"001010000",
  65399=>"111000000",
  65400=>"010010111",
  65401=>"111010101",
  65402=>"110101010",
  65403=>"101000001",
  65404=>"010000000",
  65405=>"001000011",
  65406=>"010001011",
  65407=>"000011000",
  65408=>"001101001",
  65409=>"000110000",
  65410=>"010010100",
  65411=>"000110111",
  65412=>"011010110",
  65413=>"011000100",
  65414=>"100111111",
  65415=>"011100000",
  65416=>"111101011",
  65417=>"000111111",
  65418=>"110010100",
  65419=>"010100111",
  65420=>"000110000",
  65421=>"100111111",
  65422=>"110101010",
  65423=>"101101111",
  65424=>"000001111",
  65425=>"000010010",
  65426=>"000010010",
  65427=>"001100110",
  65428=>"001001111",
  65429=>"110001000",
  65430=>"111000110",
  65431=>"111001100",
  65432=>"101001001",
  65433=>"010100100",
  65434=>"000111000",
  65435=>"111111111",
  65436=>"000001100",
  65437=>"010100100",
  65438=>"111100000",
  65439=>"011000001",
  65440=>"001011100",
  65441=>"000111000",
  65442=>"110110100",
  65443=>"101011011",
  65444=>"101011011",
  65445=>"001001001",
  65446=>"011110100",
  65447=>"101100001",
  65448=>"011111111",
  65449=>"100011110",
  65450=>"011111100",
  65451=>"101100001",
  65452=>"000001010",
  65453=>"001111000",
  65454=>"000111010",
  65455=>"011001100",
  65456=>"001110100",
  65457=>"001001110",
  65458=>"101101001",
  65459=>"010000111",
  65460=>"001000111",
  65461=>"100110111",
  65462=>"010000000",
  65463=>"101000010",
  65464=>"100010100",
  65465=>"011001001",
  65466=>"000100111",
  65467=>"001011101",
  65468=>"011001001",
  65469=>"110101100",
  65470=>"000000110",
  65471=>"100000000",
  65472=>"111100110",
  65473=>"111101111",
  65474=>"000110110",
  65475=>"000010001",
  65476=>"001101101",
  65477=>"111100011",
  65478=>"111111111",
  65479=>"110110010",
  65480=>"100000011",
  65481=>"011010110",
  65482=>"100001011",
  65483=>"110010110",
  65484=>"000100011",
  65485=>"001100000",
  65486=>"010110010",
  65487=>"101101000",
  65488=>"011010110",
  65489=>"011110111",
  65490=>"100011110",
  65491=>"110101011",
  65492=>"000000101",
  65493=>"011001011",
  65494=>"000000101",
  65495=>"101110111",
  65496=>"111100001",
  65497=>"011100110",
  65498=>"011100111",
  65499=>"111001000",
  65500=>"110110000",
  65501=>"001100011",
  65502=>"101101110",
  65503=>"001001110",
  65504=>"101111101",
  65505=>"001001111",
  65506=>"101011101",
  65507=>"111101100",
  65508=>"000000100",
  65509=>"100100000",
  65510=>"000101000",
  65511=>"101001110",
  65512=>"000001011",
  65513=>"011000111",
  65514=>"100010101",
  65515=>"010110011",
  65516=>"110100110",
  65517=>"001001001",
  65518=>"110001000",
  65519=>"100011110",
  65520=>"101010000",
  65521=>"011011010",
  65522=>"100000011",
  65523=>"011011011",
  65524=>"110011111",
  65525=>"010011100",
  65526=>"110111011",
  65527=>"010100111",
  65528=>"111001011",
  65529=>"011101100",
  65530=>"110000001",
  65531=>"000011001",
  65532=>"100010101",
  65533=>"100011110",
  65534=>"100010010",
  65535=>"010111111");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;