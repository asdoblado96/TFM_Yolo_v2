LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L6_1_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(6)-1 DOWNTO 0));
END L6_1_WROM;

ARCHITECTURE RTL OF L6_1_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"101100101",
  1=>"110100011",
  2=>"000100101",
  3=>"111011011",
  4=>"110110100",
  5=>"000000111",
  6=>"111100111",
  7=>"011111101",
  8=>"101101011",
  9=>"100100000",
  10=>"000010110",
  11=>"110101011",
  12=>"110111011",
  13=>"000010011",
  14=>"000100000",
  15=>"011100111",
  16=>"111100100",
  17=>"110000010",
  18=>"000111010",
  19=>"000001011",
  20=>"000110000",
  21=>"111100111",
  22=>"110100000",
  23=>"010111111",
  24=>"100000100",
  25=>"011010001",
  26=>"000010000",
  27=>"000010011",
  28=>"110100100",
  29=>"101000010",
  30=>"111100001",
  31=>"111111000",
  32=>"101100000",
  33=>"100100100",
  34=>"110011011",
  35=>"111100111",
  36=>"110100110",
  37=>"111100111",
  38=>"111100100",
  39=>"011100000",
  40=>"101111010",
  41=>"110000000",
  42=>"001101111",
  43=>"110101111",
  44=>"000111001",
  45=>"011100111",
  46=>"100110111",
  47=>"110011010",
  48=>"110000000",
  49=>"111111111",
  50=>"001111111",
  51=>"000110000",
  52=>"000111100",
  53=>"100011011",
  54=>"110100100",
  55=>"101100100",
  56=>"111111000",
  57=>"111100101",
  58=>"001010010",
  59=>"100100010",
  60=>"110010000",
  61=>"011111010",
  62=>"000000001",
  63=>"101101100",
  64=>"100110111",
  65=>"110100001",
  66=>"100110001",
  67=>"011001000",
  68=>"111000011",
  69=>"110000000",
  70=>"100100101",
  71=>"011111000",
  72=>"101100010",
  73=>"010011011",
  74=>"000011000",
  75=>"101011000",
  76=>"111100100",
  77=>"001101000",
  78=>"101101100",
  79=>"001001101",
  80=>"001011101",
  81=>"011110111",
  82=>"111000000",
  83=>"000000000",
  84=>"000100001",
  85=>"001100000",
  86=>"000110111",
  87=>"001001101",
  88=>"100010010",
  89=>"100111101",
  90=>"000000000",
  91=>"000000000",
  92=>"000111000",
  93=>"100101100",
  94=>"111111100",
  95=>"111110101",
  96=>"010110000",
  97=>"101000111",
  98=>"111100111",
  99=>"010110110",
  100=>"010010111",
  101=>"000011000",
  102=>"011011010",
  103=>"101100110",
  104=>"100110111",
  105=>"111111011",
  106=>"000100100",
  107=>"111011100",
  108=>"101100111",
  109=>"011011000",
  110=>"110100100",
  111=>"010010011",
  112=>"100111011",
  113=>"100111011",
  114=>"001100110",
  115=>"000000000",
  116=>"111100100",
  117=>"000100000",
  118=>"000001011",
  119=>"011000011",
  120=>"101011111",
  121=>"000000001",
  122=>"010010011",
  123=>"011111000",
  124=>"100100101",
  125=>"010010011",
  126=>"101100100",
  127=>"000010101",
  128=>"000101100",
  129=>"111100000",
  130=>"010111100",
  131=>"100001001",
  132=>"111101101",
  133=>"110001000",
  134=>"001001000",
  135=>"100100000",
  136=>"100111111",
  137=>"000000000",
  138=>"011010011",
  139=>"011001100",
  140=>"100111111",
  141=>"000011011",
  142=>"101101011",
  143=>"000001001",
  144=>"110111110",
  145=>"111100100",
  146=>"000001110",
  147=>"111100001",
  148=>"000011000",
  149=>"100100100",
  150=>"001011111",
  151=>"010010110",
  152=>"011011010",
  153=>"101011011",
  154=>"100100101",
  155=>"100100011",
  156=>"000000001",
  157=>"111111111",
  158=>"011111111",
  159=>"000000110",
  160=>"100100000",
  161=>"110100111",
  162=>"011011011",
  163=>"000011000",
  164=>"000011011",
  165=>"010011010",
  166=>"110101011",
  167=>"000000011",
  168=>"010000111",
  169=>"100111011",
  170=>"101100101",
  171=>"010100111",
  172=>"111000001",
  173=>"000000000",
  174=>"010010111",
  175=>"000000000",
  176=>"101000001",
  177=>"001011110",
  178=>"110000100",
  179=>"000000000",
  180=>"101000000",
  181=>"111011111",
  182=>"111001100",
  183=>"100110111",
  184=>"100001000",
  185=>"011011011",
  186=>"000010110",
  187=>"001011110",
  188=>"111011010",
  189=>"011001000",
  190=>"011001001",
  191=>"000000000",
  192=>"100000100",
  193=>"011011011",
  194=>"011011100",
  195=>"001011011",
  196=>"011011000",
  197=>"100100000",
  198=>"111000010",
  199=>"011011111",
  200=>"100111111",
  201=>"000011000",
  202=>"100001101",
  203=>"100100100",
  204=>"111100100",
  205=>"101111111",
  206=>"000100100",
  207=>"100100011",
  208=>"110000000",
  209=>"101101111",
  210=>"111100011",
  211=>"010100111",
  212=>"011100000",
  213=>"010001101",
  214=>"111010000",
  215=>"011011000",
  216=>"000011011",
  217=>"011000100",
  218=>"001001001",
  219=>"000000011",
  220=>"001101111",
  221=>"100110100",
  222=>"110011111",
  223=>"111100111",
  224=>"000011111",
  225=>"000000001",
  226=>"111001100",
  227=>"100110000",
  228=>"100000100",
  229=>"111011001",
  230=>"111111000",
  231=>"000000001",
  232=>"010000101",
  233=>"100000011",
  234=>"100001111",
  235=>"111111111",
  236=>"100100000",
  237=>"100100000",
  238=>"010110000",
  239=>"001100101",
  240=>"110100010",
  241=>"110000100",
  242=>"000000000",
  243=>"010111010",
  244=>"010110111",
  245=>"000000000",
  246=>"000000000",
  247=>"111100100",
  248=>"011100111",
  249=>"011000000",
  250=>"110110011",
  251=>"100100101",
  252=>"111111111",
  253=>"000100100",
  254=>"001100100",
  255=>"101100000",
  256=>"010011100",
  257=>"110111111",
  258=>"000000111",
  259=>"111111101",
  260=>"011001001",
  261=>"011000111",
  262=>"010010000",
  263=>"111010111",
  264=>"001001101",
  265=>"000000111",
  266=>"111011000",
  267=>"111011000",
  268=>"110010000",
  269=>"001001000",
  270=>"111011000",
  271=>"000111111",
  272=>"101000000",
  273=>"000111011",
  274=>"001000111",
  275=>"000110001",
  276=>"010110100",
  277=>"111011011",
  278=>"001000000",
  279=>"110011100",
  280=>"000011000",
  281=>"000000010",
  282=>"101101100",
  283=>"010111111",
  284=>"000001000",
  285=>"111001000",
  286=>"110100111",
  287=>"111111000",
  288=>"000000100",
  289=>"010011100",
  290=>"000110000",
  291=>"000000000",
  292=>"111001000",
  293=>"000000000",
  294=>"111111110",
  295=>"000000111",
  296=>"100100111",
  297=>"100000000",
  298=>"010000000",
  299=>"000010000",
  300=>"111111000",
  301=>"000000000",
  302=>"010010100",
  303=>"110010100",
  304=>"100100100",
  305=>"001011000",
  306=>"000111111",
  307=>"111111010",
  308=>"010111000",
  309=>"110110011",
  310=>"011011000",
  311=>"010111011",
  312=>"000000111",
  313=>"100111011",
  314=>"100100000",
  315=>"000101000",
  316=>"010011000",
  317=>"011011111",
  318=>"000000000",
  319=>"110000001",
  320=>"000111111",
  321=>"111000101",
  322=>"000000111",
  323=>"110100111",
  324=>"101010010",
  325=>"000010011",
  326=>"110110000",
  327=>"001000101",
  328=>"111111110",
  329=>"101100000",
  330=>"001111000",
  331=>"111111000",
  332=>"000000000",
  333=>"110111111",
  334=>"100100110",
  335=>"000000011",
  336=>"111101000",
  337=>"000111111",
  338=>"110011111",
  339=>"001000010",
  340=>"111110000",
  341=>"110110010",
  342=>"110100000",
  343=>"110011101",
  344=>"100111011",
  345=>"011001000",
  346=>"011000000",
  347=>"100100000",
  348=>"000010000",
  349=>"001101000",
  350=>"100100111",
  351=>"101001001",
  352=>"000000000",
  353=>"010101111",
  354=>"000111111",
  355=>"111001000",
  356=>"111101001",
  357=>"101100010",
  358=>"110111000",
  359=>"000000001",
  360=>"010011000",
  361=>"000111111",
  362=>"100100111",
  363=>"111110100",
  364=>"000111111",
  365=>"111111011",
  366=>"111111000",
  367=>"000111010",
  368=>"111010000",
  369=>"110000110",
  370=>"110110000",
  371=>"010011000",
  372=>"000000000",
  373=>"000000111",
  374=>"010111000",
  375=>"000000111",
  376=>"000000000",
  377=>"010011010",
  378=>"011111111",
  379=>"001000111",
  380=>"011110110",
  381=>"100001011",
  382=>"111111100",
  383=>"111001001",
  384=>"110000011",
  385=>"110000010",
  386=>"000100100",
  387=>"110111111",
  388=>"010000111",
  389=>"000001010",
  390=>"100100000",
  391=>"010111011",
  392=>"101101000",
  393=>"111111000",
  394=>"000000001",
  395=>"000000111",
  396=>"010101100",
  397=>"111001000",
  398=>"010000011",
  399=>"101001010",
  400=>"111100000",
  401=>"000100000",
  402=>"111111000",
  403=>"111111110",
  404=>"111110010",
  405=>"000101111",
  406=>"000010111",
  407=>"111000000",
  408=>"001000100",
  409=>"111011000",
  410=>"111111111",
  411=>"000000111",
  412=>"010111001",
  413=>"111000000",
  414=>"010000000",
  415=>"101000111",
  416=>"001011110",
  417=>"010010011",
  418=>"101010110",
  419=>"000111111",
  420=>"100111111",
  421=>"010111110",
  422=>"010000001",
  423=>"111011000",
  424=>"000001111",
  425=>"111000000",
  426=>"111101111",
  427=>"001100100",
  428=>"000000111",
  429=>"000000010",
  430=>"111011001",
  431=>"011000101",
  432=>"000000111",
  433=>"111111111",
  434=>"111111000",
  435=>"100111000",
  436=>"111111000",
  437=>"011100000",
  438=>"010100110",
  439=>"111011000",
  440=>"110111000",
  441=>"011011011",
  442=>"010111100",
  443=>"111111100",
  444=>"000011010",
  445=>"111000001",
  446=>"000001111",
  447=>"010111000",
  448=>"101100100",
  449=>"010111000",
  450=>"000000000",
  451=>"111111100",
  452=>"000000000",
  453=>"110100000",
  454=>"001011111",
  455=>"111111110",
  456=>"101000111",
  457=>"000001001",
  458=>"000010110",
  459=>"111111011",
  460=>"111100000",
  461=>"010011001",
  462=>"111000000",
  463=>"010010111",
  464=>"111000000",
  465=>"010001000",
  466=>"010010111",
  467=>"000000000",
  468=>"000000111",
  469=>"111111000",
  470=>"100000100",
  471=>"010000000",
  472=>"000000000",
  473=>"011111111",
  474=>"100100001",
  475=>"000000000",
  476=>"010000000",
  477=>"111000100",
  478=>"111111000",
  479=>"101101101",
  480=>"000001111",
  481=>"111001111",
  482=>"000000000",
  483=>"111111000",
  484=>"001001000",
  485=>"111111000",
  486=>"011000111",
  487=>"010110000",
  488=>"000000000",
  489=>"000000000",
  490=>"111111000",
  491=>"101101111",
  492=>"111011010",
  493=>"000100010",
  494=>"011011001",
  495=>"010101000",
  496=>"010000000",
  497=>"011001000",
  498=>"010111111",
  499=>"111000000",
  500=>"000001001",
  501=>"111001000",
  502=>"000101000",
  503=>"000101101",
  504=>"110111111",
  505=>"000010000",
  506=>"000111100",
  507=>"111101000",
  508=>"000000010",
  509=>"111010011",
  510=>"101101001",
  511=>"000000111",
  512=>"101000100",
  513=>"010000000",
  514=>"110110100",
  515=>"000111101",
  516=>"000101111",
  517=>"111111111",
  518=>"111011000",
  519=>"010111001",
  520=>"001000001",
  521=>"000110110",
  522=>"000000000",
  523=>"001000000",
  524=>"000000000",
  525=>"000000000",
  526=>"100000000",
  527=>"011001111",
  528=>"000000000",
  529=>"010111110",
  530=>"111100000",
  531=>"000000000",
  532=>"111101111",
  533=>"001101111",
  534=>"111011001",
  535=>"110111010",
  536=>"001001001",
  537=>"010111111",
  538=>"000000100",
  539=>"000010110",
  540=>"000010000",
  541=>"111000000",
  542=>"000001111",
  543=>"111011000",
  544=>"011111011",
  545=>"000000111",
  546=>"111001101",
  547=>"101101000",
  548=>"010000000",
  549=>"000001100",
  550=>"111001000",
  551=>"000111000",
  552=>"101111111",
  553=>"000000111",
  554=>"110000000",
  555=>"000111000",
  556=>"111111000",
  557=>"000101000",
  558=>"011010101",
  559=>"100000111",
  560=>"111000000",
  561=>"001000000",
  562=>"000000011",
  563=>"001111111",
  564=>"110000001",
  565=>"100001101",
  566=>"000000000",
  567=>"001000001",
  568=>"000001000",
  569=>"000101111",
  570=>"110111111",
  571=>"111001111",
  572=>"000000001",
  573=>"111111111",
  574=>"000000000",
  575=>"001001001",
  576=>"000010011",
  577=>"000000010",
  578=>"111111111",
  579=>"010000000",
  580=>"000000000",
  581=>"110000111",
  582=>"111111110",
  583=>"001100111",
  584=>"011111000",
  585=>"001000000",
  586=>"000100111",
  587=>"000000011",
  588=>"101100111",
  589=>"110000010",
  590=>"010000010",
  591=>"111001010",
  592=>"000011000",
  593=>"111111111",
  594=>"101000111",
  595=>"000100000",
  596=>"110010000",
  597=>"000000000",
  598=>"100100110",
  599=>"011000000",
  600=>"111001001",
  601=>"111100000",
  602=>"111110000",
  603=>"100101111",
  604=>"001000101",
  605=>"010100000",
  606=>"110111110",
  607=>"000000000",
  608=>"001001111",
  609=>"111111101",
  610=>"001101000",
  611=>"111111001",
  612=>"000000000",
  613=>"111111100",
  614=>"111000000",
  615=>"111010000",
  616=>"011001000",
  617=>"101111101",
  618=>"010111111",
  619=>"111111111",
  620=>"101000100",
  621=>"111111111",
  622=>"111000000",
  623=>"000111111",
  624=>"100000000",
  625=>"010000000",
  626=>"000000000",
  627=>"001000000",
  628=>"000111010",
  629=>"000000110",
  630=>"000111111",
  631=>"000000001",
  632=>"110111010",
  633=>"101111000",
  634=>"100000000",
  635=>"000001000",
  636=>"001001001",
  637=>"110010010",
  638=>"110110000",
  639=>"111010000",
  640=>"111111100",
  641=>"000111111",
  642=>"000111111",
  643=>"111111111",
  644=>"000000110",
  645=>"110110010",
  646=>"110100000",
  647=>"100100001",
  648=>"000001000",
  649=>"110001001",
  650=>"111101011",
  651=>"001011111",
  652=>"000111100",
  653=>"111111011",
  654=>"000000000",
  655=>"001000000",
  656=>"110100010",
  657=>"111111000",
  658=>"111111010",
  659=>"111101011",
  660=>"000100000",
  661=>"000111111",
  662=>"111101000",
  663=>"010010000",
  664=>"101000000",
  665=>"000100010",
  666=>"101000000",
  667=>"010111111",
  668=>"000000110",
  669=>"000000011",
  670=>"001101111",
  671=>"111000000",
  672=>"111111001",
  673=>"111111111",
  674=>"000000000",
  675=>"111100000",
  676=>"101000111",
  677=>"110001011",
  678=>"011000100",
  679=>"000100111",
  680=>"010101001",
  681=>"000001110",
  682=>"001100000",
  683=>"000000010",
  684=>"111111011",
  685=>"000000000",
  686=>"110100000",
  687=>"111111111",
  688=>"111111111",
  689=>"001100000",
  690=>"111011111",
  691=>"110000000",
  692=>"011000000",
  693=>"001000110",
  694=>"111100100",
  695=>"001111100",
  696=>"000000000",
  697=>"000001001",
  698=>"100100111",
  699=>"000101111",
  700=>"111010110",
  701=>"000111110",
  702=>"000000100",
  703=>"100000000",
  704=>"011111001",
  705=>"000110010",
  706=>"111011000",
  707=>"001001000",
  708=>"000000000",
  709=>"111000100",
  710=>"111111111",
  711=>"100111000",
  712=>"110001000",
  713=>"110111111",
  714=>"010000001",
  715=>"111111000",
  716=>"111011000",
  717=>"111000001",
  718=>"101000000",
  719=>"000111011",
  720=>"011110000",
  721=>"010000000",
  722=>"000000001",
  723=>"010111111",
  724=>"000010010",
  725=>"000111000",
  726=>"000000000",
  727=>"111101001",
  728=>"010000000",
  729=>"000000000",
  730=>"110111111",
  731=>"111111111",
  732=>"000000000",
  733=>"001111111",
  734=>"110000010",
  735=>"000001111",
  736=>"010111000",
  737=>"010110000",
  738=>"000110110",
  739=>"011111000",
  740=>"101010000",
  741=>"000101111",
  742=>"000000000",
  743=>"000111000",
  744=>"110110111",
  745=>"001000000",
  746=>"000000000",
  747=>"001010111",
  748=>"000000111",
  749=>"111111110",
  750=>"010110111",
  751=>"000000111",
  752=>"001000000",
  753=>"101101001",
  754=>"111111101",
  755=>"110010010",
  756=>"001001001",
  757=>"111111011",
  758=>"010010111",
  759=>"110111010",
  760=>"000111000",
  761=>"111111111",
  762=>"111111111",
  763=>"011000000",
  764=>"011000000",
  765=>"111000000",
  766=>"001000001",
  767=>"111011000",
  768=>"110011001",
  769=>"000000011",
  770=>"101000111",
  771=>"110101101",
  772=>"010111110",
  773=>"000000101",
  774=>"101000101",
  775=>"010000000",
  776=>"000000000",
  777=>"011010000",
  778=>"000111110",
  779=>"100011111",
  780=>"000000000",
  781=>"000111110",
  782=>"011011010",
  783=>"011110100",
  784=>"000010111",
  785=>"010110110",
  786=>"010001100",
  787=>"000111111",
  788=>"111100011",
  789=>"111000000",
  790=>"000000100",
  791=>"010010010",
  792=>"001000100",
  793=>"111111101",
  794=>"000000100",
  795=>"000100010",
  796=>"101001000",
  797=>"111000111",
  798=>"111110001",
  799=>"000000100",
  800=>"111001101",
  801=>"010010101",
  802=>"101101000",
  803=>"111000110",
  804=>"100100000",
  805=>"110110100",
  806=>"101000001",
  807=>"000110111",
  808=>"111000111",
  809=>"000001000",
  810=>"000111000",
  811=>"000000100",
  812=>"000011011",
  813=>"010111111",
  814=>"000101110",
  815=>"110110110",
  816=>"001000001",
  817=>"001101111",
  818=>"111000001",
  819=>"110000100",
  820=>"101111111",
  821=>"101111110",
  822=>"001011110",
  823=>"101000001",
  824=>"000001111",
  825=>"111001000",
  826=>"001000000",
  827=>"000000101",
  828=>"110100100",
  829=>"000111001",
  830=>"000000101",
  831=>"001001110",
  832=>"111111101",
  833=>"111111000",
  834=>"000100010",
  835=>"110000011",
  836=>"111111011",
  837=>"111111110",
  838=>"000000100",
  839=>"111011001",
  840=>"110010011",
  841=>"111111101",
  842=>"000001111",
  843=>"100000001",
  844=>"000000000",
  845=>"011001000",
  846=>"100100110",
  847=>"000011101",
  848=>"111111110",
  849=>"010000000",
  850=>"000000000",
  851=>"000101100",
  852=>"000000111",
  853=>"010111010",
  854=>"010100111",
  855=>"101111111",
  856=>"111100100",
  857=>"011101100",
  858=>"001001001",
  859=>"111111110",
  860=>"001000101",
  861=>"010001001",
  862=>"101000001",
  863=>"001000100",
  864=>"001000000",
  865=>"101000101",
  866=>"111111011",
  867=>"101100100",
  868=>"110110100",
  869=>"000111010",
  870=>"110111000",
  871=>"000000110",
  872=>"111111100",
  873=>"111110000",
  874=>"111000000",
  875=>"111000000",
  876=>"111001000",
  877=>"110110010",
  878=>"000010000",
  879=>"010001111",
  880=>"100100000",
  881=>"010000000",
  882=>"101110111",
  883=>"111001100",
  884=>"000101111",
  885=>"000000000",
  886=>"000111111",
  887=>"101101000",
  888=>"000100100",
  889=>"010011100",
  890=>"000000000",
  891=>"001101100",
  892=>"100110011",
  893=>"110100001",
  894=>"000000101",
  895=>"000010000",
  896=>"010010101",
  897=>"010101000",
  898=>"000000000",
  899=>"011011111",
  900=>"010111100",
  901=>"111000000",
  902=>"011011000",
  903=>"001010001",
  904=>"011001001",
  905=>"111000110",
  906=>"111000000",
  907=>"111111111",
  908=>"111001001",
  909=>"100000101",
  910=>"000000111",
  911=>"010000000",
  912=>"111100100",
  913=>"110100000",
  914=>"111110000",
  915=>"010000000",
  916=>"000111111",
  917=>"100100001",
  918=>"010111110",
  919=>"111100000",
  920=>"111111111",
  921=>"111111110",
  922=>"001111000",
  923=>"000000111",
  924=>"000000000",
  925=>"111111011",
  926=>"111100111",
  927=>"001101000",
  928=>"000101110",
  929=>"111101111",
  930=>"111001111",
  931=>"000010011",
  932=>"000001111",
  933=>"111011011",
  934=>"111001111",
  935=>"001111110",
  936=>"000000111",
  937=>"000010111",
  938=>"000000111",
  939=>"010111000",
  940=>"000000100",
  941=>"010010000",
  942=>"110100110",
  943=>"110000110",
  944=>"111001100",
  945=>"001011001",
  946=>"101101101",
  947=>"111101010",
  948=>"100100111",
  949=>"101101110",
  950=>"000010011",
  951=>"110110010",
  952=>"001111010",
  953=>"000110000",
  954=>"010010001",
  955=>"111110111",
  956=>"110010100",
  957=>"111111111",
  958=>"000110010",
  959=>"110111001",
  960=>"001000001",
  961=>"011000000",
  962=>"011011010",
  963=>"011011001",
  964=>"110111000",
  965=>"001111011",
  966=>"111000000",
  967=>"111111111",
  968=>"000111111",
  969=>"010000000",
  970=>"111110010",
  971=>"100000111",
  972=>"111100100",
  973=>"001011110",
  974=>"100000000",
  975=>"000000111",
  976=>"000010000",
  977=>"000000010",
  978=>"101010111",
  979=>"011111111",
  980=>"000000111",
  981=>"011100100",
  982=>"101000111",
  983=>"111000000",
  984=>"101001111",
  985=>"111000000",
  986=>"010001110",
  987=>"100100000",
  988=>"010101010",
  989=>"001000001",
  990=>"111010011",
  991=>"000001111",
  992=>"110000000",
  993=>"111000001",
  994=>"010000001",
  995=>"000001000",
  996=>"011000000",
  997=>"000000000",
  998=>"111111111",
  999=>"010000000",
  1000=>"000001111",
  1001=>"000010111",
  1002=>"011111011",
  1003=>"111111101",
  1004=>"000000000",
  1005=>"100000000",
  1006=>"000000000",
  1007=>"000000000",
  1008=>"000010111",
  1009=>"100100100",
  1010=>"001000111",
  1011=>"000011011",
  1012=>"010111101",
  1013=>"101000000",
  1014=>"010000100",
  1015=>"110010000",
  1016=>"111111000",
  1017=>"010111111",
  1018=>"111101111",
  1019=>"000001010",
  1020=>"001001101",
  1021=>"000000000",
  1022=>"010001101",
  1023=>"110000000",
  1024=>"011010100",
  1025=>"100000110",
  1026=>"001000100",
  1027=>"000000011",
  1028=>"000111110",
  1029=>"110010000",
  1030=>"110010011",
  1031=>"111000100",
  1032=>"100101101",
  1033=>"000000000",
  1034=>"111001100",
  1035=>"100100100",
  1036=>"011000000",
  1037=>"000100001",
  1038=>"000101001",
  1039=>"011010001",
  1040=>"100011011",
  1041=>"111100100",
  1042=>"000100000",
  1043=>"111100100",
  1044=>"111001010",
  1045=>"111100100",
  1046=>"000000110",
  1047=>"001000110",
  1048=>"100100100",
  1049=>"000000011",
  1050=>"100100100",
  1051=>"100100111",
  1052=>"000000001",
  1053=>"100100000",
  1054=>"111110110",
  1055=>"111100101",
  1056=>"111011000",
  1057=>"100111100",
  1058=>"000011001",
  1059=>"000011000",
  1060=>"000011000",
  1061=>"100100110",
  1062=>"000000101",
  1063=>"100000011",
  1064=>"011111101",
  1065=>"111011101",
  1066=>"011001000",
  1067=>"000100100",
  1068=>"011011111",
  1069=>"011000011",
  1070=>"111100111",
  1071=>"100000000",
  1072=>"000000000",
  1073=>"001001011",
  1074=>"011110101",
  1075=>"100100100",
  1076=>"000001000",
  1077=>"111011001",
  1078=>"000100100",
  1079=>"111000010",
  1080=>"111010000",
  1081=>"111100001",
  1082=>"000001000",
  1083=>"010000000",
  1084=>"011101010",
  1085=>"010111000",
  1086=>"100100100",
  1087=>"110111101",
  1088=>"011011000",
  1089=>"110100010",
  1090=>"011010010",
  1091=>"001111111",
  1092=>"111110000",
  1093=>"111111101",
  1094=>"110110000",
  1095=>"111100100",
  1096=>"000110111",
  1097=>"001000000",
  1098=>"000100111",
  1099=>"011111101",
  1100=>"100110000",
  1101=>"101100010",
  1102=>"000011101",
  1103=>"111100110",
  1104=>"100000000",
  1105=>"011111111",
  1106=>"110000011",
  1107=>"101000101",
  1108=>"101100100",
  1109=>"001010110",
  1110=>"001001000",
  1111=>"001000001",
  1112=>"111100100",
  1113=>"000000001",
  1114=>"001110110",
  1115=>"000111011",
  1116=>"000100010",
  1117=>"000000001",
  1118=>"111111111",
  1119=>"100111111",
  1120=>"010111000",
  1121=>"000111111",
  1122=>"100100101",
  1123=>"000000100",
  1124=>"111101100",
  1125=>"100100011",
  1126=>"011101000",
  1127=>"000000000",
  1128=>"011011000",
  1129=>"000101000",
  1130=>"100001100",
  1131=>"011100001",
  1132=>"011011000",
  1133=>"011000111",
  1134=>"000010011",
  1135=>"101100110",
  1136=>"011011011",
  1137=>"101001111",
  1138=>"000000010",
  1139=>"011011000",
  1140=>"000011110",
  1141=>"100100101",
  1142=>"101100010",
  1143=>"000000111",
  1144=>"011000111",
  1145=>"011100011",
  1146=>"000011011",
  1147=>"110000000",
  1148=>"110011100",
  1149=>"010000000",
  1150=>"000000101",
  1151=>"001111011",
  1152=>"001011000",
  1153=>"110111000",
  1154=>"000100000",
  1155=>"000100000",
  1156=>"110000100",
  1157=>"111000000",
  1158=>"000001011",
  1159=>"100000000",
  1160=>"000010111",
  1161=>"001000011",
  1162=>"001101001",
  1163=>"100000000",
  1164=>"000100000",
  1165=>"000000011",
  1166=>"100100010",
  1167=>"101000010",
  1168=>"100111110",
  1169=>"101100101",
  1170=>"100100110",
  1171=>"101001111",
  1172=>"100000010",
  1173=>"010000100",
  1174=>"100111111",
  1175=>"000011011",
  1176=>"011111011",
  1177=>"101100110",
  1178=>"000111111",
  1179=>"000000001",
  1180=>"000000111",
  1181=>"000100000",
  1182=>"111011111",
  1183=>"000000000",
  1184=>"000100100",
  1185=>"100000000",
  1186=>"000100111",
  1187=>"011100010",
  1188=>"110100011",
  1189=>"101000110",
  1190=>"000011011",
  1191=>"111100100",
  1192=>"111100111",
  1193=>"010110100",
  1194=>"011111110",
  1195=>"100100100",
  1196=>"000011000",
  1197=>"100100110",
  1198=>"100001001",
  1199=>"011010110",
  1200=>"011011000",
  1201=>"100100100",
  1202=>"111111111",
  1203=>"000000111",
  1204=>"011001001",
  1205=>"000100000",
  1206=>"011011001",
  1207=>"101000011",
  1208=>"110110001",
  1209=>"100000111",
  1210=>"011100111",
  1211=>"111010101",
  1212=>"011011000",
  1213=>"010111111",
  1214=>"001001011",
  1215=>"011000100",
  1216=>"101000001",
  1217=>"100100000",
  1218=>"100100000",
  1219=>"001000000",
  1220=>"000011000",
  1221=>"000110100",
  1222=>"111110000",
  1223=>"100011011",
  1224=>"111100001",
  1225=>"111111000",
  1226=>"111101110",
  1227=>"001101001",
  1228=>"111110110",
  1229=>"000011001",
  1230=>"100001001",
  1231=>"011111000",
  1232=>"111001000",
  1233=>"000110001",
  1234=>"100011011",
  1235=>"000000001",
  1236=>"001111000",
  1237=>"111001001",
  1238=>"111100111",
  1239=>"100111011",
  1240=>"011011111",
  1241=>"111100000",
  1242=>"000100010",
  1243=>"000000001",
  1244=>"110011001",
  1245=>"011000100",
  1246=>"111011000",
  1247=>"111101110",
  1248=>"000100000",
  1249=>"100100100",
  1250=>"001001001",
  1251=>"010100000",
  1252=>"000100110",
  1253=>"011111000",
  1254=>"100100111",
  1255=>"000110110",
  1256=>"000000000",
  1257=>"100011010",
  1258=>"111010111",
  1259=>"010011011",
  1260=>"000111110",
  1261=>"011011011",
  1262=>"000100000",
  1263=>"000000010",
  1264=>"001111000",
  1265=>"110011110",
  1266=>"011011111",
  1267=>"100100110",
  1268=>"001111111",
  1269=>"000000011",
  1270=>"000000000",
  1271=>"111101111",
  1272=>"001000010",
  1273=>"111011100",
  1274=>"010000000",
  1275=>"111111111",
  1276=>"100100000",
  1277=>"011000000",
  1278=>"000111011",
  1279=>"111100001",
  1280=>"101111111",
  1281=>"010010000",
  1282=>"011000101",
  1283=>"000000000",
  1284=>"000000000",
  1285=>"101101101",
  1286=>"111101101",
  1287=>"010110001",
  1288=>"011110100",
  1289=>"111000111",
  1290=>"111101101",
  1291=>"111000000",
  1292=>"000000110",
  1293=>"000011111",
  1294=>"111010010",
  1295=>"111011000",
  1296=>"000000000",
  1297=>"000101111",
  1298=>"001000111",
  1299=>"010010000",
  1300=>"101101111",
  1301=>"100111000",
  1302=>"001011010",
  1303=>"000000011",
  1304=>"101000000",
  1305=>"000111111",
  1306=>"101101000",
  1307=>"010111111",
  1308=>"010000000",
  1309=>"111110000",
  1310=>"000111111",
  1311=>"110010000",
  1312=>"010010000",
  1313=>"101010000",
  1314=>"101000111",
  1315=>"000000100",
  1316=>"000100000",
  1317=>"111110000",
  1318=>"010110010",
  1319=>"111111000",
  1320=>"111111010",
  1321=>"000001000",
  1322=>"000000110",
  1323=>"110000000",
  1324=>"111000000",
  1325=>"010101000",
  1326=>"111101101",
  1327=>"000010111",
  1328=>"101101111",
  1329=>"110001101",
  1330=>"101101000",
  1331=>"101000000",
  1332=>"011001100",
  1333=>"101101010",
  1334=>"011001111",
  1335=>"000000000",
  1336=>"001000101",
  1337=>"101101111",
  1338=>"101101000",
  1339=>"110100111",
  1340=>"000110100",
  1341=>"111110011",
  1342=>"001100000",
  1343=>"001100111",
  1344=>"011011100",
  1345=>"000100001",
  1346=>"000101001",
  1347=>"000000001",
  1348=>"011000000",
  1349=>"000001101",
  1350=>"010110000",
  1351=>"000001010",
  1352=>"011111000",
  1353=>"101001001",
  1354=>"100101000",
  1355=>"101001101",
  1356=>"000000000",
  1357=>"101000000",
  1358=>"000101101",
  1359=>"111011110",
  1360=>"000010000",
  1361=>"111010010",
  1362=>"000000000",
  1363=>"110001000",
  1364=>"000010111",
  1365=>"011010000",
  1366=>"011011011",
  1367=>"101101101",
  1368=>"011111111",
  1369=>"000001010",
  1370=>"100011001",
  1371=>"001011000",
  1372=>"101101000",
  1373=>"011001110",
  1374=>"000111111",
  1375=>"000000101",
  1376=>"000001001",
  1377=>"101111000",
  1378=>"101000111",
  1379=>"001111111",
  1380=>"000000101",
  1381=>"110011000",
  1382=>"011011000",
  1383=>"010010000",
  1384=>"001101111",
  1385=>"101101001",
  1386=>"111111101",
  1387=>"110111000",
  1388=>"111101000",
  1389=>"111101101",
  1390=>"000000100",
  1391=>"010010010",
  1392=>"000100000",
  1393=>"100101011",
  1394=>"111101001",
  1395=>"001000000",
  1396=>"001101000",
  1397=>"000001000",
  1398=>"000011110",
  1399=>"000000101",
  1400=>"000111110",
  1401=>"111011010",
  1402=>"010100110",
  1403=>"111000101",
  1404=>"100110110",
  1405=>"011110010",
  1406=>"111010101",
  1407=>"001000100",
  1408=>"010100111",
  1409=>"111111111",
  1410=>"111000101",
  1411=>"011010000",
  1412=>"001010000",
  1413=>"010111101",
  1414=>"011110100",
  1415=>"000011000",
  1416=>"101011010",
  1417=>"110101001",
  1418=>"000000100",
  1419=>"001010011",
  1420=>"000110111",
  1421=>"111001001",
  1422=>"010101111",
  1423=>"101000000",
  1424=>"011111011",
  1425=>"101101010",
  1426=>"100000100",
  1427=>"101011011",
  1428=>"000000000",
  1429=>"101100111",
  1430=>"111101111",
  1431=>"101111011",
  1432=>"111000000",
  1433=>"010010000",
  1434=>"000010010",
  1435=>"110000100",
  1436=>"101000000",
  1437=>"011010110",
  1438=>"100100110",
  1439=>"111101111",
  1440=>"010000100",
  1441=>"111110000",
  1442=>"011101101",
  1443=>"000111011",
  1444=>"110110001",
  1445=>"000110000",
  1446=>"010101011",
  1447=>"110001000",
  1448=>"011100100",
  1449=>"000011111",
  1450=>"101101000",
  1451=>"000100101",
  1452=>"011110111",
  1453=>"000000011",
  1454=>"011011001",
  1455=>"101001001",
  1456=>"010100111",
  1457=>"001111000",
  1458=>"001101101",
  1459=>"000011111",
  1460=>"111111010",
  1461=>"111100101",
  1462=>"100111011",
  1463=>"011000000",
  1464=>"001011111",
  1465=>"000010000",
  1466=>"010101000",
  1467=>"000000110",
  1468=>"110110001",
  1469=>"111111101",
  1470=>"110111111",
  1471=>"101100100",
  1472=>"110111000",
  1473=>"110000001",
  1474=>"000101010",
  1475=>"100100001",
  1476=>"111000100",
  1477=>"110001000",
  1478=>"110111100",
  1479=>"000010111",
  1480=>"111100100",
  1481=>"010010111",
  1482=>"101000101",
  1483=>"000110001",
  1484=>"000010000",
  1485=>"001011111",
  1486=>"011010111",
  1487=>"111011000",
  1488=>"110110101",
  1489=>"011000100",
  1490=>"000111111",
  1491=>"111010100",
  1492=>"000110000",
  1493=>"101100100",
  1494=>"001000101",
  1495=>"000111001",
  1496=>"110100000",
  1497=>"111100100",
  1498=>"110001000",
  1499=>"101000000",
  1500=>"000000000",
  1501=>"001000101",
  1502=>"101101111",
  1503=>"000010000",
  1504=>"010011000",
  1505=>"000101100",
  1506=>"010111000",
  1507=>"110111011",
  1508=>"000010000",
  1509=>"100010111",
  1510=>"100000100",
  1511=>"010100101",
  1512=>"110101000",
  1513=>"100000111",
  1514=>"111101100",
  1515=>"101001111",
  1516=>"010010010",
  1517=>"111110000",
  1518=>"100101010",
  1519=>"101101111",
  1520=>"011101111",
  1521=>"100100000",
  1522=>"100000010",
  1523=>"111100000",
  1524=>"000000110",
  1525=>"101000100",
  1526=>"000000111",
  1527=>"010111110",
  1528=>"010111111",
  1529=>"101101000",
  1530=>"100000110",
  1531=>"010001000",
  1532=>"000111011",
  1533=>"011000101",
  1534=>"111100100",
  1535=>"010100000",
  1536=>"011001000",
  1537=>"000010001",
  1538=>"000111000",
  1539=>"000111111",
  1540=>"101101011",
  1541=>"110101000",
  1542=>"111101011",
  1543=>"000001111",
  1544=>"111101000",
  1545=>"111111111",
  1546=>"000000000",
  1547=>"101111111",
  1548=>"101001111",
  1549=>"111110000",
  1550=>"000010011",
  1551=>"101000000",
  1552=>"000000011",
  1553=>"000000000",
  1554=>"000000111",
  1555=>"101111111",
  1556=>"000110111",
  1557=>"111110100",
  1558=>"001000001",
  1559=>"001110000",
  1560=>"000100111",
  1561=>"001010000",
  1562=>"000001000",
  1563=>"000011111",
  1564=>"000110000",
  1565=>"001000001",
  1566=>"111101000",
  1567=>"000101111",
  1568=>"000000000",
  1569=>"111111111",
  1570=>"000000110",
  1571=>"111101000",
  1572=>"100111010",
  1573=>"110111100",
  1574=>"010000000",
  1575=>"111111111",
  1576=>"000111111",
  1577=>"100100000",
  1578=>"111010000",
  1579=>"000000000",
  1580=>"111111001",
  1581=>"000111111",
  1582=>"111000000",
  1583=>"000000000",
  1584=>"111000000",
  1585=>"100110010",
  1586=>"000001010",
  1587=>"001000000",
  1588=>"000000000",
  1589=>"110010000",
  1590=>"100100100",
  1591=>"010110111",
  1592=>"111111111",
  1593=>"000010111",
  1594=>"110100100",
  1595=>"000000000",
  1596=>"110111111",
  1597=>"101111001",
  1598=>"111001100",
  1599=>"111111111",
  1600=>"001000000",
  1601=>"110001110",
  1602=>"110110110",
  1603=>"111111000",
  1604=>"111111110",
  1605=>"100000010",
  1606=>"111111111",
  1607=>"111111111",
  1608=>"111111111",
  1609=>"000000001",
  1610=>"011111011",
  1611=>"000000000",
  1612=>"111111000",
  1613=>"111001011",
  1614=>"111011110",
  1615=>"100010111",
  1616=>"000010011",
  1617=>"111111110",
  1618=>"111000101",
  1619=>"011011010",
  1620=>"000010000",
  1621=>"111110110",
  1622=>"111101100",
  1623=>"100000111",
  1624=>"111110000",
  1625=>"100100100",
  1626=>"111011010",
  1627=>"111100101",
  1628=>"010110111",
  1629=>"001001001",
  1630=>"010111111",
  1631=>"111111001",
  1632=>"111000000",
  1633=>"000001001",
  1634=>"111011000",
  1635=>"000000100",
  1636=>"000101101",
  1637=>"001101000",
  1638=>"001001001",
  1639=>"110010011",
  1640=>"011110110",
  1641=>"000100000",
  1642=>"110110111",
  1643=>"111000001",
  1644=>"011001000",
  1645=>"000000000",
  1646=>"110010001",
  1647=>"000001101",
  1648=>"101001000",
  1649=>"010000101",
  1650=>"011001000",
  1651=>"101001101",
  1652=>"000001000",
  1653=>"000000000",
  1654=>"111111111",
  1655=>"111111001",
  1656=>"000000000",
  1657=>"001100010",
  1658=>"000101000",
  1659=>"000101100",
  1660=>"000110111",
  1661=>"110100000",
  1662=>"000000000",
  1663=>"011000000",
  1664=>"101111000",
  1665=>"111101000",
  1666=>"111111000",
  1667=>"001101010",
  1668=>"111011100",
  1669=>"000011101",
  1670=>"111111011",
  1671=>"110110011",
  1672=>"001101011",
  1673=>"000000111",
  1674=>"000000000",
  1675=>"000000000",
  1676=>"111110000",
  1677=>"000000111",
  1678=>"001111111",
  1679=>"101000100",
  1680=>"001001001",
  1681=>"100110100",
  1682=>"111000111",
  1683=>"000001000",
  1684=>"101010111",
  1685=>"100010111",
  1686=>"010111011",
  1687=>"110101101",
  1688=>"111000100",
  1689=>"010000111",
  1690=>"111111000",
  1691=>"000000010",
  1692=>"001001001",
  1693=>"111110111",
  1694=>"111001111",
  1695=>"011000010",
  1696=>"110111111",
  1697=>"000000000",
  1698=>"011111000",
  1699=>"000111001",
  1700=>"010000000",
  1701=>"010010010",
  1702=>"000000000",
  1703=>"010110010",
  1704=>"011000011",
  1705=>"100100110",
  1706=>"111111000",
  1707=>"000100100",
  1708=>"001101110",
  1709=>"111011101",
  1710=>"100000000",
  1711=>"111111111",
  1712=>"101111011",
  1713=>"101001001",
  1714=>"000000100",
  1715=>"001110110",
  1716=>"100100010",
  1717=>"000000000",
  1718=>"110100000",
  1719=>"100010010",
  1720=>"011111111",
  1721=>"110111110",
  1722=>"111001001",
  1723=>"000000111",
  1724=>"000000000",
  1725=>"111111101",
  1726=>"111101000",
  1727=>"000000001",
  1728=>"000000000",
  1729=>"000000000",
  1730=>"110111101",
  1731=>"101001000",
  1732=>"000111011",
  1733=>"000111111",
  1734=>"100000011",
  1735=>"110110010",
  1736=>"111001011",
  1737=>"101111100",
  1738=>"001101000",
  1739=>"101111111",
  1740=>"011011110",
  1741=>"000011111",
  1742=>"000000000",
  1743=>"111100110",
  1744=>"110111001",
  1745=>"011001011",
  1746=>"101110111",
  1747=>"111011111",
  1748=>"110011101",
  1749=>"010100101",
  1750=>"110111001",
  1751=>"111001111",
  1752=>"000000000",
  1753=>"000001111",
  1754=>"001010010",
  1755=>"000000000",
  1756=>"011000010",
  1757=>"000101110",
  1758=>"000000010",
  1759=>"111111111",
  1760=>"001011111",
  1761=>"000000000",
  1762=>"111111111",
  1763=>"000100110",
  1764=>"010111111",
  1765=>"011110010",
  1766=>"111001000",
  1767=>"011001000",
  1768=>"011011000",
  1769=>"010000100",
  1770=>"000000000",
  1771=>"000000001",
  1772=>"101111111",
  1773=>"101000000",
  1774=>"100111000",
  1775=>"111101101",
  1776=>"001111000",
  1777=>"000111011",
  1778=>"001000011",
  1779=>"011011010",
  1780=>"110110100",
  1781=>"000000000",
  1782=>"011000001",
  1783=>"011001001",
  1784=>"111110111",
  1785=>"001011000",
  1786=>"001101101",
  1787=>"001111111",
  1788=>"000111111",
  1789=>"101000000",
  1790=>"100100111",
  1791=>"001001011",
  1792=>"110001000",
  1793=>"010001000",
  1794=>"000011011",
  1795=>"010111111",
  1796=>"111111111",
  1797=>"111010111",
  1798=>"111011000",
  1799=>"000000000",
  1800=>"000010000",
  1801=>"000010011",
  1802=>"110111110",
  1803=>"111111011",
  1804=>"000000010",
  1805=>"000100011",
  1806=>"111111100",
  1807=>"000001101",
  1808=>"000000000",
  1809=>"111000000",
  1810=>"111111000",
  1811=>"111111111",
  1812=>"111111010",
  1813=>"111000000",
  1814=>"111110011",
  1815=>"111111110",
  1816=>"010000001",
  1817=>"111111111",
  1818=>"001000010",
  1819=>"000000001",
  1820=>"100011011",
  1821=>"111101101",
  1822=>"011010110",
  1823=>"000000100",
  1824=>"110110111",
  1825=>"000000000",
  1826=>"001000001",
  1827=>"110110111",
  1828=>"001001000",
  1829=>"111010000",
  1830=>"111100111",
  1831=>"000000000",
  1832=>"111111010",
  1833=>"000000010",
  1834=>"000001101",
  1835=>"101111111",
  1836=>"001001001",
  1837=>"111111011",
  1838=>"000101001",
  1839=>"100011000",
  1840=>"000000000",
  1841=>"011111111",
  1842=>"000000111",
  1843=>"111000111",
  1844=>"000100011",
  1845=>"000000000",
  1846=>"001101001",
  1847=>"111000100",
  1848=>"111110010",
  1849=>"001100000",
  1850=>"001000000",
  1851=>"000000010",
  1852=>"001000001",
  1853=>"111100100",
  1854=>"000000110",
  1855=>"011110111",
  1856=>"110110010",
  1857=>"000001100",
  1858=>"000001000",
  1859=>"110001110",
  1860=>"000000000",
  1861=>"111000100",
  1862=>"000011010",
  1863=>"001001111",
  1864=>"000000101",
  1865=>"000000010",
  1866=>"111000100",
  1867=>"011000001",
  1868=>"100000011",
  1869=>"010111101",
  1870=>"000001100",
  1871=>"000100011",
  1872=>"100000100",
  1873=>"110000000",
  1874=>"000010001",
  1875=>"000000000",
  1876=>"000001000",
  1877=>"000000010",
  1878=>"111011011",
  1879=>"000001011",
  1880=>"111111110",
  1881=>"001010000",
  1882=>"110101111",
  1883=>"000000000",
  1884=>"000000001",
  1885=>"101100100",
  1886=>"000000000",
  1887=>"111110010",
  1888=>"000000011",
  1889=>"000000000",
  1890=>"000111001",
  1891=>"101111111",
  1892=>"101111101",
  1893=>"000001000",
  1894=>"000011111",
  1895=>"000100100",
  1896=>"001011011",
  1897=>"101000111",
  1898=>"111111010",
  1899=>"000010111",
  1900=>"111111110",
  1901=>"111111000",
  1902=>"111011001",
  1903=>"000000100",
  1904=>"100001100",
  1905=>"001101000",
  1906=>"110111010",
  1907=>"000110111",
  1908=>"000110000",
  1909=>"110010001",
  1910=>"111000000",
  1911=>"000000000",
  1912=>"000000111",
  1913=>"000000000",
  1914=>"111111111",
  1915=>"000011001",
  1916=>"111011011",
  1917=>"010010010",
  1918=>"011110000",
  1919=>"000000000",
  1920=>"000001000",
  1921=>"010110000",
  1922=>"111111111",
  1923=>"000001111",
  1924=>"000000000",
  1925=>"101000101",
  1926=>"110011111",
  1927=>"001010011",
  1928=>"011111011",
  1929=>"000001010",
  1930=>"111111111",
  1931=>"111111101",
  1932=>"000110111",
  1933=>"110001111",
  1934=>"101111111",
  1935=>"010000011",
  1936=>"111010110",
  1937=>"000110111",
  1938=>"000000000",
  1939=>"110110011",
  1940=>"111010011",
  1941=>"000011000",
  1942=>"000000000",
  1943=>"000000000",
  1944=>"000000000",
  1945=>"011011111",
  1946=>"000000000",
  1947=>"000111011",
  1948=>"111111110",
  1949=>"000000000",
  1950=>"000011101",
  1951=>"000000000",
  1952=>"001000010",
  1953=>"111110111",
  1954=>"000000000",
  1955=>"011011111",
  1956=>"110111001",
  1957=>"110010000",
  1958=>"000000000",
  1959=>"000111011",
  1960=>"111010000",
  1961=>"000000001",
  1962=>"000000000",
  1963=>"110000001",
  1964=>"111111111",
  1965=>"101010000",
  1966=>"111111000",
  1967=>"001101111",
  1968=>"001001100",
  1969=>"000000011",
  1970=>"100111111",
  1971=>"011011111",
  1972=>"111111111",
  1973=>"000000011",
  1974=>"010010000",
  1975=>"110011011",
  1976=>"000000000",
  1977=>"100100111",
  1978=>"010000000",
  1979=>"000110110",
  1980=>"111110100",
  1981=>"111111111",
  1982=>"111111100",
  1983=>"000000000",
  1984=>"000010000",
  1985=>"000100111",
  1986=>"001010010",
  1987=>"111111111",
  1988=>"000001001",
  1989=>"111110100",
  1990=>"000000001",
  1991=>"000000000",
  1992=>"111111001",
  1993=>"000000011",
  1994=>"000010010",
  1995=>"001001101",
  1996=>"000111111",
  1997=>"110111000",
  1998=>"000000000",
  1999=>"101111110",
  2000=>"100110100",
  2001=>"110111110",
  2002=>"000000001",
  2003=>"010000100",
  2004=>"000000000",
  2005=>"000000001",
  2006=>"000000000",
  2007=>"011010100",
  2008=>"010110000",
  2009=>"000000000",
  2010=>"001000100",
  2011=>"101111111",
  2012=>"000100110",
  2013=>"000000000",
  2014=>"000000000",
  2015=>"000000111",
  2016=>"100000011",
  2017=>"111111110",
  2018=>"000011010",
  2019=>"011001111",
  2020=>"000000011",
  2021=>"111111111",
  2022=>"100110101",
  2023=>"010110110",
  2024=>"111111111",
  2025=>"110100111",
  2026=>"111111111",
  2027=>"000000000",
  2028=>"000000000",
  2029=>"000000001",
  2030=>"111110000",
  2031=>"110000000",
  2032=>"100000000",
  2033=>"001001001",
  2034=>"000000000",
  2035=>"110111110",
  2036=>"000000110",
  2037=>"000000000",
  2038=>"111110110",
  2039=>"000000101",
  2040=>"000000000",
  2041=>"111100100",
  2042=>"111110111",
  2043=>"011111101",
  2044=>"111111111",
  2045=>"000001001",
  2046=>"111110100",
  2047=>"000000000",
  2048=>"001011111",
  2049=>"010000000",
  2050=>"000100000",
  2051=>"001000011",
  2052=>"100100111",
  2053=>"000111011",
  2054=>"000000000",
  2055=>"111000000",
  2056=>"000000110",
  2057=>"000000000",
  2058=>"001001000",
  2059=>"000000000",
  2060=>"000000101",
  2061=>"111111111",
  2062=>"000100100",
  2063=>"011100000",
  2064=>"101001000",
  2065=>"010000000",
  2066=>"010111100",
  2067=>"011000000",
  2068=>"000000111",
  2069=>"000000100",
  2070=>"111101000",
  2071=>"111111001",
  2072=>"000000000",
  2073=>"101011111",
  2074=>"000000111",
  2075=>"111001000",
  2076=>"111010010",
  2077=>"011001000",
  2078=>"000100111",
  2079=>"001001110",
  2080=>"011000010",
  2081=>"111000111",
  2082=>"000011111",
  2083=>"000000000",
  2084=>"000111111",
  2085=>"010111110",
  2086=>"000000111",
  2087=>"111111101",
  2088=>"100111111",
  2089=>"100000101",
  2090=>"111111000",
  2091=>"110111010",
  2092=>"000000110",
  2093=>"110001000",
  2094=>"110110111",
  2095=>"111111111",
  2096=>"000000110",
  2097=>"110100110",
  2098=>"000000010",
  2099=>"111011010",
  2100=>"010001000",
  2101=>"111001011",
  2102=>"110110100",
  2103=>"000001000",
  2104=>"011110111",
  2105=>"101001001",
  2106=>"111000000",
  2107=>"110000000",
  2108=>"000000010",
  2109=>"010001011",
  2110=>"000000010",
  2111=>"111011110",
  2112=>"000000010",
  2113=>"101111000",
  2114=>"000110110",
  2115=>"110011011",
  2116=>"111000000",
  2117=>"001001001",
  2118=>"111001001",
  2119=>"100110011",
  2120=>"010001001",
  2121=>"000110111",
  2122=>"111001001",
  2123=>"111000000",
  2124=>"000110111",
  2125=>"010100100",
  2126=>"011011111",
  2127=>"110000000",
  2128=>"001000111",
  2129=>"110111101",
  2130=>"000001001",
  2131=>"000000011",
  2132=>"001000000",
  2133=>"111110100",
  2134=>"000011011",
  2135=>"111001010",
  2136=>"011001011",
  2137=>"010100100",
  2138=>"111101000",
  2139=>"111111100",
  2140=>"000110110",
  2141=>"000000001",
  2142=>"110111111",
  2143=>"110100110",
  2144=>"000000000",
  2145=>"000000100",
  2146=>"010111001",
  2147=>"111111000",
  2148=>"101100110",
  2149=>"110101100",
  2150=>"100111110",
  2151=>"000111110",
  2152=>"011111001",
  2153=>"111110000",
  2154=>"111111001",
  2155=>"000100011",
  2156=>"000000110",
  2157=>"111000000",
  2158=>"111000101",
  2159=>"101000000",
  2160=>"100100011",
  2161=>"111011100",
  2162=>"011011000",
  2163=>"000001000",
  2164=>"001111000",
  2165=>"000000001",
  2166=>"000000000",
  2167=>"000111111",
  2168=>"101101000",
  2169=>"111100000",
  2170=>"111011011",
  2171=>"000110011",
  2172=>"000000000",
  2173=>"000000010",
  2174=>"110111111",
  2175=>"000110110",
  2176=>"111001000",
  2177=>"001000000",
  2178=>"011111111",
  2179=>"111010001",
  2180=>"101000111",
  2181=>"111111011",
  2182=>"110111111",
  2183=>"000000110",
  2184=>"011000111",
  2185=>"111000000",
  2186=>"010000000",
  2187=>"000110111",
  2188=>"000010111",
  2189=>"001000110",
  2190=>"111111110",
  2191=>"100000000",
  2192=>"111011011",
  2193=>"101101111",
  2194=>"000100000",
  2195=>"011000110",
  2196=>"000000110",
  2197=>"111001000",
  2198=>"110101000",
  2199=>"000000001",
  2200=>"111001001",
  2201=>"010111110",
  2202=>"000110110",
  2203=>"100001001",
  2204=>"111000000",
  2205=>"111110110",
  2206=>"100110000",
  2207=>"001001000",
  2208=>"100100011",
  2209=>"110001101",
  2210=>"000110111",
  2211=>"111000001",
  2212=>"000000000",
  2213=>"000001111",
  2214=>"000000110",
  2215=>"000110110",
  2216=>"111110110",
  2217=>"000000000",
  2218=>"101001000",
  2219=>"000000000",
  2220=>"111111010",
  2221=>"000010111",
  2222=>"011101101",
  2223=>"011111011",
  2224=>"010110101",
  2225=>"000001011",
  2226=>"000101000",
  2227=>"000011010",
  2228=>"000110111",
  2229=>"111101000",
  2230=>"010111111",
  2231=>"101010110",
  2232=>"000000010",
  2233=>"000000011",
  2234=>"001010111",
  2235=>"111001001",
  2236=>"100111010",
  2237=>"000110111",
  2238=>"001011001",
  2239=>"110001000",
  2240=>"000101101",
  2241=>"001001000",
  2242=>"001001001",
  2243=>"000000011",
  2244=>"111110111",
  2245=>"000000001",
  2246=>"110100000",
  2247=>"011000000",
  2248=>"110001010",
  2249=>"111101111",
  2250=>"000000011",
  2251=>"111001000",
  2252=>"100110110",
  2253=>"000000011",
  2254=>"111101001",
  2255=>"111011000",
  2256=>"010000001",
  2257=>"000000000",
  2258=>"111000011",
  2259=>"010000000",
  2260=>"000000011",
  2261=>"001001100",
  2262=>"000000100",
  2263=>"000001001",
  2264=>"111111001",
  2265=>"000000000",
  2266=>"111001000",
  2267=>"010000001",
  2268=>"111011011",
  2269=>"100001111",
  2270=>"111111010",
  2271=>"101001100",
  2272=>"111000100",
  2273=>"011111110",
  2274=>"111001001",
  2275=>"000000001",
  2276=>"000000000",
  2277=>"111001001",
  2278=>"000000010",
  2279=>"001101001",
  2280=>"000000010",
  2281=>"000001101",
  2282=>"100001000",
  2283=>"000111111",
  2284=>"000000111",
  2285=>"110001001",
  2286=>"000000100",
  2287=>"000000001",
  2288=>"000000000",
  2289=>"001010011",
  2290=>"111001101",
  2291=>"111011111",
  2292=>"100100111",
  2293=>"111100000",
  2294=>"000000010",
  2295=>"111111110",
  2296=>"111111001",
  2297=>"110111111",
  2298=>"111000000",
  2299=>"000000111",
  2300=>"111000000",
  2301=>"100000110",
  2302=>"011001001",
  2303=>"111101001",
  2304=>"001100111",
  2305=>"100000010",
  2306=>"000010111",
  2307=>"111111000",
  2308=>"100100110",
  2309=>"110111101",
  2310=>"101011000",
  2311=>"111101111",
  2312=>"101101111",
  2313=>"100100101",
  2314=>"000111100",
  2315=>"111100101",
  2316=>"101100000",
  2317=>"101000000",
  2318=>"000101101",
  2319=>"011110000",
  2320=>"111101000",
  2321=>"010000000",
  2322=>"111101000",
  2323=>"101111100",
  2324=>"000110111",
  2325=>"101100111",
  2326=>"110011001",
  2327=>"000110111",
  2328=>"000101100",
  2329=>"010000010",
  2330=>"111111101",
  2331=>"011011110",
  2332=>"101001111",
  2333=>"111111010",
  2334=>"101100111",
  2335=>"111000000",
  2336=>"101110001",
  2337=>"010101111",
  2338=>"000011101",
  2339=>"000000111",
  2340=>"110100001",
  2341=>"100100110",
  2342=>"000111110",
  2343=>"100100101",
  2344=>"111101001",
  2345=>"011111111",
  2346=>"111111110",
  2347=>"010000010",
  2348=>"110110110",
  2349=>"111100111",
  2350=>"100011111",
  2351=>"000100101",
  2352=>"000000100",
  2353=>"001000000",
  2354=>"000100101",
  2355=>"000000000",
  2356=>"101011101",
  2357=>"101001001",
  2358=>"000001100",
  2359=>"000001101",
  2360=>"111111101",
  2361=>"101101100",
  2362=>"011111000",
  2363=>"000000001",
  2364=>"100100101",
  2365=>"111111101",
  2366=>"001000000",
  2367=>"001000100",
  2368=>"101101111",
  2369=>"110100100",
  2370=>"100001000",
  2371=>"111101111",
  2372=>"011111000",
  2373=>"000111001",
  2374=>"101111101",
  2375=>"111110010",
  2376=>"100100111",
  2377=>"111010111",
  2378=>"111101110",
  2379=>"101101000",
  2380=>"100101101",
  2381=>"111100100",
  2382=>"011101000",
  2383=>"000000100",
  2384=>"000000000",
  2385=>"011000000",
  2386=>"011111111",
  2387=>"001000011",
  2388=>"000100101",
  2389=>"100101110",
  2390=>"111100000",
  2391=>"000101111",
  2392=>"000000011",
  2393=>"011001000",
  2394=>"011011011",
  2395=>"001001000",
  2396=>"001101101",
  2397=>"010110000",
  2398=>"101101111",
  2399=>"111101111",
  2400=>"010000110",
  2401=>"110111111",
  2402=>"100101101",
  2403=>"110110110",
  2404=>"001001000",
  2405=>"011000000",
  2406=>"101000011",
  2407=>"000000010",
  2408=>"010111011",
  2409=>"000000101",
  2410=>"110111101",
  2411=>"100100101",
  2412=>"000010110",
  2413=>"100101000",
  2414=>"100101001",
  2415=>"010111111",
  2416=>"100100100",
  2417=>"000101101",
  2418=>"000000001",
  2419=>"100101101",
  2420=>"000111010",
  2421=>"010101110",
  2422=>"100100000",
  2423=>"001000000",
  2424=>"111111111",
  2425=>"010010110",
  2426=>"111111101",
  2427=>"101100101",
  2428=>"001000000",
  2429=>"000101110",
  2430=>"110010010",
  2431=>"111000000",
  2432=>"111101100",
  2433=>"000000011",
  2434=>"000100111",
  2435=>"111111010",
  2436=>"111101111",
  2437=>"111010110",
  2438=>"001001101",
  2439=>"010000001",
  2440=>"000000100",
  2441=>"011010010",
  2442=>"101111011",
  2443=>"000100110",
  2444=>"001000001",
  2445=>"111111000",
  2446=>"011101111",
  2447=>"110111111",
  2448=>"011101000",
  2449=>"111000101",
  2450=>"000000000",
  2451=>"000101001",
  2452=>"111101011",
  2453=>"101101100",
  2454=>"101101001",
  2455=>"100100001",
  2456=>"111000101",
  2457=>"011000001",
  2458=>"111111001",
  2459=>"111011010",
  2460=>"101100000",
  2461=>"111101001",
  2462=>"101100001",
  2463=>"110010010",
  2464=>"001101101",
  2465=>"101111111",
  2466=>"010010010",
  2467=>"000101011",
  2468=>"011111011",
  2469=>"100001100",
  2470=>"100000100",
  2471=>"000000111",
  2472=>"000100000",
  2473=>"001010000",
  2474=>"000111111",
  2475=>"000010111",
  2476=>"100011010",
  2477=>"010000000",
  2478=>"110010110",
  2479=>"111000000",
  2480=>"111000110",
  2481=>"000100000",
  2482=>"000101000",
  2483=>"010100000",
  2484=>"001001111",
  2485=>"111010000",
  2486=>"100001000",
  2487=>"110111100",
  2488=>"001001100",
  2489=>"101100100",
  2490=>"100000000",
  2491=>"010110010",
  2492=>"000011011",
  2493=>"101101111",
  2494=>"111101001",
  2495=>"000000000",
  2496=>"100100001",
  2497=>"010000000",
  2498=>"101001101",
  2499=>"001001101",
  2500=>"000100000",
  2501=>"100100100",
  2502=>"111111011",
  2503=>"001001101",
  2504=>"111000001",
  2505=>"101010010",
  2506=>"110010001",
  2507=>"100101001",
  2508=>"011100100",
  2509=>"100000000",
  2510=>"010010101",
  2511=>"000000001",
  2512=>"101101001",
  2513=>"011001100",
  2514=>"000100011",
  2515=>"111111010",
  2516=>"101000100",
  2517=>"000010110",
  2518=>"001111011",
  2519=>"000011111",
  2520=>"110000000",
  2521=>"101100100",
  2522=>"101100011",
  2523=>"100101100",
  2524=>"010010011",
  2525=>"101100000",
  2526=>"000000000",
  2527=>"101101101",
  2528=>"000000101",
  2529=>"111101001",
  2530=>"111100000",
  2531=>"111100111",
  2532=>"000000000",
  2533=>"001101111",
  2534=>"111111000",
  2535=>"110110010",
  2536=>"011101101",
  2537=>"011011111",
  2538=>"010010000",
  2539=>"000010000",
  2540=>"000100111",
  2541=>"000111111",
  2542=>"001101101",
  2543=>"000001110",
  2544=>"111011110",
  2545=>"001001101",
  2546=>"101101100",
  2547=>"110100100",
  2548=>"110001111",
  2549=>"010110110",
  2550=>"000100100",
  2551=>"000010111",
  2552=>"000101001",
  2553=>"010010011",
  2554=>"000111011",
  2555=>"111000000",
  2556=>"000000111",
  2557=>"100111101",
  2558=>"000001001",
  2559=>"101100000",
  2560=>"011001100",
  2561=>"000000000",
  2562=>"101000111",
  2563=>"011110111",
  2564=>"100001001",
  2565=>"110101111",
  2566=>"000000110",
  2567=>"001000000",
  2568=>"111111101",
  2569=>"010000110",
  2570=>"100000100",
  2571=>"000001000",
  2572=>"110111011",
  2573=>"111100000",
  2574=>"010110100",
  2575=>"000000011",
  2576=>"101111001",
  2577=>"111100111",
  2578=>"111101011",
  2579=>"000000000",
  2580=>"011010100",
  2581=>"111110000",
  2582=>"100000000",
  2583=>"101101110",
  2584=>"000000111",
  2585=>"000110000",
  2586=>"000000001",
  2587=>"011000101",
  2588=>"111101111",
  2589=>"001000010",
  2590=>"001011000",
  2591=>"111000000",
  2592=>"001001001",
  2593=>"000010110",
  2594=>"011101110",
  2595=>"001001111",
  2596=>"001001001",
  2597=>"001000111",
  2598=>"001000000",
  2599=>"000010110",
  2600=>"111110000",
  2601=>"111010001",
  2602=>"100101100",
  2603=>"110111010",
  2604=>"000100111",
  2605=>"010111010",
  2606=>"111000000",
  2607=>"110111111",
  2608=>"101001011",
  2609=>"101001000",
  2610=>"111111111",
  2611=>"101000101",
  2612=>"001001001",
  2613=>"101110101",
  2614=>"000000101",
  2615=>"010000100",
  2616=>"110000000",
  2617=>"000000101",
  2618=>"000000000",
  2619=>"101101100",
  2620=>"010000000",
  2621=>"000000000",
  2622=>"000000001",
  2623=>"010000000",
  2624=>"111111111",
  2625=>"000000000",
  2626=>"010010100",
  2627=>"111111110",
  2628=>"111110000",
  2629=>"111110000",
  2630=>"000101111",
  2631=>"100000000",
  2632=>"001110000",
  2633=>"111110101",
  2634=>"000001111",
  2635=>"110000111",
  2636=>"000000101",
  2637=>"000100100",
  2638=>"011011000",
  2639=>"000000111",
  2640=>"010000000",
  2641=>"001001001",
  2642=>"000111100",
  2643=>"010000010",
  2644=>"000000000",
  2645=>"100101110",
  2646=>"011100010",
  2647=>"000110111",
  2648=>"100001000",
  2649=>"100100101",
  2650=>"001000000",
  2651=>"001111111",
  2652=>"000000000",
  2653=>"000000000",
  2654=>"111111111",
  2655=>"111011011",
  2656=>"010000000",
  2657=>"110010110",
  2658=>"001001001",
  2659=>"100000000",
  2660=>"010011011",
  2661=>"000000100",
  2662=>"000000111",
  2663=>"111111000",
  2664=>"100111111",
  2665=>"110010000",
  2666=>"000000101",
  2667=>"110001101",
  2668=>"110110000",
  2669=>"001001101",
  2670=>"000000111",
  2671=>"000000000",
  2672=>"110100100",
  2673=>"001010010",
  2674=>"000100000",
  2675=>"110011101",
  2676=>"111110000",
  2677=>"010001111",
  2678=>"111000000",
  2679=>"010010000",
  2680=>"111000111",
  2681=>"000000111",
  2682=>"001010000",
  2683=>"111111010",
  2684=>"100000100",
  2685=>"000000000",
  2686=>"111111101",
  2687=>"011000000",
  2688=>"100000000",
  2689=>"000000001",
  2690=>"001000000",
  2691=>"111000111",
  2692=>"000000110",
  2693=>"111100000",
  2694=>"000000100",
  2695=>"000001000",
  2696=>"001011000",
  2697=>"111000000",
  2698=>"000000111",
  2699=>"010010000",
  2700=>"110110000",
  2701=>"111001100",
  2702=>"011111101",
  2703=>"000100101",
  2704=>"100100000",
  2705=>"000000000",
  2706=>"000101101",
  2707=>"101000000",
  2708=>"000010111",
  2709=>"011010010",
  2710=>"001101111",
  2711=>"111011111",
  2712=>"000001000",
  2713=>"000000101",
  2714=>"011010111",
  2715=>"000010010",
  2716=>"100100100",
  2717=>"010011000",
  2718=>"000000111",
  2719=>"101001111",
  2720=>"101001010",
  2721=>"101010101",
  2722=>"111111110",
  2723=>"000000111",
  2724=>"000000000",
  2725=>"111000000",
  2726=>"111110000",
  2727=>"111101101",
  2728=>"001000100",
  2729=>"010001000",
  2730=>"101011111",
  2731=>"110000000",
  2732=>"111000110",
  2733=>"010010001",
  2734=>"100000101",
  2735=>"111111010",
  2736=>"100110111",
  2737=>"010110100",
  2738=>"000010000",
  2739=>"000110111",
  2740=>"111011011",
  2741=>"111111010",
  2742=>"111111111",
  2743=>"111111000",
  2744=>"101000100",
  2745=>"000101111",
  2746=>"010101001",
  2747=>"000010010",
  2748=>"111111111",
  2749=>"010110000",
  2750=>"111100100",
  2751=>"011010001",
  2752=>"101000010",
  2753=>"010010000",
  2754=>"010111000",
  2755=>"001000000",
  2756=>"000000100",
  2757=>"001001100",
  2758=>"000011011",
  2759=>"000100111",
  2760=>"101001100",
  2761=>"010000101",
  2762=>"111111111",
  2763=>"011001000",
  2764=>"000010000",
  2765=>"000000001",
  2766=>"111100100",
  2767=>"111101111",
  2768=>"000101111",
  2769=>"110110100",
  2770=>"101111111",
  2771=>"000000011",
  2772=>"000000000",
  2773=>"000110000",
  2774=>"000000100",
  2775=>"000011000",
  2776=>"000101000",
  2777=>"100111011",
  2778=>"001011001",
  2779=>"000000110",
  2780=>"011000101",
  2781=>"110010011",
  2782=>"010100111",
  2783=>"111000010",
  2784=>"111000101",
  2785=>"110010101",
  2786=>"000000110",
  2787=>"101111111",
  2788=>"011110111",
  2789=>"010110000",
  2790=>"100100000",
  2791=>"000011011",
  2792=>"111111110",
  2793=>"010000111",
  2794=>"101000001",
  2795=>"110110100",
  2796=>"111111101",
  2797=>"110000101",
  2798=>"000000000",
  2799=>"010000000",
  2800=>"111001000",
  2801=>"100100000",
  2802=>"011101111",
  2803=>"000100010",
  2804=>"110110011",
  2805=>"000000100",
  2806=>"000000010",
  2807=>"001111111",
  2808=>"000001111",
  2809=>"111110110",
  2810=>"101111001",
  2811=>"101111011",
  2812=>"100111111",
  2813=>"111110000",
  2814=>"000100000",
  2815=>"000001111",
  2816=>"101101101",
  2817=>"000000001",
  2818=>"001001111",
  2819=>"101010000",
  2820=>"100100111",
  2821=>"010010110",
  2822=>"001101101",
  2823=>"000010101",
  2824=>"010010000",
  2825=>"011111001",
  2826=>"100000001",
  2827=>"000011111",
  2828=>"001101111",
  2829=>"111111000",
  2830=>"000000100",
  2831=>"101000000",
  2832=>"000010000",
  2833=>"111010010",
  2834=>"011100000",
  2835=>"110100000",
  2836=>"111111111",
  2837=>"000110100",
  2838=>"011001000",
  2839=>"000011101",
  2840=>"010000000",
  2841=>"111000000",
  2842=>"111000000",
  2843=>"011000000",
  2844=>"000001111",
  2845=>"111001001",
  2846=>"010001000",
  2847=>"111001000",
  2848=>"110110000",
  2849=>"010000101",
  2850=>"111111111",
  2851=>"000111011",
  2852=>"110111100",
  2853=>"011101101",
  2854=>"011000000",
  2855=>"001111111",
  2856=>"110011001",
  2857=>"010001000",
  2858=>"000011011",
  2859=>"111111010",
  2860=>"101100101",
  2861=>"010110001",
  2862=>"111111011",
  2863=>"100010100",
  2864=>"010001100",
  2865=>"011001111",
  2866=>"111111100",
  2867=>"000101000",
  2868=>"000000101",
  2869=>"100001111",
  2870=>"001101111",
  2871=>"010011000",
  2872=>"100010011",
  2873=>"000000011",
  2874=>"000000000",
  2875=>"111111000",
  2876=>"000101011",
  2877=>"011001001",
  2878=>"101111111",
  2879=>"011011000",
  2880=>"111000000",
  2881=>"101111011",
  2882=>"000000001",
  2883=>"011001001",
  2884=>"000001001",
  2885=>"010011111",
  2886=>"101111000",
  2887=>"001111100",
  2888=>"001111011",
  2889=>"110100000",
  2890=>"101000100",
  2891=>"110011000",
  2892=>"111111000",
  2893=>"101100001",
  2894=>"110110011",
  2895=>"000001011",
  2896=>"000101111",
  2897=>"111111110",
  2898=>"010111001",
  2899=>"011001000",
  2900=>"101001000",
  2901=>"111110101",
  2902=>"011011001",
  2903=>"001111111",
  2904=>"000100111",
  2905=>"101111001",
  2906=>"011010011",
  2907=>"011010001",
  2908=>"000000100",
  2909=>"000000100",
  2910=>"111111000",
  2911=>"110000000",
  2912=>"000000101",
  2913=>"010000001",
  2914=>"001000111",
  2915=>"111111110",
  2916=>"100101011",
  2917=>"100010010",
  2918=>"110110000",
  2919=>"110000000",
  2920=>"110000000",
  2921=>"000000000",
  2922=>"101111101",
  2923=>"000001001",
  2924=>"111111000",
  2925=>"001100110",
  2926=>"000000000",
  2927=>"001111010",
  2928=>"100100000",
  2929=>"001000111",
  2930=>"001100111",
  2931=>"000101111",
  2932=>"111010000",
  2933=>"000000000",
  2934=>"000100111",
  2935=>"001100000",
  2936=>"000000100",
  2937=>"111110010",
  2938=>"110110111",
  2939=>"111111101",
  2940=>"101000000",
  2941=>"110000100",
  2942=>"110110010",
  2943=>"111000000",
  2944=>"110101000",
  2945=>"101101011",
  2946=>"010010000",
  2947=>"001111011",
  2948=>"110001010",
  2949=>"111111000",
  2950=>"000011011",
  2951=>"001000111",
  2952=>"011011000",
  2953=>"111101111",
  2954=>"000010000",
  2955=>"101111110",
  2956=>"010000000",
  2957=>"100010010",
  2958=>"110110000",
  2959=>"000001100",
  2960=>"011011010",
  2961=>"111100111",
  2962=>"110000000",
  2963=>"101000000",
  2964=>"001001100",
  2965=>"000000011",
  2966=>"000101111",
  2967=>"001011000",
  2968=>"001001101",
  2969=>"010111111",
  2970=>"101100101",
  2971=>"110000000",
  2972=>"000000000",
  2973=>"010000000",
  2974=>"000110111",
  2975=>"000101111",
  2976=>"001001011",
  2977=>"111111111",
  2978=>"101000100",
  2979=>"001101001",
  2980=>"010000000",
  2981=>"100100110",
  2982=>"111111001",
  2983=>"000000111",
  2984=>"001111111",
  2985=>"000010001",
  2986=>"000000110",
  2987=>"100000010",
  2988=>"000000011",
  2989=>"110111111",
  2990=>"100101111",
  2991=>"111111010",
  2992=>"111011000",
  2993=>"000001010",
  2994=>"111111101",
  2995=>"100000001",
  2996=>"110100000",
  2997=>"001000100",
  2998=>"001111011",
  2999=>"000001011",
  3000=>"010100111",
  3001=>"100001101",
  3002=>"001010100",
  3003=>"110010100",
  3004=>"110101011",
  3005=>"111110000",
  3006=>"110110001",
  3007=>"000000111",
  3008=>"000100110",
  3009=>"000000000",
  3010=>"111111101",
  3011=>"100110111",
  3012=>"000101100",
  3013=>"100010011",
  3014=>"001010111",
  3015=>"000110000",
  3016=>"000111011",
  3017=>"000110011",
  3018=>"111111101",
  3019=>"011000000",
  3020=>"011010000",
  3021=>"001100000",
  3022=>"110111111",
  3023=>"111010000",
  3024=>"011110000",
  3025=>"111110010",
  3026=>"101111011",
  3027=>"110000000",
  3028=>"010000000",
  3029=>"000000000",
  3030=>"000001111",
  3031=>"111011000",
  3032=>"000101111",
  3033=>"001111100",
  3034=>"110110100",
  3035=>"001100111",
  3036=>"110011001",
  3037=>"000111101",
  3038=>"000000000",
  3039=>"110000001",
  3040=>"001101101",
  3041=>"001111111",
  3042=>"000101111",
  3043=>"100111111",
  3044=>"000000000",
  3045=>"101111000",
  3046=>"111000001",
  3047=>"010111011",
  3048=>"011000001",
  3049=>"000000110",
  3050=>"001100100",
  3051=>"000001010",
  3052=>"000000111",
  3053=>"010110010",
  3054=>"000001011",
  3055=>"011011000",
  3056=>"110110000",
  3057=>"001101100",
  3058=>"001111001",
  3059=>"110000000",
  3060=>"001110010",
  3061=>"000000111",
  3062=>"000000111",
  3063=>"000000000",
  3064=>"000110111",
  3065=>"001111000",
  3066=>"111110000",
  3067=>"001000010",
  3068=>"000101011",
  3069=>"000000000",
  3070=>"011111100",
  3071=>"101101111",
  3072=>"101100100",
  3073=>"111011110",
  3074=>"100100110",
  3075=>"010011000",
  3076=>"011110001",
  3077=>"011011000",
  3078=>"100110111",
  3079=>"100100100",
  3080=>"011011001",
  3081=>"100100000",
  3082=>"100100110",
  3083=>"000000001",
  3084=>"100110111",
  3085=>"011001001",
  3086=>"110110110",
  3087=>"100100100",
  3088=>"001010001",
  3089=>"100110111",
  3090=>"110110110",
  3091=>"010000000",
  3092=>"110110011",
  3093=>"001011000",
  3094=>"111001111",
  3095=>"000110010",
  3096=>"100100111",
  3097=>"001000110",
  3098=>"011011001",
  3099=>"000010110",
  3100=>"100111111",
  3101=>"110110111",
  3102=>"001110110",
  3103=>"111011001",
  3104=>"011000000",
  3105=>"011111100",
  3106=>"110111000",
  3107=>"011001000",
  3108=>"100100010",
  3109=>"000011001",
  3110=>"011011000",
  3111=>"000100100",
  3112=>"001000000",
  3113=>"011011011",
  3114=>"000000110",
  3115=>"111100001",
  3116=>"011110111",
  3117=>"110111111",
  3118=>"011111101",
  3119=>"000100100",
  3120=>"110111000",
  3121=>"000000000",
  3122=>"111011001",
  3123=>"110100100",
  3124=>"100100111",
  3125=>"000000100",
  3126=>"001100110",
  3127=>"100100011",
  3128=>"011101111",
  3129=>"100100111",
  3130=>"000000000",
  3131=>"110111100",
  3132=>"001001000",
  3133=>"111111010",
  3134=>"100100110",
  3135=>"001001000",
  3136=>"100000111",
  3137=>"000111101",
  3138=>"011001001",
  3139=>"101101000",
  3140=>"011011000",
  3141=>"111011000",
  3142=>"100110011",
  3143=>"000000110",
  3144=>"011011011",
  3145=>"110000111",
  3146=>"100110111",
  3147=>"100100111",
  3148=>"001011011",
  3149=>"110111101",
  3150=>"001001010",
  3151=>"110111110",
  3152=>"100100110",
  3153=>"110111000",
  3154=>"011100011",
  3155=>"000000000",
  3156=>"100100100",
  3157=>"010100111",
  3158=>"001000000",
  3159=>"100100111",
  3160=>"111111011",
  3161=>"011111011",
  3162=>"111110110",
  3163=>"001101100",
  3164=>"000000000",
  3165=>"100100000",
  3166=>"001101111",
  3167=>"000010010",
  3168=>"011011000",
  3169=>"001011101",
  3170=>"100110010",
  3171=>"100110011",
  3172=>"011001100",
  3173=>"110110101",
  3174=>"011100110",
  3175=>"100100110",
  3176=>"011011000",
  3177=>"011110100",
  3178=>"001110011",
  3179=>"011110000",
  3180=>"001011100",
  3181=>"000000101",
  3182=>"000000001",
  3183=>"101011011",
  3184=>"110101100",
  3185=>"000101001",
  3186=>"100010011",
  3187=>"001000000",
  3188=>"011111000",
  3189=>"100100011",
  3190=>"011001011",
  3191=>"101111110",
  3192=>"000001011",
  3193=>"011011011",
  3194=>"110111000",
  3195=>"011110011",
  3196=>"011001001",
  3197=>"011011001",
  3198=>"110100100",
  3199=>"100010011",
  3200=>"011111010",
  3201=>"110110010",
  3202=>"001000000",
  3203=>"011000111",
  3204=>"100101000",
  3205=>"000100001",
  3206=>"101001101",
  3207=>"000100100",
  3208=>"111010010",
  3209=>"100100101",
  3210=>"100100100",
  3211=>"000100100",
  3212=>"011011000",
  3213=>"000100111",
  3214=>"000110100",
  3215=>"100100010",
  3216=>"111110000",
  3217=>"010111110",
  3218=>"000111111",
  3219=>"110110000",
  3220=>"010011000",
  3221=>"101101111",
  3222=>"100100111",
  3223=>"011001000",
  3224=>"001101110",
  3225=>"110001000",
  3226=>"100110111",
  3227=>"000100111",
  3228=>"110110000",
  3229=>"000100111",
  3230=>"000100100",
  3231=>"100110111",
  3232=>"000011111",
  3233=>"100001001",
  3234=>"000110110",
  3235=>"100101111",
  3236=>"011010000",
  3237=>"001011010",
  3238=>"111001001",
  3239=>"011110100",
  3240=>"000110111",
  3241=>"011001001",
  3242=>"011011001",
  3243=>"111110110",
  3244=>"011000000",
  3245=>"001011011",
  3246=>"000110110",
  3247=>"111010111",
  3248=>"111111111",
  3249=>"100100000",
  3250=>"000111001",
  3251=>"000000000",
  3252=>"011001010",
  3253=>"111001001",
  3254=>"011010000",
  3255=>"001100100",
  3256=>"100100011",
  3257=>"111000010",
  3258=>"011000000",
  3259=>"010001101",
  3260=>"010100100",
  3261=>"011011011",
  3262=>"011011001",
  3263=>"110110011",
  3264=>"100100111",
  3265=>"100110110",
  3266=>"000001101",
  3267=>"110100110",
  3268=>"100100110",
  3269=>"110000001",
  3270=>"100010010",
  3271=>"001001001",
  3272=>"101000000",
  3273=>"111000000",
  3274=>"101100011",
  3275=>"111001001",
  3276=>"100110111",
  3277=>"000000110",
  3278=>"100110110",
  3279=>"011001001",
  3280=>"100100100",
  3281=>"111111101",
  3282=>"100110011",
  3283=>"011011011",
  3284=>"000100111",
  3285=>"011011001",
  3286=>"111110110",
  3287=>"100001111",
  3288=>"100110111",
  3289=>"000000001",
  3290=>"111111001",
  3291=>"100100111",
  3292=>"110110010",
  3293=>"011001001",
  3294=>"011001001",
  3295=>"111111111",
  3296=>"000001011",
  3297=>"100100111",
  3298=>"010100101",
  3299=>"011000000",
  3300=>"000000000",
  3301=>"000110011",
  3302=>"001001001",
  3303=>"000010111",
  3304=>"001000001",
  3305=>"011101101",
  3306=>"100000011",
  3307=>"011011000",
  3308=>"001001000",
  3309=>"001001001",
  3310=>"010111000",
  3311=>"000011000",
  3312=>"011011000",
  3313=>"110110111",
  3314=>"001111010",
  3315=>"111100111",
  3316=>"011011011",
  3317=>"110111110",
  3318=>"100000000",
  3319=>"000001101",
  3320=>"100100111",
  3321=>"110110000",
  3322=>"110110000",
  3323=>"110000000",
  3324=>"100011111",
  3325=>"100100110",
  3326=>"000010000",
  3327=>"100100111",
  3328=>"010100100",
  3329=>"000000011",
  3330=>"101101001",
  3331=>"100110111",
  3332=>"000000010",
  3333=>"000000010",
  3334=>"110000010",
  3335=>"000111111",
  3336=>"000110110",
  3337=>"000010110",
  3338=>"010010000",
  3339=>"001000000",
  3340=>"000000110",
  3341=>"000000000",
  3342=>"011011101",
  3343=>"001110111",
  3344=>"000000110",
  3345=>"000000000",
  3346=>"100001001",
  3347=>"110111000",
  3348=>"111111110",
  3349=>"000000011",
  3350=>"111111111",
  3351=>"101110100",
  3352=>"001010001",
  3353=>"000000000",
  3354=>"100101101",
  3355=>"101101111",
  3356=>"101000011",
  3357=>"000001111",
  3358=>"110000100",
  3359=>"000000101",
  3360=>"000000000",
  3361=>"000101110",
  3362=>"000101111",
  3363=>"011110111",
  3364=>"010110000",
  3365=>"111000101",
  3366=>"000010000",
  3367=>"111000000",
  3368=>"001111111",
  3369=>"000010111",
  3370=>"000000000",
  3371=>"111100111",
  3372=>"011011000",
  3373=>"000110111",
  3374=>"110000000",
  3375=>"001001111",
  3376=>"010001000",
  3377=>"001011011",
  3378=>"111111111",
  3379=>"000100101",
  3380=>"110000000",
  3381=>"111110000",
  3382=>"110000000",
  3383=>"000000011",
  3384=>"111111111",
  3385=>"111000000",
  3386=>"000000000",
  3387=>"101111111",
  3388=>"110111000",
  3389=>"111111110",
  3390=>"101000001",
  3391=>"111100100",
  3392=>"001001101",
  3393=>"111011111",
  3394=>"001111010",
  3395=>"011100010",
  3396=>"111011000",
  3397=>"000000110",
  3398=>"110000000",
  3399=>"101000000",
  3400=>"001001011",
  3401=>"111000000",
  3402=>"000001010",
  3403=>"011110010",
  3404=>"010001001",
  3405=>"001011000",
  3406=>"100110010",
  3407=>"110111110",
  3408=>"010001001",
  3409=>"110001011",
  3410=>"010111000",
  3411=>"101100000",
  3412=>"111000101",
  3413=>"000001000",
  3414=>"110111100",
  3415=>"111000001",
  3416=>"001000000",
  3417=>"011011010",
  3418=>"110111110",
  3419=>"011001110",
  3420=>"000000011",
  3421=>"000001011",
  3422=>"111000010",
  3423=>"101001011",
  3424=>"010111110",
  3425=>"100001111",
  3426=>"011010000",
  3427=>"000001111",
  3428=>"100111000",
  3429=>"000100110",
  3430=>"111001110",
  3431=>"010000111",
  3432=>"001000000",
  3433=>"010000000",
  3434=>"111000111",
  3435=>"001000000",
  3436=>"010001111",
  3437=>"111010010",
  3438=>"000000011",
  3439=>"011011111",
  3440=>"111111001",
  3441=>"001111111",
  3442=>"011000000",
  3443=>"000000000",
  3444=>"101111111",
  3445=>"001101000",
  3446=>"100000010",
  3447=>"011001111",
  3448=>"001000000",
  3449=>"101111111",
  3450=>"111100000",
  3451=>"010010111",
  3452=>"100110010",
  3453=>"100000100",
  3454=>"000100111",
  3455=>"000000101",
  3456=>"111000111",
  3457=>"000000110",
  3458=>"110010000",
  3459=>"101011111",
  3460=>"000000001",
  3461=>"111101111",
  3462=>"110000111",
  3463=>"000011010",
  3464=>"011101110",
  3465=>"111011111",
  3466=>"000000010",
  3467=>"011000110",
  3468=>"000001111",
  3469=>"110100001",
  3470=>"101101110",
  3471=>"001001110",
  3472=>"110100100",
  3473=>"111101101",
  3474=>"000010000",
  3475=>"000001101",
  3476=>"111111001",
  3477=>"111111001",
  3478=>"111110011",
  3479=>"000000011",
  3480=>"111000000",
  3481=>"001111111",
  3482=>"111111000",
  3483=>"001000011",
  3484=>"111111011",
  3485=>"111101100",
  3486=>"011101101",
  3487=>"001001000",
  3488=>"101101010",
  3489=>"111000101",
  3490=>"101001100",
  3491=>"000000001",
  3492=>"111101000",
  3493=>"111001000",
  3494=>"100111111",
  3495=>"001101000",
  3496=>"101101111",
  3497=>"000101101",
  3498=>"100111111",
  3499=>"100111000",
  3500=>"000010011",
  3501=>"110111101",
  3502=>"111111111",
  3503=>"010001111",
  3504=>"111000000",
  3505=>"001100001",
  3506=>"101001101",
  3507=>"000100111",
  3508=>"100110010",
  3509=>"000101110",
  3510=>"000000000",
  3511=>"011010000",
  3512=>"001111100",
  3513=>"100110011",
  3514=>"010110000",
  3515=>"111111001",
  3516=>"010000010",
  3517=>"001000000",
  3518=>"100111001",
  3519=>"000100001",
  3520=>"110000000",
  3521=>"000001101",
  3522=>"111000000",
  3523=>"111110010",
  3524=>"111011010",
  3525=>"101101010",
  3526=>"010000000",
  3527=>"000000000",
  3528=>"100111110",
  3529=>"001001111",
  3530=>"000010000",
  3531=>"111000101",
  3532=>"011001001",
  3533=>"011011010",
  3534=>"111111111",
  3535=>"000101111",
  3536=>"111110000",
  3537=>"011000110",
  3538=>"000010111",
  3539=>"000111111",
  3540=>"011000000",
  3541=>"000000100",
  3542=>"111011010",
  3543=>"001011111",
  3544=>"000111110",
  3545=>"100000101",
  3546=>"111100000",
  3547=>"000000101",
  3548=>"101000110",
  3549=>"010111111",
  3550=>"000101111",
  3551=>"000000100",
  3552=>"000000101",
  3553=>"111110000",
  3554=>"000000111",
  3555=>"100110111",
  3556=>"000000001",
  3557=>"000001111",
  3558=>"111110000",
  3559=>"000101111",
  3560=>"110010000",
  3561=>"000000000",
  3562=>"101001000",
  3563=>"001101000",
  3564=>"000000110",
  3565=>"000000000",
  3566=>"000000000",
  3567=>"001001011",
  3568=>"000111101",
  3569=>"101010010",
  3570=>"110010000",
  3571=>"011101110",
  3572=>"010001011",
  3573=>"000001011",
  3574=>"000010101",
  3575=>"000100100",
  3576=>"010010000",
  3577=>"110001111",
  3578=>"101101111",
  3579=>"001111111",
  3580=>"111010111",
  3581=>"100100111",
  3582=>"111000010",
  3583=>"111000010",
  3584=>"010010011",
  3585=>"000011001",
  3586=>"111001001",
  3587=>"011001110",
  3588=>"001011111",
  3589=>"100100000",
  3590=>"111001001",
  3591=>"110000110",
  3592=>"000000110",
  3593=>"000001001",
  3594=>"111001000",
  3595=>"000110111",
  3596=>"000110110",
  3597=>"000110110",
  3598=>"100100110",
  3599=>"101110011",
  3600=>"000000100",
  3601=>"000001100",
  3602=>"110111000",
  3603=>"000000000",
  3604=>"000000101",
  3605=>"001001001",
  3606=>"010000011",
  3607=>"100110101",
  3608=>"011000001",
  3609=>"000110111",
  3610=>"000111011",
  3611=>"001001111",
  3612=>"110001101",
  3613=>"000000101",
  3614=>"111111001",
  3615=>"001000000",
  3616=>"000000111",
  3617=>"001111111",
  3618=>"001001000",
  3619=>"011001001",
  3620=>"011110010",
  3621=>"100100100",
  3622=>"111001001",
  3623=>"001111110",
  3624=>"001001101",
  3625=>"001111111",
  3626=>"111000000",
  3627=>"100001000",
  3628=>"000110110",
  3629=>"011000111",
  3630=>"000100111",
  3631=>"111111000",
  3632=>"000111111",
  3633=>"000110100",
  3634=>"001111000",
  3635=>"111001101",
  3636=>"010001000",
  3637=>"001101110",
  3638=>"000001001",
  3639=>"001001001",
  3640=>"011001111",
  3641=>"000000111",
  3642=>"110111001",
  3643=>"001111111",
  3644=>"010100110",
  3645=>"111111000",
  3646=>"000001000",
  3647=>"011001000",
  3648=>"001111110",
  3649=>"100001110",
  3650=>"110000100",
  3651=>"111011000",
  3652=>"011010001",
  3653=>"001111000",
  3654=>"000100110",
  3655=>"000000010",
  3656=>"001110110",
  3657=>"000110110",
  3658=>"111011011",
  3659=>"110111100",
  3660=>"000000000",
  3661=>"000111101",
  3662=>"010100110",
  3663=>"101001000",
  3664=>"011011000",
  3665=>"110000101",
  3666=>"000110111",
  3667=>"000010011",
  3668=>"111001001",
  3669=>"001110001",
  3670=>"101100000",
  3671=>"000010000",
  3672=>"000110000",
  3673=>"000000100",
  3674=>"111101101",
  3675=>"011111111",
  3676=>"010001011",
  3677=>"000011010",
  3678=>"111101001",
  3679=>"001001001",
  3680=>"000110010",
  3681=>"001011011",
  3682=>"100001001",
  3683=>"111011101",
  3684=>"000000101",
  3685=>"000110010",
  3686=>"001100000",
  3687=>"000000001",
  3688=>"000110111",
  3689=>"111110000",
  3690=>"001000000",
  3691=>"100110110",
  3692=>"101011111",
  3693=>"111011110",
  3694=>"110110000",
  3695=>"000111111",
  3696=>"111011011",
  3697=>"000111111",
  3698=>"010011001",
  3699=>"000011111",
  3700=>"000110000",
  3701=>"111001011",
  3702=>"111110110",
  3703=>"010110100",
  3704=>"111110000",
  3705=>"000100000",
  3706=>"000001011",
  3707=>"000110110",
  3708=>"011000111",
  3709=>"000100100",
  3710=>"001000111",
  3711=>"111000000",
  3712=>"000110100",
  3713=>"111111111",
  3714=>"011111010",
  3715=>"001101000",
  3716=>"000111111",
  3717=>"001001000",
  3718=>"100000100",
  3719=>"001000010",
  3720=>"000111110",
  3721=>"111001101",
  3722=>"000000101",
  3723=>"101110010",
  3724=>"010001101",
  3725=>"000000110",
  3726=>"111011011",
  3727=>"110000001",
  3728=>"011101111",
  3729=>"001010001",
  3730=>"110000001",
  3731=>"010001000",
  3732=>"000001001",
  3733=>"110001001",
  3734=>"001110011",
  3735=>"000000010",
  3736=>"000110110",
  3737=>"111001001",
  3738=>"111001001",
  3739=>"111000001",
  3740=>"000000011",
  3741=>"111011001",
  3742=>"001000001",
  3743=>"111001011",
  3744=>"001110111",
  3745=>"011011111",
  3746=>"000001110",
  3747=>"011001000",
  3748=>"001001010",
  3749=>"000101100",
  3750=>"101100000",
  3751=>"110111001",
  3752=>"000001001",
  3753=>"111111111",
  3754=>"111111001",
  3755=>"110011001",
  3756=>"000100000",
  3757=>"110111111",
  3758=>"011001110",
  3759=>"001000100",
  3760=>"101100100",
  3761=>"010011111",
  3762=>"110110111",
  3763=>"000001011",
  3764=>"000010110",
  3765=>"101111000",
  3766=>"000110110",
  3767=>"000110110",
  3768=>"100110110",
  3769=>"000000101",
  3770=>"001110100",
  3771=>"111110110",
  3772=>"111110000",
  3773=>"010011011",
  3774=>"100111011",
  3775=>"001111110",
  3776=>"001001111",
  3777=>"000000000",
  3778=>"111110000",
  3779=>"000010001",
  3780=>"111111110",
  3781=>"000100010",
  3782=>"000000110",
  3783=>"010001000",
  3784=>"001110110",
  3785=>"111001001",
  3786=>"001110100",
  3787=>"001100110",
  3788=>"000000010",
  3789=>"001000110",
  3790=>"111011000",
  3791=>"000110000",
  3792=>"111000001",
  3793=>"000101111",
  3794=>"000101101",
  3795=>"001110110",
  3796=>"111111100",
  3797=>"110110100",
  3798=>"111111000",
  3799=>"000100001",
  3800=>"000000111",
  3801=>"001001001",
  3802=>"001100110",
  3803=>"100000000",
  3804=>"001001001",
  3805=>"001000001",
  3806=>"000110110",
  3807=>"100110001",
  3808=>"110101000",
  3809=>"010000001",
  3810=>"101101111",
  3811=>"001110110",
  3812=>"000000111",
  3813=>"010110110",
  3814=>"011100110",
  3815=>"001001101",
  3816=>"000110111",
  3817=>"000011111",
  3818=>"110000000",
  3819=>"011010110",
  3820=>"111001000",
  3821=>"000000110",
  3822=>"010001000",
  3823=>"110011101",
  3824=>"101000011",
  3825=>"110000010",
  3826=>"000001001",
  3827=>"000101100",
  3828=>"000100010",
  3829=>"110011001",
  3830=>"010010110",
  3831=>"011001001",
  3832=>"001000001",
  3833=>"101110110",
  3834=>"000111111",
  3835=>"001000010",
  3836=>"100111101",
  3837=>"001001000",
  3838=>"000101001",
  3839=>"111111100",
  3840=>"111101111",
  3841=>"000011111",
  3842=>"000000010",
  3843=>"101111111",
  3844=>"000000001",
  3845=>"110110000",
  3846=>"001010011",
  3847=>"000000011",
  3848=>"001000000",
  3849=>"000000000",
  3850=>"111010010",
  3851=>"111110000",
  3852=>"010010000",
  3853=>"010111011",
  3854=>"100001011",
  3855=>"000000100",
  3856=>"111101000",
  3857=>"000000000",
  3858=>"110000000",
  3859=>"101011011",
  3860=>"111101101",
  3861=>"111010000",
  3862=>"000000011",
  3863=>"000100000",
  3864=>"000000000",
  3865=>"000101101",
  3866=>"110111110",
  3867=>"001001100",
  3868=>"000000100",
  3869=>"000000000",
  3870=>"110000011",
  3871=>"111011000",
  3872=>"111111111",
  3873=>"111111111",
  3874=>"101000000",
  3875=>"111111101",
  3876=>"100100111",
  3877=>"111111111",
  3878=>"111011010",
  3879=>"001101001",
  3880=>"000001111",
  3881=>"110111111",
  3882=>"000000000",
  3883=>"010000011",
  3884=>"111111111",
  3885=>"000010000",
  3886=>"111111111",
  3887=>"111111111",
  3888=>"111001111",
  3889=>"001001001",
  3890=>"101100110",
  3891=>"001001111",
  3892=>"011000000",
  3893=>"011111100",
  3894=>"001001000",
  3895=>"111111000",
  3896=>"111111110",
  3897=>"000000000",
  3898=>"000000000",
  3899=>"001101111",
  3900=>"011101101",
  3901=>"111111110",
  3902=>"000000000",
  3903=>"001000010",
  3904=>"101101101",
  3905=>"111111111",
  3906=>"101111111",
  3907=>"000000100",
  3908=>"000000000",
  3909=>"000000000",
  3910=>"100000111",
  3911=>"101000010",
  3912=>"111111100",
  3913=>"000000110",
  3914=>"000000000",
  3915=>"111111101",
  3916=>"011000000",
  3917=>"000000000",
  3918=>"001101011",
  3919=>"111000110",
  3920=>"000111111",
  3921=>"000110010",
  3922=>"111011011",
  3923=>"111001100",
  3924=>"000000000",
  3925=>"000001100",
  3926=>"111011110",
  3927=>"000100100",
  3928=>"111111001",
  3929=>"010110011",
  3930=>"100100101",
  3931=>"101101111",
  3932=>"111111000",
  3933=>"011001011",
  3934=>"000000000",
  3935=>"000000001",
  3936=>"100000000",
  3937=>"111101000",
  3938=>"100010101",
  3939=>"101101100",
  3940=>"110101111",
  3941=>"111101000",
  3942=>"100111000",
  3943=>"000000000",
  3944=>"000001001",
  3945=>"000010110",
  3946=>"010010111",
  3947=>"110110111",
  3948=>"111110110",
  3949=>"000011111",
  3950=>"011100000",
  3951=>"000000111",
  3952=>"111101101",
  3953=>"000111111",
  3954=>"101100001",
  3955=>"111000001",
  3956=>"010000000",
  3957=>"101000011",
  3958=>"000001111",
  3959=>"000000110",
  3960=>"000110000",
  3961=>"111111111",
  3962=>"100111000",
  3963=>"000000001",
  3964=>"100111111",
  3965=>"100100100",
  3966=>"000010110",
  3967=>"000000001",
  3968=>"001011000",
  3969=>"111010010",
  3970=>"111000000",
  3971=>"000000000",
  3972=>"110101101",
  3973=>"001101101",
  3974=>"101111111",
  3975=>"101111100",
  3976=>"111101111",
  3977=>"001101110",
  3978=>"100000000",
  3979=>"000100101",
  3980=>"000000000",
  3981=>"000100111",
  3982=>"111111110",
  3983=>"100000101",
  3984=>"010110011",
  3985=>"110111111",
  3986=>"001001111",
  3987=>"111000010",
  3988=>"001001101",
  3989=>"000000101",
  3990=>"110111000",
  3991=>"001011111",
  3992=>"111000000",
  3993=>"000000000",
  3994=>"111000000",
  3995=>"000000000",
  3996=>"010111000",
  3997=>"101111111",
  3998=>"111100100",
  3999=>"101000000",
  4000=>"000000001",
  4001=>"000000011",
  4002=>"000000000",
  4003=>"010110110",
  4004=>"010111111",
  4005=>"000000000",
  4006=>"010000000",
  4007=>"000010010",
  4008=>"000111111",
  4009=>"101110111",
  4010=>"010001111",
  4011=>"000000101",
  4012=>"110111111",
  4013=>"111001101",
  4014=>"010000011",
  4015=>"010010000",
  4016=>"000000000",
  4017=>"110101101",
  4018=>"000000000",
  4019=>"000000001",
  4020=>"000000101",
  4021=>"000000000",
  4022=>"101111111",
  4023=>"111111111",
  4024=>"111101111",
  4025=>"111101101",
  4026=>"111111111",
  4027=>"000000110",
  4028=>"111111110",
  4029=>"111111111",
  4030=>"100000101",
  4031=>"000000000",
  4032=>"000000000",
  4033=>"100111110",
  4034=>"101111111",
  4035=>"010111111",
  4036=>"000010000",
  4037=>"010010100",
  4038=>"000011010",
  4039=>"000001100",
  4040=>"101000010",
  4041=>"000000000",
  4042=>"111111111",
  4043=>"101000111",
  4044=>"000000100",
  4045=>"011111111",
  4046=>"000010011",
  4047=>"100010110",
  4048=>"000010000",
  4049=>"110100110",
  4050=>"111111110",
  4051=>"000000000",
  4052=>"101101111",
  4053=>"101100110",
  4054=>"110111000",
  4055=>"111000001",
  4056=>"000010000",
  4057=>"111111111",
  4058=>"000000110",
  4059=>"000000000",
  4060=>"000101011",
  4061=>"011000000",
  4062=>"000000111",
  4063=>"011111111",
  4064=>"000000000",
  4065=>"111000101",
  4066=>"000000000",
  4067=>"110101110",
  4068=>"000000111",
  4069=>"010111010",
  4070=>"111111110",
  4071=>"101101100",
  4072=>"110111101",
  4073=>"000000100",
  4074=>"011011011",
  4075=>"010111000",
  4076=>"000000000",
  4077=>"000001111",
  4078=>"000010010",
  4079=>"011001101",
  4080=>"000111011",
  4081=>"010101000",
  4082=>"111011000",
  4083=>"011101000",
  4084=>"111100111",
  4085=>"000000100",
  4086=>"000000000",
  4087=>"101000000",
  4088=>"000000111",
  4089=>"000000000",
  4090=>"000010011",
  4091=>"001111001",
  4092=>"000000100",
  4093=>"100110101",
  4094=>"000000000",
  4095=>"000010010",
  4096=>"010011000",
  4097=>"000000000",
  4098=>"100100101",
  4099=>"011000000",
  4100=>"001011011",
  4101=>"001000000",
  4102=>"010011000",
  4103=>"000011010",
  4104=>"110111111",
  4105=>"000000000",
  4106=>"111000011",
  4107=>"000000010",
  4108=>"010111000",
  4109=>"010101000",
  4110=>"011011001",
  4111=>"001000000",
  4112=>"010000111",
  4113=>"010000111",
  4114=>"000111000",
  4115=>"001111111",
  4116=>"010111101",
  4117=>"100000100",
  4118=>"001111101",
  4119=>"111000011",
  4120=>"001000000",
  4121=>"111100100",
  4122=>"000100101",
  4123=>"111110000",
  4124=>"111111111",
  4125=>"000100100",
  4126=>"011001101",
  4127=>"000000000",
  4128=>"000010010",
  4129=>"110000000",
  4130=>"111111000",
  4131=>"000111011",
  4132=>"001001001",
  4133=>"011000000",
  4134=>"000000110",
  4135=>"000010000",
  4136=>"100100100",
  4137=>"000111000",
  4138=>"101001111",
  4139=>"000000100",
  4140=>"001011011",
  4141=>"000010110",
  4142=>"011011111",
  4143=>"100000100",
  4144=>"000111111",
  4145=>"110100001",
  4146=>"111000011",
  4147=>"000111111",
  4148=>"010100111",
  4149=>"011000000",
  4150=>"110100111",
  4151=>"000100110",
  4152=>"100111000",
  4153=>"000000011",
  4154=>"111111000",
  4155=>"100111111",
  4156=>"110110110",
  4157=>"101101000",
  4158=>"000011001",
  4159=>"110100111",
  4160=>"010111100",
  4161=>"111000000",
  4162=>"001011000",
  4163=>"000000000",
  4164=>"000000000",
  4165=>"000011000",
  4166=>"000010000",
  4167=>"011010100",
  4168=>"000000110",
  4169=>"111011011",
  4170=>"010000000",
  4171=>"101000000",
  4172=>"000110111",
  4173=>"110110110",
  4174=>"011111110",
  4175=>"100010001",
  4176=>"000000001",
  4177=>"110000000",
  4178=>"000011111",
  4179=>"001010110",
  4180=>"011111011",
  4181=>"001100110",
  4182=>"110110100",
  4183=>"101101001",
  4184=>"100000000",
  4185=>"010110100",
  4186=>"100100100",
  4187=>"111110110",
  4188=>"000000000",
  4189=>"001001001",
  4190=>"111100111",
  4191=>"010000000",
  4192=>"000011011",
  4193=>"001101000",
  4194=>"111111000",
  4195=>"100101101",
  4196=>"000111110",
  4197=>"011000000",
  4198=>"110010000",
  4199=>"100100111",
  4200=>"101000110",
  4201=>"111000100",
  4202=>"010111000",
  4203=>"000000000",
  4204=>"000010011",
  4205=>"111100011",
  4206=>"000000011",
  4207=>"011011000",
  4208=>"101111001",
  4209=>"000000000",
  4210=>"011100110",
  4211=>"111100010",
  4212=>"011000000",
  4213=>"000100111",
  4214=>"000010001",
  4215=>"111111110",
  4216=>"111010111",
  4217=>"111011000",
  4218=>"111101100",
  4219=>"000100000",
  4220=>"100110011",
  4221=>"110100101",
  4222=>"111101111",
  4223=>"100100011",
  4224=>"001011111",
  4225=>"110100100",
  4226=>"100111000",
  4227=>"111011000",
  4228=>"000011111",
  4229=>"001011111",
  4230=>"111001000",
  4231=>"000111000",
  4232=>"110110100",
  4233=>"000110110",
  4234=>"011000111",
  4235=>"001000100",
  4236=>"101100100",
  4237=>"000111110",
  4238=>"011111000",
  4239=>"111001000",
  4240=>"001001000",
  4241=>"000000000",
  4242=>"100000111",
  4243=>"000111111",
  4244=>"000011110",
  4245=>"001111001",
  4246=>"000000101",
  4247=>"110010000",
  4248=>"000010111",
  4249=>"111001111",
  4250=>"000000100",
  4251=>"000011101",
  4252=>"000000000",
  4253=>"011011010",
  4254=>"110000000",
  4255=>"000100010",
  4256=>"100100000",
  4257=>"010000111",
  4258=>"111100000",
  4259=>"011011011",
  4260=>"100100111",
  4261=>"111001000",
  4262=>"010101101",
  4263=>"011011011",
  4264=>"010110111",
  4265=>"000011111",
  4266=>"100110111",
  4267=>"011111000",
  4268=>"111111000",
  4269=>"111111001",
  4270=>"110101001",
  4271=>"111111010",
  4272=>"100000000",
  4273=>"000001000",
  4274=>"010100100",
  4275=>"111001100",
  4276=>"111110111",
  4277=>"000000111",
  4278=>"011011000",
  4279=>"000111001",
  4280=>"001011001",
  4281=>"000111011",
  4282=>"010010000",
  4283=>"101100011",
  4284=>"100110000",
  4285=>"101111011",
  4286=>"011001001",
  4287=>"000000011",
  4288=>"101000100",
  4289=>"100100111",
  4290=>"000000010",
  4291=>"000111100",
  4292=>"111111010",
  4293=>"001100011",
  4294=>"010011111",
  4295=>"010010100",
  4296=>"100011011",
  4297=>"100100000",
  4298=>"010000000",
  4299=>"000100110",
  4300=>"111000000",
  4301=>"000011010",
  4302=>"111111101",
  4303=>"111111100",
  4304=>"000100111",
  4305=>"011111011",
  4306=>"100010000",
  4307=>"100100010",
  4308=>"010011010",
  4309=>"100100010",
  4310=>"000111111",
  4311=>"111000001",
  4312=>"110100111",
  4313=>"000000111",
  4314=>"110100011",
  4315=>"011001000",
  4316=>"110111110",
  4317=>"101000111",
  4318=>"001000100",
  4319=>"000100010",
  4320=>"111100100",
  4321=>"000100100",
  4322=>"011000000",
  4323=>"111111110",
  4324=>"011000000",
  4325=>"011011100",
  4326=>"000011000",
  4327=>"010100100",
  4328=>"000100001",
  4329=>"000100111",
  4330=>"111000001",
  4331=>"000101000",
  4332=>"010100100",
  4333=>"000101000",
  4334=>"010010000",
  4335=>"000100111",
  4336=>"111100111",
  4337=>"101001010",
  4338=>"000000011",
  4339=>"100001111",
  4340=>"010001001",
  4341=>"001001010",
  4342=>"000000010",
  4343=>"111000000",
  4344=>"000001000",
  4345=>"000011111",
  4346=>"100101000",
  4347=>"000111111",
  4348=>"100000111",
  4349=>"000100110",
  4350=>"101111111",
  4351=>"011111000",
  4352=>"000001111",
  4353=>"000100101",
  4354=>"000110111",
  4355=>"111010000",
  4356=>"011011010",
  4357=>"101111001",
  4358=>"001101001",
  4359=>"111010111",
  4360=>"000000010",
  4361=>"100000000",
  4362=>"101100101",
  4363=>"010000000",
  4364=>"000000000",
  4365=>"010000000",
  4366=>"011011010",
  4367=>"000001011",
  4368=>"111010000",
  4369=>"000000111",
  4370=>"000010010",
  4371=>"001101000",
  4372=>"000010010",
  4373=>"001101111",
  4374=>"100111111",
  4375=>"010111111",
  4376=>"000000100",
  4377=>"101000110",
  4378=>"000011010",
  4379=>"111010000",
  4380=>"000000010",
  4381=>"101100000",
  4382=>"001001001",
  4383=>"110000000",
  4384=>"000110000",
  4385=>"110000111",
  4386=>"000000110",
  4387=>"110010000",
  4388=>"111001000",
  4389=>"000011110",
  4390=>"110100000",
  4391=>"010010001",
  4392=>"010011111",
  4393=>"110000011",
  4394=>"000101111",
  4395=>"000110110",
  4396=>"011111111",
  4397=>"101111010",
  4398=>"101001000",
  4399=>"000100110",
  4400=>"110001000",
  4401=>"011000010",
  4402=>"010000101",
  4403=>"001001101",
  4404=>"110110110",
  4405=>"011010010",
  4406=>"000011011",
  4407=>"101001000",
  4408=>"000010010",
  4409=>"111001000",
  4410=>"000000000",
  4411=>"111111001",
  4412=>"111100100",
  4413=>"010000100",
  4414=>"000101001",
  4415=>"011011111",
  4416=>"111100111",
  4417=>"100000110",
  4418=>"101001000",
  4419=>"001001111",
  4420=>"001000000",
  4421=>"000000000",
  4422=>"101111100",
  4423=>"001000111",
  4424=>"111111001",
  4425=>"000000000",
  4426=>"000000000",
  4427=>"101111111",
  4428=>"000010010",
  4429=>"111001000",
  4430=>"110100000",
  4431=>"001111111",
  4432=>"000111111",
  4433=>"100111010",
  4434=>"110001101",
  4435=>"001100010",
  4436=>"000001001",
  4437=>"100000110",
  4438=>"011010000",
  4439=>"000101111",
  4440=>"001001101",
  4441=>"111000000",
  4442=>"101101111",
  4443=>"111110011",
  4444=>"001001111",
  4445=>"001110000",
  4446=>"110000000",
  4447=>"100001110",
  4448=>"101111000",
  4449=>"011111010",
  4450=>"000111110",
  4451=>"011011111",
  4452=>"110000000",
  4453=>"011000000",
  4454=>"111001000",
  4455=>"000101010",
  4456=>"111001000",
  4457=>"000011101",
  4458=>"111010011",
  4459=>"000010100",
  4460=>"110010010",
  4461=>"110000111",
  4462=>"000000110",
  4463=>"111110000",
  4464=>"111000110",
  4465=>"111010000",
  4466=>"000111011",
  4467=>"111000000",
  4468=>"111110100",
  4469=>"000111000",
  4470=>"111000000",
  4471=>"100111110",
  4472=>"000111111",
  4473=>"000101000",
  4474=>"110010001",
  4475=>"111001111",
  4476=>"110110000",
  4477=>"100001000",
  4478=>"101111011",
  4479=>"000001111",
  4480=>"111111000",
  4481=>"100000000",
  4482=>"111101000",
  4483=>"111010001",
  4484=>"000000000",
  4485=>"010001111",
  4486=>"001011011",
  4487=>"101000000",
  4488=>"011000011",
  4489=>"110101001",
  4490=>"000010001",
  4491=>"110000001",
  4492=>"000100100",
  4493=>"000001111",
  4494=>"101011110",
  4495=>"001000000",
  4496=>"000110100",
  4497=>"010111000",
  4498=>"111111001",
  4499=>"000101101",
  4500=>"111000001",
  4501=>"000001111",
  4502=>"010011101",
  4503=>"011000000",
  4504=>"001000000",
  4505=>"000000111",
  4506=>"001000010",
  4507=>"000101111",
  4508=>"101000000",
  4509=>"010010101",
  4510=>"111111111",
  4511=>"001000001",
  4512=>"111111110",
  4513=>"001001111",
  4514=>"000000010",
  4515=>"000111111",
  4516=>"000000000",
  4517=>"100000111",
  4518=>"110000000",
  4519=>"010010010",
  4520=>"000111111",
  4521=>"111000011",
  4522=>"000000111",
  4523=>"000101111",
  4524=>"000000000",
  4525=>"000100000",
  4526=>"001010011",
  4527=>"111110001",
  4528=>"010001001",
  4529=>"000011001",
  4530=>"000000000",
  4531=>"011000111",
  4532=>"101110011",
  4533=>"011111111",
  4534=>"111010000",
  4535=>"010000000",
  4536=>"111001001",
  4537=>"111000000",
  4538=>"110100010",
  4539=>"110000111",
  4540=>"110000000",
  4541=>"010111111",
  4542=>"011001011",
  4543=>"000000000",
  4544=>"101111100",
  4545=>"000100111",
  4546=>"010001000",
  4547=>"001000000",
  4548=>"010000000",
  4549=>"001011001",
  4550=>"010000000",
  4551=>"000111001",
  4552=>"111010000",
  4553=>"111101110",
  4554=>"000010100",
  4555=>"111010000",
  4556=>"100100100",
  4557=>"101010000",
  4558=>"101111010",
  4559=>"110111111",
  4560=>"011010000",
  4561=>"110010001",
  4562=>"110010000",
  4563=>"110001010",
  4564=>"000100111",
  4565=>"110111100",
  4566=>"000111101",
  4567=>"111000011",
  4568=>"111001000",
  4569=>"111010011",
  4570=>"111011111",
  4571=>"001000111",
  4572=>"011111111",
  4573=>"000000011",
  4574=>"000000111",
  4575=>"111001000",
  4576=>"000111110",
  4577=>"001001011",
  4578=>"010100101",
  4579=>"010100111",
  4580=>"001101111",
  4581=>"011000000",
  4582=>"111011101",
  4583=>"111011101",
  4584=>"111000000",
  4585=>"000110011",
  4586=>"100111111",
  4587=>"001111111",
  4588=>"000000010",
  4589=>"110000000",
  4590=>"000000000",
  4591=>"101111001",
  4592=>"110000000",
  4593=>"000110110",
  4594=>"000111000",
  4595=>"100011110",
  4596=>"111100001",
  4597=>"001001111",
  4598=>"000001010",
  4599=>"100000011",
  4600=>"101110111",
  4601=>"111000000",
  4602=>"111101010",
  4603=>"111000000",
  4604=>"000111111",
  4605=>"000000100",
  4606=>"110100110",
  4607=>"000100110",
  4608=>"001011011",
  4609=>"001100011",
  4610=>"000001101",
  4611=>"000000000",
  4612=>"011001001",
  4613=>"000000110",
  4614=>"000000101",
  4615=>"110110011",
  4616=>"111000010",
  4617=>"101100111",
  4618=>"101101100",
  4619=>"000000101",
  4620=>"100010110",
  4621=>"001000110",
  4622=>"000010000",
  4623=>"000000011",
  4624=>"001000000",
  4625=>"111111111",
  4626=>"100100111",
  4627=>"000000010",
  4628=>"010000000",
  4629=>"000010000",
  4630=>"110000000",
  4631=>"101000111",
  4632=>"110100010",
  4633=>"001101111",
  4634=>"000010110",
  4635=>"110100000",
  4636=>"100111111",
  4637=>"111111011",
  4638=>"000000000",
  4639=>"101010111",
  4640=>"101101010",
  4641=>"111011000",
  4642=>"111111111",
  4643=>"100000000",
  4644=>"011011111",
  4645=>"000101011",
  4646=>"111110000",
  4647=>"111111111",
  4648=>"110100100",
  4649=>"111110111",
  4650=>"001000101",
  4651=>"000010000",
  4652=>"101111111",
  4653=>"000000001",
  4654=>"000000101",
  4655=>"011111010",
  4656=>"001001000",
  4657=>"011000001",
  4658=>"000000000",
  4659=>"111111100",
  4660=>"000000100",
  4661=>"111000000",
  4662=>"110110011",
  4663=>"110000000",
  4664=>"111111010",
  4665=>"000000110",
  4666=>"000100000",
  4667=>"110011000",
  4668=>"010100000",
  4669=>"110111011",
  4670=>"001000100",
  4671=>"110110110",
  4672=>"101000101",
  4673=>"000110111",
  4674=>"000000000",
  4675=>"111001110",
  4676=>"000110010",
  4677=>"010000000",
  4678=>"000000000",
  4679=>"000000011",
  4680=>"110011111",
  4681=>"000000010",
  4682=>"101000111",
  4683=>"001000110",
  4684=>"111110111",
  4685=>"110000010",
  4686=>"110010100",
  4687=>"101010111",
  4688=>"001111001",
  4689=>"011001000",
  4690=>"000000011",
  4691=>"011000001",
  4692=>"001111111",
  4693=>"100111111",
  4694=>"000001111",
  4695=>"000000101",
  4696=>"000001000",
  4697=>"111110011",
  4698=>"000011001",
  4699=>"100000110",
  4700=>"101101110",
  4701=>"001011011",
  4702=>"010110111",
  4703=>"110100111",
  4704=>"110110110",
  4705=>"001000100",
  4706=>"111111101",
  4707=>"011011100",
  4708=>"010010000",
  4709=>"111111111",
  4710=>"001001101",
  4711=>"111110000",
  4712=>"000110111",
  4713=>"000001000",
  4714=>"011000111",
  4715=>"000000100",
  4716=>"111110110",
  4717=>"000001001",
  4718=>"001101000",
  4719=>"110101100",
  4720=>"011100001",
  4721=>"000001101",
  4722=>"101110111",
  4723=>"011010001",
  4724=>"000000000",
  4725=>"000000010",
  4726=>"111110111",
  4727=>"111110010",
  4728=>"110101101",
  4729=>"111101010",
  4730=>"101000110",
  4731=>"101100010",
  4732=>"001000100",
  4733=>"100100100",
  4734=>"111111100",
  4735=>"000000001",
  4736=>"110011110",
  4737=>"000011001",
  4738=>"000000000",
  4739=>"111101000",
  4740=>"000010101",
  4741=>"111111110",
  4742=>"000110110",
  4743=>"011000001",
  4744=>"000011000",
  4745=>"011011110",
  4746=>"100000100",
  4747=>"010000000",
  4748=>"010010011",
  4749=>"001000000",
  4750=>"010000000",
  4751=>"000000001",
  4752=>"001001100",
  4753=>"010111110",
  4754=>"001011111",
  4755=>"001000000",
  4756=>"111001000",
  4757=>"001100000",
  4758=>"101000111",
  4759=>"111111000",
  4760=>"101000000",
  4761=>"000000001",
  4762=>"000000111",
  4763=>"000000101",
  4764=>"000000101",
  4765=>"110110010",
  4766=>"010001000",
  4767=>"000000111",
  4768=>"110101011",
  4769=>"111101001",
  4770=>"111000111",
  4771=>"101101111",
  4772=>"010011111",
  4773=>"111010000",
  4774=>"110110000",
  4775=>"001101111",
  4776=>"000011111",
  4777=>"111110111",
  4778=>"000000101",
  4779=>"000000100",
  4780=>"111111011",
  4781=>"000011101",
  4782=>"111101111",
  4783=>"010110111",
  4784=>"000111111",
  4785=>"011011101",
  4786=>"000110100",
  4787=>"111011000",
  4788=>"111010001",
  4789=>"110000010",
  4790=>"111111111",
  4791=>"000111111",
  4792=>"010000001",
  4793=>"101100000",
  4794=>"111000000",
  4795=>"000001010",
  4796=>"001001000",
  4797=>"111111111",
  4798=>"111100000",
  4799=>"111111000",
  4800=>"000000101",
  4801=>"000000000",
  4802=>"001111110",
  4803=>"100010110",
  4804=>"010110011",
  4805=>"010110111",
  4806=>"000001011",
  4807=>"000001111",
  4808=>"101001111",
  4809=>"110010000",
  4810=>"111111110",
  4811=>"010010000",
  4812=>"111000010",
  4813=>"100000001",
  4814=>"001000100",
  4815=>"111111000",
  4816=>"111011111",
  4817=>"100100100",
  4818=>"001101111",
  4819=>"000101111",
  4820=>"101111010",
  4821=>"100111111",
  4822=>"000001111",
  4823=>"001111011",
  4824=>"101111111",
  4825=>"110000000",
  4826=>"111111111",
  4827=>"001001101",
  4828=>"011111010",
  4829=>"011000000",
  4830=>"001111000",
  4831=>"001101111",
  4832=>"000000000",
  4833=>"000000100",
  4834=>"010000000",
  4835=>"101101101",
  4836=>"101111111",
  4837=>"111110110",
  4838=>"111000000",
  4839=>"111101110",
  4840=>"111011111",
  4841=>"111111010",
  4842=>"001001101",
  4843=>"000000101",
  4844=>"110010000",
  4845=>"001001110",
  4846=>"000000000",
  4847=>"101100000",
  4848=>"000000010",
  4849=>"001000111",
  4850=>"000000000",
  4851=>"101000100",
  4852=>"101100101",
  4853=>"000100110",
  4854=>"000000000",
  4855=>"000110110",
  4856=>"101001101",
  4857=>"101111110",
  4858=>"100100000",
  4859=>"101101111",
  4860=>"000000111",
  4861=>"000111001",
  4862=>"100100100",
  4863=>"000110010",
  4864=>"000100010",
  4865=>"000000101",
  4866=>"000000001",
  4867=>"001111011",
  4868=>"001000110",
  4869=>"111111111",
  4870=>"101100111",
  4871=>"111111111",
  4872=>"110111111",
  4873=>"000000000",
  4874=>"111111100",
  4875=>"010111000",
  4876=>"000000000",
  4877=>"000010010",
  4878=>"001100101",
  4879=>"000101101",
  4880=>"111101110",
  4881=>"000000111",
  4882=>"000000010",
  4883=>"111110010",
  4884=>"111111111",
  4885=>"010010110",
  4886=>"001000101",
  4887=>"111001001",
  4888=>"000111010",
  4889=>"000000100",
  4890=>"001111110",
  4891=>"010110110",
  4892=>"100100000",
  4893=>"111111111",
  4894=>"001101001",
  4895=>"000000010",
  4896=>"100001111",
  4897=>"111001000",
  4898=>"001100000",
  4899=>"000000000",
  4900=>"000000100",
  4901=>"000000101",
  4902=>"001001110",
  4903=>"000001010",
  4904=>"000011111",
  4905=>"110100011",
  4906=>"011000101",
  4907=>"010000111",
  4908=>"111111100",
  4909=>"111011000",
  4910=>"100100110",
  4911=>"010010010",
  4912=>"000000010",
  4913=>"011101011",
  4914=>"000001010",
  4915=>"100111111",
  4916=>"101101111",
  4917=>"011111111",
  4918=>"001000101",
  4919=>"000000000",
  4920=>"110000111",
  4921=>"000000000",
  4922=>"101011011",
  4923=>"000101000",
  4924=>"100111101",
  4925=>"111011111",
  4926=>"001000111",
  4927=>"110111111",
  4928=>"000111100",
  4929=>"101000000",
  4930=>"000000000",
  4931=>"101000110",
  4932=>"000001101",
  4933=>"000000010",
  4934=>"000101111",
  4935=>"101000110",
  4936=>"011111111",
  4937=>"101101111",
  4938=>"000000111",
  4939=>"111101011",
  4940=>"000111111",
  4941=>"001001001",
  4942=>"100010000",
  4943=>"111101001",
  4944=>"000000101",
  4945=>"011001000",
  4946=>"110000000",
  4947=>"000000001",
  4948=>"000000000",
  4949=>"011011011",
  4950=>"001011010",
  4951=>"000000000",
  4952=>"101111101",
  4953=>"001000101",
  4954=>"111011011",
  4955=>"000101000",
  4956=>"000000001",
  4957=>"000000111",
  4958=>"111111111",
  4959=>"000000101",
  4960=>"101111111",
  4961=>"111111111",
  4962=>"000000000",
  4963=>"111111110",
  4964=>"000000000",
  4965=>"111111100",
  4966=>"111111010",
  4967=>"000111111",
  4968=>"101111111",
  4969=>"111111010",
  4970=>"000001111",
  4971=>"111111110",
  4972=>"111000001",
  4973=>"111111111",
  4974=>"000000111",
  4975=>"101111111",
  4976=>"111110010",
  4977=>"101101000",
  4978=>"001001111",
  4979=>"110111000",
  4980=>"000000011",
  4981=>"000000110",
  4982=>"111000010",
  4983=>"000101010",
  4984=>"010111111",
  4985=>"101000110",
  4986=>"110000001",
  4987=>"111110010",
  4988=>"000001001",
  4989=>"100000000",
  4990=>"110000111",
  4991=>"000000111",
  4992=>"001000000",
  4993=>"111000000",
  4994=>"110111111",
  4995=>"000000000",
  4996=>"111100000",
  4997=>"111111111",
  4998=>"100001111",
  4999=>"000000000",
  5000=>"100101101",
  5001=>"101100000",
  5002=>"000001111",
  5003=>"000000000",
  5004=>"000111111",
  5005=>"110111000",
  5006=>"000000010",
  5007=>"001000100",
  5008=>"111000000",
  5009=>"111000000",
  5010=>"111001111",
  5011=>"111100101",
  5012=>"010111000",
  5013=>"000000100",
  5014=>"001101111",
  5015=>"100001010",
  5016=>"111111011",
  5017=>"101110001",
  5018=>"011111101",
  5019=>"010110110",
  5020=>"111001000",
  5021=>"110111111",
  5022=>"000000011",
  5023=>"000000000",
  5024=>"110100100",
  5025=>"000101111",
  5026=>"000000100",
  5027=>"001001000",
  5028=>"101011100",
  5029=>"000000000",
  5030=>"000111011",
  5031=>"000000100",
  5032=>"111010101",
  5033=>"000001111",
  5034=>"111111010",
  5035=>"111000001",
  5036=>"001111111",
  5037=>"000000100",
  5038=>"011100111",
  5039=>"111011100",
  5040=>"101111000",
  5041=>"100000101",
  5042=>"000001011",
  5043=>"000000011",
  5044=>"111110111",
  5045=>"001001000",
  5046=>"000000000",
  5047=>"101001000",
  5048=>"011100011",
  5049=>"111101001",
  5050=>"110000011",
  5051=>"000111111",
  5052=>"111111010",
  5053=>"111000111",
  5054=>"111111110",
  5055=>"001001011",
  5056=>"000000000",
  5057=>"111111000",
  5058=>"111110011",
  5059=>"000000010",
  5060=>"010001000",
  5061=>"111011111",
  5062=>"110110100",
  5063=>"111011000",
  5064=>"100001010",
  5065=>"000001000",
  5066=>"000001101",
  5067=>"111111100",
  5068=>"100111111",
  5069=>"000100100",
  5070=>"000001111",
  5071=>"000110111",
  5072=>"010111010",
  5073=>"100000001",
  5074=>"000000111",
  5075=>"000000000",
  5076=>"000000000",
  5077=>"001000110",
  5078=>"000000000",
  5079=>"101000010",
  5080=>"000001000",
  5081=>"010010100",
  5082=>"010001001",
  5083=>"111110000",
  5084=>"010001100",
  5085=>"110010111",
  5086=>"000000000",
  5087=>"111111000",
  5088=>"000001000",
  5089=>"001000101",
  5090=>"010111111",
  5091=>"110011011",
  5092=>"000000110",
  5093=>"111111111",
  5094=>"111001000",
  5095=>"000011011",
  5096=>"010010010",
  5097=>"100000000",
  5098=>"111111101",
  5099=>"000000000",
  5100=>"011000100",
  5101=>"001100110",
  5102=>"000000000",
  5103=>"000001000",
  5104=>"111111010",
  5105=>"111100110",
  5106=>"010000000",
  5107=>"110011111",
  5108=>"100000110",
  5109=>"100110011",
  5110=>"010000000",
  5111=>"010101111",
  5112=>"000000001",
  5113=>"011101001",
  5114=>"101000111",
  5115=>"000110010",
  5116=>"010111010",
  5117=>"100110100",
  5118=>"000001010",
  5119=>"111000000",
  5120=>"000011000",
  5121=>"111111111",
  5122=>"000010000",
  5123=>"111101111",
  5124=>"000000000",
  5125=>"111110000",
  5126=>"000111011",
  5127=>"000111111",
  5128=>"000000111",
  5129=>"001000011",
  5130=>"111111011",
  5131=>"111111011",
  5132=>"000000101",
  5133=>"101011001",
  5134=>"001001000",
  5135=>"001000111",
  5136=>"001000111",
  5137=>"111110111",
  5138=>"110110000",
  5139=>"000000000",
  5140=>"110111100",
  5141=>"000110000",
  5142=>"000000011",
  5143=>"111101001",
  5144=>"000000001",
  5145=>"000000110",
  5146=>"010010000",
  5147=>"010000000",
  5148=>"011001000",
  5149=>"000010000",
  5150=>"110000000",
  5151=>"000111000",
  5152=>"111000001",
  5153=>"111111111",
  5154=>"001111000",
  5155=>"000101010",
  5156=>"000000000",
  5157=>"000011000",
  5158=>"111001011",
  5159=>"000000000",
  5160=>"000001111",
  5161=>"111010000",
  5162=>"111000000",
  5163=>"110001011",
  5164=>"000001000",
  5165=>"101011000",
  5166=>"111111111",
  5167=>"101111101",
  5168=>"101111000",
  5169=>"000000001",
  5170=>"111111011",
  5171=>"111110111",
  5172=>"110111111",
  5173=>"101001101",
  5174=>"110111111",
  5175=>"100111111",
  5176=>"111100001",
  5177=>"000000101",
  5178=>"010011010",
  5179=>"001100111",
  5180=>"110111111",
  5181=>"111111000",
  5182=>"000000000",
  5183=>"000000000",
  5184=>"000111111",
  5185=>"000000000",
  5186=>"010111110",
  5187=>"000000110",
  5188=>"011011000",
  5189=>"010000000",
  5190=>"000111111",
  5191=>"111111001",
  5192=>"000000000",
  5193=>"011111111",
  5194=>"000000100",
  5195=>"001000101",
  5196=>"111000010",
  5197=>"000000001",
  5198=>"000000000",
  5199=>"010110000",
  5200=>"111111111",
  5201=>"000000000",
  5202=>"010011111",
  5203=>"101000000",
  5204=>"110110001",
  5205=>"111111011",
  5206=>"000000000",
  5207=>"110111010",
  5208=>"001000000",
  5209=>"000000001",
  5210=>"000000000",
  5211=>"000000000",
  5212=>"000000111",
  5213=>"000000000",
  5214=>"111110000",
  5215=>"100100011",
  5216=>"111111111",
  5217=>"101111100",
  5218=>"000000111",
  5219=>"000000000",
  5220=>"000100101",
  5221=>"000000111",
  5222=>"010111101",
  5223=>"100001000",
  5224=>"100111101",
  5225=>"011100111",
  5226=>"111111101",
  5227=>"111111111",
  5228=>"010111111",
  5229=>"111111000",
  5230=>"111000000",
  5231=>"001010100",
  5232=>"000000000",
  5233=>"010111000",
  5234=>"011101110",
  5235=>"111010000",
  5236=>"111111000",
  5237=>"000000100",
  5238=>"110000110",
  5239=>"111000000",
  5240=>"111101001",
  5241=>"111111000",
  5242=>"111001101",
  5243=>"000000000",
  5244=>"101111111",
  5245=>"000000000",
  5246=>"101111000",
  5247=>"000000111",
  5248=>"111111000",
  5249=>"111000010",
  5250=>"101100111",
  5251=>"101111100",
  5252=>"111111000",
  5253=>"111111000",
  5254=>"111110010",
  5255=>"000000100",
  5256=>"000000000",
  5257=>"110111001",
  5258=>"001111000",
  5259=>"110000011",
  5260=>"101000100",
  5261=>"000011111",
  5262=>"000000000",
  5263=>"101000010",
  5264=>"000000000",
  5265=>"000000100",
  5266=>"101000111",
  5267=>"000000001",
  5268=>"000000000",
  5269=>"111000110",
  5270=>"000111111",
  5271=>"000000000",
  5272=>"101000110",
  5273=>"110111110",
  5274=>"101111110",
  5275=>"111111111",
  5276=>"000001001",
  5277=>"111010001",
  5278=>"111111111",
  5279=>"000000111",
  5280=>"100101000",
  5281=>"000111100",
  5282=>"001111000",
  5283=>"100111000",
  5284=>"101100000",
  5285=>"000000000",
  5286=>"000000000",
  5287=>"001111000",
  5288=>"111111000",
  5289=>"111111000",
  5290=>"101000111",
  5291=>"000000100",
  5292=>"111101000",
  5293=>"000000000",
  5294=>"001101100",
  5295=>"001111111",
  5296=>"001111111",
  5297=>"000000001",
  5298=>"000000011",
  5299=>"001000000",
  5300=>"000000000",
  5301=>"000110100",
  5302=>"011111000",
  5303=>"110001000",
  5304=>"111111111",
  5305=>"000000001",
  5306=>"000111000",
  5307=>"111111111",
  5308=>"111111001",
  5309=>"110000110",
  5310=>"000000000",
  5311=>"011111111",
  5312=>"000000000",
  5313=>"000000100",
  5314=>"111111000",
  5315=>"110001101",
  5316=>"000111000",
  5317=>"001011000",
  5318=>"111110111",
  5319=>"000000110",
  5320=>"000000001",
  5321=>"110010000",
  5322=>"011001110",
  5323=>"011000101",
  5324=>"001001001",
  5325=>"100111111",
  5326=>"000000111",
  5327=>"111111000",
  5328=>"000000000",
  5329=>"000000000",
  5330=>"111111111",
  5331=>"111100000",
  5332=>"101000101",
  5333=>"000000001",
  5334=>"111111011",
  5335=>"111111101",
  5336=>"001101101",
  5337=>"011111101",
  5338=>"000001001",
  5339=>"111000001",
  5340=>"111001000",
  5341=>"111111001",
  5342=>"101101110",
  5343=>"100111111",
  5344=>"000000110",
  5345=>"101100111",
  5346=>"000000001",
  5347=>"001000000",
  5348=>"001000010",
  5349=>"111111000",
  5350=>"000000000",
  5351=>"000000001",
  5352=>"111111110",
  5353=>"000000111",
  5354=>"111111110",
  5355=>"010110011",
  5356=>"111110010",
  5357=>"000000000",
  5358=>"010000000",
  5359=>"000000001",
  5360=>"111111000",
  5361=>"000000000",
  5362=>"110111000",
  5363=>"000000000",
  5364=>"000000000",
  5365=>"111111101",
  5366=>"111111000",
  5367=>"101011000",
  5368=>"000001111",
  5369=>"101111111",
  5370=>"111111111",
  5371=>"001101001",
  5372=>"000000111",
  5373=>"111111001",
  5374=>"000000000",
  5375=>"000110110",
  5376=>"101100110",
  5377=>"111111000",
  5378=>"000010000",
  5379=>"000000000",
  5380=>"000011111",
  5381=>"000000001",
  5382=>"010111111",
  5383=>"010110100",
  5384=>"101001000",
  5385=>"010000000",
  5386=>"010111111",
  5387=>"000000000",
  5388=>"100000000",
  5389=>"101100101",
  5390=>"000000000",
  5391=>"000000000",
  5392=>"000000010",
  5393=>"111111001",
  5394=>"110111000",
  5395=>"111011000",
  5396=>"110111111",
  5397=>"111101111",
  5398=>"111111010",
  5399=>"000010100",
  5400=>"111111000",
  5401=>"111000111",
  5402=>"111100000",
  5403=>"111111000",
  5404=>"000000001",
  5405=>"000001101",
  5406=>"101111111",
  5407=>"000000100",
  5408=>"010011111",
  5409=>"000000100",
  5410=>"101111110",
  5411=>"111101111",
  5412=>"110110100",
  5413=>"000001011",
  5414=>"110000100",
  5415=>"000001111",
  5416=>"000000110",
  5417=>"111100111",
  5418=>"010001111",
  5419=>"000000000",
  5420=>"111111111",
  5421=>"111100000",
  5422=>"110111011",
  5423=>"011111101",
  5424=>"001011010",
  5425=>"010110110",
  5426=>"111101111",
  5427=>"001011111",
  5428=>"111111111",
  5429=>"111111111",
  5430=>"110000000",
  5431=>"101010010",
  5432=>"000111111",
  5433=>"000000100",
  5434=>"000000000",
  5435=>"010010000",
  5436=>"000000001",
  5437=>"111010111",
  5438=>"001000000",
  5439=>"111111110",
  5440=>"000010010",
  5441=>"000011111",
  5442=>"000001111",
  5443=>"000010000",
  5444=>"100000100",
  5445=>"000001111",
  5446=>"111000000",
  5447=>"001001101",
  5448=>"011100010",
  5449=>"100100010",
  5450=>"000000000",
  5451=>"000000010",
  5452=>"110101001",
  5453=>"011110010",
  5454=>"110111011",
  5455=>"001001011",
  5456=>"100111111",
  5457=>"111000010",
  5458=>"100000000",
  5459=>"000010000",
  5460=>"001000000",
  5461=>"000110111",
  5462=>"000110011",
  5463=>"000000100",
  5464=>"001001011",
  5465=>"000001111",
  5466=>"000111100",
  5467=>"111111011",
  5468=>"100000100",
  5469=>"110110000",
  5470=>"010111110",
  5471=>"011001000",
  5472=>"111111111",
  5473=>"001101100",
  5474=>"001000000",
  5475=>"011111111",
  5476=>"010011110",
  5477=>"000000110",
  5478=>"101100100",
  5479=>"010011111",
  5480=>"111110011",
  5481=>"000010000",
  5482=>"000000000",
  5483=>"000000111",
  5484=>"101000101",
  5485=>"010111111",
  5486=>"001000001",
  5487=>"010000000",
  5488=>"011111111",
  5489=>"000000000",
  5490=>"111000100",
  5491=>"000111010",
  5492=>"000000100",
  5493=>"000000011",
  5494=>"100000000",
  5495=>"010000000",
  5496=>"000100000",
  5497=>"111111111",
  5498=>"011011010",
  5499=>"101100000",
  5500=>"011001000",
  5501=>"001011110",
  5502=>"001110110",
  5503=>"100000011",
  5504=>"001111001",
  5505=>"011011011",
  5506=>"010111111",
  5507=>"000011100",
  5508=>"000000111",
  5509=>"111110111",
  5510=>"000100110",
  5511=>"100100100",
  5512=>"111111111",
  5513=>"001101000",
  5514=>"000111000",
  5515=>"000010010",
  5516=>"100110011",
  5517=>"111010001",
  5518=>"000000100",
  5519=>"000000000",
  5520=>"011000111",
  5521=>"101010110",
  5522=>"010011011",
  5523=>"100001000",
  5524=>"111000000",
  5525=>"110000100",
  5526=>"111111111",
  5527=>"111100111",
  5528=>"111111111",
  5529=>"111000000",
  5530=>"111111000",
  5531=>"001000001",
  5532=>"100000100",
  5533=>"110111111",
  5534=>"111111001",
  5535=>"111000000",
  5536=>"111010010",
  5537=>"111111111",
  5538=>"111000110",
  5539=>"001011000",
  5540=>"000010011",
  5541=>"111011000",
  5542=>"000010010",
  5543=>"000011111",
  5544=>"111111110",
  5545=>"010010001",
  5546=>"101000000",
  5547=>"101100000",
  5548=>"000110111",
  5549=>"100000000",
  5550=>"101001110",
  5551=>"001111000",
  5552=>"111000100",
  5553=>"000100101",
  5554=>"000000000",
  5555=>"111100000",
  5556=>"111101011",
  5557=>"000110011",
  5558=>"000000011",
  5559=>"000101111",
  5560=>"000100000",
  5561=>"000000000",
  5562=>"111101000",
  5563=>"010000100",
  5564=>"000100100",
  5565=>"000010010",
  5566=>"110100000",
  5567=>"111111111",
  5568=>"000000000",
  5569=>"000000000",
  5570=>"000011000",
  5571=>"110111111",
  5572=>"000000111",
  5573=>"010111110",
  5574=>"111011111",
  5575=>"000100111",
  5576=>"000000000",
  5577=>"000100000",
  5578=>"000010001",
  5579=>"111000111",
  5580=>"011000000",
  5581=>"110100100",
  5582=>"000111111",
  5583=>"111011011",
  5584=>"011111111",
  5585=>"011101111",
  5586=>"001000100",
  5587=>"001111111",
  5588=>"101000101",
  5589=>"101111110",
  5590=>"000000000",
  5591=>"001000000",
  5592=>"000110111",
  5593=>"101111101",
  5594=>"111011111",
  5595=>"000111111",
  5596=>"000111010",
  5597=>"010111111",
  5598=>"101001111",
  5599=>"000000010",
  5600=>"101000000",
  5601=>"000011000",
  5602=>"011111110",
  5603=>"111111000",
  5604=>"111000100",
  5605=>"000011000",
  5606=>"011011001",
  5607=>"101000100",
  5608=>"111101010",
  5609=>"111101111",
  5610=>"111111110",
  5611=>"111100000",
  5612=>"000001001",
  5613=>"111111111",
  5614=>"111000000",
  5615=>"000000111",
  5616=>"000010110",
  5617=>"010111111",
  5618=>"011001000",
  5619=>"001011001",
  5620=>"011011011",
  5621=>"111111111",
  5622=>"000010111",
  5623=>"000000000",
  5624=>"000000111",
  5625=>"000000100",
  5626=>"000000000",
  5627=>"010000000",
  5628=>"101100101",
  5629=>"000000000",
  5630=>"111111011",
  5631=>"000011011",
  5632=>"011110100",
  5633=>"000100000",
  5634=>"000000110",
  5635=>"110010101",
  5636=>"100100000",
  5637=>"000000000",
  5638=>"111101000",
  5639=>"000001010",
  5640=>"110010010",
  5641=>"010110000",
  5642=>"100010011",
  5643=>"010000001",
  5644=>"000000000",
  5645=>"010111011",
  5646=>"111111111",
  5647=>"000101101",
  5648=>"001000000",
  5649=>"101000110",
  5650=>"111000110",
  5651=>"001000000",
  5652=>"000100101",
  5653=>"111111110",
  5654=>"000110100",
  5655=>"101101110",
  5656=>"000000000",
  5657=>"111111111",
  5658=>"111111111",
  5659=>"110110100",
  5660=>"111111111",
  5661=>"000000000",
  5662=>"000001001",
  5663=>"000000101",
  5664=>"000001000",
  5665=>"010101111",
  5666=>"000111011",
  5667=>"011111111",
  5668=>"001111101",
  5669=>"000000011",
  5670=>"000111111",
  5671=>"111001011",
  5672=>"010010000",
  5673=>"000111111",
  5674=>"111111111",
  5675=>"110001110",
  5676=>"001011100",
  5677=>"000000101",
  5678=>"011000101",
  5679=>"100000001",
  5680=>"000000100",
  5681=>"001111111",
  5682=>"000011110",
  5683=>"001011010",
  5684=>"100000000",
  5685=>"000000111",
  5686=>"010110100",
  5687=>"000010000",
  5688=>"011001010",
  5689=>"100000001",
  5690=>"000000000",
  5691=>"000100001",
  5692=>"110011110",
  5693=>"111111111",
  5694=>"000111000",
  5695=>"000100110",
  5696=>"000000000",
  5697=>"000000100",
  5698=>"111111111",
  5699=>"000000000",
  5700=>"000000001",
  5701=>"101001101",
  5702=>"100111000",
  5703=>"100101111",
  5704=>"101101110",
  5705=>"010000000",
  5706=>"000000000",
  5707=>"000000010",
  5708=>"111111111",
  5709=>"001111001",
  5710=>"011011011",
  5711=>"101111011",
  5712=>"101111111",
  5713=>"000011110",
  5714=>"000101011",
  5715=>"001000100",
  5716=>"000000000",
  5717=>"000001100",
  5718=>"101111011",
  5719=>"010111110",
  5720=>"110110110",
  5721=>"100110110",
  5722=>"100101101",
  5723=>"110100000",
  5724=>"001100110",
  5725=>"001001001",
  5726=>"011001100",
  5727=>"010000000",
  5728=>"110010010",
  5729=>"110000001",
  5730=>"010111011",
  5731=>"111101101",
  5732=>"111110110",
  5733=>"010101011",
  5734=>"010010010",
  5735=>"011111010",
  5736=>"100001001",
  5737=>"101000000",
  5738=>"001001000",
  5739=>"111110101",
  5740=>"111111111",
  5741=>"111111110",
  5742=>"100100100",
  5743=>"111010010",
  5744=>"000111001",
  5745=>"100000011",
  5746=>"000111001",
  5747=>"001001001",
  5748=>"001001001",
  5749=>"000000000",
  5750=>"000100010",
  5751=>"111010001",
  5752=>"001101110",
  5753=>"111001000",
  5754=>"111001111",
  5755=>"000000110",
  5756=>"100111001",
  5757=>"000000000",
  5758=>"000000010",
  5759=>"000000000",
  5760=>"101111111",
  5761=>"000100110",
  5762=>"010000000",
  5763=>"111111011",
  5764=>"101001001",
  5765=>"001100100",
  5766=>"001000000",
  5767=>"000100111",
  5768=>"001011100",
  5769=>"000000000",
  5770=>"111000000",
  5771=>"011000110",
  5772=>"110000000",
  5773=>"000000000",
  5774=>"101000111",
  5775=>"000001000",
  5776=>"100011111",
  5777=>"000001101",
  5778=>"001101110",
  5779=>"111100010",
  5780=>"000000000",
  5781=>"000010010",
  5782=>"010111111",
  5783=>"011010001",
  5784=>"110110110",
  5785=>"000001000",
  5786=>"010000010",
  5787=>"000000110",
  5788=>"010000000",
  5789=>"001010010",
  5790=>"001000000",
  5791=>"011010000",
  5792=>"100111111",
  5793=>"101100000",
  5794=>"111101111",
  5795=>"110110110",
  5796=>"001000000",
  5797=>"011011001",
  5798=>"011111111",
  5799=>"011011111",
  5800=>"000000100",
  5801=>"000000111",
  5802=>"100000111",
  5803=>"000001000",
  5804=>"011101001",
  5805=>"111111111",
  5806=>"100101001",
  5807=>"111111111",
  5808=>"000000010",
  5809=>"011011010",
  5810=>"101100100",
  5811=>"100011110",
  5812=>"100000100",
  5813=>"111110111",
  5814=>"100111010",
  5815=>"000100111",
  5816=>"011110111",
  5817=>"100000001",
  5818=>"111010011",
  5819=>"111010000",
  5820=>"111111111",
  5821=>"010111110",
  5822=>"110011011",
  5823=>"100111111",
  5824=>"000010111",
  5825=>"000000000",
  5826=>"101101100",
  5827=>"001100111",
  5828=>"010001110",
  5829=>"110100111",
  5830=>"110110000",
  5831=>"000000000",
  5832=>"001111111",
  5833=>"000000000",
  5834=>"111111001",
  5835=>"001000010",
  5836=>"011000000",
  5837=>"001110110",
  5838=>"000000000",
  5839=>"110000000",
  5840=>"000000111",
  5841=>"110110110",
  5842=>"110000110",
  5843=>"001001001",
  5844=>"001001000",
  5845=>"100100100",
  5846=>"111011011",
  5847=>"000000111",
  5848=>"111101111",
  5849=>"011011111",
  5850=>"010111110",
  5851=>"000000000",
  5852=>"000100001",
  5853=>"000011110",
  5854=>"100001010",
  5855=>"011010000",
  5856=>"110111010",
  5857=>"100100000",
  5858=>"011100111",
  5859=>"111111110",
  5860=>"101000010",
  5861=>"000000000",
  5862=>"111110000",
  5863=>"011111001",
  5864=>"000101100",
  5865=>"100000000",
  5866=>"010010110",
  5867=>"011000101",
  5868=>"010010010",
  5869=>"000101101",
  5870=>"100010010",
  5871=>"101100111",
  5872=>"000000111",
  5873=>"011111111",
  5874=>"011010000",
  5875=>"011010000",
  5876=>"110011000",
  5877=>"101101001",
  5878=>"100100001",
  5879=>"000101101",
  5880=>"000000111",
  5881=>"000000111",
  5882=>"000100100",
  5883=>"111001000",
  5884=>"101000000",
  5885=>"001000000",
  5886=>"101111111",
  5887=>"001001101",
  5888=>"000001000",
  5889=>"000011001",
  5890=>"110100101",
  5891=>"010011101",
  5892=>"000001000",
  5893=>"110110010",
  5894=>"001011111",
  5895=>"110110111",
  5896=>"110100100",
  5897=>"100100000",
  5898=>"000110100",
  5899=>"000011000",
  5900=>"001001011",
  5901=>"101111111",
  5902=>"000101001",
  5903=>"011010111",
  5904=>"100100010",
  5905=>"100110100",
  5906=>"110001100",
  5907=>"000000100",
  5908=>"010000101",
  5909=>"110111011",
  5910=>"111011000",
  5911=>"100111000",
  5912=>"100000000",
  5913=>"111001011",
  5914=>"010001110",
  5915=>"000100100",
  5916=>"001101101",
  5917=>"100110111",
  5918=>"010110111",
  5919=>"100000000",
  5920=>"000110000",
  5921=>"011001001",
  5922=>"000011101",
  5923=>"010110011",
  5924=>"000100000",
  5925=>"001011001",
  5926=>"100100110",
  5927=>"011001011",
  5928=>"100100000",
  5929=>"010001011",
  5930=>"111111011",
  5931=>"100001010",
  5932=>"000000001",
  5933=>"111111110",
  5934=>"111001011",
  5935=>"101100110",
  5936=>"110100100",
  5937=>"101111111",
  5938=>"011000011",
  5939=>"011001111",
  5940=>"010110100",
  5941=>"000001001",
  5942=>"110110100",
  5943=>"010000010",
  5944=>"001000111",
  5945=>"011001001",
  5946=>"001001001",
  5947=>"100101100",
  5948=>"011011011",
  5949=>"001011001",
  5950=>"001000001",
  5951=>"110111000",
  5952=>"111001001",
  5953=>"000111100",
  5954=>"011011111",
  5955=>"011100000",
  5956=>"011011011",
  5957=>"010010001",
  5958=>"011111000",
  5959=>"100111011",
  5960=>"011001001",
  5961=>"101100010",
  5962=>"010010110",
  5963=>"001011011",
  5964=>"101001001",
  5965=>"000001011",
  5966=>"001100101",
  5967=>"001001011",
  5968=>"001001011",
  5969=>"101000000",
  5970=>"011001011",
  5971=>"011001000",
  5972=>"100100100",
  5973=>"001000000",
  5974=>"110110010",
  5975=>"100100100",
  5976=>"101000000",
  5977=>"001011111",
  5978=>"011011011",
  5979=>"111111101",
  5980=>"111110000",
  5981=>"011111010",
  5982=>"011011111",
  5983=>"100100110",
  5984=>"011011011",
  5985=>"001111001",
  5986=>"001001111",
  5987=>"000000000",
  5988=>"000001000",
  5989=>"001000100",
  5990=>"011111001",
  5991=>"100100100",
  5992=>"110110110",
  5993=>"100110110",
  5994=>"111111011",
  5995=>"010001011",
  5996=>"100000010",
  5997=>"001111100",
  5998=>"001011111",
  5999=>"001011111",
  6000=>"100100101",
  6001=>"000011111",
  6002=>"110110100",
  6003=>"010000100",
  6004=>"011111000",
  6005=>"010000011",
  6006=>"001000000",
  6007=>"111001111",
  6008=>"110111110",
  6009=>"000000110",
  6010=>"110010010",
  6011=>"000000000",
  6012=>"011001000",
  6013=>"100000000",
  6014=>"100100000",
  6015=>"100100000",
  6016=>"011001110",
  6017=>"110110000",
  6018=>"110100100",
  6019=>"011010111",
  6020=>"110000111",
  6021=>"100110100",
  6022=>"011001111",
  6023=>"001011001",
  6024=>"101111100",
  6025=>"011010011",
  6026=>"100110000",
  6027=>"001000110",
  6028=>"100100100",
  6029=>"000010111",
  6030=>"100010000",
  6031=>"001000001",
  6032=>"111101000",
  6033=>"110100110",
  6034=>"100110100",
  6035=>"011011011",
  6036=>"001001011",
  6037=>"110100110",
  6038=>"011001111",
  6039=>"000001000",
  6040=>"010000000",
  6041=>"111001111",
  6042=>"110110000",
  6043=>"110100100",
  6044=>"001001001",
  6045=>"110100000",
  6046=>"010010000",
  6047=>"011001001",
  6048=>"011111111",
  6049=>"100111100",
  6050=>"010000001",
  6051=>"000011000",
  6052=>"000111011",
  6053=>"000000000",
  6054=>"010000010",
  6055=>"011000011",
  6056=>"100100110",
  6057=>"010000000",
  6058=>"111101001",
  6059=>"000000011",
  6060=>"011001000",
  6061=>"001100000",
  6062=>"111011001",
  6063=>"001001110",
  6064=>"000001110",
  6065=>"010001001",
  6066=>"110010100",
  6067=>"000000100",
  6068=>"000111000",
  6069=>"011011111",
  6070=>"011001011",
  6071=>"000001011",
  6072=>"000000001",
  6073=>"011001001",
  6074=>"111001000",
  6075=>"000100110",
  6076=>"001000100",
  6077=>"110100000",
  6078=>"100100000",
  6079=>"110000110",
  6080=>"011001011",
  6081=>"000001000",
  6082=>"000000000",
  6083=>"111101100",
  6084=>"001011011",
  6085=>"000011011",
  6086=>"100001101",
  6087=>"111001011",
  6088=>"111110110",
  6089=>"111000000",
  6090=>"001001010",
  6091=>"110111111",
  6092=>"100100100",
  6093=>"001000001",
  6094=>"100100000",
  6095=>"001110101",
  6096=>"100100110",
  6097=>"101101101",
  6098=>"001001011",
  6099=>"000000100",
  6100=>"000001011",
  6101=>"001011000",
  6102=>"011001001",
  6103=>"110110100",
  6104=>"000000100",
  6105=>"000100000",
  6106=>"001000101",
  6107=>"100110110",
  6108=>"111100000",
  6109=>"011110110",
  6110=>"000000011",
  6111=>"110000011",
  6112=>"000000011",
  6113=>"011000001",
  6114=>"100100000",
  6115=>"001101101",
  6116=>"000100100",
  6117=>"011011100",
  6118=>"001001001",
  6119=>"100101111",
  6120=>"111100011",
  6121=>"110110100",
  6122=>"000110000",
  6123=>"111001011",
  6124=>"011000000",
  6125=>"011101011",
  6126=>"000110000",
  6127=>"001000100",
  6128=>"110110111",
  6129=>"011011001",
  6130=>"011011011",
  6131=>"100000000",
  6132=>"110111000",
  6133=>"000010010",
  6134=>"000001100",
  6135=>"000001011",
  6136=>"011001101",
  6137=>"011110110",
  6138=>"000000000",
  6139=>"110000001",
  6140=>"011011011",
  6141=>"100110000",
  6142=>"111111001",
  6143=>"011001111",
  6144=>"011001000",
  6145=>"100011001",
  6146=>"111100100",
  6147=>"000011011",
  6148=>"111111111",
  6149=>"011011000",
  6150=>"001000000",
  6151=>"011010010",
  6152=>"000100011",
  6153=>"000000100",
  6154=>"001001000",
  6155=>"001011011",
  6156=>"100100110",
  6157=>"000011011",
  6158=>"111001001",
  6159=>"100100000",
  6160=>"011011011",
  6161=>"100000000",
  6162=>"000011000",
  6163=>"011001011",
  6164=>"111011100",
  6165=>"111100100",
  6166=>"110111110",
  6167=>"111110000",
  6168=>"000000100",
  6169=>"111000110",
  6170=>"000100100",
  6171=>"000001111",
  6172=>"111100100",
  6173=>"011101110",
  6174=>"011111000",
  6175=>"110100100",
  6176=>"011001011",
  6177=>"100111100",
  6178=>"000000100",
  6179=>"001000100",
  6180=>"101111100",
  6181=>"001011010",
  6182=>"000010111",
  6183=>"000011010",
  6184=>"111011000",
  6185=>"000000000",
  6186=>"000011000",
  6187=>"100000000",
  6188=>"100101111",
  6189=>"011001001",
  6190=>"111011100",
  6191=>"011001000",
  6192=>"000000011",
  6193=>"001001001",
  6194=>"101100000",
  6195=>"110110011",
  6196=>"011011100",
  6197=>"111100111",
  6198=>"110011000",
  6199=>"110100100",
  6200=>"000100111",
  6201=>"100100100",
  6202=>"000100010",
  6203=>"010100000",
  6204=>"000110110",
  6205=>"000100100",
  6206=>"000000000",
  6207=>"000011011",
  6208=>"101100001",
  6209=>"111111000",
  6210=>"111100000",
  6211=>"011011010",
  6212=>"000100100",
  6213=>"100000001",
  6214=>"110000011",
  6215=>"111101000",
  6216=>"100001000",
  6217=>"010011001",
  6218=>"111111111",
  6219=>"100100100",
  6220=>"111100000",
  6221=>"001001100",
  6222=>"000111111",
  6223=>"101110100",
  6224=>"101111101",
  6225=>"011100000",
  6226=>"101001000",
  6227=>"011001000",
  6228=>"100100000",
  6229=>"000100111",
  6230=>"100001000",
  6231=>"011011011",
  6232=>"110111010",
  6233=>"000000000",
  6234=>"110000000",
  6235=>"011011011",
  6236=>"100100100",
  6237=>"001000101",
  6238=>"111100000",
  6239=>"011011001",
  6240=>"000011000",
  6241=>"000011011",
  6242=>"110000100",
  6243=>"010110110",
  6244=>"000011110",
  6245=>"001111010",
  6246=>"000011000",
  6247=>"100100000",
  6248=>"010011011",
  6249=>"000001110",
  6250=>"000011011",
  6251=>"110110000",
  6252=>"000101111",
  6253=>"101101000",
  6254=>"110100000",
  6255=>"111111011",
  6256=>"000111000",
  6257=>"010011001",
  6258=>"001100100",
  6259=>"000000110",
  6260=>"111000011",
  6261=>"010000001",
  6262=>"011011011",
  6263=>"111001000",
  6264=>"001001010",
  6265=>"000000000",
  6266=>"000100111",
  6267=>"100100101",
  6268=>"111110011",
  6269=>"000010000",
  6270=>"100100000",
  6271=>"011011001",
  6272=>"100000000",
  6273=>"010110100",
  6274=>"011011011",
  6275=>"000001001",
  6276=>"011011010",
  6277=>"001011001",
  6278=>"011001100",
  6279=>"000011000",
  6280=>"000111111",
  6281=>"001001000",
  6282=>"000001001",
  6283=>"110000000",
  6284=>"111101111",
  6285=>"100100100",
  6286=>"100000111",
  6287=>"000000101",
  6288=>"111100001",
  6289=>"111110110",
  6290=>"010000011",
  6291=>"111111111",
  6292=>"000011011",
  6293=>"011001011",
  6294=>"100100100",
  6295=>"110100000",
  6296=>"010011000",
  6297=>"100111011",
  6298=>"111100000",
  6299=>"001011000",
  6300=>"100100000",
  6301=>"000011011",
  6302=>"000000010",
  6303=>"100100100",
  6304=>"111110011",
  6305=>"111110001",
  6306=>"100100000",
  6307=>"010101100",
  6308=>"111010100",
  6309=>"110101000",
  6310=>"001000011",
  6311=>"000000000",
  6312=>"000000111",
  6313=>"000011011",
  6314=>"111100100",
  6315=>"110000100",
  6316=>"110111101",
  6317=>"101001000",
  6318=>"111000010",
  6319=>"001011111",
  6320=>"000001000",
  6321=>"010011100",
  6322=>"100101010",
  6323=>"000000000",
  6324=>"011000011",
  6325=>"111111111",
  6326=>"011010010",
  6327=>"001011000",
  6328=>"100111000",
  6329=>"010111100",
  6330=>"000011000",
  6331=>"000101111",
  6332=>"000111000",
  6333=>"011011011",
  6334=>"010011000",
  6335=>"000000000",
  6336=>"101000000",
  6337=>"110000000",
  6338=>"111011011",
  6339=>"010011000",
  6340=>"000100010",
  6341=>"100101100",
  6342=>"011000001",
  6343=>"111100111",
  6344=>"000111011",
  6345=>"010100100",
  6346=>"100011011",
  6347=>"000011011",
  6348=>"000011010",
  6349=>"100001011",
  6350=>"101000100",
  6351=>"000011011",
  6352=>"000001000",
  6353=>"100110010",
  6354=>"111010100",
  6355=>"111100000",
  6356=>"000011111",
  6357=>"111110111",
  6358=>"111100100",
  6359=>"111001001",
  6360=>"111110111",
  6361=>"000000010",
  6362=>"111100111",
  6363=>"100000001",
  6364=>"110111110",
  6365=>"011001011",
  6366=>"000100101",
  6367=>"011011011",
  6368=>"111100101",
  6369=>"100100100",
  6370=>"000011000",
  6371=>"110111111",
  6372=>"001000000",
  6373=>"000000010",
  6374=>"100001000",
  6375=>"101100011",
  6376=>"011111001",
  6377=>"011011111",
  6378=>"010011000",
  6379=>"100000001",
  6380=>"110111111",
  6381=>"011010010",
  6382=>"000000000",
  6383=>"110000000",
  6384=>"011011000",
  6385=>"010110000",
  6386=>"000000000",
  6387=>"010111000",
  6388=>"011110101",
  6389=>"100000101",
  6390=>"000000000",
  6391=>"000100100",
  6392=>"000110110",
  6393=>"111011000",
  6394=>"011100100",
  6395=>"110111011",
  6396=>"100100010",
  6397=>"000011011",
  6398=>"100001000",
  6399=>"100000100",
  6400=>"100111011",
  6401=>"011001110",
  6402=>"100100100",
  6403=>"110100010",
  6404=>"000011010",
  6405=>"001001000",
  6406=>"000001001",
  6407=>"001111110",
  6408=>"010110100",
  6409=>"001000000",
  6410=>"101111100",
  6411=>"111110010",
  6412=>"100100011",
  6413=>"000000000",
  6414=>"000100011",
  6415=>"011000000",
  6416=>"001100100",
  6417=>"001100100",
  6418=>"000100100",
  6419=>"001101110",
  6420=>"000011011",
  6421=>"100111000",
  6422=>"101101100",
  6423=>"001101100",
  6424=>"011000000",
  6425=>"110111000",
  6426=>"110010000",
  6427=>"101101000",
  6428=>"011000001",
  6429=>"111100000",
  6430=>"011010110",
  6431=>"100000001",
  6432=>"101110010",
  6433=>"000100010",
  6434=>"000010010",
  6435=>"000010111",
  6436=>"110011001",
  6437=>"111001000",
  6438=>"100000001",
  6439=>"011111110",
  6440=>"010111111",
  6441=>"001000000",
  6442=>"001100010",
  6443=>"110111100",
  6444=>"000000011",
  6445=>"101001100",
  6446=>"011011011",
  6447=>"011110010",
  6448=>"011111100",
  6449=>"100110001",
  6450=>"011010110",
  6451=>"010100100",
  6452=>"000011011",
  6453=>"101011010",
  6454=>"001000111",
  6455=>"000110011",
  6456=>"000010000",
  6457=>"100100100",
  6458=>"000001000",
  6459=>"001100100",
  6460=>"110100000",
  6461=>"110000011",
  6462=>"111110100",
  6463=>"100111010",
  6464=>"001100100",
  6465=>"011011100",
  6466=>"011011100",
  6467=>"100111101",
  6468=>"000100001",
  6469=>"001011010",
  6470=>"101111111",
  6471=>"010100000",
  6472=>"111000111",
  6473=>"000111111",
  6474=>"111011111",
  6475=>"001011011",
  6476=>"000001111",
  6477=>"100010000",
  6478=>"100100011",
  6479=>"011110110",
  6480=>"110111000",
  6481=>"001000101",
  6482=>"011101001",
  6483=>"101111000",
  6484=>"011011101",
  6485=>"111110001",
  6486=>"000011001",
  6487=>"001100000",
  6488=>"001011011",
  6489=>"000000001",
  6490=>"111000000",
  6491=>"100101001",
  6492=>"001001111",
  6493=>"000001000",
  6494=>"111011110",
  6495=>"010010110",
  6496=>"110111111",
  6497=>"110010011",
  6498=>"101101111",
  6499=>"100101101",
  6500=>"100000000",
  6501=>"100000011",
  6502=>"010010001",
  6503=>"001011110",
  6504=>"100100001",
  6505=>"011011101",
  6506=>"001010000",
  6507=>"010010010",
  6508=>"000110011",
  6509=>"011001000",
  6510=>"111100001",
  6511=>"001011100",
  6512=>"011101001",
  6513=>"001110100",
  6514=>"000111100",
  6515=>"000110011",
  6516=>"011100111",
  6517=>"000000000",
  6518=>"111100100",
  6519=>"000011111",
  6520=>"011011100",
  6521=>"100111100",
  6522=>"001100111",
  6523=>"100000000",
  6524=>"110100000",
  6525=>"010000110",
  6526=>"010010000",
  6527=>"100111001",
  6528=>"001000100",
  6529=>"000100000",
  6530=>"001011110",
  6531=>"111100001",
  6532=>"110000100",
  6533=>"101111111",
  6534=>"001011011",
  6535=>"000100011",
  6536=>"101100001",
  6537=>"011000001",
  6538=>"011111111",
  6539=>"010010101",
  6540=>"110110001",
  6541=>"100110010",
  6542=>"001100000",
  6543=>"010000000",
  6544=>"000011001",
  6545=>"000010010",
  6546=>"000000001",
  6547=>"010110110",
  6548=>"000100000",
  6549=>"001100100",
  6550=>"000111100",
  6551=>"100000001",
  6552=>"000001000",
  6553=>"100111110",
  6554=>"100101101",
  6555=>"100100111",
  6556=>"110110111",
  6557=>"001011111",
  6558=>"011001111",
  6559=>"110101111",
  6560=>"100011011",
  6561=>"001110010",
  6562=>"100111111",
  6563=>"100010110",
  6564=>"111111100",
  6565=>"111001001",
  6566=>"010011000",
  6567=>"010110111",
  6568=>"001001100",
  6569=>"011010110",
  6570=>"111100100",
  6571=>"000110100",
  6572=>"111000001",
  6573=>"111101110",
  6574=>"001000000",
  6575=>"100110011",
  6576=>"010000110",
  6577=>"110110000",
  6578=>"100000001",
  6579=>"110100000",
  6580=>"111000001",
  6581=>"100111001",
  6582=>"000000011",
  6583=>"011011011",
  6584=>"100111111",
  6585=>"110100000",
  6586=>"001011001",
  6587=>"000000001",
  6588=>"010001001",
  6589=>"101001100",
  6590=>"111001011",
  6591=>"000100110",
  6592=>"000001000",
  6593=>"000000100",
  6594=>"011011111",
  6595=>"110111001",
  6596=>"011011010",
  6597=>"111010001",
  6598=>"001000110",
  6599=>"001100001",
  6600=>"100010000",
  6601=>"001011100",
  6602=>"000100110",
  6603=>"011011011",
  6604=>"100100000",
  6605=>"000110111",
  6606=>"100000000",
  6607=>"100100110",
  6608=>"111100001",
  6609=>"101101011",
  6610=>"001000100",
  6611=>"100000001",
  6612=>"101001111",
  6613=>"000111111",
  6614=>"010011111",
  6615=>"011001110",
  6616=>"011011111",
  6617=>"011000010",
  6618=>"101100011",
  6619=>"111101101",
  6620=>"010100111",
  6621=>"111001111",
  6622=>"001000001",
  6623=>"011111111",
  6624=>"100001011",
  6625=>"100100011",
  6626=>"001100011",
  6627=>"110010001",
  6628=>"000000000",
  6629=>"101011111",
  6630=>"011111100",
  6631=>"100110011",
  6632=>"101110111",
  6633=>"011001100",
  6634=>"011011001",
  6635=>"001101101",
  6636=>"000000010",
  6637=>"010010000",
  6638=>"100000100",
  6639=>"000100000",
  6640=>"000000010",
  6641=>"000000011",
  6642=>"011010110",
  6643=>"000010111",
  6644=>"010010000",
  6645=>"010000001",
  6646=>"000000001",
  6647=>"001110110",
  6648=>"001100100",
  6649=>"010010110",
  6650=>"100000001",
  6651=>"100101001",
  6652=>"111111111",
  6653=>"001001101",
  6654=>"000001011",
  6655=>"010011111",
  6656=>"100000111",
  6657=>"111111101",
  6658=>"111100100",
  6659=>"111011000",
  6660=>"111100100",
  6661=>"111101001",
  6662=>"000000000",
  6663=>"111001101",
  6664=>"111111111",
  6665=>"000000001",
  6666=>"111111001",
  6667=>"000000100",
  6668=>"000000000",
  6669=>"000010111",
  6670=>"000000101",
  6671=>"000110000",
  6672=>"000110100",
  6673=>"111000111",
  6674=>"111101101",
  6675=>"001111000",
  6676=>"100000000",
  6677=>"111111101",
  6678=>"011011100",
  6679=>"111111111",
  6680=>"000000001",
  6681=>"000000000",
  6682=>"111100111",
  6683=>"010010001",
  6684=>"111011010",
  6685=>"000000001",
  6686=>"110111111",
  6687=>"010000010",
  6688=>"000000000",
  6689=>"000000000",
  6690=>"111111011",
  6691=>"111111101",
  6692=>"000000010",
  6693=>"110001010",
  6694=>"110000000",
  6695=>"000010110",
  6696=>"100010000",
  6697=>"000001010",
  6698=>"000000000",
  6699=>"000000000",
  6700=>"100000000",
  6701=>"111111100",
  6702=>"000001111",
  6703=>"101111111",
  6704=>"000111111",
  6705=>"111110101",
  6706=>"000000000",
  6707=>"000001001",
  6708=>"110000000",
  6709=>"111010111",
  6710=>"010000001",
  6711=>"101101111",
  6712=>"101000000",
  6713=>"000000111",
  6714=>"100101100",
  6715=>"011111111",
  6716=>"101100001",
  6717=>"111111111",
  6718=>"010111011",
  6719=>"011111011",
  6720=>"110110000",
  6721=>"010101101",
  6722=>"001000000",
  6723=>"111101100",
  6724=>"000000000",
  6725=>"101101111",
  6726=>"000000000",
  6727=>"000001111",
  6728=>"000011111",
  6729=>"010000000",
  6730=>"000000101",
  6731=>"111111001",
  6732=>"111000101",
  6733=>"010110100",
  6734=>"010011111",
  6735=>"111100101",
  6736=>"000101101",
  6737=>"111111101",
  6738=>"010110010",
  6739=>"001000000",
  6740=>"111111010",
  6741=>"000100100",
  6742=>"010010100",
  6743=>"100100011",
  6744=>"001001010",
  6745=>"000000000",
  6746=>"000111010",
  6747=>"001001001",
  6748=>"010111111",
  6749=>"110110000",
  6750=>"000000111",
  6751=>"110001011",
  6752=>"000000000",
  6753=>"110111011",
  6754=>"110110100",
  6755=>"110111101",
  6756=>"001000000",
  6757=>"010011011",
  6758=>"000000111",
  6759=>"000000001",
  6760=>"000111000",
  6761=>"010011010",
  6762=>"011110111",
  6763=>"000000111",
  6764=>"101001101",
  6765=>"111111111",
  6766=>"000000101",
  6767=>"110010000",
  6768=>"010110111",
  6769=>"100010100",
  6770=>"011000010",
  6771=>"000000011",
  6772=>"000110111",
  6773=>"000000100",
  6774=>"111000000",
  6775=>"100000010",
  6776=>"101010010",
  6777=>"001000011",
  6778=>"000011000",
  6779=>"101111110",
  6780=>"011001001",
  6781=>"001001011",
  6782=>"000000000",
  6783=>"111111111",
  6784=>"000100100",
  6785=>"000011000",
  6786=>"011111110",
  6787=>"000001001",
  6788=>"000100000",
  6789=>"111111110",
  6790=>"110101100",
  6791=>"000000000",
  6792=>"010111011",
  6793=>"001000000",
  6794=>"111010011",
  6795=>"000101111",
  6796=>"000111111",
  6797=>"111111010",
  6798=>"111010110",
  6799=>"000111000",
  6800=>"000100100",
  6801=>"111011000",
  6802=>"000001111",
  6803=>"000011000",
  6804=>"100000000",
  6805=>"111000000",
  6806=>"111111010",
  6807=>"110110100",
  6808=>"010011000",
  6809=>"101111101",
  6810=>"110111000",
  6811=>"011010000",
  6812=>"001000000",
  6813=>"110111010",
  6814=>"010010000",
  6815=>"111001001",
  6816=>"011001001",
  6817=>"111010111",
  6818=>"000000111",
  6819=>"101011111",
  6820=>"000111011",
  6821=>"110100100",
  6822=>"000000100",
  6823=>"000100101",
  6824=>"111110110",
  6825=>"111111101",
  6826=>"111111111",
  6827=>"111000000",
  6828=>"111101001",
  6829=>"000111101",
  6830=>"110100111",
  6831=>"100011111",
  6832=>"001101000",
  6833=>"100110110",
  6834=>"011011001",
  6835=>"100100000",
  6836=>"111101011",
  6837=>"111101101",
  6838=>"000000000",
  6839=>"011011000",
  6840=>"101001101",
  6841=>"000000000",
  6842=>"001010000",
  6843=>"010000110",
  6844=>"001100000",
  6845=>"101000010",
  6846=>"011111010",
  6847=>"000000000",
  6848=>"100100110",
  6849=>"010111111",
  6850=>"000000000",
  6851=>"011001001",
  6852=>"001001101",
  6853=>"000010101",
  6854=>"001000000",
  6855=>"000000111",
  6856=>"001101101",
  6857=>"101000100",
  6858=>"000001000",
  6859=>"000001100",
  6860=>"011010011",
  6861=>"110100100",
  6862=>"000111010",
  6863=>"100101110",
  6864=>"111000111",
  6865=>"001011010",
  6866=>"000000000",
  6867=>"101000010",
  6868=>"011110000",
  6869=>"001011010",
  6870=>"000000001",
  6871=>"111111000",
  6872=>"011111111",
  6873=>"000010001",
  6874=>"101100100",
  6875=>"111111011",
  6876=>"100110000",
  6877=>"101100101",
  6878=>"000000000",
  6879=>"110110000",
  6880=>"001000000",
  6881=>"000111111",
  6882=>"000000110",
  6883=>"111111111",
  6884=>"000000111",
  6885=>"001000000",
  6886=>"001111110",
  6887=>"010011111",
  6888=>"011111010",
  6889=>"000000000",
  6890=>"011111100",
  6891=>"111101111",
  6892=>"100000000",
  6893=>"000010100",
  6894=>"101001000",
  6895=>"111111111",
  6896=>"111111000",
  6897=>"000000100",
  6898=>"100100111",
  6899=>"100000000",
  6900=>"001011001",
  6901=>"100111110",
  6902=>"101101101",
  6903=>"000010011",
  6904=>"000000000",
  6905=>"000111111",
  6906=>"000000000",
  6907=>"100000000",
  6908=>"110111010",
  6909=>"011111111",
  6910=>"011011011",
  6911=>"000101111",
  6912=>"101001001",
  6913=>"011010100",
  6914=>"111000001",
  6915=>"000111000",
  6916=>"111111111",
  6917=>"001111101",
  6918=>"110111110",
  6919=>"011010111",
  6920=>"000000111",
  6921=>"011111110",
  6922=>"011000000",
  6923=>"010000000",
  6924=>"001000100",
  6925=>"001110001",
  6926=>"000000100",
  6927=>"100001001",
  6928=>"101100100",
  6929=>"111001011",
  6930=>"100000000",
  6931=>"110001100",
  6932=>"110011011",
  6933=>"110011111",
  6934=>"101101001",
  6935=>"001111111",
  6936=>"111010111",
  6937=>"000100100",
  6938=>"111111100",
  6939=>"110011000",
  6940=>"111011001",
  6941=>"111010000",
  6942=>"011011000",
  6943=>"100000000",
  6944=>"111011011",
  6945=>"111111100",
  6946=>"110111111",
  6947=>"111111100",
  6948=>"000101011",
  6949=>"111000000",
  6950=>"001001111",
  6951=>"011100110",
  6952=>"110000011",
  6953=>"110111000",
  6954=>"001001101",
  6955=>"100011110",
  6956=>"100101011",
  6957=>"111000010",
  6958=>"111111011",
  6959=>"010111000",
  6960=>"100111001",
  6961=>"001000110",
  6962=>"101100111",
  6963=>"101111100",
  6964=>"011001000",
  6965=>"001011010",
  6966=>"001011001",
  6967=>"000101111",
  6968=>"110111101",
  6969=>"000001001",
  6970=>"100010011",
  6971=>"111011101",
  6972=>"100100000",
  6973=>"000001001",
  6974=>"100000000",
  6975=>"010000110",
  6976=>"110100100",
  6977=>"000011001",
  6978=>"101111111",
  6979=>"001001011",
  6980=>"000000000",
  6981=>"110100000",
  6982=>"011001110",
  6983=>"100111111",
  6984=>"110111111",
  6985=>"011111100",
  6986=>"000001001",
  6987=>"001010100",
  6988=>"101101000",
  6989=>"101101000",
  6990=>"100111111",
  6991=>"100000000",
  6992=>"000100000",
  6993=>"000100100",
  6994=>"001011011",
  6995=>"111011000",
  6996=>"101110000",
  6997=>"100000011",
  6998=>"100111100",
  6999=>"001001000",
  7000=>"000100110",
  7001=>"100010010",
  7002=>"111011000",
  7003=>"101100110",
  7004=>"000111011",
  7005=>"110010001",
  7006=>"111000111",
  7007=>"011001000",
  7008=>"011000111",
  7009=>"110100000",
  7010=>"001000111",
  7011=>"101111011",
  7012=>"000000000",
  7013=>"100110011",
  7014=>"100100100",
  7015=>"000010000",
  7016=>"010000010",
  7017=>"111001001",
  7018=>"111011110",
  7019=>"000110100",
  7020=>"111011111",
  7021=>"111011001",
  7022=>"011011101",
  7023=>"010110110",
  7024=>"001110000",
  7025=>"001000100",
  7026=>"000000001",
  7027=>"101100110",
  7028=>"111111010",
  7029=>"001011111",
  7030=>"011000101",
  7031=>"111011111",
  7032=>"110001000",
  7033=>"000111110",
  7034=>"100100110",
  7035=>"010011101",
  7036=>"000100100",
  7037=>"110000010",
  7038=>"011011111",
  7039=>"111011001",
  7040=>"100001111",
  7041=>"100000001",
  7042=>"110011011",
  7043=>"110111011",
  7044=>"000000110",
  7045=>"001101000",
  7046=>"100011011",
  7047=>"000100000",
  7048=>"000101101",
  7049=>"110100000",
  7050=>"100000011",
  7051=>"101111000",
  7052=>"001100111",
  7053=>"101011111",
  7054=>"000010110",
  7055=>"001010000",
  7056=>"111110000",
  7057=>"001011000",
  7058=>"110101001",
  7059=>"100110110",
  7060=>"000100110",
  7061=>"001001000",
  7062=>"100100100",
  7063=>"111001000",
  7064=>"110110011",
  7065=>"111001111",
  7066=>"011111011",
  7067=>"011000001",
  7068=>"000001000",
  7069=>"000100010",
  7070=>"010011000",
  7071=>"000000000",
  7072=>"011001100",
  7073=>"000001011",
  7074=>"111111001",
  7075=>"000100110",
  7076=>"000101001",
  7077=>"100100000",
  7078=>"010010101",
  7079=>"000000001",
  7080=>"101111000",
  7081=>"100000000",
  7082=>"110000000",
  7083=>"100001001",
  7084=>"110110000",
  7085=>"000010101",
  7086=>"110011000",
  7087=>"000100100",
  7088=>"110000110",
  7089=>"001111111",
  7090=>"001011110",
  7091=>"000100100",
  7092=>"101000011",
  7093=>"010011110",
  7094=>"100100000",
  7095=>"100000000",
  7096=>"110110000",
  7097=>"000110110",
  7098=>"100101001",
  7099=>"101111011",
  7100=>"111010000",
  7101=>"000001111",
  7102=>"011001111",
  7103=>"100100110",
  7104=>"000100000",
  7105=>"000000111",
  7106=>"011001010",
  7107=>"111111000",
  7108=>"000000011",
  7109=>"111100001",
  7110=>"000001001",
  7111=>"001010011",
  7112=>"111011110",
  7113=>"111000001",
  7114=>"101000111",
  7115=>"110000111",
  7116=>"010000001",
  7117=>"000110110",
  7118=>"110111000",
  7119=>"101100000",
  7120=>"011011001",
  7121=>"000100101",
  7122=>"001110110",
  7123=>"100000111",
  7124=>"001000111",
  7125=>"110111011",
  7126=>"011000000",
  7127=>"011011011",
  7128=>"000000101",
  7129=>"100000000",
  7130=>"100000111",
  7131=>"001001111",
  7132=>"110111000",
  7133=>"010000100",
  7134=>"000100000",
  7135=>"001100101",
  7136=>"000011111",
  7137=>"001001100",
  7138=>"001111111",
  7139=>"111111111",
  7140=>"010000000",
  7141=>"011111111",
  7142=>"011001001",
  7143=>"010101111",
  7144=>"101000000",
  7145=>"010000000",
  7146=>"011001001",
  7147=>"100001100",
  7148=>"101000100",
  7149=>"110110000",
  7150=>"000100000",
  7151=>"011001001",
  7152=>"110001000",
  7153=>"110001010",
  7154=>"010111000",
  7155=>"010001011",
  7156=>"001111000",
  7157=>"011001001",
  7158=>"111011000",
  7159=>"011110000",
  7160=>"001111110",
  7161=>"011001111",
  7162=>"100000000",
  7163=>"010110000",
  7164=>"000111000",
  7165=>"000010011",
  7166=>"110110000",
  7167=>"000000000",
  7168=>"001001001",
  7169=>"110000011",
  7170=>"000010000",
  7171=>"011101000",
  7172=>"100011100",
  7173=>"100000111",
  7174=>"010111111",
  7175=>"111111110",
  7176=>"011101100",
  7177=>"111110100",
  7178=>"101000000",
  7179=>"101000001",
  7180=>"010011110",
  7181=>"000000110",
  7182=>"100000100",
  7183=>"111111111",
  7184=>"000000000",
  7185=>"000000010",
  7186=>"111001000",
  7187=>"000101011",
  7188=>"111111000",
  7189=>"111101111",
  7190=>"011101011",
  7191=>"110111111",
  7192=>"100000000",
  7193=>"111111011",
  7194=>"000000101",
  7195=>"000000000",
  7196=>"000000000",
  7197=>"000000000",
  7198=>"101000000",
  7199=>"111001000",
  7200=>"000000010",
  7201=>"111010001",
  7202=>"101000100",
  7203=>"111101100",
  7204=>"100001100",
  7205=>"001000000",
  7206=>"000000001",
  7207=>"110001100",
  7208=>"000000101",
  7209=>"100000000",
  7210=>"100101110",
  7211=>"000000000",
  7212=>"111100001",
  7213=>"000001010",
  7214=>"010010111",
  7215=>"111111111",
  7216=>"111000000",
  7217=>"000000000",
  7218=>"111110111",
  7219=>"001010010",
  7220=>"000000000",
  7221=>"000000000",
  7222=>"000000011",
  7223=>"111111100",
  7224=>"111111111",
  7225=>"000000000",
  7226=>"000000100",
  7227=>"111000000",
  7228=>"111000000",
  7229=>"111111111",
  7230=>"000000000",
  7231=>"100100100",
  7232=>"111111110",
  7233=>"001000000",
  7234=>"000000000",
  7235=>"011011111",
  7236=>"100000111",
  7237=>"111001110",
  7238=>"001010111",
  7239=>"000000111",
  7240=>"000000011",
  7241=>"100000001",
  7242=>"101011111",
  7243=>"111111111",
  7244=>"000000111",
  7245=>"111100001",
  7246=>"111001001",
  7247=>"011000000",
  7248=>"000000000",
  7249=>"111111111",
  7250=>"111100110",
  7251=>"001000000",
  7252=>"000101001",
  7253=>"000100110",
  7254=>"011000000",
  7255=>"000000000",
  7256=>"000001000",
  7257=>"000100000",
  7258=>"010010010",
  7259=>"111011101",
  7260=>"011111111",
  7261=>"110000001",
  7262=>"011111110",
  7263=>"100100000",
  7264=>"000000000",
  7265=>"000100000",
  7266=>"110111000",
  7267=>"011011000",
  7268=>"010100100",
  7269=>"111011100",
  7270=>"000001110",
  7271=>"111110000",
  7272=>"111011000",
  7273=>"110000000",
  7274=>"000001111",
  7275=>"111001111",
  7276=>"000010111",
  7277=>"100000011",
  7278=>"111110001",
  7279=>"000001000",
  7280=>"000100100",
  7281=>"111001001",
  7282=>"001000110",
  7283=>"101000100",
  7284=>"000000101",
  7285=>"000000111",
  7286=>"111100101",
  7287=>"000010010",
  7288=>"010110110",
  7289=>"000000010",
  7290=>"101111111",
  7291=>"000111111",
  7292=>"001100010",
  7293=>"100100100",
  7294=>"111011000",
  7295=>"000001001",
  7296=>"101010010",
  7297=>"111000000",
  7298=>"000111000",
  7299=>"110110111",
  7300=>"000000000",
  7301=>"010101100",
  7302=>"000000001",
  7303=>"011001001",
  7304=>"000111111",
  7305=>"101000010",
  7306=>"110000101",
  7307=>"100000111",
  7308=>"010010000",
  7309=>"100000000",
  7310=>"010111111",
  7311=>"000000000",
  7312=>"101111100",
  7313=>"000000011",
  7314=>"000000010",
  7315=>"001011011",
  7316=>"110000001",
  7317=>"010000000",
  7318=>"110111111",
  7319=>"110101001",
  7320=>"100001010",
  7321=>"000010100",
  7322=>"000100100",
  7323=>"000010010",
  7324=>"000001011",
  7325=>"000000000",
  7326=>"111000011",
  7327=>"111001111",
  7328=>"000100101",
  7329=>"000000010",
  7330=>"111111111",
  7331=>"110110111",
  7332=>"000000111",
  7333=>"001101111",
  7334=>"011010000",
  7335=>"000000111",
  7336=>"111000110",
  7337=>"100110010",
  7338=>"101000000",
  7339=>"010000000",
  7340=>"111110111",
  7341=>"000000000",
  7342=>"000100100",
  7343=>"110111111",
  7344=>"111111111",
  7345=>"100000010",
  7346=>"011011011",
  7347=>"001000100",
  7348=>"010001000",
  7349=>"111111111",
  7350=>"000000100",
  7351=>"010111100",
  7352=>"101100000",
  7353=>"011000110",
  7354=>"000000000",
  7355=>"000100111",
  7356=>"100000000",
  7357=>"000000000",
  7358=>"111111010",
  7359=>"011010111",
  7360=>"000111101",
  7361=>"000000000",
  7362=>"001111111",
  7363=>"001001111",
  7364=>"100000110",
  7365=>"001100000",
  7366=>"100000011",
  7367=>"011011011",
  7368=>"000000000",
  7369=>"101000111",
  7370=>"010000110",
  7371=>"111101000",
  7372=>"111000010",
  7373=>"100001010",
  7374=>"000000010",
  7375=>"000000010",
  7376=>"101101101",
  7377=>"001001100",
  7378=>"101000011",
  7379=>"111111111",
  7380=>"011111011",
  7381=>"100100100",
  7382=>"000000100",
  7383=>"110010000",
  7384=>"111111111",
  7385=>"111100110",
  7386=>"101111111",
  7387=>"111000000",
  7388=>"000001011",
  7389=>"101110011",
  7390=>"111101100",
  7391=>"111101110",
  7392=>"111010011",
  7393=>"111111111",
  7394=>"000001111",
  7395=>"011110000",
  7396=>"000000000",
  7397=>"101110111",
  7398=>"100110000",
  7399=>"010011100",
  7400=>"000000000",
  7401=>"000010010",
  7402=>"100000010",
  7403=>"000010001",
  7404=>"101000000",
  7405=>"000000000",
  7406=>"111000001",
  7407=>"000000111",
  7408=>"000001000",
  7409=>"000001100",
  7410=>"000001110",
  7411=>"001001010",
  7412=>"100000100",
  7413=>"111101110",
  7414=>"000000000",
  7415=>"000010111",
  7416=>"011011000",
  7417=>"111011001",
  7418=>"111111111",
  7419=>"110100000",
  7420=>"011001111",
  7421=>"100110000",
  7422=>"000000001",
  7423=>"000100110",
  7424=>"100000100",
  7425=>"110011101",
  7426=>"011010101",
  7427=>"101001111",
  7428=>"000100111",
  7429=>"110100100",
  7430=>"111000000",
  7431=>"011000101",
  7432=>"111001001",
  7433=>"000000010",
  7434=>"110110000",
  7435=>"110101110",
  7436=>"001000111",
  7437=>"111000010",
  7438=>"110101010",
  7439=>"110010001",
  7440=>"101101000",
  7441=>"011010000",
  7442=>"111110111",
  7443=>"000000000",
  7444=>"101101000",
  7445=>"010011011",
  7446=>"011011111",
  7447=>"110111000",
  7448=>"010000110",
  7449=>"000101001",
  7450=>"011000110",
  7451=>"000111000",
  7452=>"000100100",
  7453=>"000000111",
  7454=>"000000111",
  7455=>"000000111",
  7456=>"010000010",
  7457=>"000101011",
  7458=>"000000010",
  7459=>"001101000",
  7460=>"111111111",
  7461=>"100001001",
  7462=>"110110000",
  7463=>"101011000",
  7464=>"001001111",
  7465=>"011001001",
  7466=>"111001000",
  7467=>"010111011",
  7468=>"000111010",
  7469=>"111110000",
  7470=>"101111010",
  7471=>"001111111",
  7472=>"011010000",
  7473=>"111111110",
  7474=>"101001101",
  7475=>"111111000",
  7476=>"011010010",
  7477=>"010011001",
  7478=>"010011011",
  7479=>"010000110",
  7480=>"101000111",
  7481=>"101100111",
  7482=>"000000111",
  7483=>"111111000",
  7484=>"110111010",
  7485=>"000111111",
  7486=>"000000101",
  7487=>"111111110",
  7488=>"011000000",
  7489=>"000000100",
  7490=>"011010000",
  7491=>"100101001",
  7492=>"000000000",
  7493=>"010010100",
  7494=>"001001111",
  7495=>"000111110",
  7496=>"100101111",
  7497=>"111100111",
  7498=>"101100111",
  7499=>"000111111",
  7500=>"000100101",
  7501=>"111110000",
  7502=>"110010111",
  7503=>"111111000",
  7504=>"000000111",
  7505=>"111111101",
  7506=>"101001111",
  7507=>"011101000",
  7508=>"111110111",
  7509=>"100100011",
  7510=>"110110011",
  7511=>"101100001",
  7512=>"000100011",
  7513=>"000001000",
  7514=>"000000000",
  7515=>"000000011",
  7516=>"000000110",
  7517=>"001000111",
  7518=>"100111001",
  7519=>"001100110",
  7520=>"011101000",
  7521=>"000100111",
  7522=>"101000111",
  7523=>"110100000",
  7524=>"111000111",
  7525=>"110110111",
  7526=>"100000110",
  7527=>"111111010",
  7528=>"000000000",
  7529=>"000000010",
  7530=>"000000000",
  7531=>"111000111",
  7532=>"010111011",
  7533=>"000010010",
  7534=>"111100111",
  7535=>"011010000",
  7536=>"011110111",
  7537=>"000000000",
  7538=>"000010110",
  7539=>"111000100",
  7540=>"000000000",
  7541=>"011000001",
  7542=>"000000000",
  7543=>"111010101",
  7544=>"000000000",
  7545=>"000010111",
  7546=>"000000000",
  7547=>"111111110",
  7548=>"011101001",
  7549=>"010000000",
  7550=>"111111010",
  7551=>"100100111",
  7552=>"111101000",
  7553=>"110000011",
  7554=>"000000101",
  7555=>"000011011",
  7556=>"000000110",
  7557=>"010111110",
  7558=>"001000000",
  7559=>"000000100",
  7560=>"111011010",
  7561=>"010110100",
  7562=>"010000010",
  7563=>"110010111",
  7564=>"111011001",
  7565=>"101011000",
  7566=>"000000100",
  7567=>"000110000",
  7568=>"101111100",
  7569=>"011011110",
  7570=>"000000101",
  7571=>"011111111",
  7572=>"100000001",
  7573=>"000000110",
  7574=>"111101100",
  7575=>"101100110",
  7576=>"000001101",
  7577=>"000000101",
  7578=>"100100101",
  7579=>"110010110",
  7580=>"111100111",
  7581=>"000100101",
  7582=>"000000000",
  7583=>"111010010",
  7584=>"111001000",
  7585=>"111111000",
  7586=>"111111010",
  7587=>"000111111",
  7588=>"000000100",
  7589=>"110100010",
  7590=>"010011101",
  7591=>"001000000",
  7592=>"110111010",
  7593=>"001111101",
  7594=>"111100111",
  7595=>"011000001",
  7596=>"001101101",
  7597=>"100101111",
  7598=>"001000011",
  7599=>"110100111",
  7600=>"110101101",
  7601=>"000001111",
  7602=>"111100011",
  7603=>"000001011",
  7604=>"110110000",
  7605=>"110111010",
  7606=>"001100111",
  7607=>"000000001",
  7608=>"100110110",
  7609=>"001001101",
  7610=>"110010100",
  7611=>"101001111",
  7612=>"001000101",
  7613=>"101000001",
  7614=>"000100111",
  7615=>"111010000",
  7616=>"010010000",
  7617=>"100000001",
  7618=>"000000110",
  7619=>"111110111",
  7620=>"101001000",
  7621=>"011000111",
  7622=>"000100111",
  7623=>"110110111",
  7624=>"111101111",
  7625=>"111010000",
  7626=>"100000001",
  7627=>"100000100",
  7628=>"011000000",
  7629=>"000100100",
  7630=>"000000000",
  7631=>"000101111",
  7632=>"010000000",
  7633=>"011011000",
  7634=>"100101111",
  7635=>"111111110",
  7636=>"000000011",
  7637=>"000111101",
  7638=>"111000000",
  7639=>"001001111",
  7640=>"111111000",
  7641=>"101000011",
  7642=>"110110000",
  7643=>"000000100",
  7644=>"011011010",
  7645=>"101101111",
  7646=>"111111100",
  7647=>"101000111",
  7648=>"010111010",
  7649=>"000010111",
  7650=>"100000111",
  7651=>"111011010",
  7652=>"001000001",
  7653=>"100101111",
  7654=>"110000111",
  7655=>"000010111",
  7656=>"000000111",
  7657=>"011111001",
  7658=>"011010010",
  7659=>"000000101",
  7660=>"101101001",
  7661=>"011111101",
  7662=>"101001010",
  7663=>"010110011",
  7664=>"000010000",
  7665=>"010001001",
  7666=>"000000110",
  7667=>"010011000",
  7668=>"001000010",
  7669=>"000111000",
  7670=>"000100100",
  7671=>"000011000",
  7672=>"000000000",
  7673=>"111011000",
  7674=>"100000100",
  7675=>"011001001",
  7676=>"111111111",
  7677=>"000000000",
  7678=>"110010011",
  7679=>"111000010",
  7680=>"011001100",
  7681=>"011011011",
  7682=>"100100011",
  7683=>"000010011",
  7684=>"111011111",
  7685=>"000000000",
  7686=>"011011011",
  7687=>"011011011",
  7688=>"000000000",
  7689=>"110100110",
  7690=>"000001011",
  7691=>"111011110",
  7692=>"000100110",
  7693=>"100100100",
  7694=>"100000001",
  7695=>"001001101",
  7696=>"000001011",
  7697=>"001001000",
  7698=>"100100110",
  7699=>"000001001",
  7700=>"001011111",
  7701=>"110100110",
  7702=>"001001001",
  7703=>"001001001",
  7704=>"000000001",
  7705=>"011000000",
  7706=>"001010111",
  7707=>"000000000",
  7708=>"011111011",
  7709=>"110110010",
  7710=>"001011110",
  7711=>"000100000",
  7712=>"000001100",
  7713=>"001101101",
  7714=>"111101010",
  7715=>"000100111",
  7716=>"111110110",
  7717=>"101111011",
  7718=>"110010010",
  7719=>"101001000",
  7720=>"000110101",
  7721=>"000100100",
  7722=>"001001011",
  7723=>"100100011",
  7724=>"111110011",
  7725=>"001011101",
  7726=>"010000000",
  7727=>"001000000",
  7728=>"001001100",
  7729=>"011111110",
  7730=>"001000000",
  7731=>"001111001",
  7732=>"000000111",
  7733=>"110011000",
  7734=>"100000000",
  7735=>"010000001",
  7736=>"000110000",
  7737=>"001000100",
  7738=>"110110111",
  7739=>"001001001",
  7740=>"000000000",
  7741=>"111110010",
  7742=>"000100110",
  7743=>"110001100",
  7744=>"111101101",
  7745=>"111110110",
  7746=>"100100000",
  7747=>"000010000",
  7748=>"100100100",
  7749=>"001000000",
  7750=>"011001001",
  7751=>"100110001",
  7752=>"011010000",
  7753=>"001111111",
  7754=>"001000100",
  7755=>"000000000",
  7756=>"000001011",
  7757=>"110110001",
  7758=>"110010101",
  7759=>"110001011",
  7760=>"110000000",
  7761=>"111110111",
  7762=>"000100001",
  7763=>"101100000",
  7764=>"110001001",
  7765=>"011001000",
  7766=>"010110100",
  7767=>"100100111",
  7768=>"001001110",
  7769=>"001011010",
  7770=>"011011110",
  7771=>"110100000",
  7772=>"100011011",
  7773=>"000100011",
  7774=>"101101111",
  7775=>"100100100",
  7776=>"010010010",
  7777=>"010110011",
  7778=>"100100101",
  7779=>"111011101",
  7780=>"001010010",
  7781=>"101010001",
  7782=>"111011110",
  7783=>"110110100",
  7784=>"001111110",
  7785=>"001011101",
  7786=>"001101101",
  7787=>"100110000",
  7788=>"000111111",
  7789=>"001011110",
  7790=>"011000011",
  7791=>"101111001",
  7792=>"001010010",
  7793=>"001001100",
  7794=>"110100000",
  7795=>"000100000",
  7796=>"000100100",
  7797=>"010000110",
  7798=>"110110101",
  7799=>"000000001",
  7800=>"011011111",
  7801=>"001001011",
  7802=>"001001001",
  7803=>"000010000",
  7804=>"110100101",
  7805=>"110000000",
  7806=>"001001001",
  7807=>"110100100",
  7808=>"100001111",
  7809=>"010011000",
  7810=>"100001001",
  7811=>"110100111",
  7812=>"001001001",
  7813=>"111110100",
  7814=>"101101000",
  7815=>"000000000",
  7816=>"000010111",
  7817=>"000000100",
  7818=>"010001000",
  7819=>"000000111",
  7820=>"000010010",
  7821=>"110110111",
  7822=>"010011101",
  7823=>"100100000",
  7824=>"000100100",
  7825=>"011010011",
  7826=>"000001000",
  7827=>"010110100",
  7828=>"000001001",
  7829=>"000000001",
  7830=>"100011111",
  7831=>"101111100",
  7832=>"100111110",
  7833=>"011001011",
  7834=>"100111111",
  7835=>"100100110",
  7836=>"101110010",
  7837=>"000001101",
  7838=>"001011100",
  7839=>"110111011",
  7840=>"010010100",
  7841=>"001010110",
  7842=>"110100011",
  7843=>"101100011",
  7844=>"011001001",
  7845=>"111111101",
  7846=>"001001001",
  7847=>"101001000",
  7848=>"011001001",
  7849=>"001001010",
  7850=>"100100100",
  7851=>"000000000",
  7852=>"000000001",
  7853=>"100000000",
  7854=>"000000110",
  7855=>"001110000",
  7856=>"100100000",
  7857=>"111111101",
  7858=>"000011011",
  7859=>"111110100",
  7860=>"011011100",
  7861=>"110011001",
  7862=>"011110110",
  7863=>"100100111",
  7864=>"110011010",
  7865=>"101111101",
  7866=>"001101101",
  7867=>"001011111",
  7868=>"001010111",
  7869=>"010110111",
  7870=>"010110110",
  7871=>"001010101",
  7872=>"010110010",
  7873=>"010000000",
  7874=>"010111000",
  7875=>"110110110",
  7876=>"001001111",
  7877=>"111011110",
  7878=>"000001001",
  7879=>"010000010",
  7880=>"011011000",
  7881=>"110000000",
  7882=>"110110100",
  7883=>"000111110",
  7884=>"001000111",
  7885=>"000110111",
  7886=>"010000110",
  7887=>"000000100",
  7888=>"100100100",
  7889=>"101110000",
  7890=>"111010100",
  7891=>"001001101",
  7892=>"100100111",
  7893=>"000000011",
  7894=>"000100100",
  7895=>"001001100",
  7896=>"011011010",
  7897=>"001100001",
  7898=>"000000100",
  7899=>"001001001",
  7900=>"000100011",
  7901=>"000001010",
  7902=>"001000010",
  7903=>"001001001",
  7904=>"000100000",
  7905=>"100100111",
  7906=>"101011111",
  7907=>"111110000",
  7908=>"000000000",
  7909=>"110110110",
  7910=>"110010110",
  7911=>"110110001",
  7912=>"110101011",
  7913=>"011011011",
  7914=>"111101100",
  7915=>"011001011",
  7916=>"000100100",
  7917=>"110000010",
  7918=>"010110011",
  7919=>"000000011",
  7920=>"101000001",
  7921=>"100001000",
  7922=>"001001001",
  7923=>"101001101",
  7924=>"000011011",
  7925=>"011011001",
  7926=>"100000001",
  7927=>"001000001",
  7928=>"001001001",
  7929=>"111100000",
  7930=>"111110110",
  7931=>"001110000",
  7932=>"110000011",
  7933=>"100100110",
  7934=>"000000000",
  7935=>"010110001",
  7936=>"000000001",
  7937=>"100000011",
  7938=>"101010010",
  7939=>"011010011",
  7940=>"011101011",
  7941=>"011001000",
  7942=>"000000010",
  7943=>"000000111",
  7944=>"101101000",
  7945=>"000000000",
  7946=>"001001011",
  7947=>"101011101",
  7948=>"100000000",
  7949=>"100100000",
  7950=>"000101001",
  7951=>"000000011",
  7952=>"000000111",
  7953=>"110110010",
  7954=>"111011000",
  7955=>"010101000",
  7956=>"111010001",
  7957=>"100100111",
  7958=>"101111110",
  7959=>"000010010",
  7960=>"111000001",
  7961=>"011101000",
  7962=>"000011101",
  7963=>"000100100",
  7964=>"111000101",
  7965=>"110101111",
  7966=>"110111000",
  7967=>"111100101",
  7968=>"111000000",
  7969=>"010010010",
  7970=>"000000010",
  7971=>"011011010",
  7972=>"100100000",
  7973=>"110100000",
  7974=>"000101000",
  7975=>"000000010",
  7976=>"010111000",
  7977=>"010000111",
  7978=>"000000111",
  7979=>"111000000",
  7980=>"000001011",
  7981=>"010011000",
  7982=>"011101001",
  7983=>"000001000",
  7984=>"010110000",
  7985=>"000100100",
  7986=>"000010000",
  7987=>"010011011",
  7988=>"000100100",
  7989=>"101000001",
  7990=>"100110100",
  7991=>"111000001",
  7992=>"000011111",
  7993=>"101000000",
  7994=>"111000000",
  7995=>"110111001",
  7996=>"011101001",
  7997=>"001100101",
  7998=>"000000010",
  7999=>"000100001",
  8000=>"001111100",
  8001=>"111111000",
  8002=>"011111111",
  8003=>"001000101",
  8004=>"111001000",
  8005=>"111111010",
  8006=>"000100111",
  8007=>"110111010",
  8008=>"000100110",
  8009=>"000110111",
  8010=>"110000000",
  8011=>"000000000",
  8012=>"000110000",
  8013=>"001001100",
  8014=>"110001100",
  8015=>"111000110",
  8016=>"000000010",
  8017=>"010110110",
  8018=>"000111010",
  8019=>"011001100",
  8020=>"001111100",
  8021=>"001101110",
  8022=>"000011100",
  8023=>"110111111",
  8024=>"011001001",
  8025=>"010110110",
  8026=>"011011100",
  8027=>"000000111",
  8028=>"101001000",
  8029=>"110111001",
  8030=>"000111111",
  8031=>"100100100",
  8032=>"010000101",
  8033=>"000010010",
  8034=>"111111111",
  8035=>"110110011",
  8036=>"001000101",
  8037=>"110100000",
  8038=>"110110001",
  8039=>"111111001",
  8040=>"001101100",
  8041=>"000011010",
  8042=>"010111100",
  8043=>"000000000",
  8044=>"011010000",
  8045=>"000010010",
  8046=>"100000100",
  8047=>"000000000",
  8048=>"111001001",
  8049=>"111111011",
  8050=>"000001001",
  8051=>"111000000",
  8052=>"011011101",
  8053=>"101000100",
  8054=>"000000001",
  8055=>"000111111",
  8056=>"111110111",
  8057=>"000101000",
  8058=>"110000110",
  8059=>"001010000",
  8060=>"000110111",
  8061=>"100100000",
  8062=>"011110000",
  8063=>"101000000",
  8064=>"001100111",
  8065=>"111111001",
  8066=>"000111111",
  8067=>"011111111",
  8068=>"000001000",
  8069=>"000110111",
  8070=>"011011001",
  8071=>"000000110",
  8072=>"101100100",
  8073=>"000111011",
  8074=>"111010000",
  8075=>"111011010",
  8076=>"101000000",
  8077=>"101010000",
  8078=>"001111011",
  8079=>"011001011",
  8080=>"000001001",
  8081=>"100101100",
  8082=>"000110001",
  8083=>"110001010",
  8084=>"000000011",
  8085=>"010111110",
  8086=>"001100010",
  8087=>"000100001",
  8088=>"111010110",
  8089=>"001000110",
  8090=>"001111000",
  8091=>"100100111",
  8092=>"011111111",
  8093=>"100010011",
  8094=>"011111001",
  8095=>"010101111",
  8096=>"100100010",
  8097=>"111010010",
  8098=>"000101101",
  8099=>"000000010",
  8100=>"110111101",
  8101=>"000001001",
  8102=>"001100000",
  8103=>"100100000",
  8104=>"111111110",
  8105=>"101111111",
  8106=>"000000101",
  8107=>"000010000",
  8108=>"111111111",
  8109=>"000111111",
  8110=>"111001000",
  8111=>"000111111",
  8112=>"111111000",
  8113=>"110110000",
  8114=>"111101011",
  8115=>"000001001",
  8116=>"110110110",
  8117=>"000010010",
  8118=>"001101100",
  8119=>"101011010",
  8120=>"010100100",
  8121=>"100000110",
  8122=>"100101010",
  8123=>"111111000",
  8124=>"000000010",
  8125=>"000011100",
  8126=>"100110100",
  8127=>"000010111",
  8128=>"011000000",
  8129=>"000001110",
  8130=>"011111111",
  8131=>"001100100",
  8132=>"000010000",
  8133=>"001000111",
  8134=>"000110100",
  8135=>"100000011",
  8136=>"111111111",
  8137=>"111000001",
  8138=>"011000000",
  8139=>"101111111",
  8140=>"001000111",
  8141=>"001011111",
  8142=>"100100110",
  8143=>"000110111",
  8144=>"000011000",
  8145=>"001001001",
  8146=>"111111010",
  8147=>"100001001",
  8148=>"000101111",
  8149=>"011001000",
  8150=>"101000011",
  8151=>"111111110",
  8152=>"100101001",
  8153=>"010101000",
  8154=>"001001000",
  8155=>"000000010",
  8156=>"100101011",
  8157=>"101000111",
  8158=>"000110111",
  8159=>"111111111",
  8160=>"000101111",
  8161=>"111001100",
  8162=>"000001111",
  8163=>"011001001",
  8164=>"010100000",
  8165=>"111111101",
  8166=>"101111000",
  8167=>"001000000",
  8168=>"111000000",
  8169=>"111000011",
  8170=>"100110110",
  8171=>"000101101",
  8172=>"000000000",
  8173=>"111100111",
  8174=>"010000000",
  8175=>"100000011",
  8176=>"100101100",
  8177=>"000001001",
  8178=>"111011000",
  8179=>"011001001",
  8180=>"100100001",
  8181=>"000000001",
  8182=>"000000111",
  8183=>"000111100",
  8184=>"001001011",
  8185=>"000100010",
  8186=>"010111111",
  8187=>"000000111",
  8188=>"101111111",
  8189=>"101111010",
  8190=>"110110000",
  8191=>"001011011",
  8192=>"111111100",
  8193=>"000011001",
  8194=>"101000101",
  8195=>"000000111",
  8196=>"001001011",
  8197=>"001000000",
  8198=>"111111111",
  8199=>"111101101",
  8200=>"010011001",
  8201=>"110100000",
  8202=>"000000110",
  8203=>"101111101",
  8204=>"000011000",
  8205=>"011000011",
  8206=>"100010011",
  8207=>"110000010",
  8208=>"011000000",
  8209=>"101000101",
  8210=>"100000100",
  8211=>"000000000",
  8212=>"111111101",
  8213=>"000000010",
  8214=>"101001001",
  8215=>"000000001",
  8216=>"000000111",
  8217=>"010000001",
  8218=>"000010111",
  8219=>"010110000",
  8220=>"000000000",
  8221=>"010000000",
  8222=>"000100001",
  8223=>"000001000",
  8224=>"111000100",
  8225=>"110100110",
  8226=>"001000000",
  8227=>"111010000",
  8228=>"000000100",
  8229=>"000100110",
  8230=>"000000000",
  8231=>"000000000",
  8232=>"100110111",
  8233=>"111111111",
  8234=>"001000000",
  8235=>"011000000",
  8236=>"011011111",
  8237=>"111111110",
  8238=>"001000010",
  8239=>"110100000",
  8240=>"101001011",
  8241=>"001011111",
  8242=>"010101000",
  8243=>"000100110",
  8244=>"000001100",
  8245=>"111110000",
  8246=>"000100000",
  8247=>"010101000",
  8248=>"101101000",
  8249=>"000001001",
  8250=>"010000100",
  8251=>"111000001",
  8252=>"101100100",
  8253=>"110111111",
  8254=>"000010000",
  8255=>"100011001",
  8256=>"101010010",
  8257=>"000011111",
  8258=>"101111110",
  8259=>"000000100",
  8260=>"111101100",
  8261=>"011000000",
  8262=>"110111000",
  8263=>"010010000",
  8264=>"111000000",
  8265=>"111011000",
  8266=>"000000000",
  8267=>"001101111",
  8268=>"000101111",
  8269=>"000000111",
  8270=>"100101011",
  8271=>"101101111",
  8272=>"001000001",
  8273=>"000011001",
  8274=>"010011000",
  8275=>"001101001",
  8276=>"000011000",
  8277=>"101001001",
  8278=>"000101001",
  8279=>"101101000",
  8280=>"110001111",
  8281=>"011101011",
  8282=>"001111111",
  8283=>"000011111",
  8284=>"001000110",
  8285=>"100000001",
  8286=>"011111111",
  8287=>"000001101",
  8288=>"000111111",
  8289=>"111101110",
  8290=>"000111011",
  8291=>"110000101",
  8292=>"001111110",
  8293=>"011001001",
  8294=>"111110110",
  8295=>"111010110",
  8296=>"000010011",
  8297=>"011001101",
  8298=>"010010000",
  8299=>"000000010",
  8300=>"111000001",
  8301=>"010000010",
  8302=>"010000010",
  8303=>"000000000",
  8304=>"001111111",
  8305=>"101111101",
  8306=>"001001100",
  8307=>"101010000",
  8308=>"000111011",
  8309=>"001100100",
  8310=>"000101011",
  8311=>"111111001",
  8312=>"111000000",
  8313=>"110010010",
  8314=>"001000000",
  8315=>"011000100",
  8316=>"011000000",
  8317=>"111111100",
  8318=>"111010000",
  8319=>"100000111",
  8320=>"001000000",
  8321=>"000101111",
  8322=>"110000000",
  8323=>"010100000",
  8324=>"110010010",
  8325=>"111111111",
  8326=>"000001111",
  8327=>"011000100",
  8328=>"111111101",
  8329=>"100101111",
  8330=>"010100011",
  8331=>"000000001",
  8332=>"000101100",
  8333=>"100110010",
  8334=>"101111001",
  8335=>"100001000",
  8336=>"110111000",
  8337=>"010111000",
  8338=>"101111010",
  8339=>"000010000",
  8340=>"010011111",
  8341=>"000000010",
  8342=>"111101010",
  8343=>"100110110",
  8344=>"110011010",
  8345=>"000000100",
  8346=>"110110000",
  8347=>"010010111",
  8348=>"001000010",
  8349=>"100010000",
  8350=>"101011111",
  8351=>"111001101",
  8352=>"000100100",
  8353=>"100011001",
  8354=>"100000111",
  8355=>"000000000",
  8356=>"010000000",
  8357=>"000010110",
  8358=>"011010111",
  8359=>"010110010",
  8360=>"101000000",
  8361=>"001000010",
  8362=>"101010001",
  8363=>"111101001",
  8364=>"111111100",
  8365=>"100000000",
  8366=>"111111000",
  8367=>"011010010",
  8368=>"000000010",
  8369=>"011000001",
  8370=>"101101101",
  8371=>"001001001",
  8372=>"011011001",
  8373=>"011111000",
  8374=>"000110110",
  8375=>"110111111",
  8376=>"100011001",
  8377=>"110110110",
  8378=>"101111111",
  8379=>"000000010",
  8380=>"111111010",
  8381=>"111111111",
  8382=>"010111100",
  8383=>"000000111",
  8384=>"101000101",
  8385=>"000011010",
  8386=>"000111100",
  8387=>"010111000",
  8388=>"010111001",
  8389=>"000001111",
  8390=>"111000101",
  8391=>"100000010",
  8392=>"111000001",
  8393=>"000100101",
  8394=>"101000101",
  8395=>"101000100",
  8396=>"100010110",
  8397=>"110000000",
  8398=>"010111000",
  8399=>"010110101",
  8400=>"010111000",
  8401=>"110110001",
  8402=>"010000110",
  8403=>"011101011",
  8404=>"001110111",
  8405=>"000001101",
  8406=>"100000110",
  8407=>"010111111",
  8408=>"101001101",
  8409=>"000000001",
  8410=>"100000001",
  8411=>"000000111",
  8412=>"101111101",
  8413=>"011010010",
  8414=>"010110110",
  8415=>"010000000",
  8416=>"000100011",
  8417=>"100101101",
  8418=>"010111101",
  8419=>"101111100",
  8420=>"000000011",
  8421=>"111111001",
  8422=>"000011010",
  8423=>"011011000",
  8424=>"000000010",
  8425=>"101000111",
  8426=>"000000111",
  8427=>"101111111",
  8428=>"000001000",
  8429=>"101011110",
  8430=>"000111000",
  8431=>"110101000",
  8432=>"110111000",
  8433=>"000100101",
  8434=>"000000110",
  8435=>"110011101",
  8436=>"110110000",
  8437=>"000000111",
  8438=>"000000111",
  8439=>"001000000",
  8440=>"101000000",
  8441=>"000000000",
  8442=>"111111011",
  8443=>"010101101",
  8444=>"101100001",
  8445=>"000111111",
  8446=>"110111000",
  8447=>"001111000",
  8448=>"011011110",
  8449=>"100000011",
  8450=>"100000100",
  8451=>"100000010",
  8452=>"100011011",
  8453=>"101100100",
  8454=>"111110110",
  8455=>"000001001",
  8456=>"110100100",
  8457=>"000011111",
  8458=>"110111000",
  8459=>"000100100",
  8460=>"100000000",
  8461=>"000111100",
  8462=>"000111011",
  8463=>"011011100",
  8464=>"111000100",
  8465=>"000000000",
  8466=>"010100000",
  8467=>"010000000",
  8468=>"111000101",
  8469=>"000110011",
  8470=>"001110001",
  8471=>"000011010",
  8472=>"001100100",
  8473=>"011100000",
  8474=>"000011000",
  8475=>"111100100",
  8476=>"010111111",
  8477=>"100000100",
  8478=>"111011000",
  8479=>"010010110",
  8480=>"000011000",
  8481=>"111100000",
  8482=>"101101011",
  8483=>"010011011",
  8484=>"000110100",
  8485=>"010011000",
  8486=>"001010000",
  8487=>"110011000",
  8488=>"101000100",
  8489=>"101100100",
  8490=>"111100100",
  8491=>"011111111",
  8492=>"010011011",
  8493=>"111101010",
  8494=>"111100000",
  8495=>"010000000",
  8496=>"000110011",
  8497=>"000110000",
  8498=>"000010011",
  8499=>"011100111",
  8500=>"111100000",
  8501=>"101111111",
  8502=>"101111110",
  8503=>"100100100",
  8504=>"111001101",
  8505=>"111100000",
  8506=>"110100111",
  8507=>"110100111",
  8508=>"010011000",
  8509=>"000111010",
  8510=>"100000000",
  8511=>"011111111",
  8512=>"100110011",
  8513=>"111001000",
  8514=>"110110000",
  8515=>"111011110",
  8516=>"111101111",
  8517=>"100000101",
  8518=>"000000011",
  8519=>"110011111",
  8520=>"001000100",
  8521=>"011011010",
  8522=>"111111111",
  8523=>"100011111",
  8524=>"000100000",
  8525=>"100101110",
  8526=>"111101000",
  8527=>"111101111",
  8528=>"110111111",
  8529=>"111100000",
  8530=>"101000100",
  8531=>"011001010",
  8532=>"111100100",
  8533=>"100110100",
  8534=>"001011000",
  8535=>"001011011",
  8536=>"011010100",
  8537=>"100100100",
  8538=>"110011011",
  8539=>"011011001",
  8540=>"000011100",
  8541=>"000101001",
  8542=>"101100101",
  8543=>"000100111",
  8544=>"011100000",
  8545=>"000000110",
  8546=>"011011010",
  8547=>"001000000",
  8548=>"100111100",
  8549=>"110100111",
  8550=>"010111011",
  8551=>"110011011",
  8552=>"000111111",
  8553=>"000000100",
  8554=>"011011011",
  8555=>"111111011",
  8556=>"111111110",
  8557=>"000000100",
  8558=>"000000011",
  8559=>"111111000",
  8560=>"100111100",
  8561=>"110000000",
  8562=>"010000000",
  8563=>"001011001",
  8564=>"111111111",
  8565=>"100000110",
  8566=>"000111011",
  8567=>"011000011",
  8568=>"111101111",
  8569=>"000000011",
  8570=>"101100101",
  8571=>"000100100",
  8572=>"000110011",
  8573=>"001110100",
  8574=>"011011011",
  8575=>"000011011",
  8576=>"000100111",
  8577=>"000011011",
  8578=>"111111011",
  8579=>"011110000",
  8580=>"110100100",
  8581=>"111100111",
  8582=>"010001110",
  8583=>"100110010",
  8584=>"000111000",
  8585=>"000111100",
  8586=>"111100011",
  8587=>"011011011",
  8588=>"100000111",
  8589=>"111111111",
  8590=>"011101001",
  8591=>"100001001",
  8592=>"100110011",
  8593=>"010000110",
  8594=>"111000000",
  8595=>"100000000",
  8596=>"011011001",
  8597=>"111000100",
  8598=>"111100110",
  8599=>"000001000",
  8600=>"011011010",
  8601=>"000010011",
  8602=>"010010010",
  8603=>"011000001",
  8604=>"110100100",
  8605=>"111100100",
  8606=>"111000111",
  8607=>"000100100",
  8608=>"100100100",
  8609=>"000100000",
  8610=>"110100100",
  8611=>"100000111",
  8612=>"111011011",
  8613=>"000100010",
  8614=>"101111111",
  8615=>"111100110",
  8616=>"100010000",
  8617=>"010100100",
  8618=>"100100111",
  8619=>"100100100",
  8620=>"101000101",
  8621=>"011100100",
  8622=>"110111110",
  8623=>"111000000",
  8624=>"000100100",
  8625=>"000011001",
  8626=>"000101100",
  8627=>"000010010",
  8628=>"011101001",
  8629=>"111111111",
  8630=>"111100100",
  8631=>"011011001",
  8632=>"101110100",
  8633=>"000011011",
  8634=>"010111111",
  8635=>"011011001",
  8636=>"000100100",
  8637=>"011011011",
  8638=>"011110111",
  8639=>"100000100",
  8640=>"110000000",
  8641=>"011010000",
  8642=>"000111111",
  8643=>"011111110",
  8644=>"000000001",
  8645=>"111001001",
  8646=>"110111101",
  8647=>"000011010",
  8648=>"101100100",
  8649=>"011011100",
  8650=>"001100111",
  8651=>"010111111",
  8652=>"110100100",
  8653=>"100011111",
  8654=>"000000010",
  8655=>"100111011",
  8656=>"111011000",
  8657=>"011101011",
  8658=>"110110100",
  8659=>"011000011",
  8660=>"011011000",
  8661=>"000000110",
  8662=>"111100000",
  8663=>"100001111",
  8664=>"011001001",
  8665=>"000100000",
  8666=>"011011001",
  8667=>"101000100",
  8668=>"111001001",
  8669=>"110101000",
  8670=>"111100100",
  8671=>"011110100",
  8672=>"000000000",
  8673=>"101100111",
  8674=>"101000000",
  8675=>"100110100",
  8676=>"000000000",
  8677=>"100000000",
  8678=>"111100000",
  8679=>"010011001",
  8680=>"011010000",
  8681=>"000000011",
  8682=>"011011000",
  8683=>"000111011",
  8684=>"011110100",
  8685=>"000000100",
  8686=>"001000000",
  8687=>"011001010",
  8688=>"110100100",
  8689=>"100000100",
  8690=>"000010011",
  8691=>"010100111",
  8692=>"111110000",
  8693=>"101010111",
  8694=>"000100000",
  8695=>"111100110",
  8696=>"000000000",
  8697=>"111101000",
  8698=>"100000000",
  8699=>"101111100",
  8700=>"010110110",
  8701=>"000000000",
  8702=>"001110111",
  8703=>"111111011",
  8704=>"001011101",
  8705=>"111100000",
  8706=>"101100100",
  8707=>"110011010",
  8708=>"010011001",
  8709=>"011010000",
  8710=>"100100100",
  8711=>"000010011",
  8712=>"000011010",
  8713=>"000000010",
  8714=>"110100101",
  8715=>"000100000",
  8716=>"111100111",
  8717=>"100100000",
  8718=>"101011011",
  8719=>"000000100",
  8720=>"010011011",
  8721=>"110100011",
  8722=>"111100100",
  8723=>"000000011",
  8724=>"101011100",
  8725=>"110111000",
  8726=>"001110110",
  8727=>"111111000",
  8728=>"101000000",
  8729=>"000111011",
  8730=>"001011000",
  8731=>"011000001",
  8732=>"100100100",
  8733=>"111001001",
  8734=>"000010000",
  8735=>"100100100",
  8736=>"110011011",
  8737=>"001011100",
  8738=>"000011100",
  8739=>"011100000",
  8740=>"001001011",
  8741=>"100101000",
  8742=>"000011011",
  8743=>"110010100",
  8744=>"101011101",
  8745=>"010011111",
  8746=>"000010010",
  8747=>"001011010",
  8748=>"000001001",
  8749=>"101110001",
  8750=>"011011011",
  8751=>"011111001",
  8752=>"100101111",
  8753=>"011011010",
  8754=>"000110111",
  8755=>"000100111",
  8756=>"111100000",
  8757=>"001011000",
  8758=>"110110001",
  8759=>"001100000",
  8760=>"000100011",
  8761=>"111100101",
  8762=>"100100111",
  8763=>"000000100",
  8764=>"000000100",
  8765=>"011111000",
  8766=>"000000000",
  8767=>"000011010",
  8768=>"100000101",
  8769=>"001011111",
  8770=>"111011110",
  8771=>"000011001",
  8772=>"111111011",
  8773=>"100000100",
  8774=>"100100000",
  8775=>"000011100",
  8776=>"110101111",
  8777=>"000100111",
  8778=>"101100100",
  8779=>"000000100",
  8780=>"000011011",
  8781=>"000101100",
  8782=>"000011101",
  8783=>"100100001",
  8784=>"101011000",
  8785=>"011111111",
  8786=>"100000100",
  8787=>"011001000",
  8788=>"111100000",
  8789=>"000100110",
  8790=>"100100111",
  8791=>"101000000",
  8792=>"011000111",
  8793=>"000100101",
  8794=>"100100100",
  8795=>"000011000",
  8796=>"000000000",
  8797=>"000001001",
  8798=>"111111100",
  8799=>"100110001",
  8800=>"000011011",
  8801=>"000010110",
  8802=>"111000001",
  8803=>"001000100",
  8804=>"000000001",
  8805=>"111111111",
  8806=>"110011111",
  8807=>"100011001",
  8808=>"000011101",
  8809=>"101100111",
  8810=>"000111110",
  8811=>"101111110",
  8812=>"000011011",
  8813=>"100100111",
  8814=>"000111011",
  8815=>"111100111",
  8816=>"100101001",
  8817=>"010011111",
  8818=>"001101110",
  8819=>"111111001",
  8820=>"011111000",
  8821=>"100000010",
  8822=>"000000011",
  8823=>"000011010",
  8824=>"100100111",
  8825=>"011010010",
  8826=>"001000101",
  8827=>"011000101",
  8828=>"011000001",
  8829=>"000110000",
  8830=>"110011110",
  8831=>"100011111",
  8832=>"000000000",
  8833=>"010010010",
  8834=>"001011011",
  8835=>"101111111",
  8836=>"000110000",
  8837=>"000011001",
  8838=>"001001001",
  8839=>"000100101",
  8840=>"000111111",
  8841=>"011101101",
  8842=>"111101111",
  8843=>"011011000",
  8844=>"000011011",
  8845=>"000110111",
  8846=>"111000101",
  8847=>"101001001",
  8848=>"000000100",
  8849=>"100110011",
  8850=>"110000000",
  8851=>"100111100",
  8852=>"000010100",
  8853=>"000000000",
  8854=>"111101101",
  8855=>"001011011",
  8856=>"011000000",
  8857=>"000011011",
  8858=>"111100100",
  8859=>"010111100",
  8860=>"011100101",
  8861=>"000000000",
  8862=>"001010100",
  8863=>"000000000",
  8864=>"000100100",
  8865=>"110100110",
  8866=>"000011001",
  8867=>"011111011",
  8868=>"011011001",
  8869=>"100111010",
  8870=>"110011000",
  8871=>"000100101",
  8872=>"111000111",
  8873=>"000011001",
  8874=>"110100100",
  8875=>"100100100",
  8876=>"101111111",
  8877=>"000000000",
  8878=>"001011101",
  8879=>"111111010",
  8880=>"000010100",
  8881=>"110101101",
  8882=>"000001000",
  8883=>"011000000",
  8884=>"000111010",
  8885=>"000100100",
  8886=>"000000111",
  8887=>"010001101",
  8888=>"111000001",
  8889=>"100010000",
  8890=>"000010100",
  8891=>"011111011",
  8892=>"101000100",
  8893=>"001111111",
  8894=>"011111001",
  8895=>"000000011",
  8896=>"000100000",
  8897=>"011000000",
  8898=>"000011011",
  8899=>"010010010",
  8900=>"000100100",
  8901=>"000110100",
  8902=>"000011011",
  8903=>"000100111",
  8904=>"011000100",
  8905=>"011111011",
  8906=>"001101111",
  8907=>"011000000",
  8908=>"100101101",
  8909=>"110101000",
  8910=>"100100000",
  8911=>"111000100",
  8912=>"000000010",
  8913=>"000110001",
  8914=>"011111001",
  8915=>"101100100",
  8916=>"000000000",
  8917=>"111100110",
  8918=>"000010011",
  8919=>"000001011",
  8920=>"100110100",
  8921=>"000000101",
  8922=>"011110100",
  8923=>"111100100",
  8924=>"000010000",
  8925=>"000011011",
  8926=>"000011001",
  8927=>"000000100",
  8928=>"111100011",
  8929=>"111100100",
  8930=>"111100000",
  8931=>"000010010",
  8932=>"101100110",
  8933=>"010011011",
  8934=>"000010111",
  8935=>"011001110",
  8936=>"110110111",
  8937=>"100000000",
  8938=>"001000100",
  8939=>"010100100",
  8940=>"001011011",
  8941=>"100100111",
  8942=>"000000000",
  8943=>"010011110",
  8944=>"000000100",
  8945=>"000001001",
  8946=>"011011000",
  8947=>"010111000",
  8948=>"001011001",
  8949=>"101000100",
  8950=>"000100000",
  8951=>"011001000",
  8952=>"011100111",
  8953=>"000100110",
  8954=>"100100010",
  8955=>"000000010",
  8956=>"111100100",
  8957=>"000000000",
  8958=>"100111001",
  8959=>"101100101",
  8960=>"011010000",
  8961=>"000111010",
  8962=>"111000110",
  8963=>"110111111",
  8964=>"101111111",
  8965=>"111001000",
  8966=>"110101000",
  8967=>"000110101",
  8968=>"000100110",
  8969=>"000000100",
  8970=>"110100100",
  8971=>"100000000",
  8972=>"000111111",
  8973=>"010100010",
  8974=>"011011110",
  8975=>"111111000",
  8976=>"111111111",
  8977=>"100100100",
  8978=>"000101101",
  8979=>"111101000",
  8980=>"101111110",
  8981=>"000111000",
  8982=>"011000111",
  8983=>"100000100",
  8984=>"000101001",
  8985=>"111010111",
  8986=>"000101110",
  8987=>"000000111",
  8988=>"100101111",
  8989=>"000111110",
  8990=>"011000100",
  8991=>"100101101",
  8992=>"111101000",
  8993=>"111111110",
  8994=>"010010000",
  8995=>"010100000",
  8996=>"001001011",
  8997=>"111010000",
  8998=>"111000101",
  8999=>"001000000",
  9000=>"100101111",
  9001=>"001011000",
  9002=>"111101100",
  9003=>"111000000",
  9004=>"011111111",
  9005=>"111010000",
  9006=>"101111100",
  9007=>"100001001",
  9008=>"010100110",
  9009=>"111010011",
  9010=>"000010000",
  9011=>"000011010",
  9012=>"010101001",
  9013=>"001110100",
  9014=>"001000000",
  9015=>"111000111",
  9016=>"111000000",
  9017=>"101001100",
  9018=>"010010000",
  9019=>"001000000",
  9020=>"101000100",
  9021=>"111111100",
  9022=>"010000101",
  9023=>"110111000",
  9024=>"000110111",
  9025=>"111000000",
  9026=>"111111111",
  9027=>"101100000",
  9028=>"110101010",
  9029=>"000110100",
  9030=>"001000101",
  9031=>"011101000",
  9032=>"000101111",
  9033=>"000001010",
  9034=>"000000101",
  9035=>"000000000",
  9036=>"111001111",
  9037=>"000010110",
  9038=>"011011011",
  9039=>"111111110",
  9040=>"110000101",
  9041=>"111000000",
  9042=>"111101000",
  9043=>"011000000",
  9044=>"111001011",
  9045=>"011010110",
  9046=>"010011011",
  9047=>"000000111",
  9048=>"010111011",
  9049=>"111000011",
  9050=>"111101100",
  9051=>"100000101",
  9052=>"001101001",
  9053=>"001001010",
  9054=>"000111110",
  9055=>"100000000",
  9056=>"111101000",
  9057=>"101111001",
  9058=>"101000111",
  9059=>"011001001",
  9060=>"111110100",
  9061=>"001000000",
  9062=>"110111111",
  9063=>"001001001",
  9064=>"011010000",
  9065=>"100101001",
  9066=>"000010111",
  9067=>"000101000",
  9068=>"111111100",
  9069=>"000010000",
  9070=>"000000000",
  9071=>"000010000",
  9072=>"000001110",
  9073=>"111000101",
  9074=>"000000000",
  9075=>"000000110",
  9076=>"110000000",
  9077=>"001000100",
  9078=>"000111110",
  9079=>"111111000",
  9080=>"010110111",
  9081=>"101101101",
  9082=>"000010110",
  9083=>"000001000",
  9084=>"100110011",
  9085=>"010000100",
  9086=>"000000111",
  9087=>"000001001",
  9088=>"000010000",
  9089=>"111100101",
  9090=>"100101000",
  9091=>"001010010",
  9092=>"100100000",
  9093=>"000000100",
  9094=>"011001100",
  9095=>"001011011",
  9096=>"011011011",
  9097=>"000000000",
  9098=>"111111001",
  9099=>"100011000",
  9100=>"111110010",
  9101=>"010100010",
  9102=>"110001100",
  9103=>"000000010",
  9104=>"111000101",
  9105=>"110111000",
  9106=>"101000111",
  9107=>"000000111",
  9108=>"000010111",
  9109=>"000000101",
  9110=>"111101010",
  9111=>"000010100",
  9112=>"110100000",
  9113=>"111110100",
  9114=>"111000111",
  9115=>"001100110",
  9116=>"111101111",
  9117=>"000000100",
  9118=>"010110110",
  9119=>"111000110",
  9120=>"000010011",
  9121=>"001100000",
  9122=>"111011010",
  9123=>"011000000",
  9124=>"101010000",
  9125=>"010110100",
  9126=>"000111010",
  9127=>"010001111",
  9128=>"111000000",
  9129=>"001001111",
  9130=>"000100000",
  9131=>"011000101",
  9132=>"000010101",
  9133=>"100001101",
  9134=>"110000101",
  9135=>"111010010",
  9136=>"010010010",
  9137=>"110101100",
  9138=>"110010111",
  9139=>"000001000",
  9140=>"000011011",
  9141=>"111111100",
  9142=>"111100000",
  9143=>"010011000",
  9144=>"000000001",
  9145=>"000110110",
  9146=>"101000000",
  9147=>"010010111",
  9148=>"000010000",
  9149=>"110111110",
  9150=>"001001010",
  9151=>"011100101",
  9152=>"000000010",
  9153=>"111111111",
  9154=>"000000100",
  9155=>"000001100",
  9156=>"000000000",
  9157=>"011111101",
  9158=>"000000000",
  9159=>"001101111",
  9160=>"000000000",
  9161=>"111101000",
  9162=>"111101000",
  9163=>"000011010",
  9164=>"111000100",
  9165=>"011000011",
  9166=>"010000111",
  9167=>"111000000",
  9168=>"100100000",
  9169=>"110000111",
  9170=>"100111111",
  9171=>"111111111",
  9172=>"101101111",
  9173=>"101000110",
  9174=>"111000000",
  9175=>"001001111",
  9176=>"001000110",
  9177=>"000111010",
  9178=>"101000010",
  9179=>"111000000",
  9180=>"010100111",
  9181=>"010101100",
  9182=>"111111000",
  9183=>"000011101",
  9184=>"010010011",
  9185=>"000100111",
  9186=>"101001000",
  9187=>"000110110",
  9188=>"100100111",
  9189=>"101000000",
  9190=>"101101111",
  9191=>"001001011",
  9192=>"111010000",
  9193=>"101111111",
  9194=>"110010001",
  9195=>"001110010",
  9196=>"010111110",
  9197=>"000000000",
  9198=>"000100000",
  9199=>"101110000",
  9200=>"000100000",
  9201=>"111111111",
  9202=>"010000011",
  9203=>"000100000",
  9204=>"011111100",
  9205=>"101001101",
  9206=>"000000010",
  9207=>"001000011",
  9208=>"000010010",
  9209=>"000000000",
  9210=>"001010110",
  9211=>"000101111",
  9212=>"001000100",
  9213=>"001011011",
  9214=>"010010011",
  9215=>"011100111",
  9216=>"000000001",
  9217=>"100111111",
  9218=>"100000100",
  9219=>"000000101",
  9220=>"111100000",
  9221=>"000000000",
  9222=>"111000101",
  9223=>"010111110",
  9224=>"101100100",
  9225=>"010110110",
  9226=>"010111010",
  9227=>"100000101",
  9228=>"000000000",
  9229=>"010000011",
  9230=>"001001001",
  9231=>"111010000",
  9232=>"111000010",
  9233=>"110010000",
  9234=>"010000000",
  9235=>"111001000",
  9236=>"000000000",
  9237=>"000000000",
  9238=>"000000011",
  9239=>"010011111",
  9240=>"001100000",
  9241=>"110111101",
  9242=>"000111100",
  9243=>"011111000",
  9244=>"000000011",
  9245=>"011110000",
  9246=>"111000010",
  9247=>"111111010",
  9248=>"111111101",
  9249=>"100111010",
  9250=>"000011011",
  9251=>"000011010",
  9252=>"110010011",
  9253=>"000000000",
  9254=>"100000101",
  9255=>"000001000",
  9256=>"011010111",
  9257=>"000000101",
  9258=>"001000000",
  9259=>"011101000",
  9260=>"011011010",
  9261=>"000101111",
  9262=>"000101111",
  9263=>"110100101",
  9264=>"000101111",
  9265=>"001111111",
  9266=>"111011010",
  9267=>"111000000",
  9268=>"111110110",
  9269=>"000000111",
  9270=>"000111110",
  9271=>"000000111",
  9272=>"000110000",
  9273=>"101001101",
  9274=>"100000100",
  9275=>"000101011",
  9276=>"000110101",
  9277=>"100111010",
  9278=>"100000101",
  9279=>"101110010",
  9280=>"111000000",
  9281=>"010000000",
  9282=>"000000111",
  9283=>"111111100",
  9284=>"101101111",
  9285=>"000000000",
  9286=>"000101111",
  9287=>"111110101",
  9288=>"001100000",
  9289=>"101011111",
  9290=>"111101000",
  9291=>"100000000",
  9292=>"110000010",
  9293=>"111100010",
  9294=>"111001111",
  9295=>"111101111",
  9296=>"010110111",
  9297=>"010111010",
  9298=>"111010101",
  9299=>"001000100",
  9300=>"010000000",
  9301=>"000000100",
  9302=>"011011000",
  9303=>"111101000",
  9304=>"110000010",
  9305=>"100100111",
  9306=>"001000000",
  9307=>"100100000",
  9308=>"000111111",
  9309=>"001001011",
  9310=>"001111000",
  9311=>"110111101",
  9312=>"111111000",
  9313=>"010111011",
  9314=>"111111000",
  9315=>"100100000",
  9316=>"101001100",
  9317=>"100001110",
  9318=>"111111000",
  9319=>"001011111",
  9320=>"101001101",
  9321=>"111111000",
  9322=>"000111111",
  9323=>"101000001",
  9324=>"000000111",
  9325=>"010010000",
  9326=>"000000111",
  9327=>"101000111",
  9328=>"100100100",
  9329=>"000101000",
  9330=>"010111011",
  9331=>"111011101",
  9332=>"101011111",
  9333=>"000000000",
  9334=>"000001001",
  9335=>"010000000",
  9336=>"001011000",
  9337=>"010010000",
  9338=>"000011001",
  9339=>"000000101",
  9340=>"100110010",
  9341=>"100000000",
  9342=>"000000000",
  9343=>"101001100",
  9344=>"111000101",
  9345=>"011000010",
  9346=>"110100110",
  9347=>"000000101",
  9348=>"111111111",
  9349=>"000000100",
  9350=>"010000010",
  9351=>"000110000",
  9352=>"001001001",
  9353=>"010010111",
  9354=>"101000100",
  9355=>"111101100",
  9356=>"000000100",
  9357=>"010000000",
  9358=>"000000100",
  9359=>"100000000",
  9360=>"011110001",
  9361=>"000100000",
  9362=>"010111000",
  9363=>"111000000",
  9364=>"000011111",
  9365=>"110011000",
  9366=>"111000000",
  9367=>"001001111",
  9368=>"111111010",
  9369=>"000111011",
  9370=>"111111111",
  9371=>"011001110",
  9372=>"101000000",
  9373=>"111111000",
  9374=>"000000101",
  9375=>"010010111",
  9376=>"000101101",
  9377=>"111000100",
  9378=>"110000000",
  9379=>"010000111",
  9380=>"000000011",
  9381=>"111101000",
  9382=>"010110000",
  9383=>"000010010",
  9384=>"110111111",
  9385=>"000111111",
  9386=>"111000000",
  9387=>"111010000",
  9388=>"011010000",
  9389=>"101101111",
  9390=>"010000100",
  9391=>"000000111",
  9392=>"000000010",
  9393=>"111011001",
  9394=>"100000000",
  9395=>"000000110",
  9396=>"110110010",
  9397=>"011101000",
  9398=>"011011001",
  9399=>"000000101",
  9400=>"100011000",
  9401=>"100111111",
  9402=>"000000000",
  9403=>"000111100",
  9404=>"000110111",
  9405=>"010010010",
  9406=>"001001000",
  9407=>"011110000",
  9408=>"000000101",
  9409=>"000100111",
  9410=>"000111111",
  9411=>"100000100",
  9412=>"011000001",
  9413=>"110110111",
  9414=>"000100100",
  9415=>"000000111",
  9416=>"111000001",
  9417=>"000110000",
  9418=>"100111111",
  9419=>"111101011",
  9420=>"101100101",
  9421=>"001111110",
  9422=>"111111011",
  9423=>"111111100",
  9424=>"000000000",
  9425=>"010110111",
  9426=>"011000101",
  9427=>"111111010",
  9428=>"000000111",
  9429=>"110110010",
  9430=>"100000110",
  9431=>"000111111",
  9432=>"000000101",
  9433=>"110100111",
  9434=>"000100100",
  9435=>"000010010",
  9436=>"000001000",
  9437=>"011010000",
  9438=>"111111001",
  9439=>"111111000",
  9440=>"000000101",
  9441=>"000000001",
  9442=>"001000000",
  9443=>"010000111",
  9444=>"111000000",
  9445=>"100000000",
  9446=>"010000111",
  9447=>"011000101",
  9448=>"000111111",
  9449=>"000111111",
  9450=>"000001000",
  9451=>"000000001",
  9452=>"000100000",
  9453=>"111101111",
  9454=>"000000000",
  9455=>"001010110",
  9456=>"111011010",
  9457=>"011001001",
  9458=>"000000111",
  9459=>"001001001",
  9460=>"110010011",
  9461=>"110000111",
  9462=>"000000111",
  9463=>"000001001",
  9464=>"010111010",
  9465=>"001000101",
  9466=>"000000000",
  9467=>"101011111",
  9468=>"111111110",
  9469=>"000000011",
  9470=>"011011010",
  9471=>"000000101",
  9472=>"010001000",
  9473=>"111011111",
  9474=>"100000101",
  9475=>"110000001",
  9476=>"000100100",
  9477=>"000011000",
  9478=>"010000010",
  9479=>"001010010",
  9480=>"110011000",
  9481=>"000100100",
  9482=>"001001001",
  9483=>"000010000",
  9484=>"000000000",
  9485=>"011111010",
  9486=>"000110001",
  9487=>"101000111",
  9488=>"000000000",
  9489=>"000000111",
  9490=>"000000000",
  9491=>"111111110",
  9492=>"001000001",
  9493=>"100000101",
  9494=>"111000100",
  9495=>"010010111",
  9496=>"000000000",
  9497=>"100001110",
  9498=>"101100100",
  9499=>"000000111",
  9500=>"000000111",
  9501=>"000100000",
  9502=>"110010000",
  9503=>"010010010",
  9504=>"101101110",
  9505=>"111110100",
  9506=>"100111011",
  9507=>"101000011",
  9508=>"100100100",
  9509=>"010010111",
  9510=>"000011010",
  9511=>"100100111",
  9512=>"100100100",
  9513=>"001010000",
  9514=>"000001000",
  9515=>"100000111",
  9516=>"000001011",
  9517=>"010011101",
  9518=>"100000000",
  9519=>"000101000",
  9520=>"010001000",
  9521=>"110100000",
  9522=>"001000111",
  9523=>"000000111",
  9524=>"000000100",
  9525=>"010101110",
  9526=>"011111000",
  9527=>"000000001",
  9528=>"111000100",
  9529=>"000110000",
  9530=>"000110010",
  9531=>"101101111",
  9532=>"000011111",
  9533=>"101111000",
  9534=>"111000001",
  9535=>"111111101",
  9536=>"101100111",
  9537=>"111101111",
  9538=>"111111000",
  9539=>"011011011",
  9540=>"111111111",
  9541=>"000000100",
  9542=>"000000000",
  9543=>"000100000",
  9544=>"010011001",
  9545=>"000000001",
  9546=>"010000001",
  9547=>"111000000",
  9548=>"001000000",
  9549=>"001001001",
  9550=>"111111110",
  9551=>"111001111",
  9552=>"111111111",
  9553=>"000110111",
  9554=>"000000000",
  9555=>"110000000",
  9556=>"111110101",
  9557=>"000001000",
  9558=>"100100111",
  9559=>"000000000",
  9560=>"100000010",
  9561=>"001011000",
  9562=>"000011000",
  9563=>"010111110",
  9564=>"000000100",
  9565=>"001001010",
  9566=>"111111110",
  9567=>"110100100",
  9568=>"100000000",
  9569=>"111101111",
  9570=>"100000000",
  9571=>"000001111",
  9572=>"111111100",
  9573=>"011011000",
  9574=>"101101111",
  9575=>"001111010",
  9576=>"010010000",
  9577=>"101000111",
  9578=>"000010111",
  9579=>"101000100",
  9580=>"001000000",
  9581=>"000101011",
  9582=>"101000111",
  9583=>"011011011",
  9584=>"001011001",
  9585=>"000010111",
  9586=>"001110100",
  9587=>"111111011",
  9588=>"100101111",
  9589=>"100000111",
  9590=>"101011111",
  9591=>"111111111",
  9592=>"000001111",
  9593=>"010000011",
  9594=>"111000101",
  9595=>"000000100",
  9596=>"110011101",
  9597=>"110100100",
  9598=>"001001010",
  9599=>"001000000",
  9600=>"111011010",
  9601=>"100100000",
  9602=>"111111011",
  9603=>"111111111",
  9604=>"111100100",
  9605=>"100001111",
  9606=>"100010110",
  9607=>"001001101",
  9608=>"001110000",
  9609=>"111011001",
  9610=>"000100100",
  9611=>"111000000",
  9612=>"010111000",
  9613=>"000000000",
  9614=>"000000000",
  9615=>"000000101",
  9616=>"100110110",
  9617=>"100101101",
  9618=>"110001111",
  9619=>"111111000",
  9620=>"000110100",
  9621=>"100111101",
  9622=>"111011000",
  9623=>"000011010",
  9624=>"111110000",
  9625=>"111111111",
  9626=>"111111010",
  9627=>"101000000",
  9628=>"000011011",
  9629=>"101101111",
  9630=>"100111111",
  9631=>"000000000",
  9632=>"001101010",
  9633=>"000100111",
  9634=>"011000010",
  9635=>"110010011",
  9636=>"100100111",
  9637=>"101111111",
  9638=>"001001101",
  9639=>"011111110",
  9640=>"000001011",
  9641=>"100100111",
  9642=>"101000000",
  9643=>"000000000",
  9644=>"011011001",
  9645=>"111110000",
  9646=>"001101001",
  9647=>"011010101",
  9648=>"000000000",
  9649=>"110110100",
  9650=>"111011000",
  9651=>"101111001",
  9652=>"100100111",
  9653=>"011110000",
  9654=>"101100010",
  9655=>"101000011",
  9656=>"001110011",
  9657=>"000110100",
  9658=>"010111011",
  9659=>"111010100",
  9660=>"111110110",
  9661=>"000000000",
  9662=>"011111100",
  9663=>"000110010",
  9664=>"000101111",
  9665=>"101101001",
  9666=>"110110111",
  9667=>"001001111",
  9668=>"100001011",
  9669=>"100111001",
  9670=>"101101100",
  9671=>"000011000",
  9672=>"000011010",
  9673=>"000010010",
  9674=>"110000100",
  9675=>"101101111",
  9676=>"111111111",
  9677=>"001011000",
  9678=>"000000011",
  9679=>"111000000",
  9680=>"111111011",
  9681=>"010110111",
  9682=>"000000101",
  9683=>"101100000",
  9684=>"000000110",
  9685=>"011011011",
  9686=>"111010000",
  9687=>"111110000",
  9688=>"111111010",
  9689=>"010000000",
  9690=>"110101101",
  9691=>"101000100",
  9692=>"001001000",
  9693=>"100000000",
  9694=>"110111111",
  9695=>"111011000",
  9696=>"111011000",
  9697=>"000000101",
  9698=>"100000010",
  9699=>"011111101",
  9700=>"000100111",
  9701=>"011100011",
  9702=>"000000011",
  9703=>"100101011",
  9704=>"100000000",
  9705=>"101111111",
  9706=>"100100101",
  9707=>"100101111",
  9708=>"110110000",
  9709=>"000000000",
  9710=>"000000000",
  9711=>"000000010",
  9712=>"000000110",
  9713=>"101010000",
  9714=>"100000010",
  9715=>"000011100",
  9716=>"010100000",
  9717=>"111111101",
  9718=>"000000000",
  9719=>"011100111",
  9720=>"101100100",
  9721=>"000000100",
  9722=>"100100010",
  9723=>"000000000",
  9724=>"111010000",
  9725=>"111100101",
  9726=>"100100100",
  9727=>"111000000",
  9728=>"011100000",
  9729=>"000000101",
  9730=>"000001000",
  9731=>"000111111",
  9732=>"011111100",
  9733=>"000001111",
  9734=>"000111101",
  9735=>"010010010",
  9736=>"000000000",
  9737=>"010010000",
  9738=>"110111011",
  9739=>"000001000",
  9740=>"000000100",
  9741=>"000000000",
  9742=>"100110100",
  9743=>"001111111",
  9744=>"001101000",
  9745=>"111100101",
  9746=>"000000000",
  9747=>"111000110",
  9748=>"111111111",
  9749=>"111000001",
  9750=>"000000111",
  9751=>"111000101",
  9752=>"000000000",
  9753=>"000101111",
  9754=>"001000000",
  9755=>"000000101",
  9756=>"111111001",
  9757=>"000000000",
  9758=>"111101000",
  9759=>"100000000",
  9760=>"111000011",
  9761=>"001000000",
  9762=>"010100110",
  9763=>"000000000",
  9764=>"001111110",
  9765=>"011011001",
  9766=>"010011011",
  9767=>"000111101",
  9768=>"010000000",
  9769=>"110000000",
  9770=>"111111101",
  9771=>"111110000",
  9772=>"110101100",
  9773=>"100000001",
  9774=>"011001000",
  9775=>"000110110",
  9776=>"010000000",
  9777=>"000011001",
  9778=>"000110011",
  9779=>"110000111",
  9780=>"111110000",
  9781=>"110111111",
  9782=>"000000001",
  9783=>"101010110",
  9784=>"111111010",
  9785=>"000000111",
  9786=>"010111000",
  9787=>"000101111",
  9788=>"100111110",
  9789=>"111111111",
  9790=>"100000100",
  9791=>"011111101",
  9792=>"100000000",
  9793=>"000000101",
  9794=>"111100110",
  9795=>"000011011",
  9796=>"111001101",
  9797=>"111110000",
  9798=>"010111111",
  9799=>"111010000",
  9800=>"000001111",
  9801=>"101001000",
  9802=>"101001111",
  9803=>"110110111",
  9804=>"111000000",
  9805=>"000110110",
  9806=>"010011010",
  9807=>"111111111",
  9808=>"111000000",
  9809=>"110110111",
  9810=>"100111001",
  9811=>"001000000",
  9812=>"000000010",
  9813=>"001000000",
  9814=>"000011111",
  9815=>"010111000",
  9816=>"001010000",
  9817=>"000010011",
  9818=>"111011011",
  9819=>"110010010",
  9820=>"011001000",
  9821=>"010010110",
  9822=>"000001000",
  9823=>"100110000",
  9824=>"100101100",
  9825=>"010011111",
  9826=>"111111111",
  9827=>"100100111",
  9828=>"000000000",
  9829=>"000010100",
  9830=>"000101100",
  9831=>"111111010",
  9832=>"000111111",
  9833=>"010000001",
  9834=>"111111110",
  9835=>"111111000",
  9836=>"111111110",
  9837=>"101111101",
  9838=>"101011011",
  9839=>"101000111",
  9840=>"010111110",
  9841=>"010000000",
  9842=>"000000000",
  9843=>"110010010",
  9844=>"111101000",
  9845=>"000000100",
  9846=>"000111111",
  9847=>"110001000",
  9848=>"011011010",
  9849=>"000111001",
  9850=>"000000111",
  9851=>"000000100",
  9852=>"000100110",
  9853=>"101000000",
  9854=>"011111000",
  9855=>"000001001",
  9856=>"001000000",
  9857=>"111100100",
  9858=>"111111000",
  9859=>"000100111",
  9860=>"111010011",
  9861=>"100111000",
  9862=>"110100100",
  9863=>"000110010",
  9864=>"000111111",
  9865=>"000000001",
  9866=>"010010000",
  9867=>"011011000",
  9868=>"000110000",
  9869=>"111110111",
  9870=>"010010000",
  9871=>"100000000",
  9872=>"011111011",
  9873=>"111111111",
  9874=>"001001101",
  9875=>"111000011",
  9876=>"000000000",
  9877=>"000100000",
  9878=>"100010010",
  9879=>"100100100",
  9880=>"111111000",
  9881=>"111000011",
  9882=>"000111000",
  9883=>"011010110",
  9884=>"100000000",
  9885=>"101000110",
  9886=>"110111110",
  9887=>"100101101",
  9888=>"000100001",
  9889=>"111000000",
  9890=>"000111000",
  9891=>"000010000",
  9892=>"110000111",
  9893=>"100011000",
  9894=>"000111111",
  9895=>"010101000",
  9896=>"000000001",
  9897=>"000000000",
  9898=>"100111000",
  9899=>"111110000",
  9900=>"011110110",
  9901=>"111000000",
  9902=>"111000001",
  9903=>"110111111",
  9904=>"000101111",
  9905=>"000000000",
  9906=>"100010010",
  9907=>"000110111",
  9908=>"011111111",
  9909=>"010010111",
  9910=>"111000000",
  9911=>"001001000",
  9912=>"000111111",
  9913=>"001000010",
  9914=>"111111101",
  9915=>"111101100",
  9916=>"111000000",
  9917=>"111111111",
  9918=>"100100000",
  9919=>"010000000",
  9920=>"010000000",
  9921=>"000000000",
  9922=>"110000100",
  9923=>"001011000",
  9924=>"000000000",
  9925=>"111000000",
  9926=>"111011110",
  9927=>"000010111",
  9928=>"100111100",
  9929=>"101000100",
  9930=>"111111000",
  9931=>"111100111",
  9932=>"101001000",
  9933=>"000011111",
  9934=>"111010000",
  9935=>"100111111",
  9936=>"001011111",
  9937=>"011110111",
  9938=>"000110111",
  9939=>"000111100",
  9940=>"100000011",
  9941=>"111110000",
  9942=>"000000000",
  9943=>"110000100",
  9944=>"111001000",
  9945=>"010111111",
  9946=>"100100110",
  9947=>"011000000",
  9948=>"000000111",
  9949=>"111111111",
  9950=>"100111101",
  9951=>"111110100",
  9952=>"000000000",
  9953=>"001000111",
  9954=>"000010010",
  9955=>"111111111",
  9956=>"100000000",
  9957=>"011001010",
  9958=>"101100000",
  9959=>"111000100",
  9960=>"100111111",
  9961=>"111111111",
  9962=>"011111110",
  9963=>"001000000",
  9964=>"111100100",
  9965=>"111001001",
  9966=>"001011001",
  9967=>"000000000",
  9968=>"011111000",
  9969=>"111001100",
  9970=>"111001001",
  9971=>"100100100",
  9972=>"110111011",
  9973=>"000100111",
  9974=>"100101000",
  9975=>"010111111",
  9976=>"000000111",
  9977=>"111000000",
  9978=>"001101101",
  9979=>"000101101",
  9980=>"111110111",
  9981=>"011000000",
  9982=>"000111100",
  9983=>"101101111",
  9984=>"001011011",
  9985=>"111111000",
  9986=>"111001000",
  9987=>"110111101",
  9988=>"000100100",
  9989=>"101001000",
  9990=>"000000000",
  9991=>"000000101",
  9992=>"000110110",
  9993=>"000100101",
  9994=>"110000100",
  9995=>"101001001",
  9996=>"111111101",
  9997=>"000010111",
  9998=>"000100100",
  9999=>"101111110",
  10000=>"010001000",
  10001=>"111000000",
  10002=>"110101001",
  10003=>"101000010",
  10004=>"000100111",
  10005=>"001000000",
  10006=>"011111001",
  10007=>"111111101",
  10008=>"101101111",
  10009=>"000001011",
  10010=>"000000000",
  10011=>"000101100",
  10012=>"111001011",
  10013=>"001001101",
  10014=>"110110000",
  10015=>"000010110",
  10016=>"111000101",
  10017=>"001101000",
  10018=>"101000010",
  10019=>"001110111",
  10020=>"111111110",
  10021=>"110110100",
  10022=>"101000001",
  10023=>"100011111",
  10024=>"101101111",
  10025=>"111001001",
  10026=>"001000001",
  10027=>"010010111",
  10028=>"100100100",
  10029=>"000101101",
  10030=>"000000000",
  10031=>"101100110",
  10032=>"011001100",
  10033=>"100100100",
  10034=>"011010000",
  10035=>"101000000",
  10036=>"110101001",
  10037=>"000111010",
  10038=>"000100100",
  10039=>"011011000",
  10040=>"111111000",
  10041=>"010010000",
  10042=>"000100000",
  10043=>"010000000",
  10044=>"000110010",
  10045=>"111111111",
  10046=>"000000000",
  10047=>"000111111",
  10048=>"110111101",
  10049=>"111111000",
  10050=>"011111110",
  10051=>"010111011",
  10052=>"010000110",
  10053=>"010000110",
  10054=>"000111001",
  10055=>"111000000",
  10056=>"100000100",
  10057=>"111111111",
  10058=>"000000000",
  10059=>"000001000",
  10060=>"101101101",
  10061=>"011111111",
  10062=>"010011011",
  10063=>"000000000",
  10064=>"000000000",
  10065=>"111111111",
  10066=>"111101010",
  10067=>"011011011",
  10068=>"100100110",
  10069=>"001011010",
  10070=>"000011101",
  10071=>"111000000",
  10072=>"000000101",
  10073=>"000110110",
  10074=>"010001100",
  10075=>"000111100",
  10076=>"000010000",
  10077=>"000000000",
  10078=>"000010111",
  10079=>"111100100",
  10080=>"000110111",
  10081=>"111000001",
  10082=>"100101110",
  10083=>"000001001",
  10084=>"000010011",
  10085=>"000010111",
  10086=>"000001111",
  10087=>"000010010",
  10088=>"001101000",
  10089=>"111111001",
  10090=>"110111111",
  10091=>"010110000",
  10092=>"111000101",
  10093=>"101001101",
  10094=>"000010000",
  10095=>"010100000",
  10096=>"000010111",
  10097=>"111111100",
  10098=>"010001001",
  10099=>"111001000",
  10100=>"000011111",
  10101=>"010101111",
  10102=>"000111110",
  10103=>"000000111",
  10104=>"101000000",
  10105=>"010111111",
  10106=>"111111111",
  10107=>"111000000",
  10108=>"001011010",
  10109=>"000110000",
  10110=>"100000111",
  10111=>"101101111",
  10112=>"111010111",
  10113=>"111111110",
  10114=>"000000111",
  10115=>"000000000",
  10116=>"000000110",
  10117=>"110110100",
  10118=>"111111111",
  10119=>"000000000",
  10120=>"000111111",
  10121=>"000000000",
  10122=>"000100101",
  10123=>"110111000",
  10124=>"111000111",
  10125=>"000000000",
  10126=>"000010111",
  10127=>"111001001",
  10128=>"000110100",
  10129=>"000111110",
  10130=>"000101101",
  10131=>"011000111",
  10132=>"000000000",
  10133=>"111011000",
  10134=>"111111111",
  10135=>"000000011",
  10136=>"011011000",
  10137=>"010000000",
  10138=>"111101000",
  10139=>"011000111",
  10140=>"000010000",
  10141=>"101111111",
  10142=>"111011000",
  10143=>"111111001",
  10144=>"000011011",
  10145=>"010000001",
  10146=>"011111101",
  10147=>"111000000",
  10148=>"000001000",
  10149=>"000110110",
  10150=>"110110100",
  10151=>"000010110",
  10152=>"111101010",
  10153=>"001010111",
  10154=>"111111111",
  10155=>"111111001",
  10156=>"101111110",
  10157=>"000111011",
  10158=>"100100100",
  10159=>"111000000",
  10160=>"001011001",
  10161=>"001000100",
  10162=>"000010010",
  10163=>"000011000",
  10164=>"101011101",
  10165=>"011010000",
  10166=>"010111110",
  10167=>"010110010",
  10168=>"011011010",
  10169=>"000000000",
  10170=>"010110100",
  10171=>"000110100",
  10172=>"110000011",
  10173=>"101101111",
  10174=>"000111111",
  10175=>"111000000",
  10176=>"010110110",
  10177=>"010010000",
  10178=>"010100100",
  10179=>"111011011",
  10180=>"000001101",
  10181=>"111101010",
  10182=>"111111010",
  10183=>"010000010",
  10184=>"001000101",
  10185=>"001010110",
  10186=>"000000110",
  10187=>"000111111",
  10188=>"000000111",
  10189=>"000100111",
  10190=>"010111111",
  10191=>"111000010",
  10192=>"110001001",
  10193=>"010011000",
  10194=>"000000111",
  10195=>"010111101",
  10196=>"001001000",
  10197=>"000000000",
  10198=>"110110100",
  10199=>"111110000",
  10200=>"001001010",
  10201=>"101000011",
  10202=>"000111000",
  10203=>"111000000",
  10204=>"100111110",
  10205=>"101000000",
  10206=>"000111101",
  10207=>"111110111",
  10208=>"101001110",
  10209=>"000000000",
  10210=>"101011111",
  10211=>"000000001",
  10212=>"111001101",
  10213=>"000000110",
  10214=>"111001000",
  10215=>"010011001",
  10216=>"111111111",
  10217=>"000000100",
  10218=>"001000000",
  10219=>"111010100",
  10220=>"001000000",
  10221=>"000001111",
  10222=>"000100001",
  10223=>"000110010",
  10224=>"111000111",
  10225=>"011111111",
  10226=>"011111000",
  10227=>"000011111",
  10228=>"000110110",
  10229=>"111000101",
  10230=>"111000000",
  10231=>"001100111",
  10232=>"000010010",
  10233=>"101010110",
  10234=>"111101000",
  10235=>"000000001",
  10236=>"000000010",
  10237=>"000000000",
  10238=>"000011001",
  10239=>"111000000",
  10240=>"001001011",
  10241=>"100101100",
  10242=>"101000001",
  10243=>"101111100",
  10244=>"011011111",
  10245=>"000000000",
  10246=>"000000001",
  10247=>"101110110",
  10248=>"110111000",
  10249=>"000101101",
  10250=>"001000100",
  10251=>"111000000",
  10252=>"111001101",
  10253=>"110100111",
  10254=>"110111001",
  10255=>"000000110",
  10256=>"110010010",
  10257=>"100101101",
  10258=>"000000101",
  10259=>"111010000",
  10260=>"101010100",
  10261=>"110000000",
  10262=>"011100100",
  10263=>"111001000",
  10264=>"111110000",
  10265=>"111110111",
  10266=>"000000001",
  10267=>"001101111",
  10268=>"000111001",
  10269=>"001111011",
  10270=>"000000000",
  10271=>"000000101",
  10272=>"111110000",
  10273=>"010010110",
  10274=>"000000000",
  10275=>"010111000",
  10276=>"100101100",
  10277=>"100100100",
  10278=>"111010000",
  10279=>"001000000",
  10280=>"010011000",
  10281=>"100111111",
  10282=>"010000000",
  10283=>"000000000",
  10284=>"111001011",
  10285=>"111010101",
  10286=>"100101110",
  10287=>"000000000",
  10288=>"000010000",
  10289=>"011000000",
  10290=>"000010011",
  10291=>"001000010",
  10292=>"000000101",
  10293=>"111000010",
  10294=>"000000000",
  10295=>"011111010",
  10296=>"111010000",
  10297=>"111100100",
  10298=>"110110010",
  10299=>"100000000",
  10300=>"000010110",
  10301=>"011011010",
  10302=>"100101111",
  10303=>"110011010",
  10304=>"000011111",
  10305=>"111000000",
  10306=>"111111100",
  10307=>"110110000",
  10308=>"101001000",
  10309=>"101010010",
  10310=>"000101101",
  10311=>"111111111",
  10312=>"110010001",
  10313=>"000010011",
  10314=>"101010000",
  10315=>"010111100",
  10316=>"000101000",
  10317=>"001101010",
  10318=>"100000101",
  10319=>"000000011",
  10320=>"000000101",
  10321=>"111000111",
  10322=>"110111000",
  10323=>"011101000",
  10324=>"001101111",
  10325=>"000100001",
  10326=>"011011000",
  10327=>"100000111",
  10328=>"000001111",
  10329=>"001011000",
  10330=>"000101101",
  10331=>"100011000",
  10332=>"101000000",
  10333=>"000001111",
  10334=>"111101111",
  10335=>"110011011",
  10336=>"100000000",
  10337=>"001000010",
  10338=>"000000000",
  10339=>"110000101",
  10340=>"111110010",
  10341=>"000100110",
  10342=>"000100110",
  10343=>"111111110",
  10344=>"101000110",
  10345=>"111000000",
  10346=>"000111111",
  10347=>"110000001",
  10348=>"000111010",
  10349=>"010110111",
  10350=>"000000011",
  10351=>"111111000",
  10352=>"001101000",
  10353=>"100010000",
  10354=>"000000000",
  10355=>"000000001",
  10356=>"111111101",
  10357=>"101100100",
  10358=>"000110111",
  10359=>"010111000",
  10360=>"011011010",
  10361=>"000100111",
  10362=>"011000101",
  10363=>"111111010",
  10364=>"100110111",
  10365=>"100101100",
  10366=>"111001010",
  10367=>"111000000",
  10368=>"111100000",
  10369=>"110111111",
  10370=>"010111000",
  10371=>"000111111",
  10372=>"000000111",
  10373=>"000001100",
  10374=>"001001000",
  10375=>"100011001",
  10376=>"100100000",
  10377=>"000000101",
  10378=>"100000000",
  10379=>"101111000",
  10380=>"010010000",
  10381=>"101001111",
  10382=>"101111000",
  10383=>"001000101",
  10384=>"100011001",
  10385=>"011001000",
  10386=>"111000100",
  10387=>"000010111",
  10388=>"000101001",
  10389=>"010010010",
  10390=>"111011000",
  10391=>"001001000",
  10392=>"100111100",
  10393=>"100110111",
  10394=>"000000101",
  10395=>"000000101",
  10396=>"111111101",
  10397=>"000101010",
  10398=>"111000111",
  10399=>"000100010",
  10400=>"101011111",
  10401=>"000000011",
  10402=>"111111111",
  10403=>"111110111",
  10404=>"010101110",
  10405=>"100110000",
  10406=>"100110001",
  10407=>"001111111",
  10408=>"111100000",
  10409=>"000010111",
  10410=>"111010110",
  10411=>"111111000",
  10412=>"010111000",
  10413=>"110000000",
  10414=>"000001101",
  10415=>"111101111",
  10416=>"010010001",
  10417=>"000100010",
  10418=>"111111110",
  10419=>"001110110",
  10420=>"000001000",
  10421=>"000001000",
  10422=>"111011011",
  10423=>"001000100",
  10424=>"000010011",
  10425=>"000111110",
  10426=>"111101111",
  10427=>"000000000",
  10428=>"010000000",
  10429=>"011010010",
  10430=>"011011000",
  10431=>"101000000",
  10432=>"101000000",
  10433=>"100000101",
  10434=>"010000000",
  10435=>"111001001",
  10436=>"011000100",
  10437=>"001001000",
  10438=>"111111000",
  10439=>"111111101",
  10440=>"011111100",
  10441=>"000101111",
  10442=>"111111100",
  10443=>"000000000",
  10444=>"000111111",
  10445=>"000011111",
  10446=>"000010010",
  10447=>"111111000",
  10448=>"000000011",
  10449=>"000110011",
  10450=>"101011111",
  10451=>"000011111",
  10452=>"000001010",
  10453=>"000000000",
  10454=>"101000000",
  10455=>"000111110",
  10456=>"111000000",
  10457=>"000000101",
  10458=>"000001010",
  10459=>"000000000",
  10460=>"001111100",
  10461=>"111111100",
  10462=>"100000100",
  10463=>"101111111",
  10464=>"001000000",
  10465=>"000000111",
  10466=>"000101111",
  10467=>"101001100",
  10468=>"111000011",
  10469=>"101000000",
  10470=>"011011111",
  10471=>"100100111",
  10472=>"000001111",
  10473=>"001011111",
  10474=>"100000000",
  10475=>"011010001",
  10476=>"000111000",
  10477=>"101000000",
  10478=>"000000000",
  10479=>"110000000",
  10480=>"010010000",
  10481=>"001011100",
  10482=>"010000000",
  10483=>"000100100",
  10484=>"100101011",
  10485=>"111000111",
  10486=>"000000100",
  10487=>"010001001",
  10488=>"000011010",
  10489=>"110010111",
  10490=>"111111101",
  10491=>"000000000",
  10492=>"010111000",
  10493=>"000000011",
  10494=>"100111111",
  10495=>"000111101",
  10496=>"100100100",
  10497=>"011010000",
  10498=>"000000000",
  10499=>"000000000",
  10500=>"100000011",
  10501=>"001011101",
  10502=>"111111001",
  10503=>"101111111",
  10504=>"001001001",
  10505=>"000000000",
  10506=>"111111111",
  10507=>"010110001",
  10508=>"001001100",
  10509=>"000000100",
  10510=>"010110111",
  10511=>"101111111",
  10512=>"111010011",
  10513=>"111111110",
  10514=>"111010010",
  10515=>"111111111",
  10516=>"111110111",
  10517=>"111111111",
  10518=>"001000010",
  10519=>"010111110",
  10520=>"110000101",
  10521=>"111011011",
  10522=>"101000111",
  10523=>"000000000",
  10524=>"011111111",
  10525=>"001111111",
  10526=>"000000011",
  10527=>"000010010",
  10528=>"000001001",
  10529=>"000000000",
  10530=>"000000010",
  10531=>"000000000",
  10532=>"110111000",
  10533=>"011001001",
  10534=>"010010011",
  10535=>"000000000",
  10536=>"000011111",
  10537=>"001110000",
  10538=>"111111111",
  10539=>"110111100",
  10540=>"110010000",
  10541=>"111000001",
  10542=>"001100010",
  10543=>"101101000",
  10544=>"100000000",
  10545=>"001000000",
  10546=>"001111000",
  10547=>"111111111",
  10548=>"111111111",
  10549=>"110101011",
  10550=>"111111111",
  10551=>"001111111",
  10552=>"110010101",
  10553=>"111010111",
  10554=>"011000111",
  10555=>"011000000",
  10556=>"000001011",
  10557=>"111011011",
  10558=>"000001001",
  10559=>"001000011",
  10560=>"111111110",
  10561=>"000000011",
  10562=>"000000000",
  10563=>"000101100",
  10564=>"000000000",
  10565=>"001011101",
  10566=>"101111000",
  10567=>"000101111",
  10568=>"110000000",
  10569=>"000000000",
  10570=>"011111101",
  10571=>"111111011",
  10572=>"111111111",
  10573=>"111111001",
  10574=>"100100000",
  10575=>"000000010",
  10576=>"111111111",
  10577=>"111011110",
  10578=>"111001000",
  10579=>"000100100",
  10580=>"100001000",
  10581=>"001000000",
  10582=>"000001011",
  10583=>"000000001",
  10584=>"011011111",
  10585=>"001110110",
  10586=>"111111111",
  10587=>"100111111",
  10588=>"110011001",
  10589=>"000000110",
  10590=>"001100001",
  10591=>"001011101",
  10592=>"111111111",
  10593=>"000000101",
  10594=>"111111111",
  10595=>"101100000",
  10596=>"000000000",
  10597=>"111111111",
  10598=>"000001111",
  10599=>"000001011",
  10600=>"000000000",
  10601=>"111101111",
  10602=>"111111111",
  10603=>"010111111",
  10604=>"011000000",
  10605=>"111111111",
  10606=>"000000000",
  10607=>"111110111",
  10608=>"110111110",
  10609=>"111111111",
  10610=>"111111111",
  10611=>"000111111",
  10612=>"000111111",
  10613=>"010111111",
  10614=>"000110010",
  10615=>"000010110",
  10616=>"000001101",
  10617=>"110000000",
  10618=>"110111111",
  10619=>"000000000",
  10620=>"011001001",
  10621=>"001001001",
  10622=>"000011000",
  10623=>"000000010",
  10624=>"000000101",
  10625=>"111111101",
  10626=>"000001000",
  10627=>"000001000",
  10628=>"101101111",
  10629=>"000111111",
  10630=>"011100010",
  10631=>"111010010",
  10632=>"111111000",
  10633=>"001000111",
  10634=>"000100001",
  10635=>"000111110",
  10636=>"100110000",
  10637=>"001101000",
  10638=>"101111011",
  10639=>"000000101",
  10640=>"111111111",
  10641=>"111111110",
  10642=>"111001000",
  10643=>"000101111",
  10644=>"000100111",
  10645=>"001011111",
  10646=>"111111001",
  10647=>"000011010",
  10648=>"000100100",
  10649=>"000111001",
  10650=>"000110110",
  10651=>"000000001",
  10652=>"101000100",
  10653=>"110110000",
  10654=>"100000101",
  10655=>"011000010",
  10656=>"000000000",
  10657=>"111000000",
  10658=>"000000000",
  10659=>"111000000",
  10660=>"111111111",
  10661=>"111011111",
  10662=>"000000111",
  10663=>"000000000",
  10664=>"111000000",
  10665=>"000000000",
  10666=>"111111111",
  10667=>"111111111",
  10668=>"001000111",
  10669=>"111000111",
  10670=>"011011011",
  10671=>"001000001",
  10672=>"000001101",
  10673=>"101111110",
  10674=>"001010010",
  10675=>"000110110",
  10676=>"010110111",
  10677=>"011110000",
  10678=>"011000000",
  10679=>"110111000",
  10680=>"000000110",
  10681=>"011111100",
  10682=>"000001111",
  10683=>"110111000",
  10684=>"000000001",
  10685=>"000110010",
  10686=>"000000001",
  10687=>"000000000",
  10688=>"001001110",
  10689=>"110111010",
  10690=>"100000101",
  10691=>"110110110",
  10692=>"110000000",
  10693=>"110111001",
  10694=>"010000000",
  10695=>"000000111",
  10696=>"000000101",
  10697=>"000001001",
  10698=>"110111001",
  10699=>"110110000",
  10700=>"011111011",
  10701=>"111110111",
  10702=>"010110111",
  10703=>"011110001",
  10704=>"010010010",
  10705=>"000000011",
  10706=>"000010010",
  10707=>"111111010",
  10708=>"000011011",
  10709=>"011011000",
  10710=>"000000001",
  10711=>"111111111",
  10712=>"011001000",
  10713=>"000000000",
  10714=>"000000000",
  10715=>"111110111",
  10716=>"000000000",
  10717=>"000000000",
  10718=>"111111111",
  10719=>"010011111",
  10720=>"001000000",
  10721=>"111111110",
  10722=>"001001101",
  10723=>"111111100",
  10724=>"101001001",
  10725=>"111111111",
  10726=>"000000111",
  10727=>"101010000",
  10728=>"000000010",
  10729=>"010001001",
  10730=>"111111111",
  10731=>"111101111",
  10732=>"111001001",
  10733=>"111111111",
  10734=>"111110000",
  10735=>"000000001",
  10736=>"000100111",
  10737=>"111111000",
  10738=>"000000000",
  10739=>"000000111",
  10740=>"000001000",
  10741=>"111111111",
  10742=>"110111111",
  10743=>"000001111",
  10744=>"000000110",
  10745=>"001000000",
  10746=>"000111100",
  10747=>"001110110",
  10748=>"111111010",
  10749=>"000101001",
  10750=>"011110110",
  10751=>"111111010",
  10752=>"011001101",
  10753=>"000000011",
  10754=>"001000001",
  10755=>"010111000",
  10756=>"111111101",
  10757=>"111111111",
  10758=>"111111001",
  10759=>"100000000",
  10760=>"011111111",
  10761=>"010010000",
  10762=>"110110100",
  10763=>"101111111",
  10764=>"000000000",
  10765=>"111011111",
  10766=>"111011110",
  10767=>"000000000",
  10768=>"111000110",
  10769=>"010000000",
  10770=>"000000111",
  10771=>"001001000",
  10772=>"101111100",
  10773=>"111101001",
  10774=>"011101101",
  10775=>"111111010",
  10776=>"000000000",
  10777=>"111111111",
  10778=>"100100000",
  10779=>"010011111",
  10780=>"010010111",
  10781=>"000000010",
  10782=>"111111000",
  10783=>"000000000",
  10784=>"000010100",
  10785=>"001110111",
  10786=>"000011111",
  10787=>"101111110",
  10788=>"000100100",
  10789=>"100100100",
  10790=>"001111010",
  10791=>"110110110",
  10792=>"111111010",
  10793=>"110111100",
  10794=>"000000000",
  10795=>"001110010",
  10796=>"000011001",
  10797=>"111111110",
  10798=>"100000000",
  10799=>"010000011",
  10800=>"000001000",
  10801=>"000000001",
  10802=>"111111111",
  10803=>"010000001",
  10804=>"011111110",
  10805=>"000010000",
  10806=>"011000000",
  10807=>"000000000",
  10808=>"101000000",
  10809=>"000000000",
  10810=>"000010011",
  10811=>"010000010",
  10812=>"001100011",
  10813=>"000000101",
  10814=>"000000000",
  10815=>"100110111",
  10816=>"000001101",
  10817=>"001000000",
  10818=>"010110111",
  10819=>"011011100",
  10820=>"000010000",
  10821=>"000001001",
  10822=>"000010000",
  10823=>"011000101",
  10824=>"100011011",
  10825=>"111111111",
  10826=>"111001001",
  10827=>"001100100",
  10828=>"000000000",
  10829=>"001001001",
  10830=>"001001100",
  10831=>"000000101",
  10832=>"000000000",
  10833=>"100100110",
  10834=>"111111100",
  10835=>"001000000",
  10836=>"000000000",
  10837=>"000000111",
  10838=>"011101111",
  10839=>"110010110",
  10840=>"000000101",
  10841=>"000000001",
  10842=>"000100000",
  10843=>"001000111",
  10844=>"000010000",
  10845=>"000110001",
  10846=>"010000000",
  10847=>"100101011",
  10848=>"111110010",
  10849=>"001111111",
  10850=>"110010010",
  10851=>"010010111",
  10852=>"000000001",
  10853=>"111111111",
  10854=>"111111111",
  10855=>"110110111",
  10856=>"111111111",
  10857=>"111111011",
  10858=>"000000100",
  10859=>"111111111",
  10860=>"001100111",
  10861=>"111111111",
  10862=>"111000000",
  10863=>"000000101",
  10864=>"100100100",
  10865=>"001001000",
  10866=>"110000000",
  10867=>"111110110",
  10868=>"001000101",
  10869=>"000000000",
  10870=>"111010101",
  10871=>"000000000",
  10872=>"000000000",
  10873=>"000000000",
  10874=>"000111111",
  10875=>"111111111",
  10876=>"011110111",
  10877=>"110100000",
  10878=>"111110110",
  10879=>"101111001",
  10880=>"000010101",
  10881=>"111101100",
  10882=>"001111011",
  10883=>"000000000",
  10884=>"101001000",
  10885=>"111110110",
  10886=>"001011001",
  10887=>"000001001",
  10888=>"011011010",
  10889=>"011000001",
  10890=>"101111010",
  10891=>"110010000",
  10892=>"101000100",
  10893=>"110110100",
  10894=>"000001000",
  10895=>"000000000",
  10896=>"110100100",
  10897=>"111000000",
  10898=>"001000001",
  10899=>"001110111",
  10900=>"001000011",
  10901=>"111000110",
  10902=>"010000000",
  10903=>"000000000",
  10904=>"110000000",
  10905=>"111111111",
  10906=>"100100100",
  10907=>"110000000",
  10908=>"111111000",
  10909=>"000000011",
  10910=>"111000000",
  10911=>"001010000",
  10912=>"000111101",
  10913=>"010010110",
  10914=>"000010111",
  10915=>"110001000",
  10916=>"000000110",
  10917=>"000000001",
  10918=>"000111001",
  10919=>"100100000",
  10920=>"111111011",
  10921=>"100101000",
  10922=>"001010011",
  10923=>"111001111",
  10924=>"111100111",
  10925=>"001001101",
  10926=>"100110011",
  10927=>"000111100",
  10928=>"011110100",
  10929=>"000100101",
  10930=>"010110010",
  10931=>"000000100",
  10932=>"101101101",
  10933=>"111111110",
  10934=>"101000000",
  10935=>"110111111",
  10936=>"000000110",
  10937=>"000000100",
  10938=>"010000001",
  10939=>"111101011",
  10940=>"000000000",
  10941=>"111000100",
  10942=>"111111110",
  10943=>"111001001",
  10944=>"111111111",
  10945=>"000000000",
  10946=>"110000000",
  10947=>"001001000",
  10948=>"111110010",
  10949=>"100010011",
  10950=>"101000010",
  10951=>"011111111",
  10952=>"010111110",
  10953=>"000000000",
  10954=>"111011100",
  10955=>"000100000",
  10956=>"000000000",
  10957=>"000001110",
  10958=>"000000100",
  10959=>"000001001",
  10960=>"101000000",
  10961=>"011111000",
  10962=>"000100001",
  10963=>"011000000",
  10964=>"000000000",
  10965=>"001011111",
  10966=>"111111000",
  10967=>"110000010",
  10968=>"000000111",
  10969=>"100100000",
  10970=>"000111001",
  10971=>"000000000",
  10972=>"110000100",
  10973=>"000101110",
  10974=>"101000000",
  10975=>"110000000",
  10976=>"011001001",
  10977=>"000110110",
  10978=>"101110111",
  10979=>"111111111",
  10980=>"111000000",
  10981=>"000010000",
  10982=>"101011111",
  10983=>"010010100",
  10984=>"001001110",
  10985=>"100010000",
  10986=>"011111011",
  10987=>"010111110",
  10988=>"000000000",
  10989=>"111001110",
  10990=>"000000000",
  10991=>"000000000",
  10992=>"101000000",
  10993=>"001110100",
  10994=>"001000001",
  10995=>"000000100",
  10996=>"100000001",
  10997=>"111111111",
  10998=>"010000000",
  10999=>"000000001",
  11000=>"000001000",
  11001=>"111111000",
  11002=>"100110110",
  11003=>"000010111",
  11004=>"010100111",
  11005=>"000111000",
  11006=>"001001001",
  11007=>"011101001",
  11008=>"011001001",
  11009=>"000000101",
  11010=>"101000001",
  11011=>"000110011",
  11012=>"011011101",
  11013=>"000000000",
  11014=>"111000000",
  11015=>"011001011",
  11016=>"000000000",
  11017=>"010111000",
  11018=>"000000000",
  11019=>"000000111",
  11020=>"101111111",
  11021=>"000100110",
  11022=>"011110001",
  11023=>"000000000",
  11024=>"111000000",
  11025=>"110111010",
  11026=>"000001000",
  11027=>"000001111",
  11028=>"111111000",
  11029=>"101001000",
  11030=>"100100001",
  11031=>"000111111",
  11032=>"111000101",
  11033=>"111001101",
  11034=>"010011001",
  11035=>"010010110",
  11036=>"000000101",
  11037=>"000001001",
  11038=>"111100001",
  11039=>"000111110",
  11040=>"000000001",
  11041=>"111111011",
  11042=>"000110010",
  11043=>"111111111",
  11044=>"001011011",
  11045=>"100111011",
  11046=>"110110110",
  11047=>"111111000",
  11048=>"010010000",
  11049=>"110110001",
  11050=>"100110000",
  11051=>"010000000",
  11052=>"001111101",
  11053=>"101111111",
  11054=>"111000000",
  11055=>"000001010",
  11056=>"111111111",
  11057=>"011011000",
  11058=>"001101101",
  11059=>"101001001",
  11060=>"100000100",
  11061=>"000110000",
  11062=>"000000011",
  11063=>"010000111",
  11064=>"111111111",
  11065=>"000000100",
  11066=>"000001000",
  11067=>"010100000",
  11068=>"110000001",
  11069=>"111111000",
  11070=>"000100100",
  11071=>"001111100",
  11072=>"111001011",
  11073=>"110010101",
  11074=>"001101101",
  11075=>"100011001",
  11076=>"000000111",
  11077=>"001000000",
  11078=>"000101000",
  11079=>"001001110",
  11080=>"000001111",
  11081=>"111111000",
  11082=>"000111111",
  11083=>"111101110",
  11084=>"110111000",
  11085=>"100100100",
  11086=>"110110100",
  11087=>"111011110",
  11088=>"000000110",
  11089=>"111111010",
  11090=>"001000101",
  11091=>"001001000",
  11092=>"010010000",
  11093=>"100100001",
  11094=>"100110111",
  11095=>"110111001",
  11096=>"101101101",
  11097=>"100001000",
  11098=>"100111110",
  11099=>"010000010",
  11100=>"010000000",
  11101=>"001001000",
  11102=>"101011011",
  11103=>"010100000",
  11104=>"111111111",
  11105=>"010011001",
  11106=>"011000001",
  11107=>"001001101",
  11108=>"000101001",
  11109=>"001001010",
  11110=>"110110000",
  11111=>"011111000",
  11112=>"011010111",
  11113=>"111001000",
  11114=>"111100111",
  11115=>"001111111",
  11116=>"000110111",
  11117=>"000011010",
  11118=>"000001111",
  11119=>"111001111",
  11120=>"111111100",
  11121=>"000111111",
  11122=>"011100100",
  11123=>"101101000",
  11124=>"010000000",
  11125=>"000000001",
  11126=>"000111111",
  11127=>"110111000",
  11128=>"000000111",
  11129=>"001111111",
  11130=>"000000111",
  11131=>"101101100",
  11132=>"000110000",
  11133=>"100100000",
  11134=>"010011001",
  11135=>"010000000",
  11136=>"111010010",
  11137=>"111110000",
  11138=>"111001001",
  11139=>"100100111",
  11140=>"111000000",
  11141=>"101111101",
  11142=>"011101100",
  11143=>"100001001",
  11144=>"011001000",
  11145=>"001010110",
  11146=>"000000000",
  11147=>"111001000",
  11148=>"000000000",
  11149=>"011000000",
  11150=>"111001110",
  11151=>"000000101",
  11152=>"111101111",
  11153=>"000110110",
  11154=>"010010000",
  11155=>"000000110",
  11156=>"000000000",
  11157=>"000000000",
  11158=>"111111111",
  11159=>"011011000",
  11160=>"010110111",
  11161=>"000101111",
  11162=>"000001011",
  11163=>"010000000",
  11164=>"100000000",
  11165=>"101000100",
  11166=>"111000000",
  11167=>"000000010",
  11168=>"110100110",
  11169=>"000000111",
  11170=>"111101100",
  11171=>"101111101",
  11172=>"010000001",
  11173=>"001000101",
  11174=>"010110000",
  11175=>"000000101",
  11176=>"111000001",
  11177=>"100111000",
  11178=>"000011010",
  11179=>"001000000",
  11180=>"001001011",
  11181=>"110000100",
  11182=>"010000110",
  11183=>"000000001",
  11184=>"000001111",
  11185=>"011101101",
  11186=>"000000000",
  11187=>"111001001",
  11188=>"100111011",
  11189=>"001111111",
  11190=>"000111110",
  11191=>"000110000",
  11192=>"000100100",
  11193=>"001110110",
  11194=>"010000010",
  11195=>"000010111",
  11196=>"011110011",
  11197=>"111101000",
  11198=>"100000000",
  11199=>"000000110",
  11200=>"000001111",
  11201=>"010010000",
  11202=>"111110111",
  11203=>"100100000",
  11204=>"111111000",
  11205=>"010110111",
  11206=>"000110111",
  11207=>"010010000",
  11208=>"101111111",
  11209=>"000010000",
  11210=>"111101000",
  11211=>"000000111",
  11212=>"010000000",
  11213=>"001011001",
  11214=>"001100101",
  11215=>"000000000",
  11216=>"000000000",
  11217=>"001111010",
  11218=>"001110011",
  11219=>"100000011",
  11220=>"110111000",
  11221=>"101001101",
  11222=>"111110000",
  11223=>"000000000",
  11224=>"000101111",
  11225=>"111000111",
  11226=>"011011000",
  11227=>"111000000",
  11228=>"011001000",
  11229=>"011111011",
  11230=>"101101101",
  11231=>"011001000",
  11232=>"010010000",
  11233=>"000000001",
  11234=>"010111000",
  11235=>"110100000",
  11236=>"111111000",
  11237=>"010010111",
  11238=>"101011100",
  11239=>"001001001",
  11240=>"111111000",
  11241=>"101111011",
  11242=>"000110001",
  11243=>"111111011",
  11244=>"111000000",
  11245=>"000111111",
  11246=>"111000000",
  11247=>"100000110",
  11248=>"101111011",
  11249=>"001001010",
  11250=>"010010000",
  11251=>"000101111",
  11252=>"110100100",
  11253=>"101000101",
  11254=>"000100000",
  11255=>"000000100",
  11256=>"000000000",
  11257=>"011000100",
  11258=>"111100111",
  11259=>"000101000",
  11260=>"000001111",
  11261=>"000000100",
  11262=>"100100110",
  11263=>"111000110",
  11264=>"000111100",
  11265=>"101111000",
  11266=>"100000100",
  11267=>"100110010",
  11268=>"000011001",
  11269=>"000000111",
  11270=>"000000000",
  11271=>"000011110",
  11272=>"111011000",
  11273=>"100000000",
  11274=>"000110100",
  11275=>"111101101",
  11276=>"111000000",
  11277=>"111101000",
  11278=>"000110001",
  11279=>"001000000",
  11280=>"000100111",
  11281=>"111000111",
  11282=>"110110100",
  11283=>"000000010",
  11284=>"010111111",
  11285=>"000010111",
  11286=>"011011111",
  11287=>"111000101",
  11288=>"101000000",
  11289=>"110010010",
  11290=>"000011001",
  11291=>"110111000",
  11292=>"100111101",
  11293=>"111001000",
  11294=>"000011010",
  11295=>"001000000",
  11296=>"000111000",
  11297=>"000111111",
  11298=>"100101111",
  11299=>"000000111",
  11300=>"011001001",
  11301=>"011111101",
  11302=>"000111111",
  11303=>"011110011",
  11304=>"100100000",
  11305=>"000010010",
  11306=>"000000000",
  11307=>"101110000",
  11308=>"110011011",
  11309=>"111111001",
  11310=>"000111111",
  11311=>"110111001",
  11312=>"100000101",
  11313=>"011100001",
  11314=>"111100000",
  11315=>"000111111",
  11316=>"000111111",
  11317=>"100000111",
  11318=>"001000001",
  11319=>"111100001",
  11320=>"010111111",
  11321=>"000000010",
  11322=>"111111110",
  11323=>"010010000",
  11324=>"110110110",
  11325=>"111111111",
  11326=>"000000101",
  11327=>"000000100",
  11328=>"001000000",
  11329=>"100011000",
  11330=>"111111111",
  11331=>"000000100",
  11332=>"000111111",
  11333=>"000000000",
  11334=>"001000000",
  11335=>"000000111",
  11336=>"111111001",
  11337=>"101111011",
  11338=>"111000000",
  11339=>"101111111",
  11340=>"000111011",
  11341=>"000100110",
  11342=>"000011111",
  11343=>"000000000",
  11344=>"001011001",
  11345=>"111111100",
  11346=>"000000011",
  11347=>"011001011",
  11348=>"000100110",
  11349=>"110111111",
  11350=>"110100100",
  11351=>"100000011",
  11352=>"000001001",
  11353=>"010110110",
  11354=>"100110100",
  11355=>"000100110",
  11356=>"000111010",
  11357=>"000001000",
  11358=>"110010110",
  11359=>"000000001",
  11360=>"000000111",
  11361=>"000001011",
  11362=>"000000000",
  11363=>"000001011",
  11364=>"001110000",
  11365=>"010100000",
  11366=>"000111110",
  11367=>"111111100",
  11368=>"000110010",
  11369=>"100100000",
  11370=>"111110100",
  11371=>"000010100",
  11372=>"000010111",
  11373=>"000000101",
  11374=>"010000101",
  11375=>"111011000",
  11376=>"100111111",
  11377=>"111111101",
  11378=>"110100110",
  11379=>"100000111",
  11380=>"111111100",
  11381=>"001000001",
  11382=>"001011000",
  11383=>"000000000",
  11384=>"111100000",
  11385=>"001111000",
  11386=>"111001111",
  11387=>"000110111",
  11388=>"001110111",
  11389=>"111000000",
  11390=>"000100111",
  11391=>"000000101",
  11392=>"110101110",
  11393=>"111001001",
  11394=>"000000001",
  11395=>"101000010",
  11396=>"000010111",
  11397=>"111001100",
  11398=>"110111011",
  11399=>"000011010",
  11400=>"100111111",
  11401=>"101111100",
  11402=>"000010000",
  11403=>"000010001",
  11404=>"111000101",
  11405=>"111000100",
  11406=>"000011100",
  11407=>"011001011",
  11408=>"001011011",
  11409=>"011111111",
  11410=>"000000000",
  11411=>"000111111",
  11412=>"010010010",
  11413=>"101000000",
  11414=>"111100000",
  11415=>"000100000",
  11416=>"100000100",
  11417=>"110100011",
  11418=>"111000000",
  11419=>"000000000",
  11420=>"111111000",
  11421=>"010000011",
  11422=>"111011011",
  11423=>"101111110",
  11424=>"011001000",
  11425=>"111111101",
  11426=>"111101000",
  11427=>"010111001",
  11428=>"110111111",
  11429=>"110100000",
  11430=>"011001100",
  11431=>"100111111",
  11432=>"101010111",
  11433=>"001000111",
  11434=>"111100100",
  11435=>"000000111",
  11436=>"111100111",
  11437=>"000111111",
  11438=>"111111101",
  11439=>"101101110",
  11440=>"101000100",
  11441=>"010101101",
  11442=>"000000000",
  11443=>"000000000",
  11444=>"111000101",
  11445=>"111111101",
  11446=>"001110000",
  11447=>"110111110",
  11448=>"011011011",
  11449=>"001000110",
  11450=>"000011101",
  11451=>"110011010",
  11452=>"010011001",
  11453=>"111000101",
  11454=>"100100000",
  11455=>"011010101",
  11456=>"000010000",
  11457=>"110000000",
  11458=>"110010000",
  11459=>"000110110",
  11460=>"000011100",
  11461=>"000110111",
  11462=>"000000011",
  11463=>"101100100",
  11464=>"000101001",
  11465=>"001111100",
  11466=>"000010111",
  11467=>"111000111",
  11468=>"000010001",
  11469=>"001011011",
  11470=>"110010100",
  11471=>"111011100",
  11472=>"111100000",
  11473=>"111011011",
  11474=>"000011000",
  11475=>"000000000",
  11476=>"000000111",
  11477=>"110000100",
  11478=>"000011011",
  11479=>"100000011",
  11480=>"110011011",
  11481=>"000000001",
  11482=>"100101000",
  11483=>"111100101",
  11484=>"011110111",
  11485=>"101101110",
  11486=>"010111111",
  11487=>"000000000",
  11488=>"000000000",
  11489=>"101100100",
  11490=>"111101000",
  11491=>"101111101",
  11492=>"111000000",
  11493=>"000000100",
  11494=>"101101101",
  11495=>"010111100",
  11496=>"101111000",
  11497=>"110000000",
  11498=>"001111010",
  11499=>"100010111",
  11500=>"011000000",
  11501=>"111001001",
  11502=>"000000000",
  11503=>"101000000",
  11504=>"101100100",
  11505=>"011011011",
  11506=>"001001110",
  11507=>"010011111",
  11508=>"011111111",
  11509=>"101000001",
  11510=>"100000000",
  11511=>"010011100",
  11512=>"010011000",
  11513=>"001101011",
  11514=>"111111111",
  11515=>"000001011",
  11516=>"101000000",
  11517=>"000100000",
  11518=>"001100001",
  11519=>"001100101",
  11520=>"111110110",
  11521=>"111110011",
  11522=>"000000101",
  11523=>"011011001",
  11524=>"000001100",
  11525=>"000111111",
  11526=>"010010010",
  11527=>"000000000",
  11528=>"000010011",
  11529=>"100001000",
  11530=>"110001000",
  11531=>"111001011",
  11532=>"111001000",
  11533=>"000000010",
  11534=>"010110011",
  11535=>"000111110",
  11536=>"011011101",
  11537=>"101111111",
  11538=>"101110000",
  11539=>"001011000",
  11540=>"000100100",
  11541=>"100100100",
  11542=>"000110011",
  11543=>"101001101",
  11544=>"000000001",
  11545=>"100010110",
  11546=>"111111110",
  11547=>"000000110",
  11548=>"000100110",
  11549=>"111000110",
  11550=>"000100100",
  11551=>"010010000",
  11552=>"011000001",
  11553=>"011010110",
  11554=>"000000101",
  11555=>"101000111",
  11556=>"101011111",
  11557=>"000011011",
  11558=>"101000100",
  11559=>"111111111",
  11560=>"011101101",
  11561=>"101111111",
  11562=>"100000011",
  11563=>"110010010",
  11564=>"110011011",
  11565=>"000010010",
  11566=>"000000100",
  11567=>"000111111",
  11568=>"000000111",
  11569=>"000110010",
  11570=>"111111110",
  11571=>"000000101",
  11572=>"010111110",
  11573=>"010100011",
  11574=>"000001011",
  11575=>"110100111",
  11576=>"010000100",
  11577=>"000001000",
  11578=>"000111000",
  11579=>"000000000",
  11580=>"000001111",
  11581=>"111111111",
  11582=>"000100000",
  11583=>"100101000",
  11584=>"111011011",
  11585=>"000000101",
  11586=>"010100100",
  11587=>"000000110",
  11588=>"111111111",
  11589=>"000000101",
  11590=>"101001011",
  11591=>"111011111",
  11592=>"000111001",
  11593=>"001011001",
  11594=>"111111100",
  11595=>"111100000",
  11596=>"100100111",
  11597=>"000111111",
  11598=>"000011011",
  11599=>"001011111",
  11600=>"100000100",
  11601=>"111111111",
  11602=>"000000011",
  11603=>"110111001",
  11604=>"000100000",
  11605=>"001111111",
  11606=>"000100011",
  11607=>"000111111",
  11608=>"000011010",
  11609=>"000110011",
  11610=>"010010010",
  11611=>"010000110",
  11612=>"000011111",
  11613=>"010110000",
  11614=>"101000000",
  11615=>"101101011",
  11616=>"100100000",
  11617=>"000000000",
  11618=>"000111011",
  11619=>"011111000",
  11620=>"111111100",
  11621=>"000101010",
  11622=>"000010010",
  11623=>"000000000",
  11624=>"111010100",
  11625=>"000000000",
  11626=>"111111000",
  11627=>"111111111",
  11628=>"100100100",
  11629=>"000011010",
  11630=>"000010000",
  11631=>"100111000",
  11632=>"000110110",
  11633=>"111000000",
  11634=>"000110100",
  11635=>"000110110",
  11636=>"101000000",
  11637=>"010010011",
  11638=>"100111101",
  11639=>"100000000",
  11640=>"011011011",
  11641=>"001011010",
  11642=>"000011000",
  11643=>"111000111",
  11644=>"011101001",
  11645=>"011011000",
  11646=>"001001000",
  11647=>"000000110",
  11648=>"111110110",
  11649=>"000011110",
  11650=>"000011011",
  11651=>"111100100",
  11652=>"111010000",
  11653=>"111111111",
  11654=>"000110110",
  11655=>"000101110",
  11656=>"011011001",
  11657=>"111000000",
  11658=>"001011000",
  11659=>"111111111",
  11660=>"000000100",
  11661=>"101101000",
  11662=>"011000100",
  11663=>"111000001",
  11664=>"100100100",
  11665=>"000000000",
  11666=>"001011000",
  11667=>"110011000",
  11668=>"100000000",
  11669=>"000000111",
  11670=>"101100110",
  11671=>"110110101",
  11672=>"000100010",
  11673=>"010111110",
  11674=>"000010000",
  11675=>"111010110",
  11676=>"000000000",
  11677=>"111000000",
  11678=>"001001000",
  11679=>"110000000",
  11680=>"100110010",
  11681=>"011010110",
  11682=>"011101100",
  11683=>"111011110",
  11684=>"000111111",
  11685=>"101101111",
  11686=>"000000000",
  11687=>"000010011",
  11688=>"000100000",
  11689=>"111111101",
  11690=>"000000000",
  11691=>"000110111",
  11692=>"110100000",
  11693=>"100101000",
  11694=>"101001001",
  11695=>"110001000",
  11696=>"000100101",
  11697=>"001110110",
  11698=>"000000000",
  11699=>"001011110",
  11700=>"011001000",
  11701=>"110001100",
  11702=>"011011111",
  11703=>"001111011",
  11704=>"100100001",
  11705=>"000000001",
  11706=>"000011111",
  11707=>"000010000",
  11708=>"101101111",
  11709=>"000111111",
  11710=>"110110100",
  11711=>"000000100",
  11712=>"000111111",
  11713=>"000111011",
  11714=>"011000000",
  11715=>"001001001",
  11716=>"000101110",
  11717=>"000100100",
  11718=>"111111011",
  11719=>"111011000",
  11720=>"000100111",
  11721=>"100100100",
  11722=>"110101111",
  11723=>"100000100",
  11724=>"110100111",
  11725=>"110111011",
  11726=>"000111010",
  11727=>"111111000",
  11728=>"010100101",
  11729=>"101111110",
  11730=>"110110100",
  11731=>"100101111",
  11732=>"000000000",
  11733=>"010011011",
  11734=>"000111011",
  11735=>"110000000",
  11736=>"001101100",
  11737=>"100000000",
  11738=>"000001110",
  11739=>"111111111",
  11740=>"110111110",
  11741=>"110110111",
  11742=>"010111010",
  11743=>"000000010",
  11744=>"000100000",
  11745=>"010000001",
  11746=>"110111111",
  11747=>"110111011",
  11748=>"111000000",
  11749=>"101000101",
  11750=>"111011111",
  11751=>"000000100",
  11752=>"111011111",
  11753=>"101100000",
  11754=>"111101000",
  11755=>"101111111",
  11756=>"101111101",
  11757=>"000000111",
  11758=>"100111001",
  11759=>"110001111",
  11760=>"111101111",
  11761=>"111001000",
  11762=>"011100110",
  11763=>"011011010",
  11764=>"011011011",
  11765=>"111100110",
  11766=>"000010111",
  11767=>"000000000",
  11768=>"010111101",
  11769=>"001000000",
  11770=>"110010011",
  11771=>"111111000",
  11772=>"100000000",
  11773=>"101000100",
  11774=>"000111111",
  11775=>"111100100",
  11776=>"110111111",
  11777=>"000000000",
  11778=>"100000100",
  11779=>"000000001",
  11780=>"111101011",
  11781=>"001000101",
  11782=>"010110111",
  11783=>"000101101",
  11784=>"010010010",
  11785=>"001100111",
  11786=>"000000000",
  11787=>"000010100",
  11788=>"010110011",
  11789=>"000000100",
  11790=>"100000010",
  11791=>"000100000",
  11792=>"100001001",
  11793=>"000001101",
  11794=>"111011011",
  11795=>"000000111",
  11796=>"111100000",
  11797=>"010010010",
  11798=>"000000001",
  11799=>"000000001",
  11800=>"101000000",
  11801=>"111111110",
  11802=>"000000001",
  11803=>"111001000",
  11804=>"101111101",
  11805=>"001111111",
  11806=>"001101001",
  11807=>"111110111",
  11808=>"010010000",
  11809=>"000000000",
  11810=>"000010100",
  11811=>"000000000",
  11812=>"111011011",
  11813=>"110010011",
  11814=>"001111000",
  11815=>"000010111",
  11816=>"010010010",
  11817=>"001111101",
  11818=>"010000010",
  11819=>"000010010",
  11820=>"110111111",
  11821=>"111001111",
  11822=>"001001101",
  11823=>"010010111",
  11824=>"000111111",
  11825=>"001001111",
  11826=>"000010000",
  11827=>"111111011",
  11828=>"000001110",
  11829=>"000000000",
  11830=>"011010101",
  11831=>"101101001",
  11832=>"001100001",
  11833=>"100001101",
  11834=>"100111011",
  11835=>"000000000",
  11836=>"001001100",
  11837=>"111111100",
  11838=>"000101000",
  11839=>"110100101",
  11840=>"101101010",
  11841=>"110101111",
  11842=>"001101111",
  11843=>"110010011",
  11844=>"010101101",
  11845=>"000001001",
  11846=>"111111111",
  11847=>"000000000",
  11848=>"011000111",
  11849=>"110101000",
  11850=>"000101111",
  11851=>"001001101",
  11852=>"001000000",
  11853=>"111111111",
  11854=>"100100111",
  11855=>"010000001",
  11856=>"111111000",
  11857=>"110111111",
  11858=>"010011111",
  11859=>"111011011",
  11860=>"000100000",
  11861=>"111011110",
  11862=>"110010010",
  11863=>"101000101",
  11864=>"111111100",
  11865=>"011011110",
  11866=>"001000000",
  11867=>"100001001",
  11868=>"010111111",
  11869=>"011001110",
  11870=>"111110111",
  11871=>"011110110",
  11872=>"001101100",
  11873=>"111111000",
  11874=>"101100100",
  11875=>"000000000",
  11876=>"011000000",
  11877=>"110111111",
  11878=>"010010010",
  11879=>"101000010",
  11880=>"101001000",
  11881=>"001000101",
  11882=>"000000100",
  11883=>"000100101",
  11884=>"000101111",
  11885=>"010101111",
  11886=>"001000001",
  11887=>"111111010",
  11888=>"100100111",
  11889=>"000000111",
  11890=>"110110111",
  11891=>"111110111",
  11892=>"011011001",
  11893=>"000101001",
  11894=>"101111111",
  11895=>"100110111",
  11896=>"010111000",
  11897=>"000000000",
  11898=>"110011111",
  11899=>"111110100",
  11900=>"111010000",
  11901=>"110100010",
  11902=>"010110000",
  11903=>"110010010",
  11904=>"000001000",
  11905=>"110100000",
  11906=>"000000010",
  11907=>"000000000",
  11908=>"000101001",
  11909=>"111111111",
  11910=>"010110100",
  11911=>"011111010",
  11912=>"001110111",
  11913=>"000001101",
  11914=>"000000101",
  11915=>"100001001",
  11916=>"100111110",
  11917=>"011100000",
  11918=>"110010000",
  11919=>"101101000",
  11920=>"111111011",
  11921=>"011000000",
  11922=>"000001001",
  11923=>"000111011",
  11924=>"100000000",
  11925=>"000101101",
  11926=>"010111011",
  11927=>"100111110",
  11928=>"011000101",
  11929=>"010110101",
  11930=>"010010010",
  11931=>"010010000",
  11932=>"001000101",
  11933=>"000001000",
  11934=>"000001101",
  11935=>"101101110",
  11936=>"011011011",
  11937=>"000000000",
  11938=>"010111110",
  11939=>"000100110",
  11940=>"001101111",
  11941=>"110110111",
  11942=>"101001001",
  11943=>"010000101",
  11944=>"111000001",
  11945=>"000000000",
  11946=>"101101101",
  11947=>"101001001",
  11948=>"110100101",
  11949=>"110100011",
  11950=>"011000001",
  11951=>"000011011",
  11952=>"000000000",
  11953=>"110110101",
  11954=>"000101000",
  11955=>"100010011",
  11956=>"111011111",
  11957=>"100101101",
  11958=>"000101111",
  11959=>"001001000",
  11960=>"110100011",
  11961=>"100010011",
  11962=>"000000000",
  11963=>"111101111",
  11964=>"111111111",
  11965=>"111110101",
  11966=>"001000010",
  11967=>"000000001",
  11968=>"110011011",
  11969=>"011111011",
  11970=>"101000000",
  11971=>"010011111",
  11972=>"000010000",
  11973=>"001101100",
  11974=>"000000100",
  11975=>"100111111",
  11976=>"010010111",
  11977=>"101011010",
  11978=>"000000000",
  11979=>"011101110",
  11980=>"110010010",
  11981=>"111011011",
  11982=>"101101000",
  11983=>"101000000",
  11984=>"100101111",
  11985=>"110111111",
  11986=>"100000000",
  11987=>"110100110",
  11988=>"011010101",
  11989=>"000000001",
  11990=>"111110000",
  11991=>"000001101",
  11992=>"010010111",
  11993=>"000000000",
  11994=>"100110010",
  11995=>"101101101",
  11996=>"000111011",
  11997=>"001000101",
  11998=>"111010111",
  11999=>"100100111",
  12000=>"000000111",
  12001=>"001110101",
  12002=>"111110111",
  12003=>"001000111",
  12004=>"101001000",
  12005=>"001011010",
  12006=>"000010001",
  12007=>"000001000",
  12008=>"000000101",
  12009=>"010011111",
  12010=>"111001000",
  12011=>"111110011",
  12012=>"010010010",
  12013=>"000001101",
  12014=>"001101010",
  12015=>"000010010",
  12016=>"101000001",
  12017=>"100000001",
  12018=>"000000010",
  12019=>"110110110",
  12020=>"011011011",
  12021=>"010000101",
  12022=>"000101001",
  12023=>"011111111",
  12024=>"000001001",
  12025=>"000000101",
  12026=>"111011010",
  12027=>"000001001",
  12028=>"010111000",
  12029=>"111011011",
  12030=>"011010110",
  12031=>"111111111",
  12032=>"101100101",
  12033=>"000000000",
  12034=>"000000100",
  12035=>"000001101",
  12036=>"000011000",
  12037=>"010000101",
  12038=>"101111111",
  12039=>"010011101",
  12040=>"000001001",
  12041=>"111110100",
  12042=>"000011011",
  12043=>"000000010",
  12044=>"101000000",
  12045=>"001000000",
  12046=>"111111100",
  12047=>"011001010",
  12048=>"010111011",
  12049=>"011000000",
  12050=>"000011110",
  12051=>"010111101",
  12052=>"001100110",
  12053=>"111111000",
  12054=>"011011101",
  12055=>"000111111",
  12056=>"101000000",
  12057=>"111110000",
  12058=>"000000000",
  12059=>"000010110",
  12060=>"000000110",
  12061=>"000110111",
  12062=>"000000000",
  12063=>"000011010",
  12064=>"000100111",
  12065=>"000010110",
  12066=>"000001101",
  12067=>"100111111",
  12068=>"100100111",
  12069=>"110010111",
  12070=>"000011011",
  12071=>"000111000",
  12072=>"001011111",
  12073=>"111000111",
  12074=>"010100000",
  12075=>"101001000",
  12076=>"100110110",
  12077=>"010001000",
  12078=>"011110000",
  12079=>"111111111",
  12080=>"111100100",
  12081=>"010001111",
  12082=>"000101100",
  12083=>"000001001",
  12084=>"000000011",
  12085=>"111010000",
  12086=>"011011111",
  12087=>"000101001",
  12088=>"000000111",
  12089=>"000000010",
  12090=>"000001111",
  12091=>"000000110",
  12092=>"100100110",
  12093=>"110010010",
  12094=>"000000100",
  12095=>"111011011",
  12096=>"110111111",
  12097=>"001100111",
  12098=>"010111111",
  12099=>"011000110",
  12100=>"010011010",
  12101=>"000101101",
  12102=>"000101000",
  12103=>"001000111",
  12104=>"010011010",
  12105=>"101000000",
  12106=>"001111001",
  12107=>"011000000",
  12108=>"000000111",
  12109=>"011001001",
  12110=>"000110011",
  12111=>"000000011",
  12112=>"000101111",
  12113=>"111111010",
  12114=>"111111111",
  12115=>"011000001",
  12116=>"101000000",
  12117=>"010011011",
  12118=>"011111110",
  12119=>"001111011",
  12120=>"111100000",
  12121=>"000011111",
  12122=>"111101000",
  12123=>"000100100",
  12124=>"111000000",
  12125=>"011000000",
  12126=>"111111100",
  12127=>"100111111",
  12128=>"100100000",
  12129=>"111101010",
  12130=>"101000100",
  12131=>"001011101",
  12132=>"001000000",
  12133=>"010010000",
  12134=>"111111111",
  12135=>"111000000",
  12136=>"111111010",
  12137=>"010111111",
  12138=>"111000000",
  12139=>"111000000",
  12140=>"000010010",
  12141=>"111101000",
  12142=>"000111100",
  12143=>"000111010",
  12144=>"011011011",
  12145=>"000010110",
  12146=>"110011111",
  12147=>"000101000",
  12148=>"000000010",
  12149=>"001000010",
  12150=>"010110000",
  12151=>"101101001",
  12152=>"011111111",
  12153=>"111000111",
  12154=>"000000000",
  12155=>"111011000",
  12156=>"000011111",
  12157=>"111100000",
  12158=>"101111100",
  12159=>"000000011",
  12160=>"101000000",
  12161=>"111111111",
  12162=>"110000001",
  12163=>"000100101",
  12164=>"010000110",
  12165=>"001000101",
  12166=>"111111011",
  12167=>"000100100",
  12168=>"100110111",
  12169=>"110111000",
  12170=>"111111100",
  12171=>"100000111",
  12172=>"111000000",
  12173=>"111100100",
  12174=>"010101001",
  12175=>"001001010",
  12176=>"001011011",
  12177=>"011011000",
  12178=>"000111111",
  12179=>"000100000",
  12180=>"111110000",
  12181=>"000110111",
  12182=>"010000010",
  12183=>"011011111",
  12184=>"100111100",
  12185=>"110001100",
  12186=>"111000111",
  12187=>"000000000",
  12188=>"100010111",
  12189=>"111111000",
  12190=>"000000000",
  12191=>"000001000",
  12192=>"011100100",
  12193=>"111101111",
  12194=>"010000000",
  12195=>"011000000",
  12196=>"010011000",
  12197=>"100001110",
  12198=>"001001111",
  12199=>"001010011",
  12200=>"000000100",
  12201=>"011000000",
  12202=>"101001000",
  12203=>"000010110",
  12204=>"101111111",
  12205=>"000000000",
  12206=>"000000111",
  12207=>"111101001",
  12208=>"111011000",
  12209=>"111001001",
  12210=>"000000000",
  12211=>"100110011",
  12212=>"011111110",
  12213=>"111000100",
  12214=>"101000000",
  12215=>"111111000",
  12216=>"101010011",
  12217=>"011001000",
  12218=>"111010111",
  12219=>"111001100",
  12220=>"011000000",
  12221=>"111111011",
  12222=>"110111001",
  12223=>"000000000",
  12224=>"010100111",
  12225=>"000000000",
  12226=>"010010011",
  12227=>"011011110",
  12228=>"000101100",
  12229=>"010001101",
  12230=>"000111000",
  12231=>"111111000",
  12232=>"111111100",
  12233=>"000011101",
  12234=>"111000000",
  12235=>"011000001",
  12236=>"111110110",
  12237=>"000101111",
  12238=>"001110111",
  12239=>"011001110",
  12240=>"000010101",
  12241=>"111110110",
  12242=>"110000000",
  12243=>"110100100",
  12244=>"111000000",
  12245=>"001100111",
  12246=>"000010010",
  12247=>"111100000",
  12248=>"000000101",
  12249=>"000011111",
  12250=>"000100011",
  12251=>"111101000",
  12252=>"110111011",
  12253=>"000101111",
  12254=>"111101100",
  12255=>"000110001",
  12256=>"000011010",
  12257=>"101000000",
  12258=>"000111000",
  12259=>"111001001",
  12260=>"010000000",
  12261=>"111000000",
  12262=>"111010000",
  12263=>"000101110",
  12264=>"000101110",
  12265=>"111000010",
  12266=>"000000110",
  12267=>"011001001",
  12268=>"111111010",
  12269=>"001111111",
  12270=>"110000000",
  12271=>"101000000",
  12272=>"010010111",
  12273=>"011110110",
  12274=>"010000000",
  12275=>"000011110",
  12276=>"101011001",
  12277=>"111111000",
  12278=>"000000000",
  12279=>"010000000",
  12280=>"000001111",
  12281=>"001111000",
  12282=>"000010010",
  12283=>"101111010",
  12284=>"111000000",
  12285=>"111001000",
  12286=>"010110010",
  12287=>"000110000",
  12288=>"011011000",
  12289=>"001000111",
  12290=>"101000000",
  12291=>"100000111",
  12292=>"000100100",
  12293=>"110000001",
  12294=>"010111111",
  12295=>"001011010",
  12296=>"000000101",
  12297=>"000000000",
  12298=>"011111010",
  12299=>"000111010",
  12300=>"010010010",
  12301=>"100000000",
  12302=>"000011011",
  12303=>"101110000",
  12304=>"011000101",
  12305=>"001100000",
  12306=>"111101001",
  12307=>"000010010",
  12308=>"011101111",
  12309=>"101000001",
  12310=>"101101001",
  12311=>"110101110",
  12312=>"100001111",
  12313=>"101111001",
  12314=>"010100000",
  12315=>"000011111",
  12316=>"110000001",
  12317=>"001100110",
  12318=>"111010001",
  12319=>"000000000",
  12320=>"111101101",
  12321=>"111101110",
  12322=>"110010010",
  12323=>"010010010",
  12324=>"100111001",
  12325=>"110110001",
  12326=>"001000000",
  12327=>"101000111",
  12328=>"111101111",
  12329=>"001011111",
  12330=>"011011000",
  12331=>"111101111",
  12332=>"110111111",
  12333=>"111111110",
  12334=>"111001001",
  12335=>"000100110",
  12336=>"100101000",
  12337=>"111101101",
  12338=>"010000000",
  12339=>"001000101",
  12340=>"011010000",
  12341=>"001110111",
  12342=>"110000001",
  12343=>"010110101",
  12344=>"010000111",
  12345=>"000101111",
  12346=>"011001000",
  12347=>"000111011",
  12348=>"001110011",
  12349=>"111111111",
  12350=>"101001111",
  12351=>"000011111",
  12352=>"000010111",
  12353=>"101111101",
  12354=>"000100111",
  12355=>"001000010",
  12356=>"000101000",
  12357=>"111101101",
  12358=>"000111010",
  12359=>"111010000",
  12360=>"111001111",
  12361=>"011000111",
  12362=>"111000111",
  12363=>"101101100",
  12364=>"100000000",
  12365=>"011101101",
  12366=>"100101101",
  12367=>"010111111",
  12368=>"000100100",
  12369=>"111001111",
  12370=>"110001010",
  12371=>"011001100",
  12372=>"000000000",
  12373=>"001111111",
  12374=>"001101101",
  12375=>"111000001",
  12376=>"111111000",
  12377=>"000100111",
  12378=>"101111100",
  12379=>"110100100",
  12380=>"001000001",
  12381=>"010001001",
  12382=>"111110001",
  12383=>"100000101",
  12384=>"011111010",
  12385=>"111100101",
  12386=>"000111110",
  12387=>"001001101",
  12388=>"001111001",
  12389=>"000101111",
  12390=>"000101111",
  12391=>"000000101",
  12392=>"101000011",
  12393=>"011011101",
  12394=>"010011110",
  12395=>"000000000",
  12396=>"111000101",
  12397=>"000111000",
  12398=>"001010010",
  12399=>"111001000",
  12400=>"000111001",
  12401=>"000111111",
  12402=>"011001100",
  12403=>"000011000",
  12404=>"111100000",
  12405=>"000000101",
  12406=>"000000111",
  12407=>"000111000",
  12408=>"011010111",
  12409=>"111111000",
  12410=>"001001000",
  12411=>"100000000",
  12412=>"000110110",
  12413=>"110100000",
  12414=>"110000000",
  12415=>"000000000",
  12416=>"000101100",
  12417=>"001000000",
  12418=>"101000111",
  12419=>"001000000",
  12420=>"111001011",
  12421=>"000000001",
  12422=>"111111100",
  12423=>"000000100",
  12424=>"110100000",
  12425=>"001000000",
  12426=>"000100000",
  12427=>"111010000",
  12428=>"001000100",
  12429=>"111111100",
  12430=>"110111111",
  12431=>"100001101",
  12432=>"111110101",
  12433=>"101111010",
  12434=>"000001111",
  12435=>"111000100",
  12436=>"101011001",
  12437=>"000000001",
  12438=>"100111111",
  12439=>"010001011",
  12440=>"000111110",
  12441=>"010000000",
  12442=>"010011000",
  12443=>"000010000",
  12444=>"111011011",
  12445=>"001111001",
  12446=>"000000011",
  12447=>"000001000",
  12448=>"111101011",
  12449=>"101000000",
  12450=>"010000000",
  12451=>"111010010",
  12452=>"000001111",
  12453=>"110010101",
  12454=>"000000001",
  12455=>"001111110",
  12456=>"000000001",
  12457=>"100000000",
  12458=>"111101101",
  12459=>"011000000",
  12460=>"001100000",
  12461=>"101001111",
  12462=>"111100011",
  12463=>"000010111",
  12464=>"110000111",
  12465=>"010101100",
  12466=>"111001101",
  12467=>"001100111",
  12468=>"001001101",
  12469=>"011111010",
  12470=>"001001110",
  12471=>"000011100",
  12472=>"000010010",
  12473=>"000110110",
  12474=>"000010010",
  12475=>"111011000",
  12476=>"010010010",
  12477=>"111110000",
  12478=>"101000000",
  12479=>"110000100",
  12480=>"100001101",
  12481=>"000011111",
  12482=>"110000000",
  12483=>"000011100",
  12484=>"100111000",
  12485=>"101100101",
  12486=>"111110111",
  12487=>"111111111",
  12488=>"111111111",
  12489=>"000000000",
  12490=>"111011111",
  12491=>"000111000",
  12492=>"100100001",
  12493=>"000011011",
  12494=>"010001001",
  12495=>"100000011",
  12496=>"110000000",
  12497=>"001111000",
  12498=>"010000111",
  12499=>"101101101",
  12500=>"000101111",
  12501=>"010111110",
  12502=>"000001001",
  12503=>"110110000",
  12504=>"000111000",
  12505=>"000000101",
  12506=>"111001100",
  12507=>"000000000",
  12508=>"001001111",
  12509=>"110000000",
  12510=>"000001101",
  12511=>"000010101",
  12512=>"101101111",
  12513=>"111000000",
  12514=>"101000100",
  12515=>"001100000",
  12516=>"101100101",
  12517=>"000110110",
  12518=>"101011110",
  12519=>"111001000",
  12520=>"010001111",
  12521=>"100100010",
  12522=>"110011011",
  12523=>"000010000",
  12524=>"000000000",
  12525=>"001110001",
  12526=>"000110000",
  12527=>"000000000",
  12528=>"010110010",
  12529=>"101011111",
  12530=>"110010100",
  12531=>"001001001",
  12532=>"110110100",
  12533=>"111000000",
  12534=>"000000000",
  12535=>"100000000",
  12536=>"000001000",
  12537=>"110111110",
  12538=>"111111110",
  12539=>"000100111",
  12540=>"000000010",
  12541=>"000000010",
  12542=>"001111010",
  12543=>"000110110",
  12544=>"011011001",
  12545=>"000000000",
  12546=>"101000000",
  12547=>"110000000",
  12548=>"000100010",
  12549=>"110110110",
  12550=>"000010010",
  12551=>"000010000",
  12552=>"111111111",
  12553=>"000000101",
  12554=>"000000001",
  12555=>"111110010",
  12556=>"000000000",
  12557=>"111111001",
  12558=>"000101101",
  12559=>"000000010",
  12560=>"111111010",
  12561=>"000000000",
  12562=>"111111000",
  12563=>"110101000",
  12564=>"000001111",
  12565=>"111110100",
  12566=>"111011011",
  12567=>"000111111",
  12568=>"100000000",
  12569=>"001010000",
  12570=>"111111111",
  12571=>"101111111",
  12572=>"001111000",
  12573=>"111011110",
  12574=>"001001110",
  12575=>"110011001",
  12576=>"011000000",
  12577=>"000001110",
  12578=>"000000000",
  12579=>"110010111",
  12580=>"011111011",
  12581=>"010001001",
  12582=>"110110000",
  12583=>"001111111",
  12584=>"000000000",
  12585=>"110111111",
  12586=>"000010010",
  12587=>"101010000",
  12588=>"111111010",
  12589=>"110100011",
  12590=>"000001111",
  12591=>"001001000",
  12592=>"111001011",
  12593=>"001011110",
  12594=>"011010000",
  12595=>"011000000",
  12596=>"000000000",
  12597=>"000000000",
  12598=>"111101111",
  12599=>"000101001",
  12600=>"011000111",
  12601=>"010011011",
  12602=>"000000000",
  12603=>"000000010",
  12604=>"111110011",
  12605=>"010111011",
  12606=>"000000000",
  12607=>"111111111",
  12608=>"110011010",
  12609=>"101101101",
  12610=>"010111111",
  12611=>"000001111",
  12612=>"000100000",
  12613=>"000000000",
  12614=>"000010111",
  12615=>"010110000",
  12616=>"111111111",
  12617=>"001111111",
  12618=>"111010111",
  12619=>"000001000",
  12620=>"111111111",
  12621=>"010110110",
  12622=>"101000110",
  12623=>"111101010",
  12624=>"111111101",
  12625=>"111111011",
  12626=>"010001001",
  12627=>"111001001",
  12628=>"000000010",
  12629=>"011111001",
  12630=>"111111111",
  12631=>"101000111",
  12632=>"010110000",
  12633=>"001111111",
  12634=>"010110100",
  12635=>"000011011",
  12636=>"001101101",
  12637=>"001001001",
  12638=>"000000000",
  12639=>"111100011",
  12640=>"110110110",
  12641=>"111111111",
  12642=>"000000000",
  12643=>"111011011",
  12644=>"010110100",
  12645=>"101000010",
  12646=>"111111101",
  12647=>"000000000",
  12648=>"111011010",
  12649=>"000000110",
  12650=>"000111110",
  12651=>"110111111",
  12652=>"111011110",
  12653=>"000000000",
  12654=>"011111001",
  12655=>"000101101",
  12656=>"001101100",
  12657=>"001001111",
  12658=>"110111111",
  12659=>"000000110",
  12660=>"011100010",
  12661=>"000000001",
  12662=>"010000111",
  12663=>"000000000",
  12664=>"000011001",
  12665=>"111011110",
  12666=>"011000000",
  12667=>"011111110",
  12668=>"010111111",
  12669=>"110100100",
  12670=>"101101000",
  12671=>"101100111",
  12672=>"100001001",
  12673=>"111111010",
  12674=>"011111011",
  12675=>"000011010",
  12676=>"110100101",
  12677=>"000011111",
  12678=>"000001001",
  12679=>"111100010",
  12680=>"111111000",
  12681=>"001001000",
  12682=>"000000100",
  12683=>"000000001",
  12684=>"111000000",
  12685=>"010110010",
  12686=>"001001000",
  12687=>"001000000",
  12688=>"100101100",
  12689=>"110100110",
  12690=>"010110101",
  12691=>"111000000",
  12692=>"111000010",
  12693=>"100000100",
  12694=>"000001001",
  12695=>"111111111",
  12696=>"000000000",
  12697=>"000000000",
  12698=>"111111000",
  12699=>"000000000",
  12700=>"001010111",
  12701=>"010000010",
  12702=>"111000011",
  12703=>"000010011",
  12704=>"100111110",
  12705=>"001000000",
  12706=>"000010001",
  12707=>"000000010",
  12708=>"011011010",
  12709=>"110110110",
  12710=>"000000100",
  12711=>"000000000",
  12712=>"000000000",
  12713=>"101001111",
  12714=>"111111000",
  12715=>"100000000",
  12716=>"000000001",
  12717=>"110000000",
  12718=>"110100001",
  12719=>"000000110",
  12720=>"110000111",
  12721=>"011011011",
  12722=>"110101000",
  12723=>"001001100",
  12724=>"010011011",
  12725=>"000000000",
  12726=>"011000010",
  12727=>"000000100",
  12728=>"110000111",
  12729=>"111011000",
  12730=>"001010000",
  12731=>"010011001",
  12732=>"000011101",
  12733=>"111111111",
  12734=>"111111111",
  12735=>"001011101",
  12736=>"000000000",
  12737=>"001000001",
  12738=>"110010110",
  12739=>"111001110",
  12740=>"000010000",
  12741=>"111011000",
  12742=>"111011110",
  12743=>"100100100",
  12744=>"000000000",
  12745=>"111110010",
  12746=>"000100111",
  12747=>"100000011",
  12748=>"101000000",
  12749=>"110110101",
  12750=>"000000110",
  12751=>"111011000",
  12752=>"011111010",
  12753=>"110110110",
  12754=>"111011000",
  12755=>"111111011",
  12756=>"000000000",
  12757=>"100000000",
  12758=>"110111101",
  12759=>"110010110",
  12760=>"010010010",
  12761=>"110100000",
  12762=>"011111010",
  12763=>"000000000",
  12764=>"111001000",
  12765=>"010011000",
  12766=>"001101001",
  12767=>"111111111",
  12768=>"000010000",
  12769=>"000000001",
  12770=>"000000000",
  12771=>"111101011",
  12772=>"000000000",
  12773=>"110111111",
  12774=>"011011000",
  12775=>"011000000",
  12776=>"000000111",
  12777=>"000000000",
  12778=>"000000000",
  12779=>"000000000",
  12780=>"101010110",
  12781=>"000100010",
  12782=>"111010000",
  12783=>"111000010",
  12784=>"110011000",
  12785=>"110100000",
  12786=>"111111111",
  12787=>"110111111",
  12788=>"011100100",
  12789=>"101101100",
  12790=>"000000000",
  12791=>"101111011",
  12792=>"101111111",
  12793=>"110110010",
  12794=>"111111111",
  12795=>"010111100",
  12796=>"000110111",
  12797=>"000000000",
  12798=>"110111111",
  12799=>"000100111",
  12800=>"001001111",
  12801=>"111011110",
  12802=>"001000001",
  12803=>"111111011",
  12804=>"000110001",
  12805=>"100110110",
  12806=>"000110000",
  12807=>"110000111",
  12808=>"010111101",
  12809=>"100100101",
  12810=>"011010000",
  12811=>"111001101",
  12812=>"100000010",
  12813=>"111111011",
  12814=>"001011111",
  12815=>"111110010",
  12816=>"111100111",
  12817=>"100110100",
  12818=>"011010110",
  12819=>"100010000",
  12820=>"100100011",
  12821=>"111111110",
  12822=>"011011010",
  12823=>"000011000",
  12824=>"000010111",
  12825=>"001110011",
  12826=>"001010000",
  12827=>"001011111",
  12828=>"000000000",
  12829=>"100001001",
  12830=>"001001001",
  12831=>"011011011",
  12832=>"011100001",
  12833=>"111101011",
  12834=>"100100100",
  12835=>"000110110",
  12836=>"101011011",
  12837=>"000000001",
  12838=>"001001011",
  12839=>"011100010",
  12840=>"000101111",
  12841=>"000001111",
  12842=>"011000000",
  12843=>"100110110",
  12844=>"001001101",
  12845=>"001011100",
  12846=>"100011011",
  12847=>"000100000",
  12848=>"010110100",
  12849=>"011111000",
  12850=>"001100100",
  12851=>"111100100",
  12852=>"011001111",
  12853=>"011111101",
  12854=>"100111111",
  12855=>"001011000",
  12856=>"111101111",
  12857=>"011001011",
  12858=>"111000010",
  12859=>"010110110",
  12860=>"001101001",
  12861=>"011011010",
  12862=>"000000000",
  12863=>"101001000",
  12864=>"011100000",
  12865=>"000000011",
  12866=>"010010000",
  12867=>"011001001",
  12868=>"110010110",
  12869=>"010000111",
  12870=>"001000000",
  12871=>"111101011",
  12872=>"111001011",
  12873=>"110100101",
  12874=>"011001011",
  12875=>"001011001",
  12876=>"111000111",
  12877=>"001000000",
  12878=>"001001011",
  12879=>"011100111",
  12880=>"011011011",
  12881=>"000001101",
  12882=>"010000000",
  12883=>"010011111",
  12884=>"100000000",
  12885=>"011110001",
  12886=>"001001101",
  12887=>"100100100",
  12888=>"010011010",
  12889=>"011011010",
  12890=>"000001000",
  12891=>"111111111",
  12892=>"000110100",
  12893=>"110000100",
  12894=>"100111110",
  12895=>"011101111",
  12896=>"010010000",
  12897=>"011100001",
  12898=>"000000001",
  12899=>"011111001",
  12900=>"101101111",
  12901=>"001011000",
  12902=>"000100101",
  12903=>"011001111",
  12904=>"111101011",
  12905=>"110110100",
  12906=>"111011001",
  12907=>"001011000",
  12908=>"000001111",
  12909=>"110110110",
  12910=>"111110000",
  12911=>"010000000",
  12912=>"000000010",
  12913=>"111111100",
  12914=>"010010100",
  12915=>"111110111",
  12916=>"100101001",
  12917=>"011001001",
  12918=>"011001000",
  12919=>"110110000",
  12920=>"100000100",
  12921=>"100000110",
  12922=>"000110100",
  12923=>"110110100",
  12924=>"000000100",
  12925=>"100000111",
  12926=>"100111001",
  12927=>"001001001",
  12928=>"011001000",
  12929=>"111001001",
  12930=>"110100100",
  12931=>"110111101",
  12932=>"001111100",
  12933=>"011000011",
  12934=>"011011001",
  12935=>"001110111",
  12936=>"111111111",
  12937=>"010101001",
  12938=>"110000000",
  12939=>"110100110",
  12940=>"100100100",
  12941=>"100100010",
  12942=>"001011100",
  12943=>"000000000",
  12944=>"011001010",
  12945=>"001011111",
  12946=>"001110010",
  12947=>"001011111",
  12948=>"001101101",
  12949=>"100100110",
  12950=>"011011001",
  12951=>"001000001",
  12952=>"000000000",
  12953=>"111000000",
  12954=>"000001000",
  12955=>"110110110",
  12956=>"000010000",
  12957=>"001001101",
  12958=>"011000001",
  12959=>"001001001",
  12960=>"111011111",
  12961=>"010111010",
  12962=>"100010110",
  12963=>"011001111",
  12964=>"111111010",
  12965=>"000000000",
  12966=>"110100000",
  12967=>"100100100",
  12968=>"010100110",
  12969=>"011111110",
  12970=>"100100111",
  12971=>"000000111",
  12972=>"000110000",
  12973=>"001001001",
  12974=>"001011000",
  12975=>"110100111",
  12976=>"101000000",
  12977=>"100100100",
  12978=>"010111100",
  12979=>"011000000",
  12980=>"111111111",
  12981=>"111011000",
  12982=>"111111111",
  12983=>"100110011",
  12984=>"010110000",
  12985=>"000000011",
  12986=>"000011101",
  12987=>"001100000",
  12988=>"100101111",
  12989=>"100110110",
  12990=>"111010111",
  12991=>"100100100",
  12992=>"001011101",
  12993=>"000001000",
  12994=>"001011011",
  12995=>"111011000",
  12996=>"110110100",
  12997=>"000001001",
  12998=>"100100110",
  12999=>"111000011",
  13000=>"100100111",
  13001=>"011011011",
  13002=>"100100000",
  13003=>"011001000",
  13004=>"011001000",
  13005=>"001011110",
  13006=>"011001000",
  13007=>"000100100",
  13008=>"000001000",
  13009=>"111011110",
  13010=>"011100101",
  13011=>"001111001",
  13012=>"001001011",
  13013=>"100110111",
  13014=>"001001111",
  13015=>"000001011",
  13016=>"111011000",
  13017=>"100100110",
  13018=>"000100000",
  13019=>"100100100",
  13020=>"011011111",
  13021=>"110111110",
  13022=>"001000000",
  13023=>"000011111",
  13024=>"001111001",
  13025=>"101100001",
  13026=>"100100000",
  13027=>"001001101",
  13028=>"000000000",
  13029=>"110111110",
  13030=>"001001001",
  13031=>"111011011",
  13032=>"100110011",
  13033=>"110000100",
  13034=>"000110111",
  13035=>"110111111",
  13036=>"110110100",
  13037=>"101110000",
  13038=>"000100100",
  13039=>"100001000",
  13040=>"011011000",
  13041=>"011111111",
  13042=>"011011001",
  13043=>"000000100",
  13044=>"000000000",
  13045=>"100000110",
  13046=>"000000010",
  13047=>"100100000",
  13048=>"111110110",
  13049=>"110100000",
  13050=>"111111011",
  13051=>"000000110",
  13052=>"111001011",
  13053=>"100110000",
  13054=>"111001011",
  13055=>"001001001",
  13056=>"110010000",
  13057=>"000110000",
  13058=>"001001111",
  13059=>"000000000",
  13060=>"100110110",
  13061=>"101001100",
  13062=>"110110000",
  13063=>"000110110",
  13064=>"010011110",
  13065=>"000111000",
  13066=>"010010011",
  13067=>"000001001",
  13068=>"110110110",
  13069=>"110000000",
  13070=>"110110000",
  13071=>"100110000",
  13072=>"011000100",
  13073=>"001000001",
  13074=>"001001000",
  13075=>"111111111",
  13076=>"111111111",
  13077=>"001001000",
  13078=>"010101011",
  13079=>"111111000",
  13080=>"000000001",
  13081=>"111111111",
  13082=>"010000000",
  13083=>"000000011",
  13084=>"101001001",
  13085=>"010111111",
  13086=>"110100000",
  13087=>"000110110",
  13088=>"111001101",
  13089=>"011001111",
  13090=>"000110110",
  13091=>"110111110",
  13092=>"100000000",
  13093=>"100100000",
  13094=>"000000110",
  13095=>"100110100",
  13096=>"011001000",
  13097=>"110111011",
  13098=>"110000000",
  13099=>"001000011",
  13100=>"000000000",
  13101=>"001111111",
  13102=>"111110000",
  13103=>"110111111",
  13104=>"000001000",
  13105=>"011011000",
  13106=>"111011111",
  13107=>"111001000",
  13108=>"000010000",
  13109=>"010011111",
  13110=>"110100000",
  13111=>"000011100",
  13112=>"111110100",
  13113=>"011011110",
  13114=>"000101111",
  13115=>"001111111",
  13116=>"100000110",
  13117=>"111111000",
  13118=>"000000001",
  13119=>"010111000",
  13120=>"110111111",
  13121=>"111110000",
  13122=>"111000100",
  13123=>"100100011",
  13124=>"000001110",
  13125=>"000110010",
  13126=>"001000000",
  13127=>"111001001",
  13128=>"000110110",
  13129=>"110110000",
  13130=>"110000111",
  13131=>"111110010",
  13132=>"001001000",
  13133=>"011001000",
  13134=>"100100101",
  13135=>"001010111",
  13136=>"110000001",
  13137=>"110000000",
  13138=>"110000000",
  13139=>"011011001",
  13140=>"110110000",
  13141=>"101110010",
  13142=>"001111010",
  13143=>"111110000",
  13144=>"110111110",
  13145=>"001011011",
  13146=>"000111100",
  13147=>"011111111",
  13148=>"001000001",
  13149=>"001001000",
  13150=>"111001011",
  13151=>"000111001",
  13152=>"110110100",
  13153=>"010100101",
  13154=>"001000111",
  13155=>"011010000",
  13156=>"000000000",
  13157=>"100001111",
  13158=>"000110110",
  13159=>"111011000",
  13160=>"000110000",
  13161=>"111000000",
  13162=>"001111111",
  13163=>"101000100",
  13164=>"011000100",
  13165=>"001010111",
  13166=>"001001111",
  13167=>"000111110",
  13168=>"110111001",
  13169=>"000010110",
  13170=>"011001000",
  13171=>"110110010",
  13172=>"011000111",
  13173=>"000000110",
  13174=>"000110110",
  13175=>"110110110",
  13176=>"001000011",
  13177=>"010010010",
  13178=>"111001001",
  13179=>"011001001",
  13180=>"000100100",
  13181=>"101000100",
  13182=>"000000001",
  13183=>"110110000",
  13184=>"110111100",
  13185=>"000111110",
  13186=>"110000110",
  13187=>"000101101",
  13188=>"111110001",
  13189=>"000001000",
  13190=>"111011011",
  13191=>"000101110",
  13192=>"110001101",
  13193=>"100100010",
  13194=>"011001111",
  13195=>"101011100",
  13196=>"001001111",
  13197=>"000000001",
  13198=>"000000111",
  13199=>"000000001",
  13200=>"101000100",
  13201=>"110110000",
  13202=>"000100101",
  13203=>"110101010",
  13204=>"000111111",
  13205=>"111001111",
  13206=>"110101101",
  13207=>"000010011",
  13208=>"111111100",
  13209=>"001010110",
  13210=>"110110000",
  13211=>"001110010",
  13212=>"000100001",
  13213=>"111001111",
  13214=>"001001000",
  13215=>"101000000",
  13216=>"110100000",
  13217=>"000000111",
  13218=>"100100100",
  13219=>"111100000",
  13220=>"000001001",
  13221=>"101100110",
  13222=>"000110100",
  13223=>"000000100",
  13224=>"101011011",
  13225=>"001100100",
  13226=>"001000000",
  13227=>"110000001",
  13228=>"000110111",
  13229=>"011000011",
  13230=>"000001011",
  13231=>"110000000",
  13232=>"000100110",
  13233=>"000000100",
  13234=>"011010000",
  13235=>"001100000",
  13236=>"001011011",
  13237=>"001111110",
  13238=>"000111111",
  13239=>"000110010",
  13240=>"010001111",
  13241=>"000100110",
  13242=>"010011111",
  13243=>"110000001",
  13244=>"000010110",
  13245=>"011001001",
  13246=>"100000011",
  13247=>"000001000",
  13248=>"000110011",
  13249=>"001000111",
  13250=>"111101001",
  13251=>"100110110",
  13252=>"001000000",
  13253=>"001001111",
  13254=>"110101000",
  13255=>"110110000",
  13256=>"000010000",
  13257=>"000110010",
  13258=>"000000101",
  13259=>"001001111",
  13260=>"100111000",
  13261=>"001111000",
  13262=>"000000000",
  13263=>"011001111",
  13264=>"001011011",
  13265=>"010110100",
  13266=>"011110000",
  13267=>"000000010",
  13268=>"100100000",
  13269=>"111000000",
  13270=>"111001111",
  13271=>"100000100",
  13272=>"000000110",
  13273=>"111111111",
  13274=>"011110111",
  13275=>"001011001",
  13276=>"000001100",
  13277=>"110111010",
  13278=>"110111010",
  13279=>"110110100",
  13280=>"001000111",
  13281=>"000000111",
  13282=>"000111110",
  13283=>"011111100",
  13284=>"001000000",
  13285=>"001000000",
  13286=>"111001000",
  13287=>"010011000",
  13288=>"111111111",
  13289=>"001000000",
  13290=>"000010010",
  13291=>"001100110",
  13292=>"011110110",
  13293=>"000000010",
  13294=>"000000001",
  13295=>"000000000",
  13296=>"110111110",
  13297=>"001000111",
  13298=>"110110010",
  13299=>"100000110",
  13300=>"000101000",
  13301=>"011111111",
  13302=>"110010000",
  13303=>"000110000",
  13304=>"110111110",
  13305=>"111110000",
  13306=>"111010111",
  13307=>"000110111",
  13308=>"001000100",
  13309=>"001001000",
  13310=>"001001101",
  13311=>"000000101",
  13312=>"110110010",
  13313=>"000001110",
  13314=>"101101101",
  13315=>"010010100",
  13316=>"111110111",
  13317=>"011011101",
  13318=>"010000111",
  13319=>"110011101",
  13320=>"101001000",
  13321=>"101101000",
  13322=>"000001001",
  13323=>"000100100",
  13324=>"110101100",
  13325=>"110000011",
  13326=>"110100110",
  13327=>"010111011",
  13328=>"101001001",
  13329=>"001111111",
  13330=>"110010000",
  13331=>"111010110",
  13332=>"011000000",
  13333=>"101101101",
  13334=>"100110001",
  13335=>"101101111",
  13336=>"100100000",
  13337=>"001001001",
  13338=>"100011000",
  13339=>"110110010",
  13340=>"000000010",
  13341=>"001000111",
  13342=>"001000000",
  13343=>"010010010",
  13344=>"101001000",
  13345=>"001000111",
  13346=>"111100110",
  13347=>"111101110",
  13348=>"010010010",
  13349=>"000000000",
  13350=>"101100100",
  13351=>"001101111",
  13352=>"111011011",
  13353=>"111011111",
  13354=>"111110101",
  13355=>"000001001",
  13356=>"110110110",
  13357=>"000000000",
  13358=>"010100000",
  13359=>"111011001",
  13360=>"000000000",
  13361=>"011010011",
  13362=>"111001111",
  13363=>"101111101",
  13364=>"101111010",
  13365=>"100010010",
  13366=>"001000010",
  13367=>"101100100",
  13368=>"000111000",
  13369=>"111000100",
  13370=>"010010111",
  13371=>"101111111",
  13372=>"111010111",
  13373=>"010010111",
  13374=>"100101001",
  13375=>"010000000",
  13376=>"000001001",
  13377=>"000010000",
  13378=>"010000111",
  13379=>"000100011",
  13380=>"010000111",
  13381=>"001001000",
  13382=>"001001010",
  13383=>"110110111",
  13384=>"110010000",
  13385=>"101001010",
  13386=>"101000101",
  13387=>"111111110",
  13388=>"001101111",
  13389=>"111010111",
  13390=>"111111101",
  13391=>"010001101",
  13392=>"000000001",
  13393=>"111000110",
  13394=>"011000000",
  13395=>"011010011",
  13396=>"000111000",
  13397=>"000001011",
  13398=>"110010010",
  13399=>"101101101",
  13400=>"001011000",
  13401=>"011010110",
  13402=>"011010010",
  13403=>"110110111",
  13404=>"101100000",
  13405=>"111010011",
  13406=>"111101111",
  13407=>"101100000",
  13408=>"100100000",
  13409=>"010010000",
  13410=>"001101001",
  13411=>"110110010",
  13412=>"111111111",
  13413=>"010010000",
  13414=>"111001111",
  13415=>"000000000",
  13416=>"000000011",
  13417=>"000001101",
  13418=>"011100000",
  13419=>"000001101",
  13420=>"000000000",
  13421=>"011111111",
  13422=>"001000000",
  13423=>"110010111",
  13424=>"110110010",
  13425=>"010000001",
  13426=>"100000011",
  13427=>"111111001",
  13428=>"000001010",
  13429=>"010010110",
  13430=>"111000110",
  13431=>"101000010",
  13432=>"001000001",
  13433=>"110010011",
  13434=>"111111000",
  13435=>"100000000",
  13436=>"110010000",
  13437=>"011010110",
  13438=>"100000111",
  13439=>"000000010",
  13440=>"101101000",
  13441=>"010000101",
  13442=>"101000000",
  13443=>"010110001",
  13444=>"011000100",
  13445=>"000100111",
  13446=>"000000000",
  13447=>"100100000",
  13448=>"010010010",
  13449=>"101100101",
  13450=>"010010111",
  13451=>"000001101",
  13452=>"111000000",
  13453=>"100001111",
  13454=>"111111111",
  13455=>"100100010",
  13456=>"011010011",
  13457=>"111110001",
  13458=>"111000000",
  13459=>"101000000",
  13460=>"111001100",
  13461=>"101101101",
  13462=>"111111011",
  13463=>"110110110",
  13464=>"111000111",
  13465=>"000001101",
  13466=>"101000110",
  13467=>"101001101",
  13468=>"000110010",
  13469=>"101100101",
  13470=>"000101110",
  13471=>"000001000",
  13472=>"001100010",
  13473=>"000101001",
  13474=>"011000001",
  13475=>"110111000",
  13476=>"010110001",
  13477=>"111011111",
  13478=>"010110010",
  13479=>"110011111",
  13480=>"101101101",
  13481=>"000001001",
  13482=>"110110110",
  13483=>"100101111",
  13484=>"010000000",
  13485=>"110010010",
  13486=>"011010110",
  13487=>"111101111",
  13488=>"100100000",
  13489=>"110110010",
  13490=>"111011111",
  13491=>"000001001",
  13492=>"011010110",
  13493=>"010010111",
  13494=>"111101000",
  13495=>"010010101",
  13496=>"110000111",
  13497=>"100000000",
  13498=>"010010011",
  13499=>"001000000",
  13500=>"111000011",
  13501=>"100101100",
  13502=>"110000100",
  13503=>"001001001",
  13504=>"101001000",
  13505=>"100101000",
  13506=>"000111110",
  13507=>"011110010",
  13508=>"010000001",
  13509=>"000011011",
  13510=>"010000111",
  13511=>"001001001",
  13512=>"000000000",
  13513=>"111111111",
  13514=>"000010000",
  13515=>"101100101",
  13516=>"111101111",
  13517=>"111000000",
  13518=>"000000000",
  13519=>"111101001",
  13520=>"101001111",
  13521=>"110010110",
  13522=>"100101000",
  13523=>"010110111",
  13524=>"101100110",
  13525=>"001000010",
  13526=>"000010111",
  13527=>"000010110",
  13528=>"111101101",
  13529=>"000101110",
  13530=>"101001101",
  13531=>"001101101",
  13532=>"010000100",
  13533=>"000111001",
  13534=>"111111000",
  13535=>"111000100",
  13536=>"100100101",
  13537=>"100110101",
  13538=>"111111101",
  13539=>"011010011",
  13540=>"101101101",
  13541=>"011010110",
  13542=>"111111010",
  13543=>"100110110",
  13544=>"101111101",
  13545=>"100000011",
  13546=>"100100100",
  13547=>"101111110",
  13548=>"100000100",
  13549=>"101001100",
  13550=>"111000000",
  13551=>"000000111",
  13552=>"000001010",
  13553=>"001001010",
  13554=>"010000000",
  13555=>"110010010",
  13556=>"011011010",
  13557=>"000010100",
  13558=>"101100001",
  13559=>"100110110",
  13560=>"101001101",
  13561=>"000000101",
  13562=>"111101100",
  13563=>"111111110",
  13564=>"111110111",
  13565=>"000111011",
  13566=>"110110111",
  13567=>"101001000",
  13568=>"001000000",
  13569=>"011001011",
  13570=>"100100100",
  13571=>"011010001",
  13572=>"110000101",
  13573=>"011110110",
  13574=>"101111001",
  13575=>"011011000",
  13576=>"011000111",
  13577=>"100100100",
  13578=>"000011101",
  13579=>"000011000",
  13580=>"011011011",
  13581=>"001001011",
  13582=>"100110101",
  13583=>"110010100",
  13584=>"101000111",
  13585=>"110100110",
  13586=>"110110001",
  13587=>"111100110",
  13588=>"110100111",
  13589=>"111100110",
  13590=>"100111011",
  13591=>"111111110",
  13592=>"100100110",
  13593=>"111010000",
  13594=>"001001011",
  13595=>"001001001",
  13596=>"100110011",
  13597=>"010000000",
  13598=>"000100001",
  13599=>"011001011",
  13600=>"100110110",
  13601=>"010001111",
  13602=>"100001001",
  13603=>"011011011",
  13604=>"000000100",
  13605=>"001011111",
  13606=>"100100110",
  13607=>"100000000",
  13608=>"110110111",
  13609=>"001001111",
  13610=>"100110110",
  13611=>"001011011",
  13612=>"000000000",
  13613=>"011100110",
  13614=>"001111111",
  13615=>"100110010",
  13616=>"101100110",
  13617=>"100100000",
  13618=>"110100110",
  13619=>"100110100",
  13620=>"001000000",
  13621=>"101011010",
  13622=>"001011011",
  13623=>"011000011",
  13624=>"001100100",
  13625=>"001000011",
  13626=>"000000000",
  13627=>"111100010",
  13628=>"011011001",
  13629=>"001011110",
  13630=>"100100000",
  13631=>"001000011",
  13632=>"100110100",
  13633=>"000100110",
  13634=>"101111010",
  13635=>"001010010",
  13636=>"010101111",
  13637=>"001001011",
  13638=>"000010000",
  13639=>"001111010",
  13640=>"011111101",
  13641=>"001000001",
  13642=>"011010001",
  13643=>"111011011",
  13644=>"000100110",
  13645=>"110110101",
  13646=>"110110110",
  13647=>"100110110",
  13648=>"001000001",
  13649=>"001100000",
  13650=>"100101111",
  13651=>"001100000",
  13652=>"001111111",
  13653=>"011001011",
  13654=>"000001101",
  13655=>"100000000",
  13656=>"001011011",
  13657=>"000110111",
  13658=>"000000000",
  13659=>"101110110",
  13660=>"000010111",
  13661=>"001001001",
  13662=>"110100110",
  13663=>"010000010",
  13664=>"000001001",
  13665=>"010001001",
  13666=>"110110001",
  13667=>"100011011",
  13668=>"010000001",
  13669=>"001001000",
  13670=>"011001001",
  13671=>"100100101",
  13672=>"100001000",
  13673=>"101110110",
  13674=>"100110000",
  13675=>"011000001",
  13676=>"001001000",
  13677=>"110111101",
  13678=>"000001000",
  13679=>"011011001",
  13680=>"101010000",
  13681=>"000001000",
  13682=>"001001000",
  13683=>"000000001",
  13684=>"001011000",
  13685=>"001110111",
  13686=>"100001000",
  13687=>"000000011",
  13688=>"101101110",
  13689=>"001001001",
  13690=>"010110100",
  13691=>"110110010",
  13692=>"011010000",
  13693=>"011010001",
  13694=>"110110110",
  13695=>"000010001",
  13696=>"110100100",
  13697=>"011001101",
  13698=>"001111111",
  13699=>"011110011",
  13700=>"101000001",
  13701=>"001111000",
  13702=>"001101001",
  13703=>"000011011",
  13704=>"010011111",
  13705=>"001111001",
  13706=>"111011001",
  13707=>"001100100",
  13708=>"000010000",
  13709=>"110110010",
  13710=>"110110110",
  13711=>"110000000",
  13712=>"011011001",
  13713=>"100000110",
  13714=>"000010100",
  13715=>"001010011",
  13716=>"000000001",
  13717=>"100100000",
  13718=>"001001011",
  13719=>"001100111",
  13720=>"001001011",
  13721=>"110000010",
  13722=>"100110100",
  13723=>"100110001",
  13724=>"001010011",
  13725=>"000110001",
  13726=>"001110110",
  13727=>"011010000",
  13728=>"100001000",
  13729=>"110111111",
  13730=>"001001111",
  13731=>"100110000",
  13732=>"001110011",
  13733=>"011000100",
  13734=>"010010010",
  13735=>"001001111",
  13736=>"000100110",
  13737=>"010100001",
  13738=>"110110111",
  13739=>"100000000",
  13740=>"010100011",
  13741=>"001010110",
  13742=>"011010111",
  13743=>"000101011",
  13744=>"110101001",
  13745=>"011001001",
  13746=>"110110011",
  13747=>"110001001",
  13748=>"001000011",
  13749=>"001011011",
  13750=>"000000001",
  13751=>"010111010",
  13752=>"001000001",
  13753=>"010000000",
  13754=>"001001011",
  13755=>"001011011",
  13756=>"000001101",
  13757=>"110111011",
  13758=>"100110101",
  13759=>"100100100",
  13760=>"110110100",
  13761=>"000110101",
  13762=>"001111011",
  13763=>"100110101",
  13764=>"000100100",
  13765=>"100101110",
  13766=>"011001000",
  13767=>"001001010",
  13768=>"011000111",
  13769=>"001001001",
  13770=>"001010110",
  13771=>"000000111",
  13772=>"001110100",
  13773=>"000011000",
  13774=>"100000101",
  13775=>"100000000",
  13776=>"100100000",
  13777=>"111011111",
  13778=>"001000001",
  13779=>"001001110",
  13780=>"110110100",
  13781=>"011011011",
  13782=>"001001011",
  13783=>"000110000",
  13784=>"011001110",
  13785=>"001001101",
  13786=>"110001100",
  13787=>"100110100",
  13788=>"011011000",
  13789=>"011001001",
  13790=>"000000010",
  13791=>"110100010",
  13792=>"100100101",
  13793=>"110110100",
  13794=>"110100111",
  13795=>"010001001",
  13796=>"111000100",
  13797=>"011011011",
  13798=>"000000011",
  13799=>"011010001",
  13800=>"000000000",
  13801=>"011000100",
  13802=>"000000100",
  13803=>"010101111",
  13804=>"001001011",
  13805=>"100001000",
  13806=>"000100001",
  13807=>"110010011",
  13808=>"011001010",
  13809=>"111111011",
  13810=>"001101110",
  13811=>"011001001",
  13812=>"011010100",
  13813=>"100100101",
  13814=>"100100100",
  13815=>"100110110",
  13816=>"110100000",
  13817=>"110110111",
  13818=>"011011011",
  13819=>"011011011",
  13820=>"110100111",
  13821=>"000110100",
  13822=>"100010111",
  13823=>"110110000",
  13824=>"011011001",
  13825=>"101101100",
  13826=>"101000101",
  13827=>"000000001",
  13828=>"011000000",
  13829=>"000100111",
  13830=>"000000000",
  13831=>"000100111",
  13832=>"111100001",
  13833=>"001010000",
  13834=>"001000111",
  13835=>"000000100",
  13836=>"011000100",
  13837=>"000111111",
  13838=>"001011001",
  13839=>"111011001",
  13840=>"011101101",
  13841=>"100001000",
  13842=>"001000000",
  13843=>"000000110",
  13844=>"111111101",
  13845=>"000000111",
  13846=>"111001101",
  13847=>"010110011",
  13848=>"000111110",
  13849=>"000001110",
  13850=>"111111100",
  13851=>"111000000",
  13852=>"000000110",
  13853=>"001111111",
  13854=>"110100000",
  13855=>"000111111",
  13856=>"111100100",
  13857=>"111011000",
  13858=>"010010000",
  13859=>"110111111",
  13860=>"001011111",
  13861=>"110000000",
  13862=>"111010000",
  13863=>"111000000",
  13864=>"100100110",
  13865=>"010100100",
  13866=>"000111101",
  13867=>"001001001",
  13868=>"111011001",
  13869=>"000001100",
  13870=>"111011111",
  13871=>"100000010",
  13872=>"110111100",
  13873=>"001100111",
  13874=>"111111111",
  13875=>"011001000",
  13876=>"000000000",
  13877=>"010001000",
  13878=>"111111111",
  13879=>"010111111",
  13880=>"111111000",
  13881=>"000000110",
  13882=>"000110111",
  13883=>"011001000",
  13884=>"110111101",
  13885=>"010111010",
  13886=>"110111101",
  13887=>"000010000",
  13888=>"100001111",
  13889=>"111101101",
  13890=>"100101010",
  13891=>"000000000",
  13892=>"111011000",
  13893=>"111110100",
  13894=>"101000110",
  13895=>"111000000",
  13896=>"101011101",
  13897=>"111111100",
  13898=>"111001101",
  13899=>"000011110",
  13900=>"111111000",
  13901=>"100001100",
  13902=>"100000001",
  13903=>"000000111",
  13904=>"001000010",
  13905=>"000111110",
  13906=>"101010101",
  13907=>"001001001",
  13908=>"000000110",
  13909=>"110110100",
  13910=>"100110110",
  13911=>"110010000",
  13912=>"000101111",
  13913=>"000111011",
  13914=>"110010001",
  13915=>"100110110",
  13916=>"110010000",
  13917=>"001001011",
  13918=>"110110011",
  13919=>"100000000",
  13920=>"111110000",
  13921=>"101110110",
  13922=>"111110000",
  13923=>"110100100",
  13924=>"110111110",
  13925=>"000011100",
  13926=>"010010001",
  13927=>"011000000",
  13928=>"110000101",
  13929=>"011000100",
  13930=>"000000011",
  13931=>"000110111",
  13932=>"111111101",
  13933=>"000100101",
  13934=>"011101011",
  13935=>"000000010",
  13936=>"111111001",
  13937=>"111111100",
  13938=>"011111011",
  13939=>"001111100",
  13940=>"010000000",
  13941=>"111000100",
  13942=>"000000010",
  13943=>"111010001",
  13944=>"111100000",
  13945=>"010100010",
  13946=>"111011100",
  13947=>"000100000",
  13948=>"100110111",
  13949=>"100100100",
  13950=>"111101101",
  13951=>"000111100",
  13952=>"111100100",
  13953=>"100011110",
  13954=>"111110000",
  13955=>"010000001",
  13956=>"010000100",
  13957=>"000010101",
  13958=>"110101100",
  13959=>"001001000",
  13960=>"111111010",
  13961=>"000000111",
  13962=>"110110111",
  13963=>"010010111",
  13964=>"110000000",
  13965=>"000101100",
  13966=>"101111101",
  13967=>"010000000",
  13968=>"101000010",
  13969=>"000000101",
  13970=>"110111101",
  13971=>"001000001",
  13972=>"000111111",
  13973=>"000000101",
  13974=>"000111000",
  13975=>"011011001",
  13976=>"101111111",
  13977=>"000000111",
  13978=>"000100111",
  13979=>"101101111",
  13980=>"111111101",
  13981=>"111000111",
  13982=>"001101111",
  13983=>"000010000",
  13984=>"101010111",
  13985=>"001000000",
  13986=>"011001111",
  13987=>"000111000",
  13988=>"100000111",
  13989=>"110111100",
  13990=>"110110000",
  13991=>"001101111",
  13992=>"100011111",
  13993=>"111111000",
  13994=>"000000100",
  13995=>"000000010",
  13996=>"110010100",
  13997=>"111000100",
  13998=>"011001010",
  13999=>"000000000",
  14000=>"110001101",
  14001=>"101000001",
  14002=>"111011011",
  14003=>"000100100",
  14004=>"111111000",
  14005=>"111111000",
  14006=>"111111111",
  14007=>"111001000",
  14008=>"011111011",
  14009=>"000110110",
  14010=>"000101010",
  14011=>"011111000",
  14012=>"000100111",
  14013=>"111111110",
  14014=>"101100010",
  14015=>"000000000",
  14016=>"011011001",
  14017=>"010010000",
  14018=>"101111010",
  14019=>"100100110",
  14020=>"000000000",
  14021=>"100110001",
  14022=>"111111111",
  14023=>"000000000",
  14024=>"101101111",
  14025=>"111000000",
  14026=>"111111111",
  14027=>"000001111",
  14028=>"000000111",
  14029=>"001111110",
  14030=>"011011010",
  14031=>"000001111",
  14032=>"000000000",
  14033=>"100111111",
  14034=>"000000100",
  14035=>"000101101",
  14036=>"011010001",
  14037=>"110111111",
  14038=>"101111000",
  14039=>"000001011",
  14040=>"000010111",
  14041=>"010110000",
  14042=>"000110101",
  14043=>"010010000",
  14044=>"111001001",
  14045=>"011000110",
  14046=>"011010000",
  14047=>"001000000",
  14048=>"000101111",
  14049=>"101100100",
  14050=>"100000111",
  14051=>"110100101",
  14052=>"000010000",
  14053=>"111010000",
  14054=>"000010111",
  14055=>"101110110",
  14056=>"010101111",
  14057=>"111010100",
  14058=>"100001111",
  14059=>"111101000",
  14060=>"000000000",
  14061=>"111000111",
  14062=>"010010000",
  14063=>"101101110",
  14064=>"000111111",
  14065=>"011111111",
  14066=>"111000000",
  14067=>"100100100",
  14068=>"110110000",
  14069=>"010000111",
  14070=>"001000000",
  14071=>"000100001",
  14072=>"000111111",
  14073=>"000001010",
  14074=>"010000011",
  14075=>"100101110",
  14076=>"000111111",
  14077=>"011011000",
  14078=>"111111110",
  14079=>"000001011",
  14080=>"001111111",
  14081=>"100111010",
  14082=>"000100100",
  14083=>"111101000",
  14084=>"001101011",
  14085=>"000001111",
  14086=>"101101011",
  14087=>"101111110",
  14088=>"111010000",
  14089=>"011010000",
  14090=>"001000000",
  14091=>"000000000",
  14092=>"101100100",
  14093=>"011110000",
  14094=>"011001000",
  14095=>"000111111",
  14096=>"010000000",
  14097=>"010000000",
  14098=>"000100011",
  14099=>"100000000",
  14100=>"100011010",
  14101=>"011000110",
  14102=>"100100001",
  14103=>"001111111",
  14104=>"101100000",
  14105=>"110001111",
  14106=>"000011000",
  14107=>"000100010",
  14108=>"000000010",
  14109=>"000000101",
  14110=>"011011111",
  14111=>"111111001",
  14112=>"110100110",
  14113=>"011111011",
  14114=>"100000000",
  14115=>"110010000",
  14116=>"001011001",
  14117=>"101011111",
  14118=>"011010110",
  14119=>"101001010",
  14120=>"000111111",
  14121=>"010111000",
  14122=>"000000000",
  14123=>"100100111",
  14124=>"001001111",
  14125=>"101111001",
  14126=>"000101111",
  14127=>"100101101",
  14128=>"101011010",
  14129=>"000001000",
  14130=>"010010000",
  14131=>"011001101",
  14132=>"000000000",
  14133=>"010011111",
  14134=>"110011010",
  14135=>"111101000",
  14136=>"110111111",
  14137=>"000000000",
  14138=>"111100000",
  14139=>"001000000",
  14140=>"010011110",
  14141=>"111111111",
  14142=>"010000000",
  14143=>"111011000",
  14144=>"101000100",
  14145=>"000100101",
  14146=>"111111000",
  14147=>"011000000",
  14148=>"100111111",
  14149=>"000000011",
  14150=>"010010000",
  14151=>"111101101",
  14152=>"000001001",
  14153=>"011010000",
  14154=>"000000000",
  14155=>"100010111",
  14156=>"010000000",
  14157=>"101101000",
  14158=>"000110110",
  14159=>"000011000",
  14160=>"001000000",
  14161=>"101110001",
  14162=>"110111111",
  14163=>"000100001",
  14164=>"000000000",
  14165=>"100100011",
  14166=>"101100100",
  14167=>"111000000",
  14168=>"010000000",
  14169=>"111011011",
  14170=>"100111011",
  14171=>"110100001",
  14172=>"111000001",
  14173=>"001001011",
  14174=>"100010010",
  14175=>"101001100",
  14176=>"011010000",
  14177=>"000000110",
  14178=>"111000000",
  14179=>"000000110",
  14180=>"010010000",
  14181=>"001001000",
  14182=>"100111011",
  14183=>"111101000",
  14184=>"101011011",
  14185=>"010000110",
  14186=>"001111111",
  14187=>"111000001",
  14188=>"000001100",
  14189=>"000010010",
  14190=>"111000000",
  14191=>"011000111",
  14192=>"001011000",
  14193=>"010110111",
  14194=>"111111011",
  14195=>"000000000",
  14196=>"001001010",
  14197=>"000010000",
  14198=>"111010010",
  14199=>"111000000",
  14200=>"000010111",
  14201=>"111100000",
  14202=>"100101111",
  14203=>"000000101",
  14204=>"110010000",
  14205=>"100001110",
  14206=>"000000010",
  14207=>"000000000",
  14208=>"110010000",
  14209=>"000000111",
  14210=>"111000100",
  14211=>"110110010",
  14212=>"111111110",
  14213=>"111000010",
  14214=>"111110111",
  14215=>"000000100",
  14216=>"101111000",
  14217=>"000000000",
  14218=>"100011011",
  14219=>"111001011",
  14220=>"111000011",
  14221=>"000100111",
  14222=>"111111010",
  14223=>"000001000",
  14224=>"100100101",
  14225=>"000001101",
  14226=>"001010000",
  14227=>"000000101",
  14228=>"101011011",
  14229=>"011000000",
  14230=>"111010010",
  14231=>"110011000",
  14232=>"000010000",
  14233=>"101111011",
  14234=>"000000100",
  14235=>"000000101",
  14236=>"011111000",
  14237=>"111011000",
  14238=>"011111111",
  14239=>"000001111",
  14240=>"000101101",
  14241=>"100110111",
  14242=>"111010011",
  14243=>"000011101",
  14244=>"111011111",
  14245=>"000000000",
  14246=>"000010100",
  14247=>"100001011",
  14248=>"110010010",
  14249=>"011011000",
  14250=>"000000111",
  14251=>"000000111",
  14252=>"111010001",
  14253=>"011000000",
  14254=>"101111100",
  14255=>"010000000",
  14256=>"001010010",
  14257=>"110110000",
  14258=>"000100000",
  14259=>"110110000",
  14260=>"010000011",
  14261=>"101001111",
  14262=>"000100100",
  14263=>"000111111",
  14264=>"000100011",
  14265=>"101111000",
  14266=>"111011011",
  14267=>"011010000",
  14268=>"010111111",
  14269=>"111111100",
  14270=>"111000000",
  14271=>"000000100",
  14272=>"000100100",
  14273=>"111100000",
  14274=>"011111000",
  14275=>"000000000",
  14276=>"100110010",
  14277=>"001100100",
  14278=>"101011010",
  14279=>"000000010",
  14280=>"000010010",
  14281=>"100100101",
  14282=>"111101110",
  14283=>"111111011",
  14284=>"001011001",
  14285=>"011011000",
  14286=>"100000011",
  14287=>"111101100",
  14288=>"010011000",
  14289=>"110110001",
  14290=>"011001000",
  14291=>"111110111",
  14292=>"000000000",
  14293=>"100110011",
  14294=>"010010010",
  14295=>"001000000",
  14296=>"000010011",
  14297=>"000000111",
  14298=>"100101000",
  14299=>"000000101",
  14300=>"001101111",
  14301=>"101011010",
  14302=>"000100101",
  14303=>"010100010",
  14304=>"001000100",
  14305=>"000101000",
  14306=>"000000010",
  14307=>"111010000",
  14308=>"010000000",
  14309=>"101111111",
  14310=>"111000111",
  14311=>"100110010",
  14312=>"111111011",
  14313=>"010011111",
  14314=>"000000000",
  14315=>"000100111",
  14316=>"111001000",
  14317=>"010101111",
  14318=>"110000110",
  14319=>"000000000",
  14320=>"000011011",
  14321=>"100100101",
  14322=>"010100000",
  14323=>"011100110",
  14324=>"101001111",
  14325=>"001100010",
  14326=>"100100000",
  14327=>"000000000",
  14328=>"101101100",
  14329=>"111011010",
  14330=>"110100111",
  14331=>"110100101",
  14332=>"011011000",
  14333=>"100011111",
  14334=>"101111100",
  14335=>"010010000",
  14336=>"000000100",
  14337=>"101101111",
  14338=>"111100000",
  14339=>"000111010",
  14340=>"000110111",
  14341=>"110110101",
  14342=>"000000111",
  14343=>"011010111",
  14344=>"000000010",
  14345=>"010000000",
  14346=>"111101000",
  14347=>"001101000",
  14348=>"000000000",
  14349=>"001001000",
  14350=>"000100101",
  14351=>"111111111",
  14352=>"111000000",
  14353=>"111000011",
  14354=>"111111111",
  14355=>"000000000",
  14356=>"101000001",
  14357=>"100100111",
  14358=>"000000100",
  14359=>"110000110",
  14360=>"100101000",
  14361=>"001111111",
  14362=>"100100110",
  14363=>"111000000",
  14364=>"101001011",
  14365=>"000101010",
  14366=>"001000100",
  14367=>"000000000",
  14368=>"111111000",
  14369=>"101010010",
  14370=>"010110010",
  14371=>"010000100",
  14372=>"000001111",
  14373=>"100000001",
  14374=>"110001100",
  14375=>"111111110",
  14376=>"111111010",
  14377=>"100100000",
  14378=>"001000000",
  14379=>"111111000",
  14380=>"011011011",
  14381=>"010010000",
  14382=>"011010111",
  14383=>"000111010",
  14384=>"000110110",
  14385=>"010001111",
  14386=>"111111101",
  14387=>"010000000",
  14388=>"001001000",
  14389=>"000111000",
  14390=>"000000000",
  14391=>"000101111",
  14392=>"001111111",
  14393=>"101000100",
  14394=>"111001111",
  14395=>"111111111",
  14396=>"001000111",
  14397=>"111000010",
  14398=>"000000100",
  14399=>"110111111",
  14400=>"000000011",
  14401=>"001101001",
  14402=>"111111110",
  14403=>"111110110",
  14404=>"110000000",
  14405=>"100000000",
  14406=>"000011111",
  14407=>"111111010",
  14408=>"000000001",
  14409=>"111111100",
  14410=>"111000000",
  14411=>"000010111",
  14412=>"111111101",
  14413=>"110100101",
  14414=>"000000110",
  14415=>"000110110",
  14416=>"101101101",
  14417=>"110010000",
  14418=>"000000100",
  14419=>"000011001",
  14420=>"101101101",
  14421=>"000010100",
  14422=>"011000100",
  14423=>"110111011",
  14424=>"010000001",
  14425=>"110100111",
  14426=>"100110100",
  14427=>"011111111",
  14428=>"100000111",
  14429=>"000100000",
  14430=>"100010111",
  14431=>"010010011",
  14432=>"111111111",
  14433=>"101101110",
  14434=>"111000000",
  14435=>"001011011",
  14436=>"000000000",
  14437=>"001011111",
  14438=>"100111110",
  14439=>"101001000",
  14440=>"000111111",
  14441=>"000000010",
  14442=>"111100100",
  14443=>"001101000",
  14444=>"101001101",
  14445=>"110010010",
  14446=>"000000011",
  14447=>"110101111",
  14448=>"011101111",
  14449=>"000010100",
  14450=>"111000000",
  14451=>"110000000",
  14452=>"011110100",
  14453=>"111101101",
  14454=>"111000000",
  14455=>"010111111",
  14456=>"101101110",
  14457=>"011011000",
  14458=>"111111111",
  14459=>"010010111",
  14460=>"000000100",
  14461=>"000110000",
  14462=>"101010000",
  14463=>"101101001",
  14464=>"011110101",
  14465=>"011011000",
  14466=>"101001010",
  14467=>"000101001",
  14468=>"101000110",
  14469=>"000110011",
  14470=>"101001111",
  14471=>"011001001",
  14472=>"100100110",
  14473=>"111111110",
  14474=>"010010010",
  14475=>"111111011",
  14476=>"000000111",
  14477=>"111111100",
  14478=>"011010000",
  14479=>"111100000",
  14480=>"001100111",
  14481=>"000000110",
  14482=>"000000000",
  14483=>"000000000",
  14484=>"010000001",
  14485=>"111001000",
  14486=>"011011111",
  14487=>"000100111",
  14488=>"111111010",
  14489=>"110001000",
  14490=>"000101001",
  14491=>"000010000",
  14492=>"100101101",
  14493=>"010000000",
  14494=>"000101111",
  14495=>"110000000",
  14496=>"001011011",
  14497=>"010011111",
  14498=>"000000100",
  14499=>"111000000",
  14500=>"111000111",
  14501=>"010111110",
  14502=>"101000000",
  14503=>"010000110",
  14504=>"111000000",
  14505=>"000010001",
  14506=>"111111001",
  14507=>"111000000",
  14508=>"000000000",
  14509=>"010000000",
  14510=>"000101011",
  14511=>"010010000",
  14512=>"111110110",
  14513=>"101000111",
  14514=>"000000010",
  14515=>"010001000",
  14516=>"100011100",
  14517=>"000000000",
  14518=>"000111111",
  14519=>"000111111",
  14520=>"101000101",
  14521=>"010001110",
  14522=>"000101000",
  14523=>"001101101",
  14524=>"000100010",
  14525=>"010110100",
  14526=>"001011000",
  14527=>"111111111",
  14528=>"001100001",
  14529=>"111000111",
  14530=>"111111001",
  14531=>"110010001",
  14532=>"010111011",
  14533=>"000110100",
  14534=>"000000000",
  14535=>"111011010",
  14536=>"000001010",
  14537=>"000000000",
  14538=>"000111111",
  14539=>"101000100",
  14540=>"000100110",
  14541=>"100100000",
  14542=>"101101101",
  14543=>"000000011",
  14544=>"101101111",
  14545=>"000111111",
  14546=>"101101000",
  14547=>"010011111",
  14548=>"101011111",
  14549=>"101001011",
  14550=>"111101101",
  14551=>"000110111",
  14552=>"000000000",
  14553=>"100000010",
  14554=>"000110110",
  14555=>"101101101",
  14556=>"111101011",
  14557=>"111111111",
  14558=>"110111101",
  14559=>"111000100",
  14560=>"001000010",
  14561=>"111011011",
  14562=>"101010010",
  14563=>"000011111",
  14564=>"111000111",
  14565=>"000111111",
  14566=>"010001001",
  14567=>"001001111",
  14568=>"111011010",
  14569=>"101100111",
  14570=>"111100000",
  14571=>"000110110",
  14572=>"000000000",
  14573=>"001111111",
  14574=>"110000000",
  14575=>"000010000",
  14576=>"111000111",
  14577=>"010001001",
  14578=>"111000100",
  14579=>"000111011",
  14580=>"000000110",
  14581=>"101101101",
  14582=>"010010000",
  14583=>"101010000",
  14584=>"000000111",
  14585=>"011111111",
  14586=>"000011000",
  14587=>"101110001",
  14588=>"000110111",
  14589=>"000000011",
  14590=>"001011110",
  14591=>"111111111",
  14592=>"000000000",
  14593=>"000010010",
  14594=>"111000000",
  14595=>"101101010",
  14596=>"111111101",
  14597=>"110000111",
  14598=>"000111110",
  14599=>"110111111",
  14600=>"010010010",
  14601=>"101010010",
  14602=>"100110111",
  14603=>"100000000",
  14604=>"000000011",
  14605=>"101111001",
  14606=>"110011011",
  14607=>"000010101",
  14608=>"000110110",
  14609=>"000010011",
  14610=>"010000000",
  14611=>"000010111",
  14612=>"111011010",
  14613=>"101111111",
  14614=>"010111100",
  14615=>"011011011",
  14616=>"111000100",
  14617=>"000010000",
  14618=>"010001001",
  14619=>"000000000",
  14620=>"000001001",
  14621=>"000010100",
  14622=>"111011001",
  14623=>"000000101",
  14624=>"000100001",
  14625=>"011110111",
  14626=>"111101111",
  14627=>"000111111",
  14628=>"011100000",
  14629=>"101100001",
  14630=>"001101001",
  14631=>"000010010",
  14632=>"101011010",
  14633=>"001111111",
  14634=>"100010011",
  14635=>"000000100",
  14636=>"000101111",
  14637=>"111111010",
  14638=>"000111111",
  14639=>"010001101",
  14640=>"111111001",
  14641=>"111111100",
  14642=>"010001001",
  14643=>"111111010",
  14644=>"000000000",
  14645=>"000000110",
  14646=>"001000000",
  14647=>"000000000",
  14648=>"000011011",
  14649=>"000001001",
  14650=>"011000101",
  14651=>"011011010",
  14652=>"010110010",
  14653=>"011001000",
  14654=>"000100000",
  14655=>"110010110",
  14656=>"111010111",
  14657=>"100100111",
  14658=>"111011111",
  14659=>"100100011",
  14660=>"111000111",
  14661=>"000011011",
  14662=>"011011111",
  14663=>"000000000",
  14664=>"110101101",
  14665=>"000111111",
  14666=>"000000000",
  14667=>"101000010",
  14668=>"101000011",
  14669=>"000001010",
  14670=>"011001101",
  14671=>"111111111",
  14672=>"001000111",
  14673=>"101111000",
  14674=>"111111100",
  14675=>"001001100",
  14676=>"101000000",
  14677=>"000000000",
  14678=>"100111101",
  14679=>"100010010",
  14680=>"111000001",
  14681=>"110101100",
  14682=>"111100111",
  14683=>"000011110",
  14684=>"000010111",
  14685=>"000001001",
  14686=>"100010010",
  14687=>"001011111",
  14688=>"111010111",
  14689=>"000110111",
  14690=>"111000111",
  14691=>"110100101",
  14692=>"000101111",
  14693=>"000011111",
  14694=>"000010001",
  14695=>"000010011",
  14696=>"000100111",
  14697=>"111010000",
  14698=>"000110000",
  14699=>"000101000",
  14700=>"110111000",
  14701=>"000110111",
  14702=>"000110011",
  14703=>"101111100",
  14704=>"010111111",
  14705=>"100011101",
  14706=>"000000010",
  14707=>"000000000",
  14708=>"111101000",
  14709=>"011000101",
  14710=>"000000010",
  14711=>"000110111",
  14712=>"111000100",
  14713=>"000111100",
  14714=>"110000011",
  14715=>"000011010",
  14716=>"010100010",
  14717=>"100100000",
  14718=>"001101111",
  14719=>"111101111",
  14720=>"100100111",
  14721=>"010000000",
  14722=>"001111010",
  14723=>"000101101",
  14724=>"000111000",
  14725=>"111101101",
  14726=>"001011110",
  14727=>"100000010",
  14728=>"100111011",
  14729=>"101011000",
  14730=>"000011001",
  14731=>"010110011",
  14732=>"100000110",
  14733=>"000000111",
  14734=>"000111111",
  14735=>"001100111",
  14736=>"011001101",
  14737=>"010000111",
  14738=>"111000000",
  14739=>"000010010",
  14740=>"000100111",
  14741=>"000010010",
  14742=>"111111000",
  14743=>"100101101",
  14744=>"100100111",
  14745=>"010000101",
  14746=>"111101101",
  14747=>"110101100",
  14748=>"000000000",
  14749=>"101000000",
  14750=>"001110000",
  14751=>"000010000",
  14752=>"100101000",
  14753=>"010010000",
  14754=>"000111010",
  14755=>"111010101",
  14756=>"000110100",
  14757=>"000000011",
  14758=>"000111011",
  14759=>"000101111",
  14760=>"100011110",
  14761=>"101000010",
  14762=>"111101101",
  14763=>"000000100",
  14764=>"111010011",
  14765=>"100011011",
  14766=>"111101111",
  14767=>"101010110",
  14768=>"111000000",
  14769=>"011001111",
  14770=>"000001111",
  14771=>"011001000",
  14772=>"000100111",
  14773=>"111101001",
  14774=>"111100101",
  14775=>"000011011",
  14776=>"000011000",
  14777=>"001011001",
  14778=>"000101000",
  14779=>"011111010",
  14780=>"001000101",
  14781=>"111000000",
  14782=>"011000011",
  14783=>"000110101",
  14784=>"000010000",
  14785=>"000110111",
  14786=>"101101011",
  14787=>"000001100",
  14788=>"111000111",
  14789=>"110110000",
  14790=>"011110000",
  14791=>"000111111",
  14792=>"100010011",
  14793=>"000000101",
  14794=>"000000001",
  14795=>"100101000",
  14796=>"000000001",
  14797=>"000010010",
  14798=>"010000110",
  14799=>"111010001",
  14800=>"010000000",
  14801=>"000001001",
  14802=>"100000000",
  14803=>"010010010",
  14804=>"110111110",
  14805=>"000000110",
  14806=>"011010000",
  14807=>"101111011",
  14808=>"001101111",
  14809=>"000000101",
  14810=>"011001101",
  14811=>"111000010",
  14812=>"010110000",
  14813=>"000010111",
  14814=>"011011111",
  14815=>"101111001",
  14816=>"101000111",
  14817=>"111011010",
  14818=>"111000111",
  14819=>"011111110",
  14820=>"000000010",
  14821=>"111001000",
  14822=>"111111001",
  14823=>"100011111",
  14824=>"001100110",
  14825=>"110110000",
  14826=>"001111111",
  14827=>"010011111",
  14828=>"101000000",
  14829=>"111100111",
  14830=>"001000000",
  14831=>"000100100",
  14832=>"011111010",
  14833=>"011011001",
  14834=>"111111111",
  14835=>"000001101",
  14836=>"000100100",
  14837=>"111101101",
  14838=>"101000010",
  14839=>"111000000",
  14840=>"100000010",
  14841=>"010110011",
  14842=>"000000100",
  14843=>"000000000",
  14844=>"111101001",
  14845=>"010111000",
  14846=>"000100111",
  14847=>"110111110",
  14848=>"000001000",
  14849=>"000000100",
  14850=>"111000000",
  14851=>"111111111",
  14852=>"000000011",
  14853=>"000001110",
  14854=>"111000101",
  14855=>"000101111",
  14856=>"101111111",
  14857=>"101101111",
  14858=>"000000000",
  14859=>"011000001",
  14860=>"111011000",
  14861=>"011011000",
  14862=>"011101001",
  14863=>"000111111",
  14864=>"001011000",
  14865=>"000000000",
  14866=>"100000000",
  14867=>"000000001",
  14868=>"101000111",
  14869=>"101100000",
  14870=>"001111111",
  14871=>"100100111",
  14872=>"000000000",
  14873=>"000010000",
  14874=>"000000000",
  14875=>"001000000",
  14876=>"000000100",
  14877=>"000000000",
  14878=>"110111001",
  14879=>"000111001",
  14880=>"111111111",
  14881=>"101111011",
  14882=>"001111001",
  14883=>"111111111",
  14884=>"000000000",
  14885=>"001101111",
  14886=>"111100000",
  14887=>"100110010",
  14888=>"000111111",
  14889=>"101111001",
  14890=>"000000000",
  14891=>"011111111",
  14892=>"001011001",
  14893=>"101111000",
  14894=>"101111111",
  14895=>"000000100",
  14896=>"000000000",
  14897=>"110110010",
  14898=>"001111111",
  14899=>"000110000",
  14900=>"000000000",
  14901=>"000000000",
  14902=>"001000000",
  14903=>"000110100",
  14904=>"111111111",
  14905=>"000000000",
  14906=>"000000000",
  14907=>"000100111",
  14908=>"111011111",
  14909=>"111111001",
  14910=>"000000100",
  14911=>"111111110",
  14912=>"000000001",
  14913=>"000111101",
  14914=>"000101011",
  14915=>"010110011",
  14916=>"111111000",
  14917=>"000000000",
  14918=>"101101000",
  14919=>"111111111",
  14920=>"010111101",
  14921=>"111111110",
  14922=>"000000000",
  14923=>"000000000",
  14924=>"111100001",
  14925=>"000010000",
  14926=>"011100101",
  14927=>"111111111",
  14928=>"000000000",
  14929=>"111111110",
  14930=>"101111111",
  14931=>"111011000",
  14932=>"111001110",
  14933=>"010100110",
  14934=>"001100000",
  14935=>"100010000",
  14936=>"010000010",
  14937=>"011001001",
  14938=>"100110000",
  14939=>"110010010",
  14940=>"111000000",
  14941=>"001011111",
  14942=>"111111111",
  14943=>"011001000",
  14944=>"010101100",
  14945=>"111110011",
  14946=>"110000000",
  14947=>"000100000",
  14948=>"100000000",
  14949=>"000000000",
  14950=>"111111111",
  14951=>"100100000",
  14952=>"100101111",
  14953=>"000000000",
  14954=>"000100111",
  14955=>"111111111",
  14956=>"111010111",
  14957=>"000000000",
  14958=>"000010010",
  14959=>"000000110",
  14960=>"001011001",
  14961=>"000000111",
  14962=>"001001000",
  14963=>"000000000",
  14964=>"111110000",
  14965=>"000000100",
  14966=>"110000000",
  14967=>"101111101",
  14968=>"101000111",
  14969=>"111011111",
  14970=>"000111010",
  14971=>"111111111",
  14972=>"110110000",
  14973=>"110111001",
  14974=>"101101110",
  14975=>"110000111",
  14976=>"000111000",
  14977=>"111111010",
  14978=>"111111111",
  14979=>"011111111",
  14980=>"010000000",
  14981=>"001000000",
  14982=>"000110101",
  14983=>"001011001",
  14984=>"101101100",
  14985=>"000000000",
  14986=>"000000000",
  14987=>"101101000",
  14988=>"001000101",
  14989=>"001111111",
  14990=>"100000000",
  14991=>"000000000",
  14992=>"000001001",
  14993=>"111111111",
  14994=>"000000000",
  14995=>"001111111",
  14996=>"001001100",
  14997=>"000110000",
  14998=>"000001001",
  14999=>"100101101",
  15000=>"101111111",
  15001=>"001001111",
  15002=>"010011000",
  15003=>"110100101",
  15004=>"111011000",
  15005=>"011000000",
  15006=>"111101111",
  15007=>"001010111",
  15008=>"011011011",
  15009=>"000000110",
  15010=>"000101111",
  15011=>"101100101",
  15012=>"100110000",
  15013=>"110110000",
  15014=>"001100000",
  15015=>"000011111",
  15016=>"000000111",
  15017=>"101100101",
  15018=>"000010010",
  15019=>"000000000",
  15020=>"111111011",
  15021=>"111101100",
  15022=>"111011111",
  15023=>"111111010",
  15024=>"111111111",
  15025=>"000010000",
  15026=>"110101111",
  15027=>"110100110",
  15028=>"100110000",
  15029=>"111111111",
  15030=>"100001101",
  15031=>"000011111",
  15032=>"111100111",
  15033=>"100100000",
  15034=>"110011000",
  15035=>"111111111",
  15036=>"000010001",
  15037=>"111111111",
  15038=>"111111111",
  15039=>"011100000",
  15040=>"011000100",
  15041=>"000001001",
  15042=>"101111011",
  15043=>"000101001",
  15044=>"000000000",
  15045=>"100101110",
  15046=>"000011111",
  15047=>"001000110",
  15048=>"100111101",
  15049=>"000000100",
  15050=>"110001101",
  15051=>"000000000",
  15052=>"101100101",
  15053=>"111001001",
  15054=>"000000000",
  15055=>"111111000",
  15056=>"111001000",
  15057=>"011111001",
  15058=>"001000010",
  15059=>"000000001",
  15060=>"111110111",
  15061=>"000000101",
  15062=>"111111010",
  15063=>"000000001",
  15064=>"001111101",
  15065=>"111111111",
  15066=>"110110101",
  15067=>"000000000",
  15068=>"000001010",
  15069=>"111110111",
  15070=>"000000000",
  15071=>"001101111",
  15072=>"111101001",
  15073=>"000000000",
  15074=>"111111110",
  15075=>"000110010",
  15076=>"000000000",
  15077=>"011001001",
  15078=>"011011101",
  15079=>"111111111",
  15080=>"110101111",
  15081=>"100101111",
  15082=>"000000000",
  15083=>"100000010",
  15084=>"110001010",
  15085=>"000000000",
  15086=>"111111110",
  15087=>"111111001",
  15088=>"000110110",
  15089=>"001011111",
  15090=>"111111111",
  15091=>"111111001",
  15092=>"001011011",
  15093=>"000000000",
  15094=>"000011111",
  15095=>"000011011",
  15096=>"010111111",
  15097=>"001111111",
  15098=>"111111111",
  15099=>"000011000",
  15100=>"000001001",
  15101=>"111111111",
  15102=>"000001101",
  15103=>"000010000",
  15104=>"001100100",
  15105=>"111001000",
  15106=>"111101111",
  15107=>"010111111",
  15108=>"011111000",
  15109=>"110101111",
  15110=>"000000000",
  15111=>"110110111",
  15112=>"100000101",
  15113=>"100111111",
  15114=>"111011100",
  15115=>"111111000",
  15116=>"111000101",
  15117=>"001000000",
  15118=>"111100000",
  15119=>"000001100",
  15120=>"010000001",
  15121=>"101000000",
  15122=>"110111001",
  15123=>"000000010",
  15124=>"111000100",
  15125=>"111001101",
  15126=>"111111011",
  15127=>"000010111",
  15128=>"001110000",
  15129=>"000111111",
  15130=>"000000010",
  15131=>"000111000",
  15132=>"111100101",
  15133=>"000000010",
  15134=>"100000010",
  15135=>"111101101",
  15136=>"111110000",
  15137=>"011010111",
  15138=>"010111100",
  15139=>"111111111",
  15140=>"010011111",
  15141=>"000111101",
  15142=>"111000000",
  15143=>"010101000",
  15144=>"010111111",
  15145=>"111000100",
  15146=>"010001001",
  15147=>"010111111",
  15148=>"011011011",
  15149=>"000001011",
  15150=>"010000010",
  15151=>"000110101",
  15152=>"000011011",
  15153=>"111111111",
  15154=>"000000100",
  15155=>"001010111",
  15156=>"000000000",
  15157=>"111111111",
  15158=>"111011001",
  15159=>"101000000",
  15160=>"000000010",
  15161=>"111001000",
  15162=>"100000000",
  15163=>"000111111",
  15164=>"111101001",
  15165=>"111111111",
  15166=>"100000000",
  15167=>"111110111",
  15168=>"000111111",
  15169=>"000001110",
  15170=>"000000111",
  15171=>"000000000",
  15172=>"100010010",
  15173=>"000101111",
  15174=>"000011010",
  15175=>"111101111",
  15176=>"000100010",
  15177=>"000000000",
  15178=>"110111111",
  15179=>"111001111",
  15180=>"000001000",
  15181=>"000111011",
  15182=>"111111111",
  15183=>"010101000",
  15184=>"000100101",
  15185=>"111110101",
  15186=>"000000101",
  15187=>"101110010",
  15188=>"000000111",
  15189=>"111001001",
  15190=>"111110110",
  15191=>"010000000",
  15192=>"000000001",
  15193=>"111001000",
  15194=>"000000000",
  15195=>"101011000",
  15196=>"111101101",
  15197=>"111010100",
  15198=>"000111111",
  15199=>"100000000",
  15200=>"111000000",
  15201=>"000111111",
  15202=>"000011011",
  15203=>"100000000",
  15204=>"011101001",
  15205=>"000100100",
  15206=>"101000000",
  15207=>"111100000",
  15208=>"111111111",
  15209=>"001011111",
  15210=>"010111111",
  15211=>"111000100",
  15212=>"101110110",
  15213=>"001111111",
  15214=>"101000000",
  15215=>"000000000",
  15216=>"000001101",
  15217=>"100000000",
  15218=>"100110000",
  15219=>"111000000",
  15220=>"000000000",
  15221=>"101100111",
  15222=>"111000000",
  15223=>"101000000",
  15224=>"111101001",
  15225=>"111111111",
  15226=>"111001000",
  15227=>"000111111",
  15228=>"000000010",
  15229=>"111011010",
  15230=>"110100111",
  15231=>"000011111",
  15232=>"000011111",
  15233=>"000000111",
  15234=>"000001000",
  15235=>"011111111",
  15236=>"001001000",
  15237=>"110001010",
  15238=>"000100110",
  15239=>"001010000",
  15240=>"100110011",
  15241=>"000111111",
  15242=>"110111000",
  15243=>"011100110",
  15244=>"111000000",
  15245=>"000101101",
  15246=>"000111111",
  15247=>"000000000",
  15248=>"001011000",
  15249=>"010000001",
  15250=>"111101000",
  15251=>"111101011",
  15252=>"000100000",
  15253=>"111000000",
  15254=>"000010000",
  15255=>"100000000",
  15256=>"001000000",
  15257=>"000010111",
  15258=>"010111111",
  15259=>"000111000",
  15260=>"111100000",
  15261=>"000111111",
  15262=>"000101111",
  15263=>"111000000",
  15264=>"011111100",
  15265=>"011010000",
  15266=>"010000000",
  15267=>"000000100",
  15268=>"101000000",
  15269=>"011011000",
  15270=>"110100101",
  15271=>"000010000",
  15272=>"000110000",
  15273=>"010111000",
  15274=>"000000000",
  15275=>"100000000",
  15276=>"011001001",
  15277=>"000011111",
  15278=>"000000010",
  15279=>"000111111",
  15280=>"000000111",
  15281=>"001100000",
  15282=>"001111111",
  15283=>"110111001",
  15284=>"111011000",
  15285=>"010000000",
  15286=>"011101000",
  15287=>"101100000",
  15288=>"111001000",
  15289=>"101011001",
  15290=>"010000000",
  15291=>"010100000",
  15292=>"111101000",
  15293=>"000111111",
  15294=>"110111011",
  15295=>"000000000",
  15296=>"000010111",
  15297=>"000000111",
  15298=>"010111000",
  15299=>"100000000",
  15300=>"111111000",
  15301=>"001001001",
  15302=>"000000001",
  15303=>"100100111",
  15304=>"001000101",
  15305=>"001101111",
  15306=>"111101001",
  15307=>"100000000",
  15308=>"010000000",
  15309=>"000010000",
  15310=>"111100000",
  15311=>"100011010",
  15312=>"111011010",
  15313=>"010111110",
  15314=>"000001000",
  15315=>"010111110",
  15316=>"001000110",
  15317=>"101000000",
  15318=>"011000000",
  15319=>"010001111",
  15320=>"111100101",
  15321=>"111111000",
  15322=>"100111001",
  15323=>"000111111",
  15324=>"111111100",
  15325=>"010011001",
  15326=>"001000000",
  15327=>"111111111",
  15328=>"011111111",
  15329=>"000000011",
  15330=>"000000000",
  15331=>"100011111",
  15332=>"101000000",
  15333=>"000111111",
  15334=>"111111101",
  15335=>"001000010",
  15336=>"111111001",
  15337=>"110111110",
  15338=>"011100000",
  15339=>"000000000",
  15340=>"111000000",
  15341=>"101101111",
  15342=>"110000010",
  15343=>"001000000",
  15344=>"111010000",
  15345=>"110100000",
  15346=>"000000100",
  15347=>"111111000",
  15348=>"101011011",
  15349=>"000000000",
  15350=>"000101010",
  15351=>"110100000",
  15352=>"011000000",
  15353=>"000010111",
  15354=>"110100000",
  15355=>"010111000",
  15356=>"100000000",
  15357=>"010111111",
  15358=>"110110110",
  15359=>"110101001",
  15360=>"000000111",
  15361=>"000000001",
  15362=>"111111000",
  15363=>"111010000",
  15364=>"000000110",
  15365=>"000001111",
  15366=>"000111111",
  15367=>"000000000",
  15368=>"000000000",
  15369=>"111111000",
  15370=>"001011011",
  15371=>"011001000",
  15372=>"011001101",
  15373=>"000000000",
  15374=>"010010100",
  15375=>"000000000",
  15376=>"110000111",
  15377=>"111000010",
  15378=>"111110110",
  15379=>"000001011",
  15380=>"111101100",
  15381=>"001000101",
  15382=>"000110010",
  15383=>"001000101",
  15384=>"000001001",
  15385=>"110111101",
  15386=>"000000000",
  15387=>"111110000",
  15388=>"011011101",
  15389=>"000000000",
  15390=>"111001010",
  15391=>"110100111",
  15392=>"111110010",
  15393=>"010100000",
  15394=>"000001001",
  15395=>"011111001",
  15396=>"010000011",
  15397=>"000000000",
  15398=>"100100101",
  15399=>"111001001",
  15400=>"111111111",
  15401=>"000000100",
  15402=>"000000111",
  15403=>"011111001",
  15404=>"010111011",
  15405=>"000000000",
  15406=>"011111111",
  15407=>"011000000",
  15408=>"000000110",
  15409=>"011000110",
  15410=>"000000000",
  15411=>"000111111",
  15412=>"101100111",
  15413=>"101101001",
  15414=>"000011001",
  15415=>"000111111",
  15416=>"000000000",
  15417=>"000000111",
  15418=>"001001000",
  15419=>"000000000",
  15420=>"000000000",
  15421=>"111111111",
  15422=>"001001101",
  15423=>"100100110",
  15424=>"000000010",
  15425=>"111001000",
  15426=>"010110010",
  15427=>"000100110",
  15428=>"000000000",
  15429=>"000000000",
  15430=>"010111111",
  15431=>"001001111",
  15432=>"000000010",
  15433=>"111000111",
  15434=>"001101101",
  15435=>"111000011",
  15436=>"010111111",
  15437=>"111011010",
  15438=>"000010110",
  15439=>"000111110",
  15440=>"110110110",
  15441=>"111111000",
  15442=>"001001111",
  15443=>"010110011",
  15444=>"110101101",
  15445=>"011000000",
  15446=>"111010010",
  15447=>"111111000",
  15448=>"000110111",
  15449=>"000010111",
  15450=>"011111111",
  15451=>"111111110",
  15452=>"111110010",
  15453=>"001011001",
  15454=>"110100111",
  15455=>"000111010",
  15456=>"010011000",
  15457=>"010010000",
  15458=>"011001101",
  15459=>"110111110",
  15460=>"000000110",
  15461=>"011010000",
  15462=>"101100110",
  15463=>"111111000",
  15464=>"000001111",
  15465=>"000000001",
  15466=>"000000000",
  15467=>"000001111",
  15468=>"000001000",
  15469=>"000000010",
  15470=>"011000000",
  15471=>"010000000",
  15472=>"010110110",
  15473=>"000001000",
  15474=>"000000110",
  15475=>"110011111",
  15476=>"101000111",
  15477=>"101001111",
  15478=>"010111111",
  15479=>"000010001",
  15480=>"111111101",
  15481=>"000000000",
  15482=>"001000000",
  15483=>"000000010",
  15484=>"010000000",
  15485=>"111111110",
  15486=>"000000000",
  15487=>"111111111",
  15488=>"100111110",
  15489=>"000000000",
  15490=>"000000000",
  15491=>"000000000",
  15492=>"011110111",
  15493=>"000000111",
  15494=>"000000000",
  15495=>"001000000",
  15496=>"001011001",
  15497=>"000001101",
  15498=>"000001010",
  15499=>"011111111",
  15500=>"111111011",
  15501=>"010111010",
  15502=>"000000000",
  15503=>"111000101",
  15504=>"111111111",
  15505=>"010010010",
  15506=>"001000101",
  15507=>"011101110",
  15508=>"000101101",
  15509=>"010000000",
  15510=>"100100100",
  15511=>"000000001",
  15512=>"110000000",
  15513=>"111111101",
  15514=>"001000101",
  15515=>"111110000",
  15516=>"110000010",
  15517=>"011110010",
  15518=>"000000111",
  15519=>"110111110",
  15520=>"000000010",
  15521=>"000000000",
  15522=>"001001000",
  15523=>"000010000",
  15524=>"000000100",
  15525=>"000000000",
  15526=>"000001001",
  15527=>"100000111",
  15528=>"000011011",
  15529=>"000001001",
  15530=>"111101100",
  15531=>"100110110",
  15532=>"111111011",
  15533=>"111111111",
  15534=>"001011011",
  15535=>"111111110",
  15536=>"111111111",
  15537=>"000000110",
  15538=>"000010010",
  15539=>"011000000",
  15540=>"010000010",
  15541=>"000000111",
  15542=>"111110100",
  15543=>"110010000",
  15544=>"000000000",
  15545=>"001010101",
  15546=>"000000000",
  15547=>"100000110",
  15548=>"001101111",
  15549=>"000111111",
  15550=>"000001001",
  15551=>"000100000",
  15552=>"111111111",
  15553=>"000010111",
  15554=>"000000000",
  15555=>"000010000",
  15556=>"001001101",
  15557=>"010000001",
  15558=>"000000001",
  15559=>"111111111",
  15560=>"001001101",
  15561=>"000000001",
  15562=>"111111111",
  15563=>"000000000",
  15564=>"011110111",
  15565=>"001011000",
  15566=>"111001100",
  15567=>"011001111",
  15568=>"111111111",
  15569=>"110110110",
  15570=>"111110101",
  15571=>"011101111",
  15572=>"111111111",
  15573=>"001011011",
  15574=>"111111111",
  15575=>"110111111",
  15576=>"001000001",
  15577=>"000110010",
  15578=>"000000100",
  15579=>"111100000",
  15580=>"001111110",
  15581=>"111111001",
  15582=>"010111111",
  15583=>"000000000",
  15584=>"110000001",
  15585=>"111111111",
  15586=>"111000000",
  15587=>"011111011",
  15588=>"001000000",
  15589=>"010111010",
  15590=>"001000000",
  15591=>"100110110",
  15592=>"000000000",
  15593=>"000101000",
  15594=>"100100110",
  15595=>"111111110",
  15596=>"000000000",
  15597=>"011111011",
  15598=>"010010000",
  15599=>"001000001",
  15600=>"001001101",
  15601=>"000000100",
  15602=>"011111111",
  15603=>"100001101",
  15604=>"001001011",
  15605=>"110111111",
  15606=>"110111110",
  15607=>"011000000",
  15608=>"001000001",
  15609=>"000101000",
  15610=>"111000001",
  15611=>"101111111",
  15612=>"111100111",
  15613=>"010000000",
  15614=>"000000000",
  15615=>"000111111",
  15616=>"011011011",
  15617=>"001111110",
  15618=>"101000000",
  15619=>"100111000",
  15620=>"001001110",
  15621=>"000000110",
  15622=>"000000010",
  15623=>"000100100",
  15624=>"000000000",
  15625=>"011001111",
  15626=>"001001011",
  15627=>"111101010",
  15628=>"101100110",
  15629=>"111111001",
  15630=>"001000001",
  15631=>"001111111",
  15632=>"000001110",
  15633=>"010000101",
  15634=>"000111100",
  15635=>"111000000",
  15636=>"110000000",
  15637=>"111110010",
  15638=>"111111011",
  15639=>"001000111",
  15640=>"001100111",
  15641=>"011000001",
  15642=>"010001111",
  15643=>"011001001",
  15644=>"001000100",
  15645=>"100000100",
  15646=>"111000000",
  15647=>"000110111",
  15648=>"000000000",
  15649=>"000001111",
  15650=>"111111111",
  15651=>"111110110",
  15652=>"001011111",
  15653=>"110010111",
  15654=>"110110010",
  15655=>"101010101",
  15656=>"110011000",
  15657=>"110110000",
  15658=>"001000111",
  15659=>"010000000",
  15660=>"111100000",
  15661=>"111011101",
  15662=>"101001000",
  15663=>"011111100",
  15664=>"000000001",
  15665=>"011100011",
  15666=>"101111001",
  15667=>"100000000",
  15668=>"000000000",
  15669=>"111101000",
  15670=>"100010111",
  15671=>"000111100",
  15672=>"111111010",
  15673=>"001000101",
  15674=>"000101000",
  15675=>"110111111",
  15676=>"110001000",
  15677=>"010111010",
  15678=>"000000101",
  15679=>"000000000",
  15680=>"100101101",
  15681=>"111110010",
  15682=>"110001000",
  15683=>"011000000",
  15684=>"011110000",
  15685=>"101000000",
  15686=>"000000001",
  15687=>"110000010",
  15688=>"111111111",
  15689=>"001001000",
  15690=>"000001001",
  15691=>"001000101",
  15692=>"111110110",
  15693=>"110111100",
  15694=>"010110001",
  15695=>"110111111",
  15696=>"000000000",
  15697=>"010011111",
  15698=>"111000001",
  15699=>"011001011",
  15700=>"001000011",
  15701=>"110111110",
  15702=>"111111011",
  15703=>"000000000",
  15704=>"000000111",
  15705=>"100001000",
  15706=>"001111101",
  15707=>"010100000",
  15708=>"100110110",
  15709=>"000011111",
  15710=>"111111111",
  15711=>"110000000",
  15712=>"000000000",
  15713=>"000000001",
  15714=>"001001011",
  15715=>"111110000",
  15716=>"100111111",
  15717=>"110011100",
  15718=>"001001111",
  15719=>"110110000",
  15720=>"000000000",
  15721=>"110000101",
  15722=>"000111101",
  15723=>"111110000",
  15724=>"110110101",
  15725=>"000000001",
  15726=>"111111000",
  15727=>"000100110",
  15728=>"011101101",
  15729=>"000000000",
  15730=>"001100111",
  15731=>"111000000",
  15732=>"001100110",
  15733=>"000001000",
  15734=>"000001001",
  15735=>"111110001",
  15736=>"011011111",
  15737=>"110010010",
  15738=>"111111001",
  15739=>"101000000",
  15740=>"010111101",
  15741=>"100100100",
  15742=>"110000000",
  15743=>"001001000",
  15744=>"110101110",
  15745=>"100100001",
  15746=>"111001011",
  15747=>"111101111",
  15748=>"011111101",
  15749=>"000000000",
  15750=>"110100111",
  15751=>"000001010",
  15752=>"100111011",
  15753=>"001000000",
  15754=>"000000111",
  15755=>"010000000",
  15756=>"000000100",
  15757=>"101000000",
  15758=>"000101011",
  15759=>"011000000",
  15760=>"111111111",
  15761=>"010110110",
  15762=>"000000010",
  15763=>"001000000",
  15764=>"000000000",
  15765=>"010000000",
  15766=>"001111111",
  15767=>"010011101",
  15768=>"111111111",
  15769=>"001110110",
  15770=>"110000000",
  15771=>"001001000",
  15772=>"000000000",
  15773=>"001001011",
  15774=>"110111111",
  15775=>"111010000",
  15776=>"100101110",
  15777=>"000110110",
  15778=>"100000001",
  15779=>"001001011",
  15780=>"110000011",
  15781=>"110111100",
  15782=>"110110000",
  15783=>"111001101",
  15784=>"110000000",
  15785=>"000110111",
  15786=>"101001111",
  15787=>"011000001",
  15788=>"001001011",
  15789=>"000000011",
  15790=>"100100100",
  15791=>"110100100",
  15792=>"000001001",
  15793=>"000111011",
  15794=>"000000000",
  15795=>"000000011",
  15796=>"111111111",
  15797=>"000000011",
  15798=>"111111111",
  15799=>"111110010",
  15800=>"011101001",
  15801=>"110011100",
  15802=>"111010110",
  15803=>"011001001",
  15804=>"100010000",
  15805=>"000110111",
  15806=>"000000001",
  15807=>"010111111",
  15808=>"000000111",
  15809=>"000000100",
  15810=>"101000010",
  15811=>"010111010",
  15812=>"011000000",
  15813=>"001001111",
  15814=>"100000000",
  15815=>"101010111",
  15816=>"101101001",
  15817=>"110111000",
  15818=>"001101111",
  15819=>"001101001",
  15820=>"001001000",
  15821=>"110101011",
  15822=>"001101010",
  15823=>"001111001",
  15824=>"111111000",
  15825=>"100111010",
  15826=>"001010000",
  15827=>"111111011",
  15828=>"111000001",
  15829=>"001100110",
  15830=>"111110110",
  15831=>"111111111",
  15832=>"111110010",
  15833=>"111111111",
  15834=>"110100000",
  15835=>"001000001",
  15836=>"110111001",
  15837=>"111010000",
  15838=>"111110000",
  15839=>"111111000",
  15840=>"001000101",
  15841=>"001001001",
  15842=>"111111101",
  15843=>"000000101",
  15844=>"001000110",
  15845=>"110010000",
  15846=>"101011000",
  15847=>"001001011",
  15848=>"111100100",
  15849=>"010010110",
  15850=>"001000001",
  15851=>"001001011",
  15852=>"010100000",
  15853=>"110110100",
  15854=>"110000000",
  15855=>"100110011",
  15856=>"000000000",
  15857=>"010100111",
  15858=>"111011110",
  15859=>"010011110",
  15860=>"100100100",
  15861=>"001001111",
  15862=>"000000010",
  15863=>"001001101",
  15864=>"001000000",
  15865=>"000001111",
  15866=>"001111111",
  15867=>"011111111",
  15868=>"001011001",
  15869=>"000000000",
  15870=>"000110111",
  15871=>"000000001",
  15872=>"011011111",
  15873=>"100101011",
  15874=>"001001011",
  15875=>"000011101",
  15876=>"100010100",
  15877=>"000000111",
  15878=>"011111010",
  15879=>"100010111",
  15880=>"000110111",
  15881=>"000100000",
  15882=>"000100100",
  15883=>"110000111",
  15884=>"110110100",
  15885=>"011001100",
  15886=>"011000110",
  15887=>"000000000",
  15888=>"000110110",
  15889=>"011000111",
  15890=>"001011100",
  15891=>"111001010",
  15892=>"011111111",
  15893=>"101001101",
  15894=>"110111111",
  15895=>"111110111",
  15896=>"001011111",
  15897=>"001110110",
  15898=>"000111010",
  15899=>"100110000",
  15900=>"001001101",
  15901=>"110100000",
  15902=>"000011001",
  15903=>"110110000",
  15904=>"001010111",
  15905=>"110111011",
  15906=>"111001010",
  15907=>"110100111",
  15908=>"111011000",
  15909=>"000000000",
  15910=>"001011111",
  15911=>"101000000",
  15912=>"011111111",
  15913=>"011111110",
  15914=>"000000001",
  15915=>"010110100",
  15916=>"100110001",
  15917=>"100110100",
  15918=>"001001101",
  15919=>"111111110",
  15920=>"111000100",
  15921=>"111011011",
  15922=>"100001000",
  15923=>"110000100",
  15924=>"110100000",
  15925=>"000100000",
  15926=>"100100100",
  15927=>"000100100",
  15928=>"000011011",
  15929=>"000000000",
  15930=>"100000000",
  15931=>"100001000",
  15932=>"110110110",
  15933=>"110011011",
  15934=>"000000001",
  15935=>"100000010",
  15936=>"011011111",
  15937=>"000010011",
  15938=>"110100100",
  15939=>"011000000",
  15940=>"001011000",
  15941=>"000000010",
  15942=>"100100000",
  15943=>"001111001",
  15944=>"000000000",
  15945=>"110010100",
  15946=>"010011111",
  15947=>"010001001",
  15948=>"001001110",
  15949=>"000000100",
  15950=>"001000000",
  15951=>"111111110",
  15952=>"011011010",
  15953=>"101111110",
  15954=>"100100000",
  15955=>"101101001",
  15956=>"111001000",
  15957=>"001101111",
  15958=>"100000101",
  15959=>"010110000",
  15960=>"010111110",
  15961=>"111100000",
  15962=>"101110100",
  15963=>"100010001",
  15964=>"000010100",
  15965=>"011100010",
  15966=>"101111010",
  15967=>"101111111",
  15968=>"000011111",
  15969=>"111011000",
  15970=>"011010101",
  15971=>"110111011",
  15972=>"100100100",
  15973=>"100100110",
  15974=>"110000000",
  15975=>"011111011",
  15976=>"011010110",
  15977=>"000000000",
  15978=>"110000110",
  15979=>"101110101",
  15980=>"011011110",
  15981=>"011000000",
  15982=>"100000000",
  15983=>"100000001",
  15984=>"001101100",
  15985=>"100100000",
  15986=>"100000110",
  15987=>"000000110",
  15988=>"000000000",
  15989=>"000011001",
  15990=>"111101001",
  15991=>"100011010",
  15992=>"110111111",
  15993=>"110100001",
  15994=>"011000111",
  15995=>"111001010",
  15996=>"110010100",
  15997=>"000000101",
  15998=>"100100111",
  15999=>"111000000",
  16000=>"001001000",
  16001=>"111001000",
  16002=>"101111000",
  16003=>"100111111",
  16004=>"110010100",
  16005=>"011100000",
  16006=>"001010110",
  16007=>"110011111",
  16008=>"010111111",
  16009=>"001100100",
  16010=>"100100010",
  16011=>"001010001",
  16012=>"000111110",
  16013=>"000000100",
  16014=>"001100000",
  16015=>"010000000",
  16016=>"100100110",
  16017=>"100100000",
  16018=>"000000001",
  16019=>"011011111",
  16020=>"110111010",
  16021=>"001000000",
  16022=>"000100000",
  16023=>"100000110",
  16024=>"110100110",
  16025=>"011111011",
  16026=>"001011111",
  16027=>"001100100",
  16028=>"110100000",
  16029=>"011011100",
  16030=>"000101100",
  16031=>"111001111",
  16032=>"100100001",
  16033=>"010010100",
  16034=>"011110111",
  16035=>"001011111",
  16036=>"011010110",
  16037=>"000100100",
  16038=>"111011010",
  16039=>"000110110",
  16040=>"111110000",
  16041=>"100111110",
  16042=>"001001001",
  16043=>"011011011",
  16044=>"001111111",
  16045=>"010100000",
  16046=>"010000000",
  16047=>"100100101",
  16048=>"010100100",
  16049=>"011110111",
  16050=>"001010000",
  16051=>"000000110",
  16052=>"111111111",
  16053=>"111100000",
  16054=>"100000100",
  16055=>"011100001",
  16056=>"111000010",
  16057=>"100110000",
  16058=>"100000000",
  16059=>"010111111",
  16060=>"100100010",
  16061=>"001001110",
  16062=>"111111111",
  16063=>"110010000",
  16064=>"001000000",
  16065=>"001001100",
  16066=>"001001000",
  16067=>"010011001",
  16068=>"000000000",
  16069=>"011101111",
  16070=>"100110010",
  16071=>"011011011",
  16072=>"100000001",
  16073=>"110010010",
  16074=>"000110100",
  16075=>"100100000",
  16076=>"011011100",
  16077=>"111000100",
  16078=>"110011111",
  16079=>"100100111",
  16080=>"101001000",
  16081=>"110100001",
  16082=>"100110100",
  16083=>"100000000",
  16084=>"001000000",
  16085=>"000100100",
  16086=>"111110010",
  16087=>"100000000",
  16088=>"000000000",
  16089=>"110100000",
  16090=>"100111011",
  16091=>"001011111",
  16092=>"100111111",
  16093=>"011011101",
  16094=>"000110100",
  16095=>"000111001",
  16096=>"100100100",
  16097=>"011001001",
  16098=>"100000000",
  16099=>"000100010",
  16100=>"000010100",
  16101=>"000110000",
  16102=>"100100000",
  16103=>"110010101",
  16104=>"010000000",
  16105=>"010010000",
  16106=>"111100000",
  16107=>"011000000",
  16108=>"110100000",
  16109=>"000010000",
  16110=>"010011010",
  16111=>"000000110",
  16112=>"010110111",
  16113=>"011011110",
  16114=>"000111111",
  16115=>"100100000",
  16116=>"100100111",
  16117=>"000111011",
  16118=>"000110011",
  16119=>"000000010",
  16120=>"011001111",
  16121=>"100110000",
  16122=>"011111100",
  16123=>"110011111",
  16124=>"001001100",
  16125=>"000000100",
  16126=>"100110110",
  16127=>"010011111",
  16128=>"111111001",
  16129=>"000111111",
  16130=>"100000100",
  16131=>"110111111",
  16132=>"001011001",
  16133=>"000001000",
  16134=>"000000110",
  16135=>"111111111",
  16136=>"010000000",
  16137=>"000000000",
  16138=>"000000011",
  16139=>"010111111",
  16140=>"110111111",
  16141=>"111111000",
  16142=>"000111111",
  16143=>"000000000",
  16144=>"110000000",
  16145=>"000000000",
  16146=>"111000000",
  16147=>"000100111",
  16148=>"111001000",
  16149=>"111111111",
  16150=>"101001100",
  16151=>"111010010",
  16152=>"000111111",
  16153=>"000000000",
  16154=>"000010000",
  16155=>"000000111",
  16156=>"111101111",
  16157=>"000001100",
  16158=>"011000010",
  16159=>"000111111",
  16160=>"000000000",
  16161=>"011111010",
  16162=>"101000101",
  16163=>"101111111",
  16164=>"101101001",
  16165=>"110110100",
  16166=>"000000001",
  16167=>"111111111",
  16168=>"111110111",
  16169=>"001101111",
  16170=>"111111111",
  16171=>"111100111",
  16172=>"000111111",
  16173=>"001011001",
  16174=>"111100111",
  16175=>"110111111",
  16176=>"000000010",
  16177=>"011011010",
  16178=>"111111111",
  16179=>"111101111",
  16180=>"001000000",
  16181=>"011101111",
  16182=>"111111111",
  16183=>"000000001",
  16184=>"111000000",
  16185=>"011001000",
  16186=>"000000010",
  16187=>"111000110",
  16188=>"100100110",
  16189=>"000111111",
  16190=>"000000111",
  16191=>"000000000",
  16192=>"100000001",
  16193=>"101111010",
  16194=>"000000111",
  16195=>"010000000",
  16196=>"110111111",
  16197=>"000001000",
  16198=>"000000000",
  16199=>"010000011",
  16200=>"111110111",
  16201=>"000000000",
  16202=>"111010000",
  16203=>"000000000",
  16204=>"000000000",
  16205=>"110000001",
  16206=>"000000111",
  16207=>"101111010",
  16208=>"111111110",
  16209=>"111111001",
  16210=>"000000000",
  16211=>"001011010",
  16212=>"000110111",
  16213=>"010110110",
  16214=>"000000000",
  16215=>"000000000",
  16216=>"000000000",
  16217=>"001001000",
  16218=>"000001100",
  16219=>"000001000",
  16220=>"111111000",
  16221=>"001011000",
  16222=>"101101000",
  16223=>"101000010",
  16224=>"000000000",
  16225=>"000100000",
  16226=>"111010010",
  16227=>"000000000",
  16228=>"000100000",
  16229=>"100000000",
  16230=>"001000010",
  16231=>"001000100",
  16232=>"000000000",
  16233=>"001001111",
  16234=>"111100010",
  16235=>"110111110",
  16236=>"111111101",
  16237=>"000000100",
  16238=>"110000000",
  16239=>"000011101",
  16240=>"100100100",
  16241=>"111000000",
  16242=>"111111110",
  16243=>"100000101",
  16244=>"111111000",
  16245=>"000000000",
  16246=>"001111111",
  16247=>"101111111",
  16248=>"000000000",
  16249=>"001111111",
  16250=>"000000000",
  16251=>"111111000",
  16252=>"100100110",
  16253=>"110110000",
  16254=>"001000001",
  16255=>"000000000",
  16256=>"110101000",
  16257=>"111111000",
  16258=>"000000001",
  16259=>"010001001",
  16260=>"111111111",
  16261=>"001000011",
  16262=>"110001011",
  16263=>"001001001",
  16264=>"011011111",
  16265=>"001000000",
  16266=>"100000000",
  16267=>"111010000",
  16268=>"000000000",
  16269=>"000000001",
  16270=>"000111101",
  16271=>"000100110",
  16272=>"011011011",
  16273=>"010111111",
  16274=>"111111000",
  16275=>"110111111",
  16276=>"000001111",
  16277=>"111110010",
  16278=>"111011000",
  16279=>"000000000",
  16280=>"000001001",
  16281=>"000110111",
  16282=>"110000000",
  16283=>"111000000",
  16284=>"111100010",
  16285=>"000110111",
  16286=>"111110000",
  16287=>"101000000",
  16288=>"011011100",
  16289=>"001111010",
  16290=>"111111111",
  16291=>"010000010",
  16292=>"111111111",
  16293=>"000000000",
  16294=>"111100101",
  16295=>"111111101",
  16296=>"000000111",
  16297=>"000111111",
  16298=>"111000100",
  16299=>"000111111",
  16300=>"001000011",
  16301=>"000010111",
  16302=>"110111100",
  16303=>"001101111",
  16304=>"000000000",
  16305=>"001000100",
  16306=>"000000000",
  16307=>"010100100",
  16308=>"000011011",
  16309=>"111111111",
  16310=>"001000100",
  16311=>"111101111",
  16312=>"011001001",
  16313=>"000100111",
  16314=>"000110101",
  16315=>"000110010",
  16316=>"000100000",
  16317=>"111000000",
  16318=>"000000000",
  16319=>"011011111",
  16320=>"000110000",
  16321=>"000000001",
  16322=>"111101011",
  16323=>"111011111",
  16324=>"000000000",
  16325=>"010101111",
  16326=>"000000011",
  16327=>"111110100",
  16328=>"111000111",
  16329=>"000000001",
  16330=>"010110111",
  16331=>"000000000",
  16332=>"000000000",
  16333=>"001001011",
  16334=>"000000011",
  16335=>"111101011",
  16336=>"000000000",
  16337=>"001000000",
  16338=>"001000001",
  16339=>"000000001",
  16340=>"100110100",
  16341=>"101011111",
  16342=>"110101000",
  16343=>"000000011",
  16344=>"111111100",
  16345=>"001100111",
  16346=>"110000001",
  16347=>"111000100",
  16348=>"000000011",
  16349=>"100110111",
  16350=>"000000000",
  16351=>"111010111",
  16352=>"000011001",
  16353=>"111001010",
  16354=>"101111111",
  16355=>"000100100",
  16356=>"111000000",
  16357=>"001111111",
  16358=>"011000000",
  16359=>"110110010",
  16360=>"111000001",
  16361=>"011111101",
  16362=>"000000000",
  16363=>"001001111",
  16364=>"111111111",
  16365=>"111111101",
  16366=>"000000000",
  16367=>"111001000",
  16368=>"000000000",
  16369=>"111111111",
  16370=>"111001001",
  16371=>"000111011",
  16372=>"110110110",
  16373=>"111000001",
  16374=>"101001001",
  16375=>"000001000",
  16376=>"110110010",
  16377=>"111111111",
  16378=>"011111110",
  16379=>"001000111",
  16380=>"000000000",
  16381=>"111111011",
  16382=>"110110101",
  16383=>"111101111",
  16384=>"000000000",
  16385=>"000000001",
  16386=>"010000001",
  16387=>"110000010",
  16388=>"011011010",
  16389=>"100000011",
  16390=>"111010110",
  16391=>"000111010",
  16392=>"110011000",
  16393=>"001000000",
  16394=>"000011110",
  16395=>"101000000",
  16396=>"111000000",
  16397=>"111101101",
  16398=>"100010110",
  16399=>"001000001",
  16400=>"000000110",
  16401=>"000110001",
  16402=>"101000000",
  16403=>"111000001",
  16404=>"111001111",
  16405=>"100000000",
  16406=>"101111000",
  16407=>"111010001",
  16408=>"000000001",
  16409=>"111111111",
  16410=>"111100101",
  16411=>"000110010",
  16412=>"000001101",
  16413=>"101000000",
  16414=>"110100100",
  16415=>"111000000",
  16416=>"110111100",
  16417=>"111111110",
  16418=>"000000001",
  16419=>"100110000",
  16420=>"111111111",
  16421=>"100001111",
  16422=>"000000111",
  16423=>"111110001",
  16424=>"000111110",
  16425=>"000110110",
  16426=>"111000001",
  16427=>"000000111",
  16428=>"011111011",
  16429=>"111000000",
  16430=>"100101011",
  16431=>"100111111",
  16432=>"110110101",
  16433=>"001111111",
  16434=>"110111101",
  16435=>"010110110",
  16436=>"110000111",
  16437=>"010110011",
  16438=>"001010000",
  16439=>"100000000",
  16440=>"010111011",
  16441=>"001000101",
  16442=>"011001001",
  16443=>"000010101",
  16444=>"010011100",
  16445=>"111011000",
  16446=>"111000000",
  16447=>"100001000",
  16448=>"010110000",
  16449=>"110000101",
  16450=>"101010010",
  16451=>"011010011",
  16452=>"100000101",
  16453=>"001000000",
  16454=>"001111010",
  16455=>"110000000",
  16456=>"101001101",
  16457=>"110010000",
  16458=>"001001000",
  16459=>"000000110",
  16460=>"111110110",
  16461=>"010011111",
  16462=>"000100110",
  16463=>"000001110",
  16464=>"000000110",
  16465=>"111001000",
  16466=>"011000010",
  16467=>"011011100",
  16468=>"101100110",
  16469=>"111100000",
  16470=>"000111111",
  16471=>"111101111",
  16472=>"000000100",
  16473=>"011000010",
  16474=>"111001001",
  16475=>"111011110",
  16476=>"100001001",
  16477=>"110001011",
  16478=>"001111111",
  16479=>"111100001",
  16480=>"001001111",
  16481=>"000100000",
  16482=>"101111111",
  16483=>"101000100",
  16484=>"000110100",
  16485=>"011100100",
  16486=>"101000010",
  16487=>"010101111",
  16488=>"000011111",
  16489=>"110000111",
  16490=>"011111000",
  16491=>"000000111",
  16492=>"110100111",
  16493=>"000110110",
  16494=>"111000000",
  16495=>"101111111",
  16496=>"100111101",
  16497=>"110110011",
  16498=>"001100000",
  16499=>"000001001",
  16500=>"000110000",
  16501=>"100000111",
  16502=>"000000010",
  16503=>"100001110",
  16504=>"111000110",
  16505=>"010110001",
  16506=>"111111001",
  16507=>"000001000",
  16508=>"100110100",
  16509=>"100100101",
  16510=>"110111011",
  16511=>"001001110",
  16512=>"011010010",
  16513=>"111000001",
  16514=>"101011100",
  16515=>"111101000",
  16516=>"110000100",
  16517=>"001111111",
  16518=>"110000100",
  16519=>"001100001",
  16520=>"001101011",
  16521=>"000110010",
  16522=>"000001001",
  16523=>"000000000",
  16524=>"000000100",
  16525=>"001001111",
  16526=>"110111000",
  16527=>"100000100",
  16528=>"101111111",
  16529=>"110000111",
  16530=>"010010101",
  16531=>"000001111",
  16532=>"000111110",
  16533=>"110110000",
  16534=>"000111111",
  16535=>"110000000",
  16536=>"001000110",
  16537=>"110001000",
  16538=>"010000000",
  16539=>"000010010",
  16540=>"101000010",
  16541=>"001010010",
  16542=>"110100000",
  16543=>"101001000",
  16544=>"101001100",
  16545=>"111110111",
  16546=>"001001111",
  16547=>"110000001",
  16548=>"110111111",
  16549=>"000011111",
  16550=>"101001001",
  16551=>"101000000",
  16552=>"001110111",
  16553=>"000000111",
  16554=>"111111001",
  16555=>"001110001",
  16556=>"111101101",
  16557=>"001000000",
  16558=>"110011011",
  16559=>"000000010",
  16560=>"111000000",
  16561=>"000001010",
  16562=>"111110000",
  16563=>"100001101",
  16564=>"111101101",
  16565=>"000001001",
  16566=>"000011100",
  16567=>"110010000",
  16568=>"011000101",
  16569=>"100010110",
  16570=>"011001110",
  16571=>"111011001",
  16572=>"011101010",
  16573=>"111111011",
  16574=>"001000001",
  16575=>"110110111",
  16576=>"101001000",
  16577=>"000010000",
  16578=>"010110000",
  16579=>"001011111",
  16580=>"000010111",
  16581=>"111110101",
  16582=>"111110011",
  16583=>"010111111",
  16584=>"101101010",
  16585=>"000010100",
  16586=>"001011000",
  16587=>"001110111",
  16588=>"000001110",
  16589=>"011110110",
  16590=>"111110000",
  16591=>"010010111",
  16592=>"000011000",
  16593=>"000111111",
  16594=>"000011010",
  16595=>"101001100",
  16596=>"100110010",
  16597=>"111000100",
  16598=>"101001101",
  16599=>"000000001",
  16600=>"101001001",
  16601=>"000000000",
  16602=>"011000000",
  16603=>"001000010",
  16604=>"011110000",
  16605=>"000000111",
  16606=>"000111101",
  16607=>"000000110",
  16608=>"001000110",
  16609=>"111111010",
  16610=>"110001001",
  16611=>"000111111",
  16612=>"001000000",
  16613=>"110110110",
  16614=>"000111110",
  16615=>"101101101",
  16616=>"111110000",
  16617=>"111000000",
  16618=>"000100100",
  16619=>"111100000",
  16620=>"110000000",
  16621=>"010001001",
  16622=>"110000100",
  16623=>"010111101",
  16624=>"000001000",
  16625=>"111011101",
  16626=>"100001000",
  16627=>"000011000",
  16628=>"100001011",
  16629=>"000000010",
  16630=>"000100111",
  16631=>"010101001",
  16632=>"101000100",
  16633=>"111101111",
  16634=>"011111101",
  16635=>"000111110",
  16636=>"111111111",
  16637=>"000010000",
  16638=>"110100100",
  16639=>"000111111",
  16640=>"100100100",
  16641=>"000000000",
  16642=>"010010010",
  16643=>"000000011",
  16644=>"111111111",
  16645=>"000001011",
  16646=>"001111011",
  16647=>"000101000",
  16648=>"001111111",
  16649=>"000100001",
  16650=>"110110100",
  16651=>"101001000",
  16652=>"101101101",
  16653=>"101111010",
  16654=>"110000100",
  16655=>"000010001",
  16656=>"100000101",
  16657=>"001011010",
  16658=>"010010000",
  16659=>"000110111",
  16660=>"111111111",
  16661=>"001111111",
  16662=>"100100100",
  16663=>"000101001",
  16664=>"110010000",
  16665=>"111111010",
  16666=>"000000100",
  16667=>"110110011",
  16668=>"110001110",
  16669=>"000000010",
  16670=>"001101111",
  16671=>"000010011",
  16672=>"111111111",
  16673=>"111111010",
  16674=>"000000101",
  16675=>"101001101",
  16676=>"010111000",
  16677=>"001001111",
  16678=>"010011111",
  16679=>"111111011",
  16680=>"111101000",
  16681=>"001111111",
  16682=>"100000100",
  16683=>"000000001",
  16684=>"000100100",
  16685=>"111101100",
  16686=>"000101111",
  16687=>"000100101",
  16688=>"101001000",
  16689=>"111110010",
  16690=>"110000000",
  16691=>"101000000",
  16692=>"001001111",
  16693=>"000101100",
  16694=>"000100100",
  16695=>"101101000",
  16696=>"000000000",
  16697=>"000000000",
  16698=>"000000000",
  16699=>"111111111",
  16700=>"001001011",
  16701=>"011011001",
  16702=>"100000000",
  16703=>"100101001",
  16704=>"111001001",
  16705=>"001101101",
  16706=>"101100000",
  16707=>"100001000",
  16708=>"111110011",
  16709=>"000001111",
  16710=>"001001000",
  16711=>"001101110",
  16712=>"011011001",
  16713=>"101101001",
  16714=>"000101101",
  16715=>"011001101",
  16716=>"000000100",
  16717=>"011011000",
  16718=>"111001000",
  16719=>"000000001",
  16720=>"101101111",
  16721=>"110000001",
  16722=>"000011000",
  16723=>"110000000",
  16724=>"010111101",
  16725=>"011101011",
  16726=>"011011010",
  16727=>"101000100",
  16728=>"010000100",
  16729=>"111110010",
  16730=>"011011011",
  16731=>"101110111",
  16732=>"101101100",
  16733=>"110110100",
  16734=>"101111111",
  16735=>"001000100",
  16736=>"010010010",
  16737=>"001101111",
  16738=>"110010101",
  16739=>"110110110",
  16740=>"011011011",
  16741=>"101100110",
  16742=>"001111001",
  16743=>"010010000",
  16744=>"101000001",
  16745=>"000000000",
  16746=>"001000001",
  16747=>"000011010",
  16748=>"111101100",
  16749=>"010000000",
  16750=>"101101100",
  16751=>"010010000",
  16752=>"101001100",
  16753=>"000111100",
  16754=>"100000000",
  16755=>"000000111",
  16756=>"000000101",
  16757=>"000100100",
  16758=>"101000000",
  16759=>"000010111",
  16760=>"100111100",
  16761=>"010100001",
  16762=>"111000000",
  16763=>"011001001",
  16764=>"011001001",
  16765=>"011001000",
  16766=>"101001111",
  16767=>"010010011",
  16768=>"101111000",
  16769=>"010010000",
  16770=>"000000110",
  16771=>"001001111",
  16772=>"101101001",
  16773=>"000111010",
  16774=>"100100110",
  16775=>"110100100",
  16776=>"110111011",
  16777=>"111010010",
  16778=>"000100100",
  16779=>"101111011",
  16780=>"000000000",
  16781=>"010010111",
  16782=>"101100111",
  16783=>"111000011",
  16784=>"111001111",
  16785=>"000010000",
  16786=>"001000001",
  16787=>"101001000",
  16788=>"111000000",
  16789=>"000000100",
  16790=>"111100101",
  16791=>"010100110",
  16792=>"001111111",
  16793=>"110111000",
  16794=>"000000110",
  16795=>"000000110",
  16796=>"100100100",
  16797=>"010110010",
  16798=>"101101000",
  16799=>"010011000",
  16800=>"100110000",
  16801=>"000010000",
  16802=>"100101011",
  16803=>"000000000",
  16804=>"000101101",
  16805=>"011111001",
  16806=>"111101110",
  16807=>"000100111",
  16808=>"101101001",
  16809=>"000000111",
  16810=>"000000000",
  16811=>"111101010",
  16812=>"101111111",
  16813=>"110010000",
  16814=>"011110100",
  16815=>"101011001",
  16816=>"000111111",
  16817=>"011100001",
  16818=>"000010010",
  16819=>"011011011",
  16820=>"000000000",
  16821=>"101101111",
  16822=>"111011011",
  16823=>"101111011",
  16824=>"110100110",
  16825=>"011001000",
  16826=>"100000000",
  16827=>"101111111",
  16828=>"110010011",
  16829=>"111010011",
  16830=>"100100100",
  16831=>"000101101",
  16832=>"001111000",
  16833=>"000100100",
  16834=>"111110010",
  16835=>"110100111",
  16836=>"111101000",
  16837=>"011011000",
  16838=>"110101000",
  16839=>"010100100",
  16840=>"111000010",
  16841=>"000010110",
  16842=>"000000111",
  16843=>"000000100",
  16844=>"100111111",
  16845=>"110100100",
  16846=>"011111111",
  16847=>"110101000",
  16848=>"111110000",
  16849=>"010011010",
  16850=>"101000001",
  16851=>"100001000",
  16852=>"111111111",
  16853=>"001111111",
  16854=>"110111001",
  16855=>"101000110",
  16856=>"001111101",
  16857=>"010000000",
  16858=>"010001000",
  16859=>"011000000",
  16860=>"000111110",
  16861=>"000100110",
  16862=>"100101111",
  16863=>"111111100",
  16864=>"101101101",
  16865=>"110000000",
  16866=>"101111111",
  16867=>"111000011",
  16868=>"000000000",
  16869=>"111111111",
  16870=>"101000000",
  16871=>"101111010",
  16872=>"000000000",
  16873=>"111111101",
  16874=>"101101001",
  16875=>"001100111",
  16876=>"100101101",
  16877=>"110111011",
  16878=>"111011011",
  16879=>"001111101",
  16880=>"000000001",
  16881=>"110110110",
  16882=>"101101111",
  16883=>"000000100",
  16884=>"001101101",
  16885=>"010010110",
  16886=>"011010111",
  16887=>"000000000",
  16888=>"111001001",
  16889=>"001000000",
  16890=>"010010011",
  16891=>"111000001",
  16892=>"000111111",
  16893=>"100100111",
  16894=>"111110111",
  16895=>"100110000",
  16896=>"011100000",
  16897=>"111111000",
  16898=>"111000101",
  16899=>"101111110",
  16900=>"001111011",
  16901=>"110111110",
  16902=>"011000000",
  16903=>"000000000",
  16904=>"000010010",
  16905=>"010010000",
  16906=>"110000000",
  16907=>"100000001",
  16908=>"101111011",
  16909=>"111111000",
  16910=>"101011100",
  16911=>"000000000",
  16912=>"001111011",
  16913=>"111000000",
  16914=>"001001111",
  16915=>"000010001",
  16916=>"000000010",
  16917=>"110110000",
  16918=>"001001101",
  16919=>"001000110",
  16920=>"101101000",
  16921=>"000000000",
  16922=>"001011010",
  16923=>"111110101",
  16924=>"101111111",
  16925=>"010111111",
  16926=>"111111011",
  16927=>"111000011",
  16928=>"001000000",
  16929=>"101111111",
  16930=>"001000101",
  16931=>"000100111",
  16932=>"001000010",
  16933=>"111010000",
  16934=>"000000111",
  16935=>"000000110",
  16936=>"101111000",
  16937=>"000101100",
  16938=>"011000010",
  16939=>"001101111",
  16940=>"000100111",
  16941=>"100111111",
  16942=>"100111111",
  16943=>"000110110",
  16944=>"001111100",
  16945=>"000011011",
  16946=>"010010010",
  16947=>"010110000",
  16948=>"000000101",
  16949=>"000000100",
  16950=>"111111100",
  16951=>"000001111",
  16952=>"111100000",
  16953=>"001000111",
  16954=>"111000100",
  16955=>"000000100",
  16956=>"100111001",
  16957=>"111111111",
  16958=>"101000101",
  16959=>"001000010",
  16960=>"111001000",
  16961=>"110010000",
  16962=>"111111000",
  16963=>"010001000",
  16964=>"000010000",
  16965=>"000000010",
  16966=>"000010010",
  16967=>"001111101",
  16968=>"000011011",
  16969=>"111111100",
  16970=>"101101101",
  16971=>"001001111",
  16972=>"111010101",
  16973=>"001100000",
  16974=>"110111110",
  16975=>"100111111",
  16976=>"110010000",
  16977=>"111111111",
  16978=>"000100111",
  16979=>"001000001",
  16980=>"101001101",
  16981=>"000010110",
  16982=>"111001000",
  16983=>"111111000",
  16984=>"100000000",
  16985=>"110000001",
  16986=>"000001111",
  16987=>"100000011",
  16988=>"011010000",
  16989=>"000001011",
  16990=>"011111000",
  16991=>"110001000",
  16992=>"000000000",
  16993=>"111110000",
  16994=>"000000000",
  16995=>"000101111",
  16996=>"101101000",
  16997=>"111101001",
  16998=>"011110000",
  16999=>"000110010",
  17000=>"100101001",
  17001=>"010000100",
  17002=>"011111111",
  17003=>"000010000",
  17004=>"111101101",
  17005=>"011011001",
  17006=>"000110011",
  17007=>"111100111",
  17008=>"110110010",
  17009=>"111000000",
  17010=>"111111001",
  17011=>"000000010",
  17012=>"001111011",
  17013=>"000100100",
  17014=>"100110101",
  17015=>"101100001",
  17016=>"110000101",
  17017=>"000000000",
  17018=>"111111111",
  17019=>"111111000",
  17020=>"110111011",
  17021=>"100000000",
  17022=>"100110111",
  17023=>"010010000",
  17024=>"010101111",
  17025=>"111010000",
  17026=>"001010101",
  17027=>"001111111",
  17028=>"000000011",
  17029=>"000000101",
  17030=>"011010011",
  17031=>"000000001",
  17032=>"001011010",
  17033=>"101101101",
  17034=>"000000000",
  17035=>"000111101",
  17036=>"111011000",
  17037=>"101000111",
  17038=>"111010000",
  17039=>"000000101",
  17040=>"000100110",
  17041=>"111000000",
  17042=>"011110000",
  17043=>"000000001",
  17044=>"000010110",
  17045=>"111111001",
  17046=>"001000101",
  17047=>"001001011",
  17048=>"000101000",
  17049=>"000000111",
  17050=>"111010000",
  17051=>"000100100",
  17052=>"000011000",
  17053=>"000001111",
  17054=>"000111111",
  17055=>"000000111",
  17056=>"110110011",
  17057=>"000000111",
  17058=>"011111000",
  17059=>"100101111",
  17060=>"111111111",
  17061=>"000001110",
  17062=>"000001111",
  17063=>"011111000",
  17064=>"111011111",
  17065=>"111111000",
  17066=>"111111000",
  17067=>"100100100",
  17068=>"111001111",
  17069=>"010010000",
  17070=>"011011100",
  17071=>"000101111",
  17072=>"000000001",
  17073=>"001100110",
  17074=>"000101000",
  17075=>"001100010",
  17076=>"110011111",
  17077=>"011110100",
  17078=>"101110110",
  17079=>"001000000",
  17080=>"100111100",
  17081=>"000110010",
  17082=>"011010100",
  17083=>"111111110",
  17084=>"000000001",
  17085=>"111111000",
  17086=>"111011100",
  17087=>"110000000",
  17088=>"010011111",
  17089=>"000000111",
  17090=>"110110011",
  17091=>"011011011",
  17092=>"000000001",
  17093=>"001010101",
  17094=>"010000000",
  17095=>"110101000",
  17096=>"010000000",
  17097=>"000000100",
  17098=>"000001000",
  17099=>"111111010",
  17100=>"100000001",
  17101=>"101111110",
  17102=>"000001111",
  17103=>"001111111",
  17104=>"000001111",
  17105=>"100110011",
  17106=>"110010011",
  17107=>"001001011",
  17108=>"001101111",
  17109=>"100001011",
  17110=>"111110000",
  17111=>"001000111",
  17112=>"000000011",
  17113=>"111111010",
  17114=>"111100100",
  17115=>"100000100",
  17116=>"001100011",
  17117=>"001111111",
  17118=>"110001110",
  17119=>"101001011",
  17120=>"111111000",
  17121=>"111111001",
  17122=>"000000111",
  17123=>"101110100",
  17124=>"101000000",
  17125=>"110111111",
  17126=>"000000010",
  17127=>"001110011",
  17128=>"100111111",
  17129=>"100100101",
  17130=>"011010000",
  17131=>"000000000",
  17132=>"111110000",
  17133=>"011100111",
  17134=>"010000000",
  17135=>"000101111",
  17136=>"100000101",
  17137=>"100110111",
  17138=>"011101011",
  17139=>"001010010",
  17140=>"010001001",
  17141=>"010000111",
  17142=>"000000000",
  17143=>"000000110",
  17144=>"000011010",
  17145=>"001110000",
  17146=>"000010010",
  17147=>"101110111",
  17148=>"000010000",
  17149=>"000000111",
  17150=>"000000000",
  17151=>"000101111",
  17152=>"000011001",
  17153=>"111000000",
  17154=>"001001000",
  17155=>"001111010",
  17156=>"010110111",
  17157=>"111000101",
  17158=>"000111111",
  17159=>"000110110",
  17160=>"111001000",
  17161=>"000001000",
  17162=>"100000110",
  17163=>"111111110",
  17164=>"111001000",
  17165=>"101000000",
  17166=>"100100000",
  17167=>"000101001",
  17168=>"000101101",
  17169=>"000001100",
  17170=>"000001110",
  17171=>"111110111",
  17172=>"110111111",
  17173=>"111001110",
  17174=>"001110000",
  17175=>"101101111",
  17176=>"101101100",
  17177=>"000111110",
  17178=>"111000000",
  17179=>"000001111",
  17180=>"100111111",
  17181=>"101010111",
  17182=>"111111000",
  17183=>"000000001",
  17184=>"000111110",
  17185=>"110000000",
  17186=>"111110001",
  17187=>"000000001",
  17188=>"001111111",
  17189=>"011110100",
  17190=>"001000111",
  17191=>"000100000",
  17192=>"110110100",
  17193=>"000100110",
  17194=>"000011110",
  17195=>"111001001",
  17196=>"000110101",
  17197=>"111111001",
  17198=>"100010011",
  17199=>"000010111",
  17200=>"111111000",
  17201=>"100110100",
  17202=>"000111000",
  17203=>"111110111",
  17204=>"000000111",
  17205=>"011011010",
  17206=>"000100000",
  17207=>"000000010",
  17208=>"111111000",
  17209=>"000000010",
  17210=>"010000101",
  17211=>"001001000",
  17212=>"100110011",
  17213=>"111010110",
  17214=>"000000101",
  17215=>"010000001",
  17216=>"111111000",
  17217=>"111100000",
  17218=>"111111111",
  17219=>"100011110",
  17220=>"111000000",
  17221=>"000001101",
  17222=>"001111110",
  17223=>"111000001",
  17224=>"000000000",
  17225=>"000110111",
  17226=>"000111111",
  17227=>"001001010",
  17228=>"000111111",
  17229=>"000110101",
  17230=>"001011111",
  17231=>"100010111",
  17232=>"111001001",
  17233=>"111111000",
  17234=>"000000101",
  17235=>"011011001",
  17236=>"111101001",
  17237=>"010000110",
  17238=>"000111100",
  17239=>"000111101",
  17240=>"111001000",
  17241=>"000100111",
  17242=>"000001101",
  17243=>"111110001",
  17244=>"000110000",
  17245=>"000011001",
  17246=>"111111000",
  17247=>"111110111",
  17248=>"000000000",
  17249=>"001000010",
  17250=>"111001000",
  17251=>"001101100",
  17252=>"000000111",
  17253=>"000010011",
  17254=>"000110110",
  17255=>"000010110",
  17256=>"001011011",
  17257=>"001101111",
  17258=>"000000111",
  17259=>"000100110",
  17260=>"000000001",
  17261=>"001000101",
  17262=>"000000111",
  17263=>"000001101",
  17264=>"011110111",
  17265=>"000010111",
  17266=>"000011001",
  17267=>"001111001",
  17268=>"111110011",
  17269=>"011001100",
  17270=>"111111110",
  17271=>"110000000",
  17272=>"101101110",
  17273=>"000000000",
  17274=>"001000000",
  17275=>"101001000",
  17276=>"001100100",
  17277=>"000100100",
  17278=>"000001011",
  17279=>"101000011",
  17280=>"101000000",
  17281=>"000111000",
  17282=>"000111011",
  17283=>"000001011",
  17284=>"000111101",
  17285=>"111011000",
  17286=>"100011001",
  17287=>"000000001",
  17288=>"000110101",
  17289=>"001000011",
  17290=>"000110111",
  17291=>"000000000",
  17292=>"011000000",
  17293=>"111011111",
  17294=>"000101001",
  17295=>"000001001",
  17296=>"000011101",
  17297=>"000000000",
  17298=>"100000111",
  17299=>"000000000",
  17300=>"000000111",
  17301=>"000001001",
  17302=>"101111000",
  17303=>"010100100",
  17304=>"000111111",
  17305=>"111111110",
  17306=>"111111111",
  17307=>"111000001",
  17308=>"000111011",
  17309=>"000010000",
  17310=>"111111100",
  17311=>"000000111",
  17312=>"001010001",
  17313=>"011010111",
  17314=>"000000000",
  17315=>"100010000",
  17316=>"010000000",
  17317=>"001111000",
  17318=>"001001011",
  17319=>"000110100",
  17320=>"000000000",
  17321=>"111111101",
  17322=>"111101001",
  17323=>"000010100",
  17324=>"100100110",
  17325=>"000100111",
  17326=>"010110110",
  17327=>"111001000",
  17328=>"000110010",
  17329=>"000001000",
  17330=>"111111000",
  17331=>"011011100",
  17332=>"000110111",
  17333=>"110101101",
  17334=>"010000001",
  17335=>"010111101",
  17336=>"000011111",
  17337=>"000000000",
  17338=>"000010100",
  17339=>"110111000",
  17340=>"000000000",
  17341=>"111001001",
  17342=>"100000000",
  17343=>"000000010",
  17344=>"001011110",
  17345=>"000001010",
  17346=>"111110001",
  17347=>"000111111",
  17348=>"000000000",
  17349=>"111111110",
  17350=>"000000000",
  17351=>"111111000",
  17352=>"001101111",
  17353=>"000100100",
  17354=>"000100110",
  17355=>"001110110",
  17356=>"000010010",
  17357=>"000001010",
  17358=>"000000001",
  17359=>"101101101",
  17360=>"101000001",
  17361=>"010011001",
  17362=>"000000000",
  17363=>"001101001",
  17364=>"001111111",
  17365=>"000000000",
  17366=>"000111110",
  17367=>"110110100",
  17368=>"000011000",
  17369=>"000110101",
  17370=>"000000100",
  17371=>"111001101",
  17372=>"110111011",
  17373=>"001101101",
  17374=>"000000000",
  17375=>"000010110",
  17376=>"001000111",
  17377=>"111001000",
  17378=>"111000000",
  17379=>"011010100",
  17380=>"000001111",
  17381=>"111000001",
  17382=>"110000000",
  17383=>"000111110",
  17384=>"000001001",
  17385=>"011111111",
  17386=>"001000011",
  17387=>"000001000",
  17388=>"111101001",
  17389=>"111101101",
  17390=>"010001000",
  17391=>"010001101",
  17392=>"001001001",
  17393=>"000111101",
  17394=>"000000000",
  17395=>"000011111",
  17396=>"000110111",
  17397=>"111001101",
  17398=>"000010110",
  17399=>"010000010",
  17400=>"111011000",
  17401=>"001001011",
  17402=>"010111111",
  17403=>"000110111",
  17404=>"000111110",
  17405=>"111000111",
  17406=>"000111111",
  17407=>"000110110",
  17408=>"110101111",
  17409=>"011011111",
  17410=>"100100111",
  17411=>"100011011",
  17412=>"000000000",
  17413=>"001000010",
  17414=>"001001100",
  17415=>"001001001",
  17416=>"111100111",
  17417=>"100001001",
  17418=>"000100110",
  17419=>"011011011",
  17420=>"111111111",
  17421=>"011010011",
  17422=>"110011001",
  17423=>"011011000",
  17424=>"011010000",
  17425=>"011001011",
  17426=>"100110111",
  17427=>"011000000",
  17428=>"100001100",
  17429=>"100100111",
  17430=>"110101100",
  17431=>"011111110",
  17432=>"000000101",
  17433=>"110000101",
  17434=>"000000111",
  17435=>"101101111",
  17436=>"000100111",
  17437=>"110010001",
  17438=>"111100100",
  17439=>"100010000",
  17440=>"111100111",
  17441=>"011111110",
  17442=>"000011100",
  17443=>"011011011",
  17444=>"000001000",
  17445=>"111000001",
  17446=>"001011000",
  17447=>"011111100",
  17448=>"110110100",
  17449=>"011001000",
  17450=>"010000111",
  17451=>"011011100",
  17452=>"011001001",
  17453=>"100001111",
  17454=>"111001000",
  17455=>"000100111",
  17456=>"110111011",
  17457=>"100001000",
  17458=>"000000000",
  17459=>"100110100",
  17460=>"101111001",
  17461=>"011011100",
  17462=>"110010000",
  17463=>"110110111",
  17464=>"111110110",
  17465=>"100100111",
  17466=>"011110000",
  17467=>"011111000",
  17468=>"011111010",
  17469=>"101011100",
  17470=>"101000001",
  17471=>"001101001",
  17472=>"100100010",
  17473=>"000000000",
  17474=>"100100001",
  17475=>"110000110",
  17476=>"001011000",
  17477=>"100110000",
  17478=>"000100010",
  17479=>"010011000",
  17480=>"000000001",
  17481=>"110111110",
  17482=>"100100111",
  17483=>"100100000",
  17484=>"100100100",
  17485=>"111110100",
  17486=>"110011110",
  17487=>"001111111",
  17488=>"111101100",
  17489=>"000111111",
  17490=>"001000000",
  17491=>"000000001",
  17492=>"111000000",
  17493=>"110111101",
  17494=>"111110011",
  17495=>"001001011",
  17496=>"000110000",
  17497=>"000110010",
  17498=>"010011001",
  17499=>"011011100",
  17500=>"100001100",
  17501=>"001001001",
  17502=>"111101100",
  17503=>"101101001",
  17504=>"011011000",
  17505=>"111100111",
  17506=>"100000011",
  17507=>"110110110",
  17508=>"111101111",
  17509=>"110100000",
  17510=>"000110100",
  17511=>"110111110",
  17512=>"011110001",
  17513=>"000001001",
  17514=>"001000000",
  17515=>"010000000",
  17516=>"000011011",
  17517=>"111101001",
  17518=>"110110011",
  17519=>"001011000",
  17520=>"111111101",
  17521=>"010111111",
  17522=>"000100110",
  17523=>"000001000",
  17524=>"011011000",
  17525=>"100000000",
  17526=>"100001000",
  17527=>"011010000",
  17528=>"000100001",
  17529=>"001101000",
  17530=>"111101000",
  17531=>"011010011",
  17532=>"100001000",
  17533=>"100000000",
  17534=>"100100111",
  17535=>"000000101",
  17536=>"001000100",
  17537=>"100100100",
  17538=>"000001000",
  17539=>"011001011",
  17540=>"011010000",
  17541=>"101100111",
  17542=>"010001010",
  17543=>"000100100",
  17544=>"111111001",
  17545=>"010111011",
  17546=>"110111111",
  17547=>"111101100",
  17548=>"111111100",
  17549=>"000000010",
  17550=>"110100110",
  17551=>"000000001",
  17552=>"000001000",
  17553=>"100111110",
  17554=>"011011001",
  17555=>"011110010",
  17556=>"000011111",
  17557=>"111100110",
  17558=>"000110001",
  17559=>"001001011",
  17560=>"000001000",
  17561=>"011011000",
  17562=>"100100110",
  17563=>"000000111",
  17564=>"110110111",
  17565=>"011000001",
  17566=>"100000111",
  17567=>"000001111",
  17568=>"000100000",
  17569=>"101101111",
  17570=>"100011110",
  17571=>"000000111",
  17572=>"100100101",
  17573=>"110011011",
  17574=>"011011000",
  17575=>"111011110",
  17576=>"111100111",
  17577=>"011011110",
  17578=>"100110111",
  17579=>"111100001",
  17580=>"011111101",
  17581=>"100110001",
  17582=>"101101101",
  17583=>"001001000",
  17584=>"101011111",
  17585=>"000001001",
  17586=>"000011000",
  17587=>"000000100",
  17588=>"000001000",
  17589=>"000100100",
  17590=>"001010010",
  17591=>"111111011",
  17592=>"100000000",
  17593=>"011011100",
  17594=>"111010011",
  17595=>"110110111",
  17596=>"100111111",
  17597=>"101111101",
  17598=>"101111110",
  17599=>"001011011",
  17600=>"110100101",
  17601=>"010110111",
  17602=>"100000000",
  17603=>"110100110",
  17604=>"000011011",
  17605=>"110111100",
  17606=>"000001001",
  17607=>"000000101",
  17608=>"000100100",
  17609=>"001000000",
  17610=>"100110100",
  17611=>"100100111",
  17612=>"110100000",
  17613=>"001001000",
  17614=>"100000000",
  17615=>"001000110",
  17616=>"110100000",
  17617=>"111011011",
  17618=>"000010011",
  17619=>"110110111",
  17620=>"000000000",
  17621=>"001011000",
  17622=>"000011000",
  17623=>"111100101",
  17624=>"111011001",
  17625=>"000100010",
  17626=>"101111110",
  17627=>"000100111",
  17628=>"101001010",
  17629=>"010011011",
  17630=>"011000000",
  17631=>"011110000",
  17632=>"111110111",
  17633=>"100100110",
  17634=>"001000000",
  17635=>"001100100",
  17636=>"110100111",
  17637=>"011011000",
  17638=>"011100000",
  17639=>"000000000",
  17640=>"000010001",
  17641=>"111111110",
  17642=>"100000000",
  17643=>"101111111",
  17644=>"011001100",
  17645=>"000010011",
  17646=>"000100000",
  17647=>"111011001",
  17648=>"011011000",
  17649=>"000110100",
  17650=>"111001100",
  17651=>"111111011",
  17652=>"110111101",
  17653=>"000010111",
  17654=>"000001001",
  17655=>"000001000",
  17656=>"000110000",
  17657=>"010000000",
  17658=>"000110000",
  17659=>"110111000",
  17660=>"100100111",
  17661=>"001001000",
  17662=>"000000000",
  17663=>"100000111",
  17664=>"111111011",
  17665=>"000110100",
  17666=>"001100100",
  17667=>"000100011",
  17668=>"101110001",
  17669=>"001101000",
  17670=>"000111111",
  17671=>"010010111",
  17672=>"000000111",
  17673=>"000100111",
  17674=>"010011100",
  17675=>"111011011",
  17676=>"101111001",
  17677=>"000010000",
  17678=>"000000000",
  17679=>"101111100",
  17680=>"100000100",
  17681=>"001001011",
  17682=>"011000000",
  17683=>"010100011",
  17684=>"101101111",
  17685=>"010000100",
  17686=>"110111001",
  17687=>"111111111",
  17688=>"101101100",
  17689=>"110111111",
  17690=>"001000010",
  17691=>"110110111",
  17692=>"000111110",
  17693=>"111110000",
  17694=>"000000000",
  17695=>"001011000",
  17696=>"011000101",
  17697=>"011011110",
  17698=>"011000000",
  17699=>"000000110",
  17700=>"101111101",
  17701=>"100000000",
  17702=>"000100101",
  17703=>"000011111",
  17704=>"001001111",
  17705=>"010110111",
  17706=>"000001111",
  17707=>"010000000",
  17708=>"000000000",
  17709=>"100110100",
  17710=>"111001001",
  17711=>"110000000",
  17712=>"011001001",
  17713=>"110111001",
  17714=>"111001000",
  17715=>"001000000",
  17716=>"000100011",
  17717=>"101000010",
  17718=>"000000000",
  17719=>"110110011",
  17720=>"011011010",
  17721=>"111110010",
  17722=>"101100110",
  17723=>"000100000",
  17724=>"000011011",
  17725=>"110011111",
  17726=>"001000000",
  17727=>"110111011",
  17728=>"110100100",
  17729=>"011001111",
  17730=>"001010001",
  17731=>"111011011",
  17732=>"111100100",
  17733=>"001000000",
  17734=>"000100011",
  17735=>"001001000",
  17736=>"000000010",
  17737=>"000111111",
  17738=>"011000001",
  17739=>"001100110",
  17740=>"000000000",
  17741=>"111111101",
  17742=>"110111111",
  17743=>"000011100",
  17744=>"011111000",
  17745=>"110100110",
  17746=>"100001010",
  17747=>"111101101",
  17748=>"011000000",
  17749=>"100011111",
  17750=>"111111111",
  17751=>"011111110",
  17752=>"100010111",
  17753=>"000000000",
  17754=>"000100110",
  17755=>"101011110",
  17756=>"001001010",
  17757=>"011000000",
  17758=>"101100111",
  17759=>"000000000",
  17760=>"100011001",
  17761=>"111110110",
  17762=>"001100100",
  17763=>"110010110",
  17764=>"010000001",
  17765=>"000001001",
  17766=>"111111111",
  17767=>"110111110",
  17768=>"100000000",
  17769=>"111001000",
  17770=>"100010011",
  17771=>"101111111",
  17772=>"110001100",
  17773=>"001100110",
  17774=>"110000100",
  17775=>"000110101",
  17776=>"111101101",
  17777=>"110110011",
  17778=>"110110001",
  17779=>"001001011",
  17780=>"001011010",
  17781=>"000000000",
  17782=>"000100111",
  17783=>"000111011",
  17784=>"111001010",
  17785=>"110111011",
  17786=>"010011001",
  17787=>"001000000",
  17788=>"111100111",
  17789=>"000000000",
  17790=>"111001100",
  17791=>"101100110",
  17792=>"011001011",
  17793=>"000000000",
  17794=>"101011011",
  17795=>"100110011",
  17796=>"011001001",
  17797=>"100001101",
  17798=>"001001001",
  17799=>"110100000",
  17800=>"000011111",
  17801=>"000001000",
  17802=>"110000001",
  17803=>"100000000",
  17804=>"110110010",
  17805=>"111001100",
  17806=>"111100110",
  17807=>"000001010",
  17808=>"111100111",
  17809=>"100100110",
  17810=>"000000001",
  17811=>"110110111",
  17812=>"000000001",
  17813=>"011110110",
  17814=>"110111010",
  17815=>"100000000",
  17816=>"100011011",
  17817=>"000000111",
  17818=>"000010100",
  17819=>"011000101",
  17820=>"100110011",
  17821=>"100100000",
  17822=>"111111110",
  17823=>"000100100",
  17824=>"111111000",
  17825=>"011000100",
  17826=>"000000000",
  17827=>"100100000",
  17828=>"110011001",
  17829=>"000001111",
  17830=>"001001100",
  17831=>"110001001",
  17832=>"001001010",
  17833=>"101100100",
  17834=>"011101110",
  17835=>"000000100",
  17836=>"100101100",
  17837=>"111001000",
  17838=>"000000000",
  17839=>"100100110",
  17840=>"000000000",
  17841=>"111111111",
  17842=>"010010000",
  17843=>"111111111",
  17844=>"110000000",
  17845=>"010010000",
  17846=>"100110000",
  17847=>"011111101",
  17848=>"100101000",
  17849=>"100110010",
  17850=>"110101110",
  17851=>"010011011",
  17852=>"101001001",
  17853=>"110110001",
  17854=>"101100011",
  17855=>"000000011",
  17856=>"010000000",
  17857=>"100111000",
  17858=>"110111111",
  17859=>"011111111",
  17860=>"000000000",
  17861=>"010111110",
  17862=>"100000000",
  17863=>"000010010",
  17864=>"000000000",
  17865=>"000000000",
  17866=>"010001110",
  17867=>"100110111",
  17868=>"110110111",
  17869=>"000000000",
  17870=>"001101111",
  17871=>"000000100",
  17872=>"100110010",
  17873=>"011110111",
  17874=>"100000000",
  17875=>"110011011",
  17876=>"011001100",
  17877=>"011010000",
  17878=>"011011110",
  17879=>"000000000",
  17880=>"110011001",
  17881=>"000000101",
  17882=>"001111111",
  17883=>"011100110",
  17884=>"000000000",
  17885=>"000000000",
  17886=>"100111000",
  17887=>"100010011",
  17888=>"000000100",
  17889=>"001000100",
  17890=>"110011001",
  17891=>"111011101",
  17892=>"000000001",
  17893=>"011110011",
  17894=>"100011111",
  17895=>"111011111",
  17896=>"000001011",
  17897=>"000000000",
  17898=>"000100011",
  17899=>"100101110",
  17900=>"100100111",
  17901=>"011000100",
  17902=>"110000000",
  17903=>"001000011",
  17904=>"000001011",
  17905=>"000000000",
  17906=>"111001011",
  17907=>"000011001",
  17908=>"000000000",
  17909=>"001000100",
  17910=>"001100011",
  17911=>"111000000",
  17912=>"010010001",
  17913=>"010000111",
  17914=>"101110101",
  17915=>"001111011",
  17916=>"111011011",
  17917=>"001001001",
  17918=>"000100000",
  17919=>"111011001",
  17920=>"111011000",
  17921=>"100110010",
  17922=>"110110110",
  17923=>"000111001",
  17924=>"110011011",
  17925=>"100000111",
  17926=>"100100000",
  17927=>"100111110",
  17928=>"011001001",
  17929=>"111110001",
  17930=>"101100000",
  17931=>"111000000",
  17932=>"000000000",
  17933=>"000000000",
  17934=>"110111110",
  17935=>"000001011",
  17936=>"111111001",
  17937=>"011000000",
  17938=>"111111101",
  17939=>"100101000",
  17940=>"111111100",
  17941=>"111111111",
  17942=>"111111001",
  17943=>"111111000",
  17944=>"111111111",
  17945=>"001000011",
  17946=>"000100000",
  17947=>"111000000",
  17948=>"001000000",
  17949=>"000000010",
  17950=>"101001110",
  17951=>"010000001",
  17952=>"100000000",
  17953=>"010000000",
  17954=>"010000100",
  17955=>"000001111",
  17956=>"100100000",
  17957=>"101010001",
  17958=>"111111011",
  17959=>"111011101",
  17960=>"111111000",
  17961=>"000000000",
  17962=>"110111111",
  17963=>"110000010",
  17964=>"110100000",
  17965=>"111111001",
  17966=>"000000101",
  17967=>"111011111",
  17968=>"111111111",
  17969=>"011000111",
  17970=>"000000010",
  17971=>"000000111",
  17972=>"111010000",
  17973=>"111011101",
  17974=>"011011000",
  17975=>"000000000",
  17976=>"111010000",
  17977=>"111111000",
  17978=>"000000001",
  17979=>"111000011",
  17980=>"000110000",
  17981=>"001001001",
  17982=>"100111000",
  17983=>"111111101",
  17984=>"110000000",
  17985=>"011000001",
  17986=>"000111100",
  17987=>"111111011",
  17988=>"000011001",
  17989=>"000000111",
  17990=>"000100100",
  17991=>"001000011",
  17992=>"000000000",
  17993=>"011111000",
  17994=>"111100101",
  17995=>"000010111",
  17996=>"001000011",
  17997=>"110000001",
  17998=>"010111001",
  17999=>"000000111",
  18000=>"000101101",
  18001=>"000111001",
  18002=>"010111111",
  18003=>"101000000",
  18004=>"111111011",
  18005=>"110111001",
  18006=>"010110011",
  18007=>"111001001",
  18008=>"110110000",
  18009=>"001001011",
  18010=>"001111110",
  18011=>"011100100",
  18012=>"111111000",
  18013=>"001010000",
  18014=>"110100111",
  18015=>"111111000",
  18016=>"100100000",
  18017=>"111111111",
  18018=>"001100111",
  18019=>"110111001",
  18020=>"010011000",
  18021=>"000100111",
  18022=>"111001111",
  18023=>"000000111",
  18024=>"111111000",
  18025=>"000000000",
  18026=>"110101101",
  18027=>"000000011",
  18028=>"000100000",
  18029=>"000011111",
  18030=>"111010110",
  18031=>"000011000",
  18032=>"100100011",
  18033=>"000110111",
  18034=>"111100000",
  18035=>"000000111",
  18036=>"100001101",
  18037=>"101010011",
  18038=>"110011000",
  18039=>"000110110",
  18040=>"011111010",
  18041=>"000000000",
  18042=>"010001100",
  18043=>"111000000",
  18044=>"111000000",
  18045=>"000000101",
  18046=>"001100000",
  18047=>"111101000",
  18048=>"111011010",
  18049=>"001000000",
  18050=>"111111100",
  18051=>"000000010",
  18052=>"000000000",
  18053=>"111111001",
  18054=>"101100000",
  18055=>"000100000",
  18056=>"000110010",
  18057=>"111111000",
  18058=>"001101111",
  18059=>"000000111",
  18060=>"001111111",
  18061=>"111101001",
  18062=>"111111100",
  18063=>"000010000",
  18064=>"001001110",
  18065=>"111111000",
  18066=>"000010000",
  18067=>"110111000",
  18068=>"111111100",
  18069=>"000101000",
  18070=>"000110110",
  18071=>"010100101",
  18072=>"111100101",
  18073=>"011111010",
  18074=>"111110100",
  18075=>"111101100",
  18076=>"111111111",
  18077=>"111100000",
  18078=>"111110101",
  18079=>"000000110",
  18080=>"111100100",
  18081=>"111111111",
  18082=>"000101110",
  18083=>"110000111",
  18084=>"111000000",
  18085=>"100110000",
  18086=>"001001111",
  18087=>"111111101",
  18088=>"101111100",
  18089=>"111110111",
  18090=>"111000111",
  18091=>"000111111",
  18092=>"000001100",
  18093=>"000000011",
  18094=>"111110000",
  18095=>"000000111",
  18096=>"100000000",
  18097=>"000000000",
  18098=>"000110000",
  18099=>"010100000",
  18100=>"001110000",
  18101=>"111101001",
  18102=>"010010010",
  18103=>"000000111",
  18104=>"010001000",
  18105=>"111111101",
  18106=>"111101111",
  18107=>"100000111",
  18108=>"000000101",
  18109=>"011111111",
  18110=>"110110000",
  18111=>"000000100",
  18112=>"111110000",
  18113=>"000000110",
  18114=>"000011110",
  18115=>"111110111",
  18116=>"000000100",
  18117=>"101011011",
  18118=>"011011110",
  18119=>"101000000",
  18120=>"100000000",
  18121=>"111001011",
  18122=>"000001011",
  18123=>"111000000",
  18124=>"111011111",
  18125=>"110011000",
  18126=>"000010110",
  18127=>"101000000",
  18128=>"111100100",
  18129=>"000000010",
  18130=>"000001010",
  18131=>"010010111",
  18132=>"111000000",
  18133=>"100010011",
  18134=>"111000000",
  18135=>"111011000",
  18136=>"111111000",
  18137=>"011111001",
  18138=>"111001010",
  18139=>"000000111",
  18140=>"001111100",
  18141=>"000101111",
  18142=>"001011111",
  18143=>"101110000",
  18144=>"111111111",
  18145=>"100000111",
  18146=>"110000100",
  18147=>"010110000",
  18148=>"000000010",
  18149=>"111000000",
  18150=>"110011000",
  18151=>"110100110",
  18152=>"000000011",
  18153=>"000000001",
  18154=>"111001000",
  18155=>"000000101",
  18156=>"111111111",
  18157=>"000000011",
  18158=>"000000011",
  18159=>"111000000",
  18160=>"100011000",
  18161=>"011111100",
  18162=>"111101101",
  18163=>"100110000",
  18164=>"001000000",
  18165=>"000111111",
  18166=>"000000111",
  18167=>"111101111",
  18168=>"111101000",
  18169=>"111101111",
  18170=>"000011011",
  18171=>"010001000",
  18172=>"111111000",
  18173=>"101101111",
  18174=>"001000110",
  18175=>"000000000",
  18176=>"000000111",
  18177=>"000011000",
  18178=>"000001001",
  18179=>"110000000",
  18180=>"010011001",
  18181=>"100000000",
  18182=>"111111111",
  18183=>"000011001",
  18184=>"100000000",
  18185=>"111111001",
  18186=>"000111001",
  18187=>"100000000",
  18188=>"111000000",
  18189=>"000111111",
  18190=>"001110100",
  18191=>"000000000",
  18192=>"111101001",
  18193=>"101111000",
  18194=>"111111110",
  18195=>"110010000",
  18196=>"000000000",
  18197=>"111111111",
  18198=>"000011110",
  18199=>"111011111",
  18200=>"111111111",
  18201=>"000000000",
  18202=>"000011000",
  18203=>"111111000",
  18204=>"000000010",
  18205=>"000000000",
  18206=>"111101111",
  18207=>"011000000",
  18208=>"000000000",
  18209=>"000111000",
  18210=>"000100000",
  18211=>"111000100",
  18212=>"111111111",
  18213=>"111001110",
  18214=>"111111111",
  18215=>"111111111",
  18216=>"111111000",
  18217=>"111111001",
  18218=>"000110000",
  18219=>"000011010",
  18220=>"110100110",
  18221=>"111010111",
  18222=>"000011100",
  18223=>"000010000",
  18224=>"111111110",
  18225=>"111011011",
  18226=>"111111100",
  18227=>"000111000",
  18228=>"110010101",
  18229=>"111111110",
  18230=>"001011101",
  18231=>"000001000",
  18232=>"010000011",
  18233=>"000110000",
  18234=>"110100111",
  18235=>"100110000",
  18236=>"100111011",
  18237=>"001111111",
  18238=>"000100000",
  18239=>"011011011",
  18240=>"000010001",
  18241=>"001111111",
  18242=>"000000000",
  18243=>"100000100",
  18244=>"110110000",
  18245=>"111101110",
  18246=>"111111111",
  18247=>"111111101",
  18248=>"000000010",
  18249=>"001000000",
  18250=>"100101110",
  18251=>"000111111",
  18252=>"111011000",
  18253=>"110000000",
  18254=>"001000010",
  18255=>"111000101",
  18256=>"111001000",
  18257=>"010111010",
  18258=>"000010000",
  18259=>"011111001",
  18260=>"000000000",
  18261=>"110110111",
  18262=>"110010010",
  18263=>"001001000",
  18264=>"001000101",
  18265=>"000010011",
  18266=>"110110001",
  18267=>"111111111",
  18268=>"000000000",
  18269=>"000111110",
  18270=>"010110000",
  18271=>"011100000",
  18272=>"101101000",
  18273=>"000110010",
  18274=>"000001000",
  18275=>"101111111",
  18276=>"111111111",
  18277=>"000000000",
  18278=>"000000000",
  18279=>"000000010",
  18280=>"010110100",
  18281=>"000100111",
  18282=>"000000001",
  18283=>"010111111",
  18284=>"000000000",
  18285=>"111010000",
  18286=>"111111011",
  18287=>"111111111",
  18288=>"011011110",
  18289=>"000000100",
  18290=>"000110110",
  18291=>"000000000",
  18292=>"000010000",
  18293=>"110000111",
  18294=>"100110100",
  18295=>"000000011",
  18296=>"100101000",
  18297=>"110111110",
  18298=>"111111111",
  18299=>"111000001",
  18300=>"001011001",
  18301=>"001011011",
  18302=>"010111111",
  18303=>"000000010",
  18304=>"000000000",
  18305=>"000111111",
  18306=>"010011011",
  18307=>"011101111",
  18308=>"111011001",
  18309=>"111101111",
  18310=>"110100110",
  18311=>"110101000",
  18312=>"111111111",
  18313=>"000101000",
  18314=>"111110111",
  18315=>"111101001",
  18316=>"000010000",
  18317=>"000011110",
  18318=>"000000000",
  18319=>"000000000",
  18320=>"110111011",
  18321=>"010111111",
  18322=>"000001001",
  18323=>"111101101",
  18324=>"000001001",
  18325=>"100101100",
  18326=>"000000000",
  18327=>"100111110",
  18328=>"111000000",
  18329=>"000001001",
  18330=>"111111111",
  18331=>"101011000",
  18332=>"000000000",
  18333=>"111000010",
  18334=>"001111110",
  18335=>"011010000",
  18336=>"111111111",
  18337=>"001011010",
  18338=>"011111110",
  18339=>"000001111",
  18340=>"000111111",
  18341=>"110100100",
  18342=>"111101010",
  18343=>"111000000",
  18344=>"101000111",
  18345=>"000101010",
  18346=>"010110000",
  18347=>"011011000",
  18348=>"111001111",
  18349=>"000001111",
  18350=>"100011000",
  18351=>"000111011",
  18352=>"010000001",
  18353=>"001100000",
  18354=>"000000000",
  18355=>"000011001",
  18356=>"011000111",
  18357=>"111111110",
  18358=>"000001001",
  18359=>"010000000",
  18360=>"001110000",
  18361=>"100111101",
  18362=>"111010001",
  18363=>"010001110",
  18364=>"110110111",
  18365=>"011111010",
  18366=>"000000000",
  18367=>"000111011",
  18368=>"000111111",
  18369=>"000000000",
  18370=>"111111101",
  18371=>"011011011",
  18372=>"000100100",
  18373=>"000110110",
  18374=>"000010000",
  18375=>"000101000",
  18376=>"111110010",
  18377=>"101101111",
  18378=>"101100101",
  18379=>"111111111",
  18380=>"010010010",
  18381=>"000101100",
  18382=>"110111010",
  18383=>"111111111",
  18384=>"010010010",
  18385=>"111111111",
  18386=>"100010000",
  18387=>"000000000",
  18388=>"000000000",
  18389=>"000000000",
  18390=>"111111000",
  18391=>"010111000",
  18392=>"000000010",
  18393=>"010010000",
  18394=>"111111111",
  18395=>"010111000",
  18396=>"110111110",
  18397=>"000001101",
  18398=>"000000100",
  18399=>"000000011",
  18400=>"000000000",
  18401=>"010010001",
  18402=>"010000111",
  18403=>"000000011",
  18404=>"000000000",
  18405=>"000010010",
  18406=>"011111111",
  18407=>"000111101",
  18408=>"111000001",
  18409=>"110110001",
  18410=>"011111000",
  18411=>"001001000",
  18412=>"001000000",
  18413=>"101101100",
  18414=>"000011000",
  18415=>"000000000",
  18416=>"000000000",
  18417=>"011011111",
  18418=>"111101111",
  18419=>"110110000",
  18420=>"010000111",
  18421=>"110010010",
  18422=>"111000111",
  18423=>"000010000",
  18424=>"000010011",
  18425=>"111101010",
  18426=>"111001000",
  18427=>"000010000",
  18428=>"111111111",
  18429=>"000011000",
  18430=>"111111011",
  18431=>"101111000",
  18432=>"101111001",
  18433=>"111011011",
  18434=>"111000001",
  18435=>"000000110",
  18436=>"010011111",
  18437=>"010100001",
  18438=>"011001001",
  18439=>"110111010",
  18440=>"111011011",
  18441=>"001111001",
  18442=>"000000001",
  18443=>"011001001",
  18444=>"000100100",
  18445=>"100100000",
  18446=>"001101110",
  18447=>"000010000",
  18448=>"001111001",
  18449=>"000000110",
  18450=>"010000000",
  18451=>"001000100",
  18452=>"111100100",
  18453=>"011000000",
  18454=>"001001011",
  18455=>"100001111",
  18456=>"011001011",
  18457=>"111011001",
  18458=>"100110001",
  18459=>"000000110",
  18460=>"001011111",
  18461=>"000000110",
  18462=>"110100010",
  18463=>"110100000",
  18464=>"001001001",
  18465=>"101110001",
  18466=>"000111111",
  18467=>"010000011",
  18468=>"111111101",
  18469=>"011010111",
  18470=>"001011001",
  18471=>"000110110",
  18472=>"100110000",
  18473=>"100100000",
  18474=>"001001001",
  18475=>"110011011",
  18476=>"001111111",
  18477=>"110010001",
  18478=>"001101101",
  18479=>"110111110",
  18480=>"000101110",
  18481=>"011111111",
  18482=>"111101101",
  18483=>"110110101",
  18484=>"000100111",
  18485=>"001000101",
  18486=>"001010000",
  18487=>"011001011",
  18488=>"100000000",
  18489=>"011001011",
  18490=>"000101110",
  18491=>"001011100",
  18492=>"110111111",
  18493=>"100011011",
  18494=>"011001001",
  18495=>"111101111",
  18496=>"001000000",
  18497=>"001111011",
  18498=>"001000001",
  18499=>"001011011",
  18500=>"100000110",
  18501=>"011000001",
  18502=>"100001011",
  18503=>"110010000",
  18504=>"010111111",
  18505=>"111110110",
  18506=>"011001011",
  18507=>"011001011",
  18508=>"011001001",
  18509=>"001111100",
  18510=>"010000000",
  18511=>"110010111",
  18512=>"001110100",
  18513=>"110101000",
  18514=>"011001000",
  18515=>"110011001",
  18516=>"010000110",
  18517=>"111010111",
  18518=>"111111011",
  18519=>"011111111",
  18520=>"110001101",
  18521=>"001101010",
  18522=>"100001011",
  18523=>"000000110",
  18524=>"001000010",
  18525=>"100100000",
  18526=>"000110110",
  18527=>"011001011",
  18528=>"011001111",
  18529=>"100010011",
  18530=>"100000001",
  18531=>"110101000",
  18532=>"111100100",
  18533=>"011001001",
  18534=>"000110110",
  18535=>"011011010",
  18536=>"011000110",
  18537=>"110100001",
  18538=>"110110100",
  18539=>"110111001",
  18540=>"001011001",
  18541=>"111100100",
  18542=>"001001001",
  18543=>"001110110",
  18544=>"100000000",
  18545=>"010001100",
  18546=>"100111011",
  18547=>"001001010",
  18548=>"000101110",
  18549=>"011001011",
  18550=>"100100100",
  18551=>"100110100",
  18552=>"110010000",
  18553=>"110110010",
  18554=>"100000001",
  18555=>"110111000",
  18556=>"000100011",
  18557=>"110000000",
  18558=>"101001011",
  18559=>"100000000",
  18560=>"001011111",
  18561=>"010000000",
  18562=>"111001111",
  18563=>"100111111",
  18564=>"100110000",
  18565=>"011000110",
  18566=>"001011110",
  18567=>"011001001",
  18568=>"110111111",
  18569=>"010000110",
  18570=>"111011011",
  18571=>"011011001",
  18572=>"011000000",
  18573=>"001000001",
  18574=>"011001000",
  18575=>"010001001",
  18576=>"001001001",
  18577=>"001111010",
  18578=>"001001000",
  18579=>"111011001",
  18580=>"001001001",
  18581=>"111100001",
  18582=>"011011011",
  18583=>"111111101",
  18584=>"011100001",
  18585=>"010100111",
  18586=>"101001000",
  18587=>"000000000",
  18588=>"111010000",
  18589=>"111011101",
  18590=>"000000111",
  18591=>"011001011",
  18592=>"001111111",
  18593=>"011111000",
  18594=>"000001001",
  18595=>"000001001",
  18596=>"100100110",
  18597=>"000001011",
  18598=>"110100110",
  18599=>"100110100",
  18600=>"111000001",
  18601=>"010100100",
  18602=>"100100000",
  18603=>"101100000",
  18604=>"101100100",
  18605=>"001100100",
  18606=>"110001110",
  18607=>"111110110",
  18608=>"011001011",
  18609=>"110110011",
  18610=>"110001111",
  18611=>"110101000",
  18612=>"111111101",
  18613=>"111011010",
  18614=>"111111001",
  18615=>"101111110",
  18616=>"000100111",
  18617=>"000100011",
  18618=>"010011100",
  18619=>"001100100",
  18620=>"011011010",
  18621=>"110110110",
  18622=>"100111111",
  18623=>"000001111",
  18624=>"011001001",
  18625=>"000001001",
  18626=>"000100110",
  18627=>"100111111",
  18628=>"011001001",
  18629=>"101100001",
  18630=>"110100100",
  18631=>"110110001",
  18632=>"100001101",
  18633=>"011001011",
  18634=>"000011001",
  18635=>"011011111",
  18636=>"111001001",
  18637=>"111111001",
  18638=>"011001011",
  18639=>"010001001",
  18640=>"111001000",
  18641=>"000000000",
  18642=>"000000000",
  18643=>"100000000",
  18644=>"011001011",
  18645=>"110011001",
  18646=>"001011000",
  18647=>"001011111",
  18648=>"011011111",
  18649=>"100100110",
  18650=>"000010100",
  18651=>"111001001",
  18652=>"001111000",
  18653=>"000110110",
  18654=>"011010010",
  18655=>"100000000",
  18656=>"011010101",
  18657=>"101110110",
  18658=>"111110100",
  18659=>"011011101",
  18660=>"111001001",
  18661=>"000001111",
  18662=>"111001101",
  18663=>"000011111",
  18664=>"100100101",
  18665=>"000100000",
  18666=>"000000101",
  18667=>"000010101",
  18668=>"110110100",
  18669=>"011001000",
  18670=>"100100100",
  18671=>"000000001",
  18672=>"011001011",
  18673=>"011010011",
  18674=>"011111111",
  18675=>"000000110",
  18676=>"011100101",
  18677=>"100001000",
  18678=>"001001001",
  18679=>"100011110",
  18680=>"000101010",
  18681=>"100001100",
  18682=>"101001001",
  18683=>"000010010",
  18684=>"011001001",
  18685=>"010000000",
  18686=>"111001001",
  18687=>"010001001",
  18688=>"000000100",
  18689=>"101000000",
  18690=>"010110110",
  18691=>"101000000",
  18692=>"110100110",
  18693=>"111100111",
  18694=>"111001000",
  18695=>"100111111",
  18696=>"000000000",
  18697=>"001111001",
  18698=>"000000000",
  18699=>"101000000",
  18700=>"100110111",
  18701=>"000000000",
  18702=>"000000000",
  18703=>"011111000",
  18704=>"100000000",
  18705=>"000000000",
  18706=>"000001000",
  18707=>"000101101",
  18708=>"111111000",
  18709=>"000011010",
  18710=>"111111111",
  18711=>"111111111",
  18712=>"000000000",
  18713=>"000000000",
  18714=>"111100101",
  18715=>"000011000",
  18716=>"101000000",
  18717=>"000000000",
  18718=>"000100111",
  18719=>"111111111",
  18720=>"010111111",
  18721=>"101000100",
  18722=>"101000000",
  18723=>"101111101",
  18724=>"110111100",
  18725=>"000000101",
  18726=>"000000000",
  18727=>"100000000",
  18728=>"011111011",
  18729=>"111111111",
  18730=>"000000110",
  18731=>"111100001",
  18732=>"110010010",
  18733=>"000000000",
  18734=>"000100000",
  18735=>"001111111",
  18736=>"111101101",
  18737=>"110100110",
  18738=>"101000101",
  18739=>"000000111",
  18740=>"000000000",
  18741=>"100000000",
  18742=>"001000000",
  18743=>"011011111",
  18744=>"011111001",
  18745=>"000000000",
  18746=>"000000111",
  18747=>"111111111",
  18748=>"100101000",
  18749=>"101111111",
  18750=>"000000000",
  18751=>"011011111",
  18752=>"111101111",
  18753=>"010010111",
  18754=>"101101100",
  18755=>"111110111",
  18756=>"000100100",
  18757=>"000010111",
  18758=>"101000000",
  18759=>"100101101",
  18760=>"000000010",
  18761=>"000000000",
  18762=>"000000000",
  18763=>"000111111",
  18764=>"010111011",
  18765=>"011001100",
  18766=>"100000111",
  18767=>"000000111",
  18768=>"100000000",
  18769=>"011011111",
  18770=>"000000000",
  18771=>"100100100",
  18772=>"111001101",
  18773=>"111111111",
  18774=>"010000000",
  18775=>"101000000",
  18776=>"000000000",
  18777=>"000000000",
  18778=>"111111111",
  18779=>"101011110",
  18780=>"000000000",
  18781=>"010000100",
  18782=>"010111111",
  18783=>"100001001",
  18784=>"101001000",
  18785=>"111000000",
  18786=>"000110000",
  18787=>"110111101",
  18788=>"001000000",
  18789=>"000000000",
  18790=>"000000000",
  18791=>"011111111",
  18792=>"010111011",
  18793=>"000000000",
  18794=>"100000111",
  18795=>"000000000",
  18796=>"011101111",
  18797=>"000000000",
  18798=>"111111010",
  18799=>"010000000",
  18800=>"011000000",
  18801=>"100111110",
  18802=>"001100000",
  18803=>"000000000",
  18804=>"000101100",
  18805=>"000000000",
  18806=>"000011010",
  18807=>"010010111",
  18808=>"111111111",
  18809=>"101001000",
  18810=>"001001001",
  18811=>"111100100",
  18812=>"011000100",
  18813=>"010001101",
  18814=>"000111111",
  18815=>"100100000",
  18816=>"000101100",
  18817=>"111111111",
  18818=>"110111000",
  18819=>"000101000",
  18820=>"000000111",
  18821=>"000000001",
  18822=>"000000001",
  18823=>"000000000",
  18824=>"001000001",
  18825=>"000100100",
  18826=>"000000000",
  18827=>"000000110",
  18828=>"011111011",
  18829=>"101110000",
  18830=>"010000000",
  18831=>"111100100",
  18832=>"000000000",
  18833=>"111111111",
  18834=>"111111111",
  18835=>"100100101",
  18836=>"000000000",
  18837=>"000111010",
  18838=>"111000000",
  18839=>"110110110",
  18840=>"001000001",
  18841=>"000111101",
  18842=>"000000011",
  18843=>"111111001",
  18844=>"000000000",
  18845=>"111111100",
  18846=>"000000101",
  18847=>"010000010",
  18848=>"111111111",
  18849=>"111101100",
  18850=>"000000000",
  18851=>"100000000",
  18852=>"000000010",
  18853=>"000000000",
  18854=>"001000001",
  18855=>"101011100",
  18856=>"100000000",
  18857=>"101001000",
  18858=>"001000111",
  18859=>"110000000",
  18860=>"111011111",
  18861=>"000100000",
  18862=>"011011110",
  18863=>"001111001",
  18864=>"111111111",
  18865=>"100000000",
  18866=>"010111111",
  18867=>"001000001",
  18868=>"110100000",
  18869=>"000000111",
  18870=>"111100000",
  18871=>"100000100",
  18872=>"001110100",
  18873=>"000000000",
  18874=>"000101000",
  18875=>"111101000",
  18876=>"000000000",
  18877=>"010111111",
  18878=>"110110110",
  18879=>"110111111",
  18880=>"000111001",
  18881=>"001001000",
  18882=>"000000000",
  18883=>"111111011",
  18884=>"000000000",
  18885=>"001101111",
  18886=>"111101100",
  18887=>"000011111",
  18888=>"100100001",
  18889=>"111111111",
  18890=>"000000000",
  18891=>"000010010",
  18892=>"000010010",
  18893=>"010000000",
  18894=>"111000110",
  18895=>"001100000",
  18896=>"000010011",
  18897=>"111010001",
  18898=>"000000000",
  18899=>"000000000",
  18900=>"000000111",
  18901=>"111000000",
  18902=>"011111000",
  18903=>"000000000",
  18904=>"011111111",
  18905=>"011100111",
  18906=>"111101101",
  18907=>"000010000",
  18908=>"011111111",
  18909=>"101001100",
  18910=>"000000000",
  18911=>"001111011",
  18912=>"000000111",
  18913=>"100000101",
  18914=>"100000000",
  18915=>"111000000",
  18916=>"110111000",
  18917=>"111111011",
  18918=>"111000000",
  18919=>"100100110",
  18920=>"100111111",
  18921=>"111111111",
  18922=>"100000000",
  18923=>"100000100",
  18924=>"101001000",
  18925=>"111111110",
  18926=>"110111000",
  18927=>"010110000",
  18928=>"000111011",
  18929=>"010000110",
  18930=>"111111111",
  18931=>"000000000",
  18932=>"000000000",
  18933=>"001111000",
  18934=>"000000000",
  18935=>"000000001",
  18936=>"000000000",
  18937=>"111001000",
  18938=>"100000000",
  18939=>"000000000",
  18940=>"111111110",
  18941=>"100110100",
  18942=>"100000110",
  18943=>"000000100",
  18944=>"011001000",
  18945=>"000000100",
  18946=>"101000101",
  18947=>"000000001",
  18948=>"000011011",
  18949=>"010010111",
  18950=>"010111010",
  18951=>"000010000",
  18952=>"000110000",
  18953=>"101011000",
  18954=>"000110010",
  18955=>"000000100",
  18956=>"000000000",
  18957=>"010011000",
  18958=>"000000110",
  18959=>"010010000",
  18960=>"110111000",
  18961=>"110111001",
  18962=>"000000100",
  18963=>"000000010",
  18964=>"000000100",
  18965=>"111101111",
  18966=>"000100101",
  18967=>"101111010",
  18968=>"101000000",
  18969=>"111101101",
  18970=>"000001101",
  18971=>"000000001",
  18972=>"100100100",
  18973=>"111110000",
  18974=>"111101111",
  18975=>"000010010",
  18976=>"010000101",
  18977=>"101100101",
  18978=>"000001111",
  18979=>"000000000",
  18980=>"001001001",
  18981=>"011010110",
  18982=>"001111111",
  18983=>"000111111",
  18984=>"111000000",
  18985=>"011000000",
  18986=>"000011000",
  18987=>"001000000",
  18988=>"010011011",
  18989=>"111011110",
  18990=>"011101100",
  18991=>"100010110",
  18992=>"000000110",
  18993=>"011101000",
  18994=>"101000000",
  18995=>"111111000",
  18996=>"000000000",
  18997=>"000000100",
  18998=>"000111110",
  18999=>"000000000",
  19000=>"111010000",
  19001=>"000111110",
  19002=>"010000000",
  19003=>"111111111",
  19004=>"001111110",
  19005=>"111111110",
  19006=>"000000000",
  19007=>"110111100",
  19008=>"001000100",
  19009=>"100000111",
  19010=>"000010010",
  19011=>"110100001",
  19012=>"111111111",
  19013=>"000101111",
  19014=>"000000000",
  19015=>"100101000",
  19016=>"000010011",
  19017=>"001011111",
  19018=>"111001100",
  19019=>"000111111",
  19020=>"100100100",
  19021=>"110110100",
  19022=>"100111111",
  19023=>"110111010",
  19024=>"111111101",
  19025=>"111000010",
  19026=>"000010111",
  19027=>"111111001",
  19028=>"000000000",
  19029=>"000011011",
  19030=>"000110110",
  19031=>"001000000",
  19032=>"100111111",
  19033=>"000010011",
  19034=>"000001100",
  19035=>"101101111",
  19036=>"001010000",
  19037=>"000000010",
  19038=>"010111111",
  19039=>"010100110",
  19040=>"101111111",
  19041=>"001001000",
  19042=>"111101101",
  19043=>"000101000",
  19044=>"000111010",
  19045=>"000011001",
  19046=>"000100101",
  19047=>"100000000",
  19048=>"000000111",
  19049=>"111000011",
  19050=>"011111000",
  19051=>"000011011",
  19052=>"000000111",
  19053=>"010110000",
  19054=>"101000000",
  19055=>"010111111",
  19056=>"100111101",
  19057=>"010000010",
  19058=>"111111011",
  19059=>"011101000",
  19060=>"111010000",
  19061=>"000001000",
  19062=>"000111111",
  19063=>"010101011",
  19064=>"001100011",
  19065=>"010000000",
  19066=>"110110111",
  19067=>"111100111",
  19068=>"110110010",
  19069=>"111100000",
  19070=>"101000001",
  19071=>"001001101",
  19072=>"111001101",
  19073=>"110100000",
  19074=>"011011111",
  19075=>"010010011",
  19076=>"111111101",
  19077=>"111101000",
  19078=>"110110001",
  19079=>"010110010",
  19080=>"110101100",
  19081=>"000110101",
  19082=>"010111000",
  19083=>"110001100",
  19084=>"101001101",
  19085=>"001010010",
  19086=>"000011110",
  19087=>"000000000",
  19088=>"001011001",
  19089=>"100101100",
  19090=>"000010000",
  19091=>"001101000",
  19092=>"000111111",
  19093=>"000111001",
  19094=>"000001111",
  19095=>"000010000",
  19096=>"000000000",
  19097=>"001101101",
  19098=>"000011011",
  19099=>"111100000",
  19100=>"000000000",
  19101=>"111101111",
  19102=>"011010000",
  19103=>"000000100",
  19104=>"001011111",
  19105=>"111011111",
  19106=>"111001000",
  19107=>"000000001",
  19108=>"000000011",
  19109=>"000000000",
  19110=>"100110110",
  19111=>"000011010",
  19112=>"011000111",
  19113=>"111111111",
  19114=>"000001101",
  19115=>"010111111",
  19116=>"111000000",
  19117=>"011011011",
  19118=>"100111111",
  19119=>"010010000",
  19120=>"000010000",
  19121=>"010111000",
  19122=>"000000010",
  19123=>"110000010",
  19124=>"000111000",
  19125=>"100011010",
  19126=>"000011111",
  19127=>"110110010",
  19128=>"000011011",
  19129=>"000111111",
  19130=>"000111110",
  19131=>"000000000",
  19132=>"110100111",
  19133=>"111101111",
  19134=>"011001111",
  19135=>"011010010",
  19136=>"001010000",
  19137=>"101000000",
  19138=>"011111000",
  19139=>"000011000",
  19140=>"000010000",
  19141=>"111110000",
  19142=>"000000111",
  19143=>"011111000",
  19144=>"111111111",
  19145=>"000101001",
  19146=>"110101101",
  19147=>"101100111",
  19148=>"000110000",
  19149=>"100011111",
  19150=>"010000101",
  19151=>"111111111",
  19152=>"111100101",
  19153=>"110111001",
  19154=>"000000111",
  19155=>"100100100",
  19156=>"000000001",
  19157=>"110100000",
  19158=>"000110000",
  19159=>"010010000",
  19160=>"100000000",
  19161=>"000010010",
  19162=>"001111011",
  19163=>"111101000",
  19164=>"000101110",
  19165=>"001001000",
  19166=>"000000000",
  19167=>"000000111",
  19168=>"000001001",
  19169=>"011011101",
  19170=>"000000000",
  19171=>"000011000",
  19172=>"010000000",
  19173=>"101000011",
  19174=>"000111111",
  19175=>"000111011",
  19176=>"100001111",
  19177=>"010010110",
  19178=>"000000100",
  19179=>"111000101",
  19180=>"111000000",
  19181=>"000100000",
  19182=>"100000000",
  19183=>"111000000",
  19184=>"010111111",
  19185=>"100011001",
  19186=>"111111011",
  19187=>"000111010",
  19188=>"000110001",
  19189=>"101000000",
  19190=>"000000000",
  19191=>"000011111",
  19192=>"000000100",
  19193=>"110111111",
  19194=>"110000000",
  19195=>"101001111",
  19196=>"111101111",
  19197=>"000000000",
  19198=>"000110000",
  19199=>"111100000",
  19200=>"001001100",
  19201=>"001000010",
  19202=>"111100101",
  19203=>"000010100",
  19204=>"000101111",
  19205=>"000000111",
  19206=>"001000111",
  19207=>"000100111",
  19208=>"011101000",
  19209=>"111001000",
  19210=>"001110110",
  19211=>"111101110",
  19212=>"111000000",
  19213=>"001000000",
  19214=>"001101101",
  19215=>"001000000",
  19216=>"000110101",
  19217=>"000000000",
  19218=>"110100000",
  19219=>"100000000",
  19220=>"111011100",
  19221=>"010100111",
  19222=>"001000000",
  19223=>"111000000",
  19224=>"000000001",
  19225=>"111100000",
  19226=>"000000010",
  19227=>"100000111",
  19228=>"000000000",
  19229=>"111111111",
  19230=>"010000101",
  19231=>"000000001",
  19232=>"011111011",
  19233=>"111011010",
  19234=>"000100010",
  19235=>"011011101",
  19236=>"110110000",
  19237=>"110100100",
  19238=>"010110110",
  19239=>"000010101",
  19240=>"010000000",
  19241=>"000001111",
  19242=>"111111101",
  19243=>"010010010",
  19244=>"111001101",
  19245=>"111111000",
  19246=>"010000111",
  19247=>"111111001",
  19248=>"000000101",
  19249=>"000100110",
  19250=>"000000010",
  19251=>"000000111",
  19252=>"010010010",
  19253=>"011010010",
  19254=>"101000000",
  19255=>"011111111",
  19256=>"110100001",
  19257=>"101100101",
  19258=>"010110100",
  19259=>"001011010",
  19260=>"000011101",
  19261=>"111111010",
  19262=>"000000000",
  19263=>"110000001",
  19264=>"111100001",
  19265=>"110000100",
  19266=>"100000010",
  19267=>"001100111",
  19268=>"001001000",
  19269=>"010000000",
  19270=>"000101111",
  19271=>"010011111",
  19272=>"100111111",
  19273=>"010111000",
  19274=>"101001111",
  19275=>"111010011",
  19276=>"111000000",
  19277=>"001100100",
  19278=>"001101001",
  19279=>"000000011",
  19280=>"000010011",
  19281=>"111110101",
  19282=>"101111111",
  19283=>"011101100",
  19284=>"000000000",
  19285=>"110110100",
  19286=>"010011000",
  19287=>"000000111",
  19288=>"000010010",
  19289=>"100101100",
  19290=>"000100011",
  19291=>"111111011",
  19292=>"111111010",
  19293=>"000011011",
  19294=>"111100100",
  19295=>"000000111",
  19296=>"000011010",
  19297=>"000001011",
  19298=>"101101101",
  19299=>"000010110",
  19300=>"001111101",
  19301=>"101011100",
  19302=>"000010011",
  19303=>"000100000",
  19304=>"010011111",
  19305=>"000000000",
  19306=>"111011101",
  19307=>"000000111",
  19308=>"000010010",
  19309=>"000111111",
  19310=>"011000000",
  19311=>"001000000",
  19312=>"111110001",
  19313=>"011000101",
  19314=>"101000001",
  19315=>"010100000",
  19316=>"000010011",
  19317=>"101000000",
  19318=>"000100001",
  19319=>"010000001",
  19320=>"111000010",
  19321=>"000010011",
  19322=>"110011101",
  19323=>"111111010",
  19324=>"011000000",
  19325=>"100001110",
  19326=>"010010010",
  19327=>"000000011",
  19328=>"111111101",
  19329=>"010100111",
  19330=>"000010010",
  19331=>"010111111",
  19332=>"100010011",
  19333=>"111111010",
  19334=>"011001001",
  19335=>"101111111",
  19336=>"001001100",
  19337=>"001010010",
  19338=>"111000001",
  19339=>"000010000",
  19340=>"000101010",
  19341=>"000101100",
  19342=>"101111100",
  19343=>"000001000",
  19344=>"100000001",
  19345=>"000000100",
  19346=>"101011010",
  19347=>"000101111",
  19348=>"000111011",
  19349=>"101100100",
  19350=>"100100110",
  19351=>"010110100",
  19352=>"000010111",
  19353=>"000000100",
  19354=>"010111000",
  19355=>"011001010",
  19356=>"100100100",
  19357=>"000011011",
  19358=>"011110111",
  19359=>"101100110",
  19360=>"101001000",
  19361=>"010000111",
  19362=>"100001111",
  19363=>"000000000",
  19364=>"010000100",
  19365=>"110110010",
  19366=>"110110001",
  19367=>"000000010",
  19368=>"010010010",
  19369=>"101010000",
  19370=>"000101100",
  19371=>"000000101",
  19372=>"011111001",
  19373=>"100100100",
  19374=>"000011111",
  19375=>"011101110",
  19376=>"000000000",
  19377=>"000111011",
  19378=>"100100000",
  19379=>"000000001",
  19380=>"001001010",
  19381=>"100001010",
  19382=>"111011000",
  19383=>"011011101",
  19384=>"100100001",
  19385=>"010110110",
  19386=>"110010010",
  19387=>"011100110",
  19388=>"010110110",
  19389=>"010111011",
  19390=>"011001000",
  19391=>"011000101",
  19392=>"110101000",
  19393=>"011101011",
  19394=>"011010001",
  19395=>"000100000",
  19396=>"011010000",
  19397=>"011110000",
  19398=>"011101000",
  19399=>"011111010",
  19400=>"110011000",
  19401=>"111000000",
  19402=>"011101000",
  19403=>"110000100",
  19404=>"100000001",
  19405=>"111100000",
  19406=>"000000000",
  19407=>"111010100",
  19408=>"111101101",
  19409=>"000001111",
  19410=>"100010111",
  19411=>"011000011",
  19412=>"100100000",
  19413=>"000000110",
  19414=>"101100111",
  19415=>"001000111",
  19416=>"000001001",
  19417=>"100000000",
  19418=>"111111010",
  19419=>"000000000",
  19420=>"001001000",
  19421=>"111100011",
  19422=>"000000011",
  19423=>"011000000",
  19424=>"101100010",
  19425=>"101100100",
  19426=>"001010111",
  19427=>"000101111",
  19428=>"000000001",
  19429=>"101111111",
  19430=>"000010111",
  19431=>"000001111",
  19432=>"111000011",
  19433=>"000000011",
  19434=>"110011111",
  19435=>"111110000",
  19436=>"111100000",
  19437=>"011010000",
  19438=>"110000000",
  19439=>"001111111",
  19440=>"001000010",
  19441=>"111001001",
  19442=>"111000000",
  19443=>"100101110",
  19444=>"011001001",
  19445=>"000000111",
  19446=>"000000011",
  19447=>"001001100",
  19448=>"111000000",
  19449=>"110110010",
  19450=>"101111101",
  19451=>"000111111",
  19452=>"000000000",
  19453=>"011011111",
  19454=>"001011000",
  19455=>"111000111",
  19456=>"000011100",
  19457=>"000100111",
  19458=>"101000100",
  19459=>"101101100",
  19460=>"101000011",
  19461=>"110000100",
  19462=>"000000000",
  19463=>"000010111",
  19464=>"001100000",
  19465=>"101000100",
  19466=>"101001001",
  19467=>"000100100",
  19468=>"111100100",
  19469=>"111100000",
  19470=>"100100000",
  19471=>"010011111",
  19472=>"100100100",
  19473=>"001001000",
  19474=>"010001011",
  19475=>"000000000",
  19476=>"111101000",
  19477=>"111000000",
  19478=>"010000101",
  19479=>"000100000",
  19480=>"100100010",
  19481=>"001111111",
  19482=>"101100000",
  19483=>"000010000",
  19484=>"000100000",
  19485=>"011111011",
  19486=>"111101100",
  19487=>"001101101",
  19488=>"101000000",
  19489=>"101010001",
  19490=>"100011000",
  19491=>"000000100",
  19492=>"101001000",
  19493=>"001011110",
  19494=>"111000000",
  19495=>"100100000",
  19496=>"101011011",
  19497=>"001100000",
  19498=>"110100100",
  19499=>"010010011",
  19500=>"111111011",
  19501=>"101000100",
  19502=>"111011111",
  19503=>"000110100",
  19504=>"000100111",
  19505=>"000101011",
  19506=>"101000000",
  19507=>"000000111",
  19508=>"000011100",
  19509=>"000010111",
  19510=>"000110110",
  19511=>"111100100",
  19512=>"011011110",
  19513=>"101100100",
  19514=>"101100100",
  19515=>"000011010",
  19516=>"011000011",
  19517=>"111101110",
  19518=>"000100000",
  19519=>"110011011",
  19520=>"000000000",
  19521=>"010111011",
  19522=>"011100000",
  19523=>"111100100",
  19524=>"111100101",
  19525=>"111101100",
  19526=>"001100100",
  19527=>"010000111",
  19528=>"010011100",
  19529=>"111011000",
  19530=>"000101101",
  19531=>"101100100",
  19532=>"010010100",
  19533=>"000000110",
  19534=>"101111111",
  19535=>"110011010",
  19536=>"111011011",
  19537=>"111010111",
  19538=>"110100100",
  19539=>"011001000",
  19540=>"100101111",
  19541=>"010010010",
  19542=>"111100111",
  19543=>"101101101",
  19544=>"000000000",
  19545=>"110100000",
  19546=>"001001000",
  19547=>"100010011",
  19548=>"100000100",
  19549=>"001001001",
  19550=>"100111111",
  19551=>"100100100",
  19552=>"111000000",
  19553=>"111111101",
  19554=>"101100100",
  19555=>"110101100",
  19556=>"000000010",
  19557=>"000100100",
  19558=>"000110001",
  19559=>"010010100",
  19560=>"111000000",
  19561=>"111011101",
  19562=>"111111101",
  19563=>"011111010",
  19564=>"100000111",
  19565=>"000000010",
  19566=>"101100100",
  19567=>"000000011",
  19568=>"100111111",
  19569=>"100111101",
  19570=>"000011001",
  19571=>"000000000",
  19572=>"111111111",
  19573=>"000100100",
  19574=>"100000111",
  19575=>"000001000",
  19576=>"111000000",
  19577=>"010000000",
  19578=>"100111011",
  19579=>"111000000",
  19580=>"000011011",
  19581=>"111000000",
  19582=>"011010000",
  19583=>"101000000",
  19584=>"000010110",
  19585=>"000011000",
  19586=>"000011001",
  19587=>"000000000",
  19588=>"111111111",
  19589=>"111100000",
  19590=>"010010011",
  19591=>"100001110",
  19592=>"100111111",
  19593=>"011100010",
  19594=>"100100111",
  19595=>"111111101",
  19596=>"100011011",
  19597=>"000011011",
  19598=>"010000000",
  19599=>"010000000",
  19600=>"001001001",
  19601=>"000111011",
  19602=>"000111011",
  19603=>"100100010",
  19604=>"000100111",
  19605=>"111100100",
  19606=>"111100111",
  19607=>"100100100",
  19608=>"001011111",
  19609=>"000011011",
  19610=>"101011011",
  19611=>"010000000",
  19612=>"011100100",
  19613=>"000000001",
  19614=>"000100100",
  19615=>"111100111",
  19616=>"000010011",
  19617=>"001000010",
  19618=>"000011011",
  19619=>"011010000",
  19620=>"000000001",
  19621=>"001111110",
  19622=>"001000101",
  19623=>"000010011",
  19624=>"000000100",
  19625=>"111000101",
  19626=>"001000000",
  19627=>"111100100",
  19628=>"100000000",
  19629=>"101100101",
  19630=>"011110101",
  19631=>"000000011",
  19632=>"101000001",
  19633=>"001011000",
  19634=>"010001011",
  19635=>"001010011",
  19636=>"110111011",
  19637=>"000000000",
  19638=>"000010011",
  19639=>"110011110",
  19640=>"010011010",
  19641=>"000000011",
  19642=>"000011011",
  19643=>"111111011",
  19644=>"111111111",
  19645=>"111111111",
  19646=>"101000000",
  19647=>"010011111",
  19648=>"000000000",
  19649=>"110000000",
  19650=>"010111011",
  19651=>"001001001",
  19652=>"111101000",
  19653=>"001000010",
  19654=>"000110111",
  19655=>"111000100",
  19656=>"111111110",
  19657=>"000000000",
  19658=>"001111111",
  19659=>"111100100",
  19660=>"100011001",
  19661=>"000011111",
  19662=>"010111111",
  19663=>"000000001",
  19664=>"011100000",
  19665=>"101001101",
  19666=>"000010011",
  19667=>"111110110",
  19668=>"101011000",
  19669=>"100100111",
  19670=>"111100100",
  19671=>"000100100",
  19672=>"000010010",
  19673=>"000100111",
  19674=>"101000011",
  19675=>"100000000",
  19676=>"111110011",
  19677=>"111111000",
  19678=>"100111000",
  19679=>"100100111",
  19680=>"111100001",
  19681=>"101100100",
  19682=>"100000000",
  19683=>"111100101",
  19684=>"100000000",
  19685=>"110111111",
  19686=>"000000011",
  19687=>"010000110",
  19688=>"010000000",
  19689=>"011111111",
  19690=>"110000000",
  19691=>"111100100",
  19692=>"000011011",
  19693=>"111100100",
  19694=>"001001001",
  19695=>"000000111",
  19696=>"000000000",
  19697=>"100110111",
  19698=>"010000000",
  19699=>"011101010",
  19700=>"101000001",
  19701=>"011000011",
  19702=>"000000000",
  19703=>"010011011",
  19704=>"000010000",
  19705=>"010010100",
  19706=>"111000001",
  19707=>"000101101",
  19708=>"111100100",
  19709=>"000011011",
  19710=>"011111111",
  19711=>"000000001",
  19712=>"011001100",
  19713=>"000000100",
  19714=>"000010000",
  19715=>"101101100",
  19716=>"111100001",
  19717=>"001001000",
  19718=>"010101101",
  19719=>"111000101",
  19720=>"111100101",
  19721=>"000001000",
  19722=>"000010110",
  19723=>"111000110",
  19724=>"000100100",
  19725=>"111111111",
  19726=>"100000001",
  19727=>"001101001",
  19728=>"000000010",
  19729=>"000000111",
  19730=>"000000000",
  19731=>"000100111",
  19732=>"001110010",
  19733=>"000110111",
  19734=>"011000010",
  19735=>"001111110",
  19736=>"000000000",
  19737=>"000001111",
  19738=>"001000100",
  19739=>"000011000",
  19740=>"111111111",
  19741=>"111000000",
  19742=>"111111010",
  19743=>"000101101",
  19744=>"000000110",
  19745=>"001101100",
  19746=>"000111100",
  19747=>"011101111",
  19748=>"100100010",
  19749=>"110111111",
  19750=>"000000111",
  19751=>"000010111",
  19752=>"111010111",
  19753=>"111111111",
  19754=>"000111011",
  19755=>"100111000",
  19756=>"110011011",
  19757=>"011111011",
  19758=>"111101000",
  19759=>"000000000",
  19760=>"011111000",
  19761=>"011110100",
  19762=>"111000000",
  19763=>"111011010",
  19764=>"000001011",
  19765=>"101111111",
  19766=>"000100111",
  19767=>"000111000",
  19768=>"111111000",
  19769=>"011111001",
  19770=>"111000000",
  19771=>"111111000",
  19772=>"001101011",
  19773=>"010010111",
  19774=>"000010010",
  19775=>"000001011",
  19776=>"111101101",
  19777=>"101101001",
  19778=>"001111000",
  19779=>"000100110",
  19780=>"110000000",
  19781=>"111000000",
  19782=>"000011110",
  19783=>"010100000",
  19784=>"111100001",
  19785=>"111001001",
  19786=>"010000101",
  19787=>"000010110",
  19788=>"000100101",
  19789=>"011000111",
  19790=>"110001000",
  19791=>"100110100",
  19792=>"000000111",
  19793=>"111100000",
  19794=>"100110111",
  19795=>"001000110",
  19796=>"101100010",
  19797=>"101111100",
  19798=>"100101111",
  19799=>"000010000",
  19800=>"111000111",
  19801=>"110011111",
  19802=>"001100110",
  19803=>"000110111",
  19804=>"000101111",
  19805=>"011000000",
  19806=>"010111111",
  19807=>"000001011",
  19808=>"100000000",
  19809=>"000010010",
  19810=>"100111011",
  19811=>"000000111",
  19812=>"010000000",
  19813=>"111011101",
  19814=>"010101101",
  19815=>"000000100",
  19816=>"010000000",
  19817=>"011111000",
  19818=>"011100010",
  19819=>"001000101",
  19820=>"011011001",
  19821=>"010010111",
  19822=>"000000000",
  19823=>"011001001",
  19824=>"110101101",
  19825=>"111111000",
  19826=>"000001111",
  19827=>"111000110",
  19828=>"000000101",
  19829=>"100000101",
  19830=>"001000110",
  19831=>"000111111",
  19832=>"000010010",
  19833=>"000111111",
  19834=>"010010101",
  19835=>"011010000",
  19836=>"110000000",
  19837=>"100100001",
  19838=>"111111011",
  19839=>"000000011",
  19840=>"101001011",
  19841=>"110000001",
  19842=>"111111001",
  19843=>"110111000",
  19844=>"011001101",
  19845=>"000000001",
  19846=>"111101100",
  19847=>"000000110",
  19848=>"001100000",
  19849=>"010000000",
  19850=>"111000011",
  19851=>"100100110",
  19852=>"110111000",
  19853=>"010111111",
  19854=>"000111101",
  19855=>"000001001",
  19856=>"111100110",
  19857=>"100000100",
  19858=>"000101111",
  19859=>"111000010",
  19860=>"000000000",
  19861=>"001000000",
  19862=>"000110000",
  19863=>"011000100",
  19864=>"000111111",
  19865=>"111010010",
  19866=>"000011000",
  19867=>"000011111",
  19868=>"111000000",
  19869=>"000111111",
  19870=>"000111000",
  19871=>"000000000",
  19872=>"100111011",
  19873=>"011110010",
  19874=>"100111000",
  19875=>"100000111",
  19876=>"111111101",
  19877=>"000000011",
  19878=>"011000001",
  19879=>"000111000",
  19880=>"011010000",
  19881=>"000000111",
  19882=>"111001111",
  19883=>"000000111",
  19884=>"100111000",
  19885=>"000111011",
  19886=>"011101101",
  19887=>"011010111",
  19888=>"100000000",
  19889=>"011010111",
  19890=>"000000000",
  19891=>"000001001",
  19892=>"110100100",
  19893=>"100011000",
  19894=>"100000110",
  19895=>"011000100",
  19896=>"101110110",
  19897=>"010100010",
  19898=>"101111011",
  19899=>"101001000",
  19900=>"110110011",
  19901=>"000000111",
  19902=>"011000100",
  19903=>"111000000",
  19904=>"000000110",
  19905=>"000000010",
  19906=>"101001100",
  19907=>"011000000",
  19908=>"001010000",
  19909=>"100011001",
  19910=>"111101000",
  19911=>"000011110",
  19912=>"000000110",
  19913=>"000100100",
  19914=>"010110010",
  19915=>"000101101",
  19916=>"010000011",
  19917=>"011000110",
  19918=>"000000010",
  19919=>"111111000",
  19920=>"011000010",
  19921=>"010001011",
  19922=>"011111101",
  19923=>"101101111",
  19924=>"000111111",
  19925=>"000000111",
  19926=>"000100111",
  19927=>"000111110",
  19928=>"111000000",
  19929=>"111111111",
  19930=>"111011110",
  19931=>"000000010",
  19932=>"101001000",
  19933=>"000000100",
  19934=>"100100010",
  19935=>"110101000",
  19936=>"111000000",
  19937=>"111000010",
  19938=>"111111011",
  19939=>"001000111",
  19940=>"000000111",
  19941=>"101101101",
  19942=>"001000111",
  19943=>"110001111",
  19944=>"010111111",
  19945=>"000110000",
  19946=>"000011011",
  19947=>"001001111",
  19948=>"000111100",
  19949=>"000000101",
  19950=>"000000000",
  19951=>"111010110",
  19952=>"011100100",
  19953=>"000111000",
  19954=>"111111000",
  19955=>"100011001",
  19956=>"100100010",
  19957=>"000000001",
  19958=>"000000111",
  19959=>"011011000",
  19960=>"111111000",
  19961=>"010000000",
  19962=>"111011111",
  19963=>"010000001",
  19964=>"100111111",
  19965=>"000000111",
  19966=>"011100100",
  19967=>"100111110",
  19968=>"000000100",
  19969=>"110110111",
  19970=>"000110111",
  19971=>"110000100",
  19972=>"110111111",
  19973=>"001101000",
  19974=>"011111111",
  19975=>"110110101",
  19976=>"000001011",
  19977=>"111000111",
  19978=>"000010000",
  19979=>"000000000",
  19980=>"001001111",
  19981=>"111001101",
  19982=>"000000000",
  19983=>"001001010",
  19984=>"111000000",
  19985=>"001001011",
  19986=>"000111111",
  19987=>"011001001",
  19988=>"111011000",
  19989=>"000100100",
  19990=>"011111011",
  19991=>"000000001",
  19992=>"000101111",
  19993=>"000001101",
  19994=>"001101001",
  19995=>"111111111",
  19996=>"110111111",
  19997=>"000000000",
  19998=>"000000000",
  19999=>"110111000",
  20000=>"000001000",
  20001=>"000001010",
  20002=>"101111111",
  20003=>"110011001",
  20004=>"100100100",
  20005=>"011000011",
  20006=>"110111001",
  20007=>"111001000",
  20008=>"010000010",
  20009=>"000000001",
  20010=>"110001000",
  20011=>"111000000",
  20012=>"001111101",
  20013=>"010000000",
  20014=>"101111001",
  20015=>"111111000",
  20016=>"000001000",
  20017=>"001000000",
  20018=>"000111110",
  20019=>"111000010",
  20020=>"101000010",
  20021=>"111011000",
  20022=>"000000010",
  20023=>"101000000",
  20024=>"000000111",
  20025=>"111001100",
  20026=>"100001010",
  20027=>"000000111",
  20028=>"011110100",
  20029=>"010010111",
  20030=>"000000000",
  20031=>"100000000",
  20032=>"000100111",
  20033=>"000000100",
  20034=>"111000001",
  20035=>"001001000",
  20036=>"111000000",
  20037=>"010000100",
  20038=>"000001011",
  20039=>"000000000",
  20040=>"111111111",
  20041=>"110111110",
  20042=>"101001111",
  20043=>"000101001",
  20044=>"000000101",
  20045=>"011001111",
  20046=>"110001001",
  20047=>"110000001",
  20048=>"000000000",
  20049=>"000111111",
  20050=>"000001001",
  20051=>"001000000",
  20052=>"010010000",
  20053=>"110111110",
  20054=>"000011010",
  20055=>"100000111",
  20056=>"000110111",
  20057=>"110000011",
  20058=>"111011000",
  20059=>"000000000",
  20060=>"110000001",
  20061=>"111110100",
  20062=>"110111111",
  20063=>"001110110",
  20064=>"000111111",
  20065=>"010000000",
  20066=>"001001111",
  20067=>"101111001",
  20068=>"001001001",
  20069=>"000110010",
  20070=>"001001110",
  20071=>"110001001",
  20072=>"110111100",
  20073=>"000111110",
  20074=>"111100011",
  20075=>"100000000",
  20076=>"111111110",
  20077=>"111111001",
  20078=>"110001011",
  20079=>"001100101",
  20080=>"000000001",
  20081=>"010000000",
  20082=>"011001000",
  20083=>"111000000",
  20084=>"101001001",
  20085=>"000101111",
  20086=>"001011100",
  20087=>"000001001",
  20088=>"101111000",
  20089=>"111110111",
  20090=>"000001001",
  20091=>"000010111",
  20092=>"011011110",
  20093=>"100000000",
  20094=>"110010110",
  20095=>"001111111",
  20096=>"010001001",
  20097=>"001110010",
  20098=>"001001001",
  20099=>"111110100",
  20100=>"101001000",
  20101=>"001110111",
  20102=>"000000100",
  20103=>"011001101",
  20104=>"001001111",
  20105=>"000000001",
  20106=>"101011001",
  20107=>"010000000",
  20108=>"111111000",
  20109=>"000101111",
  20110=>"000100101",
  20111=>"100000000",
  20112=>"111011000",
  20113=>"000100111",
  20114=>"100000100",
  20115=>"111001111",
  20116=>"111000000",
  20117=>"001000101",
  20118=>"001111111",
  20119=>"011000000",
  20120=>"011001001",
  20121=>"100110010",
  20122=>"000110111",
  20123=>"110001111",
  20124=>"011001011",
  20125=>"111100001",
  20126=>"000000111",
  20127=>"101000111",
  20128=>"001111111",
  20129=>"110110010",
  20130=>"110000000",
  20131=>"101111111",
  20132=>"001111000",
  20133=>"000000000",
  20134=>"100000000",
  20135=>"001000000",
  20136=>"010000111",
  20137=>"000000111",
  20138=>"101111111",
  20139=>"000000111",
  20140=>"111000001",
  20141=>"000000111",
  20142=>"100110011",
  20143=>"111001110",
  20144=>"000001001",
  20145=>"011000110",
  20146=>"101001001",
  20147=>"101001100",
  20148=>"110111000",
  20149=>"111111111",
  20150=>"000101111",
  20151=>"101110011",
  20152=>"110011001",
  20153=>"110001000",
  20154=>"010000010",
  20155=>"111111110",
  20156=>"011001011",
  20157=>"111111111",
  20158=>"100001011",
  20159=>"000000000",
  20160=>"010110001",
  20161=>"111000101",
  20162=>"111000000",
  20163=>"010001111",
  20164=>"000000011",
  20165=>"100001001",
  20166=>"111111000",
  20167=>"010010101",
  20168=>"010101101",
  20169=>"000011011",
  20170=>"110011111",
  20171=>"000110111",
  20172=>"000000111",
  20173=>"100100110",
  20174=>"111110000",
  20175=>"001111110",
  20176=>"111111111",
  20177=>"111100110",
  20178=>"000000101",
  20179=>"101101001",
  20180=>"000000111",
  20181=>"111111101",
  20182=>"111000001",
  20183=>"001000000",
  20184=>"111000000",
  20185=>"011000000",
  20186=>"100110111",
  20187=>"001001111",
  20188=>"111111100",
  20189=>"010110000",
  20190=>"000001001",
  20191=>"000000101",
  20192=>"001001011",
  20193=>"000000111",
  20194=>"110111111",
  20195=>"000100011",
  20196=>"111001001",
  20197=>"011111101",
  20198=>"001001000",
  20199=>"111111000",
  20200=>"001000000",
  20201=>"111111111",
  20202=>"001100100",
  20203=>"000101111",
  20204=>"011111111",
  20205=>"000001000",
  20206=>"000000111",
  20207=>"111101101",
  20208=>"111000100",
  20209=>"001000100",
  20210=>"000101001",
  20211=>"110101000",
  20212=>"111010000",
  20213=>"111111101",
  20214=>"101000010",
  20215=>"100000000",
  20216=>"001001111",
  20217=>"001111110",
  20218=>"111110010",
  20219=>"000110000",
  20220=>"101111100",
  20221=>"010000000",
  20222=>"000101011",
  20223=>"001000000",
  20224=>"001010111",
  20225=>"010000101",
  20226=>"000000101",
  20227=>"000100110",
  20228=>"011011110",
  20229=>"011111000",
  20230=>"111111001",
  20231=>"111011100",
  20232=>"011111000",
  20233=>"111100000",
  20234=>"000000000",
  20235=>"111000000",
  20236=>"111111010",
  20237=>"110011001",
  20238=>"000001001",
  20239=>"111111001",
  20240=>"011011111",
  20241=>"101000111",
  20242=>"110000000",
  20243=>"110000000",
  20244=>"111111111",
  20245=>"011001101",
  20246=>"000010111",
  20247=>"101010011",
  20248=>"100000000",
  20249=>"011101001",
  20250=>"010010100",
  20251=>"010111111",
  20252=>"111111111",
  20253=>"000101101",
  20254=>"010000000",
  20255=>"001010100",
  20256=>"100010000",
  20257=>"111111100",
  20258=>"000000100",
  20259=>"111110000",
  20260=>"111011011",
  20261=>"010100100",
  20262=>"000000101",
  20263=>"011111011",
  20264=>"000000111",
  20265=>"000111110",
  20266=>"101111101",
  20267=>"000000011",
  20268=>"111111111",
  20269=>"111111100",
  20270=>"111000100",
  20271=>"000100100",
  20272=>"000110111",
  20273=>"111011000",
  20274=>"000000000",
  20275=>"001000011",
  20276=>"000000111",
  20277=>"000000001",
  20278=>"000001011",
  20279=>"001000111",
  20280=>"000001111",
  20281=>"000000111",
  20282=>"111001000",
  20283=>"000000000",
  20284=>"110101000",
  20285=>"111111000",
  20286=>"000000000",
  20287=>"010110000",
  20288=>"111111110",
  20289=>"101011000",
  20290=>"101111111",
  20291=>"010111110",
  20292=>"111111111",
  20293=>"011111111",
  20294=>"111111010",
  20295=>"010000110",
  20296=>"110101111",
  20297=>"111000000",
  20298=>"100000001",
  20299=>"000101110",
  20300=>"110101000",
  20301=>"111111111",
  20302=>"001111001",
  20303=>"111111100",
  20304=>"000000000",
  20305=>"111111000",
  20306=>"011011010",
  20307=>"000001111",
  20308=>"111100000",
  20309=>"000000001",
  20310=>"100110111",
  20311=>"001000000",
  20312=>"011000000",
  20313=>"000011000",
  20314=>"110110110",
  20315=>"111111111",
  20316=>"100000100",
  20317=>"100110111",
  20318=>"111111111",
  20319=>"000011001",
  20320=>"000000000",
  20321=>"001000100",
  20322=>"110010000",
  20323=>"011011001",
  20324=>"001000111",
  20325=>"000011010",
  20326=>"000000110",
  20327=>"011111111",
  20328=>"111110111",
  20329=>"111010000",
  20330=>"111000000",
  20331=>"111111101",
  20332=>"000000000",
  20333=>"011111111",
  20334=>"001011000",
  20335=>"011110001",
  20336=>"110111100",
  20337=>"000010111",
  20338=>"000000100",
  20339=>"000000111",
  20340=>"110001111",
  20341=>"001100101",
  20342=>"010011111",
  20343=>"000000000",
  20344=>"010111110",
  20345=>"010000000",
  20346=>"000000101",
  20347=>"111111000",
  20348=>"000100000",
  20349=>"000000110",
  20350=>"111111111",
  20351=>"000000100",
  20352=>"000101110",
  20353=>"111111100",
  20354=>"010111000",
  20355=>"001111111",
  20356=>"010111111",
  20357=>"000000111",
  20358=>"000011011",
  20359=>"110000010",
  20360=>"101001100",
  20361=>"011111111",
  20362=>"110100111",
  20363=>"111001100",
  20364=>"000001111",
  20365=>"111111010",
  20366=>"100100000",
  20367=>"000000000",
  20368=>"100110111",
  20369=>"110000000",
  20370=>"000011111",
  20371=>"100001001",
  20372=>"010101111",
  20373=>"010000000",
  20374=>"111010111",
  20375=>"001011000",
  20376=>"000000000",
  20377=>"111111000",
  20378=>"000000000",
  20379=>"100000000",
  20380=>"111111100",
  20381=>"101001111",
  20382=>"111011111",
  20383=>"000001111",
  20384=>"111111110",
  20385=>"000000111",
  20386=>"000000101",
  20387=>"000000010",
  20388=>"101001000",
  20389=>"000100010",
  20390=>"111000101",
  20391=>"111001111",
  20392=>"000001000",
  20393=>"100000110",
  20394=>"000011111",
  20395=>"010000000",
  20396=>"110101100",
  20397=>"000000111",
  20398=>"000001010",
  20399=>"001000010",
  20400=>"000000000",
  20401=>"100100110",
  20402=>"101100010",
  20403=>"100110111",
  20404=>"101111010",
  20405=>"001000101",
  20406=>"011100000",
  20407=>"010110101",
  20408=>"011010000",
  20409=>"001110111",
  20410=>"000001001",
  20411=>"111000001",
  20412=>"111100011",
  20413=>"011111000",
  20414=>"111111000",
  20415=>"101001000",
  20416=>"111000010",
  20417=>"000000000",
  20418=>"010000110",
  20419=>"011001111",
  20420=>"000000101",
  20421=>"000000010",
  20422=>"000111111",
  20423=>"111111000",
  20424=>"111011000",
  20425=>"000101100",
  20426=>"000000111",
  20427=>"000000101",
  20428=>"000000100",
  20429=>"000101011",
  20430=>"000001111",
  20431=>"111111011",
  20432=>"111111010",
  20433=>"110000001",
  20434=>"010110100",
  20435=>"011111000",
  20436=>"101000000",
  20437=>"011001111",
  20438=>"110111110",
  20439=>"110100000",
  20440=>"000000101",
  20441=>"011010000",
  20442=>"110111111",
  20443=>"100000100",
  20444=>"100011111",
  20445=>"111111111",
  20446=>"001000100",
  20447=>"010100111",
  20448=>"111111111",
  20449=>"011011100",
  20450=>"111111000",
  20451=>"011111110",
  20452=>"101000000",
  20453=>"111111011",
  20454=>"111011010",
  20455=>"011000100",
  20456=>"111110111",
  20457=>"010000011",
  20458=>"000000000",
  20459=>"100000000",
  20460=>"000100000",
  20461=>"111011001",
  20462=>"000100000",
  20463=>"000000000",
  20464=>"000000000",
  20465=>"001000010",
  20466=>"101000110",
  20467=>"000110010",
  20468=>"111000011",
  20469=>"101000101",
  20470=>"011000000",
  20471=>"000100001",
  20472=>"111111000",
  20473=>"111111110",
  20474=>"011110011",
  20475=>"000000110",
  20476=>"001000111",
  20477=>"000000000",
  20478=>"110000101",
  20479=>"101000111",
  20480=>"001001100",
  20481=>"000111000",
  20482=>"000000101",
  20483=>"000100111",
  20484=>"001000001",
  20485=>"111000111",
  20486=>"000001000",
  20487=>"101001110",
  20488=>"000111111",
  20489=>"001111111",
  20490=>"000111011",
  20491=>"000000000",
  20492=>"010010000",
  20493=>"011000000",
  20494=>"101011001",
  20495=>"001000001",
  20496=>"111111010",
  20497=>"111111111",
  20498=>"000001000",
  20499=>"001111111",
  20500=>"111100000",
  20501=>"101111111",
  20502=>"100001111",
  20503=>"001001000",
  20504=>"000000000",
  20505=>"111111001",
  20506=>"111011111",
  20507=>"100000000",
  20508=>"000000001",
  20509=>"011010111",
  20510=>"111101111",
  20511=>"111000101",
  20512=>"011000001",
  20513=>"110010010",
  20514=>"101101100",
  20515=>"111000000",
  20516=>"111111001",
  20517=>"111100111",
  20518=>"010111111",
  20519=>"111111011",
  20520=>"000111110",
  20521=>"101111111",
  20522=>"100010000",
  20523=>"010010110",
  20524=>"001111111",
  20525=>"000010101",
  20526=>"111111111",
  20527=>"110000110",
  20528=>"010000111",
  20529=>"001011011",
  20530=>"100000111",
  20531=>"011111111",
  20532=>"000000000",
  20533=>"101011111",
  20534=>"001000100",
  20535=>"101100101",
  20536=>"111100010",
  20537=>"000000000",
  20538=>"000000001",
  20539=>"111101101",
  20540=>"110110010",
  20541=>"001111111",
  20542=>"000000000",
  20543=>"000100110",
  20544=>"111101111",
  20545=>"001000101",
  20546=>"100111111",
  20547=>"000100111",
  20548=>"101101111",
  20549=>"000111111",
  20550=>"111111101",
  20551=>"110110000",
  20552=>"110000000",
  20553=>"000110010",
  20554=>"000010111",
  20555=>"000001101",
  20556=>"000100110",
  20557=>"100100000",
  20558=>"000100110",
  20559=>"110111111",
  20560=>"111000000",
  20561=>"000111110",
  20562=>"000000101",
  20563=>"001001010",
  20564=>"000001111",
  20565=>"111110000",
  20566=>"001011001",
  20567=>"000100111",
  20568=>"000100111",
  20569=>"100011001",
  20570=>"100001011",
  20571=>"010000000",
  20572=>"111111111",
  20573=>"001001000",
  20574=>"111100000",
  20575=>"001011110",
  20576=>"000000011",
  20577=>"010001000",
  20578=>"101000000",
  20579=>"000000001",
  20580=>"001101000",
  20581=>"111111100",
  20582=>"100010000",
  20583=>"100111111",
  20584=>"000000110",
  20585=>"000000000",
  20586=>"111111001",
  20587=>"111101100",
  20588=>"111101000",
  20589=>"010110110",
  20590=>"011000000",
  20591=>"110111011",
  20592=>"001101010",
  20593=>"111010111",
  20594=>"111100000",
  20595=>"110100011",
  20596=>"111111000",
  20597=>"100100111",
  20598=>"000000011",
  20599=>"101100100",
  20600=>"000000010",
  20601=>"101100001",
  20602=>"011111101",
  20603=>"000000000",
  20604=>"100111110",
  20605=>"100101001",
  20606=>"110010011",
  20607=>"000000000",
  20608=>"111000000",
  20609=>"000000000",
  20610=>"111111111",
  20611=>"111100010",
  20612=>"000010111",
  20613=>"111111111",
  20614=>"111011110",
  20615=>"111111000",
  20616=>"000111011",
  20617=>"111101000",
  20618=>"000111111",
  20619=>"111010000",
  20620=>"000001101",
  20621=>"111111111",
  20622=>"100000001",
  20623=>"001100111",
  20624=>"111110000",
  20625=>"000000000",
  20626=>"000000000",
  20627=>"010111011",
  20628=>"111111010",
  20629=>"111110110",
  20630=>"111101000",
  20631=>"010101111",
  20632=>"000100000",
  20633=>"000000111",
  20634=>"000000010",
  20635=>"000001011",
  20636=>"000110110",
  20637=>"010000001",
  20638=>"011000000",
  20639=>"010000000",
  20640=>"011011000",
  20641=>"111100111",
  20642=>"110110000",
  20643=>"000001111",
  20644=>"111010001",
  20645=>"110010000",
  20646=>"111111111",
  20647=>"101111101",
  20648=>"111101111",
  20649=>"110110101",
  20650=>"111000000",
  20651=>"000011000",
  20652=>"111111101",
  20653=>"000001111",
  20654=>"010100001",
  20655=>"101111101",
  20656=>"000000000",
  20657=>"111111000",
  20658=>"000000001",
  20659=>"000110000",
  20660=>"000010011",
  20661=>"101101111",
  20662=>"111111100",
  20663=>"110111111",
  20664=>"011001000",
  20665=>"111111011",
  20666=>"111100111",
  20667=>"111000111",
  20668=>"010100010",
  20669=>"011101101",
  20670=>"101011101",
  20671=>"000111111",
  20672=>"010010000",
  20673=>"001000000",
  20674=>"001110111",
  20675=>"000101110",
  20676=>"000000000",
  20677=>"111110000",
  20678=>"000100000",
  20679=>"110000010",
  20680=>"111111000",
  20681=>"110101000",
  20682=>"010100000",
  20683=>"101001000",
  20684=>"000111111",
  20685=>"001111001",
  20686=>"111101000",
  20687=>"000000001",
  20688=>"000111111",
  20689=>"011110100",
  20690=>"111110110",
  20691=>"100000000",
  20692=>"111010000",
  20693=>"111100000",
  20694=>"000101101",
  20695=>"000011011",
  20696=>"000000001",
  20697=>"111111111",
  20698=>"110110110",
  20699=>"000000000",
  20700=>"111000011",
  20701=>"000111111",
  20702=>"111111111",
  20703=>"110111111",
  20704=>"000010111",
  20705=>"111000111",
  20706=>"111000001",
  20707=>"111100010",
  20708=>"000111000",
  20709=>"111101101",
  20710=>"101100110",
  20711=>"110100110",
  20712=>"010000111",
  20713=>"110110111",
  20714=>"001001000",
  20715=>"001101000",
  20716=>"000111100",
  20717=>"110000000",
  20718=>"000010010",
  20719=>"000000000",
  20720=>"010010110",
  20721=>"110010000",
  20722=>"111110111",
  20723=>"000110010",
  20724=>"100011001",
  20725=>"101101101",
  20726=>"000000000",
  20727=>"000010111",
  20728=>"000000000",
  20729=>"000000000",
  20730=>"111111001",
  20731=>"111111110",
  20732=>"011010000",
  20733=>"110000000",
  20734=>"001001000",
  20735=>"110000000",
  20736=>"100110100",
  20737=>"000000000",
  20738=>"000010000",
  20739=>"110101001",
  20740=>"001001000",
  20741=>"010000000",
  20742=>"000000000",
  20743=>"101101011",
  20744=>"101000000",
  20745=>"111101110",
  20746=>"000000111",
  20747=>"111001001",
  20748=>"101101111",
  20749=>"100101101",
  20750=>"000000010",
  20751=>"000111101",
  20752=>"000001000",
  20753=>"111000011",
  20754=>"111111010",
  20755=>"011100100",
  20756=>"011010000",
  20757=>"011000001",
  20758=>"110111011",
  20759=>"101010110",
  20760=>"111101110",
  20761=>"010011111",
  20762=>"000010010",
  20763=>"000111010",
  20764=>"010111000",
  20765=>"111101001",
  20766=>"000000100",
  20767=>"111010010",
  20768=>"111110000",
  20769=>"100001111",
  20770=>"000111111",
  20771=>"100011111",
  20772=>"100100110",
  20773=>"011011010",
  20774=>"000010110",
  20775=>"111001011",
  20776=>"101001011",
  20777=>"100001001",
  20778=>"000000000",
  20779=>"100100010",
  20780=>"010010000",
  20781=>"000000101",
  20782=>"000111110",
  20783=>"011101001",
  20784=>"111101100",
  20785=>"100100110",
  20786=>"100101111",
  20787=>"010000000",
  20788=>"100000101",
  20789=>"111011000",
  20790=>"111000010",
  20791=>"000100000",
  20792=>"101101101",
  20793=>"101101000",
  20794=>"011001010",
  20795=>"101010000",
  20796=>"110011110",
  20797=>"001010100",
  20798=>"111000100",
  20799=>"000000000",
  20800=>"111111000",
  20801=>"010010101",
  20802=>"110000000",
  20803=>"100000001",
  20804=>"111111011",
  20805=>"101101001",
  20806=>"100000001",
  20807=>"111000000",
  20808=>"110110110",
  20809=>"100100000",
  20810=>"101101101",
  20811=>"000000000",
  20812=>"011010000",
  20813=>"001001010",
  20814=>"111011011",
  20815=>"111111001",
  20816=>"000100101",
  20817=>"111110100",
  20818=>"101100100",
  20819=>"110011011",
  20820=>"111100111",
  20821=>"000000000",
  20822=>"001111010",
  20823=>"000100101",
  20824=>"100001000",
  20825=>"011011010",
  20826=>"000001000",
  20827=>"100100000",
  20828=>"000000110",
  20829=>"000100110",
  20830=>"100010000",
  20831=>"001000011",
  20832=>"011011010",
  20833=>"011001010",
  20834=>"101101111",
  20835=>"100001001",
  20836=>"101001011",
  20837=>"000100110",
  20838=>"101101110",
  20839=>"100101011",
  20840=>"000000010",
  20841=>"111000000",
  20842=>"010000111",
  20843=>"111111001",
  20844=>"111110010",
  20845=>"111001010",
  20846=>"000000101",
  20847=>"000111000",
  20848=>"101100111",
  20849=>"000000000",
  20850=>"011000000",
  20851=>"000001000",
  20852=>"000100011",
  20853=>"010000000",
  20854=>"100000010",
  20855=>"001001000",
  20856=>"010010111",
  20857=>"000011010",
  20858=>"111000111",
  20859=>"111100110",
  20860=>"111010100",
  20861=>"011100000",
  20862=>"101100111",
  20863=>"101000100",
  20864=>"111100000",
  20865=>"010100101",
  20866=>"000101101",
  20867=>"011111111",
  20868=>"100000111",
  20869=>"001001101",
  20870=>"100110111",
  20871=>"001010110",
  20872=>"000000011",
  20873=>"101111111",
  20874=>"010000000",
  20875=>"100010000",
  20876=>"100100101",
  20877=>"000011000",
  20878=>"101100000",
  20879=>"100000000",
  20880=>"111011001",
  20881=>"000100000",
  20882=>"000100111",
  20883=>"101100000",
  20884=>"000110000",
  20885=>"000100000",
  20886=>"000000000",
  20887=>"100100110",
  20888=>"111101000",
  20889=>"110000000",
  20890=>"101000100",
  20891=>"000010000",
  20892=>"110101101",
  20893=>"111100101",
  20894=>"000100101",
  20895=>"011101010",
  20896=>"110010110",
  20897=>"001111111",
  20898=>"101000000",
  20899=>"000101101",
  20900=>"110001111",
  20901=>"010011011",
  20902=>"101111111",
  20903=>"111111011",
  20904=>"000100000",
  20905=>"000001000",
  20906=>"110111000",
  20907=>"010101100",
  20908=>"111111100",
  20909=>"100101111",
  20910=>"011011001",
  20911=>"000000111",
  20912=>"000101110",
  20913=>"110001110",
  20914=>"010100010",
  20915=>"011000011",
  20916=>"110110110",
  20917=>"111010101",
  20918=>"000010011",
  20919=>"110111101",
  20920=>"011010011",
  20921=>"100011001",
  20922=>"000111110",
  20923=>"000100110",
  20924=>"111011011",
  20925=>"010101101",
  20926=>"100000000",
  20927=>"101000000",
  20928=>"111111111",
  20929=>"000000000",
  20930=>"011111000",
  20931=>"110100000",
  20932=>"011101111",
  20933=>"111110001",
  20934=>"101100000",
  20935=>"101000010",
  20936=>"010111010",
  20937=>"000010000",
  20938=>"010011110",
  20939=>"010000000",
  20940=>"001000000",
  20941=>"111110110",
  20942=>"010111000",
  20943=>"011101101",
  20944=>"011111001",
  20945=>"000001010",
  20946=>"011011111",
  20947=>"000110000",
  20948=>"101001000",
  20949=>"001001011",
  20950=>"010011001",
  20951=>"100000000",
  20952=>"100000101",
  20953=>"011000000",
  20954=>"000010001",
  20955=>"111101101",
  20956=>"110110110",
  20957=>"000101101",
  20958=>"001111111",
  20959=>"000000001",
  20960=>"110011111",
  20961=>"000100111",
  20962=>"010001011",
  20963=>"110100111",
  20964=>"000000000",
  20965=>"111101110",
  20966=>"000101000",
  20967=>"010110001",
  20968=>"100101100",
  20969=>"101011000",
  20970=>"000000001",
  20971=>"001101111",
  20972=>"101000111",
  20973=>"111101111",
  20974=>"010000011",
  20975=>"010111111",
  20976=>"010000001",
  20977=>"100100000",
  20978=>"000111011",
  20979=>"001010010",
  20980=>"001001011",
  20981=>"100100000",
  20982=>"111100101",
  20983=>"010000000",
  20984=>"001101101",
  20985=>"001111111",
  20986=>"111111110",
  20987=>"111000000",
  20988=>"111000000",
  20989=>"010010000",
  20990=>"000100100",
  20991=>"110010110",
  20992=>"011101010",
  20993=>"000001000",
  20994=>"100000111",
  20995=>"000000000",
  20996=>"011111111",
  20997=>"010000000",
  20998=>"010010110",
  20999=>"000010111",
  21000=>"111101110",
  21001=>"000001000",
  21002=>"000100100",
  21003=>"111001011",
  21004=>"000000000",
  21005=>"011111010",
  21006=>"101011010",
  21007=>"001101110",
  21008=>"000010110",
  21009=>"101000111",
  21010=>"001101000",
  21011=>"111000000",
  21012=>"111111111",
  21013=>"001000100",
  21014=>"111100011",
  21015=>"011000111",
  21016=>"101100111",
  21017=>"111101111",
  21018=>"000100100",
  21019=>"000111010",
  21020=>"110111101",
  21021=>"101000000",
  21022=>"111111000",
  21023=>"011001000",
  21024=>"111111111",
  21025=>"010111111",
  21026=>"000000000",
  21027=>"000011011",
  21028=>"000000100",
  21029=>"111100111",
  21030=>"111110101",
  21031=>"001111101",
  21032=>"010111001",
  21033=>"010110000",
  21034=>"111111101",
  21035=>"111101010",
  21036=>"001000000",
  21037=>"110010111",
  21038=>"111111011",
  21039=>"000001100",
  21040=>"001111111",
  21041=>"000100011",
  21042=>"011011111",
  21043=>"110000100",
  21044=>"000000000",
  21045=>"111110101",
  21046=>"010001011",
  21047=>"000000111",
  21048=>"111011000",
  21049=>"000000001",
  21050=>"000000011",
  21051=>"111111100",
  21052=>"110100111",
  21053=>"000001001",
  21054=>"010000001",
  21055=>"111111011",
  21056=>"111001000",
  21057=>"101101011",
  21058=>"000000000",
  21059=>"001110000",
  21060=>"110010010",
  21061=>"000000111",
  21062=>"101111111",
  21063=>"001000111",
  21064=>"110000000",
  21065=>"111111000",
  21066=>"111000000",
  21067=>"000000101",
  21068=>"000001000",
  21069=>"001100111",
  21070=>"111001111",
  21071=>"111011111",
  21072=>"111000111",
  21073=>"010111101",
  21074=>"000000010",
  21075=>"001001100",
  21076=>"111000000",
  21077=>"010100100",
  21078=>"000101001",
  21079=>"000111111",
  21080=>"110101000",
  21081=>"111100010",
  21082=>"110110111",
  21083=>"111110111",
  21084=>"000000000",
  21085=>"111001011",
  21086=>"010111100",
  21087=>"101010100",
  21088=>"100110000",
  21089=>"000111011",
  21090=>"000010100",
  21091=>"001011011",
  21092=>"111101101",
  21093=>"001001000",
  21094=>"001100000",
  21095=>"111000000",
  21096=>"111111111",
  21097=>"011111000",
  21098=>"010110111",
  21099=>"111001000",
  21100=>"111111110",
  21101=>"000000001",
  21102=>"111110000",
  21103=>"000101011",
  21104=>"000110100",
  21105=>"001000011",
  21106=>"010100110",
  21107=>"001000100",
  21108=>"000000111",
  21109=>"101000000",
  21110=>"000111111",
  21111=>"111000000",
  21112=>"111111111",
  21113=>"000000000",
  21114=>"000110111",
  21115=>"000010000",
  21116=>"000111000",
  21117=>"110100001",
  21118=>"001101111",
  21119=>"111111111",
  21120=>"000111000",
  21121=>"111000001",
  21122=>"111111110",
  21123=>"111111000",
  21124=>"110000000",
  21125=>"111111000",
  21126=>"110001110",
  21127=>"000001011",
  21128=>"011011111",
  21129=>"111000010",
  21130=>"111111111",
  21131=>"001001111",
  21132=>"000000001",
  21133=>"000000100",
  21134=>"010111111",
  21135=>"000000100",
  21136=>"110110100",
  21137=>"001000000",
  21138=>"000000101",
  21139=>"000000011",
  21140=>"100111111",
  21141=>"000111100",
  21142=>"000010000",
  21143=>"001000000",
  21144=>"010111100",
  21145=>"111000000",
  21146=>"111011000",
  21147=>"001000000",
  21148=>"111010100",
  21149=>"111000101",
  21150=>"010011111",
  21151=>"101100000",
  21152=>"010100000",
  21153=>"010010111",
  21154=>"111011010",
  21155=>"010010000",
  21156=>"000001010",
  21157=>"111111110",
  21158=>"000000010",
  21159=>"100111010",
  21160=>"111000110",
  21161=>"000000000",
  21162=>"001100101",
  21163=>"110101010",
  21164=>"001111000",
  21165=>"100000010",
  21166=>"110100000",
  21167=>"000000000",
  21168=>"011000000",
  21169=>"011000100",
  21170=>"010001000",
  21171=>"101100000",
  21172=>"101001000",
  21173=>"111111110",
  21174=>"011111111",
  21175=>"011001101",
  21176=>"001001011",
  21177=>"001111101",
  21178=>"111011001",
  21179=>"110110111",
  21180=>"000100100",
  21181=>"111111110",
  21182=>"111110011",
  21183=>"101000000",
  21184=>"010000000",
  21185=>"011010010",
  21186=>"000100011",
  21187=>"011111000",
  21188=>"000011000",
  21189=>"110110100",
  21190=>"010011101",
  21191=>"111001000",
  21192=>"101111111",
  21193=>"000000000",
  21194=>"111111111",
  21195=>"111111001",
  21196=>"111111111",
  21197=>"110111110",
  21198=>"101001110",
  21199=>"010110111",
  21200=>"010000000",
  21201=>"110000110",
  21202=>"010010111",
  21203=>"000111010",
  21204=>"001000101",
  21205=>"010000001",
  21206=>"111111000",
  21207=>"010110110",
  21208=>"111000111",
  21209=>"000000010",
  21210=>"011011011",
  21211=>"000000000",
  21212=>"010011111",
  21213=>"011111111",
  21214=>"111111000",
  21215=>"010101111",
  21216=>"000111011",
  21217=>"000010111",
  21218=>"111000001",
  21219=>"011000111",
  21220=>"111100101",
  21221=>"000100000",
  21222=>"001000010",
  21223=>"011100101",
  21224=>"000101010",
  21225=>"000000011",
  21226=>"100101001",
  21227=>"000111000",
  21228=>"111111010",
  21229=>"111101111",
  21230=>"001010001",
  21231=>"000111111",
  21232=>"000000000",
  21233=>"011001001",
  21234=>"111000000",
  21235=>"110100000",
  21236=>"010000111",
  21237=>"101110111",
  21238=>"101100111",
  21239=>"100011000",
  21240=>"000001010",
  21241=>"000111001",
  21242=>"111111111",
  21243=>"000000000",
  21244=>"000000110",
  21245=>"111111000",
  21246=>"100101010",
  21247=>"010000101",
  21248=>"010101101",
  21249=>"110110100",
  21250=>"111100100",
  21251=>"111000011",
  21252=>"110100100",
  21253=>"111101000",
  21254=>"000001010",
  21255=>"010111011",
  21256=>"000001011",
  21257=>"110100100",
  21258=>"100100110",
  21259=>"000011011",
  21260=>"000001001",
  21261=>"100101101",
  21262=>"111011001",
  21263=>"001101111",
  21264=>"111110110",
  21265=>"011100110",
  21266=>"011110000",
  21267=>"001011000",
  21268=>"000011010",
  21269=>"111100101",
  21270=>"110110010",
  21271=>"100011001",
  21272=>"000100110",
  21273=>"001011011",
  21274=>"000110100",
  21275=>"111110110",
  21276=>"011000000",
  21277=>"011110111",
  21278=>"000100000",
  21279=>"100111011",
  21280=>"111110100",
  21281=>"100101101",
  21282=>"010000000",
  21283=>"001011011",
  21284=>"100011011",
  21285=>"001000010",
  21286=>"000011011",
  21287=>"000011011",
  21288=>"111100111",
  21289=>"000100100",
  21290=>"100100001",
  21291=>"111100100",
  21292=>"000011000",
  21293=>"010001011",
  21294=>"000100100",
  21295=>"001001101",
  21296=>"000011000",
  21297=>"100000100",
  21298=>"111111011",
  21299=>"000110100",
  21300=>"111100100",
  21301=>"111111111",
  21302=>"110110110",
  21303=>"100100100",
  21304=>"000100000",
  21305=>"000000001",
  21306=>"000011011",
  21307=>"100110110",
  21308=>"001011011",
  21309=>"001011001",
  21310=>"001000000",
  21311=>"000000111",
  21312=>"111011000",
  21313=>"000100110",
  21314=>"110100110",
  21315=>"111100100",
  21316=>"000001000",
  21317=>"010011001",
  21318=>"011000011",
  21319=>"110011001",
  21320=>"110001000",
  21321=>"011011100",
  21322=>"000111011",
  21323=>"111100111",
  21324=>"110101000",
  21325=>"000000101",
  21326=>"100111111",
  21327=>"111110101",
  21328=>"111110101",
  21329=>"011111000",
  21330=>"011011011",
  21331=>"001001000",
  21332=>"111001111",
  21333=>"001110000",
  21334=>"010111111",
  21335=>"011000000",
  21336=>"101011011",
  21337=>"000001001",
  21338=>"110000001",
  21339=>"100000011",
  21340=>"110100100",
  21341=>"011000000",
  21342=>"111110110",
  21343=>"111100000",
  21344=>"000000001",
  21345=>"111110100",
  21346=>"010100100",
  21347=>"111110110",
  21348=>"000000011",
  21349=>"000001100",
  21350=>"110100001",
  21351=>"111010000",
  21352=>"000111111",
  21353=>"011000100",
  21354=>"111100111",
  21355=>"011011001",
  21356=>"011111100",
  21357=>"001100100",
  21358=>"000000001",
  21359=>"010000011",
  21360=>"000000000",
  21361=>"000100011",
  21362=>"110100100",
  21363=>"001011011",
  21364=>"000100100",
  21365=>"001100000",
  21366=>"111100001",
  21367=>"000000101",
  21368=>"010100000",
  21369=>"010101011",
  21370=>"000100001",
  21371=>"000011100",
  21372=>"111001001",
  21373=>"000010010",
  21374=>"111100110",
  21375=>"100100100",
  21376=>"001101100",
  21377=>"000110110",
  21378=>"110011000",
  21379=>"010011011",
  21380=>"000010001",
  21381=>"111010110",
  21382=>"000000001",
  21383=>"010110010",
  21384=>"101011011",
  21385=>"000100111",
  21386=>"110110110",
  21387=>"011011100",
  21388=>"110110110",
  21389=>"111100100",
  21390=>"011011000",
  21391=>"111100111",
  21392=>"110010010",
  21393=>"101110110",
  21394=>"111110011",
  21395=>"111111000",
  21396=>"001011010",
  21397=>"111100100",
  21398=>"100001111",
  21399=>"011100110",
  21400=>"110011001",
  21401=>"000011011",
  21402=>"000001001",
  21403=>"111100100",
  21404=>"000001001",
  21405=>"110100100",
  21406=>"111100010",
  21407=>"011111001",
  21408=>"100100010",
  21409=>"111110100",
  21410=>"110110110",
  21411=>"011001011",
  21412=>"000100001",
  21413=>"010011011",
  21414=>"011011010",
  21415=>"010100000",
  21416=>"011000000",
  21417=>"111110111",
  21418=>"111100100",
  21419=>"000100100",
  21420=>"110011000",
  21421=>"000001001",
  21422=>"000111110",
  21423=>"100110010",
  21424=>"000000000",
  21425=>"111100100",
  21426=>"001111110",
  21427=>"000001010",
  21428=>"101001011",
  21429=>"110101110",
  21430=>"000001000",
  21431=>"110000001",
  21432=>"110001011",
  21433=>"000010000",
  21434=>"001011011",
  21435=>"000011100",
  21436=>"100001001",
  21437=>"000111110",
  21438=>"011010000",
  21439=>"001001001",
  21440=>"100000000",
  21441=>"000100111",
  21442=>"111110110",
  21443=>"100100111",
  21444=>"000010001",
  21445=>"110100000",
  21446=>"011011011",
  21447=>"111100100",
  21448=>"000011111",
  21449=>"110100100",
  21450=>"011011110",
  21451=>"111100100",
  21452=>"100100110",
  21453=>"011100001",
  21454=>"100100001",
  21455=>"110111011",
  21456=>"000001001",
  21457=>"000000001",
  21458=>"111000001",
  21459=>"000000010",
  21460=>"011100100",
  21461=>"101000000",
  21462=>"010011011",
  21463=>"001011110",
  21464=>"001011111",
  21465=>"100001000",
  21466=>"000010110",
  21467=>"111100110",
  21468=>"101010001",
  21469=>"000011011",
  21470=>"001001011",
  21471=>"000110100",
  21472=>"100000100",
  21473=>"001011010",
  21474=>"110001000",
  21475=>"011110000",
  21476=>"011000100",
  21477=>"111100100",
  21478=>"000011011",
  21479=>"100011001",
  21480=>"100000001",
  21481=>"011000000",
  21482=>"111001001",
  21483=>"011110110",
  21484=>"100100100",
  21485=>"000001001",
  21486=>"000000010",
  21487=>"111101000",
  21488=>"001011010",
  21489=>"000010010",
  21490=>"000000000",
  21491=>"011011111",
  21492=>"001010110",
  21493=>"001100000",
  21494=>"001000001",
  21495=>"011100000",
  21496=>"010110111",
  21497=>"000111111",
  21498=>"001011011",
  21499=>"000011000",
  21500=>"000000000",
  21501=>"111110110",
  21502=>"100111100",
  21503=>"111100000",
  21504=>"001011001",
  21505=>"101001011",
  21506=>"101111111",
  21507=>"001000000",
  21508=>"110111000",
  21509=>"000000101",
  21510=>"011011010",
  21511=>"111110110",
  21512=>"001000100",
  21513=>"000000000",
  21514=>"000000100",
  21515=>"111111001",
  21516=>"111111101",
  21517=>"000000000",
  21518=>"111110011",
  21519=>"111111111",
  21520=>"101101110",
  21521=>"000000000",
  21522=>"000000000",
  21523=>"011111111",
  21524=>"000111011",
  21525=>"000000010",
  21526=>"011011000",
  21527=>"111111010",
  21528=>"000000000",
  21529=>"000011000",
  21530=>"101111111",
  21531=>"111011100",
  21532=>"111111110",
  21533=>"111111111",
  21534=>"000000111",
  21535=>"001001111",
  21536=>"100001000",
  21537=>"001000001",
  21538=>"101100000",
  21539=>"111111111",
  21540=>"110111000",
  21541=>"111111110",
  21542=>"000010111",
  21543=>"111111100",
  21544=>"000101111",
  21545=>"000001010",
  21546=>"100100100",
  21547=>"101111001",
  21548=>"111111111",
  21549=>"000000000",
  21550=>"111100101",
  21551=>"000001001",
  21552=>"101101111",
  21553=>"100100101",
  21554=>"100000010",
  21555=>"000100000",
  21556=>"000000101",
  21557=>"000111110",
  21558=>"100000100",
  21559=>"111110000",
  21560=>"000000000",
  21561=>"111000001",
  21562=>"111111111",
  21563=>"111111100",
  21564=>"111111111",
  21565=>"011111111",
  21566=>"000000000",
  21567=>"011010110",
  21568=>"101100100",
  21569=>"000001111",
  21570=>"010000000",
  21571=>"011000001",
  21572=>"111011001",
  21573=>"000000010",
  21574=>"111111111",
  21575=>"000000000",
  21576=>"111011110",
  21577=>"101101011",
  21578=>"101000111",
  21579=>"111111111",
  21580=>"000000100",
  21581=>"111111110",
  21582=>"111100010",
  21583=>"111111110",
  21584=>"000000111",
  21585=>"111111111",
  21586=>"001101001",
  21587=>"001111001",
  21588=>"000000001",
  21589=>"110111111",
  21590=>"111100000",
  21591=>"000000100",
  21592=>"100111100",
  21593=>"111111101",
  21594=>"000011011",
  21595=>"101111011",
  21596=>"000000001",
  21597=>"001001001",
  21598=>"011000100",
  21599=>"100000001",
  21600=>"000010111",
  21601=>"101101101",
  21602=>"000110111",
  21603=>"000100100",
  21604=>"110010000",
  21605=>"111111100",
  21606=>"111000000",
  21607=>"000000000",
  21608=>"110001001",
  21609=>"000110000",
  21610=>"001000000",
  21611=>"010011111",
  21612=>"111001000",
  21613=>"000000010",
  21614=>"111101000",
  21615=>"111011000",
  21616=>"011011010",
  21617=>"111100000",
  21618=>"011000001",
  21619=>"000000111",
  21620=>"000000111",
  21621=>"000000001",
  21622=>"100110111",
  21623=>"100000000",
  21624=>"111011000",
  21625=>"000011000",
  21626=>"001110110",
  21627=>"001111010",
  21628=>"110100010",
  21629=>"100100110",
  21630=>"111011010",
  21631=>"000010111",
  21632=>"111001001",
  21633=>"100100000",
  21634=>"000111111",
  21635=>"111111111",
  21636=>"000000110",
  21637=>"111111011",
  21638=>"101001001",
  21639=>"001100110",
  21640=>"100100101",
  21641=>"111110011",
  21642=>"000000001",
  21643=>"000000000",
  21644=>"100000001",
  21645=>"000111000",
  21646=>"111111001",
  21647=>"000001010",
  21648=>"100100000",
  21649=>"000000001",
  21650=>"110000101",
  21651=>"111101111",
  21652=>"111101101",
  21653=>"000000100",
  21654=>"111111101",
  21655=>"100000000",
  21656=>"111111000",
  21657=>"111111111",
  21658=>"000111111",
  21659=>"000010000",
  21660=>"011001101",
  21661=>"100000111",
  21662=>"111000010",
  21663=>"111111000",
  21664=>"001110100",
  21665=>"001001011",
  21666=>"101100101",
  21667=>"111111011",
  21668=>"001111111",
  21669=>"001011101",
  21670=>"111010010",
  21671=>"101110000",
  21672=>"000111001",
  21673=>"000000000",
  21674=>"000101010",
  21675=>"000000000",
  21676=>"101111011",
  21677=>"000110111",
  21678=>"110110110",
  21679=>"010000000",
  21680=>"101000111",
  21681=>"011001001",
  21682=>"000111111",
  21683=>"000100000",
  21684=>"111111000",
  21685=>"000000000",
  21686=>"111100111",
  21687=>"111111011",
  21688=>"111110111",
  21689=>"111100110",
  21690=>"010111111",
  21691=>"110001111",
  21692=>"000011010",
  21693=>"000000010",
  21694=>"000011011",
  21695=>"000000000",
  21696=>"000001000",
  21697=>"110110100",
  21698=>"000001001",
  21699=>"001011011",
  21700=>"110110010",
  21701=>"111011001",
  21702=>"111111111",
  21703=>"000110111",
  21704=>"111111010",
  21705=>"111010000",
  21706=>"000000111",
  21707=>"101000000",
  21708=>"000110111",
  21709=>"001111011",
  21710=>"000000110",
  21711=>"000100000",
  21712=>"011011010",
  21713=>"011000001",
  21714=>"000100101",
  21715=>"111111101",
  21716=>"010111101",
  21717=>"000100100",
  21718=>"000000101",
  21719=>"111000000",
  21720=>"111111010",
  21721=>"011000000",
  21722=>"100100001",
  21723=>"000000000",
  21724=>"111111000",
  21725=>"011100000",
  21726=>"011111100",
  21727=>"111100110",
  21728=>"000011001",
  21729=>"001000101",
  21730=>"111111111",
  21731=>"000111110",
  21732=>"000000000",
  21733=>"000111111",
  21734=>"111110100",
  21735=>"011011011",
  21736=>"000000000",
  21737=>"011000111",
  21738=>"000000001",
  21739=>"101111111",
  21740=>"100111111",
  21741=>"010000000",
  21742=>"010010010",
  21743=>"010111111",
  21744=>"111111111",
  21745=>"000100100",
  21746=>"011001001",
  21747=>"111111101",
  21748=>"110100100",
  21749=>"000000000",
  21750=>"000000111",
  21751=>"111111111",
  21752=>"111000000",
  21753=>"101001110",
  21754=>"000101000",
  21755=>"111111111",
  21756=>"000111111",
  21757=>"011101111",
  21758=>"001011101",
  21759=>"010010010",
  21760=>"000001001",
  21761=>"011111111",
  21762=>"000000000",
  21763=>"100111111",
  21764=>"001100101",
  21765=>"111101111",
  21766=>"110000100",
  21767=>"101000111",
  21768=>"000100111",
  21769=>"010000000",
  21770=>"110011001",
  21771=>"001000011",
  21772=>"011001101",
  21773=>"011010000",
  21774=>"100000100",
  21775=>"111000000",
  21776=>"111111000",
  21777=>"010010000",
  21778=>"000000000",
  21779=>"111111111",
  21780=>"000111101",
  21781=>"101111010",
  21782=>"000000100",
  21783=>"111111000",
  21784=>"111111101",
  21785=>"101111110",
  21786=>"111110010",
  21787=>"000111111",
  21788=>"000011000",
  21789=>"010010000",
  21790=>"110101101",
  21791=>"001000011",
  21792=>"000000000",
  21793=>"010101111",
  21794=>"010010100",
  21795=>"000010110",
  21796=>"110110111",
  21797=>"000010111",
  21798=>"111110010",
  21799=>"111101000",
  21800=>"101000101",
  21801=>"001101111",
  21802=>"000000000",
  21803=>"101111111",
  21804=>"100000110",
  21805=>"111111011",
  21806=>"000000001",
  21807=>"101101001",
  21808=>"110111000",
  21809=>"011101000",
  21810=>"101110111",
  21811=>"101000000",
  21812=>"111111000",
  21813=>"111001000",
  21814=>"111111110",
  21815=>"000111111",
  21816=>"000111100",
  21817=>"000000111",
  21818=>"000000110",
  21819=>"111110000",
  21820=>"001000110",
  21821=>"000101011",
  21822=>"000000100",
  21823=>"111111111",
  21824=>"111010000",
  21825=>"011101111",
  21826=>"000111000",
  21827=>"001100001",
  21828=>"111000000",
  21829=>"000000000",
  21830=>"010000001",
  21831=>"111000000",
  21832=>"001111111",
  21833=>"101001010",
  21834=>"100111101",
  21835=>"101111000",
  21836=>"000010111",
  21837=>"001001110",
  21838=>"100100000",
  21839=>"111111111",
  21840=>"001000111",
  21841=>"011111000",
  21842=>"011100010",
  21843=>"001000001",
  21844=>"110110000",
  21845=>"000101100",
  21846=>"011011001",
  21847=>"000000000",
  21848=>"000001111",
  21849=>"001001011",
  21850=>"100100011",
  21851=>"111110011",
  21852=>"000001111",
  21853=>"000000111",
  21854=>"111010000",
  21855=>"000100110",
  21856=>"111101000",
  21857=>"001000000",
  21858=>"000111111",
  21859=>"001001110",
  21860=>"001100111",
  21861=>"000000000",
  21862=>"100111101",
  21863=>"000111010",
  21864=>"111000000",
  21865=>"000000101",
  21866=>"100000111",
  21867=>"000101111",
  21868=>"111100111",
  21869=>"110110010",
  21870=>"000100001",
  21871=>"001110110",
  21872=>"100101111",
  21873=>"101100000",
  21874=>"111011001",
  21875=>"111000000",
  21876=>"111111000",
  21877=>"101111010",
  21878=>"111000000",
  21879=>"111111000",
  21880=>"111101010",
  21881=>"110001101",
  21882=>"000001000",
  21883=>"111101000",
  21884=>"000001111",
  21885=>"100000100",
  21886=>"100000000",
  21887=>"000000101",
  21888=>"000000000",
  21889=>"000001011",
  21890=>"111111111",
  21891=>"011111110",
  21892=>"000000100",
  21893=>"000010000",
  21894=>"000110011",
  21895=>"100000011",
  21896=>"001100110",
  21897=>"010111101",
  21898=>"010011111",
  21899=>"101100000",
  21900=>"000000111",
  21901=>"000000111",
  21902=>"000001111",
  21903=>"001001000",
  21904=>"001001011",
  21905=>"101001100",
  21906=>"111000010",
  21907=>"010010010",
  21908=>"000010101",
  21909=>"000101001",
  21910=>"000101111",
  21911=>"000001011",
  21912=>"111111111",
  21913=>"000001111",
  21914=>"111000000",
  21915=>"111000000",
  21916=>"000000101",
  21917=>"111001111",
  21918=>"111111011",
  21919=>"000000000",
  21920=>"101111011",
  21921=>"000000000",
  21922=>"100101110",
  21923=>"111111111",
  21924=>"110000100",
  21925=>"111110100",
  21926=>"100000000",
  21927=>"101000011",
  21928=>"001111110",
  21929=>"000000111",
  21930=>"100000101",
  21931=>"111000000",
  21932=>"010111110",
  21933=>"000000101",
  21934=>"000000110",
  21935=>"011000001",
  21936=>"101111101",
  21937=>"001001111",
  21938=>"111111110",
  21939=>"000110111",
  21940=>"111111000",
  21941=>"111000000",
  21942=>"111111000",
  21943=>"101000100",
  21944=>"100100111",
  21945=>"000000110",
  21946=>"000000110",
  21947=>"111010000",
  21948=>"000110111",
  21949=>"111110010",
  21950=>"101111011",
  21951=>"000101100",
  21952=>"111111000",
  21953=>"011111111",
  21954=>"100111001",
  21955=>"100100110",
  21956=>"111111001",
  21957=>"100000111",
  21958=>"010010110",
  21959=>"111000000",
  21960=>"000000000",
  21961=>"100000000",
  21962=>"101000110",
  21963=>"111111001",
  21964=>"011111101",
  21965=>"000100011",
  21966=>"111001101",
  21967=>"000011111",
  21968=>"111010000",
  21969=>"000100111",
  21970=>"000000111",
  21971=>"100100001",
  21972=>"000000111",
  21973=>"000110111",
  21974=>"000001111",
  21975=>"111111111",
  21976=>"111111000",
  21977=>"000010010",
  21978=>"111100100",
  21979=>"111000000",
  21980=>"000111001",
  21981=>"000000111",
  21982=>"111111100",
  21983=>"110111100",
  21984=>"111101000",
  21985=>"000101111",
  21986=>"111011000",
  21987=>"000000001",
  21988=>"000001010",
  21989=>"101111101",
  21990=>"000000111",
  21991=>"000000111",
  21992=>"111100000",
  21993=>"000000000",
  21994=>"110110100",
  21995=>"111111000",
  21996=>"111111111",
  21997=>"111010000",
  21998=>"000000000",
  21999=>"000111110",
  22000=>"000000011",
  22001=>"011001111",
  22002=>"010111111",
  22003=>"111100110",
  22004=>"100111011",
  22005=>"101100100",
  22006=>"000100111",
  22007=>"000100100",
  22008=>"111001101",
  22009=>"101000110",
  22010=>"111111111",
  22011=>"111000011",
  22012=>"011111000",
  22013=>"000000000",
  22014=>"100111011",
  22015=>"000000101",
  22016=>"001111011",
  22017=>"011000011",
  22018=>"100000000",
  22019=>"111010000",
  22020=>"000111100",
  22021=>"101001000",
  22022=>"111001000",
  22023=>"100000101",
  22024=>"000010010",
  22025=>"000000101",
  22026=>"000000101",
  22027=>"010111000",
  22028=>"000010111",
  22029=>"000111111",
  22030=>"100100100",
  22031=>"110100010",
  22032=>"110010000",
  22033=>"100000001",
  22034=>"111000100",
  22035=>"001000101",
  22036=>"111110101",
  22037=>"100100101",
  22038=>"011010110",
  22039=>"000000000",
  22040=>"001000001",
  22041=>"000100010",
  22042=>"010111110",
  22043=>"000011111",
  22044=>"110001111",
  22045=>"000000100",
  22046=>"000100000",
  22047=>"000111010",
  22048=>"111111110",
  22049=>"011111000",
  22050=>"000110111",
  22051=>"011000000",
  22052=>"001111111",
  22053=>"000010011",
  22054=>"000110111",
  22055=>"101000000",
  22056=>"110110000",
  22057=>"000101001",
  22058=>"111111101",
  22059=>"001000000",
  22060=>"100100000",
  22061=>"111000101",
  22062=>"111010100",
  22063=>"000101101",
  22064=>"000101011",
  22065=>"000001101",
  22066=>"010011010",
  22067=>"111101000",
  22068=>"001001000",
  22069=>"001010110",
  22070=>"100000101",
  22071=>"010010100",
  22072=>"111001111",
  22073=>"001001101",
  22074=>"011000000",
  22075=>"101101001",
  22076=>"010011111",
  22077=>"111011000",
  22078=>"000000000",
  22079=>"011011001",
  22080=>"000111111",
  22081=>"000001110",
  22082=>"101000000",
  22083=>"001100011",
  22084=>"011010011",
  22085=>"011000000",
  22086=>"101101101",
  22087=>"110110000",
  22088=>"100001101",
  22089=>"100000100",
  22090=>"000000000",
  22091=>"111010000",
  22092=>"111000110",
  22093=>"101111110",
  22094=>"001110011",
  22095=>"010000101",
  22096=>"101100000",
  22097=>"011011000",
  22098=>"110001111",
  22099=>"011001001",
  22100=>"010000110",
  22101=>"111100000",
  22102=>"001101011",
  22103=>"101000101",
  22104=>"001101111",
  22105=>"000100110",
  22106=>"000001111",
  22107=>"010011011",
  22108=>"000110110",
  22109=>"000001000",
  22110=>"111011000",
  22111=>"100111010",
  22112=>"001101111",
  22113=>"110111101",
  22114=>"101000101",
  22115=>"111100111",
  22116=>"011111100",
  22117=>"001101000",
  22118=>"000001000",
  22119=>"000010001",
  22120=>"111110110",
  22121=>"111100101",
  22122=>"110111000",
  22123=>"111000010",
  22124=>"000110110",
  22125=>"001001000",
  22126=>"000000011",
  22127=>"110000000",
  22128=>"100110100",
  22129=>"000000111",
  22130=>"001001101",
  22131=>"000010111",
  22132=>"111100000",
  22133=>"111101000",
  22134=>"011101000",
  22135=>"000111111",
  22136=>"000000111",
  22137=>"111011111",
  22138=>"000110011",
  22139=>"000111110",
  22140=>"001001001",
  22141=>"011101000",
  22142=>"000100000",
  22143=>"000110000",
  22144=>"000111111",
  22145=>"111000000",
  22146=>"000011111",
  22147=>"000000000",
  22148=>"111001101",
  22149=>"111001000",
  22150=>"000000000",
  22151=>"000011011",
  22152=>"000111110",
  22153=>"000000010",
  22154=>"000000100",
  22155=>"111010000",
  22156=>"010111010",
  22157=>"101111110",
  22158=>"010110111",
  22159=>"000000110",
  22160=>"101111111",
  22161=>"000111111",
  22162=>"000001000",
  22163=>"111001000",
  22164=>"110101010",
  22165=>"101001111",
  22166=>"111101111",
  22167=>"000011010",
  22168=>"111000000",
  22169=>"000000000",
  22170=>"000111011",
  22171=>"111001000",
  22172=>"111101111",
  22173=>"000000000",
  22174=>"010111000",
  22175=>"111000000",
  22176=>"011111111",
  22177=>"110110111",
  22178=>"000111110",
  22179=>"000100111",
  22180=>"110011100",
  22181=>"100110111",
  22182=>"110110000",
  22183=>"001001100",
  22184=>"101000000",
  22185=>"011111010",
  22186=>"001101111",
  22187=>"101000011",
  22188=>"101110010",
  22189=>"101001101",
  22190=>"111111000",
  22191=>"110110000",
  22192=>"000110100",
  22193=>"001011111",
  22194=>"111000010",
  22195=>"001101010",
  22196=>"011011000",
  22197=>"111111110",
  22198=>"000010100",
  22199=>"001010010",
  22200=>"001011111",
  22201=>"000000000",
  22202=>"000110001",
  22203=>"010010010",
  22204=>"100000000",
  22205=>"101111010",
  22206=>"010011010",
  22207=>"111111101",
  22208=>"101000000",
  22209=>"101001101",
  22210=>"101101111",
  22211=>"001011011",
  22212=>"011001001",
  22213=>"110110001",
  22214=>"000100100",
  22215=>"001001101",
  22216=>"001001000",
  22217=>"000110110",
  22218=>"101100111",
  22219=>"100111010",
  22220=>"010111110",
  22221=>"100100000",
  22222=>"000110000",
  22223=>"100111000",
  22224=>"001001001",
  22225=>"000111111",
  22226=>"000000100",
  22227=>"001001010",
  22228=>"111100000",
  22229=>"000100100",
  22230=>"101001111",
  22231=>"101101110",
  22232=>"110000000",
  22233=>"010010111",
  22234=>"001101111",
  22235=>"101000010",
  22236=>"001111001",
  22237=>"000000100",
  22238=>"110000110",
  22239=>"110001101",
  22240=>"000010110",
  22241=>"111101001",
  22242=>"111000000",
  22243=>"001111111",
  22244=>"000000001",
  22245=>"010111100",
  22246=>"111010010",
  22247=>"010110111",
  22248=>"111101000",
  22249=>"110111101",
  22250=>"000000000",
  22251=>"000111001",
  22252=>"000010101",
  22253=>"010110111",
  22254=>"101000000",
  22255=>"000111100",
  22256=>"110010000",
  22257=>"111011001",
  22258=>"111001000",
  22259=>"101000011",
  22260=>"110101100",
  22261=>"101011001",
  22262=>"000000111",
  22263=>"000110000",
  22264=>"111000000",
  22265=>"111001011",
  22266=>"010000110",
  22267=>"111111101",
  22268=>"111000100",
  22269=>"010010010",
  22270=>"000111011",
  22271=>"111001101",
  22272=>"010001001",
  22273=>"000000000",
  22274=>"010110010",
  22275=>"000000000",
  22276=>"000101001",
  22277=>"000000010",
  22278=>"010010000",
  22279=>"000001010",
  22280=>"111110110",
  22281=>"000000000",
  22282=>"001111111",
  22283=>"101010000",
  22284=>"111000100",
  22285=>"011011001",
  22286=>"101000011",
  22287=>"111000111",
  22288=>"001000000",
  22289=>"000000001",
  22290=>"100000110",
  22291=>"000000010",
  22292=>"000000001",
  22293=>"000000000",
  22294=>"001011010",
  22295=>"000000100",
  22296=>"000000001",
  22297=>"000001001",
  22298=>"010111111",
  22299=>"011111011",
  22300=>"011111111",
  22301=>"111110010",
  22302=>"000000000",
  22303=>"111101110",
  22304=>"000101011",
  22305=>"000101001",
  22306=>"110000111",
  22307=>"110000111",
  22308=>"011111011",
  22309=>"010000010",
  22310=>"000000100",
  22311=>"001111011",
  22312=>"111111111",
  22313=>"111111010",
  22314=>"001000001",
  22315=>"101101000",
  22316=>"111111001",
  22317=>"000000000",
  22318=>"110000010",
  22319=>"011000000",
  22320=>"000000000",
  22321=>"111111111",
  22322=>"111111010",
  22323=>"000000000",
  22324=>"000010000",
  22325=>"001111000",
  22326=>"000100100",
  22327=>"001000000",
  22328=>"000000000",
  22329=>"100000000",
  22330=>"100101111",
  22331=>"111110111",
  22332=>"100000000",
  22333=>"111111111",
  22334=>"000000010",
  22335=>"000011110",
  22336=>"001001000",
  22337=>"111111111",
  22338=>"111101001",
  22339=>"000111011",
  22340=>"111111000",
  22341=>"000000000",
  22342=>"010000000",
  22343=>"110111100",
  22344=>"000000000",
  22345=>"101111011",
  22346=>"111111001",
  22347=>"001111001",
  22348=>"000000011",
  22349=>"111111110",
  22350=>"111111111",
  22351=>"111111011",
  22352=>"000110111",
  22353=>"000010010",
  22354=>"000000000",
  22355=>"011001000",
  22356=>"010110110",
  22357=>"000000000",
  22358=>"111111111",
  22359=>"000000000",
  22360=>"111111010",
  22361=>"000111111",
  22362=>"101100101",
  22363=>"000100111",
  22364=>"111000000",
  22365=>"001000011",
  22366=>"011010110",
  22367=>"101111000",
  22368=>"010111111",
  22369=>"101111000",
  22370=>"101111000",
  22371=>"100101111",
  22372=>"110110110",
  22373=>"111111011",
  22374=>"101111111",
  22375=>"110111111",
  22376=>"010000000",
  22377=>"000000000",
  22378=>"000000000",
  22379=>"111111110",
  22380=>"110111111",
  22381=>"111111111",
  22382=>"001000000",
  22383=>"000000010",
  22384=>"000110011",
  22385=>"000000000",
  22386=>"000010010",
  22387=>"111111111",
  22388=>"000000000",
  22389=>"000000001",
  22390=>"000000000",
  22391=>"111111111",
  22392=>"010000111",
  22393=>"010000000",
  22394=>"001000001",
  22395=>"100100100",
  22396=>"000100010",
  22397=>"100100000",
  22398=>"010000000",
  22399=>"110111111",
  22400=>"000001111",
  22401=>"000100000",
  22402=>"000010010",
  22403=>"111110111",
  22404=>"000100101",
  22405=>"000100101",
  22406=>"011010111",
  22407=>"011001000",
  22408=>"001111111",
  22409=>"101111111",
  22410=>"101011111",
  22411=>"110000000",
  22412=>"111111000",
  22413=>"000000001",
  22414=>"010110110",
  22415=>"101000000",
  22416=>"100101111",
  22417=>"111111111",
  22418=>"000000000",
  22419=>"011010000",
  22420=>"111111111",
  22421=>"000000000",
  22422=>"111111111",
  22423=>"001000011",
  22424=>"010010100",
  22425=>"000001110",
  22426=>"001001011",
  22427=>"000010010",
  22428=>"000010010",
  22429=>"100111101",
  22430=>"000000000",
  22431=>"000001000",
  22432=>"001111101",
  22433=>"001000000",
  22434=>"111111111",
  22435=>"111000100",
  22436=>"000000000",
  22437=>"110110110",
  22438=>"111010000",
  22439=>"111111011",
  22440=>"000000101",
  22441=>"000000010",
  22442=>"111111110",
  22443=>"000101111",
  22444=>"111000100",
  22445=>"110110010",
  22446=>"110101111",
  22447=>"010010110",
  22448=>"010010010",
  22449=>"101001001",
  22450=>"111100000",
  22451=>"000000110",
  22452=>"111111111",
  22453=>"111110101",
  22454=>"000000000",
  22455=>"010010010",
  22456=>"011000000",
  22457=>"111110100",
  22458=>"110111110",
  22459=>"000110010",
  22460=>"001110110",
  22461=>"101111000",
  22462=>"011011011",
  22463=>"010000000",
  22464=>"010000000",
  22465=>"000010100",
  22466=>"000000010",
  22467=>"111111100",
  22468=>"010010011",
  22469=>"100001101",
  22470=>"000000000",
  22471=>"111111011",
  22472=>"111101111",
  22473=>"011001111",
  22474=>"111000000",
  22475=>"000100111",
  22476=>"001110000",
  22477=>"000000000",
  22478=>"000000000",
  22479=>"000000000",
  22480=>"000000010",
  22481=>"111111110",
  22482=>"110111111",
  22483=>"110100110",
  22484=>"010000000",
  22485=>"100000000",
  22486=>"010100100",
  22487=>"000000000",
  22488=>"111110110",
  22489=>"000000111",
  22490=>"110111111",
  22491=>"000000000",
  22492=>"000000000",
  22493=>"000000010",
  22494=>"010010001",
  22495=>"000000000",
  22496=>"011000001",
  22497=>"000111000",
  22498=>"111010110",
  22499=>"101101111",
  22500=>"001000001",
  22501=>"101111000",
  22502=>"100110000",
  22503=>"111111101",
  22504=>"000000000",
  22505=>"110111111",
  22506=>"101111110",
  22507=>"000010000",
  22508=>"000000010",
  22509=>"001001100",
  22510=>"010010010",
  22511=>"111010110",
  22512=>"010000010",
  22513=>"111000011",
  22514=>"000001100",
  22515=>"101001100",
  22516=>"110000000",
  22517=>"111111111",
  22518=>"000000010",
  22519=>"000000000",
  22520=>"000000000",
  22521=>"000000010",
  22522=>"011011000",
  22523=>"111011111",
  22524=>"111101111",
  22525=>"110000111",
  22526=>"111111101",
  22527=>"000000111",
  22528=>"001001000",
  22529=>"111101101",
  22530=>"011000111",
  22531=>"001000000",
  22532=>"000110110",
  22533=>"000100011",
  22534=>"111101101",
  22535=>"110111011",
  22536=>"000111010",
  22537=>"101100000",
  22538=>"000000000",
  22539=>"111101000",
  22540=>"001111011",
  22541=>"101000000",
  22542=>"000001100",
  22543=>"010110000",
  22544=>"011000010",
  22545=>"100000010",
  22546=>"011000100",
  22547=>"011011000",
  22548=>"111001001",
  22549=>"101100100",
  22550=>"110111001",
  22551=>"111101011",
  22552=>"101000000",
  22553=>"000001110",
  22554=>"010010000",
  22555=>"011000100",
  22556=>"000111011",
  22557=>"000100100",
  22558=>"101101111",
  22559=>"001111010",
  22560=>"000000000",
  22561=>"011101111",
  22562=>"100111000",
  22563=>"000011111",
  22564=>"000100110",
  22565=>"110100111",
  22566=>"111111111",
  22567=>"101011000",
  22568=>"111100111",
  22569=>"111101101",
  22570=>"101100100",
  22571=>"010100100",
  22572=>"101101111",
  22573=>"000110111",
  22574=>"100000110",
  22575=>"110111011",
  22576=>"000111111",
  22577=>"001111111",
  22578=>"001011011",
  22579=>"110111100",
  22580=>"000000000",
  22581=>"111111010",
  22582=>"110100100",
  22583=>"000000010",
  22584=>"010010000",
  22585=>"101100101",
  22586=>"001111111",
  22587=>"110011010",
  22588=>"101111011",
  22589=>"011111010",
  22590=>"100000100",
  22591=>"100111111",
  22592=>"111111111",
  22593=>"010000001",
  22594=>"000000010",
  22595=>"001000110",
  22596=>"111111010",
  22597=>"111111101",
  22598=>"000000000",
  22599=>"111011100",
  22600=>"000010111",
  22601=>"000000010",
  22602=>"111101101",
  22603=>"111000001",
  22604=>"111101101",
  22605=>"000010010",
  22606=>"000001111",
  22607=>"011111111",
  22608=>"001001001",
  22609=>"111000111",
  22610=>"111101101",
  22611=>"111101101",
  22612=>"101100100",
  22613=>"000000010",
  22614=>"101111010",
  22615=>"110100100",
  22616=>"111000000",
  22617=>"101100101",
  22618=>"100110111",
  22619=>"000000000",
  22620=>"000010111",
  22621=>"000000000",
  22622=>"111000010",
  22623=>"100000111",
  22624=>"111010011",
  22625=>"110101010",
  22626=>"000000010",
  22627=>"001001000",
  22628=>"100100010",
  22629=>"000100100",
  22630=>"111111111",
  22631=>"011011001",
  22632=>"111110010",
  22633=>"000000000",
  22634=>"000010011",
  22635=>"100011111",
  22636=>"000010101",
  22637=>"000000111",
  22638=>"010111011",
  22639=>"111101111",
  22640=>"111111101",
  22641=>"000000111",
  22642=>"111001000",
  22643=>"000011000",
  22644=>"000000000",
  22645=>"001100101",
  22646=>"010010111",
  22647=>"111100101",
  22648=>"010000000",
  22649=>"011010000",
  22650=>"100100000",
  22651=>"000101010",
  22652=>"010100111",
  22653=>"100100100",
  22654=>"101000011",
  22655=>"101000100",
  22656=>"111101000",
  22657=>"000000011",
  22658=>"000000011",
  22659=>"011111101",
  22660=>"111100100",
  22661=>"111111101",
  22662=>"001111111",
  22663=>"001001000",
  22664=>"001110100",
  22665=>"001000101",
  22666=>"111000101",
  22667=>"111111001",
  22668=>"000100000",
  22669=>"101000000",
  22670=>"000010001",
  22671=>"111100110",
  22672=>"100100100",
  22673=>"010011011",
  22674=>"001000010",
  22675=>"000101000",
  22676=>"000001010",
  22677=>"011100101",
  22678=>"001111011",
  22679=>"001001011",
  22680=>"000011111",
  22681=>"000010000",
  22682=>"110000001",
  22683=>"111100101",
  22684=>"011101100",
  22685=>"100001000",
  22686=>"010010110",
  22687=>"000010101",
  22688=>"000001001",
  22689=>"111101000",
  22690=>"000011010",
  22691=>"100101101",
  22692=>"010111101",
  22693=>"010101100",
  22694=>"010111000",
  22695=>"001000001",
  22696=>"111010000",
  22697=>"010010000",
  22698=>"111001011",
  22699=>"111100000",
  22700=>"110010000",
  22701=>"101101100",
  22702=>"101100001",
  22703=>"000100110",
  22704=>"010100010",
  22705=>"000000011",
  22706=>"011100100",
  22707=>"001000000",
  22708=>"000001010",
  22709=>"111111000",
  22710=>"011100100",
  22711=>"000011000",
  22712=>"000000010",
  22713=>"100010010",
  22714=>"111011001",
  22715=>"110011000",
  22716=>"000001011",
  22717=>"000000011",
  22718=>"100000100",
  22719=>"110000010",
  22720=>"011000000",
  22721=>"111000100",
  22722=>"010100011",
  22723=>"001100011",
  22724=>"101111010",
  22725=>"110000110",
  22726=>"111111010",
  22727=>"100100111",
  22728=>"000000101",
  22729=>"111101000",
  22730=>"000001100",
  22731=>"000011011",
  22732=>"011000110",
  22733=>"110111111",
  22734=>"101011000",
  22735=>"110111010",
  22736=>"010100111",
  22737=>"000110110",
  22738=>"010101110",
  22739=>"000101000",
  22740=>"010010010",
  22741=>"000000111",
  22742=>"011010111",
  22743=>"000000011",
  22744=>"011011011",
  22745=>"110000000",
  22746=>"111110110",
  22747=>"100000100",
  22748=>"101001001",
  22749=>"110000000",
  22750=>"011111000",
  22751=>"000000000",
  22752=>"111100000",
  22753=>"101100000",
  22754=>"010101100",
  22755=>"100000000",
  22756=>"111100101",
  22757=>"111111101",
  22758=>"000000000",
  22759=>"101111110",
  22760=>"000101011",
  22761=>"010010000",
  22762=>"000000000",
  22763=>"100000111",
  22764=>"111100000",
  22765=>"000101110",
  22766=>"000000001",
  22767=>"000011010",
  22768=>"000110010",
  22769=>"001000001",
  22770=>"111101101",
  22771=>"001101100",
  22772=>"111100100",
  22773=>"101000000",
  22774=>"000000010",
  22775=>"110000100",
  22776=>"011111111",
  22777=>"010100011",
  22778=>"000000000",
  22779=>"101100010",
  22780=>"000011011",
  22781=>"000011011",
  22782=>"000011011",
  22783=>"101001101",
  22784=>"000100100",
  22785=>"001000000",
  22786=>"110111010",
  22787=>"000000000",
  22788=>"001000101",
  22789=>"101101001",
  22790=>"111100101",
  22791=>"000000000",
  22792=>"000001000",
  22793=>"111111101",
  22794=>"111111111",
  22795=>"000000000",
  22796=>"111110110",
  22797=>"000100111",
  22798=>"000000000",
  22799=>"111111111",
  22800=>"010010000",
  22801=>"000000000",
  22802=>"111000000",
  22803=>"000000000",
  22804=>"111111111",
  22805=>"110110111",
  22806=>"010100101",
  22807=>"111111101",
  22808=>"000111111",
  22809=>"100010000",
  22810=>"111000111",
  22811=>"111111111",
  22812=>"111111111",
  22813=>"111001111",
  22814=>"000001111",
  22815=>"100100100",
  22816=>"111101111",
  22817=>"111101111",
  22818=>"111110000",
  22819=>"111111110",
  22820=>"000000100",
  22821=>"000000001",
  22822=>"110111110",
  22823=>"000000111",
  22824=>"111111001",
  22825=>"000000101",
  22826=>"000000101",
  22827=>"100110000",
  22828=>"000000000",
  22829=>"000110111",
  22830=>"000000000",
  22831=>"101110001",
  22832=>"000000000",
  22833=>"001101100",
  22834=>"011011011",
  22835=>"000000000",
  22836=>"100000100",
  22837=>"111111111",
  22838=>"111111111",
  22839=>"000000111",
  22840=>"101101000",
  22841=>"000011001",
  22842=>"011000101",
  22843=>"000000000",
  22844=>"000000000",
  22845=>"111111101",
  22846=>"111111111",
  22847=>"000000000",
  22848=>"010010001",
  22849=>"000000001",
  22850=>"111101001",
  22851=>"110111111",
  22852=>"111100111",
  22853=>"000000101",
  22854=>"001000101",
  22855=>"001000111",
  22856=>"010111111",
  22857=>"111111101",
  22858=>"000000001",
  22859=>"110111111",
  22860=>"000000000",
  22861=>"100000011",
  22862=>"011000001",
  22863=>"000011111",
  22864=>"111111111",
  22865=>"111111111",
  22866=>"000001000",
  22867=>"000000110",
  22868=>"110111000",
  22869=>"000000000",
  22870=>"000000000",
  22871=>"111111111",
  22872=>"001001100",
  22873=>"000000000",
  22874=>"000000000",
  22875=>"000000000",
  22876=>"000000100",
  22877=>"100000100",
  22878=>"111111110",
  22879=>"000100001",
  22880=>"000000000",
  22881=>"000000100",
  22882=>"111111100",
  22883=>"000000000",
  22884=>"001001001",
  22885=>"001010000",
  22886=>"000000111",
  22887=>"011101101",
  22888=>"000000000",
  22889=>"000000000",
  22890=>"000000111",
  22891=>"011110111",
  22892=>"000000001",
  22893=>"111111111",
  22894=>"111110000",
  22895=>"000000000",
  22896=>"000000000",
  22897=>"000000001",
  22898=>"111001001",
  22899=>"101011100",
  22900=>"000000101",
  22901=>"010010000",
  22902=>"000000001",
  22903=>"011111011",
  22904=>"111100111",
  22905=>"001000000",
  22906=>"000000101",
  22907=>"111111111",
  22908=>"000111000",
  22909=>"000000001",
  22910=>"111111111",
  22911=>"111111010",
  22912=>"000000000",
  22913=>"111111111",
  22914=>"000000000",
  22915=>"001000101",
  22916=>"100000101",
  22917=>"000111011",
  22918=>"000000010",
  22919=>"000000000",
  22920=>"000000001",
  22921=>"000000111",
  22922=>"000001001",
  22923=>"000000000",
  22924=>"111111110",
  22925=>"111101101",
  22926=>"111111011",
  22927=>"000011000",
  22928=>"000000100",
  22929=>"000000000",
  22930=>"001000000",
  22931=>"000000101",
  22932=>"000000000",
  22933=>"111111000",
  22934=>"110100100",
  22935=>"000000001",
  22936=>"000100001",
  22937=>"000010001",
  22938=>"111111110",
  22939=>"000101100",
  22940=>"000110111",
  22941=>"100110111",
  22942=>"010001110",
  22943=>"111111001",
  22944=>"111111010",
  22945=>"000000000",
  22946=>"001000101",
  22947=>"111011111",
  22948=>"001010101",
  22949=>"000000100",
  22950=>"000000100",
  22951=>"111111111",
  22952=>"000000000",
  22953=>"000001111",
  22954=>"111111111",
  22955=>"110000000",
  22956=>"001001111",
  22957=>"000000000",
  22958=>"111101101",
  22959=>"100111110",
  22960=>"000101001",
  22961=>"000000010",
  22962=>"111000111",
  22963=>"010000000",
  22964=>"000000001",
  22965=>"111101111",
  22966=>"000000000",
  22967=>"000000000",
  22968=>"000000000",
  22969=>"000000001",
  22970=>"000000000",
  22971=>"000000000",
  22972=>"000101111",
  22973=>"111110110",
  22974=>"000000000",
  22975=>"111011101",
  22976=>"110111111",
  22977=>"111111111",
  22978=>"000000010",
  22979=>"101100101",
  22980=>"000110010",
  22981=>"010010111",
  22982=>"001000000",
  22983=>"111111111",
  22984=>"000000001",
  22985=>"111110000",
  22986=>"000000010",
  22987=>"100111000",
  22988=>"000010110",
  22989=>"000010000",
  22990=>"111000000",
  22991=>"000001101",
  22992=>"110000000",
  22993=>"000000000",
  22994=>"001000000",
  22995=>"111110100",
  22996=>"000100000",
  22997=>"000000001",
  22998=>"111111110",
  22999=>"001000000",
  23000=>"111111111",
  23001=>"101110110",
  23002=>"001011011",
  23003=>"111110000",
  23004=>"000000001",
  23005=>"100000111",
  23006=>"111111111",
  23007=>"010000010",
  23008=>"111111010",
  23009=>"000101111",
  23010=>"111111111",
  23011=>"000000000",
  23012=>"000011000",
  23013=>"110110111",
  23014=>"000000000",
  23015=>"000001000",
  23016=>"010000101",
  23017=>"111111000",
  23018=>"101111111",
  23019=>"111101111",
  23020=>"111111000",
  23021=>"111111000",
  23022=>"110111000",
  23023=>"111101101",
  23024=>"111110000",
  23025=>"100100111",
  23026=>"001101111",
  23027=>"000000000",
  23028=>"000001011",
  23029=>"110110111",
  23030=>"101111111",
  23031=>"001001101",
  23032=>"111111111",
  23033=>"000001000",
  23034=>"111100101",
  23035=>"000000000",
  23036=>"111000111",
  23037=>"111000111",
  23038=>"000000100",
  23039=>"110111000",
  23040=>"110111011",
  23041=>"000000000",
  23042=>"000110111",
  23043=>"001000100",
  23044=>"001010010",
  23045=>"101000000",
  23046=>"111011110",
  23047=>"000000000",
  23048=>"000011010",
  23049=>"000110110",
  23050=>"001011011",
  23051=>"101100111",
  23052=>"100000101",
  23053=>"001100110",
  23054=>"000100110",
  23055=>"111011011",
  23056=>"111111001",
  23057=>"000000111",
  23058=>"111011100",
  23059=>"000000000",
  23060=>"111011001",
  23061=>"000111111",
  23062=>"111001100",
  23063=>"111111110",
  23064=>"101001110",
  23065=>"010000000",
  23066=>"001101011",
  23067=>"000000101",
  23068=>"000000000",
  23069=>"111000000",
  23070=>"010111111",
  23071=>"000000000",
  23072=>"000011000",
  23073=>"100111111",
  23074=>"110101101",
  23075=>"000101101",
  23076=>"111011001",
  23077=>"001011000",
  23078=>"000010010",
  23079=>"001101111",
  23080=>"011111111",
  23081=>"001010010",
  23082=>"101100110",
  23083=>"110000000",
  23084=>"000100011",
  23085=>"111011100",
  23086=>"111101110",
  23087=>"000111000",
  23088=>"001001000",
  23089=>"011100101",
  23090=>"001101101",
  23091=>"000000000",
  23092=>"000010010",
  23093=>"110111110",
  23094=>"011111110",
  23095=>"010010010",
  23096=>"111111100",
  23097=>"000010000",
  23098=>"000001100",
  23099=>"000000000",
  23100=>"001000000",
  23101=>"100111111",
  23102=>"110000010",
  23103=>"000001100",
  23104=>"111111000",
  23105=>"010001001",
  23106=>"101111111",
  23107=>"001000000",
  23108=>"111110000",
  23109=>"000100111",
  23110=>"000111111",
  23111=>"111111111",
  23112=>"101110000",
  23113=>"011001101",
  23114=>"000000111",
  23115=>"010010010",
  23116=>"111111010",
  23117=>"010100010",
  23118=>"011011111",
  23119=>"000000011",
  23120=>"000011111",
  23121=>"100111011",
  23122=>"000000110",
  23123=>"111100000",
  23124=>"000000001",
  23125=>"111111111",
  23126=>"000101110",
  23127=>"000000010",
  23128=>"111101100",
  23129=>"000110000",
  23130=>"000001101",
  23131=>"111110000",
  23132=>"000110000",
  23133=>"110101000",
  23134=>"101000000",
  23135=>"000000100",
  23136=>"010110010",
  23137=>"000000000",
  23138=>"011011011",
  23139=>"111111111",
  23140=>"000000100",
  23141=>"000000000",
  23142=>"000100111",
  23143=>"000000111",
  23144=>"100000000",
  23145=>"111111101",
  23146=>"010111111",
  23147=>"000000100",
  23148=>"100000111",
  23149=>"101000101",
  23150=>"000000000",
  23151=>"000000101",
  23152=>"011001011",
  23153=>"010000101",
  23154=>"111111011",
  23155=>"001001001",
  23156=>"111111111",
  23157=>"000000000",
  23158=>"001000000",
  23159=>"010111011",
  23160=>"101100111",
  23161=>"111100000",
  23162=>"111100100",
  23163=>"111000100",
  23164=>"000111111",
  23165=>"111100000",
  23166=>"101111011",
  23167=>"000100000",
  23168=>"111001000",
  23169=>"000000000",
  23170=>"101010000",
  23171=>"111111111",
  23172=>"000000000",
  23173=>"111101000",
  23174=>"101110000",
  23175=>"000100000",
  23176=>"000000000",
  23177=>"000010000",
  23178=>"000101111",
  23179=>"111101101",
  23180=>"010000000",
  23181=>"101101100",
  23182=>"111010000",
  23183=>"000010010",
  23184=>"001001001",
  23185=>"000000000",
  23186=>"000000000",
  23187=>"000000101",
  23188=>"100000000",
  23189=>"000010010",
  23190=>"111111100",
  23191=>"000100001",
  23192=>"001000000",
  23193=>"000001000",
  23194=>"010010010",
  23195=>"111100011",
  23196=>"000000111",
  23197=>"010110110",
  23198=>"001111111",
  23199=>"000010000",
  23200=>"101110000",
  23201=>"000111111",
  23202=>"101000000",
  23203=>"111111010",
  23204=>"011000000",
  23205=>"011011011",
  23206=>"111110100",
  23207=>"001111111",
  23208=>"001000101",
  23209=>"000000101",
  23210=>"011001101",
  23211=>"000001000",
  23212=>"111100000",
  23213=>"000000111",
  23214=>"001111111",
  23215=>"100100101",
  23216=>"110000001",
  23217=>"000001001",
  23218=>"111000000",
  23219=>"000001100",
  23220=>"101100111",
  23221=>"101010000",
  23222=>"010111111",
  23223=>"100101101",
  23224=>"000000000",
  23225=>"000000000",
  23226=>"000011111",
  23227=>"111100111",
  23228=>"000000101",
  23229=>"111011011",
  23230=>"110110000",
  23231=>"011011111",
  23232=>"001010010",
  23233=>"000000000",
  23234=>"111011111",
  23235=>"100000010",
  23236=>"110101101",
  23237=>"111111111",
  23238=>"010000011",
  23239=>"111001000",
  23240=>"111101111",
  23241=>"000000000",
  23242=>"111111101",
  23243=>"001000000",
  23244=>"000001000",
  23245=>"000000111",
  23246=>"010111010",
  23247=>"110010101",
  23248=>"000000000",
  23249=>"011011001",
  23250=>"110000101",
  23251=>"111111111",
  23252=>"000001111",
  23253=>"000110100",
  23254=>"000111011",
  23255=>"000111001",
  23256=>"111101111",
  23257=>"000000111",
  23258=>"101001000",
  23259=>"101000101",
  23260=>"111111001",
  23261=>"100101111",
  23262=>"010111011",
  23263=>"111010111",
  23264=>"000000111",
  23265=>"111000110",
  23266=>"110101001",
  23267=>"001011000",
  23268=>"000000000",
  23269=>"101111101",
  23270=>"100000000",
  23271=>"100110110",
  23272=>"000101111",
  23273=>"000100000",
  23274=>"110110010",
  23275=>"011101111",
  23276=>"000000111",
  23277=>"110111111",
  23278=>"000000000",
  23279=>"110000000",
  23280=>"000000000",
  23281=>"011111110",
  23282=>"111001101",
  23283=>"001011000",
  23284=>"101111011",
  23285=>"101001000",
  23286=>"001000011",
  23287=>"110000011",
  23288=>"111111000",
  23289=>"111111111",
  23290=>"100000000",
  23291=>"000000110",
  23292=>"111111000",
  23293=>"101000000",
  23294=>"110111011",
  23295=>"101000010",
  23296=>"100000010",
  23297=>"000000000",
  23298=>"100000100",
  23299=>"011011111",
  23300=>"110001001",
  23301=>"101000011",
  23302=>"110001010",
  23303=>"000111000",
  23304=>"100010000",
  23305=>"110000010",
  23306=>"010001011",
  23307=>"010000100",
  23308=>"110100000",
  23309=>"011011000",
  23310=>"010000000",
  23311=>"000001000",
  23312=>"000100000",
  23313=>"000101111",
  23314=>"101100001",
  23315=>"111100110",
  23316=>"100000000",
  23317=>"001011111",
  23318=>"111011001",
  23319=>"111101011",
  23320=>"000001110",
  23321=>"111110110",
  23322=>"001000000",
  23323=>"111111110",
  23324=>"110000000",
  23325=>"001000000",
  23326=>"111000000",
  23327=>"000100000",
  23328=>"001011110",
  23329=>"001111100",
  23330=>"000110101",
  23331=>"011011011",
  23332=>"110111110",
  23333=>"111100100",
  23334=>"000011110",
  23335=>"111110001",
  23336=>"110111100",
  23337=>"110110011",
  23338=>"100100100",
  23339=>"110001010",
  23340=>"110110110",
  23341=>"000000000",
  23342=>"110100110",
  23343=>"111100101",
  23344=>"111100110",
  23345=>"110100010",
  23346=>"000000000",
  23347=>"111000000",
  23348=>"010001110",
  23349=>"000111011",
  23350=>"111100000",
  23351=>"011111110",
  23352=>"100000011",
  23353=>"001001000",
  23354=>"000100010",
  23355=>"111111111",
  23356=>"111111111",
  23357=>"010110001",
  23358=>"000001001",
  23359=>"001001011",
  23360=>"110001000",
  23361=>"110101010",
  23362=>"110111111",
  23363=>"000011011",
  23364=>"111111111",
  23365=>"000101100",
  23366=>"010010011",
  23367=>"101011111",
  23368=>"000001011",
  23369=>"011011010",
  23370=>"000000000",
  23371=>"010001100",
  23372=>"100100010",
  23373=>"011111111",
  23374=>"001111000",
  23375=>"001000001",
  23376=>"011110100",
  23377=>"111100101",
  23378=>"110000000",
  23379=>"000000011",
  23380=>"111011000",
  23381=>"011100001",
  23382=>"110111110",
  23383=>"001010001",
  23384=>"110110111",
  23385=>"110110100",
  23386=>"001110110",
  23387=>"100111100",
  23388=>"100110001",
  23389=>"000000000",
  23390=>"111111111",
  23391=>"010011101",
  23392=>"011000001",
  23393=>"000010001",
  23394=>"110110010",
  23395=>"000110100",
  23396=>"000111100",
  23397=>"111100010",
  23398=>"111010010",
  23399=>"000010110",
  23400=>"000000010",
  23401=>"011101001",
  23402=>"010110110",
  23403=>"000001001",
  23404=>"100001111",
  23405=>"000001001",
  23406=>"011011011",
  23407=>"000000000",
  23408=>"110110110",
  23409=>"000101111",
  23410=>"000000111",
  23411=>"100100100",
  23412=>"011000011",
  23413=>"100100110",
  23414=>"001010010",
  23415=>"111110000",
  23416=>"000111111",
  23417=>"010010100",
  23418=>"000100100",
  23419=>"101001101",
  23420=>"001111111",
  23421=>"110100001",
  23422=>"110100100",
  23423=>"011111001",
  23424=>"111001000",
  23425=>"110100100",
  23426=>"111001011",
  23427=>"000000011",
  23428=>"001101001",
  23429=>"101011101",
  23430=>"000000000",
  23431=>"000000000",
  23432=>"110001001",
  23433=>"000001101",
  23434=>"100110101",
  23435=>"101001100",
  23436=>"100011111",
  23437=>"001001011",
  23438=>"111111111",
  23439=>"101000100",
  23440=>"010100000",
  23441=>"100100000",
  23442=>"100011010",
  23443=>"000100000",
  23444=>"000010000",
  23445=>"000000001",
  23446=>"011010110",
  23447=>"100000000",
  23448=>"011000101",
  23449=>"101010010",
  23450=>"011111110",
  23451=>"000100110",
  23452=>"111100001",
  23453=>"000111111",
  23454=>"010011001",
  23455=>"100101101",
  23456=>"100001000",
  23457=>"110110001",
  23458=>"011011000",
  23459=>"010010100",
  23460=>"011000010",
  23461=>"011111111",
  23462=>"111111010",
  23463=>"111011001",
  23464=>"011000000",
  23465=>"000000110",
  23466=>"001000000",
  23467=>"101101000",
  23468=>"011111110",
  23469=>"010011010",
  23470=>"111100000",
  23471=>"001010110",
  23472=>"000010000",
  23473=>"111111001",
  23474=>"011100000",
  23475=>"000001111",
  23476=>"001011111",
  23477=>"000010010",
  23478=>"110000011",
  23479=>"000000000",
  23480=>"000000000",
  23481=>"111111111",
  23482=>"111110100",
  23483=>"100100111",
  23484=>"001000000",
  23485=>"001001111",
  23486=>"000011000",
  23487=>"000111110",
  23488=>"000001000",
  23489=>"001000011",
  23490=>"001101111",
  23491=>"110010100",
  23492=>"000000001",
  23493=>"000001011",
  23494=>"110100011",
  23495=>"111111111",
  23496=>"101101110",
  23497=>"110110100",
  23498=>"101101100",
  23499=>"100001110",
  23500=>"000011100",
  23501=>"000000000",
  23502=>"101001000",
  23503=>"111100100",
  23504=>"000110110",
  23505=>"111111101",
  23506=>"000001000",
  23507=>"100000001",
  23508=>"011010000",
  23509=>"001111001",
  23510=>"100100001",
  23511=>"110100011",
  23512=>"110110000",
  23513=>"000100100",
  23514=>"000001111",
  23515=>"000001101",
  23516=>"110111000",
  23517=>"000000110",
  23518=>"001000100",
  23519=>"011101001",
  23520=>"000011011",
  23521=>"100100100",
  23522=>"000110110",
  23523=>"100110110",
  23524=>"000000011",
  23525=>"111110110",
  23526=>"101111100",
  23527=>"000000110",
  23528=>"011110100",
  23529=>"001111111",
  23530=>"001001010",
  23531=>"111110110",
  23532=>"011001000",
  23533=>"101111001",
  23534=>"101000000",
  23535=>"011100111",
  23536=>"110001011",
  23537=>"110111110",
  23538=>"011100100",
  23539=>"110101011",
  23540=>"111100000",
  23541=>"001111101",
  23542=>"000001011",
  23543=>"000000100",
  23544=>"000001001",
  23545=>"011001011",
  23546=>"000011011",
  23547=>"000111110",
  23548=>"110111011",
  23549=>"000000110",
  23550=>"100001000",
  23551=>"011001010",
  23552=>"000001100",
  23553=>"111011000",
  23554=>"000000111",
  23555=>"011000000",
  23556=>"110100100",
  23557=>"000000111",
  23558=>"110111001",
  23559=>"100000100",
  23560=>"000000000",
  23561=>"000000000",
  23562=>"011111000",
  23563=>"001000111",
  23564=>"110111000",
  23565=>"111011001",
  23566=>"001000000",
  23567=>"110101000",
  23568=>"100001001",
  23569=>"000000111",
  23570=>"111111011",
  23571=>"111010000",
  23572=>"010111110",
  23573=>"101000000",
  23574=>"000011000",
  23575=>"111000000",
  23576=>"111000001",
  23577=>"110111001",
  23578=>"000000001",
  23579=>"000000110",
  23580=>"111110011",
  23581=>"111111001",
  23582=>"111111111",
  23583=>"001001101",
  23584=>"000000000",
  23585=>"101111111",
  23586=>"100010010",
  23587=>"100000000",
  23588=>"101111001",
  23589=>"100000010",
  23590=>"000000011",
  23591=>"000000011",
  23592=>"000001111",
  23593=>"111111110",
  23594=>"000000011",
  23595=>"111000000",
  23596=>"011001010",
  23597=>"010101101",
  23598=>"111000111",
  23599=>"011111011",
  23600=>"000000000",
  23601=>"100100110",
  23602=>"111111111",
  23603=>"110000110",
  23604=>"000110000",
  23605=>"111111111",
  23606=>"101011011",
  23607=>"101001000",
  23608=>"111101000",
  23609=>"111111111",
  23610=>"000000000",
  23611=>"000000010",
  23612=>"000001001",
  23613=>"111111111",
  23614=>"000000000",
  23615=>"110110010",
  23616=>"111111110",
  23617=>"100000110",
  23618=>"011010000",
  23619=>"001000000",
  23620=>"111111111",
  23621=>"110000000",
  23622=>"010110010",
  23623=>"110111101",
  23624=>"001001001",
  23625=>"000000000",
  23626=>"101001011",
  23627=>"111111110",
  23628=>"001000110",
  23629=>"101111100",
  23630=>"001001011",
  23631=>"000000010",
  23632=>"000011101",
  23633=>"101111111",
  23634=>"000001000",
  23635=>"001000000",
  23636=>"111111110",
  23637=>"101111100",
  23638=>"110111011",
  23639=>"001011111",
  23640=>"001111111",
  23641=>"000111110",
  23642=>"101001000",
  23643=>"011000000",
  23644=>"010110100",
  23645=>"001000000",
  23646=>"111111111",
  23647=>"001000000",
  23648=>"010001110",
  23649=>"011111111",
  23650=>"000000111",
  23651=>"000000000",
  23652=>"000110100",
  23653=>"111111111",
  23654=>"001001001",
  23655=>"000100000",
  23656=>"111011111",
  23657=>"001010111",
  23658=>"101111111",
  23659=>"000010101",
  23660=>"111000100",
  23661=>"010000101",
  23662=>"011000000",
  23663=>"111001110",
  23664=>"000000000",
  23665=>"111111011",
  23666=>"111101111",
  23667=>"010011000",
  23668=>"000000000",
  23669=>"101100110",
  23670=>"110000001",
  23671=>"111011100",
  23672=>"000000000",
  23673=>"000110101",
  23674=>"000000000",
  23675=>"010001000",
  23676=>"100100011",
  23677=>"000000000",
  23678=>"000000000",
  23679=>"000000000",
  23680=>"010000110",
  23681=>"000011010",
  23682=>"000000111",
  23683=>"000111101",
  23684=>"111111100",
  23685=>"100010010",
  23686=>"001101001",
  23687=>"011000110",
  23688=>"001011000",
  23689=>"011100000",
  23690=>"011011000",
  23691=>"010111111",
  23692=>"111001000",
  23693=>"000000011",
  23694=>"000110111",
  23695=>"111000001",
  23696=>"101111111",
  23697=>"000111101",
  23698=>"010000000",
  23699=>"001101000",
  23700=>"011010101",
  23701=>"000000000",
  23702=>"110111111",
  23703=>"011101100",
  23704=>"111000111",
  23705=>"000000001",
  23706=>"000100010",
  23707=>"000000000",
  23708=>"111101001",
  23709=>"101100111",
  23710=>"101111111",
  23711=>"000000000",
  23712=>"000010001",
  23713=>"000011111",
  23714=>"010100000",
  23715=>"000010101",
  23716=>"111111111",
  23717=>"110111011",
  23718=>"110111110",
  23719=>"001000001",
  23720=>"111000111",
  23721=>"111001001",
  23722=>"000000110",
  23723=>"101111111",
  23724=>"111100000",
  23725=>"001001111",
  23726=>"001111011",
  23727=>"000000110",
  23728=>"000000001",
  23729=>"100100101",
  23730=>"000010111",
  23731=>"001000010",
  23732=>"011111000",
  23733=>"110100100",
  23734=>"011111110",
  23735=>"010000000",
  23736=>"001000100",
  23737=>"111100001",
  23738=>"110010111",
  23739=>"010111111",
  23740=>"111111101",
  23741=>"111111111",
  23742=>"001000110",
  23743=>"000111111",
  23744=>"110111000",
  23745=>"000000100",
  23746=>"111111110",
  23747=>"000011100",
  23748=>"110111111",
  23749=>"000001000",
  23750=>"111010100",
  23751=>"100000000",
  23752=>"000000000",
  23753=>"101000000",
  23754=>"110011111",
  23755=>"111001010",
  23756=>"101000000",
  23757=>"011011100",
  23758=>"111111111",
  23759=>"000000111",
  23760=>"111000001",
  23761=>"100110110",
  23762=>"110110110",
  23763=>"111111011",
  23764=>"000000111",
  23765=>"111111001",
  23766=>"101100000",
  23767=>"110111001",
  23768=>"000001000",
  23769=>"000000000",
  23770=>"000000000",
  23771=>"000010111",
  23772=>"001000011",
  23773=>"110111101",
  23774=>"111110111",
  23775=>"111111101",
  23776=>"001000011",
  23777=>"000001011",
  23778=>"000000000",
  23779=>"000000000",
  23780=>"000000000",
  23781=>"000001000",
  23782=>"000000000",
  23783=>"001011010",
  23784=>"000000010",
  23785=>"111110001",
  23786=>"110111111",
  23787=>"110010000",
  23788=>"001000010",
  23789=>"111011000",
  23790=>"000000000",
  23791=>"000000101",
  23792=>"101101111",
  23793=>"001000011",
  23794=>"111000101",
  23795=>"101000000",
  23796=>"100001011",
  23797=>"000000001",
  23798=>"010010111",
  23799=>"000000100",
  23800=>"000000000",
  23801=>"101001000",
  23802=>"110111111",
  23803=>"111010000",
  23804=>"111111011",
  23805=>"010000111",
  23806=>"101011011",
  23807=>"000000000",
  23808=>"011001001",
  23809=>"000001110",
  23810=>"001000001",
  23811=>"000000001",
  23812=>"011111111",
  23813=>"000100110",
  23814=>"000010010",
  23815=>"111000000",
  23816=>"000000000",
  23817=>"010000010",
  23818=>"111111111",
  23819=>"000000000",
  23820=>"000011011",
  23821=>"010001001",
  23822=>"011111001",
  23823=>"000110011",
  23824=>"001101000",
  23825=>"000110000",
  23826=>"110111100",
  23827=>"111111111",
  23828=>"111100100",
  23829=>"111111111",
  23830=>"111111111",
  23831=>"000001000",
  23832=>"000000000",
  23833=>"111001101",
  23834=>"000000101",
  23835=>"010000000",
  23836=>"111111111",
  23837=>"001101111",
  23838=>"111110010",
  23839=>"000000000",
  23840=>"000110000",
  23841=>"111111111",
  23842=>"001000000",
  23843=>"000000000",
  23844=>"011111000",
  23845=>"110110010",
  23846=>"000101111",
  23847=>"000001101",
  23848=>"110110000",
  23849=>"111110110",
  23850=>"001111000",
  23851=>"111101010",
  23852=>"111111111",
  23853=>"100000000",
  23854=>"000001000",
  23855=>"011001111",
  23856=>"000000000",
  23857=>"011111000",
  23858=>"000000000",
  23859=>"111110010",
  23860=>"111111111",
  23861=>"111111111",
  23862=>"110110101",
  23863=>"101000010",
  23864=>"111101111",
  23865=>"000000000",
  23866=>"000000001",
  23867=>"010001000",
  23868=>"001110000",
  23869=>"111111111",
  23870=>"001000100",
  23871=>"101001100",
  23872=>"011000111",
  23873=>"011111011",
  23874=>"111110000",
  23875=>"001000100",
  23876=>"111111111",
  23877=>"000000000",
  23878=>"010010010",
  23879=>"111110010",
  23880=>"000101001",
  23881=>"000000000",
  23882=>"000000001",
  23883=>"001000001",
  23884=>"001000001",
  23885=>"111011000",
  23886=>"110111110",
  23887=>"110110110",
  23888=>"111011100",
  23889=>"110010100",
  23890=>"000001111",
  23891=>"001000111",
  23892=>"000000001",
  23893=>"111111101",
  23894=>"111111000",
  23895=>"001000001",
  23896=>"010000000",
  23897=>"111110111",
  23898=>"111111111",
  23899=>"111100111",
  23900=>"111000000",
  23901=>"001001001",
  23902=>"110111010",
  23903=>"100000000",
  23904=>"001000000",
  23905=>"000001001",
  23906=>"111110010",
  23907=>"000110011",
  23908=>"000110100",
  23909=>"111000000",
  23910=>"000000001",
  23911=>"000100100",
  23912=>"001001111",
  23913=>"011101000",
  23914=>"111111110",
  23915=>"000000111",
  23916=>"011000100",
  23917=>"010111000",
  23918=>"001000010",
  23919=>"010011000",
  23920=>"110110111",
  23921=>"011111110",
  23922=>"011111111",
  23923=>"000000101",
  23924=>"000001111",
  23925=>"100000100",
  23926=>"111111111",
  23927=>"100110110",
  23928=>"000000000",
  23929=>"111111000",
  23930=>"111111100",
  23931=>"000001001",
  23932=>"111111111",
  23933=>"100110101",
  23934=>"011111111",
  23935=>"001000001",
  23936=>"001111111",
  23937=>"111111111",
  23938=>"010011010",
  23939=>"111111110",
  23940=>"001000110",
  23941=>"111101000",
  23942=>"100111100",
  23943=>"000100000",
  23944=>"011011001",
  23945=>"010010001",
  23946=>"000000000",
  23947=>"000000000",
  23948=>"000000000",
  23949=>"110010111",
  23950=>"001000011",
  23951=>"000001000",
  23952=>"101111001",
  23953=>"000111111",
  23954=>"000000111",
  23955=>"000000110",
  23956=>"011111110",
  23957=>"000110011",
  23958=>"110110000",
  23959=>"000001000",
  23960=>"111111111",
  23961=>"000110111",
  23962=>"010010010",
  23963=>"100000010",
  23964=>"000010011",
  23965=>"000110010",
  23966=>"000111010",
  23967=>"001000001",
  23968=>"001101000",
  23969=>"010111101",
  23970=>"000000101",
  23971=>"000000000",
  23972=>"001001111",
  23973=>"000011011",
  23974=>"101101001",
  23975=>"011111101",
  23976=>"110111111",
  23977=>"100110100",
  23978=>"000110100",
  23979=>"011011111",
  23980=>"011100000",
  23981=>"100100110",
  23982=>"100100101",
  23983=>"111111010",
  23984=>"000000000",
  23985=>"011101000",
  23986=>"000111011",
  23987=>"001101000",
  23988=>"001000100",
  23989=>"111111111",
  23990=>"011000000",
  23991=>"010110000",
  23992=>"110111011",
  23993=>"011010011",
  23994=>"101101010",
  23995=>"000000000",
  23996=>"000011000",
  23997=>"111111010",
  23998=>"100000000",
  23999=>"000000000",
  24000=>"000000000",
  24001=>"011000011",
  24002=>"000111111",
  24003=>"011111111",
  24004=>"000000000",
  24005=>"110111110",
  24006=>"010110110",
  24007=>"111001111",
  24008=>"000000000",
  24009=>"000000100",
  24010=>"001000000",
  24011=>"111111111",
  24012=>"001000000",
  24013=>"111111111",
  24014=>"111011111",
  24015=>"110010011",
  24016=>"000000110",
  24017=>"100110000",
  24018=>"000000000",
  24019=>"001000011",
  24020=>"000101111",
  24021=>"000100000",
  24022=>"000000000",
  24023=>"111111111",
  24024=>"000000100",
  24025=>"010101101",
  24026=>"111101100",
  24027=>"000111111",
  24028=>"111111110",
  24029=>"000000001",
  24030=>"100000011",
  24031=>"110010000",
  24032=>"010000010",
  24033=>"000000000",
  24034=>"000110000",
  24035=>"010000000",
  24036=>"000000100",
  24037=>"001110111",
  24038=>"001111111",
  24039=>"111011001",
  24040=>"101101110",
  24041=>"000101111",
  24042=>"111111111",
  24043=>"101111111",
  24044=>"000000000",
  24045=>"100101000",
  24046=>"110001010",
  24047=>"000000000",
  24048=>"111000010",
  24049=>"111111111",
  24050=>"001000010",
  24051=>"001111111",
  24052=>"100110100",
  24053=>"111011101",
  24054=>"000000111",
  24055=>"101100101",
  24056=>"000001000",
  24057=>"111000111",
  24058=>"010010000",
  24059=>"000111011",
  24060=>"110111111",
  24061=>"111111111",
  24062=>"110110010",
  24063=>"101111101",
  24064=>"001001110",
  24065=>"011011010",
  24066=>"111101101",
  24067=>"011010100",
  24068=>"000011111",
  24069=>"101010011",
  24070=>"000000010",
  24071=>"000000000",
  24072=>"000100010",
  24073=>"111011000",
  24074=>"001000100",
  24075=>"100100000",
  24076=>"101100011",
  24077=>"001111101",
  24078=>"110100000",
  24079=>"100111000",
  24080=>"010011011",
  24081=>"100000100",
  24082=>"100010000",
  24083=>"000000010",
  24084=>"111111001",
  24085=>"011100111",
  24086=>"111110111",
  24087=>"111001011",
  24088=>"100100110",
  24089=>"000010011",
  24090=>"000101100",
  24091=>"111101000",
  24092=>"100100100",
  24093=>"100100001",
  24094=>"111010000",
  24095=>"000100111",
  24096=>"001111111",
  24097=>"011000000",
  24098=>"111101101",
  24099=>"000100011",
  24100=>"000000110",
  24101=>"110110111",
  24102=>"000000111",
  24103=>"000101101",
  24104=>"010011011",
  24105=>"000011111",
  24106=>"010010111",
  24107=>"001011001",
  24108=>"000100000",
  24109=>"001101011",
  24110=>"111011111",
  24111=>"000000000",
  24112=>"000010010",
  24113=>"000000001",
  24114=>"011011101",
  24115=>"101111100",
  24116=>"100101000",
  24117=>"101101000",
  24118=>"000000001",
  24119=>"000000000",
  24120=>"000010010",
  24121=>"011000101",
  24122=>"111100100",
  24123=>"001000111",
  24124=>"011110110",
  24125=>"111111011",
  24126=>"000100100",
  24127=>"001110010",
  24128=>"111111000",
  24129=>"011111101",
  24130=>"111000000",
  24131=>"001011010",
  24132=>"011000000",
  24133=>"000011011",
  24134=>"000000010",
  24135=>"111000000",
  24136=>"000011011",
  24137=>"011000000",
  24138=>"000001111",
  24139=>"010011011",
  24140=>"111111011",
  24141=>"001111111",
  24142=>"000001100",
  24143=>"111101000",
  24144=>"000100111",
  24145=>"111011000",
  24146=>"011010011",
  24147=>"011001000",
  24148=>"111111100",
  24149=>"001001001",
  24150=>"111100111",
  24151=>"111011000",
  24152=>"101100110",
  24153=>"000100101",
  24154=>"011011101",
  24155=>"001101100",
  24156=>"010010010",
  24157=>"000000001",
  24158=>"011111001",
  24159=>"100110010",
  24160=>"000011111",
  24161=>"011011111",
  24162=>"100100110",
  24163=>"110010010",
  24164=>"000000010",
  24165=>"110111101",
  24166=>"111111000",
  24167=>"010011101",
  24168=>"100111111",
  24169=>"011000100",
  24170=>"101000000",
  24171=>"100010111",
  24172=>"000010011",
  24173=>"000000000",
  24174=>"001010000",
  24175=>"010001000",
  24176=>"000101001",
  24177=>"000110000",
  24178=>"000000010",
  24179=>"100111111",
  24180=>"110111100",
  24181=>"000000100",
  24182=>"111111011",
  24183=>"000101101",
  24184=>"111000100",
  24185=>"111000110",
  24186=>"000001111",
  24187=>"000000001",
  24188=>"110110110",
  24189=>"110100000",
  24190=>"011011011",
  24191=>"100100101",
  24192=>"011010100",
  24193=>"011100000",
  24194=>"001000000",
  24195=>"100000011",
  24196=>"101100010",
  24197=>"000111111",
  24198=>"011011011",
  24199=>"000001111",
  24200=>"000110111",
  24201=>"011010001",
  24202=>"011000100",
  24203=>"000110101",
  24204=>"000000100",
  24205=>"101101111",
  24206=>"100100100",
  24207=>"000000001",
  24208=>"001101101",
  24209=>"111111110",
  24210=>"000000100",
  24211=>"101000000",
  24212=>"000000000",
  24213=>"111011000",
  24214=>"110000000",
  24215=>"010100011",
  24216=>"111101100",
  24217=>"010001000",
  24218=>"100111111",
  24219=>"000000000",
  24220=>"111110000",
  24221=>"111011111",
  24222=>"011101100",
  24223=>"000000000",
  24224=>"100001010",
  24225=>"100101111",
  24226=>"000000111",
  24227=>"111000011",
  24228=>"100100111",
  24229=>"000111011",
  24230=>"111010111",
  24231=>"001111111",
  24232=>"111000111",
  24233=>"101001111",
  24234=>"101000000",
  24235=>"000010110",
  24236=>"111000100",
  24237=>"101000100",
  24238=>"001001000",
  24239=>"011011011",
  24240=>"000011000",
  24241=>"100111011",
  24242=>"000001011",
  24243=>"000001100",
  24244=>"100100111",
  24245=>"110111011",
  24246=>"101000111",
  24247=>"111011101",
  24248=>"110001011",
  24249=>"000100011",
  24250=>"000111111",
  24251=>"111000000",
  24252=>"011111000",
  24253=>"111111111",
  24254=>"000001001",
  24255=>"000111111",
  24256=>"100010010",
  24257=>"000000000",
  24258=>"011011011",
  24259=>"000000111",
  24260=>"000000001",
  24261=>"110000000",
  24262=>"010010011",
  24263=>"101000100",
  24264=>"000100000",
  24265=>"000000011",
  24266=>"100011011",
  24267=>"100110110",
  24268=>"000011011",
  24269=>"011000001",
  24270=>"111110000",
  24271=>"111111101",
  24272=>"011000101",
  24273=>"001001110",
  24274=>"000100111",
  24275=>"100100100",
  24276=>"100111101",
  24277=>"000100110",
  24278=>"111000000",
  24279=>"011010000",
  24280=>"000111000",
  24281=>"100111000",
  24282=>"001000100",
  24283=>"111000000",
  24284=>"001001110",
  24285=>"000001001",
  24286=>"100000000",
  24287=>"111011000",
  24288=>"000000001",
  24289=>"001001001",
  24290=>"101000111",
  24291=>"001001001",
  24292=>"000011111",
  24293=>"000010111",
  24294=>"000010011",
  24295=>"100100100",
  24296=>"011101000",
  24297=>"111000101",
  24298=>"110000001",
  24299=>"111111100",
  24300=>"010011010",
  24301=>"100100000",
  24302=>"111000000",
  24303=>"000000010",
  24304=>"000000000",
  24305=>"000100000",
  24306=>"111111101",
  24307=>"001101100",
  24308=>"100110101",
  24309=>"111000000",
  24310=>"000000000",
  24311=>"000100000",
  24312=>"000000110",
  24313=>"111111000",
  24314=>"111101101",
  24315=>"100000111",
  24316=>"111000000",
  24317=>"001111111",
  24318=>"110100111",
  24319=>"101011010",
  24320=>"100011100",
  24321=>"001000001",
  24322=>"011010010",
  24323=>"111101111",
  24324=>"011111111",
  24325=>"110101110",
  24326=>"000000111",
  24327=>"000000011",
  24328=>"110100000",
  24329=>"110110011",
  24330=>"111000000",
  24331=>"111011111",
  24332=>"111111001",
  24333=>"100000000",
  24334=>"101011011",
  24335=>"100011010",
  24336=>"011111100",
  24337=>"001111110",
  24338=>"111101100",
  24339=>"000000101",
  24340=>"010011000",
  24341=>"101100100",
  24342=>"000000011",
  24343=>"110111110",
  24344=>"000100001",
  24345=>"101101011",
  24346=>"011100111",
  24347=>"100000111",
  24348=>"111110111",
  24349=>"000100001",
  24350=>"011110110",
  24351=>"001001000",
  24352=>"011111000",
  24353=>"010111100",
  24354=>"111000001",
  24355=>"111000110",
  24356=>"010111001",
  24357=>"000100000",
  24358=>"000000000",
  24359=>"110001111",
  24360=>"001101000",
  24361=>"110100000",
  24362=>"010010110",
  24363=>"011111011",
  24364=>"100111001",
  24365=>"100000000",
  24366=>"011111000",
  24367=>"000000001",
  24368=>"111011011",
  24369=>"000001001",
  24370=>"011111110",
  24371=>"010110110",
  24372=>"001001001",
  24373=>"111110110",
  24374=>"011001011",
  24375=>"100000100",
  24376=>"010111010",
  24377=>"100000110",
  24378=>"111000000",
  24379=>"111001011",
  24380=>"000110000",
  24381=>"001001000",
  24382=>"110100000",
  24383=>"001011010",
  24384=>"101011000",
  24385=>"001000000",
  24386=>"101011000",
  24387=>"000011100",
  24388=>"111000011",
  24389=>"000111111",
  24390=>"110000001",
  24391=>"011111011",
  24392=>"111110000",
  24393=>"111110000",
  24394=>"010100100",
  24395=>"001001101",
  24396=>"000100101",
  24397=>"001011011",
  24398=>"010001000",
  24399=>"110001011",
  24400=>"001000000",
  24401=>"100111111",
  24402=>"111100010",
  24403=>"111000000",
  24404=>"001000000",
  24405=>"011000001",
  24406=>"101001001",
  24407=>"111110100",
  24408=>"111100101",
  24409=>"001011011",
  24410=>"001000001",
  24411=>"000001110",
  24412=>"111111111",
  24413=>"100000101",
  24414=>"110111010",
  24415=>"001011000",
  24416=>"111111011",
  24417=>"011001000",
  24418=>"011110011",
  24419=>"000000000",
  24420=>"110000000",
  24421=>"001111000",
  24422=>"001100001",
  24423=>"101000000",
  24424=>"001101000",
  24425=>"000010010",
  24426=>"010010111",
  24427=>"100100111",
  24428=>"111011111",
  24429=>"100100110",
  24430=>"110100000",
  24431=>"110000011",
  24432=>"001011011",
  24433=>"011111110",
  24434=>"111000001",
  24435=>"011000000",
  24436=>"111001111",
  24437=>"100100101",
  24438=>"000100110",
  24439=>"111000100",
  24440=>"011110000",
  24441=>"110001110",
  24442=>"000001111",
  24443=>"100100000",
  24444=>"000000001",
  24445=>"110000000",
  24446=>"111000100",
  24447=>"011000000",
  24448=>"000110110",
  24449=>"111000100",
  24450=>"110000001",
  24451=>"011000001",
  24452=>"110100001",
  24453=>"110100111",
  24454=>"010111000",
  24455=>"000001010",
  24456=>"001001001",
  24457=>"011000000",
  24458=>"000000100",
  24459=>"101100110",
  24460=>"111110100",
  24461=>"101100011",
  24462=>"110000001",
  24463=>"011011000",
  24464=>"010011011",
  24465=>"011110000",
  24466=>"001001000",
  24467=>"001001001",
  24468=>"001011111",
  24469=>"000110110",
  24470=>"000011010",
  24471=>"111011011",
  24472=>"100100111",
  24473=>"111110011",
  24474=>"011110011",
  24475=>"100000000",
  24476=>"000100100",
  24477=>"111110101",
  24478=>"010000110",
  24479=>"001100101",
  24480=>"110100000",
  24481=>"111110100",
  24482=>"111001000",
  24483=>"111010100",
  24484=>"110000111",
  24485=>"011001001",
  24486=>"110101001",
  24487=>"001111111",
  24488=>"100010110",
  24489=>"001001111",
  24490=>"111000000",
  24491=>"110000001",
  24492=>"000010101",
  24493=>"011000001",
  24494=>"011100100",
  24495=>"111110000",
  24496=>"010110000",
  24497=>"100111111",
  24498=>"110000011",
  24499=>"000000000",
  24500=>"111111001",
  24501=>"001100100",
  24502=>"011011111",
  24503=>"000000001",
  24504=>"100100110",
  24505=>"010000000",
  24506=>"111110100",
  24507=>"000011011",
  24508=>"000000111",
  24509=>"111111111",
  24510=>"111001000",
  24511=>"011011110",
  24512=>"110110000",
  24513=>"010000000",
  24514=>"000001011",
  24515=>"000011100",
  24516=>"000000000",
  24517=>"010000101",
  24518=>"100011001",
  24519=>"111100100",
  24520=>"001000011",
  24521=>"000000010",
  24522=>"001010000",
  24523=>"011010111",
  24524=>"000111000",
  24525=>"001001001",
  24526=>"000001100",
  24527=>"111111111",
  24528=>"011111110",
  24529=>"000001011",
  24530=>"011100000",
  24531=>"111101000",
  24532=>"010010001",
  24533=>"000000000",
  24534=>"110111111",
  24535=>"010011111",
  24536=>"111111001",
  24537=>"010010000",
  24538=>"001001001",
  24539=>"111100100",
  24540=>"001011011",
  24541=>"101101101",
  24542=>"000010000",
  24543=>"001011110",
  24544=>"110111011",
  24545=>"000010011",
  24546=>"111100110",
  24547=>"111110110",
  24548=>"000110100",
  24549=>"010100111",
  24550=>"001111000",
  24551=>"100100110",
  24552=>"110111111",
  24553=>"101110000",
  24554=>"110111010",
  24555=>"111111110",
  24556=>"001100000",
  24557=>"001011111",
  24558=>"000111100",
  24559=>"110000110",
  24560=>"111001001",
  24561=>"100101111",
  24562=>"110000010",
  24563=>"101011000",
  24564=>"001101001",
  24565=>"110000000",
  24566=>"000100110",
  24567=>"000000111",
  24568=>"011111110",
  24569=>"110111100",
  24570=>"110111101",
  24571=>"100001001",
  24572=>"000001001",
  24573=>"100010110",
  24574=>"110000001",
  24575=>"001001011",
  24576=>"100100111",
  24577=>"010010010",
  24578=>"101111111",
  24579=>"000000000",
  24580=>"000100100",
  24581=>"000111111",
  24582=>"100100100",
  24583=>"011111111",
  24584=>"101101101",
  24585=>"000000000",
  24586=>"111100100",
  24587=>"110000000",
  24588=>"000100111",
  24589=>"000000111",
  24590=>"011000000",
  24591=>"111111111",
  24592=>"000000000",
  24593=>"000000101",
  24594=>"001000000",
  24595=>"011011000",
  24596=>"111011111",
  24597=>"110000000",
  24598=>"111111011",
  24599=>"011000000",
  24600=>"100000000",
  24601=>"111111111",
  24602=>"000000000",
  24603=>"000000100",
  24604=>"111101111",
  24605=>"000000000",
  24606=>"000000111",
  24607=>"010010000",
  24608=>"010110010",
  24609=>"000010000",
  24610=>"000000000",
  24611=>"100110011",
  24612=>"110011001",
  24613=>"111001011",
  24614=>"111000000",
  24615=>"111110101",
  24616=>"010111011",
  24617=>"011101100",
  24618=>"111111000",
  24619=>"000001000",
  24620=>"111001000",
  24621=>"110011010",
  24622=>"100000000",
  24623=>"010111111",
  24624=>"110111010",
  24625=>"001000000",
  24626=>"011100001",
  24627=>"110000000",
  24628=>"111100110",
  24629=>"110000000",
  24630=>"011000000",
  24631=>"011000010",
  24632=>"000110111",
  24633=>"011101100",
  24634=>"110011100",
  24635=>"100110110",
  24636=>"010011011",
  24637=>"011000111",
  24638=>"000011111",
  24639=>"000000100",
  24640=>"011111101",
  24641=>"110101111",
  24642=>"100000001",
  24643=>"101101111",
  24644=>"111111111",
  24645=>"000000000",
  24646=>"111101111",
  24647=>"011110011",
  24648=>"110011111",
  24649=>"000010010",
  24650=>"000010000",
  24651=>"101100101",
  24652=>"100110111",
  24653=>"011111111",
  24654=>"100110010",
  24655=>"111000000",
  24656=>"110000000",
  24657=>"111111010",
  24658=>"111110111",
  24659=>"110110100",
  24660=>"010100100",
  24661=>"110101001",
  24662=>"111111000",
  24663=>"111001111",
  24664=>"101111101",
  24665=>"111001010",
  24666=>"000001000",
  24667=>"110000100",
  24668=>"100000000",
  24669=>"011011011",
  24670=>"101100101",
  24671=>"001001111",
  24672=>"000100100",
  24673=>"010010010",
  24674=>"000000000",
  24675=>"100100000",
  24676=>"111111111",
  24677=>"101111011",
  24678=>"010010110",
  24679=>"011110000",
  24680=>"000000000",
  24681=>"011011111",
  24682=>"010111101",
  24683=>"111101101",
  24684=>"001100000",
  24685=>"010111001",
  24686=>"000111110",
  24687=>"111111101",
  24688=>"110110110",
  24689=>"000000000",
  24690=>"001000000",
  24691=>"101000000",
  24692=>"000110000",
  24693=>"000011010",
  24694=>"000000000",
  24695=>"100111111",
  24696=>"000000000",
  24697=>"011000000",
  24698=>"111111010",
  24699=>"000100011",
  24700=>"111011001",
  24701=>"011011011",
  24702=>"000101000",
  24703=>"101000011",
  24704=>"000010110",
  24705=>"011111000",
  24706=>"000000000",
  24707=>"011011101",
  24708=>"000000000",
  24709=>"111101000",
  24710=>"110100110",
  24711=>"111110110",
  24712=>"011011011",
  24713=>"111101111",
  24714=>"000000000",
  24715=>"101101000",
  24716=>"111111111",
  24717=>"011010010",
  24718=>"000000000",
  24719=>"101000100",
  24720=>"110110110",
  24721=>"001000000",
  24722=>"100101000",
  24723=>"011101110",
  24724=>"000100000",
  24725=>"010111111",
  24726=>"111100000",
  24727=>"001110010",
  24728=>"111101100",
  24729=>"010111101",
  24730=>"000000000",
  24731=>"000011000",
  24732=>"010100100",
  24733=>"000000000",
  24734=>"010111111",
  24735=>"110000000",
  24736=>"111110111",
  24737=>"000011000",
  24738=>"111111000",
  24739=>"011011000",
  24740=>"000001110",
  24741=>"011011011",
  24742=>"000010010",
  24743=>"000000000",
  24744=>"100110000",
  24745=>"111101000",
  24746=>"000010111",
  24747=>"110111111",
  24748=>"110010010",
  24749=>"010111111",
  24750=>"011001001",
  24751=>"001000111",
  24752=>"100001111",
  24753=>"110110111",
  24754=>"000000000",
  24755=>"010011000",
  24756=>"111110000",
  24757=>"001000001",
  24758=>"001111000",
  24759=>"111001110",
  24760=>"110110010",
  24761=>"011001001",
  24762=>"110000000",
  24763=>"000110111",
  24764=>"000100100",
  24765=>"111111111",
  24766=>"110100000",
  24767=>"000000110",
  24768=>"111011011",
  24769=>"000010000",
  24770=>"000101110",
  24771=>"110011011",
  24772=>"101000000",
  24773=>"011111110",
  24774=>"000010000",
  24775=>"100000100",
  24776=>"111111111",
  24777=>"101101111",
  24778=>"000011000",
  24779=>"110100101",
  24780=>"110000000",
  24781=>"110110000",
  24782=>"111111100",
  24783=>"000000000",
  24784=>"010100000",
  24785=>"110110110",
  24786=>"010000000",
  24787=>"010100000",
  24788=>"000011111",
  24789=>"111111110",
  24790=>"101101000",
  24791=>"001010000",
  24792=>"000000000",
  24793=>"000000000",
  24794=>"111111101",
  24795=>"110110000",
  24796=>"101011110",
  24797=>"010000000",
  24798=>"100100000",
  24799=>"000000101",
  24800=>"000000000",
  24801=>"000011010",
  24802=>"000000000",
  24803=>"111010011",
  24804=>"111000000",
  24805=>"111100100",
  24806=>"110000100",
  24807=>"110010000",
  24808=>"110111111",
  24809=>"110100000",
  24810=>"111000000",
  24811=>"111101101",
  24812=>"000000010",
  24813=>"110000000",
  24814=>"000111010",
  24815=>"000111010",
  24816=>"010000000",
  24817=>"110101111",
  24818=>"000101111",
  24819=>"110000000",
  24820=>"100000011",
  24821=>"100100000",
  24822=>"111111111",
  24823=>"100100000",
  24824=>"000111101",
  24825=>"111111100",
  24826=>"111111110",
  24827=>"010110000",
  24828=>"101101101",
  24829=>"010010111",
  24830=>"111111111",
  24831=>"000000000",
  24832=>"010100100",
  24833=>"011111111",
  24834=>"000010111",
  24835=>"111111101",
  24836=>"010010111",
  24837=>"010011011",
  24838=>"000000000",
  24839=>"000111000",
  24840=>"010100000",
  24841=>"000000101",
  24842=>"001100100",
  24843=>"010101101",
  24844=>"000000000",
  24845=>"110100000",
  24846=>"110000000",
  24847=>"100000000",
  24848=>"110111101",
  24849=>"000111101",
  24850=>"110111110",
  24851=>"000100111",
  24852=>"101000010",
  24853=>"010011001",
  24854=>"010110111",
  24855=>"111111000",
  24856=>"000000000",
  24857=>"000000001",
  24858=>"000000111",
  24859=>"000111111",
  24860=>"011111001",
  24861=>"111110101",
  24862=>"010111111",
  24863=>"000000111",
  24864=>"111000101",
  24865=>"000001110",
  24866=>"000001100",
  24867=>"000111111",
  24868=>"110110110",
  24869=>"110000000",
  24870=>"000010100",
  24871=>"011011101",
  24872=>"111110010",
  24873=>"010000000",
  24874=>"110000000",
  24875=>"111000100",
  24876=>"110111000",
  24877=>"111101101",
  24878=>"110111101",
  24879=>"110001000",
  24880=>"100000100",
  24881=>"011111110",
  24882=>"000000000",
  24883=>"011101001",
  24884=>"110110000",
  24885=>"111111101",
  24886=>"111100000",
  24887=>"111101111",
  24888=>"001000011",
  24889=>"000000111",
  24890=>"111101000",
  24891=>"000000010",
  24892=>"011001001",
  24893=>"111111111",
  24894=>"101000100",
  24895=>"111011111",
  24896=>"111100000",
  24897=>"010000010",
  24898=>"011001000",
  24899=>"110110110",
  24900=>"110001110",
  24901=>"000101101",
  24902=>"000100000",
  24903=>"101101101",
  24904=>"111010000",
  24905=>"000000101",
  24906=>"000000000",
  24907=>"000000000",
  24908=>"111000100",
  24909=>"111010011",
  24910=>"110110011",
  24911=>"011111010",
  24912=>"101001000",
  24913=>"111111110",
  24914=>"111111101",
  24915=>"111011000",
  24916=>"010111010",
  24917=>"011110111",
  24918=>"000110011",
  24919=>"000010010",
  24920=>"011111111",
  24921=>"001001101",
  24922=>"110101100",
  24923=>"110010000",
  24924=>"000000101",
  24925=>"001001100",
  24926=>"111111010",
  24927=>"110111110",
  24928=>"000001111",
  24929=>"000111011",
  24930=>"101000000",
  24931=>"110110001",
  24932=>"010000001",
  24933=>"000100000",
  24934=>"010111000",
  24935=>"111010000",
  24936=>"000111111",
  24937=>"100000111",
  24938=>"000011111",
  24939=>"111011000",
  24940=>"111110100",
  24941=>"101111100",
  24942=>"100000000",
  24943=>"101101000",
  24944=>"000000110",
  24945=>"000000010",
  24946=>"001000000",
  24947=>"100000000",
  24948=>"010111111",
  24949=>"000101111",
  24950=>"000000010",
  24951=>"100100000",
  24952=>"000111111",
  24953=>"000111110",
  24954=>"101000101",
  24955=>"110000101",
  24956=>"111111000",
  24957=>"110001011",
  24958=>"111000001",
  24959=>"000111101",
  24960=>"010011011",
  24961=>"111101100",
  24962=>"111000001",
  24963=>"101111110",
  24964=>"010111111",
  24965=>"011001001",
  24966=>"010001110",
  24967=>"010000100",
  24968=>"010000001",
  24969=>"110000101",
  24970=>"000011011",
  24971=>"000100111",
  24972=>"101000101",
  24973=>"101000101",
  24974=>"100101000",
  24975=>"000000000",
  24976=>"111011001",
  24977=>"011001111",
  24978=>"101001100",
  24979=>"000111000",
  24980=>"110011100",
  24981=>"000000111",
  24982=>"110000111",
  24983=>"100100100",
  24984=>"100101001",
  24985=>"011111111",
  24986=>"111000000",
  24987=>"000110000",
  24988=>"010101000",
  24989=>"110100000",
  24990=>"000010111",
  24991=>"100000001",
  24992=>"111010010",
  24993=>"000110110",
  24994=>"000001000",
  24995=>"000000000",
  24996=>"110001101",
  24997=>"101110111",
  24998=>"001000110",
  24999=>"111111101",
  25000=>"101011011",
  25001=>"100101101",
  25002=>"000000101",
  25003=>"111000000",
  25004=>"100101101",
  25005=>"001000100",
  25006=>"011000100",
  25007=>"010000010",
  25008=>"110111010",
  25009=>"110100101",
  25010=>"000001011",
  25011=>"000000000",
  25012=>"000011011",
  25013=>"000000000",
  25014=>"110010110",
  25015=>"010000001",
  25016=>"110110000",
  25017=>"000010011",
  25018=>"000000000",
  25019=>"001000101",
  25020=>"011000010",
  25021=>"101000101",
  25022=>"100100100",
  25023=>"000000000",
  25024=>"000010110",
  25025=>"000000001",
  25026=>"011000000",
  25027=>"011000101",
  25028=>"110000000",
  25029=>"111100000",
  25030=>"000011100",
  25031=>"010011010",
  25032=>"110111000",
  25033=>"001111111",
  25034=>"110001111",
  25035=>"111110110",
  25036=>"000011010",
  25037=>"011110000",
  25038=>"101001100",
  25039=>"100000010",
  25040=>"111111111",
  25041=>"010011110",
  25042=>"010111011",
  25043=>"101100110",
  25044=>"011011000",
  25045=>"000001001",
  25046=>"010011111",
  25047=>"100001111",
  25048=>"010011010",
  25049=>"100000000",
  25050=>"011010000",
  25051=>"101000000",
  25052=>"111111111",
  25053=>"010111100",
  25054=>"000000000",
  25055=>"100101111",
  25056=>"010011010",
  25057=>"100000110",
  25058=>"000111111",
  25059=>"011010000",
  25060=>"000010010",
  25061=>"011111000",
  25062=>"111001000",
  25063=>"100111011",
  25064=>"111111111",
  25065=>"000000000",
  25066=>"010000000",
  25067=>"111101111",
  25068=>"000000000",
  25069=>"000000010",
  25070=>"000000100",
  25071=>"010111111",
  25072=>"010100101",
  25073=>"111000000",
  25074=>"010000000",
  25075=>"010110100",
  25076=>"001001001",
  25077=>"101110101",
  25078=>"111001001",
  25079=>"111111100",
  25080=>"111000000",
  25081=>"001000000",
  25082=>"011111111",
  25083=>"000000101",
  25084=>"010010111",
  25085=>"111111111",
  25086=>"010010100",
  25087=>"000101000",
  25088=>"010010000",
  25089=>"100110010",
  25090=>"100111000",
  25091=>"000101110",
  25092=>"100011011",
  25093=>"110000000",
  25094=>"111111111",
  25095=>"010000010",
  25096=>"000000000",
  25097=>"111111000",
  25098=>"110110100",
  25099=>"101101111",
  25100=>"100111111",
  25101=>"110011111",
  25102=>"100010011",
  25103=>"110100000",
  25104=>"110001101",
  25105=>"000000001",
  25106=>"000000000",
  25107=>"111001000",
  25108=>"000000000",
  25109=>"011010000",
  25110=>"011000000",
  25111=>"010111011",
  25112=>"100000011",
  25113=>"111111111",
  25114=>"010000111",
  25115=>"000000000",
  25116=>"100110111",
  25117=>"000000101",
  25118=>"111000000",
  25119=>"001111111",
  25120=>"111101101",
  25121=>"100111111",
  25122=>"000110111",
  25123=>"010000000",
  25124=>"000001101",
  25125=>"001010101",
  25126=>"010010010",
  25127=>"000001001",
  25128=>"111000000",
  25129=>"111101111",
  25130=>"010010000",
  25131=>"101111111",
  25132=>"011000011",
  25133=>"001000000",
  25134=>"111111011",
  25135=>"000000000",
  25136=>"000101111",
  25137=>"111111011",
  25138=>"000001001",
  25139=>"000000000",
  25140=>"000000000",
  25141=>"101110000",
  25142=>"010001011",
  25143=>"000000000",
  25144=>"000000010",
  25145=>"000000000",
  25146=>"010000000",
  25147=>"001101101",
  25148=>"000000000",
  25149=>"011111111",
  25150=>"100100101",
  25151=>"110110110",
  25152=>"111111011",
  25153=>"001001010",
  25154=>"110110000",
  25155=>"011000000",
  25156=>"000111111",
  25157=>"000001111",
  25158=>"111111000",
  25159=>"010001000",
  25160=>"100000101",
  25161=>"011001111",
  25162=>"000001000",
  25163=>"000001001",
  25164=>"000001001",
  25165=>"000001110",
  25166=>"110110100",
  25167=>"111011111",
  25168=>"000111000",
  25169=>"111111111",
  25170=>"101110000",
  25171=>"111011100",
  25172=>"111010000",
  25173=>"001000101",
  25174=>"001001000",
  25175=>"000000000",
  25176=>"011110110",
  25177=>"111001001",
  25178=>"011011010",
  25179=>"101000100",
  25180=>"000001111",
  25181=>"010001001",
  25182=>"000101111",
  25183=>"000000001",
  25184=>"111111011",
  25185=>"001001010",
  25186=>"001011010",
  25187=>"100000000",
  25188=>"111100000",
  25189=>"111111000",
  25190=>"000100010",
  25191=>"110010000",
  25192=>"111111111",
  25193=>"000000011",
  25194=>"010000111",
  25195=>"100111001",
  25196=>"000100111",
  25197=>"010111101",
  25198=>"010110000",
  25199=>"010000001",
  25200=>"111011111",
  25201=>"000000010",
  25202=>"110100110",
  25203=>"111111010",
  25204=>"110110111",
  25205=>"000000000",
  25206=>"000000110",
  25207=>"000000000",
  25208=>"100000000",
  25209=>"111101111",
  25210=>"111011001",
  25211=>"010000000",
  25212=>"001100000",
  25213=>"000000000",
  25214=>"110011111",
  25215=>"000000000",
  25216=>"110111101",
  25217=>"110100000",
  25218=>"000000111",
  25219=>"000000000",
  25220=>"111100000",
  25221=>"011000101",
  25222=>"100100100",
  25223=>"100101011",
  25224=>"111101001",
  25225=>"000001000",
  25226=>"010101010",
  25227=>"101000001",
  25228=>"000001001",
  25229=>"000101111",
  25230=>"000000111",
  25231=>"101000000",
  25232=>"000101100",
  25233=>"110110111",
  25234=>"000000111",
  25235=>"111000001",
  25236=>"100111111",
  25237=>"001000000",
  25238=>"000000111",
  25239=>"011001011",
  25240=>"101101111",
  25241=>"000000001",
  25242=>"100110111",
  25243=>"111000000",
  25244=>"001000001",
  25245=>"100001101",
  25246=>"111111101",
  25247=>"001001000",
  25248=>"111101101",
  25249=>"010000101",
  25250=>"000101101",
  25251=>"111100000",
  25252=>"110000111",
  25253=>"111110000",
  25254=>"001001000",
  25255=>"010000001",
  25256=>"111100000",
  25257=>"000010000",
  25258=>"010010000",
  25259=>"000000010",
  25260=>"000000000",
  25261=>"001000000",
  25262=>"110001000",
  25263=>"111111010",
  25264=>"001100111",
  25265=>"110111111",
  25266=>"000000101",
  25267=>"000110100",
  25268=>"111111111",
  25269=>"000000000",
  25270=>"101111011",
  25271=>"101111101",
  25272=>"000000000",
  25273=>"000110110",
  25274=>"110000010",
  25275=>"110110100",
  25276=>"101101101",
  25277=>"010001111",
  25278=>"001001110",
  25279=>"111111111",
  25280=>"000111001",
  25281=>"000111111",
  25282=>"111010001",
  25283=>"001000000",
  25284=>"000000000",
  25285=>"100100001",
  25286=>"110010011",
  25287=>"010010010",
  25288=>"001000111",
  25289=>"001111000",
  25290=>"111110111",
  25291=>"000001111",
  25292=>"111000001",
  25293=>"100111110",
  25294=>"111010001",
  25295=>"111101111",
  25296=>"000001111",
  25297=>"110010010",
  25298=>"111001011",
  25299=>"001110111",
  25300=>"110101001",
  25301=>"111110001",
  25302=>"011000000",
  25303=>"110010101",
  25304=>"000000000",
  25305=>"101001010",
  25306=>"111111101",
  25307=>"000111010",
  25308=>"100001000",
  25309=>"011111000",
  25310=>"111111110",
  25311=>"011111000",
  25312=>"000010110",
  25313=>"000000101",
  25314=>"000110111",
  25315=>"110100000",
  25316=>"010000000",
  25317=>"101111110",
  25318=>"011010111",
  25319=>"000100100",
  25320=>"100111111",
  25321=>"000101111",
  25322=>"001000011",
  25323=>"010111010",
  25324=>"111110000",
  25325=>"011111111",
  25326=>"000110000",
  25327=>"000000110",
  25328=>"110010000",
  25329=>"001001001",
  25330=>"110110000",
  25331=>"110100110",
  25332=>"001000110",
  25333=>"111111000",
  25334=>"000010001",
  25335=>"100110000",
  25336=>"000100101",
  25337=>"000001000",
  25338=>"111010111",
  25339=>"000101000",
  25340=>"000000111",
  25341=>"011111111",
  25342=>"111000000",
  25343=>"000000000",
  25344=>"000110110",
  25345=>"110100000",
  25346=>"001000100",
  25347=>"101100000",
  25348=>"111111111",
  25349=>"111111000",
  25350=>"000011011",
  25351=>"000000000",
  25352=>"100000001",
  25353=>"101000100",
  25354=>"111111111",
  25355=>"010101100",
  25356=>"111110100",
  25357=>"111110000",
  25358=>"110110100",
  25359=>"000000000",
  25360=>"100111111",
  25361=>"111111111",
  25362=>"000011111",
  25363=>"110010000",
  25364=>"100010010",
  25365=>"111111111",
  25366=>"000000001",
  25367=>"111111111",
  25368=>"101010011",
  25369=>"000000110",
  25370=>"111110000",
  25371=>"010100010",
  25372=>"000000001",
  25373=>"001000000",
  25374=>"000001111",
  25375=>"000010000",
  25376=>"001000000",
  25377=>"000010000",
  25378=>"000011100",
  25379=>"010000010",
  25380=>"001010111",
  25381=>"011011011",
  25382=>"000110010",
  25383=>"000000101",
  25384=>"000000100",
  25385=>"010100111",
  25386=>"010011011",
  25387=>"000010000",
  25388=>"011111110",
  25389=>"111010000",
  25390=>"111110011",
  25391=>"000000000",
  25392=>"000000000",
  25393=>"000110110",
  25394=>"011000000",
  25395=>"010111101",
  25396=>"111101111",
  25397=>"111101010",
  25398=>"001001000",
  25399=>"010011101",
  25400=>"111110110",
  25401=>"111010000",
  25402=>"001000000",
  25403=>"000000000",
  25404=>"001100001",
  25405=>"111011111",
  25406=>"000100000",
  25407=>"011011011",
  25408=>"110000111",
  25409=>"101000111",
  25410=>"111000000",
  25411=>"010001001",
  25412=>"111111110",
  25413=>"000000000",
  25414=>"000000001",
  25415=>"101101001",
  25416=>"110000010",
  25417=>"000111111",
  25418=>"100100101",
  25419=>"011101111",
  25420=>"001101111",
  25421=>"100010110",
  25422=>"001111111",
  25423=>"011111111",
  25424=>"111100000",
  25425=>"100101111",
  25426=>"000010000",
  25427=>"000110000",
  25428=>"011000100",
  25429=>"010011001",
  25430=>"000110011",
  25431=>"000000101",
  25432=>"111111101",
  25433=>"011011011",
  25434=>"011010000",
  25435=>"100111111",
  25436=>"000101101",
  25437=>"001100100",
  25438=>"000011010",
  25439=>"110101001",
  25440=>"111101000",
  25441=>"010000100",
  25442=>"000000110",
  25443=>"001011010",
  25444=>"011011011",
  25445=>"010100001",
  25446=>"000000111",
  25447=>"011111111",
  25448=>"000000000",
  25449=>"111011111",
  25450=>"110010001",
  25451=>"000111100",
  25452=>"010011111",
  25453=>"101111010",
  25454=>"000000000",
  25455=>"111111111",
  25456=>"111011110",
  25457=>"111111111",
  25458=>"001000000",
  25459=>"000110100",
  25460=>"010111101",
  25461=>"000000000",
  25462=>"111111101",
  25463=>"001000000",
  25464=>"101000000",
  25465=>"111111111",
  25466=>"000101111",
  25467=>"111111101",
  25468=>"000000000",
  25469=>"001001001",
  25470=>"001000100",
  25471=>"101100110",
  25472=>"000010010",
  25473=>"000010000",
  25474=>"101100100",
  25475=>"000111111",
  25476=>"000010000",
  25477=>"101000101",
  25478=>"101100001",
  25479=>"100000110",
  25480=>"100110111",
  25481=>"101101011",
  25482=>"111111110",
  25483=>"000101111",
  25484=>"111111100",
  25485=>"000101111",
  25486=>"100111111",
  25487=>"000000001",
  25488=>"001011011",
  25489=>"111111100",
  25490=>"101101111",
  25491=>"100100100",
  25492=>"000100110",
  25493=>"101101111",
  25494=>"111111111",
  25495=>"110110110",
  25496=>"010011111",
  25497=>"100000000",
  25498=>"101100101",
  25499=>"000000000",
  25500=>"110110111",
  25501=>"000000000",
  25502=>"100111111",
  25503=>"111111111",
  25504=>"011000111",
  25505=>"001111111",
  25506=>"111101111",
  25507=>"111010111",
  25508=>"000010000",
  25509=>"011011011",
  25510=>"000000001",
  25511=>"011111111",
  25512=>"100001000",
  25513=>"101000000",
  25514=>"001000000",
  25515=>"000110000",
  25516=>"100010000",
  25517=>"000111111",
  25518=>"000101111",
  25519=>"111000001",
  25520=>"100000100",
  25521=>"100110110",
  25522=>"000000000",
  25523=>"011011001",
  25524=>"010111111",
  25525=>"001100000",
  25526=>"011110000",
  25527=>"100111101",
  25528=>"100101000",
  25529=>"001001001",
  25530=>"001100101",
  25531=>"010000111",
  25532=>"101111111",
  25533=>"101001001",
  25534=>"100100100",
  25535=>"111110010",
  25536=>"000000010",
  25537=>"101000000",
  25538=>"110011001",
  25539=>"000000100",
  25540=>"111101111",
  25541=>"011001011",
  25542=>"001000100",
  25543=>"101001101",
  25544=>"000010000",
  25545=>"111111000",
  25546=>"110011011",
  25547=>"101000000",
  25548=>"100110111",
  25549=>"000000100",
  25550=>"010111101",
  25551=>"100111011",
  25552=>"010111010",
  25553=>"111110110",
  25554=>"111000101",
  25555=>"111110111",
  25556=>"001111111",
  25557=>"010001011",
  25558=>"111011010",
  25559=>"100011010",
  25560=>"100010111",
  25561=>"000011111",
  25562=>"000110100",
  25563=>"000000000",
  25564=>"000110010",
  25565=>"010000000",
  25566=>"010000001",
  25567=>"000001001",
  25568=>"011100011",
  25569=>"010101101",
  25570=>"000111111",
  25571=>"000111011",
  25572=>"001000000",
  25573=>"010111010",
  25574=>"110000101",
  25575=>"000110110",
  25576=>"000101111",
  25577=>"000100000",
  25578=>"011111100",
  25579=>"011001100",
  25580=>"111100000",
  25581=>"110100111",
  25582=>"010000011",
  25583=>"000000100",
  25584=>"101111111",
  25585=>"110100111",
  25586=>"000000010",
  25587=>"000010010",
  25588=>"000001011",
  25589=>"011111000",
  25590=>"000001000",
  25591=>"001100000",
  25592=>"000000000",
  25593=>"000111010",
  25594=>"110000000",
  25595=>"000111111",
  25596=>"000000000",
  25597=>"000101101",
  25598=>"000110110",
  25599=>"000111011",
  25600=>"000100101",
  25601=>"101111111",
  25602=>"111100100",
  25603=>"000010011",
  25604=>"111101101",
  25605=>"000111100",
  25606=>"011111101",
  25607=>"100110100",
  25608=>"000000001",
  25609=>"111101100",
  25610=>"101101100",
  25611=>"101100100",
  25612=>"000000111",
  25613=>"000000111",
  25614=>"111100100",
  25615=>"111010000",
  25616=>"000000100",
  25617=>"111000000",
  25618=>"011111000",
  25619=>"111011000",
  25620=>"111011111",
  25621=>"111100100",
  25622=>"101000111",
  25623=>"001001000",
  25624=>"000100000",
  25625=>"000000000",
  25626=>"000000111",
  25627=>"111000100",
  25628=>"000100000",
  25629=>"011100101",
  25630=>"000011111",
  25631=>"101100100",
  25632=>"000000000",
  25633=>"111011011",
  25634=>"011000100",
  25635=>"000011011",
  25636=>"000001110",
  25637=>"000000100",
  25638=>"100011011",
  25639=>"010010000",
  25640=>"001011011",
  25641=>"001001100",
  25642=>"111110101",
  25643=>"000011010",
  25644=>"100001011",
  25645=>"000010011",
  25646=>"000000111",
  25647=>"111010110",
  25648=>"001000101",
  25649=>"111001001",
  25650=>"000010011",
  25651=>"001110100",
  25652=>"010000001",
  25653=>"101111111",
  25654=>"000010110",
  25655=>"111101101",
  25656=>"011011101",
  25657=>"111101100",
  25658=>"111001100",
  25659=>"111000100",
  25660=>"011000000",
  25661=>"010111111",
  25662=>"111100000",
  25663=>"000001111",
  25664=>"000010000",
  25665=>"000000101",
  25666=>"111111110",
  25667=>"000100111",
  25668=>"111101111",
  25669=>"111100100",
  25670=>"000111111",
  25671=>"000011010",
  25672=>"000011111",
  25673=>"110100111",
  25674=>"110100101",
  25675=>"111100101",
  25676=>"111100000",
  25677=>"010110011",
  25678=>"111000010",
  25679=>"111011100",
  25680=>"111101000",
  25681=>"000010010",
  25682=>"111000111",
  25683=>"000011001",
  25684=>"111100100",
  25685=>"011011011",
  25686=>"011011011",
  25687=>"100100101",
  25688=>"100000100",
  25689=>"000000000",
  25690=>"111110000",
  25691=>"001011111",
  25692=>"001000111",
  25693=>"111100101",
  25694=>"100000011",
  25695=>"001000111",
  25696=>"000000011",
  25697=>"111111100",
  25698=>"011100100",
  25699=>"111101101",
  25700=>"111000011",
  25701=>"111111100",
  25702=>"000011011",
  25703=>"100001000",
  25704=>"010110111",
  25705=>"011111000",
  25706=>"100001000",
  25707=>"000101011",
  25708=>"000010111",
  25709=>"111000001",
  25710=>"000000101",
  25711=>"111000000",
  25712=>"110110111",
  25713=>"001011111",
  25714=>"110000000",
  25715=>"000000000",
  25716=>"100000011",
  25717=>"010101100",
  25718=>"011111100",
  25719=>"000000011",
  25720=>"000110011",
  25721=>"110011111",
  25722=>"101111111",
  25723=>"110011101",
  25724=>"110110010",
  25725=>"000010010",
  25726=>"110010010",
  25727=>"111100100",
  25728=>"000010101",
  25729=>"010111100",
  25730=>"000001001",
  25731=>"000000111",
  25732=>"010010100",
  25733=>"001011011",
  25734=>"000101001",
  25735=>"001000000",
  25736=>"010000101",
  25737=>"111111000",
  25738=>"001100100",
  25739=>"001011010",
  25740=>"100100011",
  25741=>"100101100",
  25742=>"111110100",
  25743=>"111000000",
  25744=>"011101011",
  25745=>"000000111",
  25746=>"011000000",
  25747=>"001011111",
  25748=>"001000000",
  25749=>"101100100",
  25750=>"111100100",
  25751=>"000010011",
  25752=>"001011001",
  25753=>"100100111",
  25754=>"000000011",
  25755=>"000000000",
  25756=>"111110111",
  25757=>"101111111",
  25758=>"001100110",
  25759=>"111101000",
  25760=>"000101001",
  25761=>"000000100",
  25762=>"000010101",
  25763=>"000000101",
  25764=>"111000110",
  25765=>"110100010",
  25766=>"000011111",
  25767=>"000011011",
  25768=>"110111000",
  25769=>"010110000",
  25770=>"000000100",
  25771=>"111101100",
  25772=>"000011011",
  25773=>"100000000",
  25774=>"101000000",
  25775=>"100010010",
  25776=>"110000000",
  25777=>"111001011",
  25778=>"111100110",
  25779=>"000010010",
  25780=>"010011011",
  25781=>"010011111",
  25782=>"000001011",
  25783=>"000010010",
  25784=>"110011000",
  25785=>"010000001",
  25786=>"000100100",
  25787=>"000010011",
  25788=>"111111111",
  25789=>"010000011",
  25790=>"000010001",
  25791=>"000101101",
  25792=>"001000100",
  25793=>"000000000",
  25794=>"100100111",
  25795=>"111101000",
  25796=>"111101101",
  25797=>"000110010",
  25798=>"100000000",
  25799=>"000010010",
  25800=>"010100000",
  25801=>"111100100",
  25802=>"000000000",
  25803=>"111101101",
  25804=>"111110100",
  25805=>"011010011",
  25806=>"011101100",
  25807=>"111000011",
  25808=>"111101000",
  25809=>"001000111",
  25810=>"000000010",
  25811=>"010100111",
  25812=>"111111110",
  25813=>"001001010",
  25814=>"011100100",
  25815=>"000000100",
  25816=>"001011011",
  25817=>"111100000",
  25818=>"001000100",
  25819=>"011000000",
  25820=>"000110101",
  25821=>"100100011",
  25822=>"111011111",
  25823=>"000000010",
  25824=>"111100100",
  25825=>"101100100",
  25826=>"111100000",
  25827=>"000000001",
  25828=>"000000000",
  25829=>"110000111",
  25830=>"111111000",
  25831=>"100000000",
  25832=>"011011011",
  25833=>"000000000",
  25834=>"101100001",
  25835=>"000011111",
  25836=>"000100111",
  25837=>"001000011",
  25838=>"000000000",
  25839=>"000000000",
  25840=>"001000000",
  25841=>"110001000",
  25842=>"000001101",
  25843=>"111010111",
  25844=>"000000110",
  25845=>"111111100",
  25846=>"011100000",
  25847=>"000011011",
  25848=>"011000001",
  25849=>"010111111",
  25850=>"000000001",
  25851=>"000000111",
  25852=>"111100100",
  25853=>"000000000",
  25854=>"000000001",
  25855=>"111111000",
  25856=>"011011101",
  25857=>"000000100",
  25858=>"101101101",
  25859=>"010111000",
  25860=>"011111010",
  25861=>"100000101",
  25862=>"010000011",
  25863=>"000001000",
  25864=>"000001110",
  25865=>"000010001",
  25866=>"000110111",
  25867=>"001001100",
  25868=>"000001111",
  25869=>"000001111",
  25870=>"111111001",
  25871=>"111110010",
  25872=>"000010111",
  25873=>"010010111",
  25874=>"100000110",
  25875=>"011010100",
  25876=>"000000000",
  25877=>"110010000",
  25878=>"000001100",
  25879=>"000000000",
  25880=>"000000010",
  25881=>"111000111",
  25882=>"000001011",
  25883=>"010011000",
  25884=>"000000000",
  25885=>"110010000",
  25886=>"101000111",
  25887=>"000000111",
  25888=>"111001101",
  25889=>"000000101",
  25890=>"100000010",
  25891=>"110000010",
  25892=>"001001011",
  25893=>"100010100",
  25894=>"000000011",
  25895=>"000001111",
  25896=>"010010000",
  25897=>"101001000",
  25898=>"101000110",
  25899=>"001000010",
  25900=>"111111111",
  25901=>"111101100",
  25902=>"011001000",
  25903=>"011001001",
  25904=>"000000000",
  25905=>"001101111",
  25906=>"010000100",
  25907=>"110111111",
  25908=>"101001111",
  25909=>"111111100",
  25910=>"000000100",
  25911=>"000100000",
  25912=>"000101001",
  25913=>"111111000",
  25914=>"000000110",
  25915=>"011110001",
  25916=>"001001001",
  25917=>"111111011",
  25918=>"001010000",
  25919=>"011011001",
  25920=>"000010111",
  25921=>"010000000",
  25922=>"100000111",
  25923=>"000000110",
  25924=>"000000000",
  25925=>"000000110",
  25926=>"100011010",
  25927=>"010010111",
  25928=>"111100101",
  25929=>"010010000",
  25930=>"010000000",
  25931=>"000100100",
  25932=>"000100000",
  25933=>"111111110",
  25934=>"101010000",
  25935=>"101100001",
  25936=>"101000111",
  25937=>"111010010",
  25938=>"001000100",
  25939=>"001001001",
  25940=>"001101001",
  25941=>"100001101",
  25942=>"111111100",
  25943=>"101101110",
  25944=>"101001101",
  25945=>"110110110",
  25946=>"000000101",
  25947=>"000010111",
  25948=>"000000000",
  25949=>"001000001",
  25950=>"000111111",
  25951=>"000100001",
  25952=>"000001111",
  25953=>"110000101",
  25954=>"101111111",
  25955=>"000000100",
  25956=>"111111110",
  25957=>"011000001",
  25958=>"111011001",
  25959=>"000000010",
  25960=>"110111000",
  25961=>"111111100",
  25962=>"000001111",
  25963=>"000000110",
  25964=>"111111111",
  25965=>"110111010",
  25966=>"000100000",
  25967=>"111111101",
  25968=>"101111101",
  25969=>"001000100",
  25970=>"000000001",
  25971=>"001000000",
  25972=>"010000000",
  25973=>"101100100",
  25974=>"000010110",
  25975=>"100111111",
  25976=>"000000011",
  25977=>"110010000",
  25978=>"001101111",
  25979=>"111111100",
  25980=>"111111001",
  25981=>"100100000",
  25982=>"010010111",
  25983=>"001000000",
  25984=>"010100101",
  25985=>"101000010",
  25986=>"010010010",
  25987=>"110000111",
  25988=>"111010010",
  25989=>"010111111",
  25990=>"001001001",
  25991=>"001011000",
  25992=>"111111101",
  25993=>"110010101",
  25994=>"010000000",
  25995=>"010010011",
  25996=>"000010001",
  25997=>"001011001",
  25998=>"110010110",
  25999=>"000000001",
  26000=>"111111101",
  26001=>"111101000",
  26002=>"011000001",
  26003=>"001000100",
  26004=>"011111111",
  26005=>"000000001",
  26006=>"011101111",
  26007=>"000000000",
  26008=>"010111111",
  26009=>"110111111",
  26010=>"010111000",
  26011=>"000000010",
  26012=>"000000000",
  26013=>"011111111",
  26014=>"000000000",
  26015=>"111011000",
  26016=>"101101101",
  26017=>"000110111",
  26018=>"111101101",
  26019=>"000000001",
  26020=>"000000101",
  26021=>"110000000",
  26022=>"101001111",
  26023=>"011111001",
  26024=>"111010110",
  26025=>"001010011",
  26026=>"100000000",
  26027=>"000010111",
  26028=>"110111111",
  26029=>"001001000",
  26030=>"000100101",
  26031=>"000010010",
  26032=>"011000011",
  26033=>"011001001",
  26034=>"010010010",
  26035=>"001001001",
  26036=>"011101001",
  26037=>"010010011",
  26038=>"011010000",
  26039=>"010000001",
  26040=>"100100110",
  26041=>"110110100",
  26042=>"000111110",
  26043=>"000100010",
  26044=>"111111000",
  26045=>"110111010",
  26046=>"101100101",
  26047=>"010010000",
  26048=>"001001101",
  26049=>"010010000",
  26050=>"010000101",
  26051=>"111111110",
  26052=>"010011000",
  26053=>"110110111",
  26054=>"111100000",
  26055=>"110010110",
  26056=>"101000011",
  26057=>"000101111",
  26058=>"110110011",
  26059=>"111111111",
  26060=>"000000000",
  26061=>"111100100",
  26062=>"000111111",
  26063=>"000011010",
  26064=>"011000000",
  26065=>"110101111",
  26066=>"000000100",
  26067=>"010111110",
  26068=>"001000111",
  26069=>"100100100",
  26070=>"111101000",
  26071=>"110101000",
  26072=>"111101101",
  26073=>"100000111",
  26074=>"101101001",
  26075=>"000010010",
  26076=>"000001001",
  26077=>"000000010",
  26078=>"101001101",
  26079=>"000000100",
  26080=>"000000111",
  26081=>"000100000",
  26082=>"000010110",
  26083=>"101111110",
  26084=>"001000101",
  26085=>"010110111",
  26086=>"010010010",
  26087=>"010011010",
  26088=>"000000000",
  26089=>"000000000",
  26090=>"000001111",
  26091=>"101110111",
  26092=>"101000101",
  26093=>"000000000",
  26094=>"001110000",
  26095=>"001111010",
  26096=>"111111000",
  26097=>"011101111",
  26098=>"100001100",
  26099=>"001001101",
  26100=>"110110110",
  26101=>"000000101",
  26102=>"000000000",
  26103=>"000000001",
  26104=>"000011011",
  26105=>"010000100",
  26106=>"111010010",
  26107=>"000101000",
  26108=>"110110110",
  26109=>"000000001",
  26110=>"111101110",
  26111=>"011111111",
  26112=>"111000000",
  26113=>"000010111",
  26114=>"000000110",
  26115=>"111000101",
  26116=>"110111111",
  26117=>"110100101",
  26118=>"000001101",
  26119=>"000000100",
  26120=>"011000000",
  26121=>"000100000",
  26122=>"000011001",
  26123=>"000000000",
  26124=>"110000000",
  26125=>"101011011",
  26126=>"100001000",
  26127=>"111010110",
  26128=>"000101011",
  26129=>"010111111",
  26130=>"111000000",
  26131=>"000011111",
  26132=>"010100110",
  26133=>"111111101",
  26134=>"000111011",
  26135=>"101011110",
  26136=>"111000000",
  26137=>"111111111",
  26138=>"111001000",
  26139=>"000000111",
  26140=>"000000111",
  26141=>"101011000",
  26142=>"100000001",
  26143=>"111010010",
  26144=>"000111111",
  26145=>"111100000",
  26146=>"000000010",
  26147=>"011001111",
  26148=>"011101101",
  26149=>"000000000",
  26150=>"111101101",
  26151=>"101001110",
  26152=>"111101001",
  26153=>"000010111",
  26154=>"000101101",
  26155=>"000010000",
  26156=>"000000111",
  26157=>"001100000",
  26158=>"001000100",
  26159=>"101100110",
  26160=>"011111110",
  26161=>"111111001",
  26162=>"000111111",
  26163=>"111011001",
  26164=>"000111110",
  26165=>"000000001",
  26166=>"000011010",
  26167=>"111100100",
  26168=>"000010101",
  26169=>"001001001",
  26170=>"111001000",
  26171=>"000011111",
  26172=>"001100101",
  26173=>"101111010",
  26174=>"010000000",
  26175=>"010110011",
  26176=>"001110010",
  26177=>"011000000",
  26178=>"110111000",
  26179=>"111000100",
  26180=>"111111101",
  26181=>"100010111",
  26182=>"000001101",
  26183=>"101111111",
  26184=>"110001001",
  26185=>"011000111",
  26186=>"111000100",
  26187=>"111101011",
  26188=>"000000010",
  26189=>"110001100",
  26190=>"011111111",
  26191=>"000010110",
  26192=>"010110110",
  26193=>"100111110",
  26194=>"001000101",
  26195=>"010011000",
  26196=>"000000100",
  26197=>"000100101",
  26198=>"001001100",
  26199=>"000000101",
  26200=>"000010101",
  26201=>"000000011",
  26202=>"010011001",
  26203=>"111011001",
  26204=>"100000000",
  26205=>"111101001",
  26206=>"011111111",
  26207=>"111001001",
  26208=>"000000000",
  26209=>"111101000",
  26210=>"111101000",
  26211=>"100101011",
  26212=>"111110100",
  26213=>"000011111",
  26214=>"110001011",
  26215=>"011000000",
  26216=>"111001000",
  26217=>"000110001",
  26218=>"000011111",
  26219=>"111011000",
  26220=>"111110000",
  26221=>"111000000",
  26222=>"111001100",
  26223=>"000101111",
  26224=>"010011101",
  26225=>"000000000",
  26226=>"000110011",
  26227=>"110110100",
  26228=>"110111111",
  26229=>"111000101",
  26230=>"111000000",
  26231=>"000001010",
  26232=>"000000111",
  26233=>"000000111",
  26234=>"001000000",
  26235=>"111111101",
  26236=>"100100111",
  26237=>"111111100",
  26238=>"000111010",
  26239=>"111001000",
  26240=>"010111000",
  26241=>"000111000",
  26242=>"000000000",
  26243=>"101111010",
  26244=>"011101000",
  26245=>"101000000",
  26246=>"100000000",
  26247=>"111000000",
  26248=>"110100101",
  26249=>"101010110",
  26250=>"011000101",
  26251=>"101111111",
  26252=>"001000100",
  26253=>"100111101",
  26254=>"010000000",
  26255=>"000000110",
  26256=>"011011011",
  26257=>"111001000",
  26258=>"101011011",
  26259=>"111011011",
  26260=>"101110010",
  26261=>"011000000",
  26262=>"011000000",
  26263=>"000100000",
  26264=>"010000111",
  26265=>"000000111",
  26266=>"111111111",
  26267=>"000000010",
  26268=>"111101101",
  26269=>"011100001",
  26270=>"110011000",
  26271=>"000000010",
  26272=>"001100000",
  26273=>"000011010",
  26274=>"111111001",
  26275=>"000000110",
  26276=>"100000000",
  26277=>"110101001",
  26278=>"000010001",
  26279=>"010000000",
  26280=>"000000010",
  26281=>"000101100",
  26282=>"111000000",
  26283=>"000111110",
  26284=>"001101010",
  26285=>"000000000",
  26286=>"001011011",
  26287=>"011101000",
  26288=>"000001100",
  26289=>"111011001",
  26290=>"011111100",
  26291=>"010100110",
  26292=>"010111111",
  26293=>"000111111",
  26294=>"000100111",
  26295=>"001011111",
  26296=>"000100100",
  26297=>"011011000",
  26298=>"000100000",
  26299=>"110000000",
  26300=>"110000000",
  26301=>"111111000",
  26302=>"010001001",
  26303=>"000110111",
  26304=>"101101000",
  26305=>"001000000",
  26306=>"111101111",
  26307=>"011011000",
  26308=>"111000000",
  26309=>"101100111",
  26310=>"000000100",
  26311=>"011001011",
  26312=>"111101100",
  26313=>"000100110",
  26314=>"101111110",
  26315=>"010110100",
  26316=>"000001111",
  26317=>"001001110",
  26318=>"000111010",
  26319=>"111100000",
  26320=>"000000110",
  26321=>"011011001",
  26322=>"011100100",
  26323=>"111111010",
  26324=>"111011111",
  26325=>"100000100",
  26326=>"111111101",
  26327=>"111111001",
  26328=>"000111111",
  26329=>"111111000",
  26330=>"100001101",
  26331=>"111100000",
  26332=>"000111111",
  26333=>"100000000",
  26334=>"000000111",
  26335=>"111101000",
  26336=>"111100101",
  26337=>"111111001",
  26338=>"000100100",
  26339=>"011001101",
  26340=>"000000101",
  26341=>"000101111",
  26342=>"000001111",
  26343=>"100100100",
  26344=>"111111101",
  26345=>"100111111",
  26346=>"100010110",
  26347=>"100000011",
  26348=>"101100100",
  26349=>"000000100",
  26350=>"110100000",
  26351=>"000111010",
  26352=>"000110011",
  26353=>"001011101",
  26354=>"000000101",
  26355=>"010111111",
  26356=>"000000100",
  26357=>"101000000",
  26358=>"111100000",
  26359=>"000101111",
  26360=>"111110111",
  26361=>"111011101",
  26362=>"001111001",
  26363=>"000101101",
  26364=>"011110000",
  26365=>"100111010",
  26366=>"000001111",
  26367=>"010000100",
  26368=>"110000000",
  26369=>"110000000",
  26370=>"110111010",
  26371=>"111101111",
  26372=>"001001001",
  26373=>"100000000",
  26374=>"110110010",
  26375=>"000000001",
  26376=>"000110111",
  26377=>"111011001",
  26378=>"111000110",
  26379=>"101000001",
  26380=>"000000000",
  26381=>"000010000",
  26382=>"110010001",
  26383=>"011111111",
  26384=>"000000110",
  26385=>"110111110",
  26386=>"000000000",
  26387=>"000111111",
  26388=>"010111110",
  26389=>"111001000",
  26390=>"100001001",
  26391=>"010110011",
  26392=>"000000000",
  26393=>"111100010",
  26394=>"100101110",
  26395=>"100000100",
  26396=>"000000000",
  26397=>"100000000",
  26398=>"010000000",
  26399=>"101101101",
  26400=>"100000111",
  26401=>"000000000",
  26402=>"000111001",
  26403=>"111000101",
  26404=>"111110000",
  26405=>"000000000",
  26406=>"011111010",
  26407=>"111110111",
  26408=>"111111001",
  26409=>"111111001",
  26410=>"110111110",
  26411=>"001001001",
  26412=>"111001001",
  26413=>"100100000",
  26414=>"000000000",
  26415=>"000000000",
  26416=>"000000001",
  26417=>"100001001",
  26418=>"000000000",
  26419=>"111101111",
  26420=>"010000000",
  26421=>"111111110",
  26422=>"111011011",
  26423=>"000000000",
  26424=>"000000000",
  26425=>"101000000",
  26426=>"010000100",
  26427=>"111111001",
  26428=>"001101100",
  26429=>"000101000",
  26430=>"101100001",
  26431=>"011011011",
  26432=>"111111111",
  26433=>"000000010",
  26434=>"100100000",
  26435=>"000100100",
  26436=>"110111111",
  26437=>"101000101",
  26438=>"000111111",
  26439=>"011111111",
  26440=>"000101001",
  26441=>"110000010",
  26442=>"111101001",
  26443=>"110110010",
  26444=>"101101001",
  26445=>"011011000",
  26446=>"110000000",
  26447=>"101110000",
  26448=>"001011001",
  26449=>"010000000",
  26450=>"001000111",
  26451=>"001000101",
  26452=>"000000000",
  26453=>"100100100",
  26454=>"100100100",
  26455=>"000001111",
  26456=>"001111111",
  26457=>"011011001",
  26458=>"100110110",
  26459=>"111111111",
  26460=>"001101101",
  26461=>"110000000",
  26462=>"010110110",
  26463=>"000001011",
  26464=>"001111111",
  26465=>"001101000",
  26466=>"000001101",
  26467=>"100111101",
  26468=>"101111100",
  26469=>"001100000",
  26470=>"011001100",
  26471=>"110000001",
  26472=>"110000111",
  26473=>"000000011",
  26474=>"001000101",
  26475=>"001000000",
  26476=>"011000110",
  26477=>"111111110",
  26478=>"000000000",
  26479=>"111000000",
  26480=>"100110111",
  26481=>"001111000",
  26482=>"111110110",
  26483=>"000000000",
  26484=>"000000001",
  26485=>"011000000",
  26486=>"111111100",
  26487=>"110111010",
  26488=>"111101101",
  26489=>"111001001",
  26490=>"111000111",
  26491=>"000001111",
  26492=>"001000110",
  26493=>"000000001",
  26494=>"010000000",
  26495=>"000000101",
  26496=>"010010000",
  26497=>"000000000",
  26498=>"111000010",
  26499=>"111111100",
  26500=>"101000000",
  26501=>"111111011",
  26502=>"000000010",
  26503=>"001110011",
  26504=>"011011011",
  26505=>"110010000",
  26506=>"011101000",
  26507=>"011111111",
  26508=>"111110111",
  26509=>"000001111",
  26510=>"000000111",
  26511=>"100000111",
  26512=>"001011011",
  26513=>"000100111",
  26514=>"100000000",
  26515=>"001111111",
  26516=>"000000111",
  26517=>"001000110",
  26518=>"100100000",
  26519=>"100100000",
  26520=>"000000000",
  26521=>"001101000",
  26522=>"110100111",
  26523=>"000000100",
  26524=>"100100000",
  26525=>"111111011",
  26526=>"010000001",
  26527=>"111000011",
  26528=>"111111111",
  26529=>"111111000",
  26530=>"011111111",
  26531=>"111111111",
  26532=>"011000000",
  26533=>"110110110",
  26534=>"001001001",
  26535=>"111111010",
  26536=>"111111111",
  26537=>"001000111",
  26538=>"000001111",
  26539=>"111000000",
  26540=>"001111101",
  26541=>"101101100",
  26542=>"101001000",
  26543=>"000000101",
  26544=>"000101101",
  26545=>"111100110",
  26546=>"000000000",
  26547=>"001000000",
  26548=>"111000000",
  26549=>"111111011",
  26550=>"111111110",
  26551=>"111111101",
  26552=>"100000000",
  26553=>"000000100",
  26554=>"101001000",
  26555=>"000100111",
  26556=>"010000000",
  26557=>"101101111",
  26558=>"001111110",
  26559=>"010010010",
  26560=>"000111111",
  26561=>"011111010",
  26562=>"010000010",
  26563=>"101100100",
  26564=>"010000000",
  26565=>"100100000",
  26566=>"000000000",
  26567=>"100000000",
  26568=>"111111101",
  26569=>"111111111",
  26570=>"111111011",
  26571=>"111011111",
  26572=>"111111101",
  26573=>"100111011",
  26574=>"000010010",
  26575=>"000000000",
  26576=>"101111000",
  26577=>"011000000",
  26578=>"100000000",
  26579=>"100000100",
  26580=>"001000101",
  26581=>"001000000",
  26582=>"001001101",
  26583=>"010000011",
  26584=>"000000000",
  26585=>"111001111",
  26586=>"110110110",
  26587=>"000000011",
  26588=>"101100001",
  26589=>"101000111",
  26590=>"111111110",
  26591=>"000000000",
  26592=>"111101000",
  26593=>"000000000",
  26594=>"000001101",
  26595=>"110110100",
  26596=>"000000100",
  26597=>"010010111",
  26598=>"111001111",
  26599=>"111111000",
  26600=>"011010000",
  26601=>"101100001",
  26602=>"100000101",
  26603=>"000111111",
  26604=>"000110000",
  26605=>"001001001",
  26606=>"000000000",
  26607=>"000000111",
  26608=>"000000000",
  26609=>"001001011",
  26610=>"000000111",
  26611=>"011101001",
  26612=>"011011001",
  26613=>"110111111",
  26614=>"000000000",
  26615=>"000000111",
  26616=>"010010111",
  26617=>"010000000",
  26618=>"111000000",
  26619=>"000000000",
  26620=>"011111100",
  26621=>"100000111",
  26622=>"111110110",
  26623=>"000000000",
  26624=>"111100110",
  26625=>"001011000",
  26626=>"111000000",
  26627=>"111010101",
  26628=>"110100110",
  26629=>"111111111",
  26630=>"111100100",
  26631=>"000001000",
  26632=>"000001001",
  26633=>"111001011",
  26634=>"000001000",
  26635=>"100000000",
  26636=>"110111111",
  26637=>"001101000",
  26638=>"110100000",
  26639=>"111111010",
  26640=>"110100010",
  26641=>"000000001",
  26642=>"100000000",
  26643=>"011111000",
  26644=>"000010000",
  26645=>"000000001",
  26646=>"111011000",
  26647=>"011111000",
  26648=>"101000101",
  26649=>"101000000",
  26650=>"011001111",
  26651=>"111000110",
  26652=>"001101101",
  26653=>"101000000",
  26654=>"111111111",
  26655=>"110000000",
  26656=>"111111110",
  26657=>"111111101",
  26658=>"001100000",
  26659=>"010111010",
  26660=>"100110010",
  26661=>"011001101",
  26662=>"000111111",
  26663=>"000001000",
  26664=>"000111010",
  26665=>"111001111",
  26666=>"111000000",
  26667=>"101000001",
  26668=>"110100010",
  26669=>"001000000",
  26670=>"011111111",
  26671=>"111001001",
  26672=>"011011000",
  26673=>"010111111",
  26674=>"101101010",
  26675=>"111101001",
  26676=>"101000000",
  26677=>"111001111",
  26678=>"111111111",
  26679=>"000000000",
  26680=>"010111001",
  26681=>"000000100",
  26682=>"000011000",
  26683=>"111000010",
  26684=>"001000000",
  26685=>"100111111",
  26686=>"111000010",
  26687=>"000000100",
  26688=>"101111000",
  26689=>"000001110",
  26690=>"111111000",
  26691=>"001000111",
  26692=>"000111011",
  26693=>"000101111",
  26694=>"011111010",
  26695=>"100101000",
  26696=>"101111010",
  26697=>"100000000",
  26698=>"011101111",
  26699=>"000000000",
  26700=>"000000111",
  26701=>"011110111",
  26702=>"001111111",
  26703=>"000000111",
  26704=>"000101001",
  26705=>"111111111",
  26706=>"000001010",
  26707=>"000110000",
  26708=>"000000000",
  26709=>"111011010",
  26710=>"011011001",
  26711=>"000000000",
  26712=>"011111000",
  26713=>"001111010",
  26714=>"011001000",
  26715=>"010001011",
  26716=>"111111011",
  26717=>"000110000",
  26718=>"101111101",
  26719=>"100100111",
  26720=>"100000101",
  26721=>"010101011",
  26722=>"000100101",
  26723=>"010000000",
  26724=>"111011001",
  26725=>"010000001",
  26726=>"111101101",
  26727=>"111000111",
  26728=>"111111100",
  26729=>"011111111",
  26730=>"000000111",
  26731=>"110101111",
  26732=>"111111111",
  26733=>"011011001",
  26734=>"101100101",
  26735=>"000000111",
  26736=>"000110111",
  26737=>"000011111",
  26738=>"011111111",
  26739=>"111101000",
  26740=>"000111111",
  26741=>"111100111",
  26742=>"011101000",
  26743=>"111101111",
  26744=>"001000000",
  26745=>"010110100",
  26746=>"000000000",
  26747=>"010110011",
  26748=>"000011000",
  26749=>"100001000",
  26750=>"001111110",
  26751=>"000000000",
  26752=>"010111101",
  26753=>"001000000",
  26754=>"001010111",
  26755=>"010111111",
  26756=>"000111011",
  26757=>"100000001",
  26758=>"000100001",
  26759=>"000000110",
  26760=>"000001111",
  26761=>"000000000",
  26762=>"110000000",
  26763=>"101011010",
  26764=>"000000000",
  26765=>"000000000",
  26766=>"000010010",
  26767=>"001000000",
  26768=>"111100011",
  26769=>"110000000",
  26770=>"000000110",
  26771=>"101000110",
  26772=>"100110000",
  26773=>"000111101",
  26774=>"111011000",
  26775=>"000100000",
  26776=>"101000000",
  26777=>"101111000",
  26778=>"010011011",
  26779=>"111000000",
  26780=>"010111000",
  26781=>"111011001",
  26782=>"111011000",
  26783=>"000000000",
  26784=>"011011110",
  26785=>"100010000",
  26786=>"000010011",
  26787=>"111111001",
  26788=>"101111100",
  26789=>"000000000",
  26790=>"001111000",
  26791=>"001000100",
  26792=>"000000111",
  26793=>"111011000",
  26794=>"111111000",
  26795=>"010010000",
  26796=>"101010000",
  26797=>"101101111",
  26798=>"000001001",
  26799=>"000000001",
  26800=>"000010000",
  26801=>"000110110",
  26802=>"101010011",
  26803=>"011010010",
  26804=>"111001000",
  26805=>"001000000",
  26806=>"110000101",
  26807=>"001100101",
  26808=>"110010000",
  26809=>"011001001",
  26810=>"010000100",
  26811=>"111111111",
  26812=>"000100001",
  26813=>"010000000",
  26814=>"100000000",
  26815=>"000100111",
  26816=>"000101100",
  26817=>"101000000",
  26818=>"010111000",
  26819=>"010110110",
  26820=>"000111011",
  26821=>"110011111",
  26822=>"010111001",
  26823=>"101000111",
  26824=>"010000010",
  26825=>"000000000",
  26826=>"011100110",
  26827=>"011111010",
  26828=>"100000000",
  26829=>"000110000",
  26830=>"110111000",
  26831=>"111111001",
  26832=>"000101101",
  26833=>"010110011",
  26834=>"011000000",
  26835=>"111010110",
  26836=>"101000000",
  26837=>"000011000",
  26838=>"110000000",
  26839=>"100001111",
  26840=>"000000000",
  26841=>"000000000",
  26842=>"110100011",
  26843=>"111111000",
  26844=>"111111000",
  26845=>"110000000",
  26846=>"100100000",
  26847=>"101111111",
  26848=>"000100000",
  26849=>"011111111",
  26850=>"110101111",
  26851=>"011001001",
  26852=>"000000000",
  26853=>"111111111",
  26854=>"000000000",
  26855=>"000110010",
  26856=>"000000100",
  26857=>"000000000",
  26858=>"000000000",
  26859=>"100000011",
  26860=>"011000000",
  26861=>"001101011",
  26862=>"000001000",
  26863=>"000000000",
  26864=>"000000110",
  26865=>"010100110",
  26866=>"101000111",
  26867=>"001111000",
  26868=>"011001011",
  26869=>"111110000",
  26870=>"000100111",
  26871=>"111111000",
  26872=>"000111010",
  26873=>"000111101",
  26874=>"000000000",
  26875=>"000000000",
  26876=>"111111011",
  26877=>"111111111",
  26878=>"000000000",
  26879=>"000000000",
  26880=>"100100110",
  26881=>"111101000",
  26882=>"100000111",
  26883=>"111101010",
  26884=>"000000000",
  26885=>"000000000",
  26886=>"011000100",
  26887=>"111111000",
  26888=>"000101110",
  26889=>"011011000",
  26890=>"110011001",
  26891=>"111000000",
  26892=>"010111000",
  26893=>"000000000",
  26894=>"110100010",
  26895=>"111111111",
  26896=>"010011000",
  26897=>"010010010",
  26898=>"010000000",
  26899=>"000100000",
  26900=>"010011000",
  26901=>"000000100",
  26902=>"000011111",
  26903=>"110111111",
  26904=>"111000000",
  26905=>"011011111",
  26906=>"101100000",
  26907=>"111111111",
  26908=>"000001111",
  26909=>"000000000",
  26910=>"001111110",
  26911=>"100000011",
  26912=>"111111100",
  26913=>"000000000",
  26914=>"100000000",
  26915=>"000000011",
  26916=>"000000001",
  26917=>"000001111",
  26918=>"000000010",
  26919=>"000011100",
  26920=>"000111111",
  26921=>"000101000",
  26922=>"010000100",
  26923=>"110010000",
  26924=>"111111001",
  26925=>"011001111",
  26926=>"100111010",
  26927=>"000000000",
  26928=>"111110001",
  26929=>"001000011",
  26930=>"101000111",
  26931=>"111010000",
  26932=>"000101000",
  26933=>"011111010",
  26934=>"100100000",
  26935=>"000000001",
  26936=>"111111010",
  26937=>"110100111",
  26938=>"110000000",
  26939=>"111101111",
  26940=>"001111101",
  26941=>"111000111",
  26942=>"100000000",
  26943=>"111100100",
  26944=>"111100010",
  26945=>"000110011",
  26946=>"000000111",
  26947=>"111000111",
  26948=>"000000000",
  26949=>"100011001",
  26950=>"111000111",
  26951=>"001000000",
  26952=>"010101110",
  26953=>"011111111",
  26954=>"100100100",
  26955=>"111111110",
  26956=>"000000000",
  26957=>"100110100",
  26958=>"001010100",
  26959=>"101100100",
  26960=>"000000000",
  26961=>"010111111",
  26962=>"111110101",
  26963=>"101000100",
  26964=>"000100111",
  26965=>"001000100",
  26966=>"101010000",
  26967=>"111011011",
  26968=>"000000010",
  26969=>"000000100",
  26970=>"001000000",
  26971=>"111011111",
  26972=>"000000110",
  26973=>"110010000",
  26974=>"000111100",
  26975=>"111011011",
  26976=>"111111111",
  26977=>"000000100",
  26978=>"000010010",
  26979=>"100000000",
  26980=>"100101111",
  26981=>"011011010",
  26982=>"000000000",
  26983=>"101000111",
  26984=>"101011111",
  26985=>"000000000",
  26986=>"010000000",
  26987=>"010111111",
  26988=>"111111101",
  26989=>"011111011",
  26990=>"000000000",
  26991=>"111000000",
  26992=>"000111001",
  26993=>"110000000",
  26994=>"000000000",
  26995=>"010011011",
  26996=>"010010000",
  26997=>"111001011",
  26998=>"100000001",
  26999=>"010111000",
  27000=>"100000001",
  27001=>"000011111",
  27002=>"101000101",
  27003=>"000011011",
  27004=>"001001101",
  27005=>"101001000",
  27006=>"111010010",
  27007=>"111100111",
  27008=>"101101100",
  27009=>"111111011",
  27010=>"000000011",
  27011=>"000101000",
  27012=>"011000000",
  27013=>"100000000",
  27014=>"100100101",
  27015=>"110000000",
  27016=>"010110100",
  27017=>"000100111",
  27018=>"011111001",
  27019=>"000001111",
  27020=>"000000011",
  27021=>"111010000",
  27022=>"000000111",
  27023=>"000000100",
  27024=>"110010010",
  27025=>"000000000",
  27026=>"001000000",
  27027=>"111100000",
  27028=>"000000100",
  27029=>"110110000",
  27030=>"111111000",
  27031=>"110100110",
  27032=>"010010001",
  27033=>"010000011",
  27034=>"010010000",
  27035=>"111000000",
  27036=>"111111111",
  27037=>"111111000",
  27038=>"100000000",
  27039=>"111111111",
  27040=>"000000010",
  27041=>"111110111",
  27042=>"111111111",
  27043=>"110011000",
  27044=>"101000000",
  27045=>"100000000",
  27046=>"010000110",
  27047=>"111101100",
  27048=>"000000000",
  27049=>"001101000",
  27050=>"000001000",
  27051=>"000000000",
  27052=>"011001010",
  27053=>"100100100",
  27054=>"110100101",
  27055=>"011010000",
  27056=>"111000001",
  27057=>"101101010",
  27058=>"000010111",
  27059=>"100000000",
  27060=>"111011000",
  27061=>"001000000",
  27062=>"000000000",
  27063=>"000001001",
  27064=>"010000011",
  27065=>"010011101",
  27066=>"000010011",
  27067=>"111111111",
  27068=>"001111111",
  27069=>"011111111",
  27070=>"111111001",
  27071=>"111010000",
  27072=>"011000100",
  27073=>"000000000",
  27074=>"111111111",
  27075=>"000000000",
  27076=>"000111111",
  27077=>"010111100",
  27078=>"011111011",
  27079=>"111000000",
  27080=>"011111010",
  27081=>"100000000",
  27082=>"000000100",
  27083=>"000000000",
  27084=>"111100101",
  27085=>"110110001",
  27086=>"100100100",
  27087=>"111111111",
  27088=>"111111111",
  27089=>"100011011",
  27090=>"100100101",
  27091=>"101111011",
  27092=>"101000100",
  27093=>"111111111",
  27094=>"100000000",
  27095=>"011010000",
  27096=>"000101101",
  27097=>"000110101",
  27098=>"000100101",
  27099=>"011010000",
  27100=>"100110101",
  27101=>"011111001",
  27102=>"101001000",
  27103=>"111111011",
  27104=>"000000000",
  27105=>"101011011",
  27106=>"111111111",
  27107=>"111011000",
  27108=>"000001100",
  27109=>"011011010",
  27110=>"000000000",
  27111=>"000100100",
  27112=>"000000011",
  27113=>"111111000",
  27114=>"110110110",
  27115=>"011011000",
  27116=>"001111011",
  27117=>"000000100",
  27118=>"100010111",
  27119=>"000000000",
  27120=>"101111111",
  27121=>"000000100",
  27122=>"000100111",
  27123=>"100100000",
  27124=>"001001111",
  27125=>"000000000",
  27126=>"011011010",
  27127=>"100010111",
  27128=>"000010000",
  27129=>"111111101",
  27130=>"000000000",
  27131=>"000110111",
  27132=>"000000111",
  27133=>"000011111",
  27134=>"001000001",
  27135=>"111111000",
  27136=>"000000100",
  27137=>"000000011",
  27138=>"111000000",
  27139=>"110000111",
  27140=>"000001001",
  27141=>"010011001",
  27142=>"001000001",
  27143=>"000001110",
  27144=>"000011001",
  27145=>"100000000",
  27146=>"000100011",
  27147=>"101101111",
  27148=>"000100101",
  27149=>"100110110",
  27150=>"000001000",
  27151=>"011011001",
  27152=>"100101000",
  27153=>"110111001",
  27154=>"111101000",
  27155=>"011111111",
  27156=>"011011101",
  27157=>"111111011",
  27158=>"111111001",
  27159=>"111111101",
  27160=>"001010000",
  27161=>"101000000",
  27162=>"100011011",
  27163=>"000000000",
  27164=>"011011010",
  27165=>"011010010",
  27166=>"110001000",
  27167=>"000000111",
  27168=>"000010110",
  27169=>"111010011",
  27170=>"001000111",
  27171=>"001111111",
  27172=>"000000000",
  27173=>"011011111",
  27174=>"100010010",
  27175=>"001000001",
  27176=>"001000010",
  27177=>"000000111",
  27178=>"101111101",
  27179=>"000001111",
  27180=>"000000111",
  27181=>"011111111",
  27182=>"010010111",
  27183=>"000000001",
  27184=>"111111110",
  27185=>"101101000",
  27186=>"000000101",
  27187=>"111001000",
  27188=>"000000010",
  27189=>"000111110",
  27190=>"011011110",
  27191=>"110111100",
  27192=>"111101000",
  27193=>"000001000",
  27194=>"000000101",
  27195=>"111111011",
  27196=>"000111011",
  27197=>"111010110",
  27198=>"000001000",
  27199=>"111011011",
  27200=>"111001000",
  27201=>"010111010",
  27202=>"111000100",
  27203=>"111011100",
  27204=>"111100111",
  27205=>"000000111",
  27206=>"000000000",
  27207=>"001000000",
  27208=>"000111110",
  27209=>"000001111",
  27210=>"000000000",
  27211=>"100111010",
  27212=>"011000000",
  27213=>"000111011",
  27214=>"001001000",
  27215=>"110111111",
  27216=>"011010111",
  27217=>"111010000",
  27218=>"011111111",
  27219=>"011011101",
  27220=>"001000110",
  27221=>"111111000",
  27222=>"000010010",
  27223=>"111000000",
  27224=>"000000000",
  27225=>"000000011",
  27226=>"000000111",
  27227=>"110000110",
  27228=>"100111000",
  27229=>"000001001",
  27230=>"111010111",
  27231=>"111101001",
  27232=>"110000000",
  27233=>"000010011",
  27234=>"110000000",
  27235=>"000001110",
  27236=>"000100111",
  27237=>"101000111",
  27238=>"000111111",
  27239=>"001110111",
  27240=>"001001111",
  27241=>"000000000",
  27242=>"110100101",
  27243=>"010000000",
  27244=>"010011010",
  27245=>"000000111",
  27246=>"000100101",
  27247=>"000000001",
  27248=>"011101111",
  27249=>"000000000",
  27250=>"110110011",
  27251=>"101110010",
  27252=>"111001010",
  27253=>"011000000",
  27254=>"000000000",
  27255=>"111110010",
  27256=>"000000100",
  27257=>"000101101",
  27258=>"000001000",
  27259=>"101100111",
  27260=>"011001100",
  27261=>"010100100",
  27262=>"111110110",
  27263=>"111001100",
  27264=>"111010000",
  27265=>"111111101",
  27266=>"010010000",
  27267=>"000011110",
  27268=>"011111101",
  27269=>"111111111",
  27270=>"110110110",
  27271=>"000100000",
  27272=>"100111011",
  27273=>"101110110",
  27274=>"000011110",
  27275=>"001000110",
  27276=>"111000000",
  27277=>"011110110",
  27278=>"111111000",
  27279=>"111101000",
  27280=>"001011101",
  27281=>"000100000",
  27282=>"001000000",
  27283=>"000001000",
  27284=>"000111000",
  27285=>"111100000",
  27286=>"111010111",
  27287=>"000011111",
  27288=>"000000111",
  27289=>"100000100",
  27290=>"111101001",
  27291=>"111100100",
  27292=>"111000010",
  27293=>"111110100",
  27294=>"111101011",
  27295=>"000001000",
  27296=>"000000001",
  27297=>"011000110",
  27298=>"000111101",
  27299=>"100100101",
  27300=>"100001100",
  27301=>"011010111",
  27302=>"111111111",
  27303=>"001010001",
  27304=>"111010111",
  27305=>"111101111",
  27306=>"111111101",
  27307=>"111101110",
  27308=>"000000110",
  27309=>"111001000",
  27310=>"000000011",
  27311=>"100100101",
  27312=>"011111100",
  27313=>"000001001",
  27314=>"000000000",
  27315=>"001101100",
  27316=>"000111111",
  27317=>"000110111",
  27318=>"000011000",
  27319=>"000001100",
  27320=>"000111111",
  27321=>"000001001",
  27322=>"011110110",
  27323=>"001101000",
  27324=>"000001010",
  27325=>"111111100",
  27326=>"100000001",
  27327=>"000111111",
  27328=>"000000000",
  27329=>"000111110",
  27330=>"011111111",
  27331=>"000000110",
  27332=>"001000000",
  27333=>"001010101",
  27334=>"000000000",
  27335=>"111000100",
  27336=>"000001101",
  27337=>"110010000",
  27338=>"011010000",
  27339=>"111100010",
  27340=>"000000000",
  27341=>"100100101",
  27342=>"000000101",
  27343=>"111000000",
  27344=>"000010111",
  27345=>"110110111",
  27346=>"000001011",
  27347=>"000000000",
  27348=>"111101000",
  27349=>"000100111",
  27350=>"110110111",
  27351=>"001101111",
  27352=>"000000111",
  27353=>"000111111",
  27354=>"011000000",
  27355=>"111101000",
  27356=>"111110000",
  27357=>"111001111",
  27358=>"101111001",
  27359=>"000100000",
  27360=>"111111000",
  27361=>"110000111",
  27362=>"001000100",
  27363=>"101111111",
  27364=>"000100111",
  27365=>"000110111",
  27366=>"010011100",
  27367=>"000000111",
  27368=>"001010110",
  27369=>"000010111",
  27370=>"001001111",
  27371=>"001101101",
  27372=>"000000000",
  27373=>"000010000",
  27374=>"111000000",
  27375=>"000101101",
  27376=>"011011110",
  27377=>"111011111",
  27378=>"100000000",
  27379=>"010011101",
  27380=>"000011001",
  27381=>"100000111",
  27382=>"001000000",
  27383=>"101010110",
  27384=>"100000000",
  27385=>"001000011",
  27386=>"010110111",
  27387=>"000010110",
  27388=>"110110100",
  27389=>"111111111",
  27390=>"100111001",
  27391=>"001100000",
  27392=>"011000101",
  27393=>"100000000",
  27394=>"111111111",
  27395=>"110010000",
  27396=>"010111111",
  27397=>"010100111",
  27398=>"101100100",
  27399=>"000000000",
  27400=>"110111100",
  27401=>"000100000",
  27402=>"000001000",
  27403=>"000000000",
  27404=>"111100000",
  27405=>"000000000",
  27406=>"100100100",
  27407=>"010111111",
  27408=>"111111000",
  27409=>"101111001",
  27410=>"111111110",
  27411=>"101011111",
  27412=>"000000100",
  27413=>"110110010",
  27414=>"000011111",
  27415=>"111000010",
  27416=>"100000000",
  27417=>"000000000",
  27418=>"100000000",
  27419=>"000011111",
  27420=>"001111111",
  27421=>"011101011",
  27422=>"000000100",
  27423=>"101101101",
  27424=>"010111111",
  27425=>"000000000",
  27426=>"111101000",
  27427=>"110101010",
  27428=>"010110000",
  27429=>"000011011",
  27430=>"111000000",
  27431=>"000111010",
  27432=>"000000000",
  27433=>"111111110",
  27434=>"111011111",
  27435=>"000111100",
  27436=>"000100100",
  27437=>"111001000",
  27438=>"000111111",
  27439=>"001011010",
  27440=>"111001000",
  27441=>"100100101",
  27442=>"000000000",
  27443=>"000000000",
  27444=>"000111110",
  27445=>"111011011",
  27446=>"100100001",
  27447=>"000011011",
  27448=>"000011000",
  27449=>"000000000",
  27450=>"000100000",
  27451=>"111111111",
  27452=>"110011011",
  27453=>"111111011",
  27454=>"000100111",
  27455=>"111010011",
  27456=>"111111000",
  27457=>"011000111",
  27458=>"000001000",
  27459=>"010011011",
  27460=>"010011010",
  27461=>"100111111",
  27462=>"000000110",
  27463=>"000000101",
  27464=>"000001000",
  27465=>"000000101",
  27466=>"110100001",
  27467=>"101000000",
  27468=>"111111111",
  27469=>"011011011",
  27470=>"011011101",
  27471=>"101001111",
  27472=>"101101111",
  27473=>"001111010",
  27474=>"000100101",
  27475=>"010110110",
  27476=>"100000001",
  27477=>"000110110",
  27478=>"001001001",
  27479=>"111000001",
  27480=>"110000000",
  27481=>"110111100",
  27482=>"001011011",
  27483=>"110111011",
  27484=>"000000100",
  27485=>"100110000",
  27486=>"000111110",
  27487=>"110110111",
  27488=>"000000000",
  27489=>"111101101",
  27490=>"101000000",
  27491=>"000110110",
  27492=>"011111111",
  27493=>"000111110",
  27494=>"000000000",
  27495=>"000010010",
  27496=>"101010100",
  27497=>"111010000",
  27498=>"000000010",
  27499=>"000001111",
  27500=>"111010010",
  27501=>"000000111",
  27502=>"000110111",
  27503=>"010000010",
  27504=>"000111100",
  27505=>"111001000",
  27506=>"001010110",
  27507=>"001000000",
  27508=>"101011000",
  27509=>"000000011",
  27510=>"101001000",
  27511=>"011011111",
  27512=>"000010100",
  27513=>"111011111",
  27514=>"111101001",
  27515=>"000001100",
  27516=>"011101111",
  27517=>"000000010",
  27518=>"111111111",
  27519=>"101000001",
  27520=>"111101111",
  27521=>"010100000",
  27522=>"111111010",
  27523=>"011111111",
  27524=>"000000000",
  27525=>"000111110",
  27526=>"000111111",
  27527=>"110100000",
  27528=>"000111010",
  27529=>"010111001",
  27530=>"001011010",
  27531=>"000101111",
  27532=>"000000000",
  27533=>"011111000",
  27534=>"000111110",
  27535=>"010001011",
  27536=>"011011111",
  27537=>"000000111",
  27538=>"000010101",
  27539=>"111101100",
  27540=>"111111111",
  27541=>"111111011",
  27542=>"000111100",
  27543=>"111100000",
  27544=>"011101001",
  27545=>"101000100",
  27546=>"000000011",
  27547=>"111111010",
  27548=>"000000000",
  27549=>"010011010",
  27550=>"100101111",
  27551=>"101000000",
  27552=>"100101001",
  27553=>"010110111",
  27554=>"000100101",
  27555=>"111101101",
  27556=>"111000001",
  27557=>"010111011",
  27558=>"010001011",
  27559=>"000000000",
  27560=>"000000011",
  27561=>"110101000",
  27562=>"111001001",
  27563=>"000000101",
  27564=>"111111000",
  27565=>"000011001",
  27566=>"110111111",
  27567=>"111111111",
  27568=>"100100000",
  27569=>"111001000",
  27570=>"011011001",
  27571=>"111000000",
  27572=>"110010011",
  27573=>"100101010",
  27574=>"011101110",
  27575=>"000000011",
  27576=>"110111100",
  27577=>"111111100",
  27578=>"000001110",
  27579=>"100010111",
  27580=>"000100000",
  27581=>"110111111",
  27582=>"111110100",
  27583=>"111100000",
  27584=>"111111111",
  27585=>"000011110",
  27586=>"011000000",
  27587=>"110000011",
  27588=>"000000001",
  27589=>"100011010",
  27590=>"010010001",
  27591=>"011111111",
  27592=>"000010100",
  27593=>"110000111",
  27594=>"111111111",
  27595=>"000101001",
  27596=>"000111111",
  27597=>"110111111",
  27598=>"100111111",
  27599=>"110011000",
  27600=>"111111111",
  27601=>"011110110",
  27602=>"111100101",
  27603=>"101110000",
  27604=>"001101101",
  27605=>"000000000",
  27606=>"000000000",
  27607=>"111100000",
  27608=>"000000000",
  27609=>"111000000",
  27610=>"010110100",
  27611=>"001000000",
  27612=>"111110111",
  27613=>"111101000",
  27614=>"111101011",
  27615=>"111111010",
  27616=>"101000001",
  27617=>"101101111",
  27618=>"000001101",
  27619=>"111111100",
  27620=>"000000100",
  27621=>"111001001",
  27622=>"110111011",
  27623=>"110110111",
  27624=>"100101001",
  27625=>"000000000",
  27626=>"000100011",
  27627=>"111101000",
  27628=>"111100100",
  27629=>"000011001",
  27630=>"111010000",
  27631=>"101000000",
  27632=>"111011000",
  27633=>"000101111",
  27634=>"000000100",
  27635=>"010111001",
  27636=>"010000011",
  27637=>"000000000",
  27638=>"000111110",
  27639=>"110100001",
  27640=>"111111111",
  27641=>"111011001",
  27642=>"000100111",
  27643=>"110110010",
  27644=>"001000011",
  27645=>"011000111",
  27646=>"000110111",
  27647=>"010111011",
  27648=>"111000001",
  27649=>"000010111",
  27650=>"100100110",
  27651=>"010000110",
  27652=>"100001001",
  27653=>"011110000",
  27654=>"111101000",
  27655=>"001000001",
  27656=>"000111111",
  27657=>"000101011",
  27658=>"001011001",
  27659=>"111111101",
  27660=>"101001001",
  27661=>"001111010",
  27662=>"000101001",
  27663=>"001011000",
  27664=>"111110111",
  27665=>"000111000",
  27666=>"010110011",
  27667=>"110101111",
  27668=>"111100011",
  27669=>"010100100",
  27670=>"100100100",
  27671=>"100011011",
  27672=>"111110011",
  27673=>"001011000",
  27674=>"001100010",
  27675=>"000101100",
  27676=>"111111100",
  27677=>"111111000",
  27678=>"111100100",
  27679=>"110001001",
  27680=>"011000001",
  27681=>"111111111",
  27682=>"111110011",
  27683=>"111101100",
  27684=>"011001010",
  27685=>"101011001",
  27686=>"111110111",
  27687=>"000011001",
  27688=>"000110011",
  27689=>"100110111",
  27690=>"111110000",
  27691=>"100010000",
  27692=>"100111100",
  27693=>"001010111",
  27694=>"000110000",
  27695=>"111100000",
  27696=>"011010001",
  27697=>"000100100",
  27698=>"001000110",
  27699=>"111100101",
  27700=>"111011011",
  27701=>"000000000",
  27702=>"000000001",
  27703=>"000001000",
  27704=>"110110111",
  27705=>"101000011",
  27706=>"000001000",
  27707=>"000001100",
  27708=>"100100100",
  27709=>"111111111",
  27710=>"000000100",
  27711=>"101111110",
  27712=>"000110100",
  27713=>"100001011",
  27714=>"010110001",
  27715=>"011001110",
  27716=>"001111100",
  27717=>"000000010",
  27718=>"000001001",
  27719=>"111110111",
  27720=>"111110011",
  27721=>"001001011",
  27722=>"011000011",
  27723=>"000011011",
  27724=>"000100010",
  27725=>"100100110",
  27726=>"110111111",
  27727=>"111111111",
  27728=>"100100100",
  27729=>"011111100",
  27730=>"001001001",
  27731=>"001001000",
  27732=>"010111110",
  27733=>"001010101",
  27734=>"001011100",
  27735=>"011100011",
  27736=>"111111111",
  27737=>"101000000",
  27738=>"011101001",
  27739=>"000001101",
  27740=>"000011011",
  27741=>"010000011",
  27742=>"110111100",
  27743=>"111010000",
  27744=>"000110111",
  27745=>"000100100",
  27746=>"110110010",
  27747=>"101011000",
  27748=>"000000011",
  27749=>"100001001",
  27750=>"000001000",
  27751=>"010100000",
  27752=>"011111111",
  27753=>"001000000",
  27754=>"000010110",
  27755=>"000011001",
  27756=>"010100100",
  27757=>"101100000",
  27758=>"110000100",
  27759=>"100101010",
  27760=>"000110100",
  27761=>"000000001",
  27762=>"110101111",
  27763=>"111101011",
  27764=>"001001000",
  27765=>"110000000",
  27766=>"100011101",
  27767=>"111100110",
  27768=>"110100010",
  27769=>"011111001",
  27770=>"100000101",
  27771=>"101101001",
  27772=>"110110110",
  27773=>"011011011",
  27774=>"001000001",
  27775=>"100010011",
  27776=>"010001000",
  27777=>"111110100",
  27778=>"011011011",
  27779=>"000101111",
  27780=>"001101111",
  27781=>"111011011",
  27782=>"110001001",
  27783=>"000000001",
  27784=>"101101111",
  27785=>"100100000",
  27786=>"000001011",
  27787=>"000001010",
  27788=>"100110110",
  27789=>"100000001",
  27790=>"111011011",
  27791=>"100000010",
  27792=>"101110101",
  27793=>"000001111",
  27794=>"000001011",
  27795=>"111101111",
  27796=>"001011010",
  27797=>"010100000",
  27798=>"000000000",
  27799=>"011010101",
  27800=>"001000001",
  27801=>"110100000",
  27802=>"111110111",
  27803=>"111110011",
  27804=>"000000110",
  27805=>"111110111",
  27806=>"000000000",
  27807=>"100101001",
  27808=>"010001101",
  27809=>"110000100",
  27810=>"011110011",
  27811=>"101110111",
  27812=>"111100001",
  27813=>"000011111",
  27814=>"011000000",
  27815=>"000001001",
  27816=>"000100011",
  27817=>"100111100",
  27818=>"001111100",
  27819=>"001110110",
  27820=>"110100111",
  27821=>"010010011",
  27822=>"001110000",
  27823=>"011000001",
  27824=>"001011000",
  27825=>"000000010",
  27826=>"011011000",
  27827=>"111100110",
  27828=>"000001001",
  27829=>"001010000",
  27830=>"000000001",
  27831=>"000000010",
  27832=>"100000001",
  27833=>"011101011",
  27834=>"001101000",
  27835=>"011000011",
  27836=>"000011000",
  27837=>"001111011",
  27838=>"000000001",
  27839=>"000001101",
  27840=>"111100001",
  27841=>"000100111",
  27842=>"111111111",
  27843=>"101101111",
  27844=>"000001001",
  27845=>"010010111",
  27846=>"000001001",
  27847=>"101110100",
  27848=>"001001000",
  27849=>"111000011",
  27850=>"101110111",
  27851=>"000011001",
  27852=>"111101000",
  27853=>"000110110",
  27854=>"000001001",
  27855=>"000000011",
  27856=>"111101100",
  27857=>"011000000",
  27858=>"100001111",
  27859=>"001001000",
  27860=>"111010000",
  27861=>"010111110",
  27862=>"101010110",
  27863=>"001001000",
  27864=>"001010011",
  27865=>"001001001",
  27866=>"100111110",
  27867=>"001000000",
  27868=>"011110100",
  27869=>"000111110",
  27870=>"100010000",
  27871=>"111101001",
  27872=>"110110100",
  27873=>"010100110",
  27874=>"011011000",
  27875=>"000110110",
  27876=>"110100101",
  27877=>"000111000",
  27878=>"101111111",
  27879=>"000101100",
  27880=>"001000000",
  27881=>"001011001",
  27882=>"110001011",
  27883=>"111110110",
  27884=>"001001011",
  27885=>"001011000",
  27886=>"001001001",
  27887=>"111010000",
  27888=>"101000011",
  27889=>"111100101",
  27890=>"011111000",
  27891=>"110111001",
  27892=>"001110110",
  27893=>"001101100",
  27894=>"011010011",
  27895=>"111000000",
  27896=>"110100111",
  27897=>"111011000",
  27898=>"111110000",
  27899=>"000011000",
  27900=>"010011000",
  27901=>"000001000",
  27902=>"001001011",
  27903=>"111110100",
  27904=>"000000000",
  27905=>"100100001",
  27906=>"101000000",
  27907=>"000000000",
  27908=>"010111101",
  27909=>"001011110",
  27910=>"111111000",
  27911=>"000000111",
  27912=>"010010100",
  27913=>"000000000",
  27914=>"110001000",
  27915=>"111101101",
  27916=>"110111101",
  27917=>"111111001",
  27918=>"000100111",
  27919=>"100001010",
  27920=>"111111111",
  27921=>"001111000",
  27922=>"000111000",
  27923=>"111111111",
  27924=>"010110111",
  27925=>"000001011",
  27926=>"111110100",
  27927=>"101110111",
  27928=>"000000000",
  27929=>"111111101",
  27930=>"000000000",
  27931=>"000000010",
  27932=>"111111101",
  27933=>"101101000",
  27934=>"111000000",
  27935=>"000101101",
  27936=>"111111111",
  27937=>"111111010",
  27938=>"000000000",
  27939=>"000000110",
  27940=>"111111011",
  27941=>"010100110",
  27942=>"111101000",
  27943=>"001000011",
  27944=>"010111111",
  27945=>"101110111",
  27946=>"000110110",
  27947=>"110111111",
  27948=>"111111111",
  27949=>"000110011",
  27950=>"111111111",
  27951=>"000000000",
  27952=>"111001000",
  27953=>"110110110",
  27954=>"001000000",
  27955=>"010010111",
  27956=>"100000000",
  27957=>"110101010",
  27958=>"110111011",
  27959=>"000000000",
  27960=>"011001100",
  27961=>"000000000",
  27962=>"000000000",
  27963=>"000000000",
  27964=>"110000110",
  27965=>"010111000",
  27966=>"110000000",
  27967=>"100100111",
  27968=>"100110101",
  27969=>"111101000",
  27970=>"111110100",
  27971=>"111100000",
  27972=>"010111000",
  27973=>"001101111",
  27974=>"111111011",
  27975=>"000111111",
  27976=>"000000011",
  27977=>"000010111",
  27978=>"111010000",
  27979=>"110110111",
  27980=>"101000000",
  27981=>"000110110",
  27982=>"010110111",
  27983=>"111110011",
  27984=>"111000001",
  27985=>"111110000",
  27986=>"000010011",
  27987=>"001000000",
  27988=>"111000000",
  27989=>"100100010",
  27990=>"100110000",
  27991=>"111101000",
  27992=>"000000001",
  27993=>"110110111",
  27994=>"000100000",
  27995=>"111111011",
  27996=>"111101101",
  27997=>"000000000",
  27998=>"000000000",
  27999=>"111111001",
  28000=>"111111111",
  28001=>"000111111",
  28002=>"110111111",
  28003=>"100000000",
  28004=>"000000000",
  28005=>"111010000",
  28006=>"110111000",
  28007=>"000000101",
  28008=>"111111111",
  28009=>"000000111",
  28010=>"010110110",
  28011=>"110010010",
  28012=>"110111011",
  28013=>"000000000",
  28014=>"111111000",
  28015=>"111010000",
  28016=>"010110110",
  28017=>"000000101",
  28018=>"111101110",
  28019=>"111111111",
  28020=>"011000000",
  28021=>"000000001",
  28022=>"000111111",
  28023=>"000101001",
  28024=>"100111111",
  28025=>"110110000",
  28026=>"000110111",
  28027=>"010010010",
  28028=>"011000100",
  28029=>"000000000",
  28030=>"000010110",
  28031=>"010000000",
  28032=>"110011000",
  28033=>"111100000",
  28034=>"000111101",
  28035=>"001010000",
  28036=>"010000000",
  28037=>"110111011",
  28038=>"111100001",
  28039=>"010011101",
  28040=>"001011111",
  28041=>"000001000",
  28042=>"000000010",
  28043=>"101111111",
  28044=>"000000000",
  28045=>"011001001",
  28046=>"000000000",
  28047=>"000000101",
  28048=>"000010000",
  28049=>"000000111",
  28050=>"100000010",
  28051=>"111110111",
  28052=>"000110111",
  28053=>"000000100",
  28054=>"010000000",
  28055=>"010110001",
  28056=>"000000100",
  28057=>"111111111",
  28058=>"111111110",
  28059=>"010110000",
  28060=>"000010000",
  28061=>"011111111",
  28062=>"000110110",
  28063=>"000000000",
  28064=>"001011100",
  28065=>"110110000",
  28066=>"111100110",
  28067=>"000000000",
  28068=>"010011010",
  28069=>"110110100",
  28070=>"001000000",
  28071=>"000111000",
  28072=>"000000110",
  28073=>"000001000",
  28074=>"000110100",
  28075=>"000110110",
  28076=>"010111001",
  28077=>"101000111",
  28078=>"110011011",
  28079=>"011111111",
  28080=>"000010000",
  28081=>"011100100",
  28082=>"000000011",
  28083=>"011111100",
  28084=>"100100001",
  28085=>"011111010",
  28086=>"110110000",
  28087=>"000101111",
  28088=>"001000011",
  28089=>"001110100",
  28090=>"000000000",
  28091=>"011111100",
  28092=>"010011111",
  28093=>"011111110",
  28094=>"001011011",
  28095=>"111000000",
  28096=>"101000000",
  28097=>"001000111",
  28098=>"111111101",
  28099=>"110001000",
  28100=>"101000000",
  28101=>"010100100",
  28102=>"000111111",
  28103=>"000001011",
  28104=>"111111101",
  28105=>"000111011",
  28106=>"101111111",
  28107=>"111111100",
  28108=>"100010110",
  28109=>"110001000",
  28110=>"110110111",
  28111=>"100111110",
  28112=>"101111111",
  28113=>"111110011",
  28114=>"011111101",
  28115=>"101000001",
  28116=>"001000111",
  28117=>"100001000",
  28118=>"000000000",
  28119=>"110000000",
  28120=>"111000111",
  28121=>"110000111",
  28122=>"110111001",
  28123=>"000010000",
  28124=>"110011001",
  28125=>"000111111",
  28126=>"110010000",
  28127=>"000010111",
  28128=>"000010010",
  28129=>"101000100",
  28130=>"001000000",
  28131=>"100110110",
  28132=>"100000000",
  28133=>"000001001",
  28134=>"000110111",
  28135=>"011001001",
  28136=>"111111111",
  28137=>"111101111",
  28138=>"010010000",
  28139=>"000010110",
  28140=>"101111111",
  28141=>"110100000",
  28142=>"000110000",
  28143=>"000011101",
  28144=>"000101000",
  28145=>"000011000",
  28146=>"101101000",
  28147=>"010011010",
  28148=>"000100010",
  28149=>"000010000",
  28150=>"000101011",
  28151=>"111000101",
  28152=>"010000000",
  28153=>"001111101",
  28154=>"010010101",
  28155=>"010000000",
  28156=>"010010100",
  28157=>"000000000",
  28158=>"000110100",
  28159=>"010010000",
  28160=>"011001101",
  28161=>"000000011",
  28162=>"101101001",
  28163=>"100000100",
  28164=>"000000101",
  28165=>"000000100",
  28166=>"111111111",
  28167=>"001010000",
  28168=>"111000000",
  28169=>"111000100",
  28170=>"000110110",
  28171=>"000000000",
  28172=>"001000101",
  28173=>"110000000",
  28174=>"011000000",
  28175=>"111111111",
  28176=>"000011111",
  28177=>"000000000",
  28178=>"111000000",
  28179=>"000100000",
  28180=>"000000110",
  28181=>"000000000",
  28182=>"000111011",
  28183=>"100000010",
  28184=>"100000100",
  28185=>"011111111",
  28186=>"001000110",
  28187=>"000011011",
  28188=>"111111010",
  28189=>"110010000",
  28190=>"001111100",
  28191=>"000000000",
  28192=>"011010000",
  28193=>"111101100",
  28194=>"101111111",
  28195=>"101000000",
  28196=>"110110000",
  28197=>"110101100",
  28198=>"000000000",
  28199=>"000000110",
  28200=>"000011000",
  28201=>"000000000",
  28202=>"110100010",
  28203=>"111111110",
  28204=>"011010000",
  28205=>"011001111",
  28206=>"010000111",
  28207=>"101100101",
  28208=>"001000110",
  28209=>"000111111",
  28210=>"101000111",
  28211=>"011111010",
  28212=>"010111111",
  28213=>"000000000",
  28214=>"001011110",
  28215=>"111111101",
  28216=>"011000111",
  28217=>"100000000",
  28218=>"111111010",
  28219=>"111111111",
  28220=>"000111000",
  28221=>"111111100",
  28222=>"000000000",
  28223=>"100011001",
  28224=>"111111111",
  28225=>"011010010",
  28226=>"111111101",
  28227=>"000000011",
  28228=>"000000000",
  28229=>"000000000",
  28230=>"000100010",
  28231=>"010000000",
  28232=>"001001100",
  28233=>"010111110",
  28234=>"101000111",
  28235=>"111111111",
  28236=>"111100000",
  28237=>"000000001",
  28238=>"000001111",
  28239=>"000000011",
  28240=>"111111010",
  28241=>"111111010",
  28242=>"100000111",
  28243=>"011001001",
  28244=>"000010110",
  28245=>"111111111",
  28246=>"011111010",
  28247=>"100101111",
  28248=>"000000010",
  28249=>"010100000",
  28250=>"001011111",
  28251=>"000100011",
  28252=>"111111000",
  28253=>"001011011",
  28254=>"111111111",
  28255=>"011011110",
  28256=>"010000000",
  28257=>"101011010",
  28258=>"101000101",
  28259=>"110111110",
  28260=>"000001011",
  28261=>"010111011",
  28262=>"010010010",
  28263=>"011000000",
  28264=>"001111111",
  28265=>"000001011",
  28266=>"111111010",
  28267=>"010000000",
  28268=>"000000000",
  28269=>"000100001",
  28270=>"000000101",
  28271=>"001001101",
  28272=>"000100100",
  28273=>"000000000",
  28274=>"010110010",
  28275=>"000101111",
  28276=>"110001000",
  28277=>"111000100",
  28278=>"100101000",
  28279=>"000001000",
  28280=>"000011000",
  28281=>"111111000",
  28282=>"100111111",
  28283=>"101000101",
  28284=>"111111111",
  28285=>"100100101",
  28286=>"110111111",
  28287=>"010000000",
  28288=>"111001100",
  28289=>"011111000",
  28290=>"000000010",
  28291=>"111111111",
  28292=>"000101000",
  28293=>"101001111",
  28294=>"000110001",
  28295=>"011011011",
  28296=>"101001010",
  28297=>"000000100",
  28298=>"001011111",
  28299=>"000000000",
  28300=>"000100100",
  28301=>"101000100",
  28302=>"100000000",
  28303=>"101001101",
  28304=>"001000011",
  28305=>"000010010",
  28306=>"000000111",
  28307=>"111010000",
  28308=>"001111011",
  28309=>"101100000",
  28310=>"111111100",
  28311=>"000000000",
  28312=>"001000000",
  28313=>"101100111",
  28314=>"101101000",
  28315=>"111011101",
  28316=>"101000000",
  28317=>"001101101",
  28318=>"000000111",
  28319=>"101000000",
  28320=>"101001011",
  28321=>"110111111",
  28322=>"100000100",
  28323=>"000000000",
  28324=>"000000011",
  28325=>"001001110",
  28326=>"110000001",
  28327=>"000000000",
  28328=>"010011111",
  28329=>"000000000",
  28330=>"101101101",
  28331=>"111001110",
  28332=>"111110100",
  28333=>"111000101",
  28334=>"111111110",
  28335=>"010001011",
  28336=>"000000100",
  28337=>"001101010",
  28338=>"110111111",
  28339=>"000100110",
  28340=>"011101111",
  28341=>"000000101",
  28342=>"000110000",
  28343=>"100000000",
  28344=>"001011000",
  28345=>"100110111",
  28346=>"111011101",
  28347=>"111110110",
  28348=>"000101001",
  28349=>"011111111",
  28350=>"001100000",
  28351=>"000000000",
  28352=>"000000000",
  28353=>"000000000",
  28354=>"010000111",
  28355=>"100000000",
  28356=>"000000011",
  28357=>"111110100",
  28358=>"010111111",
  28359=>"011111010",
  28360=>"111100001",
  28361=>"011011010",
  28362=>"111000001",
  28363=>"001000011",
  28364=>"110110010",
  28365=>"110111111",
  28366=>"111111010",
  28367=>"001010010",
  28368=>"000000100",
  28369=>"111111111",
  28370=>"101000100",
  28371=>"111111111",
  28372=>"000100101",
  28373=>"000010001",
  28374=>"101000000",
  28375=>"000010111",
  28376=>"000000000",
  28377=>"000000000",
  28378=>"101001010",
  28379=>"100100101",
  28380=>"111111110",
  28381=>"100000101",
  28382=>"111111111",
  28383=>"000000001",
  28384=>"010111010",
  28385=>"100111111",
  28386=>"101101111",
  28387=>"101101101",
  28388=>"000100000",
  28389=>"101000101",
  28390=>"000000000",
  28391=>"111111111",
  28392=>"100101001",
  28393=>"000100011",
  28394=>"010011011",
  28395=>"001000000",
  28396=>"000000000",
  28397=>"000000010",
  28398=>"110000000",
  28399=>"100000000",
  28400=>"001000000",
  28401=>"111011011",
  28402=>"010000011",
  28403=>"000011011",
  28404=>"000101111",
  28405=>"000111111",
  28406=>"000000000",
  28407=>"111101111",
  28408=>"000101111",
  28409=>"001111111",
  28410=>"000100100",
  28411=>"111100100",
  28412=>"011011001",
  28413=>"000111111",
  28414=>"011001001",
  28415=>"100000000",
  28416=>"111001100",
  28417=>"001000111",
  28418=>"000011011",
  28419=>"000001000",
  28420=>"111111111",
  28421=>"101001100",
  28422=>"010010000",
  28423=>"000011111",
  28424=>"111100000",
  28425=>"001000010",
  28426=>"001011110",
  28427=>"011111101",
  28428=>"000000000",
  28429=>"111100000",
  28430=>"110111111",
  28431=>"000010111",
  28432=>"000000000",
  28433=>"000111111",
  28434=>"111110010",
  28435=>"000100111",
  28436=>"010010000",
  28437=>"000010111",
  28438=>"111111111",
  28439=>"111010011",
  28440=>"000000000",
  28441=>"111000000",
  28442=>"001000000",
  28443=>"011011010",
  28444=>"001001000",
  28445=>"000101000",
  28446=>"000111100",
  28447=>"000000001",
  28448=>"111000010",
  28449=>"111000111",
  28450=>"010000000",
  28451=>"111111111",
  28452=>"011011011",
  28453=>"000001000",
  28454=>"110111000",
  28455=>"111000111",
  28456=>"100000101",
  28457=>"100100010",
  28458=>"111000000",
  28459=>"001101111",
  28460=>"010000110",
  28461=>"000000100",
  28462=>"011000100",
  28463=>"000010000",
  28464=>"000000010",
  28465=>"010111111",
  28466=>"111000010",
  28467=>"011111111",
  28468=>"101111001",
  28469=>"000010101",
  28470=>"111111011",
  28471=>"111111000",
  28472=>"001111101",
  28473=>"111111010",
  28474=>"000000001",
  28475=>"111111000",
  28476=>"000001001",
  28477=>"111111000",
  28478=>"001000000",
  28479=>"001111011",
  28480=>"110111000",
  28481=>"000000010",
  28482=>"111111111",
  28483=>"100100100",
  28484=>"101000001",
  28485=>"100101111",
  28486=>"010111000",
  28487=>"001000101",
  28488=>"000000110",
  28489=>"000001111",
  28490=>"110000000",
  28491=>"000010000",
  28492=>"000000000",
  28493=>"110011110",
  28494=>"110111010",
  28495=>"000010111",
  28496=>"110000000",
  28497=>"111111110",
  28498=>"000000000",
  28499=>"001100111",
  28500=>"000000000",
  28501=>"001011111",
  28502=>"111100100",
  28503=>"101000001",
  28504=>"000000001",
  28505=>"100101010",
  28506=>"001011011",
  28507=>"110110110",
  28508=>"011010000",
  28509=>"100000011",
  28510=>"001111000",
  28511=>"101001001",
  28512=>"100100000",
  28513=>"000101101",
  28514=>"000000101",
  28515=>"110110110",
  28516=>"000111010",
  28517=>"000000111",
  28518=>"010000000",
  28519=>"010010110",
  28520=>"101110000",
  28521=>"001001101",
  28522=>"111111111",
  28523=>"000000101",
  28524=>"000100110",
  28525=>"111011011",
  28526=>"000000000",
  28527=>"001001111",
  28528=>"010000001",
  28529=>"111111100",
  28530=>"111110110",
  28531=>"000000101",
  28532=>"111000000",
  28533=>"000100101",
  28534=>"000111111",
  28535=>"111111111",
  28536=>"111111011",
  28537=>"111000000",
  28538=>"111000000",
  28539=>"000101101",
  28540=>"101000010",
  28541=>"100001101",
  28542=>"011010011",
  28543=>"000000000",
  28544=>"011100110",
  28545=>"000000000",
  28546=>"011111110",
  28547=>"001110111",
  28548=>"000000110",
  28549=>"001101101",
  28550=>"000000000",
  28551=>"111000110",
  28552=>"000101000",
  28553=>"101101000",
  28554=>"000011011",
  28555=>"000101111",
  28556=>"000000000",
  28557=>"000000000",
  28558=>"000111001",
  28559=>"001000000",
  28560=>"001011111",
  28561=>"000011111",
  28562=>"111100111",
  28563=>"101101111",
  28564=>"100010000",
  28565=>"001111111",
  28566=>"001000000",
  28567=>"100010010",
  28568=>"000000111",
  28569=>"101100111",
  28570=>"101101110",
  28571=>"011111010",
  28572=>"100100111",
  28573=>"110000100",
  28574=>"111000000",
  28575=>"000000000",
  28576=>"100011101",
  28577=>"111111111",
  28578=>"000001111",
  28579=>"111111001",
  28580=>"011000111",
  28581=>"010011111",
  28582=>"001000101",
  28583=>"101110110",
  28584=>"000111111",
  28585=>"000000100",
  28586=>"111111101",
  28587=>"111111111",
  28588=>"001101101",
  28589=>"010101111",
  28590=>"111011010",
  28591=>"011111101",
  28592=>"000111000",
  28593=>"111000101",
  28594=>"001111001",
  28595=>"011100000",
  28596=>"001011111",
  28597=>"111111111",
  28598=>"100111111",
  28599=>"001000000",
  28600=>"000110100",
  28601=>"101011100",
  28602=>"101100000",
  28603=>"101000000",
  28604=>"001101001",
  28605=>"011100111",
  28606=>"111011001",
  28607=>"111000000",
  28608=>"111111000",
  28609=>"011111000",
  28610=>"010111111",
  28611=>"000110000",
  28612=>"000000100",
  28613=>"001001000",
  28614=>"000101111",
  28615=>"111000000",
  28616=>"111111001",
  28617=>"000001000",
  28618=>"111111011",
  28619=>"010111111",
  28620=>"010111011",
  28621=>"000001111",
  28622=>"111000000",
  28623=>"110100000",
  28624=>"101010010",
  28625=>"100110011",
  28626=>"101100100",
  28627=>"000000111",
  28628=>"000000000",
  28629=>"111000000",
  28630=>"110111011",
  28631=>"101100111",
  28632=>"000000000",
  28633=>"000000000",
  28634=>"011010100",
  28635=>"000000100",
  28636=>"111110111",
  28637=>"000000111",
  28638=>"000000000",
  28639=>"000000000",
  28640=>"000111011",
  28641=>"000000100",
  28642=>"000000111",
  28643=>"111110110",
  28644=>"101000000",
  28645=>"010110000",
  28646=>"101111111",
  28647=>"111110010",
  28648=>"000000000",
  28649=>"010000010",
  28650=>"111110011",
  28651=>"000000000",
  28652=>"000000000",
  28653=>"111001101",
  28654=>"010011010",
  28655=>"100000100",
  28656=>"000000100",
  28657=>"100100100",
  28658=>"001001100",
  28659=>"010111111",
  28660=>"110010001",
  28661=>"111111101",
  28662=>"000000101",
  28663=>"100000111",
  28664=>"111000000",
  28665=>"111011111",
  28666=>"101000000",
  28667=>"010010000",
  28668=>"111111011",
  28669=>"110000011",
  28670=>"101111001",
  28671=>"110111111",
  28672=>"100100111",
  28673=>"000000111",
  28674=>"101000000",
  28675=>"000010111",
  28676=>"000011011",
  28677=>"101000001",
  28678=>"100000110",
  28679=>"001000000",
  28680=>"000101000",
  28681=>"101101001",
  28682=>"110011011",
  28683=>"000000000",
  28684=>"010000101",
  28685=>"000100101",
  28686=>"010000010",
  28687=>"110001000",
  28688=>"010010000",
  28689=>"000000110",
  28690=>"101000111",
  28691=>"000000000",
  28692=>"000011111",
  28693=>"111000000",
  28694=>"000000011",
  28695=>"001111111",
  28696=>"000101110",
  28697=>"000000110",
  28698=>"001001001",
  28699=>"000111000",
  28700=>"110101111",
  28701=>"111111011",
  28702=>"011011011",
  28703=>"110000000",
  28704=>"100111111",
  28705=>"000010000",
  28706=>"110110000",
  28707=>"101101111",
  28708=>"111001001",
  28709=>"000001111",
  28710=>"000000111",
  28711=>"110111111",
  28712=>"011000000",
  28713=>"000000110",
  28714=>"101000001",
  28715=>"011001100",
  28716=>"000111111",
  28717=>"111101101",
  28718=>"111001111",
  28719=>"100010001",
  28720=>"111100000",
  28721=>"010011011",
  28722=>"111111001",
  28723=>"000010010",
  28724=>"000011111",
  28725=>"000110111",
  28726=>"100000011",
  28727=>"111101101",
  28728=>"000000100",
  28729=>"111111101",
  28730=>"001000000",
  28731=>"101111010",
  28732=>"111011111",
  28733=>"111111111",
  28734=>"001000111",
  28735=>"100111111",
  28736=>"011000100",
  28737=>"001000000",
  28738=>"000100101",
  28739=>"011001111",
  28740=>"000011010",
  28741=>"111100000",
  28742=>"000000000",
  28743=>"010000000",
  28744=>"111111001",
  28745=>"000111111",
  28746=>"111000000",
  28747=>"101101001",
  28748=>"101001111",
  28749=>"111101000",
  28750=>"001110110",
  28751=>"010010111",
  28752=>"000000001",
  28753=>"111001000",
  28754=>"110101111",
  28755=>"010011011",
  28756=>"100010000",
  28757=>"000111110",
  28758=>"010100100",
  28759=>"000110010",
  28760=>"110000000",
  28761=>"000010011",
  28762=>"110000011",
  28763=>"001000000",
  28764=>"111000001",
  28765=>"110000000",
  28766=>"111111111",
  28767=>"001001101",
  28768=>"010111111",
  28769=>"111000001",
  28770=>"100101111",
  28771=>"100000110",
  28772=>"001011001",
  28773=>"100100011",
  28774=>"010101111",
  28775=>"110111111",
  28776=>"111111000",
  28777=>"100011000",
  28778=>"010111111",
  28779=>"111000000",
  28780=>"111000110",
  28781=>"010111110",
  28782=>"111000000",
  28783=>"000100000",
  28784=>"000000011",
  28785=>"000000000",
  28786=>"001010110",
  28787=>"110110011",
  28788=>"111111111",
  28789=>"001000000",
  28790=>"111010000",
  28791=>"000111111",
  28792=>"000010111",
  28793=>"100111111",
  28794=>"000111111",
  28795=>"110111000",
  28796=>"110010110",
  28797=>"010101000",
  28798=>"000111000",
  28799=>"001001011",
  28800=>"000100000",
  28801=>"010101001",
  28802=>"000111111",
  28803=>"010110000",
  28804=>"001001010",
  28805=>"000000010",
  28806=>"100100110",
  28807=>"101001011",
  28808=>"100101000",
  28809=>"111011011",
  28810=>"000000000",
  28811=>"111000000",
  28812=>"111111000",
  28813=>"000000000",
  28814=>"000000000",
  28815=>"101000000",
  28816=>"111111011",
  28817=>"110000100",
  28818=>"001011000",
  28819=>"101011111",
  28820=>"101000100",
  28821=>"000000000",
  28822=>"110111101",
  28823=>"010110100",
  28824=>"111111111",
  28825=>"000000000",
  28826=>"111000000",
  28827=>"000100011",
  28828=>"111110100",
  28829=>"111101100",
  28830=>"001010100",
  28831=>"000111111",
  28832=>"011011101",
  28833=>"011010000",
  28834=>"011000000",
  28835=>"110010111",
  28836=>"101111111",
  28837=>"000000100",
  28838=>"000001001",
  28839=>"111000001",
  28840=>"000101111",
  28841=>"000111111",
  28842=>"111100000",
  28843=>"011000110",
  28844=>"101000001",
  28845=>"001001001",
  28846=>"110011011",
  28847=>"110111111",
  28848=>"111110000",
  28849=>"111111101",
  28850=>"000101101",
  28851=>"110000100",
  28852=>"011000001",
  28853=>"000011011",
  28854=>"010101011",
  28855=>"000010000",
  28856=>"111110111",
  28857=>"000000110",
  28858=>"010000111",
  28859=>"001000011",
  28860=>"111100111",
  28861=>"111101101",
  28862=>"001111111",
  28863=>"000110111",
  28864=>"000010111",
  28865=>"111000000",
  28866=>"111000101",
  28867=>"110110110",
  28868=>"000111011",
  28869=>"100110110",
  28870=>"000000001",
  28871=>"000000000",
  28872=>"111111110",
  28873=>"010110000",
  28874=>"000110010",
  28875=>"111001000",
  28876=>"000111011",
  28877=>"001000101",
  28878=>"001000110",
  28879=>"100110111",
  28880=>"000111111",
  28881=>"010011001",
  28882=>"001010110",
  28883=>"110000000",
  28884=>"111111011",
  28885=>"011001010",
  28886=>"100000001",
  28887=>"000000000",
  28888=>"100111000",
  28889=>"010111001",
  28890=>"010101100",
  28891=>"000000001",
  28892=>"000000110",
  28893=>"110000000",
  28894=>"011000000",
  28895=>"000000001",
  28896=>"000010010",
  28897=>"011000000",
  28898=>"111111111",
  28899=>"000110110",
  28900=>"100111110",
  28901=>"000010111",
  28902=>"001000101",
  28903=>"110100100",
  28904=>"111001001",
  28905=>"111111111",
  28906=>"000110110",
  28907=>"000110111",
  28908=>"000000000",
  28909=>"101000110",
  28910=>"111101101",
  28911=>"100111101",
  28912=>"100111000",
  28913=>"101001001",
  28914=>"000000111",
  28915=>"000110111",
  28916=>"101011111",
  28917=>"111001001",
  28918=>"111000000",
  28919=>"000010000",
  28920=>"000010000",
  28921=>"111111001",
  28922=>"111111100",
  28923=>"000000111",
  28924=>"100000000",
  28925=>"000010000",
  28926=>"011111110",
  28927=>"111000000",
  28928=>"000000000",
  28929=>"000000010",
  28930=>"111101101",
  28931=>"110000000",
  28932=>"001100100",
  28933=>"011101101",
  28934=>"000111000",
  28935=>"111010010",
  28936=>"011101100",
  28937=>"000100101",
  28938=>"110101111",
  28939=>"000011111",
  28940=>"000000000",
  28941=>"111101111",
  28942=>"011000010",
  28943=>"010011000",
  28944=>"000110110",
  28945=>"011000100",
  28946=>"100100110",
  28947=>"000101101",
  28948=>"100101001",
  28949=>"101111100",
  28950=>"001001010",
  28951=>"001000001",
  28952=>"101001000",
  28953=>"101110111",
  28954=>"010101010",
  28955=>"000000111",
  28956=>"100000000",
  28957=>"000011010",
  28958=>"010000100",
  28959=>"000010010",
  28960=>"111001101",
  28961=>"111101111",
  28962=>"101110101",
  28963=>"001010000",
  28964=>"101000001",
  28965=>"001001100",
  28966=>"010000101",
  28967=>"000000111",
  28968=>"111101111",
  28969=>"011100111",
  28970=>"000000000",
  28971=>"100001000",
  28972=>"100111111",
  28973=>"111111111",
  28974=>"010111101",
  28975=>"111111000",
  28976=>"111111101",
  28977=>"101100001",
  28978=>"111111111",
  28979=>"111001101",
  28980=>"010000011",
  28981=>"000111001",
  28982=>"011110100",
  28983=>"101100101",
  28984=>"001111101",
  28985=>"111101101",
  28986=>"000101000",
  28987=>"000111111",
  28988=>"110110011",
  28989=>"110111111",
  28990=>"101101101",
  28991=>"011000101",
  28992=>"101101101",
  28993=>"000111101",
  28994=>"110011001",
  28995=>"010000000",
  28996=>"010101001",
  28997=>"000100101",
  28998=>"000100101",
  28999=>"100111111",
  29000=>"111111111",
  29001=>"010000010",
  29002=>"111101101",
  29003=>"011101111",
  29004=>"010000000",
  29005=>"111000000",
  29006=>"111100000",
  29007=>"101111111",
  29008=>"000000000",
  29009=>"110111111",
  29010=>"100000101",
  29011=>"010011001",
  29012=>"000000000",
  29013=>"100010110",
  29014=>"000001110",
  29015=>"101100101",
  29016=>"011100110",
  29017=>"100010110",
  29018=>"010000011",
  29019=>"000000100",
  29020=>"111101101",
  29021=>"010000010",
  29022=>"111111011",
  29023=>"100000000",
  29024=>"011111000",
  29025=>"100101010",
  29026=>"110101101",
  29027=>"001001111",
  29028=>"110100000",
  29029=>"000010111",
  29030=>"111110111",
  29031=>"101100000",
  29032=>"100101000",
  29033=>"111110100",
  29034=>"111000101",
  29035=>"111111001",
  29036=>"000011001",
  29037=>"111101111",
  29038=>"001000100",
  29039=>"000111110",
  29040=>"101001001",
  29041=>"000001000",
  29042=>"000001001",
  29043=>"000000111",
  29044=>"111111101",
  29045=>"000000001",
  29046=>"110000001",
  29047=>"010111111",
  29048=>"110111110",
  29049=>"001111110",
  29050=>"111000000",
  29051=>"111010100",
  29052=>"011100000",
  29053=>"010110110",
  29054=>"000000010",
  29055=>"111101000",
  29056=>"010011101",
  29057=>"111111001",
  29058=>"111000101",
  29059=>"011110101",
  29060=>"000000000",
  29061=>"111111111",
  29062=>"100101011",
  29063=>"111001110",
  29064=>"101111110",
  29065=>"111001110",
  29066=>"000000111",
  29067=>"111111101",
  29068=>"000101101",
  29069=>"111100010",
  29070=>"000010000",
  29071=>"000000001",
  29072=>"011001010",
  29073=>"000110111",
  29074=>"000010111",
  29075=>"011111111",
  29076=>"000101000",
  29077=>"111100101",
  29078=>"000010111",
  29079=>"100100000",
  29080=>"101111111",
  29081=>"111010001",
  29082=>"100100100",
  29083=>"111100000",
  29084=>"010000100",
  29085=>"111000000",
  29086=>"011000100",
  29087=>"010000011",
  29088=>"100111011",
  29089=>"111100011",
  29090=>"000011011",
  29091=>"000000101",
  29092=>"111000111",
  29093=>"111110001",
  29094=>"101000101",
  29095=>"110101111",
  29096=>"000011001",
  29097=>"110000000",
  29098=>"111101101",
  29099=>"111000000",
  29100=>"001110101",
  29101=>"010101010",
  29102=>"001001010",
  29103=>"100101110",
  29104=>"000101111",
  29105=>"100111011",
  29106=>"111111100",
  29107=>"001001001",
  29108=>"000011111",
  29109=>"110011000",
  29110=>"000011011",
  29111=>"011000010",
  29112=>"000011010",
  29113=>"001101001",
  29114=>"010010011",
  29115=>"000111111",
  29116=>"101011000",
  29117=>"111111001",
  29118=>"010000000",
  29119=>"100101000",
  29120=>"010111111",
  29121=>"111101100",
  29122=>"111100100",
  29123=>"110000100",
  29124=>"100010110",
  29125=>"010011010",
  29126=>"000000100",
  29127=>"111100110",
  29128=>"000000111",
  29129=>"111101100",
  29130=>"110010100",
  29131=>"001001001",
  29132=>"111111110",
  29133=>"100100011",
  29134=>"000100011",
  29135=>"111101101",
  29136=>"111010001",
  29137=>"000111010",
  29138=>"100110100",
  29139=>"000010000",
  29140=>"111000111",
  29141=>"001110110",
  29142=>"001000010",
  29143=>"000110111",
  29144=>"000011111",
  29145=>"011100100",
  29146=>"111111110",
  29147=>"101100000",
  29148=>"100000000",
  29149=>"111101000",
  29150=>"000010010",
  29151=>"110101101",
  29152=>"111101001",
  29153=>"011101010",
  29154=>"101000000",
  29155=>"000001011",
  29156=>"010000000",
  29157=>"101111011",
  29158=>"111000000",
  29159=>"000100000",
  29160=>"011101001",
  29161=>"101000000",
  29162=>"111000011",
  29163=>"010010111",
  29164=>"111100101",
  29165=>"111000101",
  29166=>"000000111",
  29167=>"000110010",
  29168=>"000010111",
  29169=>"110111110",
  29170=>"000000000",
  29171=>"000110111",
  29172=>"010000000",
  29173=>"011000000",
  29174=>"010000100",
  29175=>"000010010",
  29176=>"111100100",
  29177=>"000000001",
  29178=>"111111000",
  29179=>"011110000",
  29180=>"110000000",
  29181=>"000111001",
  29182=>"110111111",
  29183=>"111101111",
  29184=>"101001000",
  29185=>"000011011",
  29186=>"000000000",
  29187=>"000011111",
  29188=>"101101100",
  29189=>"011011001",
  29190=>"010001000",
  29191=>"010011110",
  29192=>"001001011",
  29193=>"011001001",
  29194=>"010011001",
  29195=>"010111000",
  29196=>"001001001",
  29197=>"111110100",
  29198=>"101001101",
  29199=>"010100110",
  29200=>"111011001",
  29201=>"000001001",
  29202=>"101100101",
  29203=>"101011011",
  29204=>"010001000",
  29205=>"111111111",
  29206=>"100101110",
  29207=>"100111111",
  29208=>"001001000",
  29209=>"011011111",
  29210=>"011011101",
  29211=>"010011011",
  29212=>"000100100",
  29213=>"111010110",
  29214=>"011001001",
  29215=>"000010110",
  29216=>"000000000",
  29217=>"001000011",
  29218=>"000100110",
  29219=>"000001011",
  29220=>"011111110",
  29221=>"000000010",
  29222=>"001001111",
  29223=>"000001000",
  29224=>"111110110",
  29225=>"000001011",
  29226=>"000000101",
  29227=>"110110010",
  29228=>"111100100",
  29229=>"001001001",
  29230=>"011010001",
  29231=>"100110000",
  29232=>"001011111",
  29233=>"000000011",
  29234=>"000000011",
  29235=>"011001001",
  29236=>"000001001",
  29237=>"000000000",
  29238=>"000000000",
  29239=>"101001001",
  29240=>"011111000",
  29241=>"011011011",
  29242=>"100100100",
  29243=>"011011000",
  29244=>"011001111",
  29245=>"110110110",
  29246=>"000000001",
  29247=>"011011000",
  29248=>"111011001",
  29249=>"011001011",
  29250=>"000111010",
  29251=>"101000011",
  29252=>"011010000",
  29253=>"001101000",
  29254=>"100011000",
  29255=>"000100111",
  29256=>"100000110",
  29257=>"110111111",
  29258=>"111101111",
  29259=>"001101001",
  29260=>"001000100",
  29261=>"001001001",
  29262=>"000001001",
  29263=>"000000000",
  29264=>"000000000",
  29265=>"110000110",
  29266=>"111111011",
  29267=>"010000010",
  29268=>"000011110",
  29269=>"010000000",
  29270=>"100110111",
  29271=>"011011000",
  29272=>"000000111",
  29273=>"010000011",
  29274=>"010110110",
  29275=>"101101111",
  29276=>"011011001",
  29277=>"000010111",
  29278=>"001011001",
  29279=>"010010000",
  29280=>"000010010",
  29281=>"110110000",
  29282=>"011010000",
  29283=>"100101100",
  29284=>"000010110",
  29285=>"000111100",
  29286=>"111000111",
  29287=>"001000110",
  29288=>"011011111",
  29289=>"010001001",
  29290=>"110110011",
  29291=>"010011111",
  29292=>"110101111",
  29293=>"110110100",
  29294=>"001000000",
  29295=>"000000100",
  29296=>"101000001",
  29297=>"011111111",
  29298=>"001010001",
  29299=>"000000000",
  29300=>"011000010",
  29301=>"001001001",
  29302=>"000011011",
  29303=>"111100001",
  29304=>"000000000",
  29305=>"010100110",
  29306=>"000100110",
  29307=>"111011111",
  29308=>"111011000",
  29309=>"111001000",
  29310=>"100110111",
  29311=>"000110110",
  29312=>"001001001",
  29313=>"110110011",
  29314=>"001001011",
  29315=>"001000000",
  29316=>"111111110",
  29317=>"100110000",
  29318=>"011110100",
  29319=>"100100100",
  29320=>"011011010",
  29321=>"100110111",
  29322=>"011111001",
  29323=>"000001000",
  29324=>"001111011",
  29325=>"111111000",
  29326=>"011000011",
  29327=>"000001011",
  29328=>"101100101",
  29329=>"111101110",
  29330=>"000000001",
  29331=>"000111011",
  29332=>"000101111",
  29333=>"001001001",
  29334=>"001000010",
  29335=>"101100100",
  29336=>"000010101",
  29337=>"000000111",
  29338=>"001000010",
  29339=>"001000010",
  29340=>"001101111",
  29341=>"000000000",
  29342=>"000111001",
  29343=>"100100001",
  29344=>"100000001",
  29345=>"011111011",
  29346=>"000010110",
  29347=>"000000001",
  29348=>"110011011",
  29349=>"101001111",
  29350=>"011111010",
  29351=>"100000110",
  29352=>"001011001",
  29353=>"001101101",
  29354=>"101001001",
  29355=>"000001000",
  29356=>"001111100",
  29357=>"101000000",
  29358=>"010010000",
  29359=>"011010001",
  29360=>"011001001",
  29361=>"110011001",
  29362=>"000000000",
  29363=>"000001011",
  29364=>"010011011",
  29365=>"010100010",
  29366=>"101000101",
  29367=>"010011000",
  29368=>"100100100",
  29369=>"010010010",
  29370=>"001000110",
  29371=>"011110111",
  29372=>"110110100",
  29373=>"100110110",
  29374=>"100010000",
  29375=>"000001010",
  29376=>"001001001",
  29377=>"011000001",
  29378=>"011111111",
  29379=>"000011010",
  29380=>"000001111",
  29381=>"000110010",
  29382=>"110100111",
  29383=>"011000111",
  29384=>"100000110",
  29385=>"111010010",
  29386=>"110000011",
  29387=>"000100101",
  29388=>"100101101",
  29389=>"000000000",
  29390=>"001001001",
  29391=>"111101100",
  29392=>"101000000",
  29393=>"100100110",
  29394=>"111001001",
  29395=>"110110110",
  29396=>"001001111",
  29397=>"100110110",
  29398=>"000011000",
  29399=>"011111001",
  29400=>"000010010",
  29401=>"110010110",
  29402=>"011000000",
  29403=>"001001001",
  29404=>"011111111",
  29405=>"100100111",
  29406=>"111111111",
  29407=>"000111011",
  29408=>"000000001",
  29409=>"001001001",
  29410=>"100110111",
  29411=>"110110011",
  29412=>"001001001",
  29413=>"110110110",
  29414=>"111111010",
  29415=>"101111010",
  29416=>"000100111",
  29417=>"100010000",
  29418=>"001111101",
  29419=>"011011000",
  29420=>"001000011",
  29421=>"001111110",
  29422=>"100000100",
  29423=>"000100111",
  29424=>"000000000",
  29425=>"101100101",
  29426=>"001001001",
  29427=>"101101100",
  29428=>"011000001",
  29429=>"100110110",
  29430=>"000001110",
  29431=>"110110100",
  29432=>"001001001",
  29433=>"001111010",
  29434=>"101100001",
  29435=>"111110110",
  29436=>"111111111",
  29437=>"110110111",
  29438=>"001110110",
  29439=>"001111000",
  29440=>"110110011",
  29441=>"001001001",
  29442=>"111000000",
  29443=>"111010000",
  29444=>"001000001",
  29445=>"000000000",
  29446=>"110010010",
  29447=>"010000010",
  29448=>"000000000",
  29449=>"000110010",
  29450=>"001011000",
  29451=>"000110100",
  29452=>"001000111",
  29453=>"000000000",
  29454=>"100111011",
  29455=>"111111101",
  29456=>"001000000",
  29457=>"110110011",
  29458=>"111000000",
  29459=>"000000011",
  29460=>"111111010",
  29461=>"000100111",
  29462=>"100100100",
  29463=>"010000000",
  29464=>"000000000",
  29465=>"000000110",
  29466=>"100101011",
  29467=>"011000111",
  29468=>"100101000",
  29469=>"001100000",
  29470=>"111110000",
  29471=>"101101000",
  29472=>"000111100",
  29473=>"011011000",
  29474=>"110111111",
  29475=>"101101000",
  29476=>"001001000",
  29477=>"000100110",
  29478=>"100101111",
  29479=>"101111101",
  29480=>"101010111",
  29481=>"111101101",
  29482=>"110111101",
  29483=>"111111001",
  29484=>"011111111",
  29485=>"011100111",
  29486=>"111111111",
  29487=>"110100000",
  29488=>"000011011",
  29489=>"010101001",
  29490=>"000011010",
  29491=>"000111111",
  29492=>"001101111",
  29493=>"000111000",
  29494=>"001001001",
  29495=>"000111110",
  29496=>"001010111",
  29497=>"010000011",
  29498=>"011001000",
  29499=>"000000101",
  29500=>"001001001",
  29501=>"111101000",
  29502=>"000010001",
  29503=>"010110001",
  29504=>"101111000",
  29505=>"100111011",
  29506=>"111000111",
  29507=>"001001001",
  29508=>"101001011",
  29509=>"000000000",
  29510=>"000000000",
  29511=>"010011010",
  29512=>"001001100",
  29513=>"000110110",
  29514=>"000010110",
  29515=>"000110001",
  29516=>"001101011",
  29517=>"000001001",
  29518=>"000000001",
  29519=>"011111101",
  29520=>"111000000",
  29521=>"000000000",
  29522=>"000001111",
  29523=>"011011101",
  29524=>"101000000",
  29525=>"101101000",
  29526=>"010000001",
  29527=>"111111010",
  29528=>"111111101",
  29529=>"010100101",
  29530=>"011001000",
  29531=>"000011011",
  29532=>"001000000",
  29533=>"010011001",
  29534=>"000011111",
  29535=>"001110100",
  29536=>"101111111",
  29537=>"111010111",
  29538=>"101001000",
  29539=>"110010000",
  29540=>"010010100",
  29541=>"111101111",
  29542=>"011011000",
  29543=>"011110000",
  29544=>"000011111",
  29545=>"110110110",
  29546=>"010001000",
  29547=>"001110010",
  29548=>"111101010",
  29549=>"110010011",
  29550=>"111111010",
  29551=>"000000010",
  29552=>"000001000",
  29553=>"000000111",
  29554=>"100100100",
  29555=>"000001000",
  29556=>"100111000",
  29557=>"111010111",
  29558=>"111111110",
  29559=>"000000000",
  29560=>"111011010",
  29561=>"011101101",
  29562=>"000001101",
  29563=>"000111111",
  29564=>"000110100",
  29565=>"110110001",
  29566=>"101111010",
  29567=>"000000110",
  29568=>"000000101",
  29569=>"000000000",
  29570=>"111100000",
  29571=>"111111001",
  29572=>"101001000",
  29573=>"000110010",
  29574=>"001001011",
  29575=>"110000000",
  29576=>"001001001",
  29577=>"110000110",
  29578=>"010010111",
  29579=>"000000000",
  29580=>"000101111",
  29581=>"011111011",
  29582=>"010001001",
  29583=>"000000000",
  29584=>"000100101",
  29585=>"101111111",
  29586=>"000110111",
  29587=>"111111101",
  29588=>"000000011",
  29589=>"001000000",
  29590=>"111111001",
  29591=>"000000001",
  29592=>"011010011",
  29593=>"001001111",
  29594=>"101001111",
  29595=>"000110000",
  29596=>"010110000",
  29597=>"001001101",
  29598=>"001110000",
  29599=>"111100001",
  29600=>"101100100",
  29601=>"000101111",
  29602=>"101111111",
  29603=>"000000000",
  29604=>"100110011",
  29605=>"100100100",
  29606=>"000000100",
  29607=>"100111100",
  29608=>"111000100",
  29609=>"000101101",
  29610=>"111101110",
  29611=>"111101000",
  29612=>"001000000",
  29613=>"000000001",
  29614=>"011011001",
  29615=>"010011110",
  29616=>"000100000",
  29617=>"011010000",
  29618=>"000011111",
  29619=>"011001000",
  29620=>"000001001",
  29621=>"001101000",
  29622=>"000010011",
  29623=>"000110111",
  29624=>"100100100",
  29625=>"000100110",
  29626=>"000100101",
  29627=>"010110010",
  29628=>"111111111",
  29629=>"110010010",
  29630=>"000100010",
  29631=>"101011111",
  29632=>"001101011",
  29633=>"111011000",
  29634=>"010000010",
  29635=>"001011001",
  29636=>"000000011",
  29637=>"110110101",
  29638=>"001000000",
  29639=>"110111110",
  29640=>"111000000",
  29641=>"100000111",
  29642=>"000110010",
  29643=>"101000111",
  29644=>"100111010",
  29645=>"001011000",
  29646=>"111101001",
  29647=>"011111001",
  29648=>"011101111",
  29649=>"000000011",
  29650=>"000000110",
  29651=>"101101110",
  29652=>"111000110",
  29653=>"111010000",
  29654=>"111111001",
  29655=>"110111100",
  29656=>"000000111",
  29657=>"000000000",
  29658=>"111011011",
  29659=>"000000110",
  29660=>"001001001",
  29661=>"001000000",
  29662=>"001111111",
  29663=>"011111110",
  29664=>"000000000",
  29665=>"101001111",
  29666=>"101101111",
  29667=>"011111101",
  29668=>"000000000",
  29669=>"101010000",
  29670=>"000000010",
  29671=>"100100100",
  29672=>"010110010",
  29673=>"110111101",
  29674=>"100110000",
  29675=>"111111011",
  29676=>"000000110",
  29677=>"000000111",
  29678=>"100000010",
  29679=>"001000111",
  29680=>"001101001",
  29681=>"101111101",
  29682=>"101101111",
  29683=>"111111001",
  29684=>"011001110",
  29685=>"010110101",
  29686=>"010000000",
  29687=>"011111111",
  29688=>"101001000",
  29689=>"101101111",
  29690=>"011111000",
  29691=>"010000101",
  29692=>"010111101",
  29693=>"001000000",
  29694=>"010000100",
  29695=>"111111000",
  29696=>"000000011",
  29697=>"100000000",
  29698=>"010010000",
  29699=>"010000011",
  29700=>"100101111",
  29701=>"110110000",
  29702=>"111011111",
  29703=>"000010110",
  29704=>"000001101",
  29705=>"000111111",
  29706=>"100100101",
  29707=>"101110110",
  29708=>"111001000",
  29709=>"110111000",
  29710=>"000011010",
  29711=>"000010000",
  29712=>"000001000",
  29713=>"000010000",
  29714=>"000000000",
  29715=>"101111111",
  29716=>"001100010",
  29717=>"000110010",
  29718=>"010000000",
  29719=>"001011110",
  29720=>"000000000",
  29721=>"101001111",
  29722=>"001001111",
  29723=>"000000000",
  29724=>"000000111",
  29725=>"101001111",
  29726=>"000000000",
  29727=>"000001111",
  29728=>"111000000",
  29729=>"000101000",
  29730=>"000000000",
  29731=>"000000000",
  29732=>"101111111",
  29733=>"001000110",
  29734=>"111010000",
  29735=>"111000011",
  29736=>"010111111",
  29737=>"000100110",
  29738=>"110111101",
  29739=>"111111111",
  29740=>"001001111",
  29741=>"000000011",
  29742=>"101001000",
  29743=>"010001001",
  29744=>"010000101",
  29745=>"111111111",
  29746=>"000101000",
  29747=>"000000000",
  29748=>"111110011",
  29749=>"111010110",
  29750=>"110001001",
  29751=>"000111111",
  29752=>"111000000",
  29753=>"000000000",
  29754=>"001000000",
  29755=>"111000000",
  29756=>"101111111",
  29757=>"111111000",
  29758=>"000000010",
  29759=>"110110110",
  29760=>"001000000",
  29761=>"100101101",
  29762=>"111000010",
  29763=>"110111111",
  29764=>"010000111",
  29765=>"000001000",
  29766=>"001101100",
  29767=>"111111001",
  29768=>"101111111",
  29769=>"000001000",
  29770=>"000000001",
  29771=>"000000001",
  29772=>"001011111",
  29773=>"111011111",
  29774=>"011111111",
  29775=>"110000000",
  29776=>"001100000",
  29777=>"111000000",
  29778=>"111000111",
  29779=>"011001101",
  29780=>"101000010",
  29781=>"101100111",
  29782=>"011011001",
  29783=>"110111100",
  29784=>"001011001",
  29785=>"111101111",
  29786=>"100100000",
  29787=>"101101101",
  29788=>"000000100",
  29789=>"000000001",
  29790=>"111111111",
  29791=>"110111011",
  29792=>"010110010",
  29793=>"000000000",
  29794=>"000000000",
  29795=>"010111000",
  29796=>"000000000",
  29797=>"111101000",
  29798=>"111001111",
  29799=>"101111111",
  29800=>"010000000",
  29801=>"000101111",
  29802=>"000000011",
  29803=>"111111110",
  29804=>"110000110",
  29805=>"110010000",
  29806=>"001001111",
  29807=>"000100000",
  29808=>"101011011",
  29809=>"001101101",
  29810=>"011100101",
  29811=>"010000000",
  29812=>"111111111",
  29813=>"000000101",
  29814=>"111111101",
  29815=>"111111000",
  29816=>"110111100",
  29817=>"001000000",
  29818=>"100000110",
  29819=>"111001001",
  29820=>"100000110",
  29821=>"100000000",
  29822=>"111000010",
  29823=>"001001001",
  29824=>"001000100",
  29825=>"111101000",
  29826=>"000100110",
  29827=>"111101110",
  29828=>"001000010",
  29829=>"111001010",
  29830=>"101101111",
  29831=>"010001101",
  29832=>"001001001",
  29833=>"111100000",
  29834=>"101000001",
  29835=>"001000100",
  29836=>"010111111",
  29837=>"000000110",
  29838=>"110111011",
  29839=>"001000000",
  29840=>"001001011",
  29841=>"110010110",
  29842=>"110000001",
  29843=>"010100110",
  29844=>"000010010",
  29845=>"111111110",
  29846=>"110011110",
  29847=>"000001001",
  29848=>"111111111",
  29849=>"111101111",
  29850=>"111111111",
  29851=>"010000100",
  29852=>"100111010",
  29853=>"111111011",
  29854=>"000010111",
  29855=>"101000101",
  29856=>"111100100",
  29857=>"000000000",
  29858=>"110111010",
  29859=>"111101111",
  29860=>"101000101",
  29861=>"001001100",
  29862=>"000000000",
  29863=>"111101001",
  29864=>"101010011",
  29865=>"000000000",
  29866=>"111001000",
  29867=>"000000000",
  29868=>"000001000",
  29869=>"000110000",
  29870=>"000000100",
  29871=>"010001011",
  29872=>"111110110",
  29873=>"110100001",
  29874=>"111111101",
  29875=>"000000100",
  29876=>"100100100",
  29877=>"000000000",
  29878=>"111111111",
  29879=>"000101101",
  29880=>"001011111",
  29881=>"100100100",
  29882=>"110110011",
  29883=>"000000110",
  29884=>"100111111",
  29885=>"111111111",
  29886=>"011011011",
  29887=>"011000000",
  29888=>"000010010",
  29889=>"000000000",
  29890=>"101110100",
  29891=>"011101101",
  29892=>"001111000",
  29893=>"101000001",
  29894=>"000000111",
  29895=>"001000000",
  29896=>"101111110",
  29897=>"110010101",
  29898=>"011111011",
  29899=>"111011111",
  29900=>"011111000",
  29901=>"010011011",
  29902=>"000000000",
  29903=>"111111111",
  29904=>"000000000",
  29905=>"110000010",
  29906=>"001001110",
  29907=>"001011110",
  29908=>"101010000",
  29909=>"001000000",
  29910=>"000000000",
  29911=>"101111111",
  29912=>"111111111",
  29913=>"000100111",
  29914=>"111001001",
  29915=>"001000000",
  29916=>"000000000",
  29917=>"101001001",
  29918=>"101111111",
  29919=>"110000111",
  29920=>"000000001",
  29921=>"000000000",
  29922=>"111111111",
  29923=>"100000000",
  29924=>"001000000",
  29925=>"001000000",
  29926=>"101111111",
  29927=>"100010000",
  29928=>"111111111",
  29929=>"101000001",
  29930=>"000000001",
  29931=>"110010010",
  29932=>"000000000",
  29933=>"101111111",
  29934=>"000000000",
  29935=>"000000111",
  29936=>"101111111",
  29937=>"111011000",
  29938=>"000000100",
  29939=>"001001001",
  29940=>"000000100",
  29941=>"000000000",
  29942=>"001000111",
  29943=>"111111101",
  29944=>"101100111",
  29945=>"001010010",
  29946=>"101111011",
  29947=>"100010001",
  29948=>"000000000",
  29949=>"111111111",
  29950=>"000000101",
  29951=>"111110000",
  29952=>"000001001",
  29953=>"100111111",
  29954=>"000000100",
  29955=>"101101101",
  29956=>"110011101",
  29957=>"100010110",
  29958=>"111011011",
  29959=>"100111111",
  29960=>"000000000",
  29961=>"000000110",
  29962=>"000000100",
  29963=>"110100010",
  29964=>"011000000",
  29965=>"110010011",
  29966=>"001001110",
  29967=>"001101001",
  29968=>"100000000",
  29969=>"111000110",
  29970=>"000000000",
  29971=>"011000111",
  29972=>"100100111",
  29973=>"000011000",
  29974=>"010110011",
  29975=>"001001011",
  29976=>"001101000",
  29977=>"010100100",
  29978=>"100000111",
  29979=>"000000100",
  29980=>"110000011",
  29981=>"100111110",
  29982=>"000010000",
  29983=>"101101100",
  29984=>"111100011",
  29985=>"100110010",
  29986=>"000010001",
  29987=>"111111011",
  29988=>"001001110",
  29989=>"011100111",
  29990=>"011000100",
  29991=>"001100111",
  29992=>"000000101",
  29993=>"110010011",
  29994=>"001100001",
  29995=>"101100010",
  29996=>"001111011",
  29997=>"110111111",
  29998=>"100101111",
  29999=>"000100011",
  30000=>"000111111",
  30001=>"110010001",
  30002=>"110110100",
  30003=>"000011111",
  30004=>"000000000",
  30005=>"000111011",
  30006=>"000001111",
  30007=>"000011111",
  30008=>"011111010",
  30009=>"101000011",
  30010=>"000100001",
  30011=>"111011111",
  30012=>"010001100",
  30013=>"111111000",
  30014=>"000000101",
  30015=>"001100001",
  30016=>"111111001",
  30017=>"001000010",
  30018=>"011011001",
  30019=>"110000100",
  30020=>"011011000",
  30021=>"000010101",
  30022=>"000100111",
  30023=>"011111110",
  30024=>"001111111",
  30025=>"000000011",
  30026=>"101100101",
  30027=>"111100111",
  30028=>"000000100",
  30029=>"110110011",
  30030=>"011001010",
  30031=>"011111111",
  30032=>"000010111",
  30033=>"000100100",
  30034=>"001000000",
  30035=>"000110110",
  30036=>"110100000",
  30037=>"111101100",
  30038=>"010001011",
  30039=>"111000110",
  30040=>"000100100",
  30041=>"110010000",
  30042=>"110111110",
  30043=>"001100000",
  30044=>"011010000",
  30045=>"000000101",
  30046=>"011011000",
  30047=>"001100100",
  30048=>"011000000",
  30049=>"000000110",
  30050=>"111000000",
  30051=>"100101001",
  30052=>"100110011",
  30053=>"100100011",
  30054=>"000101111",
  30055=>"000100111",
  30056=>"000011000",
  30057=>"100000000",
  30058=>"110111000",
  30059=>"000011110",
  30060=>"111110100",
  30061=>"101000111",
  30062=>"000000001",
  30063=>"011001111",
  30064=>"110100111",
  30065=>"100100110",
  30066=>"100110110",
  30067=>"011011000",
  30068=>"111110001",
  30069=>"000000011",
  30070=>"100111000",
  30071=>"011000000",
  30072=>"000000000",
  30073=>"011000101",
  30074=>"100110000",
  30075=>"111101011",
  30076=>"100111111",
  30077=>"100100111",
  30078=>"111001000",
  30079=>"000000100",
  30080=>"001011011",
  30081=>"000011111",
  30082=>"011000011",
  30083=>"001000010",
  30084=>"000010111",
  30085=>"001101011",
  30086=>"010000001",
  30087=>"010001000",
  30088=>"101111000",
  30089=>"100011011",
  30090=>"100100011",
  30091=>"100011000",
  30092=>"001000111",
  30093=>"000111111",
  30094=>"001000000",
  30095=>"000000000",
  30096=>"110111111",
  30097=>"000011001",
  30098=>"000000010",
  30099=>"010000000",
  30100=>"001101010",
  30101=>"001000100",
  30102=>"011111000",
  30103=>"001001011",
  30104=>"100001111",
  30105=>"001100000",
  30106=>"000100111",
  30107=>"000000110",
  30108=>"011000011",
  30109=>"000000011",
  30110=>"000111011",
  30111=>"101000100",
  30112=>"000111111",
  30113=>"100100111",
  30114=>"000000111",
  30115=>"100100000",
  30116=>"100000000",
  30117=>"000011110",
  30118=>"100010000",
  30119=>"011110110",
  30120=>"111001111",
  30121=>"111111111",
  30122=>"111100111",
  30123=>"011000000",
  30124=>"101000011",
  30125=>"000100100",
  30126=>"001101100",
  30127=>"111011011",
  30128=>"000000011",
  30129=>"000101110",
  30130=>"000100110",
  30131=>"100000000",
  30132=>"110101100",
  30133=>"111011111",
  30134=>"011000001",
  30135=>"011011000",
  30136=>"101000000",
  30137=>"110101101",
  30138=>"000010000",
  30139=>"011100000",
  30140=>"111010001",
  30141=>"111111101",
  30142=>"110100100",
  30143=>"000000111",
  30144=>"000100101",
  30145=>"100000000",
  30146=>"001111011",
  30147=>"110110001",
  30148=>"000110110",
  30149=>"010111111",
  30150=>"110010110",
  30151=>"001001111",
  30152=>"111111011",
  30153=>"011011000",
  30154=>"000101010",
  30155=>"111001100",
  30156=>"000000100",
  30157=>"011001010",
  30158=>"000001000",
  30159=>"111011000",
  30160=>"111100100",
  30161=>"111110100",
  30162=>"010000001",
  30163=>"000000000",
  30164=>"000100111",
  30165=>"100110111",
  30166=>"101011001",
  30167=>"100111111",
  30168=>"111101011",
  30169=>"011000100",
  30170=>"111101111",
  30171=>"001000111",
  30172=>"111000110",
  30173=>"111000100",
  30174=>"011000000",
  30175=>"000111110",
  30176=>"011011000",
  30177=>"000100000",
  30178=>"100000000",
  30179=>"010100111",
  30180=>"111000000",
  30181=>"001010000",
  30182=>"111101011",
  30183=>"100100111",
  30184=>"011000010",
  30185=>"101001000",
  30186=>"010000001",
  30187=>"111011000",
  30188=>"011011000",
  30189=>"011011011",
  30190=>"000010000",
  30191=>"111100100",
  30192=>"100111011",
  30193=>"000101001",
  30194=>"011010000",
  30195=>"001101101",
  30196=>"100110110",
  30197=>"000001011",
  30198=>"000000000",
  30199=>"100100111",
  30200=>"000111010",
  30201=>"000101011",
  30202=>"100000111",
  30203=>"100100010",
  30204=>"111100001",
  30205=>"101000000",
  30206=>"000000001",
  30207=>"100100011",
  30208=>"000100000",
  30209=>"001001010",
  30210=>"100000000",
  30211=>"000101101",
  30212=>"110111011",
  30213=>"001001101",
  30214=>"101111111",
  30215=>"111000000",
  30216=>"000001001",
  30217=>"100000000",
  30218=>"100100111",
  30219=>"000111111",
  30220=>"101111111",
  30221=>"000011111",
  30222=>"100010101",
  30223=>"111110111",
  30224=>"100010111",
  30225=>"111000111",
  30226=>"010000110",
  30227=>"111000000",
  30228=>"101111001",
  30229=>"000000110",
  30230=>"110110101",
  30231=>"110111011",
  30232=>"000000000",
  30233=>"100000000",
  30234=>"001100100",
  30235=>"000010111",
  30236=>"000000011",
  30237=>"010101000",
  30238=>"101010000",
  30239=>"001000101",
  30240=>"111101111",
  30241=>"110111111",
  30242=>"001000000",
  30243=>"000000000",
  30244=>"110011100",
  30245=>"100000000",
  30246=>"111000111",
  30247=>"111000101",
  30248=>"111111000",
  30249=>"101111011",
  30250=>"100000101",
  30251=>"111000000",
  30252=>"101100010",
  30253=>"111000110",
  30254=>"101000000",
  30255=>"111111111",
  30256=>"000111111",
  30257=>"011111001",
  30258=>"111101111",
  30259=>"100000000",
  30260=>"111001000",
  30261=>"000111111",
  30262=>"110100011",
  30263=>"000111111",
  30264=>"110000000",
  30265=>"000000001",
  30266=>"001000000",
  30267=>"111111111",
  30268=>"001011101",
  30269=>"000010001",
  30270=>"000000101",
  30271=>"000001101",
  30272=>"101011111",
  30273=>"111010010",
  30274=>"000011110",
  30275=>"000000000",
  30276=>"111101000",
  30277=>"000101011",
  30278=>"000110011",
  30279=>"111000111",
  30280=>"000001101",
  30281=>"000000100",
  30282=>"101000000",
  30283=>"000001011",
  30284=>"111000001",
  30285=>"111000000",
  30286=>"111111110",
  30287=>"000000001",
  30288=>"100000000",
  30289=>"000111001",
  30290=>"100100000",
  30291=>"100000000",
  30292=>"000000000",
  30293=>"011110111",
  30294=>"111000000",
  30295=>"110000010",
  30296=>"101000001",
  30297=>"111000001",
  30298=>"101111111",
  30299=>"010100100",
  30300=>"000000000",
  30301=>"100100000",
  30302=>"111111111",
  30303=>"100000000",
  30304=>"111101101",
  30305=>"000000000",
  30306=>"000000000",
  30307=>"110110111",
  30308=>"000001101",
  30309=>"011001011",
  30310=>"000000000",
  30311=>"000000000",
  30312=>"001001000",
  30313=>"111111011",
  30314=>"111000000",
  30315=>"000100011",
  30316=>"011000110",
  30317=>"111111100",
  30318=>"000100111",
  30319=>"010101111",
  30320=>"100110000",
  30321=>"000000111",
  30322=>"011000110",
  30323=>"111000000",
  30324=>"011011111",
  30325=>"100000000",
  30326=>"110111111",
  30327=>"000111101",
  30328=>"101010101",
  30329=>"111001001",
  30330=>"110111110",
  30331=>"111101000",
  30332=>"001001001",
  30333=>"001000000",
  30334=>"111111111",
  30335=>"000100000",
  30336=>"001000100",
  30337=>"000011011",
  30338=>"000001111",
  30339=>"001001100",
  30340=>"000000010",
  30341=>"010000000",
  30342=>"010011000",
  30343=>"000000100",
  30344=>"001111110",
  30345=>"011000100",
  30346=>"111111000",
  30347=>"100111111",
  30348=>"011111000",
  30349=>"000000000",
  30350=>"111111111",
  30351=>"101000101",
  30352=>"001101001",
  30353=>"111011111",
  30354=>"010111111",
  30355=>"000011101",
  30356=>"000000100",
  30357=>"000000000",
  30358=>"111111100",
  30359=>"110111111",
  30360=>"111001000",
  30361=>"001000000",
  30362=>"010000001",
  30363=>"110000111",
  30364=>"000000000",
  30365=>"010111000",
  30366=>"001100101",
  30367=>"111000111",
  30368=>"110100011",
  30369=>"111000101",
  30370=>"001000011",
  30371=>"000000000",
  30372=>"101001101",
  30373=>"011000001",
  30374=>"101100111",
  30375=>"111111101",
  30376=>"000000000",
  30377=>"111011101",
  30378=>"000000000",
  30379=>"111000000",
  30380=>"000101110",
  30381=>"000000000",
  30382=>"101010110",
  30383=>"001000010",
  30384=>"000110111",
  30385=>"100000110",
  30386=>"100000011",
  30387=>"000000100",
  30388=>"100110001",
  30389=>"010100111",
  30390=>"111100100",
  30391=>"011111101",
  30392=>"000000000",
  30393=>"010110001",
  30394=>"101000000",
  30395=>"000001111",
  30396=>"000101010",
  30397=>"011111010",
  30398=>"111110101",
  30399=>"111000000",
  30400=>"000000001",
  30401=>"000000111",
  30402=>"110010110",
  30403=>"011111111",
  30404=>"111111111",
  30405=>"001011111",
  30406=>"110110011",
  30407=>"111000001",
  30408=>"111100110",
  30409=>"000010110",
  30410=>"101111111",
  30411=>"100000000",
  30412=>"100000000",
  30413=>"000000000",
  30414=>"111111111",
  30415=>"010111101",
  30416=>"001000001",
  30417=>"111111001",
  30418=>"000100111",
  30419=>"111111100",
  30420=>"000000000",
  30421=>"001011011",
  30422=>"000000000",
  30423=>"000000111",
  30424=>"111111111",
  30425=>"011000000",
  30426=>"011000000",
  30427=>"111111000",
  30428=>"000001111",
  30429=>"111000001",
  30430=>"111000100",
  30431=>"000000111",
  30432=>"000000100",
  30433=>"000010010",
  30434=>"000111111",
  30435=>"111100000",
  30436=>"000000101",
  30437=>"101111011",
  30438=>"000000111",
  30439=>"011101001",
  30440=>"111001000",
  30441=>"111111011",
  30442=>"111100111",
  30443=>"000000001",
  30444=>"011111111",
  30445=>"111001110",
  30446=>"000000000",
  30447=>"100001111",
  30448=>"011000010",
  30449=>"000010110",
  30450=>"000001011",
  30451=>"001000001",
  30452=>"101001000",
  30453=>"010110111",
  30454=>"100000000",
  30455=>"000010111",
  30456=>"110111000",
  30457=>"111011011",
  30458=>"000000000",
  30459=>"111111111",
  30460=>"111000101",
  30461=>"001110111",
  30462=>"000000000",
  30463=>"110000000",
  30464=>"011111100",
  30465=>"010111111",
  30466=>"000000101",
  30467=>"101111000",
  30468=>"000000010",
  30469=>"000000000",
  30470=>"000000010",
  30471=>"111111111",
  30472=>"111111111",
  30473=>"111100000",
  30474=>"111010100",
  30475=>"101011001",
  30476=>"001011000",
  30477=>"000000000",
  30478=>"000000100",
  30479=>"111111110",
  30480=>"111110101",
  30481=>"101101000",
  30482=>"111111111",
  30483=>"111101000",
  30484=>"110110010",
  30485=>"111000001",
  30486=>"000010110",
  30487=>"110100001",
  30488=>"100100111",
  30489=>"100111001",
  30490=>"000001011",
  30491=>"111111111",
  30492=>"110101010",
  30493=>"000010000",
  30494=>"111001011",
  30495=>"110000000",
  30496=>"000010110",
  30497=>"111111000",
  30498=>"111010001",
  30499=>"000000000",
  30500=>"100100101",
  30501=>"111111011",
  30502=>"000101011",
  30503=>"001110010",
  30504=>"111111111",
  30505=>"111010111",
  30506=>"000000000",
  30507=>"001110000",
  30508=>"000110000",
  30509=>"111111000",
  30510=>"010010000",
  30511=>"001000010",
  30512=>"000000110",
  30513=>"101011011",
  30514=>"101000011",
  30515=>"111111000",
  30516=>"000000010",
  30517=>"110110010",
  30518=>"001011011",
  30519=>"111101100",
  30520=>"110011011",
  30521=>"000000001",
  30522=>"011001001",
  30523=>"100111111",
  30524=>"111111011",
  30525=>"111111111",
  30526=>"000000000",
  30527=>"000000110",
  30528=>"010000101",
  30529=>"101100101",
  30530=>"001101111",
  30531=>"010000001",
  30532=>"111111111",
  30533=>"010000000",
  30534=>"010111110",
  30535=>"010000000",
  30536=>"111110001",
  30537=>"011010011",
  30538=>"000111111",
  30539=>"011111011",
  30540=>"000000101",
  30541=>"000000110",
  30542=>"000110111",
  30543=>"111110111",
  30544=>"110101111",
  30545=>"111111110",
  30546=>"111111111",
  30547=>"111001001",
  30548=>"110111011",
  30549=>"111110100",
  30550=>"111110101",
  30551=>"110100111",
  30552=>"100001000",
  30553=>"011011000",
  30554=>"000101011",
  30555=>"000011011",
  30556=>"000000111",
  30557=>"001001011",
  30558=>"111000111",
  30559=>"111000100",
  30560=>"110100000",
  30561=>"111011110",
  30562=>"000000000",
  30563=>"000001101",
  30564=>"000101111",
  30565=>"100011010",
  30566=>"010111011",
  30567=>"111000110",
  30568=>"010111111",
  30569=>"010000000",
  30570=>"000001110",
  30571=>"010000100",
  30572=>"110110111",
  30573=>"001000000",
  30574=>"010010000",
  30575=>"000101111",
  30576=>"000100110",
  30577=>"000011101",
  30578=>"110110110",
  30579=>"110000111",
  30580=>"111111000",
  30581=>"100000011",
  30582=>"000000000",
  30583=>"110000000",
  30584=>"111111000",
  30585=>"000110010",
  30586=>"111111111",
  30587=>"101111111",
  30588=>"110110101",
  30589=>"100000000",
  30590=>"101000100",
  30591=>"100000110",
  30592=>"000101000",
  30593=>"111000000",
  30594=>"100000000",
  30595=>"001001111",
  30596=>"111111111",
  30597=>"101111111",
  30598=>"100010000",
  30599=>"001000000",
  30600=>"000010110",
  30601=>"000010101",
  30602=>"111101110",
  30603=>"010000000",
  30604=>"111000111",
  30605=>"000000000",
  30606=>"111010111",
  30607=>"001000100",
  30608=>"000111111",
  30609=>"111000010",
  30610=>"000100111",
  30611=>"001010000",
  30612=>"000110000",
  30613=>"011111000",
  30614=>"000000101",
  30615=>"111111111",
  30616=>"010110011",
  30617=>"111000000",
  30618=>"101000001",
  30619=>"011111110",
  30620=>"111111100",
  30621=>"111011110",
  30622=>"111010000",
  30623=>"000001000",
  30624=>"100010000",
  30625=>"001000111",
  30626=>"000000000",
  30627=>"001010011",
  30628=>"000000000",
  30629=>"100101100",
  30630=>"110101011",
  30631=>"000100010",
  30632=>"011111110",
  30633=>"011111101",
  30634=>"101111110",
  30635=>"111111101",
  30636=>"000000010",
  30637=>"010000111",
  30638=>"101111101",
  30639=>"000111010",
  30640=>"000101111",
  30641=>"011101101",
  30642=>"001000000",
  30643=>"101101111",
  30644=>"000011011",
  30645=>"000000010",
  30646=>"010000011",
  30647=>"010000000",
  30648=>"111100110",
  30649=>"111010011",
  30650=>"110110111",
  30651=>"000000000",
  30652=>"000111010",
  30653=>"111010000",
  30654=>"111100110",
  30655=>"000000010",
  30656=>"010001111",
  30657=>"000000000",
  30658=>"110111100",
  30659=>"000001011",
  30660=>"011010000",
  30661=>"101111100",
  30662=>"011111010",
  30663=>"100000111",
  30664=>"111100000",
  30665=>"110000100",
  30666=>"000010000",
  30667=>"111000001",
  30668=>"010000000",
  30669=>"011111110",
  30670=>"000000101",
  30671=>"000000010",
  30672=>"111111000",
  30673=>"100111111",
  30674=>"111011011",
  30675=>"111111111",
  30676=>"111111111",
  30677=>"000011111",
  30678=>"000100101",
  30679=>"110010100",
  30680=>"010000000",
  30681=>"001110001",
  30682=>"101110000",
  30683=>"101100101",
  30684=>"110110010",
  30685=>"000111000",
  30686=>"010010110",
  30687=>"100000101",
  30688=>"111101111",
  30689=>"000001100",
  30690=>"101010010",
  30691=>"000101111",
  30692=>"111111011",
  30693=>"010000000",
  30694=>"000000000",
  30695=>"100000000",
  30696=>"010110000",
  30697=>"000000100",
  30698=>"101011001",
  30699=>"111111111",
  30700=>"110000000",
  30701=>"011110100",
  30702=>"111001000",
  30703=>"111001001",
  30704=>"111111000",
  30705=>"111111001",
  30706=>"110111011",
  30707=>"111111110",
  30708=>"110001011",
  30709=>"000100101",
  30710=>"001001001",
  30711=>"101111111",
  30712=>"111110001",
  30713=>"111111100",
  30714=>"111111110",
  30715=>"000111010",
  30716=>"001001101",
  30717=>"000101010",
  30718=>"001011011",
  30719=>"000101001",
  30720=>"010111101",
  30721=>"101111111",
  30722=>"000101010",
  30723=>"000000010",
  30724=>"100111000",
  30725=>"000111101",
  30726=>"111011011",
  30727=>"011011000",
  30728=>"001000100",
  30729=>"010010111",
  30730=>"011110100",
  30731=>"101011101",
  30732=>"101101101",
  30733=>"101101101",
  30734=>"011011010",
  30735=>"111111111",
  30736=>"000000000",
  30737=>"000000011",
  30738=>"101101111",
  30739=>"000011000",
  30740=>"111111111",
  30741=>"110100001",
  30742=>"000001001",
  30743=>"000000000",
  30744=>"010000000",
  30745=>"100101111",
  30746=>"101101010",
  30747=>"010010000",
  30748=>"100000101",
  30749=>"011110010",
  30750=>"100111011",
  30751=>"000000101",
  30752=>"101100100",
  30753=>"101100111",
  30754=>"101010001",
  30755=>"000000000",
  30756=>"110100100",
  30757=>"100111111",
  30758=>"100101100",
  30759=>"101010101",
  30760=>"101101100",
  30761=>"011011000",
  30762=>"000000000",
  30763=>"010000001",
  30764=>"011011011",
  30765=>"110010010",
  30766=>"000101111",
  30767=>"111111101",
  30768=>"010101000",
  30769=>"100011011",
  30770=>"000000000",
  30771=>"010111010",
  30772=>"011111101",
  30773=>"010111101",
  30774=>"001001100",
  30775=>"011111101",
  30776=>"001101100",
  30777=>"001000000",
  30778=>"100100110",
  30779=>"010010010",
  30780=>"000001001",
  30781=>"111111101",
  30782=>"010000001",
  30783=>"000100000",
  30784=>"001001000",
  30785=>"110110100",
  30786=>"000110110",
  30787=>"000010110",
  30788=>"111001010",
  30789=>"011101001",
  30790=>"111010100",
  30791=>"000000000",
  30792=>"101100010",
  30793=>"010101010",
  30794=>"011101111",
  30795=>"010011011",
  30796=>"000100101",
  30797=>"101001000",
  30798=>"000100100",
  30799=>"010010010",
  30800=>"001000111",
  30801=>"000000111",
  30802=>"111010101",
  30803=>"001001000",
  30804=>"001001000",
  30805=>"001011100",
  30806=>"011000100",
  30807=>"101100000",
  30808=>"000111100",
  30809=>"110011000",
  30810=>"000000001",
  30811=>"001111111",
  30812=>"000000000",
  30813=>"001001001",
  30814=>"000100111",
  30815=>"001110101",
  30816=>"111111111",
  30817=>"111000000",
  30818=>"000100001",
  30819=>"110000000",
  30820=>"110111100",
  30821=>"001110100",
  30822=>"111010101",
  30823=>"110110010",
  30824=>"000010110",
  30825=>"010110111",
  30826=>"001010111",
  30827=>"110110010",
  30828=>"010010011",
  30829=>"010110000",
  30830=>"010010000",
  30831=>"110101101",
  30832=>"001001111",
  30833=>"111111110",
  30834=>"000000101",
  30835=>"111100000",
  30836=>"111111111",
  30837=>"100101101",
  30838=>"101000100",
  30839=>"111101111",
  30840=>"000100100",
  30841=>"010000000",
  30842=>"111110111",
  30843=>"000000000",
  30844=>"110111011",
  30845=>"100100001",
  30846=>"000000000",
  30847=>"001000111",
  30848=>"000000110",
  30849=>"000101000",
  30850=>"010011100",
  30851=>"111111111",
  30852=>"111111001",
  30853=>"110010101",
  30854=>"001110111",
  30855=>"100001011",
  30856=>"101101111",
  30857=>"110111111",
  30858=>"010010000",
  30859=>"100000000",
  30860=>"000001001",
  30861=>"010110010",
  30862=>"111001000",
  30863=>"101101101",
  30864=>"111101111",
  30865=>"101111101",
  30866=>"000001101",
  30867=>"101100000",
  30868=>"011011011",
  30869=>"000010111",
  30870=>"111100101",
  30871=>"100100110",
  30872=>"010010111",
  30873=>"000111000",
  30874=>"010010000",
  30875=>"000000000",
  30876=>"111111000",
  30877=>"000001001",
  30878=>"010000100",
  30879=>"011101001",
  30880=>"111011001",
  30881=>"100000000",
  30882=>"001000010",
  30883=>"000000000",
  30884=>"000010000",
  30885=>"101101111",
  30886=>"000001011",
  30887=>"010010011",
  30888=>"011000111",
  30889=>"001001000",
  30890=>"000101111",
  30891=>"011001001",
  30892=>"110011101",
  30893=>"010000000",
  30894=>"111111111",
  30895=>"010011010",
  30896=>"000000111",
  30897=>"011111001",
  30898=>"101101100",
  30899=>"100110010",
  30900=>"100101000",
  30901=>"010011110",
  30902=>"111100100",
  30903=>"100101101",
  30904=>"000100100",
  30905=>"111110110",
  30906=>"000000011",
  30907=>"111111000",
  30908=>"111111010",
  30909=>"000000000",
  30910=>"101001110",
  30911=>"010101110",
  30912=>"101001101",
  30913=>"011010000",
  30914=>"000110101",
  30915=>"111011011",
  30916=>"011001000",
  30917=>"110100100",
  30918=>"000001000",
  30919=>"000000000",
  30920=>"001101111",
  30921=>"101101001",
  30922=>"100111100",
  30923=>"111110100",
  30924=>"101000111",
  30925=>"001011110",
  30926=>"010001101",
  30927=>"100111111",
  30928=>"000000101",
  30929=>"111011000",
  30930=>"111110110",
  30931=>"111110101",
  30932=>"101111111",
  30933=>"100000100",
  30934=>"101100000",
  30935=>"010110111",
  30936=>"101011010",
  30937=>"001011001",
  30938=>"110000000",
  30939=>"010000000",
  30940=>"000001000",
  30941=>"000100000",
  30942=>"111111011",
  30943=>"000000100",
  30944=>"000100011",
  30945=>"000001110",
  30946=>"100000001",
  30947=>"111111111",
  30948=>"000100010",
  30949=>"101011111",
  30950=>"111110101",
  30951=>"011111111",
  30952=>"000010001",
  30953=>"111000101",
  30954=>"110111001",
  30955=>"100000000",
  30956=>"111101101",
  30957=>"101000000",
  30958=>"000000000",
  30959=>"000011111",
  30960=>"111111111",
  30961=>"101001101",
  30962=>"000010010",
  30963=>"000000000",
  30964=>"010001001",
  30965=>"110011101",
  30966=>"100000110",
  30967=>"000000011",
  30968=>"000000000",
  30969=>"111010110",
  30970=>"111111111",
  30971=>"000000100",
  30972=>"111111000",
  30973=>"101011101",
  30974=>"011011000",
  30975=>"011110111",
  30976=>"011001001",
  30977=>"000000111",
  30978=>"000000111",
  30979=>"111100010",
  30980=>"000000100",
  30981=>"010000000",
  30982=>"111011110",
  30983=>"111111110",
  30984=>"011100100",
  30985=>"100001101",
  30986=>"110111000",
  30987=>"000000011",
  30988=>"101001110",
  30989=>"001110000",
  30990=>"111001001",
  30991=>"100000000",
  30992=>"110110010",
  30993=>"000101000",
  30994=>"000000000",
  30995=>"000000011",
  30996=>"111111000",
  30997=>"001001000",
  30998=>"000001000",
  30999=>"000000010",
  31000=>"110010000",
  31001=>"010111000",
  31002=>"011000000",
  31003=>"000111110",
  31004=>"111110110",
  31005=>"000000000",
  31006=>"111001000",
  31007=>"000101111",
  31008=>"010110010",
  31009=>"001001111",
  31010=>"111001101",
  31011=>"100000100",
  31012=>"000101100",
  31013=>"100011110",
  31014=>"111111000",
  31015=>"101110100",
  31016=>"110110111",
  31017=>"111111111",
  31018=>"000010011",
  31019=>"110001000",
  31020=>"000000100",
  31021=>"111111110",
  31022=>"110000111",
  31023=>"000001001",
  31024=>"000000000",
  31025=>"000011001",
  31026=>"111100000",
  31027=>"000001010",
  31028=>"111111000",
  31029=>"111111010",
  31030=>"000000100",
  31031=>"011000000",
  31032=>"110001111",
  31033=>"111001101",
  31034=>"000000100",
  31035=>"111111100",
  31036=>"100111111",
  31037=>"100111111",
  31038=>"001000101",
  31039=>"110110000",
  31040=>"010011101",
  31041=>"000001111",
  31042=>"111111000",
  31043=>"110110000",
  31044=>"000000101",
  31045=>"011001000",
  31046=>"010000111",
  31047=>"101101101",
  31048=>"101111111",
  31049=>"110110000",
  31050=>"101100000",
  31051=>"111110111",
  31052=>"001000111",
  31053=>"001111011",
  31054=>"100101101",
  31055=>"101101111",
  31056=>"001000001",
  31057=>"010000000",
  31058=>"111110100",
  31059=>"100001000",
  31060=>"000000101",
  31061=>"110000011",
  31062=>"100101110",
  31063=>"111111000",
  31064=>"110100111",
  31065=>"110100110",
  31066=>"001000001",
  31067=>"000001001",
  31068=>"001011011",
  31069=>"001001011",
  31070=>"001101111",
  31071=>"011010000",
  31072=>"000001101",
  31073=>"110110000",
  31074=>"101000100",
  31075=>"100010100",
  31076=>"100000100",
  31077=>"001000001",
  31078=>"110110000",
  31079=>"010111110",
  31080=>"111101000",
  31081=>"000111100",
  31082=>"111000100",
  31083=>"110001101",
  31084=>"100110111",
  31085=>"000110000",
  31086=>"111000000",
  31087=>"001101111",
  31088=>"100110101",
  31089=>"111001000",
  31090=>"100000000",
  31091=>"011000000",
  31092=>"111111000",
  31093=>"011000000",
  31094=>"001000010",
  31095=>"000010010",
  31096=>"000100111",
  31097=>"000100111",
  31098=>"000001000",
  31099=>"101000000",
  31100=>"110010110",
  31101=>"100101000",
  31102=>"110110010",
  31103=>"110110110",
  31104=>"001000000",
  31105=>"010000000",
  31106=>"011110101",
  31107=>"010011111",
  31108=>"111010000",
  31109=>"110000000",
  31110=>"011100111",
  31111=>"000000011",
  31112=>"011011010",
  31113=>"001101001",
  31114=>"011111010",
  31115=>"111000000",
  31116=>"000000000",
  31117=>"000000111",
  31118=>"000000000",
  31119=>"000000110",
  31120=>"010011001",
  31121=>"110000001",
  31122=>"001001001",
  31123=>"111011111",
  31124=>"011100011",
  31125=>"010000110",
  31126=>"111000000",
  31127=>"100100110",
  31128=>"011100101",
  31129=>"101111111",
  31130=>"001001111",
  31131=>"010110010",
  31132=>"111101111",
  31133=>"101111000",
  31134=>"111100011",
  31135=>"000000000",
  31136=>"001101110",
  31137=>"001000000",
  31138=>"001101010",
  31139=>"110111100",
  31140=>"010000101",
  31141=>"101100101",
  31142=>"000000001",
  31143=>"001000100",
  31144=>"110000001",
  31145=>"110111000",
  31146=>"111111111",
  31147=>"111000000",
  31148=>"001000010",
  31149=>"101100101",
  31150=>"000000100",
  31151=>"111111010",
  31152=>"000000010",
  31153=>"001001110",
  31154=>"000111111",
  31155=>"100000010",
  31156=>"011111010",
  31157=>"111111111",
  31158=>"000000100",
  31159=>"000000000",
  31160=>"001111111",
  31161=>"010101110",
  31162=>"011010011",
  31163=>"100010000",
  31164=>"110110111",
  31165=>"011010000",
  31166=>"011011001",
  31167=>"111111101",
  31168=>"110010111",
  31169=>"000000111",
  31170=>"000111110",
  31171=>"110111100",
  31172=>"000111000",
  31173=>"100100011",
  31174=>"000000010",
  31175=>"100000111",
  31176=>"111001001",
  31177=>"001000001",
  31178=>"001001001",
  31179=>"011111101",
  31180=>"000010111",
  31181=>"011000011",
  31182=>"010000111",
  31183=>"000100000",
  31184=>"000000100",
  31185=>"111111111",
  31186=>"001001000",
  31187=>"010100000",
  31188=>"000001111",
  31189=>"100101111",
  31190=>"111000000",
  31191=>"111000100",
  31192=>"100100111",
  31193=>"001110000",
  31194=>"101100100",
  31195=>"010010000",
  31196=>"001100011",
  31197=>"111101000",
  31198=>"010101001",
  31199=>"000000010",
  31200=>"101000111",
  31201=>"111000000",
  31202=>"000000000",
  31203=>"101100101",
  31204=>"010010000",
  31205=>"101101111",
  31206=>"000101111",
  31207=>"100000010",
  31208=>"001000000",
  31209=>"001110010",
  31210=>"011111001",
  31211=>"010110001",
  31212=>"101001000",
  31213=>"001111000",
  31214=>"000000000",
  31215=>"111101111",
  31216=>"000010010",
  31217=>"011010111",
  31218=>"111111000",
  31219=>"111101000",
  31220=>"111101110",
  31221=>"111000000",
  31222=>"000000001",
  31223=>"000000101",
  31224=>"111000110",
  31225=>"101000000",
  31226=>"011111110",
  31227=>"100101110",
  31228=>"000000101",
  31229=>"001111110",
  31230=>"000000001",
  31231=>"000011111",
  31232=>"001101100",
  31233=>"111000001",
  31234=>"000110000",
  31235=>"110101010",
  31236=>"111110010",
  31237=>"100001110",
  31238=>"001001111",
  31239=>"110100010",
  31240=>"100101111",
  31241=>"000001101",
  31242=>"000000001",
  31243=>"000101101",
  31244=>"111110010",
  31245=>"010011010",
  31246=>"011011011",
  31247=>"000001000",
  31248=>"110110000",
  31249=>"000100000",
  31250=>"000110111",
  31251=>"111111000",
  31252=>"111010000",
  31253=>"111111101",
  31254=>"011100011",
  31255=>"100110010",
  31256=>"111111101",
  31257=>"001000000",
  31258=>"000000101",
  31259=>"000001000",
  31260=>"000001010",
  31261=>"001101111",
  31262=>"001101110",
  31263=>"010000000",
  31264=>"000101011",
  31265=>"100111111",
  31266=>"000001000",
  31267=>"000000000",
  31268=>"011011000",
  31269=>"100100101",
  31270=>"000000000",
  31271=>"000001010",
  31272=>"111111111",
  31273=>"110110010",
  31274=>"000000000",
  31275=>"001000100",
  31276=>"111011011",
  31277=>"000100100",
  31278=>"000001001",
  31279=>"001011001",
  31280=>"000101101",
  31281=>"111111111",
  31282=>"000001000",
  31283=>"001001000",
  31284=>"000000011",
  31285=>"110000110",
  31286=>"000000001",
  31287=>"010111101",
  31288=>"001000001",
  31289=>"000110010",
  31290=>"100100011",
  31291=>"111111000",
  31292=>"100110000",
  31293=>"000001111",
  31294=>"000000000",
  31295=>"011001011",
  31296=>"110111110",
  31297=>"111001101",
  31298=>"111011010",
  31299=>"011001001",
  31300=>"000000000",
  31301=>"100010010",
  31302=>"000001001",
  31303=>"000101111",
  31304=>"011100111",
  31305=>"010011011",
  31306=>"000000000",
  31307=>"111000011",
  31308=>"000000100",
  31309=>"111111101",
  31310=>"111111011",
  31311=>"111111000",
  31312=>"001010000",
  31313=>"110110111",
  31314=>"100111010",
  31315=>"011110101",
  31316=>"000010110",
  31317=>"110100011",
  31318=>"000100000",
  31319=>"000000111",
  31320=>"011101011",
  31321=>"101100000",
  31322=>"111000010",
  31323=>"110110000",
  31324=>"000101001",
  31325=>"001001000",
  31326=>"111111001",
  31327=>"000000000",
  31328=>"111111110",
  31329=>"000000100",
  31330=>"001111110",
  31331=>"111010010",
  31332=>"100110110",
  31333=>"000000100",
  31334=>"000001101",
  31335=>"001101111",
  31336=>"000001100",
  31337=>"001000101",
  31338=>"000000111",
  31339=>"111111101",
  31340=>"000001000",
  31341=>"111110101",
  31342=>"001100001",
  31343=>"100010000",
  31344=>"101011110",
  31345=>"000001101",
  31346=>"010000100",
  31347=>"000010000",
  31348=>"010000101",
  31349=>"000101000",
  31350=>"010110111",
  31351=>"110110001",
  31352=>"000000000",
  31353=>"111110100",
  31354=>"100001011",
  31355=>"001101000",
  31356=>"110110101",
  31357=>"100100101",
  31358=>"000000111",
  31359=>"000010110",
  31360=>"111000000",
  31361=>"110110111",
  31362=>"000101101",
  31363=>"111111001",
  31364=>"100111110",
  31365=>"100010010",
  31366=>"011001001",
  31367=>"111110010",
  31368=>"011011111",
  31369=>"111001111",
  31370=>"101100000",
  31371=>"001011101",
  31372=>"011001001",
  31373=>"011001111",
  31374=>"000000000",
  31375=>"000001110",
  31376=>"101011010",
  31377=>"000001111",
  31378=>"100011101",
  31379=>"110111101",
  31380=>"111111101",
  31381=>"000000111",
  31382=>"011010110",
  31383=>"011011000",
  31384=>"000000100",
  31385=>"110000010",
  31386=>"000000101",
  31387=>"000000000",
  31388=>"011000000",
  31389=>"111111100",
  31390=>"001111111",
  31391=>"010010010",
  31392=>"111010111",
  31393=>"000000001",
  31394=>"111111000",
  31395=>"000000000",
  31396=>"001011100",
  31397=>"110110111",
  31398=>"100111110",
  31399=>"011000001",
  31400=>"111000000",
  31401=>"110110110",
  31402=>"101101101",
  31403=>"110110111",
  31404=>"111111111",
  31405=>"001001101",
  31406=>"001011001",
  31407=>"101111111",
  31408=>"000000000",
  31409=>"011011011",
  31410=>"101101101",
  31411=>"100000000",
  31412=>"111110110",
  31413=>"101111111",
  31414=>"101110000",
  31415=>"001001001",
  31416=>"011011011",
  31417=>"111110100",
  31418=>"000000100",
  31419=>"000001000",
  31420=>"001001101",
  31421=>"000010000",
  31422=>"000000000",
  31423=>"000001111",
  31424=>"000001111",
  31425=>"000100111",
  31426=>"000010011",
  31427=>"100100100",
  31428=>"111011001",
  31429=>"100111111",
  31430=>"000111010",
  31431=>"000000000",
  31432=>"000000000",
  31433=>"111010000",
  31434=>"000111111",
  31435=>"111110000",
  31436=>"001000100",
  31437=>"011011001",
  31438=>"000110110",
  31439=>"111111101",
  31440=>"000000111",
  31441=>"111110011",
  31442=>"000110110",
  31443=>"111111111",
  31444=>"000111111",
  31445=>"000000000",
  31446=>"000001001",
  31447=>"010101101",
  31448=>"110111011",
  31449=>"000101101",
  31450=>"111110111",
  31451=>"101001000",
  31452=>"110111111",
  31453=>"011001100",
  31454=>"000101000",
  31455=>"000001111",
  31456=>"011010010",
  31457=>"001001011",
  31458=>"101111110",
  31459=>"111100100",
  31460=>"000010010",
  31461=>"110011000",
  31462=>"101100011",
  31463=>"110100100",
  31464=>"000101000",
  31465=>"110111000",
  31466=>"000000000",
  31467=>"000001000",
  31468=>"111110000",
  31469=>"100111110",
  31470=>"000000000",
  31471=>"001001000",
  31472=>"101101100",
  31473=>"111100100",
  31474=>"000101001",
  31475=>"001001111",
  31476=>"011101110",
  31477=>"000000000",
  31478=>"001000000",
  31479=>"100101110",
  31480=>"000000000",
  31481=>"000000000",
  31482=>"111111101",
  31483=>"010111111",
  31484=>"000101101",
  31485=>"000000001",
  31486=>"110110101",
  31487=>"101111110",
  31488=>"000000000",
  31489=>"001101101",
  31490=>"111111001",
  31491=>"001000000",
  31492=>"010010001",
  31493=>"000111111",
  31494=>"011110111",
  31495=>"111000000",
  31496=>"000000000",
  31497=>"101000111",
  31498=>"000100011",
  31499=>"000000000",
  31500=>"001001011",
  31501=>"111101101",
  31502=>"011011011",
  31503=>"101111010",
  31504=>"000000000",
  31505=>"000000000",
  31506=>"110110000",
  31507=>"000000100",
  31508=>"111111011",
  31509=>"111111111",
  31510=>"010111111",
  31511=>"111111110",
  31512=>"001110000",
  31513=>"111001101",
  31514=>"111011100",
  31515=>"000111111",
  31516=>"111111110",
  31517=>"111111111",
  31518=>"000001111",
  31519=>"000010000",
  31520=>"000000000",
  31521=>"000001011",
  31522=>"001111111",
  31523=>"011001001",
  31524=>"111100100",
  31525=>"100001000",
  31526=>"001000000",
  31527=>"111110101",
  31528=>"111111111",
  31529=>"110110111",
  31530=>"000000001",
  31531=>"111111101",
  31532=>"011110010",
  31533=>"110000101",
  31534=>"000000000",
  31535=>"110011111",
  31536=>"000000000",
  31537=>"110000011",
  31538=>"000001001",
  31539=>"000010000",
  31540=>"101010000",
  31541=>"010111110",
  31542=>"110111110",
  31543=>"000001001",
  31544=>"000000000",
  31545=>"000000000",
  31546=>"100000111",
  31547=>"111111111",
  31548=>"100011011",
  31549=>"101101000",
  31550=>"000000111",
  31551=>"011111111",
  31552=>"000000000",
  31553=>"101000001",
  31554=>"010010011",
  31555=>"000000000",
  31556=>"111101111",
  31557=>"000110000",
  31558=>"101000000",
  31559=>"111111100",
  31560=>"111101100",
  31561=>"011111101",
  31562=>"101010010",
  31563=>"000000111",
  31564=>"000000110",
  31565=>"000000000",
  31566=>"100000100",
  31567=>"101000111",
  31568=>"001000000",
  31569=>"100010000",
  31570=>"000000111",
  31571=>"001001001",
  31572=>"111111111",
  31573=>"110101111",
  31574=>"111111111",
  31575=>"001000001",
  31576=>"001010110",
  31577=>"111111001",
  31578=>"111111111",
  31579=>"000001000",
  31580=>"000000000",
  31581=>"000001001",
  31582=>"111000000",
  31583=>"000000001",
  31584=>"000001011",
  31585=>"000000111",
  31586=>"011011000",
  31587=>"110111110",
  31588=>"000000000",
  31589=>"111001011",
  31590=>"010000011",
  31591=>"111111111",
  31592=>"000010000",
  31593=>"001000000",
  31594=>"000010000",
  31595=>"010010001",
  31596=>"011111011",
  31597=>"111110010",
  31598=>"110111101",
  31599=>"110101111",
  31600=>"000000000",
  31601=>"000000000",
  31602=>"001111011",
  31603=>"000000110",
  31604=>"000110110",
  31605=>"111000001",
  31606=>"000000000",
  31607=>"110111101",
  31608=>"111111001",
  31609=>"000001100",
  31610=>"000000000",
  31611=>"111111000",
  31612=>"000000000",
  31613=>"100100000",
  31614=>"111111110",
  31615=>"001000000",
  31616=>"111010111",
  31617=>"001000000",
  31618=>"111111000",
  31619=>"111100111",
  31620=>"011001000",
  31621=>"111111111",
  31622=>"111101011",
  31623=>"011011111",
  31624=>"000000000",
  31625=>"111001111",
  31626=>"000000000",
  31627=>"000101101",
  31628=>"111101110",
  31629=>"101111111",
  31630=>"000000010",
  31631=>"000000001",
  31632=>"110011000",
  31633=>"000111001",
  31634=>"111011000",
  31635=>"000001001",
  31636=>"000010010",
  31637=>"000000011",
  31638=>"010000000",
  31639=>"000000000",
  31640=>"000111001",
  31641=>"111111101",
  31642=>"110110000",
  31643=>"000110010",
  31644=>"000000000",
  31645=>"000000101",
  31646=>"000000000",
  31647=>"000000000",
  31648=>"111111011",
  31649=>"100111111",
  31650=>"111000000",
  31651=>"011111111",
  31652=>"000000111",
  31653=>"111101000",
  31654=>"000000000",
  31655=>"000000011",
  31656=>"111100110",
  31657=>"000001000",
  31658=>"000001000",
  31659=>"000000000",
  31660=>"110100101",
  31661=>"000000000",
  31662=>"000110000",
  31663=>"111111111",
  31664=>"001101111",
  31665=>"010000100",
  31666=>"110110110",
  31667=>"100100111",
  31668=>"111111111",
  31669=>"010110111",
  31670=>"111100101",
  31671=>"000000110",
  31672=>"001110110",
  31673=>"010100000",
  31674=>"001111111",
  31675=>"000001001",
  31676=>"111111111",
  31677=>"111010000",
  31678=>"000110111",
  31679=>"000000101",
  31680=>"111111100",
  31681=>"111111111",
  31682=>"110111111",
  31683=>"000001111",
  31684=>"111000000",
  31685=>"001010111",
  31686=>"000000100",
  31687=>"111111100",
  31688=>"111000000",
  31689=>"111001000",
  31690=>"000100011",
  31691=>"001000000",
  31692=>"000010011",
  31693=>"000100100",
  31694=>"111111111",
  31695=>"101111111",
  31696=>"010110110",
  31697=>"011011000",
  31698=>"000001000",
  31699=>"010010000",
  31700=>"000000000",
  31701=>"000000011",
  31702=>"000010000",
  31703=>"000000100",
  31704=>"111101111",
  31705=>"000000000",
  31706=>"111111111",
  31707=>"111000000",
  31708=>"000000010",
  31709=>"000000001",
  31710=>"111000101",
  31711=>"100000000",
  31712=>"111111111",
  31713=>"000000000",
  31714=>"110111110",
  31715=>"010100110",
  31716=>"000000000",
  31717=>"000100111",
  31718=>"000000000",
  31719=>"010111111",
  31720=>"000010000",
  31721=>"001100110",
  31722=>"000000101",
  31723=>"001111000",
  31724=>"000000001",
  31725=>"000000111",
  31726=>"000000000",
  31727=>"000000111",
  31728=>"111111111",
  31729=>"100111111",
  31730=>"000000000",
  31731=>"001011000",
  31732=>"101100111",
  31733=>"111111111",
  31734=>"000011001",
  31735=>"111111111",
  31736=>"000000111",
  31737=>"101111111",
  31738=>"100100000",
  31739=>"000100001",
  31740=>"111111111",
  31741=>"111101001",
  31742=>"010010000",
  31743=>"111110110",
  31744=>"010110010",
  31745=>"001001001",
  31746=>"110110110",
  31747=>"000011111",
  31748=>"101111111",
  31749=>"000000110",
  31750=>"000101001",
  31751=>"001001001",
  31752=>"000001001",
  31753=>"000000111",
  31754=>"110110100",
  31755=>"001000011",
  31756=>"110110111",
  31757=>"010000010",
  31758=>"100101000",
  31759=>"110111111",
  31760=>"010001011",
  31761=>"110000111",
  31762=>"000110000",
  31763=>"000001001",
  31764=>"011011011",
  31765=>"001100100",
  31766=>"001000000",
  31767=>"110110100",
  31768=>"110110010",
  31769=>"010110110",
  31770=>"000000010",
  31771=>"000001011",
  31772=>"010011110",
  31773=>"100000000",
  31774=>"001111111",
  31775=>"001000000",
  31776=>"110110110",
  31777=>"001001000",
  31778=>"101010000",
  31779=>"000010000",
  31780=>"000001001",
  31781=>"100010010",
  31782=>"011110110",
  31783=>"011011011",
  31784=>"111111101",
  31785=>"000000110",
  31786=>"011000011",
  31787=>"010111011",
  31788=>"001010010",
  31789=>"111001100",
  31790=>"010000001",
  31791=>"011011011",
  31792=>"011001000",
  31793=>"100100101",
  31794=>"101000000",
  31795=>"111111010",
  31796=>"111000001",
  31797=>"011000010",
  31798=>"111111001",
  31799=>"011011011",
  31800=>"001011001",
  31801=>"011001000",
  31802=>"001111000",
  31803=>"011011010",
  31804=>"000011001",
  31805=>"111011101",
  31806=>"100100011",
  31807=>"000001001",
  31808=>"111110110",
  31809=>"010011111",
  31810=>"110100000",
  31811=>"010110100",
  31812=>"000100111",
  31813=>"001111110",
  31814=>"011000001",
  31815=>"100100100",
  31816=>"011111111",
  31817=>"001001001",
  31818=>"011010111",
  31819=>"001011000",
  31820=>"110100000",
  31821=>"011011010",
  31822=>"010010110",
  31823=>"111011010",
  31824=>"011000000",
  31825=>"001110000",
  31826=>"001001000",
  31827=>"001000000",
  31828=>"001000111",
  31829=>"110010011",
  31830=>"101111011",
  31831=>"100100110",
  31832=>"100100110",
  31833=>"000000000",
  31834=>"000011001",
  31835=>"001000000",
  31836=>"000001011",
  31837=>"000100000",
  31838=>"101101100",
  31839=>"110100110",
  31840=>"111100110",
  31841=>"111111010",
  31842=>"100110110",
  31843=>"001011011",
  31844=>"011011001",
  31845=>"011001001",
  31846=>"000001001",
  31847=>"011001001",
  31848=>"001001011",
  31849=>"101100111",
  31850=>"111111000",
  31851=>"100111100",
  31852=>"110111000",
  31853=>"100110100",
  31854=>"011100001",
  31855=>"011001011",
  31856=>"011111000",
  31857=>"011000011",
  31858=>"011001111",
  31859=>"100110110",
  31860=>"111010010",
  31861=>"000110001",
  31862=>"011000000",
  31863=>"001101000",
  31864=>"001111011",
  31865=>"001001001",
  31866=>"111001000",
  31867=>"100100110",
  31868=>"111011100",
  31869=>"000000001",
  31870=>"110101001",
  31871=>"001000100",
  31872=>"011110100",
  31873=>"111110110",
  31874=>"001001001",
  31875=>"000111011",
  31876=>"011011011",
  31877=>"011011111",
  31878=>"011001011",
  31879=>"000000000",
  31880=>"000000000",
  31881=>"000011000",
  31882=>"000001011",
  31883=>"100000010",
  31884=>"111110100",
  31885=>"011001100",
  31886=>"000001001",
  31887=>"010000011",
  31888=>"010010010",
  31889=>"010111011",
  31890=>"011000000",
  31891=>"010000010",
  31892=>"000001001",
  31893=>"110110110",
  31894=>"000001000",
  31895=>"001111011",
  31896=>"111011000",
  31897=>"101001001",
  31898=>"100100111",
  31899=>"111111111",
  31900=>"001001001",
  31901=>"000000111",
  31902=>"001001001",
  31903=>"110110111",
  31904=>"010000000",
  31905=>"111000111",
  31906=>"111111110",
  31907=>"000010010",
  31908=>"111011001",
  31909=>"111111100",
  31910=>"010000011",
  31911=>"011001000",
  31912=>"110000010",
  31913=>"000001000",
  31914=>"111110111",
  31915=>"100110110",
  31916=>"111000000",
  31917=>"000001001",
  31918=>"001001011",
  31919=>"001101101",
  31920=>"111011001",
  31921=>"111111000",
  31922=>"111100100",
  31923=>"110001100",
  31924=>"100000101",
  31925=>"101001001",
  31926=>"000010010",
  31927=>"001010011",
  31928=>"001001000",
  31929=>"000011010",
  31930=>"010011001",
  31931=>"100100001",
  31932=>"001001000",
  31933=>"110110110",
  31934=>"000000000",
  31935=>"001110111",
  31936=>"010011001",
  31937=>"000000001",
  31938=>"111100000",
  31939=>"100101001",
  31940=>"001000000",
  31941=>"111011111",
  31942=>"000010011",
  31943=>"100110010",
  31944=>"010001000",
  31945=>"100100110",
  31946=>"100100000",
  31947=>"000101101",
  31948=>"001001011",
  31949=>"001001001",
  31950=>"001000001",
  31951=>"111110100",
  31952=>"111110110",
  31953=>"100001101",
  31954=>"010001011",
  31955=>"100000011",
  31956=>"111111011",
  31957=>"111010111",
  31958=>"101100110",
  31959=>"000001011",
  31960=>"011011001",
  31961=>"000011001",
  31962=>"111111111",
  31963=>"110110110",
  31964=>"111111011",
  31965=>"111110110",
  31966=>"001001000",
  31967=>"011001001",
  31968=>"100100111",
  31969=>"111110110",
  31970=>"100101100",
  31971=>"000000000",
  31972=>"000001000",
  31973=>"100100100",
  31974=>"001000100",
  31975=>"101111001",
  31976=>"100101111",
  31977=>"100110110",
  31978=>"110100100",
  31979=>"110100000",
  31980=>"100100110",
  31981=>"001000011",
  31982=>"000110010",
  31983=>"001011011",
  31984=>"000110010",
  31985=>"010000111",
  31986=>"000011011",
  31987=>"011011111",
  31988=>"000000011",
  31989=>"000101000",
  31990=>"100100011",
  31991=>"000001011",
  31992=>"011110111",
  31993=>"001001011",
  31994=>"110110110",
  31995=>"011110100",
  31996=>"011011111",
  31997=>"100001101",
  31998=>"001001000",
  31999=>"001101001",
  32000=>"011001000",
  32001=>"000000111",
  32002=>"000000000",
  32003=>"000110111",
  32004=>"000000100",
  32005=>"000011010",
  32006=>"001001101",
  32007=>"101000110",
  32008=>"000001011",
  32009=>"000001111",
  32010=>"010100110",
  32011=>"110101101",
  32012=>"011011100",
  32013=>"110001000",
  32014=>"101001001",
  32015=>"000000011",
  32016=>"110111000",
  32017=>"110000000",
  32018=>"001000010",
  32019=>"101111111",
  32020=>"001111010",
  32021=>"111111111",
  32022=>"011100001",
  32023=>"111111010",
  32024=>"000100100",
  32025=>"101000000",
  32026=>"000000000",
  32027=>"011010100",
  32028=>"000100111",
  32029=>"000111111",
  32030=>"111000000",
  32031=>"001111111",
  32032=>"110111000",
  32033=>"000100000",
  32034=>"111000101",
  32035=>"110110111",
  32036=>"110111111",
  32037=>"110100000",
  32038=>"010111010",
  32039=>"010000001",
  32040=>"111111000",
  32041=>"111111000",
  32042=>"101001000",
  32043=>"101000101",
  32044=>"110100111",
  32045=>"000000110",
  32046=>"000111110",
  32047=>"001001011",
  32048=>"101101011",
  32049=>"001101001",
  32050=>"000110111",
  32051=>"101000001",
  32052=>"001000101",
  32053=>"000101110",
  32054=>"110111111",
  32055=>"000000111",
  32056=>"110010101",
  32057=>"001110100",
  32058=>"100100100",
  32059=>"111101111",
  32060=>"000010000",
  32061=>"111111000",
  32062=>"011000001",
  32063=>"011111111",
  32064=>"100000000",
  32065=>"100000000",
  32066=>"101111111",
  32067=>"101110100",
  32068=>"100100010",
  32069=>"011000010",
  32070=>"001000110",
  32071=>"100111100",
  32072=>"000000011",
  32073=>"110111010",
  32074=>"000000000",
  32075=>"001000001",
  32076=>"001000111",
  32077=>"011111010",
  32078=>"101101110",
  32079=>"000000111",
  32080=>"111111000",
  32081=>"001011000",
  32082=>"011111010",
  32083=>"011000100",
  32084=>"101101000",
  32085=>"001000011",
  32086=>"011001001",
  32087=>"111110010",
  32088=>"110100100",
  32089=>"111111111",
  32090=>"100101001",
  32091=>"111011110",
  32092=>"000000000",
  32093=>"001001001",
  32094=>"111111110",
  32095=>"110011011",
  32096=>"000000000",
  32097=>"011010010",
  32098=>"010000000",
  32099=>"100111001",
  32100=>"110111000",
  32101=>"010011011",
  32102=>"000001111",
  32103=>"000101111",
  32104=>"000010001",
  32105=>"000110010",
  32106=>"010000111",
  32107=>"010000000",
  32108=>"000000000",
  32109=>"000000000",
  32110=>"001001010",
  32111=>"000001010",
  32112=>"100100101",
  32113=>"010000101",
  32114=>"000111111",
  32115=>"101000101",
  32116=>"010010111",
  32117=>"000000000",
  32118=>"000110111",
  32119=>"111111111",
  32120=>"000000010",
  32121=>"111001000",
  32122=>"000000110",
  32123=>"110111000",
  32124=>"000110111",
  32125=>"110100100",
  32126=>"010101101",
  32127=>"111111001",
  32128=>"100000111",
  32129=>"111000000",
  32130=>"111000010",
  32131=>"001010010",
  32132=>"011010010",
  32133=>"111101001",
  32134=>"000011000",
  32135=>"011000000",
  32136=>"101101011",
  32137=>"111000000",
  32138=>"000010110",
  32139=>"110000111",
  32140=>"001000000",
  32141=>"101111011",
  32142=>"011111010",
  32143=>"101001101",
  32144=>"100111110",
  32145=>"010000000",
  32146=>"101000101",
  32147=>"111000000",
  32148=>"111111001",
  32149=>"110110000",
  32150=>"010111101",
  32151=>"111011011",
  32152=>"000000111",
  32153=>"000000010",
  32154=>"000001101",
  32155=>"111111111",
  32156=>"111011010",
  32157=>"100111010",
  32158=>"000010111",
  32159=>"001000101",
  32160=>"100110110",
  32161=>"111010100",
  32162=>"110111000",
  32163=>"011100101",
  32164=>"111000000",
  32165=>"111001011",
  32166=>"111110110",
  32167=>"010000111",
  32168=>"010100000",
  32169=>"101000110",
  32170=>"110111111",
  32171=>"000000000",
  32172=>"001000000",
  32173=>"111110000",
  32174=>"110101110",
  32175=>"010111110",
  32176=>"000000000",
  32177=>"110000000",
  32178=>"111000000",
  32179=>"000100110",
  32180=>"011011111",
  32181=>"101100010",
  32182=>"010000000",
  32183=>"011010000",
  32184=>"000010010",
  32185=>"110110100",
  32186=>"111101000",
  32187=>"110011111",
  32188=>"000000000",
  32189=>"100110000",
  32190=>"110110110",
  32191=>"000110100",
  32192=>"000010010",
  32193=>"000000001",
  32194=>"110110100",
  32195=>"100110110",
  32196=>"101000000",
  32197=>"001001011",
  32198=>"000100000",
  32199=>"101000000",
  32200=>"011110001",
  32201=>"101000001",
  32202=>"000000100",
  32203=>"000111000",
  32204=>"000000000",
  32205=>"000011011",
  32206=>"011101111",
  32207=>"111110000",
  32208=>"010010010",
  32209=>"110110110",
  32210=>"111111101",
  32211=>"000000111",
  32212=>"011000001",
  32213=>"000000110",
  32214=>"000110011",
  32215=>"000111111",
  32216=>"000000111",
  32217=>"011111111",
  32218=>"011001000",
  32219=>"100000000",
  32220=>"000001100",
  32221=>"001000011",
  32222=>"000000000",
  32223=>"110100000",
  32224=>"001001111",
  32225=>"000000001",
  32226=>"110111010",
  32227=>"110010000",
  32228=>"101000001",
  32229=>"000000111",
  32230=>"000000100",
  32231=>"010011001",
  32232=>"000001100",
  32233=>"000000000",
  32234=>"100001001",
  32235=>"111001001",
  32236=>"010010010",
  32237=>"111000000",
  32238=>"000000000",
  32239=>"001000000",
  32240=>"111111111",
  32241=>"100100000",
  32242=>"011101100",
  32243=>"001001110",
  32244=>"110000001",
  32245=>"000111000",
  32246=>"110000000",
  32247=>"101101111",
  32248=>"011000111",
  32249=>"010000110",
  32250=>"000010010",
  32251=>"000000010",
  32252=>"011111010",
  32253=>"100111110",
  32254=>"110111111",
  32255=>"111000000",
  32256=>"000000110",
  32257=>"111000010",
  32258=>"000100110",
  32259=>"111000100",
  32260=>"111011011",
  32261=>"000010011",
  32262=>"000000111",
  32263=>"110111011",
  32264=>"000101001",
  32265=>"101000000",
  32266=>"100001000",
  32267=>"101001011",
  32268=>"000110111",
  32269=>"011001111",
  32270=>"100011001",
  32271=>"000000000",
  32272=>"100010110",
  32273=>"001000000",
  32274=>"000111000",
  32275=>"111111001",
  32276=>"000100011",
  32277=>"111111010",
  32278=>"100111001",
  32279=>"010010010",
  32280=>"111001101",
  32281=>"111111111",
  32282=>"000101111",
  32283=>"101101101",
  32284=>"101101101",
  32285=>"000000000",
  32286=>"000000000",
  32287=>"000000000",
  32288=>"110111000",
  32289=>"101101111",
  32290=>"000010000",
  32291=>"001011010",
  32292=>"001101111",
  32293=>"101101110",
  32294=>"011001000",
  32295=>"110000001",
  32296=>"101101011",
  32297=>"110011000",
  32298=>"000000000",
  32299=>"111111101",
  32300=>"001111110",
  32301=>"000000110",
  32302=>"000111111",
  32303=>"111101010",
  32304=>"000111010",
  32305=>"001100101",
  32306=>"000010100",
  32307=>"000000010",
  32308=>"000000000",
  32309=>"111111110",
  32310=>"100000000",
  32311=>"011110000",
  32312=>"000011101",
  32313=>"000000101",
  32314=>"111010000",
  32315=>"000001011",
  32316=>"110110111",
  32317=>"000111011",
  32318=>"100000101",
  32319=>"100000111",
  32320=>"000000000",
  32321=>"111101111",
  32322=>"111101111",
  32323=>"101000000",
  32324=>"000000011",
  32325=>"000010000",
  32326=>"000000001",
  32327=>"001000101",
  32328=>"000100111",
  32329=>"000101111",
  32330=>"010111101",
  32331=>"010011000",
  32332=>"000001101",
  32333=>"110100110",
  32334=>"101001011",
  32335=>"111110111",
  32336=>"001000000",
  32337=>"011111111",
  32338=>"100101001",
  32339=>"001111111",
  32340=>"101000000",
  32341=>"001111110",
  32342=>"000011011",
  32343=>"111000010",
  32344=>"000001000",
  32345=>"000100100",
  32346=>"111110000",
  32347=>"111101001",
  32348=>"000000101",
  32349=>"000000000",
  32350=>"000001010",
  32351=>"000011001",
  32352=>"111101101",
  32353=>"000000111",
  32354=>"101101101",
  32355=>"111000000",
  32356=>"000100000",
  32357=>"101100110",
  32358=>"010010000",
  32359=>"111101000",
  32360=>"111000001",
  32361=>"000000100",
  32362=>"000100101",
  32363=>"000001111",
  32364=>"110111011",
  32365=>"001100110",
  32366=>"000100010",
  32367=>"011010001",
  32368=>"001001111",
  32369=>"000000100",
  32370=>"001000001",
  32371=>"110010000",
  32372=>"001000000",
  32373=>"000000001",
  32374=>"010101101",
  32375=>"001110111",
  32376=>"111000000",
  32377=>"000111111",
  32378=>"000000000",
  32379=>"000000001",
  32380=>"001110100",
  32381=>"000001111",
  32382=>"000000011",
  32383=>"100110111",
  32384=>"111000010",
  32385=>"000111111",
  32386=>"001111111",
  32387=>"111000001",
  32388=>"000000100",
  32389=>"111001111",
  32390=>"101101011",
  32391=>"111100011",
  32392=>"100100110",
  32393=>"000101000",
  32394=>"111011011",
  32395=>"000001111",
  32396=>"000000000",
  32397=>"111010000",
  32398=>"000100100",
  32399=>"001000000",
  32400=>"100111010",
  32401=>"111101000",
  32402=>"000000101",
  32403=>"000000000",
  32404=>"110100100",
  32405=>"000000111",
  32406=>"000010110",
  32407=>"010011000",
  32408=>"111111001",
  32409=>"111101000",
  32410=>"100000100",
  32411=>"111000000",
  32412=>"000111011",
  32413=>"111100000",
  32414=>"100101011",
  32415=>"010111101",
  32416=>"101111111",
  32417=>"010100000",
  32418=>"000111111",
  32419=>"111101101",
  32420=>"111011000",
  32421=>"101111111",
  32422=>"111110100",
  32423=>"111001011",
  32424=>"111000011",
  32425=>"000000100",
  32426=>"111100010",
  32427=>"000000000",
  32428=>"011010000",
  32429=>"101101101",
  32430=>"100001001",
  32431=>"000111111",
  32432=>"110100000",
  32433=>"111111110",
  32434=>"101111111",
  32435=>"001001000",
  32436=>"001011001",
  32437=>"010010000",
  32438=>"111111111",
  32439=>"101001100",
  32440=>"111111111",
  32441=>"111011110",
  32442=>"111110011",
  32443=>"010000010",
  32444=>"101101111",
  32445=>"111111010",
  32446=>"000001011",
  32447=>"110100000",
  32448=>"000000100",
  32449=>"000000101",
  32450=>"101101111",
  32451=>"100100110",
  32452=>"000111110",
  32453=>"100100001",
  32454=>"000000011",
  32455=>"000010101",
  32456=>"000000111",
  32457=>"110011010",
  32458=>"111111111",
  32459=>"111111010",
  32460=>"111111000",
  32461=>"100101001",
  32462=>"100010000",
  32463=>"111101001",
  32464=>"100110100",
  32465=>"111111010",
  32466=>"011000101",
  32467=>"000111111",
  32468=>"000000000",
  32469=>"110110110",
  32470=>"000000101",
  32471=>"101111000",
  32472=>"010000000",
  32473=>"000000101",
  32474=>"101110111",
  32475=>"010000000",
  32476=>"100100001",
  32477=>"111111010",
  32478=>"111101001",
  32479=>"000000111",
  32480=>"111000011",
  32481=>"101101101",
  32482=>"101001000",
  32483=>"001001110",
  32484=>"010111111",
  32485=>"000110010",
  32486=>"000000000",
  32487=>"010111000",
  32488=>"000100100",
  32489=>"010111101",
  32490=>"000000000",
  32491=>"000010111",
  32492=>"100111111",
  32493=>"111101111",
  32494=>"000000001",
  32495=>"000110000",
  32496=>"000110000",
  32497=>"000000100",
  32498=>"110011001",
  32499=>"100000010",
  32500=>"000011000",
  32501=>"101101000",
  32502=>"010000100",
  32503=>"111101000",
  32504=>"001101110",
  32505=>"111000000",
  32506=>"111101111",
  32507=>"000110101",
  32508=>"000100111",
  32509=>"101101010",
  32510=>"011011011",
  32511=>"110111111",
  32512=>"000001001",
  32513=>"111000000",
  32514=>"001000001",
  32515=>"000000001",
  32516=>"110111111",
  32517=>"111111110",
  32518=>"000010011",
  32519=>"110101000",
  32520=>"111111111",
  32521=>"101001000",
  32522=>"110110010",
  32523=>"101010110",
  32524=>"000000000",
  32525=>"000000101",
  32526=>"100111111",
  32527=>"100000000",
  32528=>"111100000",
  32529=>"000111111",
  32530=>"000100101",
  32531=>"111001100",
  32532=>"111111000",
  32533=>"101001111",
  32534=>"000010000",
  32535=>"110111111",
  32536=>"101000111",
  32537=>"111110001",
  32538=>"101101111",
  32539=>"000000000",
  32540=>"110101000",
  32541=>"110000001",
  32542=>"001101110",
  32543=>"010010000",
  32544=>"010110000",
  32545=>"000010000",
  32546=>"010010111",
  32547=>"111111111",
  32548=>"011111110",
  32549=>"001011001",
  32550=>"100001000",
  32551=>"001111011",
  32552=>"000010000",
  32553=>"000001001",
  32554=>"111000010",
  32555=>"111111110",
  32556=>"111110111",
  32557=>"111110001",
  32558=>"010110010",
  32559=>"010010010",
  32560=>"011010111",
  32561=>"111111100",
  32562=>"000000000",
  32563=>"010011000",
  32564=>"110111101",
  32565=>"001100011",
  32566=>"111111000",
  32567=>"000000000",
  32568=>"111111111",
  32569=>"000001111",
  32570=>"010000101",
  32571=>"011111111",
  32572=>"110111011",
  32573=>"110111111",
  32574=>"001000101",
  32575=>"000111111",
  32576=>"000101001",
  32577=>"101001111",
  32578=>"000101000",
  32579=>"100111011",
  32580=>"001000101",
  32581=>"000101101",
  32582=>"110101111",
  32583=>"000000100",
  32584=>"000001111",
  32585=>"011110111",
  32586=>"001101111",
  32587=>"101000000",
  32588=>"000000000",
  32589=>"010101001",
  32590=>"001111111",
  32591=>"010000000",
  32592=>"101100101",
  32593=>"010111111",
  32594=>"010011111",
  32595=>"011001000",
  32596=>"101000000",
  32597=>"111000000",
  32598=>"110111011",
  32599=>"101110101",
  32600=>"101001101",
  32601=>"001001000",
  32602=>"111111101",
  32603=>"111111011",
  32604=>"000000001",
  32605=>"000000111",
  32606=>"000000000",
  32607=>"011111100",
  32608=>"101101111",
  32609=>"000010110",
  32610=>"000000000",
  32611=>"110111100",
  32612=>"000110010",
  32613=>"000000011",
  32614=>"110111111",
  32615=>"111111000",
  32616=>"010010111",
  32617=>"000010111",
  32618=>"000100000",
  32619=>"110110111",
  32620=>"000110111",
  32621=>"010111010",
  32622=>"000000111",
  32623=>"000011111",
  32624=>"010110010",
  32625=>"001000111",
  32626=>"111111001",
  32627=>"100111000",
  32628=>"111011010",
  32629=>"000000000",
  32630=>"101101111",
  32631=>"000000111",
  32632=>"001001000",
  32633=>"000001111",
  32634=>"111111111",
  32635=>"111000111",
  32636=>"011011111",
  32637=>"010100000",
  32638=>"001010010",
  32639=>"111010101",
  32640=>"110101010",
  32641=>"111100110",
  32642=>"111110000",
  32643=>"001000111",
  32644=>"000000000",
  32645=>"011111111",
  32646=>"101110100",
  32647=>"000110111",
  32648=>"011111101",
  32649=>"010111001",
  32650=>"000000000",
  32651=>"000111001",
  32652=>"000110111",
  32653=>"010110110",
  32654=>"101100100",
  32655=>"000001011",
  32656=>"111001101",
  32657=>"011010110",
  32658=>"011111010",
  32659=>"100100111",
  32660=>"111111010",
  32661=>"111110001",
  32662=>"000000000",
  32663=>"110110110",
  32664=>"111001111",
  32665=>"001000001",
  32666=>"111010000",
  32667=>"111111000",
  32668=>"110101001",
  32669=>"100110101",
  32670=>"110000010",
  32671=>"101000101",
  32672=>"101100010",
  32673=>"000000110",
  32674=>"101000101",
  32675=>"000000001",
  32676=>"000000000",
  32677=>"110111111",
  32678=>"011011011",
  32679=>"000000101",
  32680=>"111111011",
  32681=>"000100111",
  32682=>"101000100",
  32683=>"111000000",
  32684=>"101010000",
  32685=>"000101111",
  32686=>"000000100",
  32687=>"000000000",
  32688=>"000101101",
  32689=>"000011111",
  32690=>"000100000",
  32691=>"100111111",
  32692=>"110110111",
  32693=>"000000000",
  32694=>"111111101",
  32695=>"000101000",
  32696=>"110110110",
  32697=>"110011011",
  32698=>"011010100",
  32699=>"000110111",
  32700=>"010111111",
  32701=>"111111100",
  32702=>"000101111",
  32703=>"001000111",
  32704=>"000011110",
  32705=>"001000111",
  32706=>"001111110",
  32707=>"000010010",
  32708=>"010111111",
  32709=>"011000000",
  32710=>"111111111",
  32711=>"001000000",
  32712=>"111101111",
  32713=>"100001000",
  32714=>"111111011",
  32715=>"001101111",
  32716=>"000010000",
  32717=>"010111101",
  32718=>"111111111",
  32719=>"111110100",
  32720=>"010000000",
  32721=>"111011011",
  32722=>"110011011",
  32723=>"001001000",
  32724=>"111110000",
  32725=>"000001011",
  32726=>"100000001",
  32727=>"111111110",
  32728=>"001111011",
  32729=>"000111000",
  32730=>"100000000",
  32731=>"000000110",
  32732=>"000000000",
  32733=>"101101111",
  32734=>"111111011",
  32735=>"001000111",
  32736=>"000000000",
  32737=>"100001101",
  32738=>"000010000",
  32739=>"101101111",
  32740=>"011111011",
  32741=>"000111011",
  32742=>"010111111",
  32743=>"000000000",
  32744=>"000011111",
  32745=>"111110000",
  32746=>"001011011",
  32747=>"001111111",
  32748=>"101100101",
  32749=>"101100101",
  32750=>"000010010",
  32751=>"111010110",
  32752=>"111111111",
  32753=>"111001000",
  32754=>"000010010",
  32755=>"110100000",
  32756=>"010010110",
  32757=>"111011111",
  32758=>"110000011",
  32759=>"111111111",
  32760=>"101100011",
  32761=>"010010000",
  32762=>"011111111",
  32763=>"010011101",
  32764=>"000000000",
  32765=>"110111100",
  32766=>"001000001",
  32767=>"010101000",
  32768=>"010010101",
  32769=>"010111011",
  32770=>"111000001",
  32771=>"111111001",
  32772=>"001001001",
  32773=>"111110001",
  32774=>"000010000",
  32775=>"000111111",
  32776=>"000000110",
  32777=>"000100100",
  32778=>"101101111",
  32779=>"101000001",
  32780=>"000100100",
  32781=>"010000000",
  32782=>"111111101",
  32783=>"110110001",
  32784=>"100110110",
  32785=>"110000000",
  32786=>"000000000",
  32787=>"101101101",
  32788=>"111100000",
  32789=>"000000000",
  32790=>"110111011",
  32791=>"110010000",
  32792=>"000000000",
  32793=>"010100000",
  32794=>"110111111",
  32795=>"111111010",
  32796=>"000000000",
  32797=>"000010000",
  32798=>"111111111",
  32799=>"000000000",
  32800=>"100001000",
  32801=>"111111101",
  32802=>"000000001",
  32803=>"010011111",
  32804=>"001011001",
  32805=>"100111001",
  32806=>"010111110",
  32807=>"111101111",
  32808=>"101111101",
  32809=>"000111111",
  32810=>"111111110",
  32811=>"000000000",
  32812=>"111111110",
  32813=>"001000000",
  32814=>"010010111",
  32815=>"011001101",
  32816=>"111011111",
  32817=>"100100100",
  32818=>"000110110",
  32819=>"110110111",
  32820=>"111111011",
  32821=>"000000000",
  32822=>"000111101",
  32823=>"111111010",
  32824=>"111000000",
  32825=>"000000010",
  32826=>"000001000",
  32827=>"111101100",
  32828=>"010000001",
  32829=>"101111111",
  32830=>"001000001",
  32831=>"100111000",
  32832=>"111000110",
  32833=>"110101111",
  32834=>"011111111",
  32835=>"011011110",
  32836=>"000000110",
  32837=>"000000010",
  32838=>"101000001",
  32839=>"111000000",
  32840=>"000001000",
  32841=>"101001000",
  32842=>"000000000",
  32843=>"111111110",
  32844=>"111000000",
  32845=>"000000100",
  32846=>"001000000",
  32847=>"111000000",
  32848=>"110110000",
  32849=>"000111111",
  32850=>"000001100",
  32851=>"000000000",
  32852=>"010010000",
  32853=>"100111100",
  32854=>"011001100",
  32855=>"000001000",
  32856=>"000000001",
  32857=>"010100100",
  32858=>"111111001",
  32859=>"100100100",
  32860=>"010110110",
  32861=>"111001001",
  32862=>"111000000",
  32863=>"110100111",
  32864=>"010110110",
  32865=>"110000000",
  32866=>"000001000",
  32867=>"110110000",
  32868=>"101101110",
  32869=>"000000001",
  32870=>"101101111",
  32871=>"111111000",
  32872=>"111110111",
  32873=>"000000111",
  32874=>"111111010",
  32875=>"010100110",
  32876=>"010111111",
  32877=>"111111111",
  32878=>"111000101",
  32879=>"111111011",
  32880=>"001001001",
  32881=>"111001111",
  32882=>"000111111",
  32883=>"001001000",
  32884=>"010111000",
  32885=>"000000111",
  32886=>"111111101",
  32887=>"010000000",
  32888=>"111101001",
  32889=>"110000000",
  32890=>"001111101",
  32891=>"000000101",
  32892=>"101001100",
  32893=>"000100010",
  32894=>"101000000",
  32895=>"011110110",
  32896=>"000000000",
  32897=>"000000000",
  32898=>"100000111",
  32899=>"111111000",
  32900=>"000110110",
  32901=>"000000110",
  32902=>"011111000",
  32903=>"000001000",
  32904=>"100100100",
  32905=>"000000101",
  32906=>"111101111",
  32907=>"010111111",
  32908=>"111000000",
  32909=>"000000000",
  32910=>"011011000",
  32911=>"110011100",
  32912=>"010111011",
  32913=>"100110110",
  32914=>"110010010",
  32915=>"110010111",
  32916=>"010010111",
  32917=>"101001000",
  32918=>"110111111",
  32919=>"111010011",
  32920=>"111111111",
  32921=>"110010001",
  32922=>"101101011",
  32923=>"001001100",
  32924=>"111010000",
  32925=>"000001000",
  32926=>"111111011",
  32927=>"100111110",
  32928=>"110100010",
  32929=>"111000010",
  32930=>"010110111",
  32931=>"110001001",
  32932=>"100001111",
  32933=>"000000000",
  32934=>"010111000",
  32935=>"111111111",
  32936=>"110000100",
  32937=>"111111111",
  32938=>"001000101",
  32939=>"111010001",
  32940=>"111100000",
  32941=>"110111000",
  32942=>"000000011",
  32943=>"111001000",
  32944=>"111111111",
  32945=>"100110101",
  32946=>"011010000",
  32947=>"011001100",
  32948=>"110010000",
  32949=>"111101111",
  32950=>"000000000",
  32951=>"011111111",
  32952=>"001000000",
  32953=>"100110100",
  32954=>"111000000",
  32955=>"111011000",
  32956=>"011000110",
  32957=>"000110111",
  32958=>"110110010",
  32959=>"000000000",
  32960=>"000000000",
  32961=>"111001010",
  32962=>"111010111",
  32963=>"100101110",
  32964=>"000000010",
  32965=>"011010001",
  32966=>"000000000",
  32967=>"101000000",
  32968=>"000000000",
  32969=>"000000000",
  32970=>"000000001",
  32971=>"100001101",
  32972=>"111111110",
  32973=>"011000000",
  32974=>"110110001",
  32975=>"000000000",
  32976=>"010000000",
  32977=>"110110010",
  32978=>"010000000",
  32979=>"000000000",
  32980=>"011001000",
  32981=>"111110000",
  32982=>"111110100",
  32983=>"000000101",
  32984=>"000000000",
  32985=>"001000100",
  32986=>"011001010",
  32987=>"111111000",
  32988=>"010101000",
  32989=>"000000000",
  32990=>"000000000",
  32991=>"111111000",
  32992=>"111000000",
  32993=>"000000000",
  32994=>"000001000",
  32995=>"011001001",
  32996=>"101101000",
  32997=>"000010000",
  32998=>"000010010",
  32999=>"000100010",
  33000=>"000111111",
  33001=>"110010001",
  33002=>"001011100",
  33003=>"011000101",
  33004=>"000010010",
  33005=>"000000000",
  33006=>"000000000",
  33007=>"000000000",
  33008=>"000000111",
  33009=>"111000000",
  33010=>"011001111",
  33011=>"011010010",
  33012=>"000100011",
  33013=>"111111111",
  33014=>"100000000",
  33015=>"000001000",
  33016=>"111000000",
  33017=>"001111111",
  33018=>"111100100",
  33019=>"000010001",
  33020=>"001000000",
  33021=>"000111111",
  33022=>"011111111",
  33023=>"100111111",
  33024=>"011011111",
  33025=>"011010100",
  33026=>"100000111",
  33027=>"000000111",
  33028=>"000100101",
  33029=>"111000000",
  33030=>"100100111",
  33031=>"000111110",
  33032=>"000000000",
  33033=>"001000000",
  33034=>"011010011",
  33035=>"000100000",
  33036=>"111111101",
  33037=>"000011111",
  33038=>"100100111",
  33039=>"101000000",
  33040=>"000000011",
  33041=>"000111111",
  33042=>"100000100",
  33043=>"110000000",
  33044=>"001000011",
  33045=>"000111000",
  33046=>"011001000",
  33047=>"010111111",
  33048=>"011010000",
  33049=>"011101001",
  33050=>"001011010",
  33051=>"001000000",
  33052=>"111000111",
  33053=>"101010000",
  33054=>"110010000",
  33055=>"100101100",
  33056=>"000111010",
  33057=>"001101000",
  33058=>"000000000",
  33059=>"000101011",
  33060=>"111111110",
  33061=>"110110001",
  33062=>"000011010",
  33063=>"101000010",
  33064=>"000010010",
  33065=>"010111000",
  33066=>"100000000",
  33067=>"111111000",
  33068=>"111111100",
  33069=>"111000000",
  33070=>"111011111",
  33071=>"001000010",
  33072=>"010011010",
  33073=>"000010011",
  33074=>"101111010",
  33075=>"111111000",
  33076=>"000010000",
  33077=>"000100000",
  33078=>"111110100",
  33079=>"000000110",
  33080=>"011010011",
  33081=>"000000000",
  33082=>"000000010",
  33083=>"101010011",
  33084=>"100100000",
  33085=>"010101000",
  33086=>"000101101",
  33087=>"000001011",
  33088=>"011110001",
  33089=>"111001000",
  33090=>"010011000",
  33091=>"001001011",
  33092=>"111111100",
  33093=>"000000000",
  33094=>"111010000",
  33095=>"100111111",
  33096=>"000001110",
  33097=>"000110011",
  33098=>"000101100",
  33099=>"001000001",
  33100=>"100000010",
  33101=>"100100110",
  33102=>"001001111",
  33103=>"111100110",
  33104=>"010000100",
  33105=>"010000000",
  33106=>"111001101",
  33107=>"011011011",
  33108=>"000011111",
  33109=>"011111001",
  33110=>"001111011",
  33111=>"000000000",
  33112=>"111000001",
  33113=>"010000001",
  33114=>"000000010",
  33115=>"011011001",
  33116=>"111111111",
  33117=>"000001000",
  33118=>"111101000",
  33119=>"100000011",
  33120=>"111111011",
  33121=>"001000111",
  33122=>"111101001",
  33123=>"110010000",
  33124=>"001101101",
  33125=>"000000000",
  33126=>"000010111",
  33127=>"000000000",
  33128=>"111111111",
  33129=>"010000010",
  33130=>"111000001",
  33131=>"110000101",
  33132=>"000111000",
  33133=>"100111111",
  33134=>"000000100",
  33135=>"000000000",
  33136=>"000100110",
  33137=>"111011000",
  33138=>"011011000",
  33139=>"011110100",
  33140=>"110100111",
  33141=>"001000000",
  33142=>"010000010",
  33143=>"111101000",
  33144=>"111111010",
  33145=>"110000111",
  33146=>"111101000",
  33147=>"001011111",
  33148=>"010001111",
  33149=>"010110010",
  33150=>"001111111",
  33151=>"000011111",
  33152=>"111011000",
  33153=>"010010010",
  33154=>"000000010",
  33155=>"101001000",
  33156=>"000000000",
  33157=>"100010111",
  33158=>"011001100",
  33159=>"011000110",
  33160=>"100001011",
  33161=>"000010111",
  33162=>"000011011",
  33163=>"000111110",
  33164=>"000000110",
  33165=>"000111111",
  33166=>"111101000",
  33167=>"111001001",
  33168=>"001001001",
  33169=>"101111010",
  33170=>"100111111",
  33171=>"000001010",
  33172=>"111111111",
  33173=>"100000000",
  33174=>"111100000",
  33175=>"000110110",
  33176=>"010111000",
  33177=>"101010101",
  33178=>"000010010",
  33179=>"111111010",
  33180=>"111100111",
  33181=>"111111000",
  33182=>"011111000",
  33183=>"001001010",
  33184=>"001000000",
  33185=>"111110000",
  33186=>"000011100",
  33187=>"000011011",
  33188=>"110111000",
  33189=>"110100000",
  33190=>"010000001",
  33191=>"110110100",
  33192=>"111000000",
  33193=>"001011010",
  33194=>"001101110",
  33195=>"000001101",
  33196=>"111101100",
  33197=>"101001011",
  33198=>"010101001",
  33199=>"011000000",
  33200=>"001101000",
  33201=>"110110110",
  33202=>"100000000",
  33203=>"000000000",
  33204=>"000111111",
  33205=>"010000100",
  33206=>"010011101",
  33207=>"111000100",
  33208=>"001000001",
  33209=>"010111011",
  33210=>"111010000",
  33211=>"000011011",
  33212=>"001001101",
  33213=>"111111111",
  33214=>"000110111",
  33215=>"111111000",
  33216=>"100100100",
  33217=>"010011111",
  33218=>"111111000",
  33219=>"110111110",
  33220=>"111011010",
  33221=>"100111001",
  33222=>"110011010",
  33223=>"001111111",
  33224=>"111000000",
  33225=>"000010000",
  33226=>"111010100",
  33227=>"010011101",
  33228=>"000010011",
  33229=>"110100010",
  33230=>"000101000",
  33231=>"010000111",
  33232=>"000000010",
  33233=>"110111010",
  33234=>"010010000",
  33235=>"111100100",
  33236=>"111111010",
  33237=>"011011011",
  33238=>"111111111",
  33239=>"000000011",
  33240=>"101001000",
  33241=>"000011111",
  33242=>"100100000",
  33243=>"000000010",
  33244=>"111100000",
  33245=>"000100110",
  33246=>"011011101",
  33247=>"001000000",
  33248=>"001001111",
  33249=>"111011000",
  33250=>"100000000",
  33251=>"011110110",
  33252=>"111011011",
  33253=>"111111000",
  33254=>"000000000",
  33255=>"000011000",
  33256=>"000111001",
  33257=>"110110101",
  33258=>"010011110",
  33259=>"101101001",
  33260=>"011001000",
  33261=>"111111110",
  33262=>"000000010",
  33263=>"000000000",
  33264=>"000111011",
  33265=>"011001100",
  33266=>"111011000",
  33267=>"100111111",
  33268=>"010111011",
  33269=>"111101111",
  33270=>"000000001",
  33271=>"100000000",
  33272=>"001001101",
  33273=>"011100000",
  33274=>"010111101",
  33275=>"111110111",
  33276=>"111000000",
  33277=>"000110111",
  33278=>"001101100",
  33279=>"010000000",
  33280=>"111000000",
  33281=>"000000100",
  33282=>"000100111",
  33283=>"000000000",
  33284=>"100110101",
  33285=>"000000111",
  33286=>"000010111",
  33287=>"100110111",
  33288=>"001001001",
  33289=>"111000000",
  33290=>"100110000",
  33291=>"000000000",
  33292=>"111001000",
  33293=>"000000000",
  33294=>"110011000",
  33295=>"001000000",
  33296=>"111010110",
  33297=>"000010110",
  33298=>"100010111",
  33299=>"000111111",
  33300=>"000010011",
  33301=>"000100111",
  33302=>"111001110",
  33303=>"010010000",
  33304=>"101000000",
  33305=>"011010011",
  33306=>"100100000",
  33307=>"000110111",
  33308=>"110000111",
  33309=>"110110110",
  33310=>"111010110",
  33311=>"000100100",
  33312=>"000000010",
  33313=>"000000000",
  33314=>"000000111",
  33315=>"111101111",
  33316=>"011000000",
  33317=>"011000000",
  33318=>"101111100",
  33319=>"111111111",
  33320=>"111111010",
  33321=>"100100000",
  33322=>"101111001",
  33323=>"110111111",
  33324=>"010011001",
  33325=>"110101111",
  33326=>"111111111",
  33327=>"000011001",
  33328=>"000000000",
  33329=>"110010110",
  33330=>"000001111",
  33331=>"011000000",
  33332=>"000111111",
  33333=>"000101000",
  33334=>"011011011",
  33335=>"000000111",
  33336=>"000000000",
  33337=>"000001011",
  33338=>"000011011",
  33339=>"011000000",
  33340=>"111100100",
  33341=>"010000001",
  33342=>"111100000",
  33343=>"000011001",
  33344=>"111000111",
  33345=>"010010011",
  33346=>"000111111",
  33347=>"000000000",
  33348=>"000011010",
  33349=>"111100000",
  33350=>"010000011",
  33351=>"110001101",
  33352=>"110101110",
  33353=>"111111100",
  33354=>"100110001",
  33355=>"101110010",
  33356=>"111000000",
  33357=>"110000011",
  33358=>"011000001",
  33359=>"010100111",
  33360=>"111001111",
  33361=>"111001101",
  33362=>"000010011",
  33363=>"011001000",
  33364=>"101000000",
  33365=>"111011000",
  33366=>"100110011",
  33367=>"000001111",
  33368=>"111011010",
  33369=>"111100000",
  33370=>"001010000",
  33371=>"000000100",
  33372=>"111011000",
  33373=>"011110000",
  33374=>"011111111",
  33375=>"001100101",
  33376=>"001001000",
  33377=>"011110111",
  33378=>"101000000",
  33379=>"100000100",
  33380=>"011111000",
  33381=>"000101001",
  33382=>"000110010",
  33383=>"000110100",
  33384=>"111010000",
  33385=>"000100110",
  33386=>"111111010",
  33387=>"000010111",
  33388=>"000111000",
  33389=>"000011111",
  33390=>"000000111",
  33391=>"000000000",
  33392=>"111100000",
  33393=>"000000100",
  33394=>"110110110",
  33395=>"001000110",
  33396=>"011111111",
  33397=>"100000000",
  33398=>"000010000",
  33399=>"100000101",
  33400=>"000000010",
  33401=>"111111111",
  33402=>"000111101",
  33403=>"011010000",
  33404=>"001010001",
  33405=>"111110000",
  33406=>"100111111",
  33407=>"000000010",
  33408=>"110110000",
  33409=>"000000000",
  33410=>"100100100",
  33411=>"000110111",
  33412=>"011001000",
  33413=>"000100110",
  33414=>"110000001",
  33415=>"000100100",
  33416=>"010010010",
  33417=>"000011011",
  33418=>"110011010",
  33419=>"000100111",
  33420=>"000101101",
  33421=>"000000000",
  33422=>"111000000",
  33423=>"010001001",
  33424=>"110011111",
  33425=>"111010110",
  33426=>"100000010",
  33427=>"111111100",
  33428=>"010111011",
  33429=>"111000000",
  33430=>"111011000",
  33431=>"111000000",
  33432=>"101111000",
  33433=>"101000111",
  33434=>"000000000",
  33435=>"011001001",
  33436=>"111101100",
  33437=>"111011000",
  33438=>"000000000",
  33439=>"110111010",
  33440=>"011010010",
  33441=>"110100010",
  33442=>"000111111",
  33443=>"101010111",
  33444=>"111011111",
  33445=>"110011011",
  33446=>"110000101",
  33447=>"000111111",
  33448=>"010110111",
  33449=>"000100000",
  33450=>"111000000",
  33451=>"000010100",
  33452=>"000000011",
  33453=>"111101001",
  33454=>"111010001",
  33455=>"000000010",
  33456=>"111000000",
  33457=>"010110111",
  33458=>"111000000",
  33459=>"100101001",
  33460=>"111100100",
  33461=>"000100000",
  33462=>"001000000",
  33463=>"000000000",
  33464=>"011001011",
  33465=>"100001010",
  33466=>"111100000",
  33467=>"000101000",
  33468=>"010010111",
  33469=>"111011111",
  33470=>"110100100",
  33471=>"000100011",
  33472=>"000111111",
  33473=>"010001101",
  33474=>"101101101",
  33475=>"110011111",
  33476=>"000100100",
  33477=>"011011100",
  33478=>"000100000",
  33479=>"111111111",
  33480=>"110001111",
  33481=>"000000000",
  33482=>"000010111",
  33483=>"111000000",
  33484=>"000100010",
  33485=>"010011001",
  33486=>"110110000",
  33487=>"111000000",
  33488=>"000111111",
  33489=>"111110001",
  33490=>"000100000",
  33491=>"011111101",
  33492=>"000000110",
  33493=>"001001001",
  33494=>"111101111",
  33495=>"000100001",
  33496=>"100111000",
  33497=>"000011000",
  33498=>"010010001",
  33499=>"111000000",
  33500=>"111100001",
  33501=>"011000101",
  33502=>"001001001",
  33503=>"000000000",
  33504=>"000100111",
  33505=>"000110111",
  33506=>"010000000",
  33507=>"001011111",
  33508=>"100000000",
  33509=>"000000001",
  33510=>"000011111",
  33511=>"111101000",
  33512=>"111110100",
  33513=>"000110010",
  33514=>"001011110",
  33515=>"000000111",
  33516=>"000101111",
  33517=>"000000000",
  33518=>"000000101",
  33519=>"111001000",
  33520=>"101110000",
  33521=>"111010100",
  33522=>"110000100",
  33523=>"111001000",
  33524=>"011100100",
  33525=>"000000111",
  33526=>"111101101",
  33527=>"011111000",
  33528=>"100111110",
  33529=>"010111011",
  33530=>"111000111",
  33531=>"000001001",
  33532=>"111000000",
  33533=>"010000000",
  33534=>"011010010",
  33535=>"011111111",
  33536=>"100001010",
  33537=>"110011011",
  33538=>"111001001",
  33539=>"000000110",
  33540=>"110000000",
  33541=>"010110000",
  33542=>"100110110",
  33543=>"000001111",
  33544=>"001111011",
  33545=>"011001001",
  33546=>"000100000",
  33547=>"110100100",
  33548=>"000100110",
  33549=>"011001000",
  33550=>"101001000",
  33551=>"111100100",
  33552=>"001001001",
  33553=>"000000111",
  33554=>"110011000",
  33555=>"110110010",
  33556=>"110001101",
  33557=>"001100110",
  33558=>"011000011",
  33559=>"110011001",
  33560=>"011001001",
  33561=>"001000011",
  33562=>"000010010",
  33563=>"000011111",
  33564=>"000010010",
  33565=>"010111110",
  33566=>"101111000",
  33567=>"001110110",
  33568=>"001001101",
  33569=>"011111010",
  33570=>"111101110",
  33571=>"000110110",
  33572=>"100100000",
  33573=>"001001011",
  33574=>"001110110",
  33575=>"000000011",
  33576=>"001111110",
  33577=>"000100110",
  33578=>"001110011",
  33579=>"001001001",
  33580=>"000101110",
  33581=>"100100111",
  33582=>"010111001",
  33583=>"000001111",
  33584=>"100110110",
  33585=>"001111111",
  33586=>"011011010",
  33587=>"111001000",
  33588=>"101001110",
  33589=>"110110110",
  33590=>"101001001",
  33591=>"110001111",
  33592=>"111001100",
  33593=>"111001011",
  33594=>"000111100",
  33595=>"000011011",
  33596=>"001110101",
  33597=>"111111000",
  33598=>"000000001",
  33599=>"000110110",
  33600=>"001001001",
  33601=>"001001011",
  33602=>"111001000",
  33603=>"001111111",
  33604=>"011001010",
  33605=>"000110011",
  33606=>"110000110",
  33607=>"110110000",
  33608=>"111100100",
  33609=>"110011100",
  33610=>"000000111",
  33611=>"001001000",
  33612=>"111001111",
  33613=>"000101100",
  33614=>"000100100",
  33615=>"001101101",
  33616=>"011001001",
  33617=>"010101000",
  33618=>"110000110",
  33619=>"110011011",
  33620=>"111001001",
  33621=>"110000011",
  33622=>"111110110",
  33623=>"111001001",
  33624=>"010110100",
  33625=>"110111111",
  33626=>"000001001",
  33627=>"000100000",
  33628=>"000001000",
  33629=>"000010011",
  33630=>"111001011",
  33631=>"000101000",
  33632=>"000110110",
  33633=>"010110111",
  33634=>"001001001",
  33635=>"111111001",
  33636=>"010001110",
  33637=>"000000100",
  33638=>"110100000",
  33639=>"011000011",
  33640=>"000100110",
  33641=>"110110001",
  33642=>"000101101",
  33643=>"010001110",
  33644=>"110011111",
  33645=>"000000001",
  33646=>"001001100",
  33647=>"000111111",
  33648=>"111111011",
  33649=>"000000000",
  33650=>"000001001",
  33651=>"000110000",
  33652=>"001001011",
  33653=>"010001001",
  33654=>"101000000",
  33655=>"001001001",
  33656=>"000011001",
  33657=>"111110010",
  33658=>"111001000",
  33659=>"000111100",
  33660=>"111000011",
  33661=>"101000000",
  33662=>"001001001",
  33663=>"001100100",
  33664=>"110111001",
  33665=>"000110000",
  33666=>"000110100",
  33667=>"000110001",
  33668=>"000110010",
  33669=>"110001000",
  33670=>"000001111",
  33671=>"111001101",
  33672=>"110110110",
  33673=>"001000000",
  33674=>"000001001",
  33675=>"110100001",
  33676=>"011001001",
  33677=>"011001001",
  33678=>"100000000",
  33679=>"001001111",
  33680=>"101101110",
  33681=>"001000111",
  33682=>"001001000",
  33683=>"111110011",
  33684=>"101000000",
  33685=>"011001100",
  33686=>"001110010",
  33687=>"000110111",
  33688=>"000110000",
  33689=>"001111000",
  33690=>"100110100",
  33691=>"111011001",
  33692=>"111111000",
  33693=>"111001001",
  33694=>"111110111",
  33695=>"001110000",
  33696=>"111111101",
  33697=>"011001001",
  33698=>"011001001",
  33699=>"110111011",
  33700=>"110110000",
  33701=>"000000111",
  33702=>"100100000",
  33703=>"000000100",
  33704=>"110100110",
  33705=>"110100110",
  33706=>"000100100",
  33707=>"001111001",
  33708=>"110110010",
  33709=>"011001000",
  33710=>"010000011",
  33711=>"101001001",
  33712=>"000010100",
  33713=>"000010111",
  33714=>"000011001",
  33715=>"101011001",
  33716=>"010110100",
  33717=>"111011111",
  33718=>"110110101",
  33719=>"001001011",
  33720=>"000110100",
  33721=>"110010011",
  33722=>"010011000",
  33723=>"110110001",
  33724=>"110110110",
  33725=>"111111110",
  33726=>"000111101",
  33727=>"000111001",
  33728=>"111001001",
  33729=>"101001011",
  33730=>"111110110",
  33731=>"001100100",
  33732=>"000100010",
  33733=>"000110110",
  33734=>"110001001",
  33735=>"000110001",
  33736=>"000110001",
  33737=>"000000110",
  33738=>"110011011",
  33739=>"000000110",
  33740=>"011001001",
  33741=>"111001001",
  33742=>"011001001",
  33743=>"010111111",
  33744=>"100100000",
  33745=>"000100100",
  33746=>"111100011",
  33747=>"000100010",
  33748=>"001001001",
  33749=>"011001100",
  33750=>"011000101",
  33751=>"000111110",
  33752=>"100100110",
  33753=>"110110110",
  33754=>"001101001",
  33755=>"110001001",
  33756=>"001001000",
  33757=>"001111010",
  33758=>"110111110",
  33759=>"010101001",
  33760=>"001001111",
  33761=>"111011001",
  33762=>"101100000",
  33763=>"011111111",
  33764=>"101001101",
  33765=>"011001001",
  33766=>"000110110",
  33767=>"000110011",
  33768=>"010010000",
  33769=>"100100111",
  33770=>"001000000",
  33771=>"100001011",
  33772=>"001010100",
  33773=>"000110110",
  33774=>"010001111",
  33775=>"000110110",
  33776=>"110110110",
  33777=>"110000101",
  33778=>"100101000",
  33779=>"100100000",
  33780=>"000110101",
  33781=>"111001001",
  33782=>"000000010",
  33783=>"110000000",
  33784=>"111001011",
  33785=>"110000010",
  33786=>"110001001",
  33787=>"000111110",
  33788=>"000110110",
  33789=>"011001001",
  33790=>"110101001",
  33791=>"111001001",
  33792=>"000001100",
  33793=>"010000000",
  33794=>"001001111",
  33795=>"000000110",
  33796=>"001001101",
  33797=>"010001011",
  33798=>"110101111",
  33799=>"000000001",
  33800=>"000010100",
  33801=>"001100111",
  33802=>"010101001",
  33803=>"110100010",
  33804=>"000000001",
  33805=>"001001001",
  33806=>"011011011",
  33807=>"111001000",
  33808=>"010110100",
  33809=>"000000100",
  33810=>"001111110",
  33811=>"000110110",
  33812=>"111111111",
  33813=>"010010110",
  33814=>"000000001",
  33815=>"000110110",
  33816=>"110111111",
  33817=>"111111011",
  33818=>"000000000",
  33819=>"000000001",
  33820=>"110110000",
  33821=>"000101110",
  33822=>"000000011",
  33823=>"001001101",
  33824=>"001101111",
  33825=>"000001010",
  33826=>"001000000",
  33827=>"001000100",
  33828=>"101100100",
  33829=>"111101010",
  33830=>"000101111",
  33831=>"111000101",
  33832=>"001001111",
  33833=>"011100011",
  33834=>"000000000",
  33835=>"001000100",
  33836=>"010001000",
  33837=>"111111111",
  33838=>"010100011",
  33839=>"110001010",
  33840=>"000000000",
  33841=>"101111011",
  33842=>"000001111",
  33843=>"001001011",
  33844=>"110110100",
  33845=>"111101110",
  33846=>"111011111",
  33847=>"110111000",
  33848=>"011000110",
  33849=>"001001000",
  33850=>"111111100",
  33851=>"000000100",
  33852=>"010000000",
  33853=>"111011010",
  33854=>"000000011",
  33855=>"100101111",
  33856=>"110111111",
  33857=>"110110000",
  33858=>"001000000",
  33859=>"011000100",
  33860=>"000001000",
  33861=>"001101111",
  33862=>"110110000",
  33863=>"001111111",
  33864=>"101011010",
  33865=>"111101001",
  33866=>"000001011",
  33867=>"110110000",
  33868=>"111001111",
  33869=>"011111011",
  33870=>"100111101",
  33871=>"001010110",
  33872=>"000010010",
  33873=>"101000111",
  33874=>"011111111",
  33875=>"011011010",
  33876=>"010110000",
  33877=>"000001010",
  33878=>"010011010",
  33879=>"000010111",
  33880=>"011011000",
  33881=>"000001001",
  33882=>"000101000",
  33883=>"011111000",
  33884=>"000000000",
  33885=>"001000001",
  33886=>"110010110",
  33887=>"100001011",
  33888=>"101101111",
  33889=>"000000000",
  33890=>"001000101",
  33891=>"000001110",
  33892=>"000000000",
  33893=>"111111101",
  33894=>"100101011",
  33895=>"001101111",
  33896=>"111101111",
  33897=>"000111111",
  33898=>"001111111",
  33899=>"000000100",
  33900=>"000001000",
  33901=>"110110111",
  33902=>"000100110",
  33903=>"010000000",
  33904=>"001011001",
  33905=>"000000000",
  33906=>"001000100",
  33907=>"111111000",
  33908=>"000000000",
  33909=>"101001000",
  33910=>"111010010",
  33911=>"111000001",
  33912=>"001000110",
  33913=>"011111111",
  33914=>"111010000",
  33915=>"110001011",
  33916=>"110010010",
  33917=>"100000010",
  33918=>"111110110",
  33919=>"001001001",
  33920=>"111100000",
  33921=>"010000000",
  33922=>"111000100",
  33923=>"110010111",
  33924=>"001001100",
  33925=>"111111101",
  33926=>"011011001",
  33927=>"011001000",
  33928=>"000000000",
  33929=>"000000001",
  33930=>"010111101",
  33931=>"000000110",
  33932=>"000000100",
  33933=>"110110110",
  33934=>"111011000",
  33935=>"111000000",
  33936=>"111010110",
  33937=>"011111100",
  33938=>"000000010",
  33939=>"000110111",
  33940=>"110111101",
  33941=>"001000110",
  33942=>"111111000",
  33943=>"100100010",
  33944=>"111101111",
  33945=>"010001111",
  33946=>"111010111",
  33947=>"111111111",
  33948=>"011111111",
  33949=>"010010000",
  33950=>"110110000",
  33951=>"000100111",
  33952=>"101100110",
  33953=>"111001111",
  33954=>"000000010",
  33955=>"101111001",
  33956=>"010110110",
  33957=>"110111000",
  33958=>"000000111",
  33959=>"111101000",
  33960=>"010110010",
  33961=>"101010110",
  33962=>"111111010",
  33963=>"001000110",
  33964=>"111111111",
  33965=>"000000010",
  33966=>"110000000",
  33967=>"111111110",
  33968=>"110000011",
  33969=>"010111001",
  33970=>"111001001",
  33971=>"001000100",
  33972=>"000001010",
  33973=>"000011000",
  33974=>"111101000",
  33975=>"100000000",
  33976=>"011010010",
  33977=>"110110010",
  33978=>"111101110",
  33979=>"101111111",
  33980=>"000100101",
  33981=>"111111111",
  33982=>"010011111",
  33983=>"000000000",
  33984=>"110110110",
  33985=>"010110000",
  33986=>"110000000",
  33987=>"011110100",
  33988=>"110001001",
  33989=>"001101001",
  33990=>"000111110",
  33991=>"000000001",
  33992=>"111100110",
  33993=>"001001001",
  33994=>"001000000",
  33995=>"111111000",
  33996=>"000101000",
  33997=>"011101100",
  33998=>"000010000",
  33999=>"101101111",
  34000=>"010110010",
  34001=>"011011111",
  34002=>"110000000",
  34003=>"111110000",
  34004=>"010000101",
  34005=>"000000010",
  34006=>"001001111",
  34007=>"110011010",
  34008=>"000100110",
  34009=>"000110110",
  34010=>"011001001",
  34011=>"000110000",
  34012=>"000000001",
  34013=>"101101010",
  34014=>"111111000",
  34015=>"001101100",
  34016=>"001001101",
  34017=>"101001001",
  34018=>"010000000",
  34019=>"110110001",
  34020=>"001001111",
  34021=>"000000001",
  34022=>"110110111",
  34023=>"010110111",
  34024=>"001001111",
  34025=>"010110110",
  34026=>"010100100",
  34027=>"011110010",
  34028=>"000001101",
  34029=>"110100000",
  34030=>"000000000",
  34031=>"000000001",
  34032=>"000000000",
  34033=>"000011100",
  34034=>"001000011",
  34035=>"000001111",
  34036=>"000111011",
  34037=>"011000000",
  34038=>"110100010",
  34039=>"010000010",
  34040=>"110010000",
  34041=>"000001111",
  34042=>"010110000",
  34043=>"010111110",
  34044=>"111111110",
  34045=>"010111111",
  34046=>"111111011",
  34047=>"111111001",
  34048=>"000000000",
  34049=>"000000000",
  34050=>"111000111",
  34051=>"010000111",
  34052=>"000000000",
  34053=>"111111011",
  34054=>"000000100",
  34055=>"000000000",
  34056=>"000010011",
  34057=>"000000111",
  34058=>"000000100",
  34059=>"011100100",
  34060=>"011011111",
  34061=>"101000101",
  34062=>"110000100",
  34063=>"110000000",
  34064=>"111011011",
  34065=>"101111000",
  34066=>"100000110",
  34067=>"011111000",
  34068=>"111011001",
  34069=>"000001001",
  34070=>"000000000",
  34071=>"111111100",
  34072=>"000010011",
  34073=>"101000000",
  34074=>"000000010",
  34075=>"000000111",
  34076=>"011111011",
  34077=>"000101000",
  34078=>"100111010",
  34079=>"101100100",
  34080=>"111000101",
  34081=>"000000000",
  34082=>"000100001",
  34083=>"111100111",
  34084=>"100110110",
  34085=>"100000010",
  34086=>"111110000",
  34087=>"000101011",
  34088=>"111111111",
  34089=>"001111111",
  34090=>"000000000",
  34091=>"001111111",
  34092=>"000011011",
  34093=>"111010100",
  34094=>"100111000",
  34095=>"000000000",
  34096=>"101111010",
  34097=>"011000100",
  34098=>"000000000",
  34099=>"101111000",
  34100=>"000000111",
  34101=>"100110000",
  34102=>"010000011",
  34103=>"000100111",
  34104=>"100111111",
  34105=>"000000000",
  34106=>"111000000",
  34107=>"100111111",
  34108=>"100001101",
  34109=>"111101101",
  34110=>"000110010",
  34111=>"000010011",
  34112=>"001111011",
  34113=>"000001010",
  34114=>"001011000",
  34115=>"000100110",
  34116=>"101000000",
  34117=>"000111111",
  34118=>"000000000",
  34119=>"100100000",
  34120=>"010011111",
  34121=>"100000011",
  34122=>"110010110",
  34123=>"010111011",
  34124=>"011111111",
  34125=>"000001011",
  34126=>"100000000",
  34127=>"111111100",
  34128=>"000000111",
  34129=>"101100101",
  34130=>"000111000",
  34131=>"100010110",
  34132=>"110000100",
  34133=>"001001111",
  34134=>"011110100",
  34135=>"101101101",
  34136=>"001001000",
  34137=>"000011001",
  34138=>"011011011",
  34139=>"000111011",
  34140=>"000111010",
  34141=>"111000100",
  34142=>"101000101",
  34143=>"100000011",
  34144=>"111011111",
  34145=>"100100000",
  34146=>"010010111",
  34147=>"111110110",
  34148=>"010111101",
  34149=>"010010010",
  34150=>"100000000",
  34151=>"100100111",
  34152=>"001000110",
  34153=>"000000110",
  34154=>"000111111",
  34155=>"010000010",
  34156=>"111111000",
  34157=>"000111000",
  34158=>"111111010",
  34159=>"000000000",
  34160=>"010011011",
  34161=>"111111011",
  34162=>"001000110",
  34163=>"000100000",
  34164=>"000111111",
  34165=>"110100111",
  34166=>"000000000",
  34167=>"111111111",
  34168=>"101001000",
  34169=>"000111111",
  34170=>"111111000",
  34171=>"101000100",
  34172=>"011001100",
  34173=>"000001001",
  34174=>"101100111",
  34175=>"011100111",
  34176=>"100011111",
  34177=>"111111000",
  34178=>"000011010",
  34179=>"100100111",
  34180=>"000010000",
  34181=>"111111111",
  34182=>"001010110",
  34183=>"110100001",
  34184=>"111010010",
  34185=>"000000000",
  34186=>"111111101",
  34187=>"001001111",
  34188=>"111111011",
  34189=>"000111010",
  34190=>"000110111",
  34191=>"011000000",
  34192=>"001000011",
  34193=>"100111111",
  34194=>"101000000",
  34195=>"000000000",
  34196=>"010000010",
  34197=>"001111011",
  34198=>"111000001",
  34199=>"110111111",
  34200=>"000111011",
  34201=>"101101101",
  34202=>"111000100",
  34203=>"100011111",
  34204=>"000011011",
  34205=>"100111000",
  34206=>"010111111",
  34207=>"111111111",
  34208=>"101111111",
  34209=>"111111000",
  34210=>"010000111",
  34211=>"111000000",
  34212=>"000111110",
  34213=>"000110110",
  34214=>"000111011",
  34215=>"010111011",
  34216=>"000111111",
  34217=>"111011111",
  34218=>"101000001",
  34219=>"010111111",
  34220=>"101101001",
  34221=>"010110011",
  34222=>"100101101",
  34223=>"111111000",
  34224=>"100111101",
  34225=>"110011100",
  34226=>"000010000",
  34227=>"011011000",
  34228=>"100010110",
  34229=>"000010000",
  34230=>"000000100",
  34231=>"010000011",
  34232=>"100100101",
  34233=>"010000000",
  34234=>"100001000",
  34235=>"001111111",
  34236=>"100111000",
  34237=>"111100101",
  34238=>"000010000",
  34239=>"101000111",
  34240=>"111111011",
  34241=>"010110010",
  34242=>"111001000",
  34243=>"111110111",
  34244=>"001100000",
  34245=>"110111011",
  34246=>"100111000",
  34247=>"001000001",
  34248=>"001000000",
  34249=>"011011111",
  34250=>"000000000",
  34251=>"111000000",
  34252=>"111111111",
  34253=>"111100101",
  34254=>"010000000",
  34255=>"001111110",
  34256=>"110111011",
  34257=>"001011011",
  34258=>"111111000",
  34259=>"111110010",
  34260=>"000000000",
  34261=>"001000001",
  34262=>"011010010",
  34263=>"011011011",
  34264=>"001000100",
  34265=>"100011111",
  34266=>"111010010",
  34267=>"010111010",
  34268=>"000000110",
  34269=>"100111001",
  34270=>"000010000",
  34271=>"100000110",
  34272=>"000101010",
  34273=>"111111110",
  34274=>"100000100",
  34275=>"100110111",
  34276=>"010000001",
  34277=>"000101100",
  34278=>"010011010",
  34279=>"000001101",
  34280=>"011010000",
  34281=>"110000111",
  34282=>"000000000",
  34283=>"000000001",
  34284=>"111111111",
  34285=>"000100000",
  34286=>"100111111",
  34287=>"111000100",
  34288=>"000000000",
  34289=>"001110011",
  34290=>"000101111",
  34291=>"000011011",
  34292=>"000100000",
  34293=>"010010010",
  34294=>"010011010",
  34295=>"011000000",
  34296=>"101101101",
  34297=>"100000100",
  34298=>"111111011",
  34299=>"000100101",
  34300=>"101111101",
  34301=>"000011010",
  34302=>"000010110",
  34303=>"111011111",
  34304=>"111001100",
  34305=>"000000000",
  34306=>"111101100",
  34307=>"101010100",
  34308=>"000000010",
  34309=>"001011100",
  34310=>"000001001",
  34311=>"000000001",
  34312=>"000000000",
  34313=>"010100000",
  34314=>"000100110",
  34315=>"000011110",
  34316=>"110010000",
  34317=>"100001001",
  34318=>"100010000",
  34319=>"101010011",
  34320=>"101000000",
  34321=>"111000100",
  34322=>"001110100",
  34323=>"011001111",
  34324=>"111100110",
  34325=>"111000110",
  34326=>"001110111",
  34327=>"111101111",
  34328=>"111010000",
  34329=>"100000011",
  34330=>"000110011",
  34331=>"000100110",
  34332=>"000000011",
  34333=>"000000100",
  34334=>"010111100",
  34335=>"111100011",
  34336=>"001000111",
  34337=>"001001001",
  34338=>"110000011",
  34339=>"000000000",
  34340=>"000000101",
  34341=>"100001001",
  34342=>"111100100",
  34343=>"000000011",
  34344=>"111110100",
  34345=>"111011110",
  34346=>"000011111",
  34347=>"111111100",
  34348=>"000010011",
  34349=>"000010000",
  34350=>"000000110",
  34351=>"000001011",
  34352=>"110100100",
  34353=>"101011011",
  34354=>"111000100",
  34355=>"101111111",
  34356=>"001011111",
  34357=>"110111111",
  34358=>"000110000",
  34359=>"100110100",
  34360=>"000011011",
  34361=>"111100000",
  34362=>"111100000",
  34363=>"001110110",
  34364=>"100100001",
  34365=>"010011111",
  34366=>"111100100",
  34367=>"000001000",
  34368=>"100100100",
  34369=>"010111111",
  34370=>"000011011",
  34371=>"010110100",
  34372=>"111000000",
  34373=>"000001001",
  34374=>"001100100",
  34375=>"111001001",
  34376=>"000110111",
  34377=>"000011111",
  34378=>"001111110",
  34379=>"010110111",
  34380=>"010100110",
  34381=>"110111010",
  34382=>"110100101",
  34383=>"100001111",
  34384=>"111110001",
  34385=>"011100111",
  34386=>"111011110",
  34387=>"001011001",
  34388=>"000000000",
  34389=>"001000111",
  34390=>"100000010",
  34391=>"010011000",
  34392=>"100100111",
  34393=>"010001011",
  34394=>"100111101",
  34395=>"010000101",
  34396=>"000000000",
  34397=>"010100100",
  34398=>"111010110",
  34399=>"111100100",
  34400=>"110100000",
  34401=>"100110111",
  34402=>"111110100",
  34403=>"000000110",
  34404=>"100010001",
  34405=>"100100110",
  34406=>"000000001",
  34407=>"111011000",
  34408=>"011110100",
  34409=>"000000111",
  34410=>"011010000",
  34411=>"111110111",
  34412=>"111110100",
  34413=>"010111111",
  34414=>"010001001",
  34415=>"011011111",
  34416=>"000011111",
  34417=>"000100000",
  34418=>"111000100",
  34419=>"000101001",
  34420=>"010100111",
  34421=>"101100100",
  34422=>"000010011",
  34423=>"100111100",
  34424=>"101000010",
  34425=>"010001111",
  34426=>"011111111",
  34427=>"000000101",
  34428=>"110011011",
  34429=>"100101010",
  34430=>"001100100",
  34431=>"011010000",
  34432=>"110011000",
  34433=>"001011100",
  34434=>"011001001",
  34435=>"000001000",
  34436=>"000100111",
  34437=>"011110000",
  34438=>"010010011",
  34439=>"000000010",
  34440=>"110101110",
  34441=>"111000000",
  34442=>"101111000",
  34443=>"000001111",
  34444=>"111110100",
  34445=>"000000000",
  34446=>"100111001",
  34447=>"000100000",
  34448=>"110010011",
  34449=>"101111011",
  34450=>"100000011",
  34451=>"111111100",
  34452=>"000100011",
  34453=>"011100100",
  34454=>"110010111",
  34455=>"110111111",
  34456=>"001111111",
  34457=>"100110011",
  34458=>"000010011",
  34459=>"111100101",
  34460=>"000000000",
  34461=>"111110000",
  34462=>"000011000",
  34463=>"111110000",
  34464=>"000010001",
  34465=>"111111111",
  34466=>"100101011",
  34467=>"010010000",
  34468=>"000000011",
  34469=>"000100111",
  34470=>"100000000",
  34471=>"000001011",
  34472=>"111111100",
  34473=>"001011001",
  34474=>"110100100",
  34475=>"111011000",
  34476=>"100011111",
  34477=>"000011011",
  34478=>"111111110",
  34479=>"011101000",
  34480=>"001011000",
  34481=>"000100100",
  34482=>"001111110",
  34483=>"000001000",
  34484=>"100000011",
  34485=>"010111011",
  34486=>"000011011",
  34487=>"010011011",
  34488=>"000111001",
  34489=>"000000111",
  34490=>"000011011",
  34491=>"010011001",
  34492=>"000111011",
  34493=>"011110111",
  34494=>"000001010",
  34495=>"010000001",
  34496=>"111100100",
  34497=>"000001001",
  34498=>"000011011",
  34499=>"000011011",
  34500=>"000000011",
  34501=>"100100111",
  34502=>"111011011",
  34503=>"000001111",
  34504=>"000001010",
  34505=>"011111000",
  34506=>"100110011",
  34507=>"111100100",
  34508=>"110111110",
  34509=>"011110011",
  34510=>"001001001",
  34511=>"100001000",
  34512=>"010110000",
  34513=>"000010110",
  34514=>"110100000",
  34515=>"010110111",
  34516=>"111100100",
  34517=>"110100010",
  34518=>"001001100",
  34519=>"110011011",
  34520=>"000010011",
  34521=>"110000000",
  34522=>"100110111",
  34523=>"011100100",
  34524=>"110111010",
  34525=>"011000111",
  34526=>"000011011",
  34527=>"000000100",
  34528=>"111000001",
  34529=>"111110100",
  34530=>"011000100",
  34531=>"111011110",
  34532=>"010111010",
  34533=>"001000011",
  34534=>"000011011",
  34535=>"111111110",
  34536=>"000100110",
  34537=>"000100011",
  34538=>"000100000",
  34539=>"101011011",
  34540=>"110011011",
  34541=>"011111110",
  34542=>"010000000",
  34543=>"000001100",
  34544=>"110100100",
  34545=>"000010111",
  34546=>"011001100",
  34547=>"000010010",
  34548=>"001001110",
  34549=>"100100100",
  34550=>"011100000",
  34551=>"000000000",
  34552=>"000000111",
  34553=>"000001001",
  34554=>"011011111",
  34555=>"011000111",
  34556=>"111100100",
  34557=>"001000110",
  34558=>"000011111",
  34559=>"010111100",
  34560=>"111110110",
  34561=>"000000001",
  34562=>"111111110",
  34563=>"100111001",
  34564=>"111111100",
  34565=>"110010001",
  34566=>"000010110",
  34567=>"110111110",
  34568=>"111111000",
  34569=>"111001001",
  34570=>"001001011",
  34571=>"111111001",
  34572=>"111010000",
  34573=>"000101000",
  34574=>"111011000",
  34575=>"000000010",
  34576=>"000110010",
  34577=>"000000000",
  34578=>"000000001",
  34579=>"010000010",
  34580=>"000011010",
  34581=>"111111110",
  34582=>"000000110",
  34583=>"111110010",
  34584=>"010000011",
  34585=>"000100111",
  34586=>"001000000",
  34587=>"000000011",
  34588=>"101011111",
  34589=>"101000011",
  34590=>"111011101",
  34591=>"101000000",
  34592=>"000111111",
  34593=>"111011001",
  34594=>"111011000",
  34595=>"111000111",
  34596=>"011101100",
  34597=>"101011010",
  34598=>"000000101",
  34599=>"000000000",
  34600=>"000100110",
  34601=>"111111111",
  34602=>"111000000",
  34603=>"000110111",
  34604=>"011011000",
  34605=>"100111101",
  34606=>"000000000",
  34607=>"001101111",
  34608=>"011111111",
  34609=>"101101001",
  34610=>"000101000",
  34611=>"000111111",
  34612=>"010110000",
  34613=>"111111111",
  34614=>"000001010",
  34615=>"111001100",
  34616=>"110111111",
  34617=>"111001000",
  34618=>"101011000",
  34619=>"000111110",
  34620=>"011000011",
  34621=>"001011011",
  34622=>"000000000",
  34623=>"101000000",
  34624=>"110010110",
  34625=>"110011001",
  34626=>"010010101",
  34627=>"001000100",
  34628=>"010000000",
  34629=>"010010001",
  34630=>"011000000",
  34631=>"000001100",
  34632=>"111011111",
  34633=>"000011111",
  34634=>"110111101",
  34635=>"111111000",
  34636=>"111111111",
  34637=>"101001000",
  34638=>"111101010",
  34639=>"111110000",
  34640=>"001001001",
  34641=>"100111010",
  34642=>"111000000",
  34643=>"111100111",
  34644=>"000000001",
  34645=>"100101001",
  34646=>"000010011",
  34647=>"000001111",
  34648=>"111101001",
  34649=>"001001000",
  34650=>"111000001",
  34651=>"001010000",
  34652=>"100010110",
  34653=>"100000100",
  34654=>"011111110",
  34655=>"000011111",
  34656=>"010000000",
  34657=>"001000000",
  34658=>"100000000",
  34659=>"011000000",
  34660=>"111000000",
  34661=>"111001000",
  34662=>"001111111",
  34663=>"001111111",
  34664=>"110011111",
  34665=>"000000101",
  34666=>"001001011",
  34667=>"111111000",
  34668=>"000110100",
  34669=>"000011111",
  34670=>"000000101",
  34671=>"000000000",
  34672=>"011111110",
  34673=>"001111111",
  34674=>"000100111",
  34675=>"111010011",
  34676=>"101000110",
  34677=>"001101001",
  34678=>"011111100",
  34679=>"111111100",
  34680=>"000000111",
  34681=>"000000111",
  34682=>"001101010",
  34683=>"101111000",
  34684=>"101100010",
  34685=>"110100011",
  34686=>"000111111",
  34687=>"110000000",
  34688=>"000010001",
  34689=>"111111000",
  34690=>"000010110",
  34691=>"111111000",
  34692=>"111000011",
  34693=>"101111111",
  34694=>"010100001",
  34695=>"011011010",
  34696=>"011111011",
  34697=>"000001101",
  34698=>"000111111",
  34699=>"010010011",
  34700=>"000101111",
  34701=>"000011111",
  34702=>"001000100",
  34703=>"001000000",
  34704=>"000001011",
  34705=>"101000000",
  34706=>"000111011",
  34707=>"111101000",
  34708=>"111101100",
  34709=>"000101001",
  34710=>"110000000",
  34711=>"100111100",
  34712=>"111101100",
  34713=>"000000111",
  34714=>"000100111",
  34715=>"100000000",
  34716=>"111111000",
  34717=>"101000000",
  34718=>"000001001",
  34719=>"110110000",
  34720=>"000000010",
  34721=>"000111011",
  34722=>"000111000",
  34723=>"110000101",
  34724=>"110111101",
  34725=>"001000000",
  34726=>"111110000",
  34727=>"000010110",
  34728=>"000111111",
  34729=>"000010101",
  34730=>"011111101",
  34731=>"010000000",
  34732=>"001111000",
  34733=>"110100000",
  34734=>"101011011",
  34735=>"011110000",
  34736=>"111100110",
  34737=>"111101010",
  34738=>"100011000",
  34739=>"001001100",
  34740=>"100111001",
  34741=>"111110110",
  34742=>"111111000",
  34743=>"111111111",
  34744=>"100000110",
  34745=>"001000001",
  34746=>"111011011",
  34747=>"000001110",
  34748=>"111101101",
  34749=>"111000111",
  34750=>"111100000",
  34751=>"001111111",
  34752=>"111010000",
  34753=>"011000000",
  34754=>"011011101",
  34755=>"111001100",
  34756=>"100000111",
  34757=>"001100111",
  34758=>"110100111",
  34759=>"111011000",
  34760=>"011111100",
  34761=>"111001001",
  34762=>"110000001",
  34763=>"111000001",
  34764=>"000000000",
  34765=>"010001010",
  34766=>"001000000",
  34767=>"100000100",
  34768=>"010000001",
  34769=>"001001000",
  34770=>"111000001",
  34771=>"100111011",
  34772=>"111000000",
  34773=>"001000010",
  34774=>"110000000",
  34775=>"000000100",
  34776=>"110111111",
  34777=>"100000111",
  34778=>"001000001",
  34779=>"001100111",
  34780=>"000111110",
  34781=>"111111101",
  34782=>"111111000",
  34783=>"111110100",
  34784=>"111000000",
  34785=>"111011000",
  34786=>"111011000",
  34787=>"110000000",
  34788=>"101000010",
  34789=>"111111000",
  34790=>"100110000",
  34791=>"110110010",
  34792=>"000000000",
  34793=>"000110111",
  34794=>"100000010",
  34795=>"011000000",
  34796=>"110111000",
  34797=>"000000000",
  34798=>"010010000",
  34799=>"111000000",
  34800=>"000000111",
  34801=>"001001010",
  34802=>"111001001",
  34803=>"011000000",
  34804=>"111010111",
  34805=>"001000101",
  34806=>"111000000",
  34807=>"001000111",
  34808=>"010111000",
  34809=>"001111110",
  34810=>"000000000",
  34811=>"001000101",
  34812=>"111010111",
  34813=>"001111111",
  34814=>"111000000",
  34815=>"011000000",
  34816=>"001100100",
  34817=>"011100000",
  34818=>"110100100",
  34819=>"111111111",
  34820=>"011000000",
  34821=>"001111111",
  34822=>"000111000",
  34823=>"110111111",
  34824=>"000000000",
  34825=>"000001010",
  34826=>"000000111",
  34827=>"101000000",
  34828=>"111010000",
  34829=>"000000000",
  34830=>"101000000",
  34831=>"000000110",
  34832=>"000000000",
  34833=>"011111000",
  34834=>"111000000",
  34835=>"111111000",
  34836=>"001000000",
  34837=>"111000010",
  34838=>"010000111",
  34839=>"111111001",
  34840=>"001010000",
  34841=>"000000000",
  34842=>"011000100",
  34843=>"101100110",
  34844=>"100000001",
  34845=>"000000000",
  34846=>"001100111",
  34847=>"000111110",
  34848=>"111111111",
  34849=>"010000100",
  34850=>"001101000",
  34851=>"011111111",
  34852=>"110111111",
  34853=>"000101001",
  34854=>"010111001",
  34855=>"110110000",
  34856=>"000001110",
  34857=>"111000000",
  34858=>"100000000",
  34859=>"010100101",
  34860=>"001010000",
  34861=>"011000001",
  34862=>"111100100",
  34863=>"000110111",
  34864=>"111000010",
  34865=>"111111110",
  34866=>"000000110",
  34867=>"100110011",
  34868=>"101000110",
  34869=>"111111000",
  34870=>"000001111",
  34871=>"000000111",
  34872=>"001111111",
  34873=>"101100000",
  34874=>"000010111",
  34875=>"111111111",
  34876=>"111100100",
  34877=>"111111111",
  34878=>"000000000",
  34879=>"111010011",
  34880=>"010001111",
  34881=>"000101011",
  34882=>"000111111",
  34883=>"000000001",
  34884=>"111000000",
  34885=>"111000000",
  34886=>"000000000",
  34887=>"011011000",
  34888=>"001111111",
  34889=>"110110000",
  34890=>"000000000",
  34891=>"111010000",
  34892=>"111000111",
  34893=>"011000110",
  34894=>"110111011",
  34895=>"101111000",
  34896=>"111110110",
  34897=>"100111010",
  34898=>"111111111",
  34899=>"000000000",
  34900=>"110000001",
  34901=>"111110110",
  34902=>"111011000",
  34903=>"010111001",
  34904=>"010011001",
  34905=>"101011110",
  34906=>"000010110",
  34907=>"001011000",
  34908=>"001111000",
  34909=>"000000010",
  34910=>"000111111",
  34911=>"000000010",
  34912=>"000000101",
  34913=>"111000000",
  34914=>"100000111",
  34915=>"001011001",
  34916=>"110100010",
  34917=>"100000010",
  34918=>"111000100",
  34919=>"111111000",
  34920=>"000100111",
  34921=>"100110010",
  34922=>"001001000",
  34923=>"000100111",
  34924=>"100100111",
  34925=>"111111111",
  34926=>"011011100",
  34927=>"111100000",
  34928=>"100100011",
  34929=>"000000000",
  34930=>"000000011",
  34931=>"110000000",
  34932=>"000111100",
  34933=>"100000000",
  34934=>"100101001",
  34935=>"000000000",
  34936=>"000001011",
  34937=>"111111111",
  34938=>"000000000",
  34939=>"111111111",
  34940=>"100100100",
  34941=>"000000000",
  34942=>"000011110",
  34943=>"010000000",
  34944=>"011100000",
  34945=>"010101011",
  34946=>"010000000",
  34947=>"011111111",
  34948=>"111001000",
  34949=>"000000010",
  34950=>"010111100",
  34951=>"111110010",
  34952=>"111100110",
  34953=>"111000000",
  34954=>"111011000",
  34955=>"000000000",
  34956=>"000000011",
  34957=>"110000111",
  34958=>"000111011",
  34959=>"111000000",
  34960=>"111110001",
  34961=>"000000111",
  34962=>"000111111",
  34963=>"000000000",
  34964=>"000011000",
  34965=>"000111011",
  34966=>"000000000",
  34967=>"110000011",
  34968=>"000111101",
  34969=>"010011000",
  34970=>"000010000",
  34971=>"000000000",
  34972=>"111111000",
  34973=>"101101000",
  34974=>"001100000",
  34975=>"000100000",
  34976=>"011100011",
  34977=>"000000111",
  34978=>"010000000",
  34979=>"111111111",
  34980=>"000000111",
  34981=>"111001000",
  34982=>"111000110",
  34983=>"000111110",
  34984=>"111000000",
  34985=>"000000111",
  34986=>"000000000",
  34987=>"000100110",
  34988=>"110011000",
  34989=>"110000000",
  34990=>"100001011",
  34991=>"111111111",
  34992=>"100000100",
  34993=>"001000111",
  34994=>"100000110",
  34995=>"000000000",
  34996=>"011001011",
  34997=>"010000000",
  34998=>"001100010",
  34999=>"001000000",
  35000=>"111100010",
  35001=>"001000000",
  35002=>"010101111",
  35003=>"100010000",
  35004=>"111111010",
  35005=>"100001111",
  35006=>"111111100",
  35007=>"111010000",
  35008=>"111000100",
  35009=>"110100101",
  35010=>"000000000",
  35011=>"001011100",
  35012=>"000000000",
  35013=>"010000000",
  35014=>"000110000",
  35015=>"111111111",
  35016=>"111111101",
  35017=>"000000110",
  35018=>"110110101",
  35019=>"111110100",
  35020=>"011110000",
  35021=>"110101000",
  35022=>"000000100",
  35023=>"101111111",
  35024=>"111101000",
  35025=>"001110110",
  35026=>"000100000",
  35027=>"001000000",
  35028=>"110111110",
  35029=>"100000101",
  35030=>"100100111",
  35031=>"000000010",
  35032=>"111111100",
  35033=>"000000011",
  35034=>"110010001",
  35035=>"100000000",
  35036=>"111101100",
  35037=>"111111000",
  35038=>"000001000",
  35039=>"001110110",
  35040=>"000100000",
  35041=>"000000000",
  35042=>"011001011",
  35043=>"111011011",
  35044=>"010010100",
  35045=>"111000000",
  35046=>"010101101",
  35047=>"000110110",
  35048=>"000001000",
  35049=>"111110001",
  35050=>"010000100",
  35051=>"000100111",
  35052=>"000100111",
  35053=>"100000000",
  35054=>"010110000",
  35055=>"000000000",
  35056=>"111100000",
  35057=>"011000000",
  35058=>"011000000",
  35059=>"000110000",
  35060=>"001001000",
  35061=>"100000000",
  35062=>"100000000",
  35063=>"000011111",
  35064=>"000000000",
  35065=>"001011100",
  35066=>"111010000",
  35067=>"000000010",
  35068=>"111011000",
  35069=>"010111111",
  35070=>"000000001",
  35071=>"100111101",
  35072=>"011111011",
  35073=>"000111111",
  35074=>"001000101",
  35075=>"000000000",
  35076=>"001011011",
  35077=>"000000100",
  35078=>"000000000",
  35079=>"000111111",
  35080=>"110010111",
  35081=>"000000000",
  35082=>"110111000",
  35083=>"000001111",
  35084=>"000000011",
  35085=>"000000001",
  35086=>"111111010",
  35087=>"000001011",
  35088=>"111001000",
  35089=>"011111000",
  35090=>"101000100",
  35091=>"000111111",
  35092=>"101010100",
  35093=>"000101100",
  35094=>"111001100",
  35095=>"000010010",
  35096=>"010010000",
  35097=>"111001101",
  35098=>"110011000",
  35099=>"000000000",
  35100=>"000000100",
  35101=>"000010010",
  35102=>"111110000",
  35103=>"000010111",
  35104=>"111000111",
  35105=>"110110000",
  35106=>"000000000",
  35107=>"011000000",
  35108=>"000000000",
  35109=>"011011110",
  35110=>"010011000",
  35111=>"111110001",
  35112=>"111001101",
  35113=>"010010000",
  35114=>"001000000",
  35115=>"000110101",
  35116=>"001011011",
  35117=>"110000011",
  35118=>"111011000",
  35119=>"000001001",
  35120=>"010000100",
  35121=>"011011001",
  35122=>"111101001",
  35123=>"000000000",
  35124=>"111010000",
  35125=>"000000001",
  35126=>"011111100",
  35127=>"000000101",
  35128=>"000111111",
  35129=>"111111111",
  35130=>"101000100",
  35131=>"000000111",
  35132=>"100110000",
  35133=>"111111000",
  35134=>"000000101",
  35135=>"110011011",
  35136=>"111000000",
  35137=>"011111111",
  35138=>"111111000",
  35139=>"000100110",
  35140=>"111011010",
  35141=>"000111111",
  35142=>"001101000",
  35143=>"111100111",
  35144=>"000011011",
  35145=>"110010010",
  35146=>"101000111",
  35147=>"000010000",
  35148=>"001111111",
  35149=>"101111000",
  35150=>"110110110",
  35151=>"000111111",
  35152=>"110111111",
  35153=>"011111111",
  35154=>"011000001",
  35155=>"001000000",
  35156=>"000000010",
  35157=>"010000011",
  35158=>"111110010",
  35159=>"001001000",
  35160=>"000110000",
  35161=>"001000011",
  35162=>"000011011",
  35163=>"110110110",
  35164=>"111101000",
  35165=>"001011010",
  35166=>"010000111",
  35167=>"000001110",
  35168=>"110010000",
  35169=>"100100101",
  35170=>"111001110",
  35171=>"000110100",
  35172=>"101110000",
  35173=>"111100111",
  35174=>"111111001",
  35175=>"110000111",
  35176=>"001100000",
  35177=>"000111000",
  35178=>"111010000",
  35179=>"000001000",
  35180=>"100110111",
  35181=>"110110101",
  35182=>"101101111",
  35183=>"000010111",
  35184=>"011011000",
  35185=>"010000000",
  35186=>"110111011",
  35187=>"000001111",
  35188=>"111110000",
  35189=>"110111100",
  35190=>"111111111",
  35191=>"011000001",
  35192=>"000101111",
  35193=>"111000000",
  35194=>"111101000",
  35195=>"000100001",
  35196=>"100110111",
  35197=>"110100000",
  35198=>"000010110",
  35199=>"110000010",
  35200=>"111111101",
  35201=>"000000000",
  35202=>"001010111",
  35203=>"110000101",
  35204=>"111110010",
  35205=>"111101111",
  35206=>"100110111",
  35207=>"111110000",
  35208=>"111110000",
  35209=>"000110000",
  35210=>"100000001",
  35211=>"110111001",
  35212=>"100100001",
  35213=>"000000011",
  35214=>"001000101",
  35215=>"110111001",
  35216=>"011011000",
  35217=>"010011010",
  35218=>"000000100",
  35219=>"010000000",
  35220=>"111011001",
  35221=>"111111000",
  35222=>"010010001",
  35223=>"011000001",
  35224=>"111011101",
  35225=>"000111111",
  35226=>"000000101",
  35227=>"100000111",
  35228=>"101100111",
  35229=>"110100111",
  35230=>"010000111",
  35231=>"000000011",
  35232=>"001100100",
  35233=>"101000111",
  35234=>"111011000",
  35235=>"111101101",
  35236=>"111010000",
  35237=>"111111110",
  35238=>"110111111",
  35239=>"010111111",
  35240=>"000111111",
  35241=>"001111111",
  35242=>"000000111",
  35243=>"010111111",
  35244=>"111101111",
  35245=>"111000111",
  35246=>"100010010",
  35247=>"110100101",
  35248=>"000101001",
  35249=>"000011000",
  35250=>"000110100",
  35251=>"100110010",
  35252=>"110010011",
  35253=>"111111010",
  35254=>"011010100",
  35255=>"011110000",
  35256=>"001001111",
  35257=>"110110001",
  35258=>"010010000",
  35259=>"010010000",
  35260=>"100100000",
  35261=>"111111000",
  35262=>"010000010",
  35263=>"111110000",
  35264=>"001001101",
  35265=>"001101100",
  35266=>"111111000",
  35267=>"100100100",
  35268=>"111101101",
  35269=>"110011000",
  35270=>"000111111",
  35271=>"111101000",
  35272=>"011111001",
  35273=>"000100111",
  35274=>"011011000",
  35275=>"101101110",
  35276=>"011110011",
  35277=>"011011111",
  35278=>"000000100",
  35279=>"110110000",
  35280=>"000111000",
  35281=>"100100000",
  35282=>"000000101",
  35283=>"111101111",
  35284=>"101101011",
  35285=>"110110110",
  35286=>"000001111",
  35287=>"000111111",
  35288=>"000000111",
  35289=>"101111111",
  35290=>"001001001",
  35291=>"000000111",
  35292=>"011100010",
  35293=>"000111111",
  35294=>"010010000",
  35295=>"000110111",
  35296=>"111001010",
  35297=>"011000000",
  35298=>"110000000",
  35299=>"101111000",
  35300=>"010000110",
  35301=>"010010000",
  35302=>"111110111",
  35303=>"011100110",
  35304=>"111000000",
  35305=>"001111111",
  35306=>"011111001",
  35307=>"111111000",
  35308=>"111101111",
  35309=>"000000111",
  35310=>"101100000",
  35311=>"001100000",
  35312=>"000000111",
  35313=>"011010000",
  35314=>"000101111",
  35315=>"000000000",
  35316=>"110011100",
  35317=>"010010010",
  35318=>"111000111",
  35319=>"111100111",
  35320=>"111001010",
  35321=>"000001001",
  35322=>"110010000",
  35323=>"101011000",
  35324=>"100101110",
  35325=>"100000100",
  35326=>"100100000",
  35327=>"100111000",
  35328=>"110111111",
  35329=>"101000000",
  35330=>"101000000",
  35331=>"000000000",
  35332=>"001111101",
  35333=>"111011111",
  35334=>"000000000",
  35335=>"101111111",
  35336=>"000111001",
  35337=>"001001000",
  35338=>"100000100",
  35339=>"101001111",
  35340=>"110110111",
  35341=>"000000000",
  35342=>"110100011",
  35343=>"000101110",
  35344=>"010110111",
  35345=>"000000000",
  35346=>"010100001",
  35347=>"111100000",
  35348=>"111111101",
  35349=>"111101001",
  35350=>"011100000",
  35351=>"111000000",
  35352=>"100000101",
  35353=>"001110011",
  35354=>"000111101",
  35355=>"000000111",
  35356=>"010111110",
  35357=>"010000001",
  35358=>"111011111",
  35359=>"110111001",
  35360=>"000000110",
  35361=>"010111001",
  35362=>"111101100",
  35363=>"010110111",
  35364=>"110111101",
  35365=>"011111111",
  35366=>"111001001",
  35367=>"100011110",
  35368=>"111111111",
  35369=>"001111111",
  35370=>"001000010",
  35371=>"011000000",
  35372=>"111111100",
  35373=>"101101100",
  35374=>"000000000",
  35375=>"000000000",
  35376=>"000111111",
  35377=>"000110111",
  35378=>"111111111",
  35379=>"000111111",
  35380=>"101000000",
  35381=>"000000000",
  35382=>"001010011",
  35383=>"111111010",
  35384=>"111111111",
  35385=>"010100110",
  35386=>"001000000",
  35387=>"000000000",
  35388=>"011011001",
  35389=>"000111101",
  35390=>"000000100",
  35391=>"000001110",
  35392=>"111001111",
  35393=>"101011111",
  35394=>"011011010",
  35395=>"011011001",
  35396=>"000000000",
  35397=>"101110000",
  35398=>"111000101",
  35399=>"011000000",
  35400=>"101110111",
  35401=>"110111111",
  35402=>"000010101",
  35403=>"100111011",
  35404=>"111000101",
  35405=>"010110001",
  35406=>"000110111",
  35407=>"000000010",
  35408=>"101000100",
  35409=>"101111111",
  35410=>"111111111",
  35411=>"000000110",
  35412=>"000000100",
  35413=>"111110110",
  35414=>"000111111",
  35415=>"111000010",
  35416=>"000000000",
  35417=>"011111101",
  35418=>"011111100",
  35419=>"111111111",
  35420=>"000000100",
  35421=>"100000000",
  35422=>"111111111",
  35423=>"000110000",
  35424=>"000011000",
  35425=>"110111111",
  35426=>"000000000",
  35427=>"100000000",
  35428=>"011111111",
  35429=>"011011111",
  35430=>"110011111",
  35431=>"000011101",
  35432=>"011001000",
  35433=>"111011110",
  35434=>"000001100",
  35435=>"111111101",
  35436=>"000000001",
  35437=>"000000000",
  35438=>"010011000",
  35439=>"101010111",
  35440=>"000011001",
  35441=>"001001101",
  35442=>"100000100",
  35443=>"100111111",
  35444=>"010001100",
  35445=>"111111000",
  35446=>"110000000",
  35447=>"101110111",
  35448=>"010000000",
  35449=>"000000000",
  35450=>"001111101",
  35451=>"000101111",
  35452=>"001110100",
  35453=>"000100000",
  35454=>"100000010",
  35455=>"001101111",
  35456=>"000010010",
  35457=>"000110000",
  35458=>"000001101",
  35459=>"110010101",
  35460=>"101001111",
  35461=>"001000000",
  35462=>"110100101",
  35463=>"000000100",
  35464=>"000101100",
  35465=>"001001000",
  35466=>"111000000",
  35467=>"100000100",
  35468=>"000111000",
  35469=>"111000000",
  35470=>"000001111",
  35471=>"001001010",
  35472=>"111101000",
  35473=>"111101101",
  35474=>"000000011",
  35475=>"000000110",
  35476=>"000000010",
  35477=>"100111111",
  35478=>"111101111",
  35479=>"100111101",
  35480=>"111111110",
  35481=>"111001000",
  35482=>"100000000",
  35483=>"001000000",
  35484=>"110110010",
  35485=>"000000000",
  35486=>"010111001",
  35487=>"101001101",
  35488=>"000001111",
  35489=>"001000000",
  35490=>"000000000",
  35491=>"111101111",
  35492=>"010111111",
  35493=>"110110000",
  35494=>"111110110",
  35495=>"111110111",
  35496=>"111011100",
  35497=>"010000000",
  35498=>"101101111",
  35499=>"110001101",
  35500=>"000000100",
  35501=>"101011111",
  35502=>"001101000",
  35503=>"111101011",
  35504=>"000001100",
  35505=>"001111011",
  35506=>"000100011",
  35507=>"001001111",
  35508=>"110011101",
  35509=>"111111000",
  35510=>"100100010",
  35511=>"111010101",
  35512=>"110111110",
  35513=>"000000110",
  35514=>"111000111",
  35515=>"110001001",
  35516=>"100111001",
  35517=>"101111110",
  35518=>"111111111",
  35519=>"111000100",
  35520=>"111000011",
  35521=>"101000000",
  35522=>"111111101",
  35523=>"010110100",
  35524=>"111010000",
  35525=>"000000000",
  35526=>"111111011",
  35527=>"100111110",
  35528=>"000000101",
  35529=>"000101000",
  35530=>"100000000",
  35531=>"000010000",
  35532=>"000000000",
  35533=>"000011111",
  35534=>"101000000",
  35535=>"010100100",
  35536=>"110111000",
  35537=>"010111101",
  35538=>"101000001",
  35539=>"100111000",
  35540=>"111101100",
  35541=>"001011001",
  35542=>"001001001",
  35543=>"111111111",
  35544=>"111001000",
  35545=>"000000000",
  35546=>"000000000",
  35547=>"001000100",
  35548=>"111011001",
  35549=>"110000101",
  35550=>"101111110",
  35551=>"111111111",
  35552=>"100010001",
  35553=>"111111111",
  35554=>"001001011",
  35555=>"000001100",
  35556=>"010100000",
  35557=>"111111101",
  35558=>"111001000",
  35559=>"000011011",
  35560=>"000001011",
  35561=>"100011110",
  35562=>"101000001",
  35563=>"101101001",
  35564=>"111111101",
  35565=>"101110111",
  35566=>"000011000",
  35567=>"000100110",
  35568=>"101000100",
  35569=>"001000010",
  35570=>"111111111",
  35571=>"000111111",
  35572=>"000110011",
  35573=>"000000001",
  35574=>"100001001",
  35575=>"110000111",
  35576=>"101111111",
  35577=>"111111111",
  35578=>"000111101",
  35579=>"000000000",
  35580=>"000111111",
  35581=>"000000100",
  35582=>"101101111",
  35583=>"011000000",
  35584=>"001010011",
  35585=>"000100000",
  35586=>"101000000",
  35587=>"001111010",
  35588=>"010011111",
  35589=>"110110000",
  35590=>"110110110",
  35591=>"111001001",
  35592=>"000110111",
  35593=>"000000001",
  35594=>"111001111",
  35595=>"001001001",
  35596=>"000110110",
  35597=>"000111111",
  35598=>"100000100",
  35599=>"110111110",
  35600=>"111001001",
  35601=>"111101111",
  35602=>"010110010",
  35603=>"111101100",
  35604=>"111101101",
  35605=>"001000110",
  35606=>"101000111",
  35607=>"101101000",
  35608=>"110101111",
  35609=>"010001001",
  35610=>"000001001",
  35611=>"000000100",
  35612=>"000101111",
  35613=>"110111111",
  35614=>"000000000",
  35615=>"110000010",
  35616=>"110111100",
  35617=>"010110111",
  35618=>"000000111",
  35619=>"000110110",
  35620=>"111011001",
  35621=>"101000000",
  35622=>"000001011",
  35623=>"111001111",
  35624=>"000000000",
  35625=>"001001001",
  35626=>"100000000",
  35627=>"110111000",
  35628=>"100001001",
  35629=>"111000111",
  35630=>"111000001",
  35631=>"000000000",
  35632=>"001100111",
  35633=>"011111011",
  35634=>"000110111",
  35635=>"101101111",
  35636=>"000000101",
  35637=>"000001110",
  35638=>"000110111",
  35639=>"111101001",
  35640=>"111111101",
  35641=>"111000000",
  35642=>"111000000",
  35643=>"111000000",
  35644=>"011100000",
  35645=>"110110111",
  35646=>"001000000",
  35647=>"000110010",
  35648=>"001000011",
  35649=>"000001000",
  35650=>"000111111",
  35651=>"010110000",
  35652=>"000110110",
  35653=>"111110000",
  35654=>"000110110",
  35655=>"110100000",
  35656=>"110110111",
  35657=>"001000101",
  35658=>"110001101",
  35659=>"111101001",
  35660=>"101101111",
  35661=>"110111010",
  35662=>"110111001",
  35663=>"011000001",
  35664=>"000011111",
  35665=>"111010000",
  35666=>"111000000",
  35667=>"011001001",
  35668=>"001000001",
  35669=>"111110110",
  35670=>"101011111",
  35671=>"101000000",
  35672=>"110010000",
  35673=>"011110111",
  35674=>"111000000",
  35675=>"101100100",
  35676=>"100000000",
  35677=>"011000010",
  35678=>"111111110",
  35679=>"010110100",
  35680=>"000000111",
  35681=>"000000000",
  35682=>"001001001",
  35683=>"111011001",
  35684=>"111000000",
  35685=>"000011111",
  35686=>"101001000",
  35687=>"001000001",
  35688=>"111001001",
  35689=>"111010111",
  35690=>"000010000",
  35691=>"110100001",
  35692=>"111111101",
  35693=>"111001000",
  35694=>"110110010",
  35695=>"001001111",
  35696=>"011100101",
  35697=>"001000111",
  35698=>"001010111",
  35699=>"111001111",
  35700=>"110001000",
  35701=>"000001001",
  35702=>"111111001",
  35703=>"000111110",
  35704=>"101001001",
  35705=>"110111001",
  35706=>"001001101",
  35707=>"010111111",
  35708=>"111100000",
  35709=>"100100000",
  35710=>"111110001",
  35711=>"000110110",
  35712=>"000000111",
  35713=>"111000000",
  35714=>"000111111",
  35715=>"000100000",
  35716=>"011001000",
  35717=>"000001001",
  35718=>"011111011",
  35719=>"111001000",
  35720=>"110011011",
  35721=>"111001001",
  35722=>"111001000",
  35723=>"111110000",
  35724=>"000110110",
  35725=>"011111111",
  35726=>"010010010",
  35727=>"111001001",
  35728=>"110110100",
  35729=>"001111111",
  35730=>"000111111",
  35731=>"000000001",
  35732=>"111010000",
  35733=>"001111110",
  35734=>"110001001",
  35735=>"000011011",
  35736=>"010110001",
  35737=>"110000000",
  35738=>"011111111",
  35739=>"010010110",
  35740=>"000110110",
  35741=>"111111010",
  35742=>"001001111",
  35743=>"001001001",
  35744=>"011110111",
  35745=>"000001000",
  35746=>"010000000",
  35747=>"000000110",
  35748=>"000110111",
  35749=>"100001011",
  35750=>"001000000",
  35751=>"000010110",
  35752=>"111111111",
  35753=>"001010100",
  35754=>"101101000",
  35755=>"001001000",
  35756=>"101100001",
  35757=>"111111010",
  35758=>"111100100",
  35759=>"111110110",
  35760=>"111110000",
  35761=>"100010000",
  35762=>"111000000",
  35763=>"110000000",
  35764=>"011001111",
  35765=>"000000110",
  35766=>"000000110",
  35767=>"000110011",
  35768=>"000100111",
  35769=>"010010001",
  35770=>"000000000",
  35771=>"100000000",
  35772=>"111111111",
  35773=>"011110110",
  35774=>"001111011",
  35775=>"111110111",
  35776=>"001000001",
  35777=>"011101111",
  35778=>"000111111",
  35779=>"011111011",
  35780=>"000000000",
  35781=>"111000000",
  35782=>"010110101",
  35783=>"011000001",
  35784=>"000000001",
  35785=>"101000001",
  35786=>"000010110",
  35787=>"111011111",
  35788=>"111001000",
  35789=>"010000000",
  35790=>"011001101",
  35791=>"000000000",
  35792=>"010000010",
  35793=>"010110110",
  35794=>"001000001",
  35795=>"110010010",
  35796=>"101001101",
  35797=>"110001110",
  35798=>"100000100",
  35799=>"110110000",
  35800=>"111001001",
  35801=>"000000110",
  35802=>"110111011",
  35803=>"101001001",
  35804=>"001001111",
  35805=>"111001010",
  35806=>"000001101",
  35807=>"111111111",
  35808=>"101000000",
  35809=>"001010011",
  35810=>"001000000",
  35811=>"000011001",
  35812=>"000101101",
  35813=>"110000000",
  35814=>"000110110",
  35815=>"000001011",
  35816=>"110111111",
  35817=>"111111101",
  35818=>"111100101",
  35819=>"000000111",
  35820=>"000000000",
  35821=>"010111111",
  35822=>"111011000",
  35823=>"000000000",
  35824=>"010000001",
  35825=>"111000011",
  35826=>"001000000",
  35827=>"110000111",
  35828=>"000101100",
  35829=>"101000000",
  35830=>"011000101",
  35831=>"111101000",
  35832=>"000000000",
  35833=>"110101100",
  35834=>"111010000",
  35835=>"000101100",
  35836=>"111110101",
  35837=>"000000000",
  35838=>"110110110",
  35839=>"111001101",
  35840=>"100010000",
  35841=>"000000001",
  35842=>"011001111",
  35843=>"011111000",
  35844=>"000100000",
  35845=>"000010001",
  35846=>"000010010",
  35847=>"101110011",
  35848=>"000110100",
  35849=>"111101110",
  35850=>"011000001",
  35851=>"000000000",
  35852=>"000111010",
  35853=>"111101001",
  35854=>"101001000",
  35855=>"000000011",
  35856=>"110111001",
  35857=>"111100111",
  35858=>"111100000",
  35859=>"111101101",
  35860=>"010101111",
  35861=>"111101111",
  35862=>"101000101",
  35863=>"011100101",
  35864=>"110101010",
  35865=>"000110110",
  35866=>"000111111",
  35867=>"000010000",
  35868=>"111011001",
  35869=>"101101111",
  35870=>"011011000",
  35871=>"101000000",
  35872=>"011101001",
  35873=>"010000100",
  35874=>"111000000",
  35875=>"000111010",
  35876=>"110000011",
  35877=>"000000000",
  35878=>"000100111",
  35879=>"110100010",
  35880=>"000010110",
  35881=>"010111011",
  35882=>"111010100",
  35883=>"010010011",
  35884=>"000011000",
  35885=>"000001000",
  35886=>"101111111",
  35887=>"100010000",
  35888=>"010001001",
  35889=>"111100110",
  35890=>"111110100",
  35891=>"101101000",
  35892=>"000001101",
  35893=>"100000000",
  35894=>"110001111",
  35895=>"001111000",
  35896=>"111001100",
  35897=>"000000000",
  35898=>"000110111",
  35899=>"100101001",
  35900=>"011110110",
  35901=>"111111111",
  35902=>"100000111",
  35903=>"111110111",
  35904=>"111011110",
  35905=>"000000001",
  35906=>"101111010",
  35907=>"111001000",
  35908=>"000100111",
  35909=>"000000000",
  35910=>"111111111",
  35911=>"010000101",
  35912=>"101000000",
  35913=>"110011001",
  35914=>"101001101",
  35915=>"111101001",
  35916=>"111000100",
  35917=>"011110000",
  35918=>"111100101",
  35919=>"110111010",
  35920=>"101101101",
  35921=>"111111111",
  35922=>"101000001",
  35923=>"000000000",
  35924=>"011010000",
  35925=>"111000001",
  35926=>"110011001",
  35927=>"000000011",
  35928=>"101001001",
  35929=>"111100110",
  35930=>"111100100",
  35931=>"000100010",
  35932=>"000000000",
  35933=>"000001111",
  35934=>"111010110",
  35935=>"100000001",
  35936=>"111111111",
  35937=>"000011111",
  35938=>"100100111",
  35939=>"110101111",
  35940=>"000111000",
  35941=>"001001000",
  35942=>"110111000",
  35943=>"000000000",
  35944=>"101111011",
  35945=>"100000111",
  35946=>"101111111",
  35947=>"111111001",
  35948=>"000001111",
  35949=>"110101000",
  35950=>"000001000",
  35951=>"000010000",
  35952=>"001011001",
  35953=>"010001001",
  35954=>"111100100",
  35955=>"000101000",
  35956=>"101111000",
  35957=>"001000000",
  35958=>"000100000",
  35959=>"011000000",
  35960=>"010000100",
  35961=>"001100000",
  35962=>"101010011",
  35963=>"100100101",
  35964=>"101110110",
  35965=>"010000000",
  35966=>"100101111",
  35967=>"000001101",
  35968=>"101001011",
  35969=>"010000000",
  35970=>"000100100",
  35971=>"001110111",
  35972=>"100011010",
  35973=>"111110001",
  35974=>"000000000",
  35975=>"101001001",
  35976=>"000110110",
  35977=>"001100000",
  35978=>"010001000",
  35979=>"010110111",
  35980=>"101000101",
  35981=>"111101000",
  35982=>"111110110",
  35983=>"001000110",
  35984=>"000100000",
  35985=>"101000000",
  35986=>"101000000",
  35987=>"011000011",
  35988=>"100000000",
  35989=>"000000001",
  35990=>"110111000",
  35991=>"110110000",
  35992=>"110111010",
  35993=>"011000011",
  35994=>"100011101",
  35995=>"000000011",
  35996=>"011001011",
  35997=>"111111111",
  35998=>"010010010",
  35999=>"101100001",
  36000=>"101100110",
  36001=>"110001111",
  36002=>"110111010",
  36003=>"001011000",
  36004=>"110011010",
  36005=>"100110100",
  36006=>"011001001",
  36007=>"000010010",
  36008=>"110000011",
  36009=>"110101111",
  36010=>"101100111",
  36011=>"010000101",
  36012=>"111110100",
  36013=>"000000010",
  36014=>"000000000",
  36015=>"101000000",
  36016=>"111001101",
  36017=>"101000100",
  36018=>"000010010",
  36019=>"010010000",
  36020=>"111011101",
  36021=>"100101110",
  36022=>"111111000",
  36023=>"111111001",
  36024=>"101011000",
  36025=>"101100000",
  36026=>"010000100",
  36027=>"010111100",
  36028=>"010010000",
  36029=>"111000111",
  36030=>"000011011",
  36031=>"111101111",
  36032=>"001101011",
  36033=>"000000000",
  36034=>"111111000",
  36035=>"110011100",
  36036=>"000001011",
  36037=>"110100001",
  36038=>"000111011",
  36039=>"000100000",
  36040=>"111111111",
  36041=>"100000010",
  36042=>"001101111",
  36043=>"001000101",
  36044=>"111100100",
  36045=>"101011011",
  36046=>"111111011",
  36047=>"111101101",
  36048=>"111101111",
  36049=>"011110000",
  36050=>"000010111",
  36051=>"010000000",
  36052=>"001000000",
  36053=>"011100010",
  36054=>"000100100",
  36055=>"100010001",
  36056=>"000000000",
  36057=>"000011111",
  36058=>"110001011",
  36059=>"111100111",
  36060=>"000100100",
  36061=>"001111011",
  36062=>"010011010",
  36063=>"111010000",
  36064=>"000101111",
  36065=>"011000000",
  36066=>"111010111",
  36067=>"000001011",
  36068=>"001000101",
  36069=>"010000011",
  36070=>"101001000",
  36071=>"000000000",
  36072=>"000101011",
  36073=>"000000101",
  36074=>"110000110",
  36075=>"000110111",
  36076=>"101111111",
  36077=>"111100111",
  36078=>"000010100",
  36079=>"000000000",
  36080=>"000000100",
  36081=>"110000000",
  36082=>"101011010",
  36083=>"001100011",
  36084=>"000011011",
  36085=>"111101111",
  36086=>"000000000",
  36087=>"110110111",
  36088=>"111111111",
  36089=>"110110001",
  36090=>"101101101",
  36091=>"000001001",
  36092=>"000010011",
  36093=>"111000000",
  36094=>"000011001",
  36095=>"111011000",
  36096=>"110110110",
  36097=>"000101110",
  36098=>"101101000",
  36099=>"000000110",
  36100=>"011011010",
  36101=>"010010010",
  36102=>"100001111",
  36103=>"011000000",
  36104=>"010110111",
  36105=>"001010000",
  36106=>"011110110",
  36107=>"111111010",
  36108=>"000111111",
  36109=>"101000000",
  36110=>"000000001",
  36111=>"100000111",
  36112=>"000000000",
  36113=>"110010111",
  36114=>"000000000",
  36115=>"000000000",
  36116=>"111011000",
  36117=>"011011000",
  36118=>"110110110",
  36119=>"111010010",
  36120=>"101001110",
  36121=>"100001000",
  36122=>"110110000",
  36123=>"000100110",
  36124=>"100000101",
  36125=>"111010000",
  36126=>"111110000",
  36127=>"111111111",
  36128=>"111111000",
  36129=>"010111000",
  36130=>"000000111",
  36131=>"110100000",
  36132=>"001001001",
  36133=>"111101001",
  36134=>"000000101",
  36135=>"000000000",
  36136=>"101000100",
  36137=>"010111000",
  36138=>"001001000",
  36139=>"010011110",
  36140=>"000101001",
  36141=>"111100000",
  36142=>"110111111",
  36143=>"010001001",
  36144=>"111111111",
  36145=>"001011001",
  36146=>"110000101",
  36147=>"001000001",
  36148=>"000010111",
  36149=>"111111010",
  36150=>"010010000",
  36151=>"100100101",
  36152=>"010100100",
  36153=>"001000100",
  36154=>"111101111",
  36155=>"110100010",
  36156=>"011010000",
  36157=>"111111111",
  36158=>"000111101",
  36159=>"011011011",
  36160=>"100101100",
  36161=>"010010010",
  36162=>"000000000",
  36163=>"010011110",
  36164=>"101111010",
  36165=>"000101111",
  36166=>"101000000",
  36167=>"101111000",
  36168=>"000101001",
  36169=>"111101111",
  36170=>"101001101",
  36171=>"100101100",
  36172=>"101011111",
  36173=>"110011011",
  36174=>"000110110",
  36175=>"111011010",
  36176=>"111111010",
  36177=>"010010000",
  36178=>"001011000",
  36179=>"111001000",
  36180=>"111110010",
  36181=>"000110110",
  36182=>"110100110",
  36183=>"000010010",
  36184=>"110111110",
  36185=>"001001000",
  36186=>"000100000",
  36187=>"000100110",
  36188=>"100000101",
  36189=>"001001001",
  36190=>"001000000",
  36191=>"010010001",
  36192=>"000110011",
  36193=>"011010010",
  36194=>"000110100",
  36195=>"101001001",
  36196=>"110111111",
  36197=>"000100100",
  36198=>"111111011",
  36199=>"011111011",
  36200=>"111111101",
  36201=>"011000000",
  36202=>"010111111",
  36203=>"000111111",
  36204=>"101001001",
  36205=>"000000010",
  36206=>"000000000",
  36207=>"011000110",
  36208=>"101000001",
  36209=>"000000010",
  36210=>"010010000",
  36211=>"000000000",
  36212=>"111111000",
  36213=>"100100111",
  36214=>"110011000",
  36215=>"111111110",
  36216=>"100100010",
  36217=>"111000110",
  36218=>"100111100",
  36219=>"010000000",
  36220=>"000110010",
  36221=>"111100100",
  36222=>"010110001",
  36223=>"010110010",
  36224=>"000000000",
  36225=>"010111000",
  36226=>"111000000",
  36227=>"101101111",
  36228=>"010011101",
  36229=>"101101111",
  36230=>"110011011",
  36231=>"000000000",
  36232=>"100111101",
  36233=>"110010000",
  36234=>"001000000",
  36235=>"011010000",
  36236=>"010010010",
  36237=>"111111010",
  36238=>"101001001",
  36239=>"111001001",
  36240=>"110110100",
  36241=>"000000000",
  36242=>"000000010",
  36243=>"111111000",
  36244=>"100001111",
  36245=>"000011000",
  36246=>"000000000",
  36247=>"010111111",
  36248=>"011111011",
  36249=>"010011011",
  36250=>"101000100",
  36251=>"101111101",
  36252=>"001111111",
  36253=>"100000001",
  36254=>"111001000",
  36255=>"111100001",
  36256=>"000000011",
  36257=>"000010010",
  36258=>"000000100",
  36259=>"000111101",
  36260=>"111011000",
  36261=>"100001100",
  36262=>"111111101",
  36263=>"100000000",
  36264=>"010000111",
  36265=>"000100010",
  36266=>"000000000",
  36267=>"000100100",
  36268=>"101011101",
  36269=>"101110111",
  36270=>"110110100",
  36271=>"000000010",
  36272=>"000000101",
  36273=>"001011000",
  36274=>"111010110",
  36275=>"100010010",
  36276=>"111111011",
  36277=>"010000000",
  36278=>"000001111",
  36279=>"000101010",
  36280=>"000001000",
  36281=>"000110101",
  36282=>"100110000",
  36283=>"111111111",
  36284=>"010000111",
  36285=>"111111111",
  36286=>"110110110",
  36287=>"011010010",
  36288=>"001000101",
  36289=>"000010010",
  36290=>"101011111",
  36291=>"110110100",
  36292=>"001000000",
  36293=>"110110100",
  36294=>"000011111",
  36295=>"000000101",
  36296=>"000000000",
  36297=>"100000001",
  36298=>"000000111",
  36299=>"110111010",
  36300=>"011111001",
  36301=>"000010000",
  36302=>"010100100",
  36303=>"111011101",
  36304=>"111110110",
  36305=>"010000011",
  36306=>"000000000",
  36307=>"111100000",
  36308=>"101000100",
  36309=>"111101110",
  36310=>"000000011",
  36311=>"000000000",
  36312=>"000000000",
  36313=>"000000000",
  36314=>"000100101",
  36315=>"101001000",
  36316=>"011110110",
  36317=>"011111110",
  36318=>"111111111",
  36319=>"111111000",
  36320=>"110010011",
  36321=>"111111100",
  36322=>"011111000",
  36323=>"111000000",
  36324=>"000000111",
  36325=>"110111010",
  36326=>"000110010",
  36327=>"001111100",
  36328=>"111100000",
  36329=>"011001000",
  36330=>"011011011",
  36331=>"000110010",
  36332=>"010111111",
  36333=>"000010111",
  36334=>"100010000",
  36335=>"100111111",
  36336=>"110100100",
  36337=>"011010001",
  36338=>"000100111",
  36339=>"100100100",
  36340=>"010110010",
  36341=>"111101000",
  36342=>"000000000",
  36343=>"111010000",
  36344=>"100111011",
  36345=>"000100000",
  36346=>"011000000",
  36347=>"111111100",
  36348=>"101000101",
  36349=>"010111010",
  36350=>"110111000",
  36351=>"000000000",
  36352=>"110100111",
  36353=>"110010111",
  36354=>"101000100",
  36355=>"001000001",
  36356=>"010000000",
  36357=>"110101111",
  36358=>"001000111",
  36359=>"000000111",
  36360=>"110001001",
  36361=>"010000000",
  36362=>"100110111",
  36363=>"111101100",
  36364=>"000000110",
  36365=>"010001100",
  36366=>"111101100",
  36367=>"111111000",
  36368=>"010000000",
  36369=>"000000111",
  36370=>"111101111",
  36371=>"000000011",
  36372=>"011110111",
  36373=>"001110100",
  36374=>"010000011",
  36375=>"010010101",
  36376=>"101100000",
  36377=>"000110000",
  36378=>"000000001",
  36379=>"100010111",
  36380=>"110011011",
  36381=>"000110100",
  36382=>"010101111",
  36383=>"000000000",
  36384=>"000111000",
  36385=>"010100111",
  36386=>"101101100",
  36387=>"010111000",
  36388=>"100000001",
  36389=>"111110010",
  36390=>"000011010",
  36391=>"000000001",
  36392=>"111001011",
  36393=>"000000111",
  36394=>"010000111",
  36395=>"000010010",
  36396=>"111101100",
  36397=>"100000001",
  36398=>"110010000",
  36399=>"010000000",
  36400=>"110001000",
  36401=>"110000100",
  36402=>"000000011",
  36403=>"000001001",
  36404=>"010101111",
  36405=>"100110110",
  36406=>"000110010",
  36407=>"111110000",
  36408=>"011101110",
  36409=>"101000011",
  36410=>"111100010",
  36411=>"000100100",
  36412=>"011110110",
  36413=>"111110110",
  36414=>"101000000",
  36415=>"111100101",
  36416=>"011000000",
  36417=>"011010111",
  36418=>"101000101",
  36419=>"111110010",
  36420=>"111011010",
  36421=>"001000000",
  36422=>"010000101",
  36423=>"000111011",
  36424=>"000011110",
  36425=>"111111010",
  36426=>"101101001",
  36427=>"111000110",
  36428=>"000000100",
  36429=>"101000011",
  36430=>"010000000",
  36431=>"111111101",
  36432=>"000000111",
  36433=>"010010000",
  36434=>"000000110",
  36435=>"110001010",
  36436=>"000010010",
  36437=>"111010010",
  36438=>"111100110",
  36439=>"001000000",
  36440=>"000000011",
  36441=>"001000000",
  36442=>"101101011",
  36443=>"110000110",
  36444=>"101000110",
  36445=>"100101110",
  36446=>"111111111",
  36447=>"001101010",
  36448=>"010000111",
  36449=>"000111111",
  36450=>"111000010",
  36451=>"000110111",
  36452=>"111001011",
  36453=>"010001011",
  36454=>"010111100",
  36455=>"110111000",
  36456=>"001101100",
  36457=>"011100011",
  36458=>"000000010",
  36459=>"010111000",
  36460=>"000111111",
  36461=>"101111101",
  36462=>"000000101",
  36463=>"110001111",
  36464=>"000001011",
  36465=>"000101101",
  36466=>"000011001",
  36467=>"000011000",
  36468=>"011101001",
  36469=>"010001000",
  36470=>"101001101",
  36471=>"000000000",
  36472=>"111000001",
  36473=>"000000110",
  36474=>"101000001",
  36475=>"101100100",
  36476=>"100110011",
  36477=>"111100010",
  36478=>"000111011",
  36479=>"101101111",
  36480=>"111110000",
  36481=>"111000000",
  36482=>"000110000",
  36483=>"000111111",
  36484=>"100000111",
  36485=>"110111100",
  36486=>"110011001",
  36487=>"100100100",
  36488=>"000000100",
  36489=>"101101101",
  36490=>"100000000",
  36491=>"000010000",
  36492=>"111110000",
  36493=>"000000100",
  36494=>"101111001",
  36495=>"000000001",
  36496=>"011011100",
  36497=>"000010111",
  36498=>"100001000",
  36499=>"010110000",
  36500=>"101101000",
  36501=>"000000100",
  36502=>"011011001",
  36503=>"110100100",
  36504=>"000100101",
  36505=>"001110000",
  36506=>"000010000",
  36507=>"100000111",
  36508=>"111100100",
  36509=>"000000111",
  36510=>"000001000",
  36511=>"000010010",
  36512=>"011111110",
  36513=>"001111010",
  36514=>"010011000",
  36515=>"000110010",
  36516=>"101000111",
  36517=>"111100001",
  36518=>"000000000",
  36519=>"100100111",
  36520=>"010010101",
  36521=>"101000101",
  36522=>"111101011",
  36523=>"100000111",
  36524=>"010111111",
  36525=>"001000000",
  36526=>"001011011",
  36527=>"000111011",
  36528=>"111111000",
  36529=>"100001100",
  36530=>"111101101",
  36531=>"000111011",
  36532=>"111111110",
  36533=>"000110110",
  36534=>"000101000",
  36535=>"111000000",
  36536=>"100011011",
  36537=>"001001001",
  36538=>"000111111",
  36539=>"111111100",
  36540=>"010010110",
  36541=>"010001101",
  36542=>"000000111",
  36543=>"000010010",
  36544=>"000110010",
  36545=>"000111111",
  36546=>"111010000",
  36547=>"111001100",
  36548=>"001000101",
  36549=>"011011000",
  36550=>"100100000",
  36551=>"010111011",
  36552=>"000001001",
  36553=>"111010110",
  36554=>"011011000",
  36555=>"001001101",
  36556=>"000010000",
  36557=>"101011010",
  36558=>"000000000",
  36559=>"000111111",
  36560=>"111000000",
  36561=>"110011010",
  36562=>"010000001",
  36563=>"000000100",
  36564=>"110000101",
  36565=>"001100111",
  36566=>"101000011",
  36567=>"010101010",
  36568=>"010010000",
  36569=>"000000100",
  36570=>"110111001",
  36571=>"101000101",
  36572=>"000000110",
  36573=>"100000000",
  36574=>"000000000",
  36575=>"111101111",
  36576=>"010000101",
  36577=>"001000001",
  36578=>"011111000",
  36579=>"010101011",
  36580=>"000000001",
  36581=>"000011010",
  36582=>"000000001",
  36583=>"000101111",
  36584=>"111000010",
  36585=>"000111101",
  36586=>"000001111",
  36587=>"001001000",
  36588=>"000100111",
  36589=>"000101100",
  36590=>"001111111",
  36591=>"010111011",
  36592=>"011000000",
  36593=>"111010000",
  36594=>"000000001",
  36595=>"001100100",
  36596=>"001000011",
  36597=>"111000111",
  36598=>"010000000",
  36599=>"110101101",
  36600=>"110001000",
  36601=>"001110010",
  36602=>"011111001",
  36603=>"111001110",
  36604=>"110011100",
  36605=>"000111010",
  36606=>"000001010",
  36607=>"110000111",
  36608=>"000001100",
  36609=>"000010000",
  36610=>"000000100",
  36611=>"000000100",
  36612=>"111101100",
  36613=>"010101001",
  36614=>"100111111",
  36615=>"001000011",
  36616=>"101111011",
  36617=>"000101111",
  36618=>"000000001",
  36619=>"010111000",
  36620=>"000011111",
  36621=>"111111110",
  36622=>"100000011",
  36623=>"011111000",
  36624=>"101000001",
  36625=>"000000001",
  36626=>"000000101",
  36627=>"101100111",
  36628=>"101101011",
  36629=>"111111000",
  36630=>"111100100",
  36631=>"000001001",
  36632=>"000100001",
  36633=>"111111111",
  36634=>"000101000",
  36635=>"100100011",
  36636=>"101101011",
  36637=>"111111111",
  36638=>"110100000",
  36639=>"101000000",
  36640=>"111101000",
  36641=>"111111010",
  36642=>"000010100",
  36643=>"000000011",
  36644=>"100100110",
  36645=>"011011011",
  36646=>"111011000",
  36647=>"000100111",
  36648=>"010000000",
  36649=>"111111111",
  36650=>"110111011",
  36651=>"001000010",
  36652=>"011111000",
  36653=>"100011111",
  36654=>"011110000",
  36655=>"000000000",
  36656=>"101100000",
  36657=>"000000100",
  36658=>"000100010",
  36659=>"001001000",
  36660=>"100100001",
  36661=>"111111111",
  36662=>"110100001",
  36663=>"000000000",
  36664=>"001011010",
  36665=>"100000000",
  36666=>"000000000",
  36667=>"000111101",
  36668=>"010001101",
  36669=>"100111101",
  36670=>"101101000",
  36671=>"011011010",
  36672=>"101011111",
  36673=>"111101111",
  36674=>"000000001",
  36675=>"111111101",
  36676=>"111110110",
  36677=>"100010111",
  36678=>"101100100",
  36679=>"011111111",
  36680=>"011001110",
  36681=>"101111111",
  36682=>"100100111",
  36683=>"111000000",
  36684=>"111111010",
  36685=>"011011011",
  36686=>"010100100",
  36687=>"111111011",
  36688=>"111000100",
  36689=>"010111111",
  36690=>"000000000",
  36691=>"001010110",
  36692=>"000000000",
  36693=>"110100000",
  36694=>"011111111",
  36695=>"000000101",
  36696=>"010000000",
  36697=>"000000011",
  36698=>"110010001",
  36699=>"111111010",
  36700=>"100000101",
  36701=>"000000000",
  36702=>"010010000",
  36703=>"111111001",
  36704=>"111111010",
  36705=>"110110010",
  36706=>"111101111",
  36707=>"110100000",
  36708=>"000000110",
  36709=>"001000111",
  36710=>"000000100",
  36711=>"100000111",
  36712=>"011011000",
  36713=>"111100000",
  36714=>"010011010",
  36715=>"110100000",
  36716=>"000000000",
  36717=>"000000000",
  36718=>"000000000",
  36719=>"000000111",
  36720=>"111111100",
  36721=>"000101111",
  36722=>"011000100",
  36723=>"000000110",
  36724=>"101111111",
  36725=>"100100000",
  36726=>"110111100",
  36727=>"111110100",
  36728=>"011111001",
  36729=>"011110100",
  36730=>"111011011",
  36731=>"000000011",
  36732=>"001000010",
  36733=>"100100000",
  36734=>"100000000",
  36735=>"111111111",
  36736=>"111111010",
  36737=>"110101000",
  36738=>"111010011",
  36739=>"111111000",
  36740=>"111101011",
  36741=>"111111110",
  36742=>"111100111",
  36743=>"011110110",
  36744=>"101001000",
  36745=>"001011110",
  36746=>"100000111",
  36747=>"000000000",
  36748=>"010010000",
  36749=>"011111111",
  36750=>"000000001",
  36751=>"000001101",
  36752=>"100101101",
  36753=>"111011011",
  36754=>"101101000",
  36755=>"101001001",
  36756=>"101111101",
  36757=>"000000111",
  36758=>"010111011",
  36759=>"000111010",
  36760=>"111101101",
  36761=>"111111111",
  36762=>"111011111",
  36763=>"000000001",
  36764=>"000000000",
  36765=>"011111111",
  36766=>"101111111",
  36767=>"000000000",
  36768=>"111111110",
  36769=>"011111000",
  36770=>"101111100",
  36771=>"000001100",
  36772=>"000000000",
  36773=>"110011011",
  36774=>"011111011",
  36775=>"000000000",
  36776=>"000010111",
  36777=>"101000000",
  36778=>"111111010",
  36779=>"100100111",
  36780=>"110011100",
  36781=>"100000101",
  36782=>"000001001",
  36783=>"010011111",
  36784=>"011110001",
  36785=>"001100110",
  36786=>"011111011",
  36787=>"001000100",
  36788=>"100111010",
  36789=>"011101000",
  36790=>"011111100",
  36791=>"111111000",
  36792=>"011100111",
  36793=>"111101000",
  36794=>"000010111",
  36795=>"000101111",
  36796=>"111101000",
  36797=>"111111111",
  36798=>"111111111",
  36799=>"100101011",
  36800=>"000000100",
  36801=>"000000000",
  36802=>"000001011",
  36803=>"100010110",
  36804=>"000100010",
  36805=>"000000110",
  36806=>"111010111",
  36807=>"111011010",
  36808=>"000000111",
  36809=>"010111100",
  36810=>"100101101",
  36811=>"011111111",
  36812=>"000000000",
  36813=>"110100000",
  36814=>"100101101",
  36815=>"000000000",
  36816=>"110110110",
  36817=>"111111111",
  36818=>"111011010",
  36819=>"111111111",
  36820=>"000000000",
  36821=>"000100100",
  36822=>"100100011",
  36823=>"011011010",
  36824=>"101000011",
  36825=>"000110000",
  36826=>"111111111",
  36827=>"000000011",
  36828=>"001011001",
  36829=>"011100000",
  36830=>"011111010",
  36831=>"100111010",
  36832=>"000000000",
  36833=>"000000100",
  36834=>"000011111",
  36835=>"001100110",
  36836=>"000000000",
  36837=>"101111000",
  36838=>"111111011",
  36839=>"011100100",
  36840=>"000100111",
  36841=>"100101001",
  36842=>"000000000",
  36843=>"011001100",
  36844=>"000000110",
  36845=>"010000000",
  36846=>"111111000",
  36847=>"001000000",
  36848=>"110111011",
  36849=>"000011111",
  36850=>"000111100",
  36851=>"101001100",
  36852=>"110110000",
  36853=>"101000011",
  36854=>"000000000",
  36855=>"001111011",
  36856=>"000010111",
  36857=>"100000000",
  36858=>"111111111",
  36859=>"011101111",
  36860=>"111100000",
  36861=>"001111011",
  36862=>"111111001",
  36863=>"000000000",
  36864=>"111111100",
  36865=>"111111000",
  36866=>"000000100",
  36867=>"010111000",
  36868=>"111111111",
  36869=>"000000001",
  36870=>"110100011",
  36871=>"000000000",
  36872=>"000010000",
  36873=>"000000000",
  36874=>"011011111",
  36875=>"001001000",
  36876=>"000000000",
  36877=>"111111001",
  36878=>"100111100",
  36879=>"100000001",
  36880=>"000000100",
  36881=>"000111111",
  36882=>"110110001",
  36883=>"000010010",
  36884=>"010111110",
  36885=>"111111111",
  36886=>"111111111",
  36887=>"111111010",
  36888=>"100000000",
  36889=>"000000000",
  36890=>"000000000",
  36891=>"111100111",
  36892=>"000000000",
  36893=>"110111111",
  36894=>"011101111",
  36895=>"010011101",
  36896=>"000000000",
  36897=>"111010111",
  36898=>"010001111",
  36899=>"011000000",
  36900=>"011001011",
  36901=>"000000001",
  36902=>"110010000",
  36903=>"011001001",
  36904=>"111111000",
  36905=>"110001100",
  36906=>"000000001",
  36907=>"000001000",
  36908=>"001010111",
  36909=>"111111111",
  36910=>"111111111",
  36911=>"000101100",
  36912=>"000000000",
  36913=>"001000010",
  36914=>"001010111",
  36915=>"100111111",
  36916=>"111111101",
  36917=>"111010001",
  36918=>"111111000",
  36919=>"011011111",
  36920=>"010111110",
  36921=>"000000110",
  36922=>"010000011",
  36923=>"001000000",
  36924=>"000000000",
  36925=>"111111111",
  36926=>"000000001",
  36927=>"110101001",
  36928=>"000000110",
  36929=>"000000000",
  36930=>"011000000",
  36931=>"011000100",
  36932=>"111111111",
  36933=>"001001001",
  36934=>"100101111",
  36935=>"111111101",
  36936=>"011111111",
  36937=>"111001000",
  36938=>"000000000",
  36939=>"000000000",
  36940=>"000000011",
  36941=>"000100100",
  36942=>"000011111",
  36943=>"000000111",
  36944=>"010010110",
  36945=>"111111111",
  36946=>"000010111",
  36947=>"001000000",
  36948=>"010111100",
  36949=>"111111111",
  36950=>"000011000",
  36951=>"000000000",
  36952=>"010110110",
  36953=>"111110110",
  36954=>"000011111",
  36955=>"111011000",
  36956=>"111111111",
  36957=>"000000000",
  36958=>"111111111",
  36959=>"000000110",
  36960=>"000000000",
  36961=>"010111011",
  36962=>"000000001",
  36963=>"000100011",
  36964=>"010011111",
  36965=>"011111101",
  36966=>"011001010",
  36967=>"110111101",
  36968=>"111000010",
  36969=>"001110010",
  36970=>"011111110",
  36971=>"111001000",
  36972=>"110111001",
  36973=>"111111111",
  36974=>"011001000",
  36975=>"000000000",
  36976=>"100111101",
  36977=>"111111010",
  36978=>"111101100",
  36979=>"000000000",
  36980=>"001100000",
  36981=>"000000000",
  36982=>"111101000",
  36983=>"000000010",
  36984=>"000000101",
  36985=>"111011111",
  36986=>"111111011",
  36987=>"111100100",
  36988=>"111100100",
  36989=>"110000000",
  36990=>"111111111",
  36991=>"001000000",
  36992=>"000000000",
  36993=>"000000000",
  36994=>"111010100",
  36995=>"110111111",
  36996=>"000010111",
  36997=>"100101001",
  36998=>"000000000",
  36999=>"000000000",
  37000=>"100001001",
  37001=>"000001001",
  37002=>"010110010",
  37003=>"000000000",
  37004=>"101000001",
  37005=>"000001011",
  37006=>"000110111",
  37007=>"000000000",
  37008=>"100010111",
  37009=>"000010111",
  37010=>"111101111",
  37011=>"000000000",
  37012=>"000000010",
  37013=>"000100111",
  37014=>"010110000",
  37015=>"000100111",
  37016=>"000000010",
  37017=>"000111111",
  37018=>"000110010",
  37019=>"000000000",
  37020=>"100111110",
  37021=>"001101000",
  37022=>"000011111",
  37023=>"101100101",
  37024=>"100110111",
  37025=>"111111111",
  37026=>"111000000",
  37027=>"111111000",
  37028=>"011110001",
  37029=>"000000000",
  37030=>"000000101",
  37031=>"100111011",
  37032=>"000110100",
  37033=>"000000001",
  37034=>"000000000",
  37035=>"000000000",
  37036=>"000000101",
  37037=>"110011001",
  37038=>"110111111",
  37039=>"011001011",
  37040=>"000000000",
  37041=>"000110010",
  37042=>"111000001",
  37043=>"111110000",
  37044=>"111111110",
  37045=>"110100000",
  37046=>"000000000",
  37047=>"000000000",
  37048=>"000000000",
  37049=>"000000000",
  37050=>"000000000",
  37051=>"000101010",
  37052=>"000100010",
  37053=>"100101101",
  37054=>"001001000",
  37055=>"111000011",
  37056=>"011011001",
  37057=>"000000000",
  37058=>"000100010",
  37059=>"011111110",
  37060=>"000000111",
  37061=>"111111111",
  37062=>"111000000",
  37063=>"101101111",
  37064=>"100100100",
  37065=>"000000011",
  37066=>"000000000",
  37067=>"011111010",
  37068=>"111000000",
  37069=>"000000001",
  37070=>"000000000",
  37071=>"000001000",
  37072=>"010111111",
  37073=>"000000100",
  37074=>"000000000",
  37075=>"111111110",
  37076=>"000000000",
  37077=>"000100000",
  37078=>"010011110",
  37079=>"111001001",
  37080=>"111111111",
  37081=>"011111010",
  37082=>"010111011",
  37083=>"000000000",
  37084=>"111111111",
  37085=>"000000000",
  37086=>"000000000",
  37087=>"111110110",
  37088=>"000000111",
  37089=>"011010010",
  37090=>"110000100",
  37091=>"000000000",
  37092=>"000000000",
  37093=>"010001100",
  37094=>"000000001",
  37095=>"011011111",
  37096=>"000000010",
  37097=>"000001000",
  37098=>"110110110",
  37099=>"000000100",
  37100=>"000111111",
  37101=>"101111000",
  37102=>"000010000",
  37103=>"001000100",
  37104=>"001000111",
  37105=>"111111111",
  37106=>"000001000",
  37107=>"111111000",
  37108=>"111011000",
  37109=>"010111111",
  37110=>"011000000",
  37111=>"000000000",
  37112=>"001000000",
  37113=>"111000010",
  37114=>"000000111",
  37115=>"100011101",
  37116=>"000000010",
  37117=>"011011000",
  37118=>"101000011",
  37119=>"011011000",
  37120=>"100100111",
  37121=>"101100001",
  37122=>"101001001",
  37123=>"111000111",
  37124=>"100100110",
  37125=>"001101011",
  37126=>"111110111",
  37127=>"011110011",
  37128=>"011011001",
  37129=>"001001101",
  37130=>"101011111",
  37131=>"001001101",
  37132=>"111000000",
  37133=>"111011001",
  37134=>"000000001",
  37135=>"111101001",
  37136=>"000000000",
  37137=>"000000110",
  37138=>"000000000",
  37139=>"111000000",
  37140=>"101101111",
  37141=>"101100111",
  37142=>"000000000",
  37143=>"000010010",
  37144=>"101000010",
  37145=>"111101111",
  37146=>"000100101",
  37147=>"000001001",
  37148=>"100101010",
  37149=>"111110100",
  37150=>"000000000",
  37151=>"110110010",
  37152=>"000000000",
  37153=>"000000101",
  37154=>"000010010",
  37155=>"101000000",
  37156=>"111110011",
  37157=>"001001111",
  37158=>"001000010",
  37159=>"000010011",
  37160=>"000111111",
  37161=>"111111111",
  37162=>"111110111",
  37163=>"001000011",
  37164=>"111100010",
  37165=>"010001010",
  37166=>"000000011",
  37167=>"111111100",
  37168=>"111101001",
  37169=>"000111111",
  37170=>"001110000",
  37171=>"101101101",
  37172=>"001111111",
  37173=>"100111111",
  37174=>"001001001",
  37175=>"111111011",
  37176=>"100001110",
  37177=>"111001000",
  37178=>"111101000",
  37179=>"000111111",
  37180=>"111011011",
  37181=>"011111111",
  37182=>"000000001",
  37183=>"000111010",
  37184=>"011101000",
  37185=>"000101111",
  37186=>"001000011",
  37187=>"100110100",
  37188=>"011000000",
  37189=>"000000100",
  37190=>"001100110",
  37191=>"011111101",
  37192=>"111011111",
  37193=>"000000001",
  37194=>"111000001",
  37195=>"111100101",
  37196=>"101001111",
  37197=>"010011101",
  37198=>"110111011",
  37199=>"001000111",
  37200=>"001001000",
  37201=>"111111111",
  37202=>"000000000",
  37203=>"001101100",
  37204=>"100000000",
  37205=>"110011011",
  37206=>"111011111",
  37207=>"100000000",
  37208=>"001111111",
  37209=>"011001001",
  37210=>"011011011",
  37211=>"000001100",
  37212=>"000000000",
  37213=>"110000101",
  37214=>"111111000",
  37215=>"001110000",
  37216=>"000010011",
  37217=>"001000011",
  37218=>"000000000",
  37219=>"101011111",
  37220=>"011001010",
  37221=>"111100100",
  37222=>"010000110",
  37223=>"111010110",
  37224=>"111100001",
  37225=>"000010110",
  37226=>"001010111",
  37227=>"011011111",
  37228=>"010001011",
  37229=>"001001001",
  37230=>"011111000",
  37231=>"101001101",
  37232=>"010010011",
  37233=>"101000010",
  37234=>"100100100",
  37235=>"010110110",
  37236=>"100111111",
  37237=>"000000111",
  37238=>"111101111",
  37239=>"000001111",
  37240=>"000000000",
  37241=>"000000000",
  37242=>"001000101",
  37243=>"111111010",
  37244=>"001000001",
  37245=>"101000001",
  37246=>"101000000",
  37247=>"001001101",
  37248=>"010001100",
  37249=>"010000011",
  37250=>"101001110",
  37251=>"111101110",
  37252=>"111111111",
  37253=>"011110100",
  37254=>"100100111",
  37255=>"010100101",
  37256=>"110010110",
  37257=>"010001001",
  37258=>"000010000",
  37259=>"011000000",
  37260=>"000000011",
  37261=>"111001001",
  37262=>"011111100",
  37263=>"000001000",
  37264=>"111100100",
  37265=>"001111111",
  37266=>"000001110",
  37267=>"111111000",
  37268=>"111101000",
  37269=>"001000000",
  37270=>"110111000",
  37271=>"010000101",
  37272=>"111010000",
  37273=>"000010001",
  37274=>"111111111",
  37275=>"000010000",
  37276=>"111101101",
  37277=>"001111100",
  37278=>"000010111",
  37279=>"011101111",
  37280=>"011111110",
  37281=>"000000100",
  37282=>"011000001",
  37283=>"001001111",
  37284=>"000000101",
  37285=>"101101011",
  37286=>"000111110",
  37287=>"000000000",
  37288=>"101000000",
  37289=>"000101000",
  37290=>"001001000",
  37291=>"000000000",
  37292=>"000111111",
  37293=>"000100101",
  37294=>"100010000",
  37295=>"000111000",
  37296=>"000100001",
  37297=>"010100000",
  37298=>"111101111",
  37299=>"100000111",
  37300=>"111011010",
  37301=>"010100000",
  37302=>"001000110",
  37303=>"111100111",
  37304=>"111100110",
  37305=>"111001101",
  37306=>"101111111",
  37307=>"111001101",
  37308=>"100110110",
  37309=>"000011011",
  37310=>"000110000",
  37311=>"000101111",
  37312=>"000000101",
  37313=>"000000010",
  37314=>"100000010",
  37315=>"011111000",
  37316=>"010110010",
  37317=>"001001000",
  37318=>"110111100",
  37319=>"001000100",
  37320=>"111011011",
  37321=>"111000111",
  37322=>"000000101",
  37323=>"000111111",
  37324=>"110111111",
  37325=>"000000100",
  37326=>"011101101",
  37327=>"101101010",
  37328=>"000010000",
  37329=>"001110011",
  37330=>"111101101",
  37331=>"111111000",
  37332=>"100010000",
  37333=>"011001100",
  37334=>"100000000",
  37335=>"110101010",
  37336=>"010110010",
  37337=>"000110000",
  37338=>"001101000",
  37339=>"000000001",
  37340=>"110110010",
  37341=>"100000010",
  37342=>"110110111",
  37343=>"100000000",
  37344=>"000000000",
  37345=>"000000100",
  37346=>"110110110",
  37347=>"000000000",
  37348=>"101000001",
  37349=>"000101111",
  37350=>"101001000",
  37351=>"111110001",
  37352=>"111010110",
  37353=>"101000111",
  37354=>"110110110",
  37355=>"101000101",
  37356=>"000000000",
  37357=>"000110001",
  37358=>"111000110",
  37359=>"010111010",
  37360=>"111111110",
  37361=>"101000110",
  37362=>"000000001",
  37363=>"111101001",
  37364=>"010000110",
  37365=>"000000011",
  37366=>"101000110",
  37367=>"100111111",
  37368=>"000000111",
  37369=>"110110111",
  37370=>"101100111",
  37371=>"011001000",
  37372=>"111011000",
  37373=>"000000100",
  37374=>"101111001",
  37375=>"000000010",
  37376=>"001001100",
  37377=>"000001010",
  37378=>"110010000",
  37379=>"111101101",
  37380=>"111011111",
  37381=>"001000111",
  37382=>"111111010",
  37383=>"010001111",
  37384=>"101001010",
  37385=>"000000000",
  37386=>"011110010",
  37387=>"000000001",
  37388=>"000000101",
  37389=>"100000101",
  37390=>"000001011",
  37391=>"110001101",
  37392=>"000101111",
  37393=>"100111111",
  37394=>"101110000",
  37395=>"110111011",
  37396=>"111111110",
  37397=>"000000000",
  37398=>"110110001",
  37399=>"001110110",
  37400=>"100000101",
  37401=>"000000001",
  37402=>"000000100",
  37403=>"001111111",
  37404=>"101101000",
  37405=>"011000000",
  37406=>"000000101",
  37407=>"010000000",
  37408=>"111111101",
  37409=>"000100111",
  37410=>"111111010",
  37411=>"000111110",
  37412=>"111001011",
  37413=>"100001000",
  37414=>"110110111",
  37415=>"000000000",
  37416=>"111010000",
  37417=>"101000001",
  37418=>"100110111",
  37419=>"000000000",
  37420=>"111111110",
  37421=>"001111000",
  37422=>"000110100",
  37423=>"110000000",
  37424=>"111111001",
  37425=>"001111111",
  37426=>"111011001",
  37427=>"000011010",
  37428=>"000111011",
  37429=>"000000000",
  37430=>"000001111",
  37431=>"011000110",
  37432=>"110111111",
  37433=>"000111010",
  37434=>"001000000",
  37435=>"100000000",
  37436=>"000001001",
  37437=>"010010010",
  37438=>"000100100",
  37439=>"110001100",
  37440=>"011010101",
  37441=>"101000000",
  37442=>"000000110",
  37443=>"011011001",
  37444=>"111000111",
  37445=>"111100000",
  37446=>"111000000",
  37447=>"111101100",
  37448=>"101011011",
  37449=>"101101111",
  37450=>"101001011",
  37451=>"000010111",
  37452=>"000000001",
  37453=>"101111111",
  37454=>"000010111",
  37455=>"111100111",
  37456=>"000100000",
  37457=>"111111010",
  37458=>"000111101",
  37459=>"011000110",
  37460=>"000000111",
  37461=>"100100000",
  37462=>"111011000",
  37463=>"000000111",
  37464=>"000000111",
  37465=>"001000001",
  37466=>"011000001",
  37467=>"001111100",
  37468=>"111111010",
  37469=>"110000001",
  37470=>"010111111",
  37471=>"110100000",
  37472=>"011101111",
  37473=>"001000100",
  37474=>"001111111",
  37475=>"100000000",
  37476=>"000000001",
  37477=>"000111000",
  37478=>"111000000",
  37479=>"111101100",
  37480=>"010000100",
  37481=>"111010000",
  37482=>"111011111",
  37483=>"111000111",
  37484=>"111110110",
  37485=>"111111110",
  37486=>"111000000",
  37487=>"000100010",
  37488=>"101110111",
  37489=>"111000111",
  37490=>"001110111",
  37491=>"111111100",
  37492=>"111000000",
  37493=>"000000101",
  37494=>"001000111",
  37495=>"000001100",
  37496=>"111001000",
  37497=>"010000110",
  37498=>"111111010",
  37499=>"110000000",
  37500=>"011101110",
  37501=>"110000001",
  37502=>"111111000",
  37503=>"000001101",
  37504=>"100010000",
  37505=>"000000000",
  37506=>"101011000",
  37507=>"011111000",
  37508=>"010111111",
  37509=>"011010000",
  37510=>"001000000",
  37511=>"000000000",
  37512=>"000101111",
  37513=>"000000000",
  37514=>"011111101",
  37515=>"110111001",
  37516=>"000010000",
  37517=>"010001000",
  37518=>"111000000",
  37519=>"000001101",
  37520=>"101111011",
  37521=>"000000110",
  37522=>"101100001",
  37523=>"100111111",
  37524=>"011111101",
  37525=>"100000111",
  37526=>"000001000",
  37527=>"100000000",
  37528=>"010000000",
  37529=>"110111111",
  37530=>"110110101",
  37531=>"011001000",
  37532=>"110000110",
  37533=>"000000111",
  37534=>"000111010",
  37535=>"000000000",
  37536=>"111001000",
  37537=>"000000010",
  37538=>"010000001",
  37539=>"100000011",
  37540=>"111010011",
  37541=>"100000000",
  37542=>"111010000",
  37543=>"000010010",
  37544=>"001000111",
  37545=>"000110000",
  37546=>"000000000",
  37547=>"000111111",
  37548=>"111011100",
  37549=>"001101001",
  37550=>"000000001",
  37551=>"111011011",
  37552=>"010000000",
  37553=>"000001010",
  37554=>"111000000",
  37555=>"101000100",
  37556=>"111011110",
  37557=>"111111100",
  37558=>"010111111",
  37559=>"001000000",
  37560=>"000101010",
  37561=>"100100101",
  37562=>"000000111",
  37563=>"111000000",
  37564=>"001010000",
  37565=>"111011111",
  37566=>"000100001",
  37567=>"101110011",
  37568=>"100000010",
  37569=>"000111010",
  37570=>"101101111",
  37571=>"011101100",
  37572=>"111110000",
  37573=>"100100110",
  37574=>"111110110",
  37575=>"000000000",
  37576=>"111111001",
  37577=>"101111101",
  37578=>"111111110",
  37579=>"111001000",
  37580=>"111000100",
  37581=>"100101011",
  37582=>"000111011",
  37583=>"011111110",
  37584=>"000111111",
  37585=>"000001111",
  37586=>"000101111",
  37587=>"010000000",
  37588=>"000000111",
  37589=>"101000010",
  37590=>"000000111",
  37591=>"110100111",
  37592=>"111000000",
  37593=>"011111111",
  37594=>"010110000",
  37595=>"111010000",
  37596=>"011111100",
  37597=>"110110000",
  37598=>"001001100",
  37599=>"000100111",
  37600=>"101110111",
  37601=>"111010011",
  37602=>"010000101",
  37603=>"000111110",
  37604=>"110100101",
  37605=>"110100111",
  37606=>"000111111",
  37607=>"010111100",
  37608=>"001001100",
  37609=>"110000001",
  37610=>"100100100",
  37611=>"000100111",
  37612=>"000000110",
  37613=>"000000001",
  37614=>"000000010",
  37615=>"111000000",
  37616=>"000000001",
  37617=>"001011001",
  37618=>"010011000",
  37619=>"110011011",
  37620=>"100111111",
  37621=>"010000011",
  37622=>"000010111",
  37623=>"111011000",
  37624=>"001111000",
  37625=>"111000000",
  37626=>"111001001",
  37627=>"000001111",
  37628=>"111111000",
  37629=>"111111111",
  37630=>"000001100",
  37631=>"101101110",
  37632=>"001110100",
  37633=>"100111010",
  37634=>"111000101",
  37635=>"001111111",
  37636=>"000000100",
  37637=>"000010000",
  37638=>"000101110",
  37639=>"010010100",
  37640=>"100001111",
  37641=>"111100000",
  37642=>"011011000",
  37643=>"011011001",
  37644=>"010011001",
  37645=>"000000111",
  37646=>"011011000",
  37647=>"001000000",
  37648=>"000100100",
  37649=>"100111010",
  37650=>"001000010",
  37651=>"000000000",
  37652=>"111000011",
  37653=>"001000000",
  37654=>"101011100",
  37655=>"001111110",
  37656=>"100101100",
  37657=>"001101101",
  37658=>"000111111",
  37659=>"011011000",
  37660=>"101111011",
  37661=>"100100000",
  37662=>"111111100",
  37663=>"000011111",
  37664=>"010000110",
  37665=>"000100111",
  37666=>"111000100",
  37667=>"111111001",
  37668=>"111001110",
  37669=>"010000000",
  37670=>"100000000",
  37671=>"111011001",
  37672=>"011011000",
  37673=>"101101111",
  37674=>"000110111",
  37675=>"000000000",
  37676=>"100111110",
  37677=>"000111011",
  37678=>"011010000",
  37679=>"110100001",
  37680=>"111111110",
  37681=>"011011011",
  37682=>"100100111",
  37683=>"110111111",
  37684=>"011011000",
  37685=>"000000000",
  37686=>"001001010",
  37687=>"000101111",
  37688=>"110100001",
  37689=>"000000111",
  37690=>"000100100",
  37691=>"111111010",
  37692=>"111111001",
  37693=>"111111001",
  37694=>"011000000",
  37695=>"111111100",
  37696=>"000010101",
  37697=>"001111111",
  37698=>"000110110",
  37699=>"111110100",
  37700=>"000100101",
  37701=>"100001101",
  37702=>"010000100",
  37703=>"100100111",
  37704=>"001001111",
  37705=>"011010000",
  37706=>"101100101",
  37707=>"100101111",
  37708=>"100100111",
  37709=>"010110110",
  37710=>"111111000",
  37711=>"000000100",
  37712=>"111100000",
  37713=>"101100111",
  37714=>"000100101",
  37715=>"011110000",
  37716=>"011011000",
  37717=>"101111000",
  37718=>"111110000",
  37719=>"111010000",
  37720=>"110000100",
  37721=>"101111001",
  37722=>"111100011",
  37723=>"011011011",
  37724=>"000111101",
  37725=>"001001011",
  37726=>"101100111",
  37727=>"111000100",
  37728=>"001111111",
  37729=>"111111000",
  37730=>"010100100",
  37731=>"111011110",
  37732=>"000000000",
  37733=>"001000011",
  37734=>"001011000",
  37735=>"000100110",
  37736=>"101100000",
  37737=>"010111111",
  37738=>"000000111",
  37739=>"000000101",
  37740=>"100000111",
  37741=>"110100010",
  37742=>"111100110",
  37743=>"111011011",
  37744=>"110110010",
  37745=>"000000000",
  37746=>"100111011",
  37747=>"110111110",
  37748=>"001101000",
  37749=>"000100111",
  37750=>"111111000",
  37751=>"000000001",
  37752=>"111110111",
  37753=>"000111111",
  37754=>"000010010",
  37755=>"000000100",
  37756=>"110010010",
  37757=>"110111100",
  37758=>"000000100",
  37759=>"111010000",
  37760=>"101111010",
  37761=>"100011100",
  37762=>"100101000",
  37763=>"100111111",
  37764=>"011001000",
  37765=>"110000111",
  37766=>"010100101",
  37767=>"010010000",
  37768=>"111011000",
  37769=>"000000000",
  37770=>"111110011",
  37771=>"000000000",
  37772=>"111111000",
  37773=>"110000000",
  37774=>"011011111",
  37775=>"110000010",
  37776=>"110110100",
  37777=>"000010111",
  37778=>"100000000",
  37779=>"011111001",
  37780=>"011011000",
  37781=>"010000101",
  37782=>"000111111",
  37783=>"100100111",
  37784=>"100111011",
  37785=>"101011111",
  37786=>"000100111",
  37787=>"100100101",
  37788=>"000000111",
  37789=>"000100010",
  37790=>"110111111",
  37791=>"100000100",
  37792=>"100110111",
  37793=>"000000000",
  37794=>"000000111",
  37795=>"100000101",
  37796=>"000010001",
  37797=>"010110100",
  37798=>"100101011",
  37799=>"000100111",
  37800=>"000111111",
  37801=>"110000010",
  37802=>"111100000",
  37803=>"010100000",
  37804=>"100100111",
  37805=>"011010000",
  37806=>"111101000",
  37807=>"010000001",
  37808=>"100110101",
  37809=>"001110111",
  37810=>"100101010",
  37811=>"000010100",
  37812=>"001001000",
  37813=>"101111010",
  37814=>"100100100",
  37815=>"000000000",
  37816=>"111011011",
  37817=>"110110100",
  37818=>"010101000",
  37819=>"100010111",
  37820=>"000001101",
  37821=>"110100000",
  37822=>"101111011",
  37823=>"000011100",
  37824=>"000100100",
  37825=>"000101010",
  37826=>"111111111",
  37827=>"110110000",
  37828=>"011000000",
  37829=>"101001011",
  37830=>"000010111",
  37831=>"011000110",
  37832=>"000000100",
  37833=>"100101110",
  37834=>"000100101",
  37835=>"111100000",
  37836=>"000000110",
  37837=>"011011100",
  37838=>"011011011",
  37839=>"111111111",
  37840=>"100100111",
  37841=>"001011110",
  37842=>"010000111",
  37843=>"100101110",
  37844=>"011000000",
  37845=>"111001110",
  37846=>"100100111",
  37847=>"000011110",
  37848=>"000000011",
  37849=>"100100100",
  37850=>"001101101",
  37851=>"110000000",
  37852=>"110100100",
  37853=>"100000011",
  37854=>"000111010",
  37855=>"111011111",
  37856=>"000001111",
  37857=>"011011100",
  37858=>"011011010",
  37859=>"110110000",
  37860=>"101110000",
  37861=>"100100000",
  37862=>"000100101",
  37863=>"110110111",
  37864=>"111011010",
  37865=>"010100111",
  37866=>"111110000",
  37867=>"111111100",
  37868=>"010010000",
  37869=>"011010000",
  37870=>"010010000",
  37871=>"000110011",
  37872=>"101001000",
  37873=>"001001101",
  37874=>"100111100",
  37875=>"100100110",
  37876=>"100111011",
  37877=>"010101110",
  37878=>"011100000",
  37879=>"110011110",
  37880=>"000000100",
  37881=>"110100100",
  37882=>"000001001",
  37883=>"100101010",
  37884=>"101011010",
  37885=>"011000000",
  37886=>"001011000",
  37887=>"011000000",
  37888=>"010011001",
  37889=>"001010000",
  37890=>"111100100",
  37891=>"011001010",
  37892=>"100110110",
  37893=>"010000011",
  37894=>"000101111",
  37895=>"100111110",
  37896=>"101000100",
  37897=>"000000111",
  37898=>"000110010",
  37899=>"100010011",
  37900=>"111100100",
  37901=>"000101011",
  37902=>"101111001",
  37903=>"001111111",
  37904=>"000010010",
  37905=>"000011010",
  37906=>"011000000",
  37907=>"000000011",
  37908=>"111100101",
  37909=>"001000000",
  37910=>"111000000",
  37911=>"110010111",
  37912=>"010010100",
  37913=>"001000111",
  37914=>"111100000",
  37915=>"000100000",
  37916=>"000000000",
  37917=>"100101011",
  37918=>"000010011",
  37919=>"111000011",
  37920=>"011101100",
  37921=>"111100000",
  37922=>"011111100",
  37923=>"101101001",
  37924=>"010110110",
  37925=>"000110100",
  37926=>"110100100",
  37927=>"001110111",
  37928=>"000010100",
  37929=>"010011011",
  37930=>"000011111",
  37931=>"101111110",
  37932=>"011111100",
  37933=>"111111111",
  37934=>"010010111",
  37935=>"111111011",
  37936=>"111111101",
  37937=>"111111111",
  37938=>"111000001",
  37939=>"111010011",
  37940=>"000110111",
  37941=>"011011001",
  37942=>"000000010",
  37943=>"000010000",
  37944=>"000000011",
  37945=>"001111011",
  37946=>"000011010",
  37947=>"000111000",
  37948=>"000110110",
  37949=>"011101110",
  37950=>"010000000",
  37951=>"110110101",
  37952=>"010000000",
  37953=>"111111000",
  37954=>"111000100",
  37955=>"111100111",
  37956=>"111101101",
  37957=>"000000101",
  37958=>"000111101",
  37959=>"000010000",
  37960=>"110111001",
  37961=>"000111011",
  37962=>"111001111",
  37963=>"000010010",
  37964=>"111000001",
  37965=>"111011011",
  37966=>"010111111",
  37967=>"111111000",
  37968=>"011001011",
  37969=>"011111111",
  37970=>"111011000",
  37971=>"011001000",
  37972=>"000010010",
  37973=>"000111011",
  37974=>"011011001",
  37975=>"000100101",
  37976=>"100001011",
  37977=>"011111011",
  37978=>"101110111",
  37979=>"000001111",
  37980=>"111000000",
  37981=>"101000000",
  37982=>"101111011",
  37983=>"001001001",
  37984=>"111111001",
  37985=>"110111011",
  37986=>"110100101",
  37987=>"010100000",
  37988=>"000101111",
  37989=>"100111111",
  37990=>"111111111",
  37991=>"101100101",
  37992=>"111011110",
  37993=>"000010110",
  37994=>"000000000",
  37995=>"011010001",
  37996=>"111111001",
  37997=>"100111111",
  37998=>"011101100",
  37999=>"100110111",
  38000=>"001001101",
  38001=>"101111111",
  38002=>"000001011",
  38003=>"101100100",
  38004=>"000101111",
  38005=>"000000101",
  38006=>"011100111",
  38007=>"111111111",
  38008=>"010111000",
  38009=>"000000100",
  38010=>"001000100",
  38011=>"111111101",
  38012=>"000110010",
  38013=>"111100000",
  38014=>"111101101",
  38015=>"101000111",
  38016=>"110000000",
  38017=>"010000000",
  38018=>"000111010",
  38019=>"000000110",
  38020=>"100101000",
  38021=>"000101000",
  38022=>"100011111",
  38023=>"100000011",
  38024=>"111101111",
  38025=>"101011101",
  38026=>"000001001",
  38027=>"100000111",
  38028=>"111100101",
  38029=>"000000000",
  38030=>"000011111",
  38031=>"100001001",
  38032=>"011111111",
  38033=>"111011011",
  38034=>"000011100",
  38035=>"000000000",
  38036=>"000000000",
  38037=>"000000100",
  38038=>"000010011",
  38039=>"110110100",
  38040=>"101000010",
  38041=>"111111000",
  38042=>"000111011",
  38043=>"000000100",
  38044=>"101000000",
  38045=>"001010010",
  38046=>"001100011",
  38047=>"111101000",
  38048=>"110101011",
  38049=>"111011011",
  38050=>"010000101",
  38051=>"111000000",
  38052=>"011110100",
  38053=>"100100111",
  38054=>"001001001",
  38055=>"000000000",
  38056=>"000000000",
  38057=>"111001000",
  38058=>"011101101",
  38059=>"000000010",
  38060=>"000010000",
  38061=>"110000000",
  38062=>"011111100",
  38063=>"111001000",
  38064=>"011011000",
  38065=>"001000110",
  38066=>"100011111",
  38067=>"001000000",
  38068=>"000110111",
  38069=>"010010111",
  38070=>"111111110",
  38071=>"001010010",
  38072=>"000011111",
  38073=>"000000011",
  38074=>"000110111",
  38075=>"111111010",
  38076=>"000000111",
  38077=>"110111111",
  38078=>"001001000",
  38079=>"111000000",
  38080=>"000010010",
  38081=>"000110111",
  38082=>"111110101",
  38083=>"001110110",
  38084=>"000111101",
  38085=>"010110101",
  38086=>"111111100",
  38087=>"000101100",
  38088=>"101110111",
  38089=>"111101000",
  38090=>"111101000",
  38091=>"111111111",
  38092=>"000010010",
  38093=>"000001010",
  38094=>"010010010",
  38095=>"111100100",
  38096=>"000011111",
  38097=>"011111001",
  38098=>"101000000",
  38099=>"000111011",
  38100=>"101000100",
  38101=>"100000000",
  38102=>"111100000",
  38103=>"000111111",
  38104=>"010011000",
  38105=>"101000000",
  38106=>"000001000",
  38107=>"111000111",
  38108=>"011100100",
  38109=>"111100000",
  38110=>"000011111",
  38111=>"000010110",
  38112=>"111100000",
  38113=>"011101101",
  38114=>"000111111",
  38115=>"110100101",
  38116=>"101000000",
  38117=>"000000000",
  38118=>"010000000",
  38119=>"110001000",
  38120=>"111111100",
  38121=>"011111110",
  38122=>"000111011",
  38123=>"010111101",
  38124=>"111100000",
  38125=>"101111110",
  38126=>"010000000",
  38127=>"000000011",
  38128=>"000100111",
  38129=>"100011001",
  38130=>"010000000",
  38131=>"110011001",
  38132=>"000110011",
  38133=>"110111111",
  38134=>"000000010",
  38135=>"011101100",
  38136=>"000111000",
  38137=>"111111111",
  38138=>"010100101",
  38139=>"010001101",
  38140=>"000010010",
  38141=>"000000000",
  38142=>"011000101",
  38143=>"111111000",
  38144=>"011011100",
  38145=>"111110010",
  38146=>"000000010",
  38147=>"000010111",
  38148=>"010001001",
  38149=>"000100000",
  38150=>"000111111",
  38151=>"111111011",
  38152=>"000000101",
  38153=>"111011111",
  38154=>"100100100",
  38155=>"100101000",
  38156=>"111000000",
  38157=>"000000111",
  38158=>"100001100",
  38159=>"000101010",
  38160=>"000111011",
  38161=>"000001000",
  38162=>"101000010",
  38163=>"011010000",
  38164=>"000011111",
  38165=>"000010010",
  38166=>"011011111",
  38167=>"000010111",
  38168=>"101010010",
  38169=>"101111111",
  38170=>"000110100",
  38171=>"111010110",
  38172=>"101101000",
  38173=>"110000000",
  38174=>"001001010",
  38175=>"001001000",
  38176=>"000000010",
  38177=>"101101110",
  38178=>"010000000",
  38179=>"111111011",
  38180=>"001001000",
  38181=>"001101000",
  38182=>"010010100",
  38183=>"010010101",
  38184=>"111101101",
  38185=>"010000001",
  38186=>"101001111",
  38187=>"010000010",
  38188=>"110100000",
  38189=>"011010000",
  38190=>"000000110",
  38191=>"110110001",
  38192=>"000101111",
  38193=>"101101100",
  38194=>"100100001",
  38195=>"000110111",
  38196=>"111000000",
  38197=>"011010111",
  38198=>"111110010",
  38199=>"010000101",
  38200=>"111001001",
  38201=>"000111000",
  38202=>"000000010",
  38203=>"001110010",
  38204=>"110111010",
  38205=>"011101000",
  38206=>"000001100",
  38207=>"011011011",
  38208=>"111011000",
  38209=>"001101100",
  38210=>"001111001",
  38211=>"011001000",
  38212=>"000001000",
  38213=>"000001000",
  38214=>"010110000",
  38215=>"010000100",
  38216=>"111110001",
  38217=>"111111111",
  38218=>"000000000",
  38219=>"101110111",
  38220=>"000010111",
  38221=>"100100100",
  38222=>"011001001",
  38223=>"000000001",
  38224=>"111100000",
  38225=>"000000111",
  38226=>"101101010",
  38227=>"001000010",
  38228=>"111111101",
  38229=>"011111110",
  38230=>"100101100",
  38231=>"000010000",
  38232=>"111111111",
  38233=>"011100100",
  38234=>"111100000",
  38235=>"110101111",
  38236=>"000011011",
  38237=>"000000010",
  38238=>"000011111",
  38239=>"110100100",
  38240=>"111100000",
  38241=>"101000000",
  38242=>"000000111",
  38243=>"001001100",
  38244=>"100100000",
  38245=>"111001001",
  38246=>"100111000",
  38247=>"000001101",
  38248=>"111010011",
  38249=>"111000111",
  38250=>"000000111",
  38251=>"000111111",
  38252=>"110000000",
  38253=>"000000111",
  38254=>"100110111",
  38255=>"101000100",
  38256=>"111101010",
  38257=>"000111111",
  38258=>"111011010",
  38259=>"101000000",
  38260=>"100000000",
  38261=>"000100100",
  38262=>"000011111",
  38263=>"000000100",
  38264=>"000010111",
  38265=>"111011111",
  38266=>"100100101",
  38267=>"011001101",
  38268=>"001001011",
  38269=>"110100010",
  38270=>"111100001",
  38271=>"101101101",
  38272=>"010111111",
  38273=>"100000000",
  38274=>"000000011",
  38275=>"000000011",
  38276=>"100111010",
  38277=>"111101111",
  38278=>"100100000",
  38279=>"000001001",
  38280=>"111100100",
  38281=>"000000000",
  38282=>"100110011",
  38283=>"110010010",
  38284=>"010110101",
  38285=>"000101100",
  38286=>"011101000",
  38287=>"100100100",
  38288=>"101101100",
  38289=>"011111000",
  38290=>"101111111",
  38291=>"110000101",
  38292=>"000001101",
  38293=>"000010111",
  38294=>"010111011",
  38295=>"010011110",
  38296=>"111111100",
  38297=>"010111111",
  38298=>"111101111",
  38299=>"001000000",
  38300=>"000000000",
  38301=>"111111000",
  38302=>"111111111",
  38303=>"111111100",
  38304=>"111001001",
  38305=>"111111111",
  38306=>"000000000",
  38307=>"011101101",
  38308=>"001110111",
  38309=>"011001000",
  38310=>"101000101",
  38311=>"011111100",
  38312=>"100000111",
  38313=>"011000000",
  38314=>"101101111",
  38315=>"101010010",
  38316=>"111000010",
  38317=>"111001100",
  38318=>"110100000",
  38319=>"111111101",
  38320=>"111110000",
  38321=>"001101100",
  38322=>"010000111",
  38323=>"011000000",
  38324=>"011111110",
  38325=>"100100000",
  38326=>"111011111",
  38327=>"101110010",
  38328=>"001011010",
  38329=>"000000111",
  38330=>"011010000",
  38331=>"100100111",
  38332=>"111100000",
  38333=>"100111111",
  38334=>"010010110",
  38335=>"111000000",
  38336=>"101111111",
  38337=>"000010010",
  38338=>"000110010",
  38339=>"011001000",
  38340=>"000011111",
  38341=>"011001001",
  38342=>"111011011",
  38343=>"000000110",
  38344=>"000111111",
  38345=>"010010110",
  38346=>"010011011",
  38347=>"100100000",
  38348=>"001100000",
  38349=>"000100110",
  38350=>"101000000",
  38351=>"010010000",
  38352=>"001000000",
  38353=>"111101001",
  38354=>"000000101",
  38355=>"001000000",
  38356=>"110101101",
  38357=>"110100000",
  38358=>"000010010",
  38359=>"010011010",
  38360=>"011111000",
  38361=>"010000000",
  38362=>"110101100",
  38363=>"100000110",
  38364=>"111110111",
  38365=>"111111111",
  38366=>"111111101",
  38367=>"000000001",
  38368=>"000000111",
  38369=>"000000111",
  38370=>"111111001",
  38371=>"001001001",
  38372=>"000010110",
  38373=>"010100000",
  38374=>"101000000",
  38375=>"111011001",
  38376=>"110000000",
  38377=>"111001010",
  38378=>"001001000",
  38379=>"101110111",
  38380=>"000000000",
  38381=>"000111111",
  38382=>"000000000",
  38383=>"100010000",
  38384=>"111000000",
  38385=>"000100000",
  38386=>"001000111",
  38387=>"111001011",
  38388=>"110110000",
  38389=>"101000000",
  38390=>"000000010",
  38391=>"101111101",
  38392=>"000110101",
  38393=>"000001010",
  38394=>"111001110",
  38395=>"010000100",
  38396=>"010000000",
  38397=>"000111111",
  38398=>"110100000",
  38399=>"010010000",
  38400=>"001000100",
  38401=>"000011000",
  38402=>"000000101",
  38403=>"101110100",
  38404=>"111111011",
  38405=>"001000011",
  38406=>"000000110",
  38407=>"000101000",
  38408=>"111111010",
  38409=>"111110100",
  38410=>"111110111",
  38411=>"000000100",
  38412=>"000000000",
  38413=>"101111111",
  38414=>"011011000",
  38415=>"001001101",
  38416=>"111101011",
  38417=>"110000000",
  38418=>"000000000",
  38419=>"010000001",
  38420=>"111111010",
  38421=>"111110000",
  38422=>"111001000",
  38423=>"000111000",
  38424=>"000000111",
  38425=>"000000000",
  38426=>"100100000",
  38427=>"110111111",
  38428=>"100000000",
  38429=>"000000101",
  38430=>"000000111",
  38431=>"010000001",
  38432=>"000000010",
  38433=>"111111010",
  38434=>"111101010",
  38435=>"011111111",
  38436=>"010110111",
  38437=>"011011011",
  38438=>"110000000",
  38439=>"111111001",
  38440=>"110111100",
  38441=>"111111111",
  38442=>"100000001",
  38443=>"101111111",
  38444=>"000000001",
  38445=>"111100000",
  38446=>"000100100",
  38447=>"101111010",
  38448=>"000111000",
  38449=>"000100100",
  38450=>"000111110",
  38451=>"010110100",
  38452=>"010000000",
  38453=>"000000000",
  38454=>"111111000",
  38455=>"000000101",
  38456=>"111111111",
  38457=>"000000000",
  38458=>"000000111",
  38459=>"110000010",
  38460=>"000000000",
  38461=>"111111011",
  38462=>"100001111",
  38463=>"111111100",
  38464=>"001111111",
  38465=>"000011000",
  38466=>"000100000",
  38467=>"011111011",
  38468=>"111001111",
  38469=>"000000000",
  38470=>"111111110",
  38471=>"111111111",
  38472=>"110110010",
  38473=>"000000001",
  38474=>"000000000",
  38475=>"101100000",
  38476=>"000000011",
  38477=>"111111110",
  38478=>"000011001",
  38479=>"000000000",
  38480=>"111111000",
  38481=>"111111111",
  38482=>"111011111",
  38483=>"001100111",
  38484=>"000000000",
  38485=>"111110000",
  38486=>"111011000",
  38487=>"001000011",
  38488=>"011100000",
  38489=>"000100100",
  38490=>"011011000",
  38491=>"111111111",
  38492=>"010111111",
  38493=>"011001100",
  38494=>"111111000",
  38495=>"111110110",
  38496=>"111111111",
  38497=>"111111100",
  38498=>"101000111",
  38499=>"100000001",
  38500=>"101101000",
  38501=>"010000101",
  38502=>"000000111",
  38503=>"111001111",
  38504=>"101010101",
  38505=>"111111111",
  38506=>"100000010",
  38507=>"001111000",
  38508=>"111111111",
  38509=>"110000110",
  38510=>"101101111",
  38511=>"000000111",
  38512=>"011001011",
  38513=>"111111111",
  38514=>"111111000",
  38515=>"111000001",
  38516=>"000000110",
  38517=>"000001111",
  38518=>"101000111",
  38519=>"111111111",
  38520=>"000000101",
  38521=>"111001101",
  38522=>"101100001",
  38523=>"111111000",
  38524=>"111010100",
  38525=>"100001110",
  38526=>"110111111",
  38527=>"001001001",
  38528=>"000111111",
  38529=>"000000101",
  38530=>"111111111",
  38531=>"101101111",
  38532=>"000000000",
  38533=>"111111010",
  38534=>"100110000",
  38535=>"110110110",
  38536=>"110110000",
  38537=>"110111100",
  38538=>"111111110",
  38539=>"001110001",
  38540=>"000000010",
  38541=>"000101000",
  38542=>"001001000",
  38543=>"011110000",
  38544=>"001001111",
  38545=>"101111111",
  38546=>"000000000",
  38547=>"000000000",
  38548=>"111011000",
  38549=>"010110000",
  38550=>"111111111",
  38551=>"001011011",
  38552=>"000000000",
  38553=>"011010001",
  38554=>"101111011",
  38555=>"000000000",
  38556=>"101110011",
  38557=>"010111111",
  38558=>"111111000",
  38559=>"000000000",
  38560=>"001101011",
  38561=>"000000111",
  38562=>"000101011",
  38563=>"000010000",
  38564=>"111111011",
  38565=>"001011011",
  38566=>"110100000",
  38567=>"001001111",
  38568=>"111001010",
  38569=>"111111111",
  38570=>"111111110",
  38571=>"000001000",
  38572=>"101101110",
  38573=>"000000111",
  38574=>"100100111",
  38575=>"111111110",
  38576=>"000000100",
  38577=>"011010011",
  38578=>"000000000",
  38579=>"100010001",
  38580=>"001000000",
  38581=>"111111111",
  38582=>"000000111",
  38583=>"100000000",
  38584=>"100000100",
  38585=>"011101000",
  38586=>"001111111",
  38587=>"001000000",
  38588=>"000000000",
  38589=>"000000000",
  38590=>"110110010",
  38591=>"010000101",
  38592=>"000010000",
  38593=>"000000000",
  38594=>"011111110",
  38595=>"000000000",
  38596=>"000000111",
  38597=>"111001000",
  38598=>"000001111",
  38599=>"111110000",
  38600=>"000101001",
  38601=>"000000000",
  38602=>"100110111",
  38603=>"000000010",
  38604=>"000000000",
  38605=>"111100000",
  38606=>"000100101",
  38607=>"111111000",
  38608=>"110011010",
  38609=>"110111111",
  38610=>"000000001",
  38611=>"000000000",
  38612=>"000000100",
  38613=>"100000000",
  38614=>"111111111",
  38615=>"001111111",
  38616=>"000000001",
  38617=>"111000000",
  38618=>"000001110",
  38619=>"000000111",
  38620=>"111110010",
  38621=>"111111000",
  38622=>"000001101",
  38623=>"111111000",
  38624=>"010010001",
  38625=>"100110000",
  38626=>"010000000",
  38627=>"111111000",
  38628=>"001000001",
  38629=>"100111111",
  38630=>"101101010",
  38631=>"000010010",
  38632=>"001000101",
  38633=>"100101000",
  38634=>"111111110",
  38635=>"001111100",
  38636=>"010010000",
  38637=>"000000101",
  38638=>"111111000",
  38639=>"111101000",
  38640=>"000000001",
  38641=>"111000100",
  38642=>"111111110",
  38643=>"000001000",
  38644=>"001011011",
  38645=>"111110000",
  38646=>"100101111",
  38647=>"000000000",
  38648=>"000111111",
  38649=>"000100000",
  38650=>"110000000",
  38651=>"110000000",
  38652=>"000001000",
  38653=>"000000011",
  38654=>"111111110",
  38655=>"000000100",
  38656=>"000000100",
  38657=>"000011111",
  38658=>"000000110",
  38659=>"111111011",
  38660=>"100001001",
  38661=>"111100111",
  38662=>"101101111",
  38663=>"000111111",
  38664=>"001001001",
  38665=>"000001010",
  38666=>"100100000",
  38667=>"110110111",
  38668=>"111110010",
  38669=>"000000001",
  38670=>"000010000",
  38671=>"000100110",
  38672=>"000110111",
  38673=>"100011100",
  38674=>"111101011",
  38675=>"010000001",
  38676=>"000000110",
  38677=>"000101111",
  38678=>"000000000",
  38679=>"111111111",
  38680=>"111010010",
  38681=>"010000101",
  38682=>"111001000",
  38683=>"100111000",
  38684=>"100111110",
  38685=>"101100000",
  38686=>"000000111",
  38687=>"000000000",
  38688=>"000010010",
  38689=>"000001111",
  38690=>"111000110",
  38691=>"001111111",
  38692=>"010000110",
  38693=>"001000000",
  38694=>"011111111",
  38695=>"101000111",
  38696=>"001001000",
  38697=>"000111111",
  38698=>"000000000",
  38699=>"110111110",
  38700=>"000011000",
  38701=>"100111001",
  38702=>"111110111",
  38703=>"000000011",
  38704=>"000000000",
  38705=>"000000000",
  38706=>"000000110",
  38707=>"000000011",
  38708=>"011000001",
  38709=>"010111111",
  38710=>"011011000",
  38711=>"000000001",
  38712=>"111100010",
  38713=>"000101000",
  38714=>"010010010",
  38715=>"111010001",
  38716=>"010000000",
  38717=>"111000111",
  38718=>"010000001",
  38719=>"011001000",
  38720=>"111110111",
  38721=>"001111010",
  38722=>"000001010",
  38723=>"111011000",
  38724=>"000000001",
  38725=>"000000000",
  38726=>"010011011",
  38727=>"101100111",
  38728=>"001110110",
  38729=>"010101011",
  38730=>"000000000",
  38731=>"001001101",
  38732=>"110111100",
  38733=>"100100100",
  38734=>"001001001",
  38735=>"011001011",
  38736=>"000001001",
  38737=>"111111111",
  38738=>"111111111",
  38739=>"000010011",
  38740=>"001001101",
  38741=>"011000000",
  38742=>"010001000",
  38743=>"000000111",
  38744=>"010001001",
  38745=>"110110011",
  38746=>"000100100",
  38747=>"111010110",
  38748=>"101001001",
  38749=>"000000100",
  38750=>"111111111",
  38751=>"000000010",
  38752=>"010111001",
  38753=>"000001000",
  38754=>"111110000",
  38755=>"110111111",
  38756=>"010001000",
  38757=>"110000000",
  38758=>"000001100",
  38759=>"101111111",
  38760=>"000000000",
  38761=>"000000111",
  38762=>"000000000",
  38763=>"001101111",
  38764=>"000000000",
  38765=>"000001111",
  38766=>"011001001",
  38767=>"000000010",
  38768=>"111011000",
  38769=>"000010010",
  38770=>"110100000",
  38771=>"000110011",
  38772=>"111110000",
  38773=>"010010000",
  38774=>"000000001",
  38775=>"001010000",
  38776=>"111111100",
  38777=>"110111111",
  38778=>"000000000",
  38779=>"111111111",
  38780=>"000001000",
  38781=>"000010010",
  38782=>"111010110",
  38783=>"111111010",
  38784=>"000000000",
  38785=>"000110000",
  38786=>"000101011",
  38787=>"001101111",
  38788=>"111111111",
  38789=>"000000000",
  38790=>"000000000",
  38791=>"000000000",
  38792=>"111110000",
  38793=>"000000000",
  38794=>"000111111",
  38795=>"000101111",
  38796=>"000000010",
  38797=>"111111111",
  38798=>"111111111",
  38799=>"011010011",
  38800=>"110100000",
  38801=>"111101000",
  38802=>"011001110",
  38803=>"000000000",
  38804=>"110101100",
  38805=>"110010010",
  38806=>"111111111",
  38807=>"110010101",
  38808=>"111111101",
  38809=>"000000101",
  38810=>"111000000",
  38811=>"111010010",
  38812=>"110110000",
  38813=>"100101111",
  38814=>"010100010",
  38815=>"000000000",
  38816=>"110110011",
  38817=>"011000111",
  38818=>"011000000",
  38819=>"000001111",
  38820=>"000110110",
  38821=>"110110110",
  38822=>"011001011",
  38823=>"101001101",
  38824=>"000000001",
  38825=>"111101111",
  38826=>"111000000",
  38827=>"001001101",
  38828=>"111000000",
  38829=>"000000110",
  38830=>"111111111",
  38831=>"100110111",
  38832=>"111000010",
  38833=>"000100010",
  38834=>"010010000",
  38835=>"010010000",
  38836=>"111010100",
  38837=>"101000011",
  38838=>"000010001",
  38839=>"001101110",
  38840=>"100000000",
  38841=>"110000000",
  38842=>"010101100",
  38843=>"000001000",
  38844=>"010000010",
  38845=>"110000000",
  38846=>"100100100",
  38847=>"000010000",
  38848=>"001001011",
  38849=>"000000000",
  38850=>"001011111",
  38851=>"101110110",
  38852=>"000000000",
  38853=>"111011111",
  38854=>"000000101",
  38855=>"111111010",
  38856=>"111101101",
  38857=>"111010000",
  38858=>"011001110",
  38859=>"000001001",
  38860=>"110111111",
  38861=>"010000001",
  38862=>"111111110",
  38863=>"111111110",
  38864=>"111000111",
  38865=>"111111110",
  38866=>"000000001",
  38867=>"000000010",
  38868=>"111111001",
  38869=>"000000001",
  38870=>"111101101",
  38871=>"100000000",
  38872=>"001001000",
  38873=>"000000010",
  38874=>"111011111",
  38875=>"000111111",
  38876=>"000111010",
  38877=>"000000111",
  38878=>"000000101",
  38879=>"110111100",
  38880=>"111001101",
  38881=>"101001111",
  38882=>"110110110",
  38883=>"001000001",
  38884=>"111001110",
  38885=>"000000111",
  38886=>"110100001",
  38887=>"000101101",
  38888=>"111000100",
  38889=>"000111000",
  38890=>"011001000",
  38891=>"111111111",
  38892=>"000001001",
  38893=>"110111100",
  38894=>"110010010",
  38895=>"000010000",
  38896=>"000000000",
  38897=>"100100011",
  38898=>"111110111",
  38899=>"110111101",
  38900=>"011111111",
  38901=>"000101111",
  38902=>"110101000",
  38903=>"111111111",
  38904=>"110111000",
  38905=>"000111111",
  38906=>"111101101",
  38907=>"001000000",
  38908=>"111111110",
  38909=>"111011111",
  38910=>"001011000",
  38911=>"111111011",
  38912=>"011011001",
  38913=>"000100111",
  38914=>"101101001",
  38915=>"000010111",
  38916=>"100000110",
  38917=>"111110000",
  38918=>"001000000",
  38919=>"101101111",
  38920=>"111111111",
  38921=>"111111001",
  38922=>"001100000",
  38923=>"011111111",
  38924=>"000010011",
  38925=>"000000001",
  38926=>"100100101",
  38927=>"000110000",
  38928=>"000001111",
  38929=>"000111100",
  38930=>"110011010",
  38931=>"111111111",
  38932=>"111000000",
  38933=>"000000011",
  38934=>"100000100",
  38935=>"010010010",
  38936=>"000000011",
  38937=>"001010011",
  38938=>"111111101",
  38939=>"110000000",
  38940=>"111111000",
  38941=>"000000101",
  38942=>"110110000",
  38943=>"000000100",
  38944=>"111111000",
  38945=>"111011001",
  38946=>"111000000",
  38947=>"000011111",
  38948=>"011011001",
  38949=>"111110101",
  38950=>"111101000",
  38951=>"000010000",
  38952=>"000000000",
  38953=>"001111111",
  38954=>"011111101",
  38955=>"011000000",
  38956=>"001011011",
  38957=>"000000010",
  38958=>"111011111",
  38959=>"000111001",
  38960=>"000010010",
  38961=>"001111111",
  38962=>"111111011",
  38963=>"000001000",
  38964=>"111000000",
  38965=>"000010011",
  38966=>"101001000",
  38967=>"000010010",
  38968=>"000000001",
  38969=>"000000000",
  38970=>"001010111",
  38971=>"000100111",
  38972=>"000110110",
  38973=>"011001010",
  38974=>"000000100",
  38975=>"011011001",
  38976=>"101111011",
  38977=>"111111000",
  38978=>"011111111",
  38979=>"101001011",
  38980=>"010010000",
  38981=>"100110011",
  38982=>"111111011",
  38983=>"111000110",
  38984=>"000000100",
  38985=>"010010011",
  38986=>"000000111",
  38987=>"110100010",
  38988=>"001111111",
  38989=>"110100111",
  38990=>"000111011",
  38991=>"000111110",
  38992=>"010000101",
  38993=>"000000000",
  38994=>"010111101",
  38995=>"011011001",
  38996=>"101111111",
  38997=>"000000001",
  38998=>"011111001",
  38999=>"111111101",
  39000=>"000001000",
  39001=>"100111111",
  39002=>"010111110",
  39003=>"111010111",
  39004=>"111111001",
  39005=>"001011000",
  39006=>"101000110",
  39007=>"110111111",
  39008=>"110111111",
  39009=>"110110000",
  39010=>"111101100",
  39011=>"100100101",
  39012=>"010110010",
  39013=>"101111100",
  39014=>"111111101",
  39015=>"000010001",
  39016=>"111010010",
  39017=>"111111010",
  39018=>"101111111",
  39019=>"000010000",
  39020=>"000010000",
  39021=>"000100100",
  39022=>"000010010",
  39023=>"101111100",
  39024=>"111110010",
  39025=>"000000010",
  39026=>"101000100",
  39027=>"101111011",
  39028=>"111011011",
  39029=>"101000101",
  39030=>"000001111",
  39031=>"111111111",
  39032=>"110111101",
  39033=>"011110000",
  39034=>"010010000",
  39035=>"000000000",
  39036=>"100110110",
  39037=>"110110100",
  39038=>"000000000",
  39039=>"111000100",
  39040=>"010110101",
  39041=>"111111000",
  39042=>"111111111",
  39043=>"000000100",
  39044=>"000111111",
  39045=>"000000111",
  39046=>"111111001",
  39047=>"100101111",
  39048=>"011111100",
  39049=>"111100010",
  39050=>"011111110",
  39051=>"010011000",
  39052=>"110010100",
  39053=>"100111111",
  39054=>"111111000",
  39055=>"111001001",
  39056=>"010111011",
  39057=>"100000000",
  39058=>"010010111",
  39059=>"111000011",
  39060=>"001011111",
  39061=>"101111111",
  39062=>"010011000",
  39063=>"001011011",
  39064=>"100111111",
  39065=>"100111111",
  39066=>"111000101",
  39067=>"011111101",
  39068=>"100101100",
  39069=>"010011000",
  39070=>"111111101",
  39071=>"000000000",
  39072=>"101001000",
  39073=>"000101000",
  39074=>"000000000",
  39075=>"001011100",
  39076=>"111111110",
  39077=>"001000110",
  39078=>"111110110",
  39079=>"010010000",
  39080=>"000000101",
  39081=>"000011111",
  39082=>"000111111",
  39083=>"111100000",
  39084=>"111011110",
  39085=>"111111111",
  39086=>"111100000",
  39087=>"101101111",
  39088=>"111000111",
  39089=>"001101001",
  39090=>"111111111",
  39091=>"101010000",
  39092=>"000000100",
  39093=>"000110011",
  39094=>"111011001",
  39095=>"010010111",
  39096=>"010111011",
  39097=>"000100111",
  39098=>"111111100",
  39099=>"000110111",
  39100=>"010011001",
  39101=>"011111111",
  39102=>"111111111",
  39103=>"001000000",
  39104=>"111001111",
  39105=>"110111111",
  39106=>"011101101",
  39107=>"000010011",
  39108=>"101000000",
  39109=>"000000001",
  39110=>"000011010",
  39111=>"111100111",
  39112=>"000111111",
  39113=>"010000111",
  39114=>"111000000",
  39115=>"000000011",
  39116=>"100000100",
  39117=>"000011011",
  39118=>"111010110",
  39119=>"000111011",
  39120=>"010000010",
  39121=>"101110011",
  39122=>"111011111",
  39123=>"111111011",
  39124=>"001000101",
  39125=>"110000110",
  39126=>"000000100",
  39127=>"000011111",
  39128=>"100101101",
  39129=>"010000000",
  39130=>"010100000",
  39131=>"000111000",
  39132=>"001001101",
  39133=>"010111111",
  39134=>"011101111",
  39135=>"000000111",
  39136=>"000000110",
  39137=>"111000100",
  39138=>"000000111",
  39139=>"001111000",
  39140=>"111111100",
  39141=>"000011010",
  39142=>"111111111",
  39143=>"000001000",
  39144=>"110010010",
  39145=>"101000101",
  39146=>"100000000",
  39147=>"011010010",
  39148=>"000000101",
  39149=>"011111111",
  39150=>"010010010",
  39151=>"010110000",
  39152=>"010111100",
  39153=>"000000000",
  39154=>"011011111",
  39155=>"000111011",
  39156=>"110110100",
  39157=>"111010010",
  39158=>"000000000",
  39159=>"000000011",
  39160=>"001000111",
  39161=>"111100110",
  39162=>"000010101",
  39163=>"100100111",
  39164=>"000000000",
  39165=>"000000000",
  39166=>"000111101",
  39167=>"110110111",
  39168=>"011011001",
  39169=>"110100110",
  39170=>"111000100",
  39171=>"011000000",
  39172=>"000000110",
  39173=>"101101000",
  39174=>"010110000",
  39175=>"000101101",
  39176=>"000000000",
  39177=>"100000000",
  39178=>"001001101",
  39179=>"111111010",
  39180=>"111101101",
  39181=>"110111001",
  39182=>"010101011",
  39183=>"011110000",
  39184=>"000000010",
  39185=>"000000000",
  39186=>"010111000",
  39187=>"000000111",
  39188=>"000000100",
  39189=>"111100100",
  39190=>"100010011",
  39191=>"111000000",
  39192=>"000000000",
  39193=>"000110110",
  39194=>"010111000",
  39195=>"111000111",
  39196=>"110010111",
  39197=>"111000000",
  39198=>"110010000",
  39199=>"111111011",
  39200=>"001000000",
  39201=>"001010010",
  39202=>"001001000",
  39203=>"101101000",
  39204=>"110110110",
  39205=>"000100100",
  39206=>"101000111",
  39207=>"000010010",
  39208=>"010010000",
  39209=>"000011011",
  39210=>"000001000",
  39211=>"000110111",
  39212=>"100111101",
  39213=>"111111110",
  39214=>"010001101",
  39215=>"000110000",
  39216=>"101000001",
  39217=>"110000110",
  39218=>"000000000",
  39219=>"000111111",
  39220=>"100000100",
  39221=>"000000000",
  39222=>"110111111",
  39223=>"111111101",
  39224=>"010111010",
  39225=>"111011011",
  39226=>"000000000",
  39227=>"000010000",
  39228=>"110100100",
  39229=>"001010001",
  39230=>"010101001",
  39231=>"001001101",
  39232=>"000011111",
  39233=>"101000000",
  39234=>"111111000",
  39235=>"101001001",
  39236=>"110000000",
  39237=>"001000000",
  39238=>"010111111",
  39239=>"010110000",
  39240=>"011101001",
  39241=>"111101000",
  39242=>"111000000",
  39243=>"001001000",
  39244=>"000000000",
  39245=>"110110111",
  39246=>"001001111",
  39247=>"100000000",
  39248=>"001010010",
  39249=>"111111111",
  39250=>"000011010",
  39251=>"010010000",
  39252=>"000000000",
  39253=>"101101111",
  39254=>"000001010",
  39255=>"111000111",
  39256=>"010000100",
  39257=>"011010111",
  39258=>"000101111",
  39259=>"001011000",
  39260=>"000010000",
  39261=>"001001000",
  39262=>"111111101",
  39263=>"100000110",
  39264=>"000010000",
  39265=>"010000001",
  39266=>"111101000",
  39267=>"000000100",
  39268=>"011101010",
  39269=>"000011000",
  39270=>"000000101",
  39271=>"011000000",
  39272=>"000010110",
  39273=>"111011001",
  39274=>"000010011",
  39275=>"111101100",
  39276=>"010010001",
  39277=>"111000110",
  39278=>"111101000",
  39279=>"101000100",
  39280=>"000111101",
  39281=>"010000000",
  39282=>"001011011",
  39283=>"000000000",
  39284=>"100010111",
  39285=>"101100010",
  39286=>"011111110",
  39287=>"101000000",
  39288=>"000000001",
  39289=>"110011010",
  39290=>"111111111",
  39291=>"011101101",
  39292=>"000100100",
  39293=>"000010000",
  39294=>"110000001",
  39295=>"000001001",
  39296=>"010110000",
  39297=>"010101100",
  39298=>"111010000",
  39299=>"000001101",
  39300=>"111100000",
  39301=>"110110000",
  39302=>"010011001",
  39303=>"000001011",
  39304=>"000111000",
  39305=>"111011000",
  39306=>"111000111",
  39307=>"101001010",
  39308=>"111000000",
  39309=>"000111111",
  39310=>"111111000",
  39311=>"000000000",
  39312=>"111101011",
  39313=>"010000111",
  39314=>"000010000",
  39315=>"101000000",
  39316=>"000000111",
  39317=>"000000010",
  39318=>"101001000",
  39319=>"100100110",
  39320=>"110010100",
  39321=>"011000000",
  39322=>"110111000",
  39323=>"100100100",
  39324=>"010100000",
  39325=>"001000000",
  39326=>"010010010",
  39327=>"111000010",
  39328=>"110101111",
  39329=>"000000110",
  39330=>"110101111",
  39331=>"000100001",
  39332=>"110110110",
  39333=>"100110110",
  39334=>"000000110",
  39335=>"000110000",
  39336=>"010110011",
  39337=>"011111110",
  39338=>"101110110",
  39339=>"000000000",
  39340=>"000001101",
  39341=>"110000010",
  39342=>"001110100",
  39343=>"110011000",
  39344=>"100101101",
  39345=>"100101101",
  39346=>"111101000",
  39347=>"011000000",
  39348=>"001011110",
  39349=>"010011000",
  39350=>"000011011",
  39351=>"010011001",
  39352=>"011001001",
  39353=>"000100110",
  39354=>"110110010",
  39355=>"111111000",
  39356=>"010010000",
  39357=>"111111111",
  39358=>"001000100",
  39359=>"110000011",
  39360=>"000000000",
  39361=>"010000001",
  39362=>"111101001",
  39363=>"001010110",
  39364=>"011000000",
  39365=>"110101111",
  39366=>"110110110",
  39367=>"001000001",
  39368=>"000000101",
  39369=>"101000000",
  39370=>"010110000",
  39371=>"101001111",
  39372=>"000000001",
  39373=>"100011001",
  39374=>"000000000",
  39375=>"001111101",
  39376=>"111000000",
  39377=>"010111011",
  39378=>"000100011",
  39379=>"111000000",
  39380=>"101000000",
  39381=>"111111001",
  39382=>"110101000",
  39383=>"110010000",
  39384=>"000000000",
  39385=>"101000000",
  39386=>"111001111",
  39387=>"011001111",
  39388=>"001100010",
  39389=>"001111000",
  39390=>"010110000",
  39391=>"100110011",
  39392=>"111000101",
  39393=>"101101100",
  39394=>"111111111",
  39395=>"001001000",
  39396=>"111000010",
  39397=>"011011010",
  39398=>"000111111",
  39399=>"010000011",
  39400=>"100101000",
  39401=>"000000101",
  39402=>"110000001",
  39403=>"001111111",
  39404=>"101001000",
  39405=>"000000011",
  39406=>"010000000",
  39407=>"000001010",
  39408=>"111001000",
  39409=>"011001100",
  39410=>"101101101",
  39411=>"010110001",
  39412=>"010110111",
  39413=>"011000011",
  39414=>"010000000",
  39415=>"000010110",
  39416=>"010010011",
  39417=>"111000000",
  39418=>"010010011",
  39419=>"001011000",
  39420=>"111100101",
  39421=>"111111111",
  39422=>"000011011",
  39423=>"010001111",
  39424=>"011001000",
  39425=>"000000100",
  39426=>"101001101",
  39427=>"011101001",
  39428=>"011011010",
  39429=>"100000001",
  39430=>"010000000",
  39431=>"000011010",
  39432=>"000100010",
  39433=>"111101111",
  39434=>"101001011",
  39435=>"011011000",
  39436=>"010000000",
  39437=>"100000101",
  39438=>"000011001",
  39439=>"010110111",
  39440=>"000110010",
  39441=>"111101000",
  39442=>"000001001",
  39443=>"000010000",
  39444=>"000111101",
  39445=>"110000000",
  39446=>"001100101",
  39447=>"101101111",
  39448=>"101000011",
  39449=>"111010110",
  39450=>"000000000",
  39451=>"101101000",
  39452=>"000000000",
  39453=>"000001111",
  39454=>"111000000",
  39455=>"111111101",
  39456=>"000110111",
  39457=>"010011111",
  39458=>"000011000",
  39459=>"000011010",
  39460=>"000001011",
  39461=>"000000000",
  39462=>"011110000",
  39463=>"011000100",
  39464=>"000000001",
  39465=>"111110111",
  39466=>"001011000",
  39467=>"111011000",
  39468=>"000000001",
  39469=>"100000011",
  39470=>"011111111",
  39471=>"111101110",
  39472=>"000010111",
  39473=>"001011110",
  39474=>"000000010",
  39475=>"000110111",
  39476=>"010010000",
  39477=>"010110100",
  39478=>"100001001",
  39479=>"000000110",
  39480=>"100111111",
  39481=>"000000100",
  39482=>"000000000",
  39483=>"101100100",
  39484=>"110110100",
  39485=>"010111001",
  39486=>"000000000",
  39487=>"111011111",
  39488=>"111011111",
  39489=>"010010110",
  39490=>"000000111",
  39491=>"001000000",
  39492=>"010111101",
  39493=>"010010000",
  39494=>"000000111",
  39495=>"010010111",
  39496=>"011001100",
  39497=>"010000000",
  39498=>"000000001",
  39499=>"111101001",
  39500=>"111111110",
  39501=>"001110110",
  39502=>"100110010",
  39503=>"100101001",
  39504=>"100000100",
  39505=>"000000010",
  39506=>"000100111",
  39507=>"011000000",
  39508=>"001000001",
  39509=>"111100100",
  39510=>"001001011",
  39511=>"000110000",
  39512=>"111111000",
  39513=>"000000111",
  39514=>"111111000",
  39515=>"000100000",
  39516=>"111011010",
  39517=>"000000000",
  39518=>"000000110",
  39519=>"000001000",
  39520=>"110111111",
  39521=>"010111101",
  39522=>"010001100",
  39523=>"111011001",
  39524=>"000000000",
  39525=>"000100111",
  39526=>"111010111",
  39527=>"000010111",
  39528=>"000001111",
  39529=>"000000111",
  39530=>"000000000",
  39531=>"011010011",
  39532=>"100111111",
  39533=>"101101111",
  39534=>"000000000",
  39535=>"000000110",
  39536=>"001001010",
  39537=>"000000010",
  39538=>"001100010",
  39539=>"111111111",
  39540=>"000000000",
  39541=>"000100000",
  39542=>"010010011",
  39543=>"111101000",
  39544=>"111000000",
  39545=>"111111000",
  39546=>"000000100",
  39547=>"000001001",
  39548=>"100111011",
  39549=>"110000100",
  39550=>"010001001",
  39551=>"100011000",
  39552=>"000000000",
  39553=>"000010010",
  39554=>"110000100",
  39555=>"010100000",
  39556=>"001000110",
  39557=>"000000000",
  39558=>"011000000",
  39559=>"000111000",
  39560=>"110110110",
  39561=>"101010011",
  39562=>"111101111",
  39563=>"111011001",
  39564=>"111000111",
  39565=>"011111101",
  39566=>"100111010",
  39567=>"001001110",
  39568=>"100111011",
  39569=>"101010000",
  39570=>"111000010",
  39571=>"011101111",
  39572=>"000011011",
  39573=>"010110111",
  39574=>"000111111",
  39575=>"000011001",
  39576=>"000000101",
  39577=>"000000000",
  39578=>"000000111",
  39579=>"000101111",
  39580=>"110010100",
  39581=>"000000010",
  39582=>"000000110",
  39583=>"111111000",
  39584=>"111100000",
  39585=>"111000000",
  39586=>"010111101",
  39587=>"000110101",
  39588=>"111000000",
  39589=>"110010000",
  39590=>"000110000",
  39591=>"000000010",
  39592=>"000000010",
  39593=>"000010111",
  39594=>"111111100",
  39595=>"111000000",
  39596=>"111111000",
  39597=>"100110110",
  39598=>"111101111",
  39599=>"101101110",
  39600=>"000001000",
  39601=>"100000101",
  39602=>"000000000",
  39603=>"000000000",
  39604=>"111000100",
  39605=>"001011111",
  39606=>"011011111",
  39607=>"011011001",
  39608=>"011110000",
  39609=>"000110111",
  39610=>"110000001",
  39611=>"111011000",
  39612=>"011001101",
  39613=>"000100111",
  39614=>"011010010",
  39615=>"011001000",
  39616=>"100000000",
  39617=>"101000000",
  39618=>"001001101",
  39619=>"111110111",
  39620=>"000111000",
  39621=>"101011111",
  39622=>"000010010",
  39623=>"100000101",
  39624=>"000111111",
  39625=>"110000000",
  39626=>"011011111",
  39627=>"000001111",
  39628=>"000000000",
  39629=>"001011110",
  39630=>"111110110",
  39631=>"110111111",
  39632=>"111101000",
  39633=>"110110110",
  39634=>"100010111",
  39635=>"111011111",
  39636=>"000000011",
  39637=>"001100100",
  39638=>"010011111",
  39639=>"000011110",
  39640=>"111101101",
  39641=>"000000111",
  39642=>"111011001",
  39643=>"000001101",
  39644=>"111100101",
  39645=>"000111011",
  39646=>"111010000",
  39647=>"000001101",
  39648=>"101000100",
  39649=>"011001101",
  39650=>"111111101",
  39651=>"101111110",
  39652=>"101000011",
  39653=>"110110000",
  39654=>"111011111",
  39655=>"011111111",
  39656=>"001000000",
  39657=>"010000100",
  39658=>"100100111",
  39659=>"110111111",
  39660=>"111110000",
  39661=>"111010000",
  39662=>"000000000",
  39663=>"011111100",
  39664=>"111111100",
  39665=>"111111101",
  39666=>"011010000",
  39667=>"000001001",
  39668=>"110110000",
  39669=>"110100111",
  39670=>"000000000",
  39671=>"000000000",
  39672=>"010000000",
  39673=>"000000001",
  39674=>"111100000",
  39675=>"100111111",
  39676=>"000000011",
  39677=>"000010111",
  39678=>"100011001",
  39679=>"000000101",
  39680=>"111111111",
  39681=>"010000101",
  39682=>"000000000",
  39683=>"000001111",
  39684=>"000111111",
  39685=>"001001000",
  39686=>"000101101",
  39687=>"101001111",
  39688=>"111001010",
  39689=>"001001111",
  39690=>"001000000",
  39691=>"001000111",
  39692=>"000000000",
  39693=>"011001001",
  39694=>"111101101",
  39695=>"111011111",
  39696=>"110000111",
  39697=>"000000000",
  39698=>"110000100",
  39699=>"000000000",
  39700=>"111111111",
  39701=>"010000110",
  39702=>"001011001",
  39703=>"101010000",
  39704=>"000000000",
  39705=>"111111111",
  39706=>"111011011",
  39707=>"111111000",
  39708=>"000000000",
  39709=>"111001001",
  39710=>"001011111",
  39711=>"001000000",
  39712=>"111111110",
  39713=>"101111111",
  39714=>"000000000",
  39715=>"000011011",
  39716=>"000100000",
  39717=>"011011011",
  39718=>"001011110",
  39719=>"000001000",
  39720=>"111111010",
  39721=>"011111111",
  39722=>"000000011",
  39723=>"100000111",
  39724=>"010111100",
  39725=>"111111100",
  39726=>"000001000",
  39727=>"010111011",
  39728=>"101111000",
  39729=>"100100001",
  39730=>"001010001",
  39731=>"010111101",
  39732=>"000000000",
  39733=>"101111111",
  39734=>"000000001",
  39735=>"111101101",
  39736=>"100011111",
  39737=>"111001000",
  39738=>"111000111",
  39739=>"000011111",
  39740=>"011011010",
  39741=>"001111111",
  39742=>"000000000",
  39743=>"001101110",
  39744=>"010100111",
  39745=>"001111110",
  39746=>"000000000",
  39747=>"100000100",
  39748=>"111100000",
  39749=>"000000000",
  39750=>"100110111",
  39751=>"001001011",
  39752=>"011110001",
  39753=>"011111001",
  39754=>"101001000",
  39755=>"111100000",
  39756=>"111000000",
  39757=>"000010001",
  39758=>"110001111",
  39759=>"001001011",
  39760=>"000000000",
  39761=>"101111111",
  39762=>"111111010",
  39763=>"101111010",
  39764=>"000001111",
  39765=>"000010011",
  39766=>"000111110",
  39767=>"101001111",
  39768=>"111000010",
  39769=>"110000001",
  39770=>"101011011",
  39771=>"010101000",
  39772=>"000111111",
  39773=>"100000101",
  39774=>"111111100",
  39775=>"001000001",
  39776=>"001000000",
  39777=>"010000101",
  39778=>"000001000",
  39779=>"011000000",
  39780=>"111110111",
  39781=>"101111000",
  39782=>"110110001",
  39783=>"111010010",
  39784=>"011101000",
  39785=>"110010101",
  39786=>"000111100",
  39787=>"001000111",
  39788=>"010001111",
  39789=>"000000001",
  39790=>"000000111",
  39791=>"111101000",
  39792=>"001011010",
  39793=>"111111111",
  39794=>"000000001",
  39795=>"000000000",
  39796=>"001000000",
  39797=>"011000110",
  39798=>"001111001",
  39799=>"000000111",
  39800=>"111011001",
  39801=>"100101111",
  39802=>"111111110",
  39803=>"100000000",
  39804=>"001011011",
  39805=>"011000000",
  39806=>"000000001",
  39807=>"001000000",
  39808=>"010100000",
  39809=>"001001000",
  39810=>"000011011",
  39811=>"111000111",
  39812=>"000110000",
  39813=>"010110110",
  39814=>"100111100",
  39815=>"111100101",
  39816=>"001101000",
  39817=>"110111010",
  39818=>"001111111",
  39819=>"001000101",
  39820=>"111000000",
  39821=>"001001001",
  39822=>"001111111",
  39823=>"110000000",
  39824=>"111110010",
  39825=>"011111000",
  39826=>"111111001",
  39827=>"111111111",
  39828=>"111101001",
  39829=>"000000001",
  39830=>"000000000",
  39831=>"101100111",
  39832=>"001000010",
  39833=>"000100111",
  39834=>"001111111",
  39835=>"001001011",
  39836=>"111101100",
  39837=>"000100000",
  39838=>"011111110",
  39839=>"111000000",
  39840=>"000010011",
  39841=>"000000000",
  39842=>"001000000",
  39843=>"000000000",
  39844=>"000111111",
  39845=>"101000010",
  39846=>"011111111",
  39847=>"000111011",
  39848=>"000000100",
  39849=>"101001111",
  39850=>"000000001",
  39851=>"100000000",
  39852=>"000101111",
  39853=>"000000000",
  39854=>"000000000",
  39855=>"000000110",
  39856=>"000001000",
  39857=>"000100101",
  39858=>"111111101",
  39859=>"011010011",
  39860=>"111010000",
  39861=>"110111011",
  39862=>"010000001",
  39863=>"111111111",
  39864=>"100100100",
  39865=>"011110011",
  39866=>"110110110",
  39867=>"000000011",
  39868=>"111111111",
  39869=>"110000010",
  39870=>"010001000",
  39871=>"000001011",
  39872=>"010000000",
  39873=>"000000111",
  39874=>"111010011",
  39875=>"000000000",
  39876=>"111111111",
  39877=>"011010111",
  39878=>"000001001",
  39879=>"001001111",
  39880=>"000000111",
  39881=>"000000000",
  39882=>"000000000",
  39883=>"000001111",
  39884=>"000000000",
  39885=>"100100100",
  39886=>"111111111",
  39887=>"110001111",
  39888=>"000000000",
  39889=>"001001100",
  39890=>"110100111",
  39891=>"111001001",
  39892=>"000001001",
  39893=>"000001000",
  39894=>"011000000",
  39895=>"001001011",
  39896=>"011111000",
  39897=>"111111000",
  39898=>"111101111",
  39899=>"000000000",
  39900=>"111101100",
  39901=>"000000111",
  39902=>"000000110",
  39903=>"111110000",
  39904=>"111001001",
  39905=>"101001001",
  39906=>"110000001",
  39907=>"111010011",
  39908=>"011000001",
  39909=>"111001100",
  39910=>"000100111",
  39911=>"001000000",
  39912=>"000110000",
  39913=>"111001001",
  39914=>"000001000",
  39915=>"001011111",
  39916=>"101011000",
  39917=>"000000000",
  39918=>"100000101",
  39919=>"000000111",
  39920=>"000110110",
  39921=>"101111111",
  39922=>"001001110",
  39923=>"010101000",
  39924=>"110111000",
  39925=>"110000001",
  39926=>"000000000",
  39927=>"111111110",
  39928=>"111000000",
  39929=>"001010110",
  39930=>"111111111",
  39931=>"111110111",
  39932=>"111010011",
  39933=>"110111111",
  39934=>"000111111",
  39935=>"010000000",
  39936=>"011001100",
  39937=>"000001000",
  39938=>"101100111",
  39939=>"101101011",
  39940=>"111101110",
  39941=>"011000111",
  39942=>"101100000",
  39943=>"001010010",
  39944=>"000000000",
  39945=>"000000010",
  39946=>"001001101",
  39947=>"101000000",
  39948=>"111000000",
  39949=>"010010000",
  39950=>"001011000",
  39951=>"100100101",
  39952=>"000000000",
  39953=>"111000010",
  39954=>"001011000",
  39955=>"111011000",
  39956=>"111011101",
  39957=>"100100111",
  39958=>"100101100",
  39959=>"111101000",
  39960=>"001000010",
  39961=>"011011111",
  39962=>"011111111",
  39963=>"111111100",
  39964=>"100000000",
  39965=>"000000011",
  39966=>"101010010",
  39967=>"000001111",
  39968=>"000001101",
  39969=>"111111111",
  39970=>"111100000",
  39971=>"111000000",
  39972=>"011011011",
  39973=>"011000111",
  39974=>"111011111",
  39975=>"000101111",
  39976=>"111110000",
  39977=>"010010000",
  39978=>"000100000",
  39979=>"011000000",
  39980=>"001011111",
  39981=>"001010011",
  39982=>"111111111",
  39983=>"000101100",
  39984=>"001000111",
  39985=>"111110100",
  39986=>"010111011",
  39987=>"100000111",
  39988=>"011010001",
  39989=>"000111000",
  39990=>"000000001",
  39991=>"000000010",
  39992=>"101000000",
  39993=>"001000100",
  39994=>"000100000",
  39995=>"101101111",
  39996=>"111111111",
  39997=>"001101101",
  39998=>"010000000",
  39999=>"011011110",
  40000=>"111000000",
  40001=>"111010000",
  40002=>"010111111",
  40003=>"111110000",
  40004=>"000000111",
  40005=>"000000000",
  40006=>"010001111",
  40007=>"111111000",
  40008=>"010111111",
  40009=>"100100000",
  40010=>"001000000",
  40011=>"000100111",
  40012=>"000000000",
  40013=>"101010000",
  40014=>"111111111",
  40015=>"100000001",
  40016=>"000111111",
  40017=>"011000000",
  40018=>"011101111",
  40019=>"011000100",
  40020=>"111001111",
  40021=>"011011111",
  40022=>"111011000",
  40023=>"100111110",
  40024=>"111000000",
  40025=>"100100100",
  40026=>"100000011",
  40027=>"111100000",
  40028=>"000010000",
  40029=>"000001111",
  40030=>"010010010",
  40031=>"011011000",
  40032=>"111111010",
  40033=>"000000111",
  40034=>"010000101",
  40035=>"000000100",
  40036=>"000000000",
  40037=>"111111100",
  40038=>"110111100",
  40039=>"100111100",
  40040=>"000001011",
  40041=>"111001111",
  40042=>"011111010",
  40043=>"011111000",
  40044=>"000110111",
  40045=>"001001000",
  40046=>"000000111",
  40047=>"011000011",
  40048=>"001011110",
  40049=>"010010110",
  40050=>"010100100",
  40051=>"111111111",
  40052=>"100111100",
  40053=>"001000000",
  40054=>"100000000",
  40055=>"111000000",
  40056=>"111111000",
  40057=>"111111000",
  40058=>"000000101",
  40059=>"101001011",
  40060=>"000010011",
  40061=>"110100001",
  40062=>"110000001",
  40063=>"000000000",
  40064=>"101010000",
  40065=>"000000011",
  40066=>"110000001",
  40067=>"000000000",
  40068=>"111011100",
  40069=>"011100000",
  40070=>"011101111",
  40071=>"010000110",
  40072=>"100000011",
  40073=>"000000111",
  40074=>"111101100",
  40075=>"111111000",
  40076=>"000000111",
  40077=>"000001111",
  40078=>"000000010",
  40079=>"000000000",
  40080=>"000000001",
  40081=>"001001010",
  40082=>"101101111",
  40083=>"111101100",
  40084=>"100100100",
  40085=>"111000000",
  40086=>"000101111",
  40087=>"011001000",
  40088=>"101100000",
  40089=>"000111011",
  40090=>"111010010",
  40091=>"100100011",
  40092=>"000000000",
  40093=>"111111111",
  40094=>"111000110",
  40095=>"000000000",
  40096=>"000010011",
  40097=>"100100111",
  40098=>"111000000",
  40099=>"111111111",
  40100=>"000101000",
  40101=>"010001001",
  40102=>"111111000",
  40103=>"001111110",
  40104=>"000010111",
  40105=>"000111011",
  40106=>"101100000",
  40107=>"101000010",
  40108=>"111011000",
  40109=>"111000100",
  40110=>"101001010",
  40111=>"110010000",
  40112=>"000000000",
  40113=>"100001001",
  40114=>"000101111",
  40115=>"000100000",
  40116=>"100101000",
  40117=>"100100011",
  40118=>"000000000",
  40119=>"110111111",
  40120=>"001111110",
  40121=>"011001001",
  40122=>"101110111",
  40123=>"111110011",
  40124=>"001010001",
  40125=>"000011110",
  40126=>"001001100",
  40127=>"001000011",
  40128=>"000000111",
  40129=>"101000101",
  40130=>"101111111",
  40131=>"000010000",
  40132=>"000101000",
  40133=>"001011111",
  40134=>"000010000",
  40135=>"000100111",
  40136=>"000011000",
  40137=>"000000000",
  40138=>"111101110",
  40139=>"101100010",
  40140=>"101100101",
  40141=>"010000111",
  40142=>"000000111",
  40143=>"111111000",
  40144=>"111001101",
  40145=>"110110110",
  40146=>"111100000",
  40147=>"101100000",
  40148=>"000000111",
  40149=>"000100111",
  40150=>"111111111",
  40151=>"111000000",
  40152=>"111011100",
  40153=>"001011000",
  40154=>"000100100",
  40155=>"001000001",
  40156=>"010010111",
  40157=>"100011010",
  40158=>"110100011",
  40159=>"110010010",
  40160=>"010000000",
  40161=>"100000111",
  40162=>"111100000",
  40163=>"101111000",
  40164=>"111000111",
  40165=>"000111111",
  40166=>"011000000",
  40167=>"000100111",
  40168=>"111000101",
  40169=>"000010111",
  40170=>"001001111",
  40171=>"000000110",
  40172=>"011010000",
  40173=>"111000001",
  40174=>"000000000",
  40175=>"000000110",
  40176=>"000110000",
  40177=>"100011010",
  40178=>"001110000",
  40179=>"101101011",
  40180=>"110001000",
  40181=>"111100110",
  40182=>"001111011",
  40183=>"101000000",
  40184=>"000000111",
  40185=>"100001000",
  40186=>"111001111",
  40187=>"100101000",
  40188=>"000010000",
  40189=>"001101000",
  40190=>"110101000",
  40191=>"101011000",
  40192=>"000111111",
  40193=>"111000111",
  40194=>"000100011",
  40195=>"111010000",
  40196=>"110111111",
  40197=>"001000000",
  40198=>"000110111",
  40199=>"100111010",
  40200=>"000110111",
  40201=>"100010111",
  40202=>"000000000",
  40203=>"100001111",
  40204=>"000000101",
  40205=>"000010101",
  40206=>"011101001",
  40207=>"011100111",
  40208=>"111000010",
  40209=>"000000011",
  40210=>"110101101",
  40211=>"001011111",
  40212=>"111101001",
  40213=>"001001001",
  40214=>"101100100",
  40215=>"000100100",
  40216=>"000000111",
  40217=>"010111111",
  40218=>"000000000",
  40219=>"000011011",
  40220=>"001001100",
  40221=>"110010000",
  40222=>"101101000",
  40223=>"111000000",
  40224=>"001000001",
  40225=>"101111111",
  40226=>"100111111",
  40227=>"000100000",
  40228=>"000100101",
  40229=>"100000100",
  40230=>"000000000",
  40231=>"000001111",
  40232=>"111111110",
  40233=>"000101111",
  40234=>"111000000",
  40235=>"110000001",
  40236=>"110000001",
  40237=>"111101101",
  40238=>"000101111",
  40239=>"000111010",
  40240=>"001010011",
  40241=>"001011101",
  40242=>"000000110",
  40243=>"001111110",
  40244=>"010000101",
  40245=>"111010110",
  40246=>"000000000",
  40247=>"100000000",
  40248=>"101101010",
  40249=>"001101000",
  40250=>"010000000",
  40251=>"101111110",
  40252=>"000000000",
  40253=>"000010101",
  40254=>"001000000",
  40255=>"100000000",
  40256=>"000111111",
  40257=>"100101000",
  40258=>"111010010",
  40259=>"100101000",
  40260=>"011000111",
  40261=>"010001111",
  40262=>"010010000",
  40263=>"010010111",
  40264=>"101100100",
  40265=>"011111101",
  40266=>"101001000",
  40267=>"000111011",
  40268=>"000000000",
  40269=>"001101000",
  40270=>"100100101",
  40271=>"001100111",
  40272=>"111000000",
  40273=>"000011111",
  40274=>"000010111",
  40275=>"000001000",
  40276=>"100000001",
  40277=>"100100100",
  40278=>"101101100",
  40279=>"100000100",
  40280=>"110110000",
  40281=>"110000011",
  40282=>"111001000",
  40283=>"100100100",
  40284=>"000101100",
  40285=>"011101100",
  40286=>"011101101",
  40287=>"011100000",
  40288=>"110101100",
  40289=>"000101111",
  40290=>"101000100",
  40291=>"111110000",
  40292=>"111110000",
  40293=>"001100000",
  40294=>"000110001",
  40295=>"111010010",
  40296=>"110111110",
  40297=>"111111011",
  40298=>"101101110",
  40299=>"010000000",
  40300=>"000100001",
  40301=>"110010110",
  40302=>"011111011",
  40303=>"000101001",
  40304=>"101101101",
  40305=>"111100010",
  40306=>"000000000",
  40307=>"000000100",
  40308=>"101011010",
  40309=>"001000000",
  40310=>"111011010",
  40311=>"000101101",
  40312=>"111100010",
  40313=>"111101101",
  40314=>"110110111",
  40315=>"101111101",
  40316=>"111000111",
  40317=>"000110000",
  40318=>"111110110",
  40319=>"000000000",
  40320=>"101101011",
  40321=>"100101111",
  40322=>"000101100",
  40323=>"010000010",
  40324=>"111111000",
  40325=>"010111011",
  40326=>"001001001",
  40327=>"001001111",
  40328=>"001101101",
  40329=>"001010010",
  40330=>"101010011",
  40331=>"000000010",
  40332=>"011010000",
  40333=>"000010011",
  40334=>"110011011",
  40335=>"100000010",
  40336=>"101101100",
  40337=>"111001010",
  40338=>"100000000",
  40339=>"000001101",
  40340=>"011010011",
  40341=>"101000010",
  40342=>"011011100",
  40343=>"011000000",
  40344=>"010010011",
  40345=>"111110000",
  40346=>"000010111",
  40347=>"000000011",
  40348=>"011000010",
  40349=>"000000100",
  40350=>"111000100",
  40351=>"010010111",
  40352=>"101101001",
  40353=>"111010000",
  40354=>"110000100",
  40355=>"101001010",
  40356=>"110101000",
  40357=>"001100100",
  40358=>"010010011",
  40359=>"001010110",
  40360=>"110000110",
  40361=>"010010110",
  40362=>"010100000",
  40363=>"101000000",
  40364=>"111100101",
  40365=>"010000000",
  40366=>"000011000",
  40367=>"000000000",
  40368=>"011011011",
  40369=>"010001111",
  40370=>"010110101",
  40371=>"111001110",
  40372=>"010011001",
  40373=>"000000011",
  40374=>"011100100",
  40375=>"011101000",
  40376=>"000001101",
  40377=>"110010110",
  40378=>"010010010",
  40379=>"001111101",
  40380=>"111111111",
  40381=>"010001110",
  40382=>"000001101",
  40383=>"000010010",
  40384=>"101101101",
  40385=>"000000000",
  40386=>"110111000",
  40387=>"001001001",
  40388=>"110111111",
  40389=>"100011001",
  40390=>"111110000",
  40391=>"000010111",
  40392=>"111010111",
  40393=>"000101000",
  40394=>"011111111",
  40395=>"110101110",
  40396=>"100111111",
  40397=>"111000011",
  40398=>"010000101",
  40399=>"010111010",
  40400=>"011011000",
  40401=>"111101100",
  40402=>"010111111",
  40403=>"011110000",
  40404=>"100101101",
  40405=>"110000101",
  40406=>"101101000",
  40407=>"111100000",
  40408=>"101101000",
  40409=>"000010101",
  40410=>"101110111",
  40411=>"000010010",
  40412=>"101001001",
  40413=>"010000000",
  40414=>"010000010",
  40415=>"001001111",
  40416=>"001000100",
  40417=>"011010111",
  40418=>"010010010",
  40419=>"111001000",
  40420=>"000000000",
  40421=>"111111011",
  40422=>"011011111",
  40423=>"010110000",
  40424=>"100101101",
  40425=>"010000000",
  40426=>"000000000",
  40427=>"010000001",
  40428=>"000000000",
  40429=>"000000011",
  40430=>"000000110",
  40431=>"101101101",
  40432=>"000010011",
  40433=>"001100100",
  40434=>"000101011",
  40435=>"110100000",
  40436=>"100110110",
  40437=>"111010000",
  40438=>"000000111",
  40439=>"111111111",
  40440=>"100101101",
  40441=>"111110111",
  40442=>"010111101",
  40443=>"101011011",
  40444=>"001100100",
  40445=>"110111100",
  40446=>"100001101",
  40447=>"101011000",
  40448=>"000000000",
  40449=>"000001000",
  40450=>"101101101",
  40451=>"000001000",
  40452=>"111100000",
  40453=>"111001000",
  40454=>"011011000",
  40455=>"010111111",
  40456=>"001110110",
  40457=>"000010110",
  40458=>"011001100",
  40459=>"000010101",
  40460=>"111000101",
  40461=>"111010000",
  40462=>"011000000",
  40463=>"010000000",
  40464=>"010000000",
  40465=>"010000111",
  40466=>"010101100",
  40467=>"011000000",
  40468=>"000111011",
  40469=>"000101111",
  40470=>"011101001",
  40471=>"011010100",
  40472=>"000000000",
  40473=>"100000101",
  40474=>"101101001",
  40475=>"001001010",
  40476=>"000000110",
  40477=>"111110010",
  40478=>"001101000",
  40479=>"101111011",
  40480=>"000101000",
  40481=>"110110000",
  40482=>"101101100",
  40483=>"110100000",
  40484=>"100111000",
  40485=>"100100100",
  40486=>"000000000",
  40487=>"110110000",
  40488=>"001111111",
  40489=>"000000100",
  40490=>"000000111",
  40491=>"000110000",
  40492=>"011110110",
  40493=>"010000011",
  40494=>"100000000",
  40495=>"000111010",
  40496=>"101100100",
  40497=>"010100000",
  40498=>"101101100",
  40499=>"101101000",
  40500=>"001000101",
  40501=>"101101111",
  40502=>"010111110",
  40503=>"000001011",
  40504=>"000000000",
  40505=>"000000000",
  40506=>"000101100",
  40507=>"110111101",
  40508=>"110101011",
  40509=>"111111111",
  40510=>"100001000",
  40511=>"011110100",
  40512=>"111111101",
  40513=>"010100100",
  40514=>"111010011",
  40515=>"011100100",
  40516=>"010000001",
  40517=>"000100000",
  40518=>"111000011",
  40519=>"000101010",
  40520=>"011111101",
  40521=>"001001010",
  40522=>"101101000",
  40523=>"010110000",
  40524=>"110000011",
  40525=>"110110000",
  40526=>"001000100",
  40527=>"010101000",
  40528=>"000101000",
  40529=>"111111011",
  40530=>"101101111",
  40531=>"011011000",
  40532=>"000000101",
  40533=>"111111111",
  40534=>"000100111",
  40535=>"101010010",
  40536=>"001101101",
  40537=>"001000001",
  40538=>"100011011",
  40539=>"001011000",
  40540=>"000010000",
  40541=>"001001001",
  40542=>"111011001",
  40543=>"000001001",
  40544=>"000000100",
  40545=>"000100110",
  40546=>"111100101",
  40547=>"000111110",
  40548=>"111110000",
  40549=>"001001111",
  40550=>"010000001",
  40551=>"000010010",
  40552=>"100100000",
  40553=>"111101000",
  40554=>"000010111",
  40555=>"111111101",
  40556=>"000110111",
  40557=>"011000000",
  40558=>"000001010",
  40559=>"010000111",
  40560=>"100001001",
  40561=>"001000110",
  40562=>"010011011",
  40563=>"001000000",
  40564=>"111010000",
  40565=>"000001000",
  40566=>"111001000",
  40567=>"000010110",
  40568=>"000100100",
  40569=>"101111110",
  40570=>"111100101",
  40571=>"111101101",
  40572=>"111110011",
  40573=>"010100000",
  40574=>"010110011",
  40575=>"000101101",
  40576=>"010000000",
  40577=>"000101000",
  40578=>"010111101",
  40579=>"111101000",
  40580=>"011000000",
  40581=>"111111111",
  40582=>"000011000",
  40583=>"000010000",
  40584=>"110001111",
  40585=>"111000000",
  40586=>"010000110",
  40587=>"010010111",
  40588=>"000111110",
  40589=>"100101000",
  40590=>"011100110",
  40591=>"000000000",
  40592=>"101100000",
  40593=>"101101101",
  40594=>"010111111",
  40595=>"000000000",
  40596=>"000000000",
  40597=>"001010110",
  40598=>"100101101",
  40599=>"001000000",
  40600=>"111000000",
  40601=>"101111011",
  40602=>"100000111",
  40603=>"111010000",
  40604=>"000010001",
  40605=>"011001101",
  40606=>"000000111",
  40607=>"110000000",
  40608=>"010110111",
  40609=>"000101111",
  40610=>"101101001",
  40611=>"111101000",
  40612=>"001000001",
  40613=>"100110000",
  40614=>"111111000",
  40615=>"000000010",
  40616=>"001001001",
  40617=>"000000001",
  40618=>"101101111",
  40619=>"111000000",
  40620=>"111110000",
  40621=>"101110111",
  40622=>"001001100",
  40623=>"101001111",
  40624=>"000000000",
  40625=>"100100001",
  40626=>"001101011",
  40627=>"000110110",
  40628=>"110111101",
  40629=>"010001011",
  40630=>"111111001",
  40631=>"110000111",
  40632=>"001101010",
  40633=>"000000000",
  40634=>"010001111",
  40635=>"000111011",
  40636=>"000010000",
  40637=>"111001111",
  40638=>"111011001",
  40639=>"000000001",
  40640=>"001000110",
  40641=>"000000000",
  40642=>"101000011",
  40643=>"110111001",
  40644=>"011000000",
  40645=>"110011001",
  40646=>"010001111",
  40647=>"000111111",
  40648=>"111100111",
  40649=>"011011000",
  40650=>"101101010",
  40651=>"100100101",
  40652=>"000011000",
  40653=>"101110110",
  40654=>"000010111",
  40655=>"111111111",
  40656=>"001101111",
  40657=>"101011011",
  40658=>"000000000",
  40659=>"101101001",
  40660=>"111011001",
  40661=>"001000100",
  40662=>"111001101",
  40663=>"000010101",
  40664=>"001000000",
  40665=>"000000111",
  40666=>"101000100",
  40667=>"111000101",
  40668=>"111100000",
  40669=>"111011111",
  40670=>"111101000",
  40671=>"010111011",
  40672=>"110000000",
  40673=>"001000000",
  40674=>"011011011",
  40675=>"111100001",
  40676=>"001011011",
  40677=>"101111110",
  40678=>"111000000",
  40679=>"000001010",
  40680=>"110110000",
  40681=>"000110110",
  40682=>"100000001",
  40683=>"101001000",
  40684=>"000010100",
  40685=>"110110110",
  40686=>"100000101",
  40687=>"110111111",
  40688=>"110010010",
  40689=>"111111110",
  40690=>"000001100",
  40691=>"111110000",
  40692=>"100100001",
  40693=>"000011000",
  40694=>"000010011",
  40695=>"100010111",
  40696=>"111001110",
  40697=>"101001111",
  40698=>"111101000",
  40699=>"001010000",
  40700=>"100101101",
  40701=>"011010111",
  40702=>"011001001",
  40703=>"110000000",
  40704=>"000000000",
  40705=>"000001010",
  40706=>"000000001",
  40707=>"111111101",
  40708=>"111111111",
  40709=>"111011011",
  40710=>"000000010",
  40711=>"000000000",
  40712=>"110000000",
  40713=>"000001101",
  40714=>"111110000",
  40715=>"010110111",
  40716=>"000000001",
  40717=>"111111111",
  40718=>"110000000",
  40719=>"000000000",
  40720=>"010010010",
  40721=>"110110111",
  40722=>"001111000",
  40723=>"000101111",
  40724=>"000100000",
  40725=>"111111111",
  40726=>"000000001",
  40727=>"000000000",
  40728=>"100111000",
  40729=>"111110000",
  40730=>"110000110",
  40731=>"000000010",
  40732=>"001001111",
  40733=>"000101101",
  40734=>"000001000",
  40735=>"000000100",
  40736=>"000000000",
  40737=>"111111000",
  40738=>"000000101",
  40739=>"100001111",
  40740=>"100100101",
  40741=>"111111111",
  40742=>"111111001",
  40743=>"000000111",
  40744=>"110110010",
  40745=>"000010000",
  40746=>"000000000",
  40747=>"010110100",
  40748=>"000000010",
  40749=>"111000000",
  40750=>"111110000",
  40751=>"001000001",
  40752=>"000000000",
  40753=>"100111110",
  40754=>"100001000",
  40755=>"110111111",
  40756=>"110010110",
  40757=>"000000011",
  40758=>"100000110",
  40759=>"000000101",
  40760=>"111011000",
  40761=>"000000000",
  40762=>"000000000",
  40763=>"110111111",
  40764=>"111011011",
  40765=>"111111011",
  40766=>"000000100",
  40767=>"111011011",
  40768=>"110111110",
  40769=>"111111100",
  40770=>"110111111",
  40771=>"001010110",
  40772=>"000000011",
  40773=>"000110111",
  40774=>"000000000",
  40775=>"000000111",
  40776=>"001101100",
  40777=>"111111000",
  40778=>"000000000",
  40779=>"111111111",
  40780=>"010011010",
  40781=>"111111110",
  40782=>"001111111",
  40783=>"000000001",
  40784=>"111001111",
  40785=>"110110010",
  40786=>"000100111",
  40787=>"001000001",
  40788=>"010000000",
  40789=>"001101101",
  40790=>"001000000",
  40791=>"111110100",
  40792=>"000000001",
  40793=>"000000011",
  40794=>"111111110",
  40795=>"010110000",
  40796=>"111111000",
  40797=>"001001000",
  40798=>"111111110",
  40799=>"001011111",
  40800=>"111111000",
  40801=>"000000000",
  40802=>"001001101",
  40803=>"111111000",
  40804=>"110110000",
  40805=>"110010000",
  40806=>"000110000",
  40807=>"000010001",
  40808=>"000000111",
  40809=>"000111010",
  40810=>"110111111",
  40811=>"111111010",
  40812=>"000000001",
  40813=>"110010000",
  40814=>"000000001",
  40815=>"110010010",
  40816=>"001110110",
  40817=>"111111000",
  40818=>"010100110",
  40819=>"000110111",
  40820=>"001111111",
  40821=>"000000001",
  40822=>"111110100",
  40823=>"111111000",
  40824=>"111111010",
  40825=>"000110010",
  40826=>"001001001",
  40827=>"111111111",
  40828=>"110000100",
  40829=>"100100000",
  40830=>"000000010",
  40831=>"101000100",
  40832=>"001001000",
  40833=>"101000000",
  40834=>"010011000",
  40835=>"011100101",
  40836=>"111001010",
  40837=>"000001000",
  40838=>"110110110",
  40839=>"110110111",
  40840=>"011011011",
  40841=>"000000000",
  40842=>"010111011",
  40843=>"110111111",
  40844=>"110111010",
  40845=>"000001001",
  40846=>"000000000",
  40847=>"001000000",
  40848=>"111111111",
  40849=>"110010011",
  40850=>"111000010",
  40851=>"000010000",
  40852=>"110110110",
  40853=>"001000000",
  40854=>"010110001",
  40855=>"110010110",
  40856=>"011111000",
  40857=>"000000001",
  40858=>"111111110",
  40859=>"000001110",
  40860=>"000000000",
  40861=>"110110000",
  40862=>"100101000",
  40863=>"000000000",
  40864=>"001001001",
  40865=>"010110010",
  40866=>"110111010",
  40867=>"000000001",
  40868=>"110000001",
  40869=>"000000000",
  40870=>"111011111",
  40871=>"000111110",
  40872=>"110110001",
  40873=>"000111111",
  40874=>"001001100",
  40875=>"100101110",
  40876=>"000000000",
  40877=>"111110110",
  40878=>"000000000",
  40879=>"111001111",
  40880=>"111111010",
  40881=>"010110100",
  40882=>"111111011",
  40883=>"000100101",
  40884=>"110101111",
  40885=>"000000000",
  40886=>"111010101",
  40887=>"111111111",
  40888=>"111100101",
  40889=>"111111101",
  40890=>"111111011",
  40891=>"110111110",
  40892=>"000111110",
  40893=>"011111111",
  40894=>"101100100",
  40895=>"110110000",
  40896=>"111010000",
  40897=>"001001000",
  40898=>"110000100",
  40899=>"100100110",
  40900=>"110000000",
  40901=>"100100000",
  40902=>"000000000",
  40903=>"111111000",
  40904=>"110001111",
  40905=>"111111000",
  40906=>"101001000",
  40907=>"000000101",
  40908=>"010111110",
  40909=>"011010111",
  40910=>"010111110",
  40911=>"101101011",
  40912=>"000000010",
  40913=>"101110110",
  40914=>"111110010",
  40915=>"000000010",
  40916=>"111010000",
  40917=>"001101001",
  40918=>"000000101",
  40919=>"000001000",
  40920=>"000000000",
  40921=>"111101111",
  40922=>"000001100",
  40923=>"001001111",
  40924=>"101111100",
  40925=>"101111111",
  40926=>"010110000",
  40927=>"111111111",
  40928=>"111000111",
  40929=>"110000000",
  40930=>"011110111",
  40931=>"000000010",
  40932=>"110110010",
  40933=>"101111111",
  40934=>"100100111",
  40935=>"010000000",
  40936=>"111111011",
  40937=>"010000110",
  40938=>"111011000",
  40939=>"001000000",
  40940=>"110110110",
  40941=>"111111111",
  40942=>"110010001",
  40943=>"001001000",
  40944=>"000001111",
  40945=>"011010100",
  40946=>"000000111",
  40947=>"001001111",
  40948=>"000001001",
  40949=>"110111110",
  40950=>"110110100",
  40951=>"000001011",
  40952=>"011011000",
  40953=>"000110110",
  40954=>"000000000",
  40955=>"010010010",
  40956=>"111010000",
  40957=>"101101100",
  40958=>"100110110",
  40959=>"000000000",
  40960=>"100101111",
  40961=>"101101000",
  40962=>"000000000",
  40963=>"011000000",
  40964=>"010010011",
  40965=>"111100100",
  40966=>"010011111",
  40967=>"011111000",
  40968=>"010000101",
  40969=>"000101000",
  40970=>"010111000",
  40971=>"101000000",
  40972=>"101000000",
  40973=>"000000110",
  40974=>"100000111",
  40975=>"111110010",
  40976=>"100111011",
  40977=>"100111111",
  40978=>"000000101",
  40979=>"000000000",
  40980=>"001000000",
  40981=>"111100000",
  40982=>"110101000",
  40983=>"010111111",
  40984=>"111001000",
  40985=>"111111111",
  40986=>"110100101",
  40987=>"011101101",
  40988=>"110000000",
  40989=>"011111110",
  40990=>"111111100",
  40991=>"000000110",
  40992=>"111001001",
  40993=>"010000000",
  40994=>"000010010",
  40995=>"111001101",
  40996=>"000000011",
  40997=>"001111001",
  40998=>"111010000",
  40999=>"000101101",
  41000=>"000000000",
  41001=>"111111111",
  41002=>"100111000",
  41003=>"000000101",
  41004=>"011111000",
  41005=>"000101000",
  41006=>"111101000",
  41007=>"111111111",
  41008=>"111010001",
  41009=>"010000111",
  41010=>"101101001",
  41011=>"010011010",
  41012=>"000000000",
  41013=>"000111111",
  41014=>"111110111",
  41015=>"010111111",
  41016=>"101000000",
  41017=>"000000010",
  41018=>"000000000",
  41019=>"000010111",
  41020=>"100110001",
  41021=>"010111010",
  41022=>"010000011",
  41023=>"100000111",
  41024=>"111101100",
  41025=>"111010001",
  41026=>"101101111",
  41027=>"001100111",
  41028=>"100111010",
  41029=>"000101111",
  41030=>"011011011",
  41031=>"000001111",
  41032=>"010000001",
  41033=>"000000111",
  41034=>"001000000",
  41035=>"101000000",
  41036=>"000111000",
  41037=>"110011000",
  41038=>"111111111",
  41039=>"000010011",
  41040=>"111000000",
  41041=>"010111000",
  41042=>"011010000",
  41043=>"111000111",
  41044=>"111111000",
  41045=>"001000001",
  41046=>"000000110",
  41047=>"000111100",
  41048=>"100011010",
  41049=>"010010010",
  41050=>"000110010",
  41051=>"100000110",
  41052=>"111110000",
  41053=>"100100000",
  41054=>"000111111",
  41055=>"100001111",
  41056=>"111101111",
  41057=>"111000000",
  41058=>"000010000",
  41059=>"000010110",
  41060=>"110000000",
  41061=>"011011111",
  41062=>"100000111",
  41063=>"001111111",
  41064=>"000100101",
  41065=>"101111111",
  41066=>"111001101",
  41067=>"010010111",
  41068=>"010000000",
  41069=>"000111011",
  41070=>"101000000",
  41071=>"100000010",
  41072=>"000000011",
  41073=>"010000111",
  41074=>"111111011",
  41075=>"000111000",
  41076=>"111010011",
  41077=>"101000101",
  41078=>"000000000",
  41079=>"000000000",
  41080=>"000100000",
  41081=>"111111000",
  41082=>"000111111",
  41083=>"111000000",
  41084=>"000100001",
  41085=>"111101111",
  41086=>"000100111",
  41087=>"101000000",
  41088=>"011001000",
  41089=>"000000000",
  41090=>"111111010",
  41091=>"011010111",
  41092=>"111111000",
  41093=>"010001000",
  41094=>"110111100",
  41095=>"110011110",
  41096=>"110010000",
  41097=>"000000111",
  41098=>"111111100",
  41099=>"000100111",
  41100=>"000101010",
  41101=>"001100101",
  41102=>"101000100",
  41103=>"001000010",
  41104=>"111001111",
  41105=>"100100000",
  41106=>"110000001",
  41107=>"011000010",
  41108=>"100000110",
  41109=>"000000010",
  41110=>"000110010",
  41111=>"011011111",
  41112=>"111111111",
  41113=>"100111001",
  41114=>"101011000",
  41115=>"110101111",
  41116=>"010000010",
  41117=>"001111111",
  41118=>"010000111",
  41119=>"001000000",
  41120=>"000000100",
  41121=>"000100111",
  41122=>"111000101",
  41123=>"111010000",
  41124=>"000000101",
  41125=>"111000011",
  41126=>"011000000",
  41127=>"000000000",
  41128=>"011111110",
  41129=>"000000000",
  41130=>"111100100",
  41131=>"101000000",
  41132=>"001000001",
  41133=>"000000001",
  41134=>"010010110",
  41135=>"000001011",
  41136=>"011000100",
  41137=>"001110111",
  41138=>"111101100",
  41139=>"000100100",
  41140=>"100100101",
  41141=>"010001110",
  41142=>"111000000",
  41143=>"000010101",
  41144=>"000010110",
  41145=>"001000011",
  41146=>"111111000",
  41147=>"110110111",
  41148=>"000000011",
  41149=>"000111111",
  41150=>"101111011",
  41151=>"000100000",
  41152=>"000000010",
  41153=>"000010011",
  41154=>"000000111",
  41155=>"010001101",
  41156=>"000000101",
  41157=>"000011101",
  41158=>"111010000",
  41159=>"000000111",
  41160=>"111000010",
  41161=>"111101101",
  41162=>"111011011",
  41163=>"001000101",
  41164=>"011100111",
  41165=>"000011000",
  41166=>"010111111",
  41167=>"111111111",
  41168=>"001111111",
  41169=>"111011011",
  41170=>"000010111",
  41171=>"111100000",
  41172=>"000000111",
  41173=>"000111000",
  41174=>"000000000",
  41175=>"111110111",
  41176=>"000000010",
  41177=>"000000001",
  41178=>"011100001",
  41179=>"101000011",
  41180=>"101100000",
  41181=>"000101111",
  41182=>"101000101",
  41183=>"000000111",
  41184=>"111000101",
  41185=>"000000101",
  41186=>"000101101",
  41187=>"111100111",
  41188=>"000000101",
  41189=>"010000111",
  41190=>"111000000",
  41191=>"100001001",
  41192=>"111000000",
  41193=>"111111000",
  41194=>"011111100",
  41195=>"111111111",
  41196=>"000000100",
  41197=>"000111000",
  41198=>"000000001",
  41199=>"111000000",
  41200=>"000111001",
  41201=>"010110000",
  41202=>"000000100",
  41203=>"010011001",
  41204=>"111110111",
  41205=>"101111010",
  41206=>"100011010",
  41207=>"111001101",
  41208=>"000000010",
  41209=>"000001000",
  41210=>"111111111",
  41211=>"010111111",
  41212=>"111111100",
  41213=>"000001111",
  41214=>"100000011",
  41215=>"111000000",
  41216=>"101100100",
  41217=>"001110010",
  41218=>"000001111",
  41219=>"111000110",
  41220=>"111101101",
  41221=>"100001110",
  41222=>"000100111",
  41223=>"000010000",
  41224=>"111010010",
  41225=>"100101111",
  41226=>"101100101",
  41227=>"000100000",
  41228=>"000101110",
  41229=>"110010000",
  41230=>"000000000",
  41231=>"000111111",
  41232=>"111000111",
  41233=>"100100111",
  41234=>"111111011",
  41235=>"000000000",
  41236=>"101101111",
  41237=>"011011100",
  41238=>"011111011",
  41239=>"110110000",
  41240=>"101111000",
  41241=>"000000100",
  41242=>"110001000",
  41243=>"000101111",
  41244=>"110000010",
  41245=>"000000000",
  41246=>"111000000",
  41247=>"000000000",
  41248=>"100001111",
  41249=>"011111000",
  41250=>"110000100",
  41251=>"010010000",
  41252=>"001001001",
  41253=>"111011111",
  41254=>"010110000",
  41255=>"100001000",
  41256=>"111001000",
  41257=>"000000000",
  41258=>"000101111",
  41259=>"010011000",
  41260=>"101111001",
  41261=>"011000000",
  41262=>"111010000",
  41263=>"000010101",
  41264=>"100101010",
  41265=>"111011101",
  41266=>"101010001",
  41267=>"101000000",
  41268=>"110101111",
  41269=>"010110111",
  41270=>"111001101",
  41271=>"100000000",
  41272=>"101100111",
  41273=>"000000111",
  41274=>"101001000",
  41275=>"101100000",
  41276=>"111111001",
  41277=>"111010111",
  41278=>"001000101",
  41279=>"101000000",
  41280=>"100010111",
  41281=>"101101011",
  41282=>"101101001",
  41283=>"111101100",
  41284=>"100101111",
  41285=>"111000100",
  41286=>"001001000",
  41287=>"011100100",
  41288=>"111110010",
  41289=>"111101100",
  41290=>"001000111",
  41291=>"011010111",
  41292=>"000000000",
  41293=>"111100010",
  41294=>"111100110",
  41295=>"101010111",
  41296=>"111101101",
  41297=>"011111111",
  41298=>"111101110",
  41299=>"010001000",
  41300=>"000010001",
  41301=>"010010000",
  41302=>"111100000",
  41303=>"101000111",
  41304=>"001010000",
  41305=>"000001001",
  41306=>"000000000",
  41307=>"101011100",
  41308=>"000000001",
  41309=>"011001000",
  41310=>"011111111",
  41311=>"100101001",
  41312=>"010010000",
  41313=>"010010101",
  41314=>"001101111",
  41315=>"110010000",
  41316=>"101001000",
  41317=>"100101101",
  41318=>"111110000",
  41319=>"000000111",
  41320=>"010010000",
  41321=>"111111000",
  41322=>"101111110",
  41323=>"110000110",
  41324=>"100010000",
  41325=>"001101001",
  41326=>"011010010",
  41327=>"101111000",
  41328=>"101100000",
  41329=>"001101000",
  41330=>"111100000",
  41331=>"000000101",
  41332=>"101010000",
  41333=>"000000110",
  41334=>"001101110",
  41335=>"000000000",
  41336=>"000010000",
  41337=>"000000001",
  41338=>"101100111",
  41339=>"000101001",
  41340=>"100001100",
  41341=>"010010000",
  41342=>"010111100",
  41343=>"100101101",
  41344=>"111101001",
  41345=>"101100000",
  41346=>"100000001",
  41347=>"100010111",
  41348=>"111000100",
  41349=>"000000101",
  41350=>"100100010",
  41351=>"000000100",
  41352=>"101100011",
  41353=>"001100111",
  41354=>"101000101",
  41355=>"000100111",
  41356=>"011111101",
  41357=>"111111101",
  41358=>"000111101",
  41359=>"000000000",
  41360=>"111001000",
  41361=>"000000000",
  41362=>"010000000",
  41363=>"010110000",
  41364=>"111100000",
  41365=>"101001111",
  41366=>"111000101",
  41367=>"111001000",
  41368=>"011000011",
  41369=>"011010011",
  41370=>"101100101",
  41371=>"000000001",
  41372=>"001100010",
  41373=>"000000111",
  41374=>"100100011",
  41375=>"000101100",
  41376=>"011011001",
  41377=>"100010011",
  41378=>"011111000",
  41379=>"000011111",
  41380=>"001011000",
  41381=>"101100001",
  41382=>"111001101",
  41383=>"011011000",
  41384=>"011101100",
  41385=>"010100000",
  41386=>"000101111",
  41387=>"101000111",
  41388=>"011111000",
  41389=>"101101111",
  41390=>"011011001",
  41391=>"000000111",
  41392=>"010010111",
  41393=>"110000000",
  41394=>"100101000",
  41395=>"100001000",
  41396=>"111011000",
  41397=>"010010100",
  41398=>"111100100",
  41399=>"110100000",
  41400=>"011111110",
  41401=>"110001000",
  41402=>"111010110",
  41403=>"011000101",
  41404=>"111110101",
  41405=>"101111101",
  41406=>"111000000",
  41407=>"010000000",
  41408=>"001100000",
  41409=>"000000111",
  41410=>"111111000",
  41411=>"100101100",
  41412=>"000000100",
  41413=>"111111100",
  41414=>"100011011",
  41415=>"101101111",
  41416=>"010010101",
  41417=>"001010100",
  41418=>"000000000",
  41419=>"111010110",
  41420=>"100101111",
  41421=>"111110001",
  41422=>"000101110",
  41423=>"001010011",
  41424=>"000000111",
  41425=>"111100000",
  41426=>"000000000",
  41427=>"001010000",
  41428=>"000000111",
  41429=>"110110000",
  41430=>"111000000",
  41431=>"001000101",
  41432=>"010011100",
  41433=>"111111110",
  41434=>"100110100",
  41435=>"000100111",
  41436=>"110100000",
  41437=>"011011001",
  41438=>"111101101",
  41439=>"101101001",
  41440=>"100101100",
  41441=>"000000011",
  41442=>"110010101",
  41443=>"111101001",
  41444=>"101000001",
  41445=>"111111000",
  41446=>"100101110",
  41447=>"000110000",
  41448=>"101101111",
  41449=>"000010000",
  41450=>"101100110",
  41451=>"111000101",
  41452=>"000010110",
  41453=>"101100111",
  41454=>"100111010",
  41455=>"101111000",
  41456=>"100000000",
  41457=>"111011000",
  41458=>"101101010",
  41459=>"110110000",
  41460=>"111000100",
  41461=>"000001101",
  41462=>"010000111",
  41463=>"000111000",
  41464=>"100111011",
  41465=>"100010000",
  41466=>"111011001",
  41467=>"101111000",
  41468=>"000101111",
  41469=>"000010110",
  41470=>"100000101",
  41471=>"000101111",
  41472=>"011001100",
  41473=>"111111101",
  41474=>"000000000",
  41475=>"001000000",
  41476=>"100011011",
  41477=>"111000111",
  41478=>"111111111",
  41479=>"011111111",
  41480=>"111111111",
  41481=>"001000111",
  41482=>"001000001",
  41483=>"011101001",
  41484=>"000010000",
  41485=>"101001001",
  41486=>"000000100",
  41487=>"001011011",
  41488=>"101000111",
  41489=>"001000111",
  41490=>"111001111",
  41491=>"111100000",
  41492=>"111111000",
  41493=>"001101111",
  41494=>"100011001",
  41495=>"111111010",
  41496=>"101101111",
  41497=>"100111110",
  41498=>"110010111",
  41499=>"000000101",
  41500=>"000000001",
  41501=>"111101000",
  41502=>"110101111",
  41503=>"000000000",
  41504=>"000000000",
  41505=>"011111011",
  41506=>"000011110",
  41507=>"001011010",
  41508=>"111111001",
  41509=>"011001001",
  41510=>"000111111",
  41511=>"101010011",
  41512=>"010010000",
  41513=>"110111111",
  41514=>"101100111",
  41515=>"010010000",
  41516=>"111111111",
  41517=>"001111011",
  41518=>"110000010",
  41519=>"111000111",
  41520=>"111111010",
  41521=>"111111000",
  41522=>"000010111",
  41523=>"111101101",
  41524=>"000000000",
  41525=>"100110001",
  41526=>"111011000",
  41527=>"100001000",
  41528=>"011010000",
  41529=>"000000111",
  41530=>"001000111",
  41531=>"101111110",
  41532=>"001000000",
  41533=>"111010000",
  41534=>"000000001",
  41535=>"110011011",
  41536=>"111111111",
  41537=>"001101101",
  41538=>"111000000",
  41539=>"011000000",
  41540=>"111111010",
  41541=>"001000000",
  41542=>"100100000",
  41543=>"111011111",
  41544=>"111011111",
  41545=>"001101111",
  41546=>"101000101",
  41547=>"101110000",
  41548=>"000000000",
  41549=>"000110110",
  41550=>"101110010",
  41551=>"100011000",
  41552=>"000100100",
  41553=>"111111111",
  41554=>"111000111",
  41555=>"011000000",
  41556=>"000000111",
  41557=>"100110110",
  41558=>"001010000",
  41559=>"000000000",
  41560=>"000100101",
  41561=>"110001001",
  41562=>"000110110",
  41563=>"000011011",
  41564=>"111110111",
  41565=>"100000110",
  41566=>"111111110",
  41567=>"100000000",
  41568=>"000000000",
  41569=>"010000101",
  41570=>"000000000",
  41571=>"001001001",
  41572=>"001000001",
  41573=>"011001000",
  41574=>"000001101",
  41575=>"000000101",
  41576=>"111111000",
  41577=>"111000100",
  41578=>"010110111",
  41579=>"111010111",
  41580=>"001001011",
  41581=>"000000101",
  41582=>"101101110",
  41583=>"000101011",
  41584=>"111111100",
  41585=>"111000011",
  41586=>"011011000",
  41587=>"000000000",
  41588=>"000011000",
  41589=>"111000100",
  41590=>"111001011",
  41591=>"111111110",
  41592=>"000000000",
  41593=>"100001001",
  41594=>"000010111",
  41595=>"000111110",
  41596=>"000011001",
  41597=>"110000011",
  41598=>"011010000",
  41599=>"000000000",
  41600=>"111011100",
  41601=>"000010001",
  41602=>"101101101",
  41603=>"100111001",
  41604=>"101000011",
  41605=>"111111000",
  41606=>"110100100",
  41607=>"100001110",
  41608=>"100111001",
  41609=>"000000000",
  41610=>"100000000",
  41611=>"111010111",
  41612=>"011000000",
  41613=>"100011111",
  41614=>"111000000",
  41615=>"000000000",
  41616=>"010110101",
  41617=>"000000000",
  41618=>"111000010",
  41619=>"111111110",
  41620=>"010110100",
  41621=>"111000111",
  41622=>"111001110",
  41623=>"100111111",
  41624=>"101011000",
  41625=>"111101001",
  41626=>"010011010",
  41627=>"010000101",
  41628=>"000000110",
  41629=>"111100001",
  41630=>"111000100",
  41631=>"011000111",
  41632=>"001011111",
  41633=>"010000111",
  41634=>"000111010",
  41635=>"000000000",
  41636=>"111111111",
  41637=>"000100110",
  41638=>"101110100",
  41639=>"000000111",
  41640=>"110101000",
  41641=>"000000001",
  41642=>"010000000",
  41643=>"000000111",
  41644=>"101111010",
  41645=>"000000111",
  41646=>"000000001",
  41647=>"010000001",
  41648=>"001011001",
  41649=>"111111111",
  41650=>"010000000",
  41651=>"001000011",
  41652=>"101001011",
  41653=>"101011000",
  41654=>"111001101",
  41655=>"001111000",
  41656=>"000000000",
  41657=>"111011001",
  41658=>"000000000",
  41659=>"111000000",
  41660=>"000000001",
  41661=>"110111110",
  41662=>"110111000",
  41663=>"000000000",
  41664=>"000000111",
  41665=>"101000000",
  41666=>"110111001",
  41667=>"110001000",
  41668=>"010111101",
  41669=>"101111111",
  41670=>"001000000",
  41671=>"110010000",
  41672=>"111111100",
  41673=>"000011000",
  41674=>"010011000",
  41675=>"101111000",
  41676=>"011101101",
  41677=>"000010110",
  41678=>"101101101",
  41679=>"111010011",
  41680=>"111000000",
  41681=>"000111011",
  41682=>"001000000",
  41683=>"001111011",
  41684=>"000000000",
  41685=>"011001001",
  41686=>"000000000",
  41687=>"011000100",
  41688=>"111111000",
  41689=>"000110000",
  41690=>"100110010",
  41691=>"110000101",
  41692=>"000000110",
  41693=>"111000101",
  41694=>"010100000",
  41695=>"111111000",
  41696=>"100000000",
  41697=>"000000011",
  41698=>"111010010",
  41699=>"001111111",
  41700=>"000000001",
  41701=>"000111000",
  41702=>"010111101",
  41703=>"000001100",
  41704=>"011000111",
  41705=>"000001000",
  41706=>"100000100",
  41707=>"000110000",
  41708=>"111111001",
  41709=>"010000110",
  41710=>"010000000",
  41711=>"000011010",
  41712=>"001111000",
  41713=>"111011111",
  41714=>"111111111",
  41715=>"111110110",
  41716=>"110011111",
  41717=>"101101101",
  41718=>"000000101",
  41719=>"001000000",
  41720=>"001111010",
  41721=>"000110111",
  41722=>"110011000",
  41723=>"000011111",
  41724=>"010010000",
  41725=>"111011111",
  41726=>"001011111",
  41727=>"110110111",
  41728=>"111010000",
  41729=>"000000111",
  41730=>"101000001",
  41731=>"111000101",
  41732=>"011101111",
  41733=>"101000000",
  41734=>"010011011",
  41735=>"001000101",
  41736=>"011110111",
  41737=>"111011001",
  41738=>"010000111",
  41739=>"101001101",
  41740=>"000010000",
  41741=>"101100000",
  41742=>"100011011",
  41743=>"011111001",
  41744=>"000010110",
  41745=>"010000000",
  41746=>"000001000",
  41747=>"000000110",
  41748=>"111111101",
  41749=>"011000000",
  41750=>"100100111",
  41751=>"000000110",
  41752=>"000001101",
  41753=>"101011101",
  41754=>"111111010",
  41755=>"111111000",
  41756=>"110110101",
  41757=>"000000000",
  41758=>"110010000",
  41759=>"011000000",
  41760=>"000110000",
  41761=>"000111011",
  41762=>"000111011",
  41763=>"111000000",
  41764=>"110111000",
  41765=>"110110000",
  41766=>"000000000",
  41767=>"111111111",
  41768=>"110110111",
  41769=>"110111111",
  41770=>"000100111",
  41771=>"011000000",
  41772=>"000011011",
  41773=>"101010011",
  41774=>"111111111",
  41775=>"000000000",
  41776=>"111000000",
  41777=>"000100000",
  41778=>"000000110",
  41779=>"001110111",
  41780=>"110000000",
  41781=>"111111000",
  41782=>"100011011",
  41783=>"000000101",
  41784=>"010000000",
  41785=>"101000001",
  41786=>"011000101",
  41787=>"000000010",
  41788=>"110110110",
  41789=>"010111110",
  41790=>"000010000",
  41791=>"110011010",
  41792=>"001101111",
  41793=>"111010001",
  41794=>"000000101",
  41795=>"000110110",
  41796=>"000111111",
  41797=>"101000110",
  41798=>"011111000",
  41799=>"111000000",
  41800=>"000001000",
  41801=>"011000111",
  41802=>"101000001",
  41803=>"111111100",
  41804=>"010010110",
  41805=>"001001000",
  41806=>"000101100",
  41807=>"010111110",
  41808=>"101000000",
  41809=>"000000001",
  41810=>"111101111",
  41811=>"011100100",
  41812=>"111111111",
  41813=>"000110110",
  41814=>"111011001",
  41815=>"111010000",
  41816=>"111100011",
  41817=>"100110110",
  41818=>"001110000",
  41819=>"111111000",
  41820=>"000110111",
  41821=>"111001000",
  41822=>"011111011",
  41823=>"000011011",
  41824=>"000111111",
  41825=>"001010000",
  41826=>"111110101",
  41827=>"000111111",
  41828=>"111111000",
  41829=>"011001000",
  41830=>"101111111",
  41831=>"011001001",
  41832=>"000000001",
  41833=>"011010001",
  41834=>"110010111",
  41835=>"000101101",
  41836=>"011000110",
  41837=>"101000111",
  41838=>"011001000",
  41839=>"111010111",
  41840=>"000101000",
  41841=>"010010111",
  41842=>"001100100",
  41843=>"110000000",
  41844=>"000100111",
  41845=>"000000101",
  41846=>"000000000",
  41847=>"111111111",
  41848=>"000111111",
  41849=>"111001001",
  41850=>"000101111",
  41851=>"100000000",
  41852=>"000110110",
  41853=>"110100000",
  41854=>"011101000",
  41855=>"011000000",
  41856=>"001000000",
  41857=>"010000000",
  41858=>"111111000",
  41859=>"111110101",
  41860=>"011111111",
  41861=>"110111000",
  41862=>"110011000",
  41863=>"001010000",
  41864=>"100101100",
  41865=>"010000000",
  41866=>"000000000",
  41867=>"101000000",
  41868=>"000111001",
  41869=>"011111110",
  41870=>"010010010",
  41871=>"000001000",
  41872=>"001001000",
  41873=>"010010000",
  41874=>"011001101",
  41875=>"011001111",
  41876=>"000011111",
  41877=>"000010111",
  41878=>"111101111",
  41879=>"000011011",
  41880=>"000000000",
  41881=>"001010111",
  41882=>"000111111",
  41883=>"000000101",
  41884=>"000010000",
  41885=>"010111110",
  41886=>"000000110",
  41887=>"000000100",
  41888=>"000000000",
  41889=>"000010000",
  41890=>"000000000",
  41891=>"111111101",
  41892=>"111010000",
  41893=>"000000000",
  41894=>"101111111",
  41895=>"110111000",
  41896=>"001000010",
  41897=>"000111000",
  41898=>"111110101",
  41899=>"000000000",
  41900=>"101001111",
  41901=>"101001000",
  41902=>"110000000",
  41903=>"101110011",
  41904=>"000101000",
  41905=>"101011100",
  41906=>"000000010",
  41907=>"001100100",
  41908=>"111101000",
  41909=>"101010010",
  41910=>"111101100",
  41911=>"111111010",
  41912=>"001011010",
  41913=>"000100111",
  41914=>"000100101",
  41915=>"111010011",
  41916=>"111111000",
  41917=>"000111111",
  41918=>"011111100",
  41919=>"111000000",
  41920=>"111010000",
  41921=>"111001000",
  41922=>"010101111",
  41923=>"000100100",
  41924=>"010000000",
  41925=>"000001001",
  41926=>"010001010",
  41927=>"000000000",
  41928=>"111101000",
  41929=>"000000000",
  41930=>"011001101",
  41931=>"000000001",
  41932=>"000000000",
  41933=>"000011011",
  41934=>"001101101",
  41935=>"000111100",
  41936=>"111001000",
  41937=>"111110100",
  41938=>"111000111",
  41939=>"000001001",
  41940=>"100010010",
  41941=>"111100000",
  41942=>"000000110",
  41943=>"010010110",
  41944=>"000001011",
  41945=>"000000111",
  41946=>"001000101",
  41947=>"001000101",
  41948=>"001011111",
  41949=>"100011000",
  41950=>"111111010",
  41951=>"100000110",
  41952=>"000010001",
  41953=>"111000111",
  41954=>"111101000",
  41955=>"111111100",
  41956=>"000010000",
  41957=>"000000111",
  41958=>"111000000",
  41959=>"011000000",
  41960=>"000000101",
  41961=>"001111111",
  41962=>"010000111",
  41963=>"001111110",
  41964=>"000000101",
  41965=>"000000000",
  41966=>"000010000",
  41967=>"000000000",
  41968=>"000000011",
  41969=>"000000110",
  41970=>"110000000",
  41971=>"011011001",
  41972=>"100111001",
  41973=>"000101000",
  41974=>"000000000",
  41975=>"000101111",
  41976=>"000010110",
  41977=>"101101111",
  41978=>"010111100",
  41979=>"000101011",
  41980=>"000010110",
  41981=>"000000001",
  41982=>"000100011",
  41983=>"000000000",
  41984=>"000001100",
  41985=>"000100101",
  41986=>"100100010",
  41987=>"111101111",
  41988=>"001101010",
  41989=>"100101100",
  41990=>"100010111",
  41991=>"011011111",
  41992=>"001001101",
  41993=>"100111111",
  41994=>"100100101",
  41995=>"000000011",
  41996=>"011011011",
  41997=>"011011001",
  41998=>"101101001",
  41999=>"000000001",
  42000=>"010011000",
  42001=>"110100000",
  42002=>"101000101",
  42003=>"100000010",
  42004=>"111000000",
  42005=>"111111111",
  42006=>"000011111",
  42007=>"100100000",
  42008=>"100100100",
  42009=>"000000001",
  42010=>"000011100",
  42011=>"100111011",
  42012=>"100110011",
  42013=>"000001111",
  42014=>"111001111",
  42015=>"011001000",
  42016=>"110010110",
  42017=>"000111110",
  42018=>"000011011",
  42019=>"000101111",
  42020=>"100100110",
  42021=>"110101011",
  42022=>"000100011",
  42023=>"100110110",
  42024=>"111111011",
  42025=>"011001010",
  42026=>"100100110",
  42027=>"000100101",
  42028=>"111011011",
  42029=>"101011111",
  42030=>"111000001",
  42031=>"000000100",
  42032=>"111101111",
  42033=>"111110110",
  42034=>"000001000",
  42035=>"000011001",
  42036=>"000000000",
  42037=>"011010011",
  42038=>"000101101",
  42039=>"011110000",
  42040=>"111101011",
  42041=>"000100100",
  42042=>"000000000",
  42043=>"100011011",
  42044=>"011011101",
  42045=>"011011001",
  42046=>"000000011",
  42047=>"101001011",
  42048=>"011011001",
  42049=>"000011001",
  42050=>"100110000",
  42051=>"000000101",
  42052=>"000000000",
  42053=>"011000000",
  42054=>"100100111",
  42055=>"110111011",
  42056=>"111110110",
  42057=>"001111000",
  42058=>"000110100",
  42059=>"011011001",
  42060=>"000000000",
  42061=>"011111111",
  42062=>"111001101",
  42063=>"111011001",
  42064=>"100100100",
  42065=>"000111111",
  42066=>"011000000",
  42067=>"000000000",
  42068=>"100010011",
  42069=>"110111111",
  42070=>"100100000",
  42071=>"100100100",
  42072=>"111011000",
  42073=>"010010011",
  42074=>"110000110",
  42075=>"011111100",
  42076=>"110111110",
  42077=>"000000000",
  42078=>"111100000",
  42079=>"110101100",
  42080=>"000110110",
  42081=>"010110100",
  42082=>"100110111",
  42083=>"100000101",
  42084=>"010000010",
  42085=>"000100100",
  42086=>"111111000",
  42087=>"111010011",
  42088=>"000111111",
  42089=>"110100001",
  42090=>"111010011",
  42091=>"011101000",
  42092=>"101111001",
  42093=>"111000000",
  42094=>"100110111",
  42095=>"011111000",
  42096=>"000111010",
  42097=>"100101000",
  42098=>"000110100",
  42099=>"011000100",
  42100=>"101100000",
  42101=>"100100000",
  42102=>"011011011",
  42103=>"011111101",
  42104=>"100100110",
  42105=>"000100000",
  42106=>"011110000",
  42107=>"110001111",
  42108=>"110010111",
  42109=>"110110111",
  42110=>"000011111",
  42111=>"100110011",
  42112=>"000100000",
  42113=>"100111111",
  42114=>"110110000",
  42115=>"011101000",
  42116=>"111011011",
  42117=>"000011111",
  42118=>"000100010",
  42119=>"000110001",
  42120=>"110101001",
  42121=>"001000100",
  42122=>"110110011",
  42123=>"000110000",
  42124=>"111011010",
  42125=>"111110111",
  42126=>"000000010",
  42127=>"000001010",
  42128=>"010000100",
  42129=>"000000011",
  42130=>"100110011",
  42131=>"010111101",
  42132=>"001001101",
  42133=>"100000111",
  42134=>"000001111",
  42135=>"001001000",
  42136=>"010100011",
  42137=>"000000011",
  42138=>"100100111",
  42139=>"100010010",
  42140=>"101100100",
  42141=>"000110111",
  42142=>"100110111",
  42143=>"000011000",
  42144=>"000011101",
  42145=>"000000000",
  42146=>"011000111",
  42147=>"000000010",
  42148=>"100000110",
  42149=>"011011000",
  42150=>"011101110",
  42151=>"000100100",
  42152=>"100000111",
  42153=>"011011101",
  42154=>"111101111",
  42155=>"000100111",
  42156=>"011001000",
  42157=>"100100100",
  42158=>"100101111",
  42159=>"000010111",
  42160=>"000111101",
  42161=>"000001101",
  42162=>"011001000",
  42163=>"100000000",
  42164=>"011011010",
  42165=>"011010111",
  42166=>"001000001",
  42167=>"001100110",
  42168=>"101010110",
  42169=>"011011111",
  42170=>"000011000",
  42171=>"110110000",
  42172=>"011001101",
  42173=>"111110111",
  42174=>"000000011",
  42175=>"001111101",
  42176=>"100111011",
  42177=>"100000111",
  42178=>"000111110",
  42179=>"100101100",
  42180=>"011000100",
  42181=>"110110000",
  42182=>"011001011",
  42183=>"100011011",
  42184=>"100000101",
  42185=>"011011011",
  42186=>"000000010",
  42187=>"011111011",
  42188=>"000010100",
  42189=>"001000111",
  42190=>"011011000",
  42191=>"011011000",
  42192=>"000101001",
  42193=>"011101001",
  42194=>"011011000",
  42195=>"011001110",
  42196=>"100110011",
  42197=>"010111100",
  42198=>"100111101",
  42199=>"100000111",
  42200=>"011100100",
  42201=>"011001000",
  42202=>"010001000",
  42203=>"100100100",
  42204=>"111110000",
  42205=>"001011101",
  42206=>"111000000",
  42207=>"111101011",
  42208=>"001111001",
  42209=>"100110101",
  42210=>"101001101",
  42211=>"100010110",
  42212=>"100100100",
  42213=>"110011010",
  42214=>"000111111",
  42215=>"100000000",
  42216=>"100011011",
  42217=>"110110000",
  42218=>"000000000",
  42219=>"000000100",
  42220=>"001011011",
  42221=>"100111000",
  42222=>"101001001",
  42223=>"000000011",
  42224=>"011011000",
  42225=>"111101101",
  42226=>"111011101",
  42227=>"111000100",
  42228=>"011111111",
  42229=>"100100100",
  42230=>"100000001",
  42231=>"110110000",
  42232=>"000000110",
  42233=>"111001000",
  42234=>"011001000",
  42235=>"011000001",
  42236=>"100100101",
  42237=>"000100001",
  42238=>"111011011",
  42239=>"100110111",
  42240=>"011010110",
  42241=>"010011101",
  42242=>"101000111",
  42243=>"110111011",
  42244=>"001001110",
  42245=>"110000111",
  42246=>"010111111",
  42247=>"001111111",
  42248=>"001101111",
  42249=>"000000111",
  42250=>"000100000",
  42251=>"110101000",
  42252=>"010000110",
  42253=>"000000110",
  42254=>"000000100",
  42255=>"001011000",
  42256=>"000110111",
  42257=>"000000011",
  42258=>"000000110",
  42259=>"011010000",
  42260=>"111011001",
  42261=>"111101101",
  42262=>"001011001",
  42263=>"111111101",
  42264=>"100000100",
  42265=>"101101101",
  42266=>"110101111",
  42267=>"101101101",
  42268=>"111010000",
  42269=>"000000000",
  42270=>"110010100",
  42271=>"000000000",
  42272=>"001101000",
  42273=>"011111011",
  42274=>"010101100",
  42275=>"010110000",
  42276=>"001110110",
  42277=>"111010001",
  42278=>"101000000",
  42279=>"000001110",
  42280=>"010011111",
  42281=>"000001001",
  42282=>"000000010",
  42283=>"000111000",
  42284=>"100111000",
  42285=>"101001101",
  42286=>"111011000",
  42287=>"001011000",
  42288=>"110010101",
  42289=>"000110010",
  42290=>"000100000",
  42291=>"111101000",
  42292=>"011000001",
  42293=>"010001001",
  42294=>"110110010",
  42295=>"010011001",
  42296=>"110010011",
  42297=>"000000000",
  42298=>"000000000",
  42299=>"111101000",
  42300=>"100000001",
  42301=>"111000000",
  42302=>"000000011",
  42303=>"000000000",
  42304=>"111101101",
  42305=>"111011000",
  42306=>"001100101",
  42307=>"011010000",
  42308=>"100010010",
  42309=>"000010000",
  42310=>"000101101",
  42311=>"000000111",
  42312=>"110111110",
  42313=>"010010000",
  42314=>"000001001",
  42315=>"111100111",
  42316=>"011000100",
  42317=>"110111011",
  42318=>"100101011",
  42319=>"111111100",
  42320=>"000111011",
  42321=>"000111111",
  42322=>"010010100",
  42323=>"011001010",
  42324=>"110001100",
  42325=>"100000100",
  42326=>"001011010",
  42327=>"100000110",
  42328=>"100110011",
  42329=>"000011011",
  42330=>"000000001",
  42331=>"011011111",
  42332=>"011000000",
  42333=>"000100110",
  42334=>"111010111",
  42335=>"100110101",
  42336=>"000000000",
  42337=>"100010010",
  42338=>"001000111",
  42339=>"000010100",
  42340=>"000001011",
  42341=>"011000000",
  42342=>"000011010",
  42343=>"000010111",
  42344=>"000000000",
  42345=>"111000100",
  42346=>"111010111",
  42347=>"111110110",
  42348=>"100111110",
  42349=>"001011111",
  42350=>"100101000",
  42351=>"110111111",
  42352=>"000101100",
  42353=>"010100101",
  42354=>"011011101",
  42355=>"000000101",
  42356=>"111100000",
  42357=>"100000101",
  42358=>"100111111",
  42359=>"001001001",
  42360=>"011000111",
  42361=>"010000000",
  42362=>"100101101",
  42363=>"000100010",
  42364=>"101001001",
  42365=>"100100010",
  42366=>"000000101",
  42367=>"000000111",
  42368=>"010111001",
  42369=>"011001000",
  42370=>"101011101",
  42371=>"000101111",
  42372=>"011000000",
  42373=>"101100101",
  42374=>"111010100",
  42375=>"101100110",
  42376=>"100110011",
  42377=>"010011101",
  42378=>"111111111",
  42379=>"010111100",
  42380=>"100101111",
  42381=>"100000001",
  42382=>"010010101",
  42383=>"000100111",
  42384=>"101011111",
  42385=>"001010000",
  42386=>"101101101",
  42387=>"001111000",
  42388=>"001100110",
  42389=>"010101110",
  42390=>"111111111",
  42391=>"000110110",
  42392=>"111110000",
  42393=>"101111000",
  42394=>"101011000",
  42395=>"101000111",
  42396=>"111100100",
  42397=>"111111010",
  42398=>"010010101",
  42399=>"001111010",
  42400=>"000001001",
  42401=>"000010011",
  42402=>"000001110",
  42403=>"111111100",
  42404=>"100001000",
  42405=>"100001011",
  42406=>"110110000",
  42407=>"010111110",
  42408=>"101011000",
  42409=>"010111101",
  42410=>"111001110",
  42411=>"000100010",
  42412=>"101111100",
  42413=>"000011111",
  42414=>"100110011",
  42415=>"110101111",
  42416=>"110000101",
  42417=>"111001001",
  42418=>"000010011",
  42419=>"001001011",
  42420=>"101111100",
  42421=>"111011011",
  42422=>"011101111",
  42423=>"000000010",
  42424=>"001000100",
  42425=>"101101001",
  42426=>"000010010",
  42427=>"010000111",
  42428=>"010000000",
  42429=>"111001011",
  42430=>"101100010",
  42431=>"000000000",
  42432=>"000010001",
  42433=>"100000000",
  42434=>"110010000",
  42435=>"000011000",
  42436=>"000001100",
  42437=>"000100110",
  42438=>"011010110",
  42439=>"000110111",
  42440=>"000000101",
  42441=>"010000001",
  42442=>"111111000",
  42443=>"000001111",
  42444=>"000100100",
  42445=>"000100100",
  42446=>"000001011",
  42447=>"000100000",
  42448=>"101010010",
  42449=>"001011011",
  42450=>"011111001",
  42451=>"000101111",
  42452=>"100000001",
  42453=>"101111001",
  42454=>"000000010",
  42455=>"111111111",
  42456=>"000000000",
  42457=>"001010000",
  42458=>"010110100",
  42459=>"101000101",
  42460=>"001101001",
  42461=>"111010100",
  42462=>"111101000",
  42463=>"010000001",
  42464=>"100000101",
  42465=>"111000011",
  42466=>"010000101",
  42467=>"000010010",
  42468=>"000000001",
  42469=>"111111000",
  42470=>"111001000",
  42471=>"000110110",
  42472=>"000000101",
  42473=>"000011000",
  42474=>"100111010",
  42475=>"010101010",
  42476=>"000000111",
  42477=>"111010100",
  42478=>"001000000",
  42479=>"011100110",
  42480=>"101100000",
  42481=>"001001011",
  42482=>"111011001",
  42483=>"001110110",
  42484=>"100110110",
  42485=>"000000100",
  42486=>"100000111",
  42487=>"000000100",
  42488=>"000111111",
  42489=>"000110111",
  42490=>"000111111",
  42491=>"100001000",
  42492=>"010100000",
  42493=>"000000000",
  42494=>"101011111",
  42495=>"001010000",
  42496=>"111111111",
  42497=>"000010010",
  42498=>"000000101",
  42499=>"000110101",
  42500=>"000001000",
  42501=>"001000100",
  42502=>"011111011",
  42503=>"111111000",
  42504=>"101000000",
  42505=>"000000001",
  42506=>"011011010",
  42507=>"111010101",
  42508=>"000000000",
  42509=>"000000100",
  42510=>"110100000",
  42511=>"111111111",
  42512=>"001000000",
  42513=>"011111110",
  42514=>"000111000",
  42515=>"010010010",
  42516=>"111111010",
  42517=>"100100111",
  42518=>"000011010",
  42519=>"000111011",
  42520=>"101100000",
  42521=>"111011011",
  42522=>"000101100",
  42523=>"000000000",
  42524=>"001111001",
  42525=>"000011111",
  42526=>"111101000",
  42527=>"000000000",
  42528=>"000100100",
  42529=>"000000000",
  42530=>"000000111",
  42531=>"010001001",
  42532=>"101111111",
  42533=>"100101000",
  42534=>"000010010",
  42535=>"100010000",
  42536=>"101111110",
  42537=>"111111000",
  42538=>"000000110",
  42539=>"001100000",
  42540=>"001111111",
  42541=>"011110000",
  42542=>"010000000",
  42543=>"101000100",
  42544=>"000011010",
  42545=>"010101000",
  42546=>"001101100",
  42547=>"011111001",
  42548=>"000111011",
  42549=>"111111011",
  42550=>"000011011",
  42551=>"100111010",
  42552=>"111100000",
  42553=>"000111111",
  42554=>"000000101",
  42555=>"011011011",
  42556=>"110010000",
  42557=>"111111011",
  42558=>"000000100",
  42559=>"000111111",
  42560=>"001011010",
  42561=>"101010100",
  42562=>"111000000",
  42563=>"111101111",
  42564=>"000000000",
  42565=>"101101111",
  42566=>"001111011",
  42567=>"011011111",
  42568=>"000000000",
  42569=>"000101100",
  42570=>"111111101",
  42571=>"110111111",
  42572=>"101111110",
  42573=>"001111101",
  42574=>"101001001",
  42575=>"111000000",
  42576=>"000000010",
  42577=>"111111111",
  42578=>"111011111",
  42579=>"001111000",
  42580=>"000000111",
  42581=>"100111100",
  42582=>"001111011",
  42583=>"011000000",
  42584=>"010011111",
  42585=>"010111010",
  42586=>"000111000",
  42587=>"000111010",
  42588=>"101101000",
  42589=>"110000000",
  42590=>"101111000",
  42591=>"111101001",
  42592=>"101000001",
  42593=>"000000000",
  42594=>"000000101",
  42595=>"011111100",
  42596=>"010000101",
  42597=>"010010010",
  42598=>"000000000",
  42599=>"110111010",
  42600=>"111111111",
  42601=>"011011110",
  42602=>"000000000",
  42603=>"100111011",
  42604=>"000001000",
  42605=>"000111000",
  42606=>"100000000",
  42607=>"101100000",
  42608=>"110110100",
  42609=>"010111110",
  42610=>"010010010",
  42611=>"111100000",
  42612=>"101111000",
  42613=>"000000111",
  42614=>"001011000",
  42615=>"000000011",
  42616=>"000111111",
  42617=>"000000000",
  42618=>"101011110",
  42619=>"111100000",
  42620=>"101101100",
  42621=>"101001000",
  42622=>"100000000",
  42623=>"111100101",
  42624=>"101100000",
  42625=>"111111111",
  42626=>"000000010",
  42627=>"000000011",
  42628=>"111101010",
  42629=>"010010111",
  42630=>"011111000",
  42631=>"000000000",
  42632=>"001011011",
  42633=>"111111000",
  42634=>"111100000",
  42635=>"111110000",
  42636=>"111100100",
  42637=>"111111111",
  42638=>"000111111",
  42639=>"100000000",
  42640=>"000110110",
  42641=>"000011010",
  42642=>"000000010",
  42643=>"100011010",
  42644=>"000011011",
  42645=>"101000000",
  42646=>"011011000",
  42647=>"111111100",
  42648=>"000000011",
  42649=>"011111111",
  42650=>"000011010",
  42651=>"101000110",
  42652=>"100111111",
  42653=>"000001000",
  42654=>"111010001",
  42655=>"010111111",
  42656=>"111000110",
  42657=>"101111001",
  42658=>"010101001",
  42659=>"000011011",
  42660=>"000111011",
  42661=>"010010011",
  42662=>"011101100",
  42663=>"000111110",
  42664=>"010000010",
  42665=>"011000001",
  42666=>"000000000",
  42667=>"000000111",
  42668=>"110000101",
  42669=>"000000101",
  42670=>"110111101",
  42671=>"111000000",
  42672=>"100100101",
  42673=>"010010000",
  42674=>"111111111",
  42675=>"011110110",
  42676=>"100111011",
  42677=>"000011010",
  42678=>"000000000",
  42679=>"000000000",
  42680=>"000011100",
  42681=>"000000010",
  42682=>"000000011",
  42683=>"000111001",
  42684=>"100011010",
  42685=>"111111111",
  42686=>"110100100",
  42687=>"000111011",
  42688=>"000000000",
  42689=>"000111000",
  42690=>"011111010",
  42691=>"010001001",
  42692=>"000111010",
  42693=>"111101011",
  42694=>"100010010",
  42695=>"000101111",
  42696=>"000010111",
  42697=>"100111111",
  42698=>"000010011",
  42699=>"000011000",
  42700=>"100101110",
  42701=>"111111010",
  42702=>"000011110",
  42703=>"110100100",
  42704=>"000111010",
  42705=>"111111101",
  42706=>"010000000",
  42707=>"111111000",
  42708=>"101000101",
  42709=>"000001000",
  42710=>"100000000",
  42711=>"000111000",
  42712=>"000011000",
  42713=>"000000100",
  42714=>"010111000",
  42715=>"010000000",
  42716=>"000111010",
  42717=>"000100100",
  42718=>"100000010",
  42719=>"000000000",
  42720=>"101000100",
  42721=>"001000000",
  42722=>"111111101",
  42723=>"000010000",
  42724=>"100000000",
  42725=>"111011000",
  42726=>"100111001",
  42727=>"001110110",
  42728=>"000001010",
  42729=>"010111000",
  42730=>"000111010",
  42731=>"010000011",
  42732=>"000000000",
  42733=>"100011000",
  42734=>"101101111",
  42735=>"011000101",
  42736=>"010111011",
  42737=>"011101111",
  42738=>"010000000",
  42739=>"100111100",
  42740=>"100101011",
  42741=>"011010000",
  42742=>"111000000",
  42743=>"110000111",
  42744=>"000111000",
  42745=>"011110010",
  42746=>"000011000",
  42747=>"101110100",
  42748=>"000111010",
  42749=>"111111000",
  42750=>"100111001",
  42751=>"010111000",
  42752=>"100001111",
  42753=>"110100110",
  42754=>"001011001",
  42755=>"000011101",
  42756=>"110111000",
  42757=>"001011000",
  42758=>"001000000",
  42759=>"100000000",
  42760=>"100110111",
  42761=>"011011001",
  42762=>"110100000",
  42763=>"100010100",
  42764=>"011011000",
  42765=>"000001111",
  42766=>"111000000",
  42767=>"100111010",
  42768=>"100010011",
  42769=>"011011011",
  42770=>"010010100",
  42771=>"100100000",
  42772=>"100100100",
  42773=>"001011001",
  42774=>"101100100",
  42775=>"001001010",
  42776=>"010011011",
  42777=>"001101100",
  42778=>"001011011",
  42779=>"001101100",
  42780=>"000110110",
  42781=>"110100100",
  42782=>"010011011",
  42783=>"100100100",
  42784=>"011010011",
  42785=>"010011111",
  42786=>"011001000",
  42787=>"010110110",
  42788=>"111000100",
  42789=>"100101000",
  42790=>"010011000",
  42791=>"111011000",
  42792=>"010100100",
  42793=>"010110000",
  42794=>"110010110",
  42795=>"100100100",
  42796=>"100100100",
  42797=>"000011111",
  42798=>"110111001",
  42799=>"111100110",
  42800=>"110110110",
  42801=>"110110110",
  42802=>"011011001",
  42803=>"001011011",
  42804=>"100100111",
  42805=>"110100100",
  42806=>"110100000",
  42807=>"100100111",
  42808=>"101011011",
  42809=>"100000100",
  42810=>"100100000",
  42811=>"010000111",
  42812=>"010000000",
  42813=>"100100100",
  42814=>"001011001",
  42815=>"010011011",
  42816=>"111011011",
  42817=>"100010111",
  42818=>"101001001",
  42819=>"000011011",
  42820=>"011001001",
  42821=>"001011001",
  42822=>"000010000",
  42823=>"000000000",
  42824=>"110100000",
  42825=>"000110110",
  42826=>"110011110",
  42827=>"001001111",
  42828=>"001001001",
  42829=>"000000001",
  42830=>"100001101",
  42831=>"011100111",
  42832=>"110000100",
  42833=>"100100111",
  42834=>"001011001",
  42835=>"100100111",
  42836=>"110100100",
  42837=>"100100100",
  42838=>"010000000",
  42839=>"001011001",
  42840=>"111011001",
  42841=>"111110100",
  42842=>"100100110",
  42843=>"011010010",
  42844=>"001001011",
  42845=>"110100100",
  42846=>"011011011",
  42847=>"010110100",
  42848=>"011011011",
  42849=>"001010101",
  42850=>"001011001",
  42851=>"110000000",
  42852=>"000000101",
  42853=>"110100010",
  42854=>"110100100",
  42855=>"100100111",
  42856=>"000101101",
  42857=>"001011011",
  42858=>"111011000",
  42859=>"101111111",
  42860=>"011011111",
  42861=>"111011001",
  42862=>"001001000",
  42863=>"110100000",
  42864=>"110101101",
  42865=>"010011011",
  42866=>"100100110",
  42867=>"000011000",
  42868=>"101111111",
  42869=>"000011011",
  42870=>"001111001",
  42871=>"001001001",
  42872=>"100010110",
  42873=>"110000100",
  42874=>"000001101",
  42875=>"011011001",
  42876=>"100101110",
  42877=>"100000000",
  42878=>"100100100",
  42879=>"111111100",
  42880=>"001011001",
  42881=>"110010110",
  42882=>"000011000",
  42883=>"111011101",
  42884=>"011001101",
  42885=>"000101101",
  42886=>"000100011",
  42887=>"011011000",
  42888=>"100100100",
  42889=>"110111101",
  42890=>"000100111",
  42891=>"101011110",
  42892=>"011100000",
  42893=>"101111110",
  42894=>"000011101",
  42895=>"011001001",
  42896=>"111101101",
  42897=>"010010110",
  42898=>"000010010",
  42899=>"100100100",
  42900=>"000000000",
  42901=>"011011001",
  42902=>"111101101",
  42903=>"000001000",
  42904=>"000100100",
  42905=>"101101111",
  42906=>"001001001",
  42907=>"001001011",
  42908=>"100111001",
  42909=>"000001111",
  42910=>"000011111",
  42911=>"110110100",
  42912=>"010110111",
  42913=>"101111111",
  42914=>"110101111",
  42915=>"001001001",
  42916=>"100001000",
  42917=>"001001001",
  42918=>"001111000",
  42919=>"110101001",
  42920=>"111001011",
  42921=>"001000110",
  42922=>"011011011",
  42923=>"100010001",
  42924=>"011100011",
  42925=>"000010110",
  42926=>"110100100",
  42927=>"011111101",
  42928=>"011011011",
  42929=>"000100010",
  42930=>"110000100",
  42931=>"000011110",
  42932=>"110000110",
  42933=>"100100000",
  42934=>"011011010",
  42935=>"000110110",
  42936=>"000100110",
  42937=>"101101100",
  42938=>"100110110",
  42939=>"000000100",
  42940=>"000110110",
  42941=>"000001001",
  42942=>"000010010",
  42943=>"000111110",
  42944=>"001111011",
  42945=>"100001001",
  42946=>"000011111",
  42947=>"100100110",
  42948=>"001011001",
  42949=>"110111110",
  42950=>"111011001",
  42951=>"000010000",
  42952=>"110101000",
  42953=>"011000110",
  42954=>"001111110",
  42955=>"001011000",
  42956=>"110100100",
  42957=>"110100000",
  42958=>"100000000",
  42959=>"011011011",
  42960=>"100100111",
  42961=>"100100100",
  42962=>"001101100",
  42963=>"001100111",
  42964=>"111011011",
  42965=>"100100100",
  42966=>"101111111",
  42967=>"111011111",
  42968=>"100100100",
  42969=>"011110010",
  42970=>"010000000",
  42971=>"011011011",
  42972=>"000000100",
  42973=>"001011001",
  42974=>"100000000",
  42975=>"111011011",
  42976=>"000010011",
  42977=>"001011001",
  42978=>"111101100",
  42979=>"011111101",
  42980=>"110110000",
  42981=>"100100110",
  42982=>"100110000",
  42983=>"000100100",
  42984=>"000011001",
  42985=>"110110110",
  42986=>"100100101",
  42987=>"011011000",
  42988=>"001011011",
  42989=>"011010100",
  42990=>"000000000",
  42991=>"111011110",
  42992=>"000110110",
  42993=>"100001011",
  42994=>"010011011",
  42995=>"100000000",
  42996=>"111110100",
  42997=>"011011011",
  42998=>"011011011",
  42999=>"111000110",
  43000=>"100001000",
  43001=>"100111110",
  43002=>"111111101",
  43003=>"111011111",
  43004=>"111110110",
  43005=>"110011011",
  43006=>"111110001",
  43007=>"000010100",
  43008=>"011001100",
  43009=>"111101000",
  43010=>"000010010",
  43011=>"000001011",
  43012=>"001011010",
  43013=>"100001111",
  43014=>"110111111",
  43015=>"100010010",
  43016=>"001101001",
  43017=>"110000111",
  43018=>"111111110",
  43019=>"001111111",
  43020=>"000110110",
  43021=>"000000000",
  43022=>"101011011",
  43023=>"000000001",
  43024=>"000010010",
  43025=>"001001000",
  43026=>"101001000",
  43027=>"110001111",
  43028=>"111000000",
  43029=>"000010011",
  43030=>"011101100",
  43031=>"111001111",
  43032=>"010000001",
  43033=>"011001101",
  43034=>"000000000",
  43035=>"000110110",
  43036=>"111101111",
  43037=>"000000000",
  43038=>"110100000",
  43039=>"001111101",
  43040=>"000111111",
  43041=>"111000101",
  43042=>"000000100",
  43043=>"000000111",
  43044=>"111111011",
  43045=>"110000100",
  43046=>"010111011",
  43047=>"000000000",
  43048=>"111111000",
  43049=>"011000000",
  43050=>"111011001",
  43051=>"111101001",
  43052=>"100000001",
  43053=>"110000000",
  43054=>"101100110",
  43055=>"101000000",
  43056=>"111010010",
  43057=>"111101101",
  43058=>"000000000",
  43059=>"111001000",
  43060=>"111111101",
  43061=>"111111111",
  43062=>"010110110",
  43063=>"000000000",
  43064=>"111010110",
  43065=>"000111011",
  43066=>"010000000",
  43067=>"111100000",
  43068=>"000001000",
  43069=>"111101111",
  43070=>"000010000",
  43071=>"000011001",
  43072=>"111001000",
  43073=>"000100110",
  43074=>"101101111",
  43075=>"001111110",
  43076=>"111101000",
  43077=>"000010010",
  43078=>"101011110",
  43079=>"101000000",
  43080=>"000000000",
  43081=>"111101100",
  43082=>"010010010",
  43083=>"000100100",
  43084=>"110000101",
  43085=>"011111111",
  43086=>"100111110",
  43087=>"000010111",
  43088=>"001111101",
  43089=>"111111111",
  43090=>"111111111",
  43091=>"011001110",
  43092=>"000111110",
  43093=>"001001000",
  43094=>"111011010",
  43095=>"100010010",
  43096=>"001111001",
  43097=>"011111111",
  43098=>"000111100",
  43099=>"101101000",
  43100=>"011101101",
  43101=>"000111001",
  43102=>"010111111",
  43103=>"100110011",
  43104=>"001101101",
  43105=>"010010000",
  43106=>"010111000",
  43107=>"000010001",
  43108=>"001101101",
  43109=>"111001001",
  43110=>"001000111",
  43111=>"111001111",
  43112=>"111000010",
  43113=>"111000000",
  43114=>"110011000",
  43115=>"000000101",
  43116=>"011011011",
  43117=>"100001011",
  43118=>"111111001",
  43119=>"010100101",
  43120=>"110100000",
  43121=>"111000000",
  43122=>"111011101",
  43123=>"000000111",
  43124=>"011111000",
  43125=>"000000111",
  43126=>"000000110",
  43127=>"111111111",
  43128=>"000011110",
  43129=>"001101111",
  43130=>"000000000",
  43131=>"101010010",
  43132=>"011101110",
  43133=>"110100000",
  43134=>"111101000",
  43135=>"000111100",
  43136=>"111101010",
  43137=>"111010010",
  43138=>"111111100",
  43139=>"000001100",
  43140=>"111110000",
  43141=>"101110111",
  43142=>"110000001",
  43143=>"011111000",
  43144=>"011101101",
  43145=>"010001011",
  43146=>"000000001",
  43147=>"000000000",
  43148=>"010111111",
  43149=>"000110111",
  43150=>"000111111",
  43151=>"001000001",
  43152=>"111101011",
  43153=>"101101001",
  43154=>"111101001",
  43155=>"001011010",
  43156=>"000001101",
  43157=>"111010110",
  43158=>"001111111",
  43159=>"000001001",
  43160=>"000110100",
  43161=>"001000000",
  43162=>"011111111",
  43163=>"001010000",
  43164=>"000001011",
  43165=>"000111100",
  43166=>"111000101",
  43167=>"111001111",
  43168=>"000000000",
  43169=>"010010000",
  43170=>"001111111",
  43171=>"011011000",
  43172=>"111111010",
  43173=>"110100100",
  43174=>"001110000",
  43175=>"101101101",
  43176=>"111011000",
  43177=>"000010001",
  43178=>"111111100",
  43179=>"111111101",
  43180=>"111000010",
  43181=>"010111000",
  43182=>"101101000",
  43183=>"001111111",
  43184=>"101000100",
  43185=>"100000000",
  43186=>"101101000",
  43187=>"001100100",
  43188=>"000011011",
  43189=>"001100111",
  43190=>"000110111",
  43191=>"000111010",
  43192=>"011001000",
  43193=>"000100000",
  43194=>"001101101",
  43195=>"110111111",
  43196=>"100000000",
  43197=>"111110000",
  43198=>"000100100",
  43199=>"000000000",
  43200=>"010000000",
  43201=>"000001111",
  43202=>"111000101",
  43203=>"111101001",
  43204=>"001111010",
  43205=>"101000000",
  43206=>"000100001",
  43207=>"111000000",
  43208=>"000000101",
  43209=>"000101111",
  43210=>"010100111",
  43211=>"010111110",
  43212=>"011001001",
  43213=>"110000011",
  43214=>"111101000",
  43215=>"000111111",
  43216=>"111111001",
  43217=>"011010000",
  43218=>"111111011",
  43219=>"000000100",
  43220=>"111111110",
  43221=>"101110000",
  43222=>"101111111",
  43223=>"110000000",
  43224=>"000111111",
  43225=>"110111001",
  43226=>"101001001",
  43227=>"111000000",
  43228=>"111011111",
  43229=>"000001101",
  43230=>"110011110",
  43231=>"111000000",
  43232=>"111110111",
  43233=>"001010010",
  43234=>"000111111",
  43235=>"001101011",
  43236=>"000000000",
  43237=>"100111110",
  43238=>"000000000",
  43239=>"011011101",
  43240=>"111100000",
  43241=>"111000101",
  43242=>"010110111",
  43243=>"000010010",
  43244=>"010111111",
  43245=>"000111111",
  43246=>"001011000",
  43247=>"010001000",
  43248=>"111111111",
  43249=>"011000000",
  43250=>"111110111",
  43251=>"000111110",
  43252=>"110100001",
  43253=>"001101101",
  43254=>"000001101",
  43255=>"101001001",
  43256=>"010111111",
  43257=>"111110000",
  43258=>"111111101",
  43259=>"001001010",
  43260=>"011111011",
  43261=>"111111111",
  43262=>"110101101",
  43263=>"000000000",
  43264=>"011100001",
  43265=>"010110111",
  43266=>"000000111",
  43267=>"100001111",
  43268=>"000001111",
  43269=>"000000000",
  43270=>"110111111",
  43271=>"111111111",
  43272=>"111000000",
  43273=>"111000111",
  43274=>"011011100",
  43275=>"010111111",
  43276=>"000000001",
  43277=>"000000000",
  43278=>"101001001",
  43279=>"000000111",
  43280=>"101100110",
  43281=>"000000000",
  43282=>"100100011",
  43283=>"111111000",
  43284=>"101101110",
  43285=>"111111100",
  43286=>"011011011",
  43287=>"111111000",
  43288=>"111111000",
  43289=>"101101111",
  43290=>"100101100",
  43291=>"111111111",
  43292=>"011111111",
  43293=>"111110000",
  43294=>"100000111",
  43295=>"110000000",
  43296=>"101111001",
  43297=>"000000111",
  43298=>"010010000",
  43299=>"000000000",
  43300=>"111110100",
  43301=>"000000010",
  43302=>"010011000",
  43303=>"000000001",
  43304=>"101000111",
  43305=>"111111110",
  43306=>"111001111",
  43307=>"011000000",
  43308=>"011110110",
  43309=>"111101111",
  43310=>"100000111",
  43311=>"001000000",
  43312=>"010000000",
  43313=>"001001000",
  43314=>"010010110",
  43315=>"111111010",
  43316=>"111111011",
  43317=>"111111010",
  43318=>"100000000",
  43319=>"100111100",
  43320=>"000011111",
  43321=>"110100111",
  43322=>"111111110",
  43323=>"011110011",
  43324=>"011001000",
  43325=>"011111011",
  43326=>"001000101",
  43327=>"111011011",
  43328=>"111000101",
  43329=>"000111000",
  43330=>"101001000",
  43331=>"100100111",
  43332=>"010111110",
  43333=>"001000000",
  43334=>"000000111",
  43335=>"111000110",
  43336=>"101111111",
  43337=>"000101111",
  43338=>"111111101",
  43339=>"100100111",
  43340=>"111110000",
  43341=>"001111000",
  43342=>"000100111",
  43343=>"010111110",
  43344=>"011000000",
  43345=>"010010011",
  43346=>"010111111",
  43347=>"111111001",
  43348=>"000000000",
  43349=>"111100110",
  43350=>"000000000",
  43351=>"100100111",
  43352=>"110111111",
  43353=>"111011001",
  43354=>"100001100",
  43355=>"000000000",
  43356=>"100101101",
  43357=>"001011111",
  43358=>"000000100",
  43359=>"000000001",
  43360=>"111111111",
  43361=>"000010000",
  43362=>"001001111",
  43363=>"001111011",
  43364=>"110011011",
  43365=>"011000000",
  43366=>"110111101",
  43367=>"111111000",
  43368=>"010111110",
  43369=>"000111111",
  43370=>"001111111",
  43371=>"000101101",
  43372=>"111111110",
  43373=>"101111100",
  43374=>"110100000",
  43375=>"000000110",
  43376=>"111001000",
  43377=>"001111111",
  43378=>"000000000",
  43379=>"000000000",
  43380=>"111011000",
  43381=>"001101111",
  43382=>"000000000",
  43383=>"000010000",
  43384=>"000000111",
  43385=>"111111111",
  43386=>"011001001",
  43387=>"000000000",
  43388=>"110000010",
  43389=>"111001100",
  43390=>"000000001",
  43391=>"000000111",
  43392=>"111111110",
  43393=>"111111111",
  43394=>"111111111",
  43395=>"010110111",
  43396=>"110110000",
  43397=>"111111111",
  43398=>"110011001",
  43399=>"011010011",
  43400=>"110100000",
  43401=>"011011000",
  43402=>"111010111",
  43403=>"001000100",
  43404=>"000000000",
  43405=>"011111111",
  43406=>"111100110",
  43407=>"000001000",
  43408=>"001001000",
  43409=>"111111101",
  43410=>"110111101",
  43411=>"000000000",
  43412=>"111100100",
  43413=>"000000101",
  43414=>"001101111",
  43415=>"000110000",
  43416=>"010010000",
  43417=>"111111111",
  43418=>"000010111",
  43419=>"000000111",
  43420=>"111111000",
  43421=>"000101011",
  43422=>"111101111",
  43423=>"010011111",
  43424=>"111111011",
  43425=>"111111111",
  43426=>"000000000",
  43427=>"111111111",
  43428=>"000111000",
  43429=>"110110110",
  43430=>"000000000",
  43431=>"111101011",
  43432=>"101000000",
  43433=>"010110111",
  43434=>"000000111",
  43435=>"010000001",
  43436=>"100110001",
  43437=>"000010101",
  43438=>"011001100",
  43439=>"111000111",
  43440=>"100100001",
  43441=>"100010100",
  43442=>"000000000",
  43443=>"000100100",
  43444=>"100010011",
  43445=>"010000000",
  43446=>"111111001",
  43447=>"101000111",
  43448=>"111010000",
  43449=>"101001000",
  43450=>"010000111",
  43451=>"111110010",
  43452=>"111111101",
  43453=>"100000100",
  43454=>"111001111",
  43455=>"000011000",
  43456=>"000000000",
  43457=>"110111001",
  43458=>"111111111",
  43459=>"100100100",
  43460=>"011011000",
  43461=>"111001111",
  43462=>"111111111",
  43463=>"000000000",
  43464=>"111111111",
  43465=>"111110010",
  43466=>"111111000",
  43467=>"000111111",
  43468=>"111111111",
  43469=>"100000110",
  43470=>"010111101",
  43471=>"001100111",
  43472=>"010011000",
  43473=>"111011000",
  43474=>"111111010",
  43475=>"001101101",
  43476=>"101111111",
  43477=>"000000001",
  43478=>"111101111",
  43479=>"000000010",
  43480=>"111011000",
  43481=>"010110010",
  43482=>"111111111",
  43483=>"010011000",
  43484=>"111000110",
  43485=>"000000110",
  43486=>"100010000",
  43487=>"000001101",
  43488=>"000000000",
  43489=>"101000111",
  43490=>"000000000",
  43491=>"001111111",
  43492=>"000011001",
  43493=>"000000000",
  43494=>"111111111",
  43495=>"101100100",
  43496=>"111111001",
  43497=>"000111001",
  43498=>"100010000",
  43499=>"000000000",
  43500=>"000011000",
  43501=>"100111000",
  43502=>"010010110",
  43503=>"010000101",
  43504=>"110111001",
  43505=>"111101111",
  43506=>"010000111",
  43507=>"111111000",
  43508=>"111111010",
  43509=>"111111000",
  43510=>"000000000",
  43511=>"110011000",
  43512=>"000000010",
  43513=>"110010000",
  43514=>"111111111",
  43515=>"000100101",
  43516=>"101100011",
  43517=>"100000000",
  43518=>"011111110",
  43519=>"010000000",
  43520=>"110100000",
  43521=>"000001000",
  43522=>"000000000",
  43523=>"000010010",
  43524=>"011011011",
  43525=>"111111001",
  43526=>"000010001",
  43527=>"111111100",
  43528=>"010111111",
  43529=>"010111111",
  43530=>"000011111",
  43531=>"000000010",
  43532=>"111111000",
  43533=>"110010111",
  43534=>"101111111",
  43535=>"111111111",
  43536=>"111111111",
  43537=>"111111111",
  43538=>"000101111",
  43539=>"111000101",
  43540=>"000101111",
  43541=>"111111111",
  43542=>"100110110",
  43543=>"011110000",
  43544=>"001001111",
  43545=>"000000000",
  43546=>"100111000",
  43547=>"011111111",
  43548=>"000001101",
  43549=>"011010000",
  43550=>"001000111",
  43551=>"111011010",
  43552=>"000000100",
  43553=>"111111111",
  43554=>"000000010",
  43555=>"111111111",
  43556=>"000000000",
  43557=>"000011001",
  43558=>"110111110",
  43559=>"000000001",
  43560=>"000000100",
  43561=>"000111101",
  43562=>"000000101",
  43563=>"111101111",
  43564=>"100110000",
  43565=>"000000000",
  43566=>"001000111",
  43567=>"000000001",
  43568=>"000111111",
  43569=>"011010100",
  43570=>"111111111",
  43571=>"000000111",
  43572=>"000000000",
  43573=>"000100000",
  43574=>"100111100",
  43575=>"000000111",
  43576=>"100111111",
  43577=>"000000000",
  43578=>"111000111",
  43579=>"001101111",
  43580=>"001001001",
  43581=>"111111010",
  43582=>"001101101",
  43583=>"101100111",
  43584=>"111111110",
  43585=>"001111111",
  43586=>"111111001",
  43587=>"111111111",
  43588=>"110111000",
  43589=>"001000010",
  43590=>"111111111",
  43591=>"000000000",
  43592=>"011000101",
  43593=>"000010111",
  43594=>"101110111",
  43595=>"001000000",
  43596=>"111111000",
  43597=>"010000000",
  43598=>"000000000",
  43599=>"111001000",
  43600=>"110111111",
  43601=>"111010000",
  43602=>"110100000",
  43603=>"000100100",
  43604=>"000000000",
  43605=>"011111111",
  43606=>"111011111",
  43607=>"011111011",
  43608=>"000110110",
  43609=>"000000100",
  43610=>"000011011",
  43611=>"000000000",
  43612=>"000111111",
  43613=>"010001001",
  43614=>"000000000",
  43615=>"111111100",
  43616=>"110110110",
  43617=>"000000001",
  43618=>"111110010",
  43619=>"001000100",
  43620=>"000000101",
  43621=>"000000001",
  43622=>"000000111",
  43623=>"000111111",
  43624=>"000001101",
  43625=>"111000011",
  43626=>"110000000",
  43627=>"111111101",
  43628=>"001101101",
  43629=>"000000110",
  43630=>"000001101",
  43631=>"000000111",
  43632=>"001001011",
  43633=>"000000111",
  43634=>"111011001",
  43635=>"111110111",
  43636=>"011000001",
  43637=>"000000100",
  43638=>"111111000",
  43639=>"111111111",
  43640=>"001010110",
  43641=>"111111000",
  43642=>"001001000",
  43643=>"110010111",
  43644=>"011001001",
  43645=>"001000000",
  43646=>"111111111",
  43647=>"110111111",
  43648=>"000111111",
  43649=>"111110010",
  43650=>"011100100",
  43651=>"101111111",
  43652=>"111000001",
  43653=>"000000000",
  43654=>"000110111",
  43655=>"100000000",
  43656=>"100010100",
  43657=>"101000111",
  43658=>"000000101",
  43659=>"111001011",
  43660=>"110111000",
  43661=>"111101110",
  43662=>"111101011",
  43663=>"001001011",
  43664=>"100100111",
  43665=>"111111111",
  43666=>"000111111",
  43667=>"111001000",
  43668=>"000001100",
  43669=>"111111111",
  43670=>"111111001",
  43671=>"000111111",
  43672=>"000000000",
  43673=>"010010110",
  43674=>"011110010",
  43675=>"111111000",
  43676=>"000000011",
  43677=>"010010011",
  43678=>"000111111",
  43679=>"000000000",
  43680=>"000110110",
  43681=>"000011110",
  43682=>"111111010",
  43683=>"100000000",
  43684=>"010111000",
  43685=>"000000010",
  43686=>"111111110",
  43687=>"000001010",
  43688=>"110010011",
  43689=>"011101011",
  43690=>"111111100",
  43691=>"000101111",
  43692=>"000000001",
  43693=>"110011011",
  43694=>"011011001",
  43695=>"001000110",
  43696=>"000000000",
  43697=>"000000001",
  43698=>"100110010",
  43699=>"101101011",
  43700=>"111000011",
  43701=>"000000000",
  43702=>"000000001",
  43703=>"001000000",
  43704=>"000100100",
  43705=>"000000000",
  43706=>"001000000",
  43707=>"011000000",
  43708=>"111000000",
  43709=>"111111011",
  43710=>"011011011",
  43711=>"000000000",
  43712=>"000000001",
  43713=>"001101111",
  43714=>"001001111",
  43715=>"000000110",
  43716=>"000000111",
  43717=>"000000001",
  43718=>"000000000",
  43719=>"110010000",
  43720=>"110000010",
  43721=>"010111001",
  43722=>"000000011",
  43723=>"001000000",
  43724=>"000000000",
  43725=>"100001100",
  43726=>"000101111",
  43727=>"110111110",
  43728=>"000000010",
  43729=>"100100111",
  43730=>"000000000",
  43731=>"111000000",
  43732=>"000001001",
  43733=>"000100100",
  43734=>"111111111",
  43735=>"000000001",
  43736=>"000000000",
  43737=>"000000010",
  43738=>"001001000",
  43739=>"110110010",
  43740=>"011111001",
  43741=>"111111010",
  43742=>"000000100",
  43743=>"000000000",
  43744=>"000111111",
  43745=>"110111000",
  43746=>"110111111",
  43747=>"101100111",
  43748=>"111001111",
  43749=>"111111001",
  43750=>"010010000",
  43751=>"000111111",
  43752=>"111110100",
  43753=>"001000111",
  43754=>"100010011",
  43755=>"111110000",
  43756=>"111111110",
  43757=>"000001010",
  43758=>"000000000",
  43759=>"110111110",
  43760=>"110000000",
  43761=>"000001000",
  43762=>"001001000",
  43763=>"101100001",
  43764=>"110000000",
  43765=>"111111111",
  43766=>"111111100",
  43767=>"100000000",
  43768=>"111111010",
  43769=>"011000000",
  43770=>"010011000",
  43771=>"010000000",
  43772=>"111111111",
  43773=>"000111001",
  43774=>"110000000",
  43775=>"001000000",
  43776=>"100100110",
  43777=>"011100001",
  43778=>"000010000",
  43779=>"101000000",
  43780=>"000111111",
  43781=>"001101111",
  43782=>"111000101",
  43783=>"010011000",
  43784=>"101001001",
  43785=>"001000000",
  43786=>"011000100",
  43787=>"111100000",
  43788=>"111001100",
  43789=>"000110000",
  43790=>"101100001",
  43791=>"001111101",
  43792=>"000000000",
  43793=>"010001000",
  43794=>"100000100",
  43795=>"111111101",
  43796=>"001001111",
  43797=>"011010001",
  43798=>"001111011",
  43799=>"110111110",
  43800=>"000000000",
  43801=>"000001111",
  43802=>"110110011",
  43803=>"101000101",
  43804=>"000101111",
  43805=>"010000000",
  43806=>"000101111",
  43807=>"000000000",
  43808=>"000111111",
  43809=>"000010111",
  43810=>"010010000",
  43811=>"000000101",
  43812=>"111110111",
  43813=>"001001011",
  43814=>"001111101",
  43815=>"001010111",
  43816=>"111111011",
  43817=>"011101111",
  43818=>"111100110",
  43819=>"011010000",
  43820=>"011100101",
  43821=>"111111111",
  43822=>"000110111",
  43823=>"000011010",
  43824=>"100001111",
  43825=>"000011001",
  43826=>"110000000",
  43827=>"010001011",
  43828=>"000000000",
  43829=>"001010111",
  43830=>"111111001",
  43831=>"100000000",
  43832=>"010100100",
  43833=>"101000000",
  43834=>"111101001",
  43835=>"110011111",
  43836=>"011001011",
  43837=>"111110111",
  43838=>"100000100",
  43839=>"000110000",
  43840=>"100101011",
  43841=>"000101111",
  43842=>"001100101",
  43843=>"000100100",
  43844=>"011101001",
  43845=>"000111111",
  43846=>"000111111",
  43847=>"101000001",
  43848=>"011111111",
  43849=>"111100101",
  43850=>"101101111",
  43851=>"101000000",
  43852=>"100000101",
  43853=>"111101010",
  43854=>"001110110",
  43855=>"010010111",
  43856=>"111101101",
  43857=>"111111111",
  43858=>"010000000",
  43859=>"010001000",
  43860=>"111000000",
  43861=>"010110010",
  43862=>"001011010",
  43863=>"100000001",
  43864=>"010000000",
  43865=>"011001001",
  43866=>"001010000",
  43867=>"010111101",
  43868=>"111000000",
  43869=>"100110000",
  43870=>"010011010",
  43871=>"000000001",
  43872=>"000000000",
  43873=>"100100100",
  43874=>"000000001",
  43875=>"000110110",
  43876=>"111001001",
  43877=>"000111111",
  43878=>"111101010",
  43879=>"000000101",
  43880=>"011011001",
  43881=>"110111101",
  43882=>"011111101",
  43883=>"111101001",
  43884=>"001000001",
  43885=>"001000000",
  43886=>"001101101",
  43887=>"000101011",
  43888=>"100110110",
  43889=>"000000010",
  43890=>"011001100",
  43891=>"000000000",
  43892=>"000001111",
  43893=>"000001101",
  43894=>"000000001",
  43895=>"011101100",
  43896=>"110111010",
  43897=>"000100111",
  43898=>"010010111",
  43899=>"011000001",
  43900=>"001001001",
  43901=>"000001000",
  43902=>"011011000",
  43903=>"101001001",
  43904=>"111000000",
  43905=>"011011010",
  43906=>"101111001",
  43907=>"101111111",
  43908=>"000101111",
  43909=>"011000000",
  43910=>"000101100",
  43911=>"100000101",
  43912=>"000011001",
  43913=>"110100100",
  43914=>"001000100",
  43915=>"111101111",
  43916=>"000111010",
  43917=>"111001011",
  43918=>"100101100",
  43919=>"001000101",
  43920=>"000100101",
  43921=>"000110110",
  43922=>"101111011",
  43923=>"100100010",
  43924=>"000010000",
  43925=>"000000110",
  43926=>"111100100",
  43927=>"011001000",
  43928=>"111101011",
  43929=>"101111111",
  43930=>"001100000",
  43931=>"000000000",
  43932=>"100100100",
  43933=>"111000000",
  43934=>"000101111",
  43935=>"111100111",
  43936=>"111011111",
  43937=>"111111011",
  43938=>"111101111",
  43939=>"100000101",
  43940=>"110011111",
  43941=>"000000001",
  43942=>"111101010",
  43943=>"111101000",
  43944=>"010010111",
  43945=>"000000000",
  43946=>"100111111",
  43947=>"100000000",
  43948=>"010011010",
  43949=>"000000101",
  43950=>"111111001",
  43951=>"011101101",
  43952=>"000001000",
  43953=>"111110100",
  43954=>"000100100",
  43955=>"000000100",
  43956=>"111111011",
  43957=>"101000100",
  43958=>"000000110",
  43959=>"000001110",
  43960=>"011100110",
  43961=>"011000010",
  43962=>"101001101",
  43963=>"100000101",
  43964=>"111111110",
  43965=>"111011000",
  43966=>"000101000",
  43967=>"000110111",
  43968=>"010111001",
  43969=>"111000000",
  43970=>"111101101",
  43971=>"110100110",
  43972=>"000000000",
  43973=>"110111110",
  43974=>"100000000",
  43975=>"000000000",
  43976=>"010000000",
  43977=>"000011011",
  43978=>"000000010",
  43979=>"000000001",
  43980=>"100000000",
  43981=>"110100101",
  43982=>"000000001",
  43983=>"000001010",
  43984=>"110111010",
  43985=>"010011101",
  43986=>"000000101",
  43987=>"000011111",
  43988=>"000010000",
  43989=>"000001011",
  43990=>"001000000",
  43991=>"111101011",
  43992=>"011011000",
  43993=>"010010100",
  43994=>"111111101",
  43995=>"101000000",
  43996=>"010011011",
  43997=>"110100000",
  43998=>"010000000",
  43999=>"000111101",
  44000=>"010000000",
  44001=>"100000101",
  44002=>"001111111",
  44003=>"001100000",
  44004=>"000010011",
  44005=>"000000000",
  44006=>"110000000",
  44007=>"011111111",
  44008=>"101000100",
  44009=>"000011111",
  44010=>"100100001",
  44011=>"000000000",
  44012=>"101000000",
  44013=>"000010111",
  44014=>"000000100",
  44015=>"000000100",
  44016=>"011010000",
  44017=>"111111011",
  44018=>"100000000",
  44019=>"110110000",
  44020=>"101001111",
  44021=>"011000000",
  44022=>"000000001",
  44023=>"000011000",
  44024=>"000111111",
  44025=>"000111111",
  44026=>"000010010",
  44027=>"111111101",
  44028=>"100100101",
  44029=>"100000000",
  44030=>"111110111",
  44031=>"010000111",
  44032=>"001100100",
  44033=>"000000000",
  44034=>"101000000",
  44035=>"011111011",
  44036=>"000011101",
  44037=>"000000001",
  44038=>"000111010",
  44039=>"000011011",
  44040=>"010001001",
  44041=>"010010000",
  44042=>"001001001",
  44043=>"110110111",
  44044=>"000000000",
  44045=>"001000000",
  44046=>"001011011",
  44047=>"001111110",
  44048=>"010000000",
  44049=>"000000000",
  44050=>"000000101",
  44051=>"000000000",
  44052=>"111111111",
  44053=>"111011000",
  44054=>"011011111",
  44055=>"111010000",
  44056=>"100100001",
  44057=>"111010101",
  44058=>"011001001",
  44059=>"011010001",
  44060=>"111000001",
  44061=>"001101001",
  44062=>"110000000",
  44063=>"000001111",
  44064=>"000000000",
  44065=>"100011001",
  44066=>"000111001",
  44067=>"111111000",
  44068=>"100101101",
  44069=>"110000001",
  44070=>"001001001",
  44071=>"010000011",
  44072=>"000000111",
  44073=>"010010000",
  44074=>"110010000",
  44075=>"010000111",
  44076=>"000000000",
  44077=>"111000100",
  44078=>"011010000",
  44079=>"111111011",
  44080=>"110000001",
  44081=>"100111101",
  44082=>"110000000",
  44083=>"010000000",
  44084=>"000000111",
  44085=>"110011011",
  44086=>"001011001",
  44087=>"000011000",
  44088=>"010000000",
  44089=>"100000000",
  44090=>"001110110",
  44091=>"000000101",
  44092=>"100110110",
  44093=>"111101110",
  44094=>"000010000",
  44095=>"000110000",
  44096=>"111011101",
  44097=>"110110000",
  44098=>"011111100",
  44099=>"000100100",
  44100=>"111100000",
  44101=>"010010101",
  44102=>"000000110",
  44103=>"001010111",
  44104=>"101011100",
  44105=>"111111001",
  44106=>"000000100",
  44107=>"000110111",
  44108=>"010000010",
  44109=>"001111101",
  44110=>"000101001",
  44111=>"111100111",
  44112=>"000001111",
  44113=>"101000000",
  44114=>"111010111",
  44115=>"011000110",
  44116=>"101110101",
  44117=>"000000000",
  44118=>"001100000",
  44119=>"000111101",
  44120=>"100100110",
  44121=>"001111110",
  44122=>"100101011",
  44123=>"011011001",
  44124=>"010010000",
  44125=>"000001001",
  44126=>"111010001",
  44127=>"000001111",
  44128=>"000111010",
  44129=>"000001000",
  44130=>"101101001",
  44131=>"111111101",
  44132=>"000110110",
  44133=>"000001100",
  44134=>"100110111",
  44135=>"001111101",
  44136=>"000000111",
  44137=>"111010000",
  44138=>"011011010",
  44139=>"011010000",
  44140=>"111000001",
  44141=>"111001111",
  44142=>"101000000",
  44143=>"111000101",
  44144=>"001111111",
  44145=>"110110000",
  44146=>"100100100",
  44147=>"101111101",
  44148=>"110111101",
  44149=>"000000000",
  44150=>"000000000",
  44151=>"000100000",
  44152=>"010010111",
  44153=>"000010011",
  44154=>"100000010",
  44155=>"111011000",
  44156=>"100110110",
  44157=>"100000000",
  44158=>"000001111",
  44159=>"111111100",
  44160=>"000000110",
  44161=>"111000110",
  44162=>"111111001",
  44163=>"101101010",
  44164=>"111000001",
  44165=>"010000110",
  44166=>"011011000",
  44167=>"000110100",
  44168=>"100111111",
  44169=>"101011010",
  44170=>"011110100",
  44171=>"000000000",
  44172=>"111111111",
  44173=>"000011010",
  44174=>"010011010",
  44175=>"000001010",
  44176=>"101100111",
  44177=>"010000100",
  44178=>"010111111",
  44179=>"101101111",
  44180=>"011100000",
  44181=>"111011000",
  44182=>"111010000",
  44183=>"000001011",
  44184=>"111011000",
  44185=>"111011011",
  44186=>"111101000",
  44187=>"000000011",
  44188=>"110001010",
  44189=>"010011000",
  44190=>"010011100",
  44191=>"000111000",
  44192=>"000001100",
  44193=>"000101111",
  44194=>"001001000",
  44195=>"001101010",
  44196=>"111001111",
  44197=>"100110000",
  44198=>"010110101",
  44199=>"000001010",
  44200=>"111010100",
  44201=>"000111111",
  44202=>"101000101",
  44203=>"000101111",
  44204=>"010001100",
  44205=>"000111111",
  44206=>"000001011",
  44207=>"010010010",
  44208=>"110110111",
  44209=>"000001001",
  44210=>"010000100",
  44211=>"100110110",
  44212=>"110111001",
  44213=>"001011000",
  44214=>"011111010",
  44215=>"111010000",
  44216=>"001011011",
  44217=>"000001000",
  44218=>"010011010",
  44219=>"010010000",
  44220=>"101101010",
  44221=>"101011010",
  44222=>"101111000",
  44223=>"010000110",
  44224=>"010110010",
  44225=>"010010000",
  44226=>"010010111",
  44227=>"100101111",
  44228=>"110100100",
  44229=>"100110111",
  44230=>"000000000",
  44231=>"111010001",
  44232=>"111011011",
  44233=>"000000100",
  44234=>"101111100",
  44235=>"111011001",
  44236=>"000001000",
  44237=>"001011000",
  44238=>"000100000",
  44239=>"010001111",
  44240=>"101010010",
  44241=>"000101111",
  44242=>"110100111",
  44243=>"000101111",
  44244=>"110110111",
  44245=>"001101110",
  44246=>"110010101",
  44247=>"110010001",
  44248=>"100000010",
  44249=>"111010001",
  44250=>"000100000",
  44251=>"111000000",
  44252=>"110111101",
  44253=>"111101001",
  44254=>"000011011",
  44255=>"010010001",
  44256=>"101111111",
  44257=>"011111101",
  44258=>"111000111",
  44259=>"100111111",
  44260=>"000111000",
  44261=>"000101111",
  44262=>"100111110",
  44263=>"000100100",
  44264=>"011010101",
  44265=>"000000000",
  44266=>"100100100",
  44267=>"111111001",
  44268=>"000000000",
  44269=>"000000000",
  44270=>"000000110",
  44271=>"010001000",
  44272=>"101001001",
  44273=>"001011101",
  44274=>"111011010",
  44275=>"000011110",
  44276=>"000001001",
  44277=>"111101001",
  44278=>"010110000",
  44279=>"010000111",
  44280=>"110000000",
  44281=>"001010010",
  44282=>"011110110",
  44283=>"101111111",
  44284=>"111111010",
  44285=>"111111111",
  44286=>"000111111",
  44287=>"000011010",
  44288=>"000000100",
  44289=>"000001011",
  44290=>"100100100",
  44291=>"010100111",
  44292=>"110000001",
  44293=>"110100000",
  44294=>"111011011",
  44295=>"000011011",
  44296=>"100100100",
  44297=>"110001001",
  44298=>"000011011",
  44299=>"000000011",
  44300=>"110100000",
  44301=>"000100001",
  44302=>"110101000",
  44303=>"111110101",
  44304=>"001011000",
  44305=>"110001011",
  44306=>"110100010",
  44307=>"001001011",
  44308=>"110110111",
  44309=>"110110111",
  44310=>"000010001",
  44311=>"101011011",
  44312=>"110000000",
  44313=>"110010110",
  44314=>"110000011",
  44315=>"001001000",
  44316=>"000000110",
  44317=>"110000100",
  44318=>"100100000",
  44319=>"110100100",
  44320=>"101101100",
  44321=>"110010001",
  44322=>"111100000",
  44323=>"000000000",
  44324=>"011111100",
  44325=>"001101101",
  44326=>"100001111",
  44327=>"001011010",
  44328=>"111010100",
  44329=>"000000000",
  44330=>"110010011",
  44331=>"001000000",
  44332=>"011110011",
  44333=>"110100100",
  44334=>"011110111",
  44335=>"111010111",
  44336=>"001111100",
  44337=>"101110000",
  44338=>"100000101",
  44339=>"001110011",
  44340=>"000011111",
  44341=>"011011110",
  44342=>"010100101",
  44343=>"000011011",
  44344=>"001100111",
  44345=>"110100000",
  44346=>"111100100",
  44347=>"001011010",
  44348=>"011110000",
  44349=>"011111111",
  44350=>"100001000",
  44351=>"001000111",
  44352=>"111000010",
  44353=>"001011010",
  44354=>"111011000",
  44355=>"100001001",
  44356=>"111100010",
  44357=>"100000001",
  44358=>"100110101",
  44359=>"111101100",
  44360=>"111111101",
  44361=>"000100011",
  44362=>"011001011",
  44363=>"000001011",
  44364=>"111100111",
  44365=>"100101100",
  44366=>"000011110",
  44367=>"011110000",
  44368=>"000000001",
  44369=>"011111111",
  44370=>"010111100",
  44371=>"001001010",
  44372=>"111100100",
  44373=>"000111110",
  44374=>"111110111",
  44375=>"110100000",
  44376=>"111011111",
  44377=>"000000000",
  44378=>"001001101",
  44379=>"000001000",
  44380=>"000001000",
  44381=>"110100000",
  44382=>"101011001",
  44383=>"010100001",
  44384=>"110110110",
  44385=>"010100001",
  44386=>"110100111",
  44387=>"111111100",
  44388=>"000110100",
  44389=>"001000000",
  44390=>"000100111",
  44391=>"000000110",
  44392=>"100100100",
  44393=>"111100110",
  44394=>"111011000",
  44395=>"111011111",
  44396=>"001000010",
  44397=>"100001011",
  44398=>"011000000",
  44399=>"110111011",
  44400=>"010111000",
  44401=>"001000011",
  44402=>"000001011",
  44403=>"100100100",
  44404=>"011011010",
  44405=>"110100011",
  44406=>"100100010",
  44407=>"000100100",
  44408=>"111101001",
  44409=>"000011111",
  44410=>"101011010",
  44411=>"111110100",
  44412=>"001011011",
  44413=>"011110000",
  44414=>"001011111",
  44415=>"110100100",
  44416=>"011010100",
  44417=>"100100000",
  44418=>"100011011",
  44419=>"000111000",
  44420=>"100100001",
  44421=>"010100100",
  44422=>"001001110",
  44423=>"000001001",
  44424=>"011111101",
  44425=>"000000000",
  44426=>"110011000",
  44427=>"101011010",
  44428=>"110001001",
  44429=>"000100111",
  44430=>"010111100",
  44431=>"110000001",
  44432=>"011010100",
  44433=>"000001011",
  44434=>"001011010",
  44435=>"000011010",
  44436=>"110001000",
  44437=>"100000011",
  44438=>"100111111",
  44439=>"111110000",
  44440=>"001011000",
  44441=>"110100000",
  44442=>"110110100",
  44443=>"100100101",
  44444=>"011001011",
  44445=>"110100100",
  44446=>"011001001",
  44447=>"000000010",
  44448=>"000000110",
  44449=>"101100001",
  44450=>"000101001",
  44451=>"000101010",
  44452=>"110010011",
  44453=>"101101001",
  44454=>"001010011",
  44455=>"000000000",
  44456=>"011001011",
  44457=>"010110110",
  44458=>"000100100",
  44459=>"111000001",
  44460=>"100100000",
  44461=>"110100100",
  44462=>"111111011",
  44463=>"001011010",
  44464=>"111000000",
  44465=>"000001111",
  44466=>"111110110",
  44467=>"001010110",
  44468=>"000110111",
  44469=>"011111000",
  44470=>"000001001",
  44471=>"011001011",
  44472=>"000001000",
  44473=>"000001100",
  44474=>"011100100",
  44475=>"011110100",
  44476=>"111111110",
  44477=>"111011001",
  44478=>"000000000",
  44479=>"001010000",
  44480=>"110100000",
  44481=>"000001001",
  44482=>"100110010",
  44483=>"000000000",
  44484=>"001010000",
  44485=>"111110110",
  44486=>"000111011",
  44487=>"110100100",
  44488=>"010110110",
  44489=>"010000011",
  44490=>"011101110",
  44491=>"100111000",
  44492=>"000001000",
  44493=>"000001000",
  44494=>"011001001",
  44495=>"110101000",
  44496=>"101000000",
  44497=>"000000000",
  44498=>"100110010",
  44499=>"011110000",
  44500=>"100100011",
  44501=>"001010000",
  44502=>"011100000",
  44503=>"011111001",
  44504=>"001011111",
  44505=>"111000000",
  44506=>"011110100",
  44507=>"111100011",
  44508=>"111011010",
  44509=>"100100100",
  44510=>"010100111",
  44511=>"110000001",
  44512=>"111010100",
  44513=>"101100000",
  44514=>"000011111",
  44515=>"000111101",
  44516=>"000010001",
  44517=>"100001111",
  44518=>"111101010",
  44519=>"001001100",
  44520=>"111111111",
  44521=>"001011001",
  44522=>"000001001",
  44523=>"000100100",
  44524=>"000010010",
  44525=>"010010011",
  44526=>"000000000",
  44527=>"111000100",
  44528=>"001000011",
  44529=>"000000010",
  44530=>"000011001",
  44531=>"111111100",
  44532=>"000011000",
  44533=>"111010001",
  44534=>"100000000",
  44535=>"001000100",
  44536=>"000011010",
  44537=>"111111110",
  44538=>"011100111",
  44539=>"100110100",
  44540=>"010111110",
  44541=>"001011110",
  44542=>"000000000",
  44543=>"000011010",
  44544=>"011000001",
  44545=>"000110111",
  44546=>"101101101",
  44547=>"000000110",
  44548=>"111000100",
  44549=>"010000000",
  44550=>"000010111",
  44551=>"000000000",
  44552=>"101111111",
  44553=>"111101000",
  44554=>"010100111",
  44555=>"000100101",
  44556=>"000011111",
  44557=>"000100111",
  44558=>"100101111",
  44559=>"110111110",
  44560=>"000000010",
  44561=>"000000010",
  44562=>"000000101",
  44563=>"010010000",
  44564=>"111101111",
  44565=>"101010111",
  44566=>"001111011",
  44567=>"000000000",
  44568=>"111000101",
  44569=>"111100010",
  44570=>"011101100",
  44571=>"000000100",
  44572=>"000001111",
  44573=>"111010011",
  44574=>"111101001",
  44575=>"000010110",
  44576=>"111101100",
  44577=>"001101111",
  44578=>"000010010",
  44579=>"010111000",
  44580=>"000110100",
  44581=>"100000000",
  44582=>"100101011",
  44583=>"001000101",
  44584=>"110010000",
  44585=>"001110110",
  44586=>"010000000",
  44587=>"100001001",
  44588=>"110010011",
  44589=>"010111101",
  44590=>"011111101",
  44591=>"111011101",
  44592=>"010001000",
  44593=>"000110111",
  44594=>"000011000",
  44595=>"000111110",
  44596=>"000000010",
  44597=>"011011110",
  44598=>"000100000",
  44599=>"000110011",
  44600=>"000000000",
  44601=>"000100101",
  44602=>"000111101",
  44603=>"001000111",
  44604=>"110000111",
  44605=>"111101101",
  44606=>"001000000",
  44607=>"000000110",
  44608=>"000000010",
  44609=>"000000010",
  44610=>"101101001",
  44611=>"000000110",
  44612=>"111101101",
  44613=>"000010000",
  44614=>"000000111",
  44615=>"010000111",
  44616=>"001101000",
  44617=>"001001111",
  44618=>"000000000",
  44619=>"111111101",
  44620=>"100101101",
  44621=>"001101001",
  44622=>"110000111",
  44623=>"010000010",
  44624=>"000101000",
  44625=>"110000100",
  44626=>"000000011",
  44627=>"001001001",
  44628=>"001010010",
  44629=>"011010111",
  44630=>"000011011",
  44631=>"000000000",
  44632=>"000111101",
  44633=>"001011111",
  44634=>"110100100",
  44635=>"001011010",
  44636=>"000101001",
  44637=>"000001111",
  44638=>"110111010",
  44639=>"000000001",
  44640=>"000101111",
  44641=>"000000110",
  44642=>"000001001",
  44643=>"001000001",
  44644=>"010000101",
  44645=>"000100000",
  44646=>"010111110",
  44647=>"101111010",
  44648=>"000001110",
  44649=>"100000101",
  44650=>"111111010",
  44651=>"111100101",
  44652=>"010101111",
  44653=>"111010110",
  44654=>"000000111",
  44655=>"011011111",
  44656=>"110111101",
  44657=>"000000110",
  44658=>"001101000",
  44659=>"011011000",
  44660=>"111110010",
  44661=>"101001001",
  44662=>"000010010",
  44663=>"111111111",
  44664=>"010000000",
  44665=>"111100011",
  44666=>"010110010",
  44667=>"111111101",
  44668=>"001001001",
  44669=>"110100100",
  44670=>"000000011",
  44671=>"101111101",
  44672=>"010000000",
  44673=>"000010111",
  44674=>"111000111",
  44675=>"010000011",
  44676=>"110000000",
  44677=>"001000000",
  44678=>"000000010",
  44679=>"000000000",
  44680=>"100110110",
  44681=>"000101000",
  44682=>"011001000",
  44683=>"010000000",
  44684=>"111110000",
  44685=>"100000111",
  44686=>"111100101",
  44687=>"001000000",
  44688=>"011000000",
  44689=>"000000000",
  44690=>"111001000",
  44691=>"000000010",
  44692=>"000000000",
  44693=>"111000000",
  44694=>"010111111",
  44695=>"000011001",
  44696=>"110010111",
  44697=>"000001101",
  44698=>"000010011",
  44699=>"101000100",
  44700=>"100101111",
  44701=>"011001000",
  44702=>"001100000",
  44703=>"110100110",
  44704=>"111111011",
  44705=>"000011000",
  44706=>"000000111",
  44707=>"000000001",
  44708=>"111100100",
  44709=>"100110110",
  44710=>"010110000",
  44711=>"000000100",
  44712=>"010000110",
  44713=>"000111110",
  44714=>"111111101",
  44715=>"101000000",
  44716=>"010010111",
  44717=>"000000000",
  44718=>"100100100",
  44719=>"000000111",
  44720=>"110100011",
  44721=>"101001111",
  44722=>"111101101",
  44723=>"000000000",
  44724=>"110011001",
  44725=>"010011001",
  44726=>"111101000",
  44727=>"001000001",
  44728=>"010000011",
  44729=>"000100000",
  44730=>"000000001",
  44731=>"110110100",
  44732=>"111000111",
  44733=>"011111101",
  44734=>"011011111",
  44735=>"000111000",
  44736=>"000001101",
  44737=>"000000101",
  44738=>"000101110",
  44739=>"001110111",
  44740=>"000000001",
  44741=>"010110100",
  44742=>"010010001",
  44743=>"000000000",
  44744=>"101111111",
  44745=>"110111000",
  44746=>"111101111",
  44747=>"101010010",
  44748=>"111100100",
  44749=>"000100000",
  44750=>"111111010",
  44751=>"000010000",
  44752=>"101000000",
  44753=>"110110110",
  44754=>"000010110",
  44755=>"111010111",
  44756=>"101000000",
  44757=>"101111111",
  44758=>"000101111",
  44759=>"100101110",
  44760=>"000010011",
  44761=>"010010000",
  44762=>"111011110",
  44763=>"100000000",
  44764=>"100011110",
  44765=>"111011111",
  44766=>"000001000",
  44767=>"000010000",
  44768=>"000000001",
  44769=>"101101100",
  44770=>"000000000",
  44771=>"001011111",
  44772=>"111001000",
  44773=>"010101011",
  44774=>"000000011",
  44775=>"001001011",
  44776=>"010000010",
  44777=>"000000001",
  44778=>"110011011",
  44779=>"010010010",
  44780=>"000010010",
  44781=>"111011000",
  44782=>"000000000",
  44783=>"000000010",
  44784=>"010010110",
  44785=>"100010001",
  44786=>"000001000",
  44787=>"110010100",
  44788=>"000110001",
  44789=>"101101101",
  44790=>"000000000",
  44791=>"000111110",
  44792=>"000000000",
  44793=>"000100000",
  44794=>"101101001",
  44795=>"010011000",
  44796=>"111111010",
  44797=>"010000100",
  44798=>"100000001",
  44799=>"010000010",
  44800=>"000010110",
  44801=>"000000000",
  44802=>"101101101",
  44803=>"111011011",
  44804=>"100000011",
  44805=>"100000101",
  44806=>"000110111",
  44807=>"111010010",
  44808=>"000010010",
  44809=>"000111011",
  44810=>"100000100",
  44811=>"101000000",
  44812=>"010100000",
  44813=>"000000001",
  44814=>"111110110",
  44815=>"000011110",
  44816=>"110110110",
  44817=>"000000110",
  44818=>"111000110",
  44819=>"000010010",
  44820=>"101111110",
  44821=>"101001111",
  44822=>"101001000",
  44823=>"101110111",
  44824=>"001000000",
  44825=>"110010000",
  44826=>"000010010",
  44827=>"000110010",
  44828=>"000101000",
  44829=>"111000010",
  44830=>"111101101",
  44831=>"111001000",
  44832=>"111000000",
  44833=>"000010110",
  44834=>"000001001",
  44835=>"000000000",
  44836=>"000111010",
  44837=>"011111111",
  44838=>"010110111",
  44839=>"110111111",
  44840=>"000010000",
  44841=>"101010110",
  44842=>"000110010",
  44843=>"100001000",
  44844=>"000011111",
  44845=>"111111111",
  44846=>"111010111",
  44847=>"001001111",
  44848=>"000101000",
  44849=>"110000101",
  44850=>"101110111",
  44851=>"110111111",
  44852=>"111000000",
  44853=>"000000010",
  44854=>"111000100",
  44855=>"110100000",
  44856=>"000010111",
  44857=>"001100001",
  44858=>"100011111",
  44859=>"000000000",
  44860=>"111111100",
  44861=>"111011001",
  44862=>"001101000",
  44863=>"000010101",
  44864=>"111000111",
  44865=>"101111111",
  44866=>"110000100",
  44867=>"000000100",
  44868=>"111000011",
  44869=>"000101111",
  44870=>"111100000",
  44871=>"111010000",
  44872=>"011110111",
  44873=>"010010010",
  44874=>"000100101",
  44875=>"100011111",
  44876=>"110000000",
  44877=>"000111111",
  44878=>"001100100",
  44879=>"100110010",
  44880=>"111001000",
  44881=>"111011101",
  44882=>"011010010",
  44883=>"110011001",
  44884=>"101000000",
  44885=>"011111111",
  44886=>"000111000",
  44887=>"001001101",
  44888=>"001111000",
  44889=>"011010000",
  44890=>"011000000",
  44891=>"000110100",
  44892=>"100111111",
  44893=>"001011111",
  44894=>"101011110",
  44895=>"000000001",
  44896=>"000000000",
  44897=>"111011001",
  44898=>"101001101",
  44899=>"110100000",
  44900=>"000111101",
  44901=>"000111000",
  44902=>"000110110",
  44903=>"100000000",
  44904=>"110011111",
  44905=>"000010111",
  44906=>"000001111",
  44907=>"110110001",
  44908=>"001110111",
  44909=>"000110111",
  44910=>"011000100",
  44911=>"000111111",
  44912=>"001111001",
  44913=>"100110110",
  44914=>"111101000",
  44915=>"101011000",
  44916=>"010010101",
  44917=>"010001001",
  44918=>"000000000",
  44919=>"111011000",
  44920=>"111000101",
  44921=>"010010000",
  44922=>"000000000",
  44923=>"100111111",
  44924=>"111110010",
  44925=>"110110100",
  44926=>"100111111",
  44927=>"111000000",
  44928=>"010110001",
  44929=>"111100000",
  44930=>"000110100",
  44931=>"010111111",
  44932=>"011110100",
  44933=>"010010000",
  44934=>"100110111",
  44935=>"011000000",
  44936=>"001110100",
  44937=>"000100011",
  44938=>"100111111",
  44939=>"010001110",
  44940=>"000001001",
  44941=>"110111111",
  44942=>"111010000",
  44943=>"110001001",
  44944=>"100011001",
  44945=>"010111111",
  44946=>"100111110",
  44947=>"000000100",
  44948=>"111000000",
  44949=>"101101111",
  44950=>"010011000",
  44951=>"000010000",
  44952=>"000100001",
  44953=>"100000000",
  44954=>"001111101",
  44955=>"111100001",
  44956=>"111111100",
  44957=>"111001001",
  44958=>"001010000",
  44959=>"111101101",
  44960=>"110111011",
  44961=>"000111101",
  44962=>"100010111",
  44963=>"000111101",
  44964=>"000111111",
  44965=>"010110000",
  44966=>"100001111",
  44967=>"000010000",
  44968=>"000000110",
  44969=>"010010010",
  44970=>"001101101",
  44971=>"101000000",
  44972=>"110101101",
  44973=>"100000000",
  44974=>"111110001",
  44975=>"010001111",
  44976=>"111000110",
  44977=>"110001001",
  44978=>"110111000",
  44979=>"110101000",
  44980=>"000011100",
  44981=>"010111111",
  44982=>"101111010",
  44983=>"100110111",
  44984=>"111111101",
  44985=>"011000000",
  44986=>"111010000",
  44987=>"000000111",
  44988=>"111111110",
  44989=>"111101111",
  44990=>"011011001",
  44991=>"000110000",
  44992=>"011001101",
  44993=>"000000000",
  44994=>"010110011",
  44995=>"000110110",
  44996=>"000010011",
  44997=>"011000110",
  44998=>"000000000",
  44999=>"011111000",
  45000=>"101111111",
  45001=>"001001000",
  45002=>"111111010",
  45003=>"101000010",
  45004=>"111010000",
  45005=>"111110010",
  45006=>"101000000",
  45007=>"000000001",
  45008=>"011101111",
  45009=>"011111100",
  45010=>"000000000",
  45011=>"101000000",
  45012=>"001001000",
  45013=>"110000000",
  45014=>"110010010",
  45015=>"000000000",
  45016=>"001000110",
  45017=>"001111110",
  45018=>"010110101",
  45019=>"000000101",
  45020=>"110010000",
  45021=>"111101101",
  45022=>"110000000",
  45023=>"100000000",
  45024=>"111000100",
  45025=>"111100000",
  45026=>"101101011",
  45027=>"011111001",
  45028=>"111000000",
  45029=>"011000000",
  45030=>"101110111",
  45031=>"000110001",
  45032=>"010111100",
  45033=>"000000000",
  45034=>"001001011",
  45035=>"100001111",
  45036=>"111100110",
  45037=>"000000000",
  45038=>"111100000",
  45039=>"111100000",
  45040=>"111000000",
  45041=>"110000011",
  45042=>"000000000",
  45043=>"110110111",
  45044=>"000111111",
  45045=>"000000000",
  45046=>"010000000",
  45047=>"000010000",
  45048=>"000100110",
  45049=>"111110101",
  45050=>"010110010",
  45051=>"000000010",
  45052=>"000110111",
  45053=>"100000000",
  45054=>"001111100",
  45055=>"101111101",
  45056=>"101000001",
  45057=>"010111111",
  45058=>"111111010",
  45059=>"000000101",
  45060=>"111000100",
  45061=>"101001000",
  45062=>"111100111",
  45063=>"100101100",
  45064=>"100101000",
  45065=>"110100101",
  45066=>"011001110",
  45067=>"000100111",
  45068=>"111111110",
  45069=>"000110110",
  45070=>"110000000",
  45071=>"111001001",
  45072=>"111111110",
  45073=>"000000111",
  45074=>"010000001",
  45075=>"000000000",
  45076=>"111000111",
  45077=>"111111111",
  45078=>"110111110",
  45079=>"111000000",
  45080=>"000001001",
  45081=>"010100111",
  45082=>"111111000",
  45083=>"001000100",
  45084=>"101110111",
  45085=>"011111111",
  45086=>"111010000",
  45087=>"111011000",
  45088=>"000100111",
  45089=>"111010111",
  45090=>"111010101",
  45091=>"111001001",
  45092=>"111100110",
  45093=>"111001100",
  45094=>"010010110",
  45095=>"000010111",
  45096=>"111110110",
  45097=>"000110001",
  45098=>"001111000",
  45099=>"001000011",
  45100=>"000000100",
  45101=>"111100001",
  45102=>"111111110",
  45103=>"111001100",
  45104=>"000010000",
  45105=>"111010110",
  45106=>"111111111",
  45107=>"001000000",
  45108=>"000110111",
  45109=>"010010111",
  45110=>"100000100",
  45111=>"111000000",
  45112=>"111001111",
  45113=>"000000000",
  45114=>"000101111",
  45115=>"101000010",
  45116=>"111110111",
  45117=>"111000001",
  45118=>"000000101",
  45119=>"111001000",
  45120=>"000111111",
  45121=>"001000001",
  45122=>"101101011",
  45123=>"111110001",
  45124=>"111111010",
  45125=>"001000000",
  45126=>"111101101",
  45127=>"011000000",
  45128=>"100111110",
  45129=>"011111101",
  45130=>"001011010",
  45131=>"100111011",
  45132=>"111111111",
  45133=>"010001001",
  45134=>"111011000",
  45135=>"111001011",
  45136=>"111111111",
  45137=>"111110000",
  45138=>"010111001",
  45139=>"000000110",
  45140=>"111000010",
  45141=>"111011110",
  45142=>"111100000",
  45143=>"001000010",
  45144=>"111111000",
  45145=>"111011111",
  45146=>"001111001",
  45147=>"000101111",
  45148=>"000000011",
  45149=>"100111111",
  45150=>"110000110",
  45151=>"111011111",
  45152=>"111101000",
  45153=>"011111111",
  45154=>"011101111",
  45155=>"110100110",
  45156=>"000011101",
  45157=>"011001010",
  45158=>"000000111",
  45159=>"111110000",
  45160=>"111111111",
  45161=>"111000100",
  45162=>"101111000",
  45163=>"111001001",
  45164=>"011000111",
  45165=>"000100101",
  45166=>"000111111",
  45167=>"110111111",
  45168=>"000010011",
  45169=>"111010111",
  45170=>"011000000",
  45171=>"011000000",
  45172=>"111111111",
  45173=>"101000001",
  45174=>"000111100",
  45175=>"000101110",
  45176=>"000111111",
  45177=>"000000100",
  45178=>"111111001",
  45179=>"001000001",
  45180=>"111011100",
  45181=>"000000101",
  45182=>"000000000",
  45183=>"000100101",
  45184=>"000000010",
  45185=>"111111101",
  45186=>"110101111",
  45187=>"000010110",
  45188=>"000000100",
  45189=>"111011010",
  45190=>"100100010",
  45191=>"111010111",
  45192=>"011001000",
  45193=>"011000110",
  45194=>"000000011",
  45195=>"000000000",
  45196=>"111111110",
  45197=>"001000011",
  45198=>"111000000",
  45199=>"000010110",
  45200=>"111110011",
  45201=>"000001011",
  45202=>"110110111",
  45203=>"000001101",
  45204=>"000000000",
  45205=>"111111111",
  45206=>"000000111",
  45207=>"000111100",
  45208=>"101100110",
  45209=>"111111111",
  45210=>"111000100",
  45211=>"101000011",
  45212=>"111110010",
  45213=>"000100111",
  45214=>"100111100",
  45215=>"111000000",
  45216=>"111110100",
  45217=>"110001000",
  45218=>"111111111",
  45219=>"010010000",
  45220=>"001000101",
  45221=>"110010110",
  45222=>"110111000",
  45223=>"000000111",
  45224=>"001000000",
  45225=>"111111000",
  45226=>"100101100",
  45227=>"000010111",
  45228=>"011000000",
  45229=>"000000000",
  45230=>"111111011",
  45231=>"010011010",
  45232=>"011001000",
  45233=>"101111101",
  45234=>"000000111",
  45235=>"110011111",
  45236=>"111101010",
  45237=>"111101111",
  45238=>"001100111",
  45239=>"100101010",
  45240=>"110111111",
  45241=>"001001000",
  45242=>"000100000",
  45243=>"000000000",
  45244=>"010000010",
  45245=>"111111000",
  45246=>"011001000",
  45247=>"011000000",
  45248=>"000110111",
  45249=>"010000001",
  45250=>"111011001",
  45251=>"110110111",
  45252=>"110111111",
  45253=>"111010110",
  45254=>"110010111",
  45255=>"011011100",
  45256=>"001101111",
  45257=>"111000000",
  45258=>"011111111",
  45259=>"001000110",
  45260=>"000100111",
  45261=>"111110000",
  45262=>"000111111",
  45263=>"111000000",
  45264=>"000000000",
  45265=>"100011011",
  45266=>"100100000",
  45267=>"111001110",
  45268=>"001101010",
  45269=>"000011011",
  45270=>"111111111",
  45271=>"110111111",
  45272=>"111010011",
  45273=>"000010010",
  45274=>"110000011",
  45275=>"111000000",
  45276=>"011110011",
  45277=>"111111100",
  45278=>"110111011",
  45279=>"111110110",
  45280=>"111010111",
  45281=>"110101000",
  45282=>"011000000",
  45283=>"111000000",
  45284=>"111111000",
  45285=>"111000001",
  45286=>"111001001",
  45287=>"110111111",
  45288=>"011111101",
  45289=>"001000100",
  45290=>"100110110",
  45291=>"010100000",
  45292=>"111001010",
  45293=>"011000001",
  45294=>"011000000",
  45295=>"111001001",
  45296=>"111000000",
  45297=>"010001001",
  45298=>"000000001",
  45299=>"000100111",
  45300=>"000100100",
  45301=>"010100000",
  45302=>"000001100",
  45303=>"111001111",
  45304=>"111111111",
  45305=>"111111111",
  45306=>"111111000",
  45307=>"000011100",
  45308=>"111000011",
  45309=>"000000000",
  45310=>"100100111",
  45311=>"000000110",
  45312=>"110100100",
  45313=>"110111100",
  45314=>"101001001",
  45315=>"010001000",
  45316=>"111101100",
  45317=>"110000110",
  45318=>"000010100",
  45319=>"111011100",
  45320=>"000000111",
  45321=>"110000011",
  45322=>"101000100",
  45323=>"111010111",
  45324=>"100001011",
  45325=>"000000100",
  45326=>"110111000",
  45327=>"000000100",
  45328=>"011010011",
  45329=>"011011100",
  45330=>"000000100",
  45331=>"011100001",
  45332=>"111110000",
  45333=>"111111111",
  45334=>"110110010",
  45335=>"101111101",
  45336=>"100000000",
  45337=>"001010100",
  45338=>"000111110",
  45339=>"101111000",
  45340=>"110100100",
  45341=>"001001011",
  45342=>"100110001",
  45343=>"001000100",
  45344=>"001110110",
  45345=>"110010010",
  45346=>"010100110",
  45347=>"011110100",
  45348=>"001000100",
  45349=>"100100110",
  45350=>"001001100",
  45351=>"100001011",
  45352=>"110111110",
  45353=>"000110100",
  45354=>"001111000",
  45355=>"011010000",
  45356=>"011111110",
  45357=>"010000100",
  45358=>"100110110",
  45359=>"011111100",
  45360=>"110111111",
  45361=>"001001010",
  45362=>"100101111",
  45363=>"000011011",
  45364=>"100100111",
  45365=>"011111110",
  45366=>"000110110",
  45367=>"000001011",
  45368=>"000010000",
  45369=>"000000011",
  45370=>"010000000",
  45371=>"101001011",
  45372=>"000001110",
  45373=>"110000110",
  45374=>"000010000",
  45375=>"000111000",
  45376=>"101000001",
  45377=>"110110100",
  45378=>"111001010",
  45379=>"101100000",
  45380=>"011000000",
  45381=>"000000011",
  45382=>"101010110",
  45383=>"000011100",
  45384=>"101111111",
  45385=>"001010001",
  45386=>"000000101",
  45387=>"110101001",
  45388=>"100100110",
  45389=>"111110100",
  45390=>"001001100",
  45391=>"110110111",
  45392=>"010110100",
  45393=>"000111111",
  45394=>"111100100",
  45395=>"010010110",
  45396=>"000001001",
  45397=>"110010100",
  45398=>"001100100",
  45399=>"100111001",
  45400=>"000000100",
  45401=>"001111110",
  45402=>"000100110",
  45403=>"100110111",
  45404=>"100001001",
  45405=>"011011001",
  45406=>"111000011",
  45407=>"000111000",
  45408=>"000000010",
  45409=>"001011001",
  45410=>"100000001",
  45411=>"011111110",
  45412=>"001100100",
  45413=>"001101001",
  45414=>"000110001",
  45415=>"000100110",
  45416=>"001001011",
  45417=>"100110000",
  45418=>"100000001",
  45419=>"100000001",
  45420=>"101111110",
  45421=>"001010000",
  45422=>"000000000",
  45423=>"100111111",
  45424=>"011001101",
  45425=>"110001001",
  45426=>"111110110",
  45427=>"101001001",
  45428=>"000000000",
  45429=>"100000100",
  45430=>"110011011",
  45431=>"000100001",
  45432=>"000110010",
  45433=>"000000001",
  45434=>"001000011",
  45435=>"100101001",
  45436=>"000001111",
  45437=>"001110100",
  45438=>"000000000",
  45439=>"011111110",
  45440=>"000110100",
  45441=>"000000100",
  45442=>"100000100",
  45443=>"100110011",
  45444=>"011001001",
  45445=>"001100110",
  45446=>"110100100",
  45447=>"011001001",
  45448=>"001101111",
  45449=>"011100100",
  45450=>"101100100",
  45451=>"000001001",
  45452=>"110001010",
  45453=>"000100101",
  45454=>"011111001",
  45455=>"000000000",
  45456=>"000010110",
  45457=>"110110110",
  45458=>"010100110",
  45459=>"001011011",
  45460=>"011011011",
  45461=>"110001000",
  45462=>"010111111",
  45463=>"000110111",
  45464=>"100100110",
  45465=>"011100110",
  45466=>"010100000",
  45467=>"001001101",
  45468=>"010100111",
  45469=>"011011111",
  45470=>"100110111",
  45471=>"001000000",
  45472=>"100111111",
  45473=>"111011101",
  45474=>"000110111",
  45475=>"110110101",
  45476=>"000000000",
  45477=>"000000100",
  45478=>"101101100",
  45479=>"001110110",
  45480=>"100001011",
  45481=>"110100001",
  45482=>"111001100",
  45483=>"111110000",
  45484=>"111001111",
  45485=>"111101011",
  45486=>"001110111",
  45487=>"001000110",
  45488=>"010011011",
  45489=>"000011110",
  45490=>"001111111",
  45491=>"000000110",
  45492=>"101011110",
  45493=>"100011110",
  45494=>"110100001",
  45495=>"111111100",
  45496=>"011011100",
  45497=>"000001011",
  45498=>"110110110",
  45499=>"000000100",
  45500=>"011100000",
  45501=>"000100110",
  45502=>"011011000",
  45503=>"011011010",
  45504=>"001000011",
  45505=>"000000000",
  45506=>"100100100",
  45507=>"001111010",
  45508=>"000010011",
  45509=>"111001000",
  45510=>"100111000",
  45511=>"100010111",
  45512=>"001001010",
  45513=>"000111010",
  45514=>"111011101",
  45515=>"110000010",
  45516=>"001000110",
  45517=>"011011001",
  45518=>"011011011",
  45519=>"000011011",
  45520=>"111110100",
  45521=>"011111100",
  45522=>"001000011",
  45523=>"110100000",
  45524=>"101000100",
  45525=>"111111000",
  45526=>"000010000",
  45527=>"100111001",
  45528=>"001001100",
  45529=>"100000100",
  45530=>"111101100",
  45531=>"111000001",
  45532=>"011011011",
  45533=>"110010110",
  45534=>"110101000",
  45535=>"101101010",
  45536=>"000000110",
  45537=>"100001111",
  45538=>"100100001",
  45539=>"001111110",
  45540=>"000000000",
  45541=>"111110111",
  45542=>"001011001",
  45543=>"101101001",
  45544=>"111000110",
  45545=>"100100001",
  45546=>"111100000",
  45547=>"110001111",
  45548=>"000000000",
  45549=>"100000000",
  45550=>"000000100",
  45551=>"000000001",
  45552=>"011001011",
  45553=>"000010111",
  45554=>"110110010",
  45555=>"111001000",
  45556=>"001001111",
  45557=>"000000000",
  45558=>"000000110",
  45559=>"011011011",
  45560=>"110011001",
  45561=>"001110000",
  45562=>"000000100",
  45563=>"001001000",
  45564=>"111110110",
  45565=>"100011000",
  45566=>"101001101",
  45567=>"001110010",
  45568=>"011001000",
  45569=>"000111110",
  45570=>"000000100",
  45571=>"010110111",
  45572=>"000101000",
  45573=>"110010010",
  45574=>"000001001",
  45575=>"011111010",
  45576=>"000111110",
  45577=>"000000001",
  45578=>"000000010",
  45579=>"000100011",
  45580=>"000000010",
  45581=>"010010000",
  45582=>"000000001",
  45583=>"000001011",
  45584=>"011111010",
  45585=>"000000000",
  45586=>"101101101",
  45587=>"000011010",
  45588=>"000001010",
  45589=>"000011010",
  45590=>"000111010",
  45591=>"111111111",
  45592=>"111000100",
  45593=>"011111011",
  45594=>"111111011",
  45595=>"010111010",
  45596=>"111001111",
  45597=>"000000000",
  45598=>"110100000",
  45599=>"000000010",
  45600=>"000000000",
  45601=>"010111111",
  45602=>"111101111",
  45603=>"010111010",
  45604=>"001111011",
  45605=>"110111001",
  45606=>"010010010",
  45607=>"000110000",
  45608=>"010011010",
  45609=>"100110110",
  45610=>"000011111",
  45611=>"010000000",
  45612=>"110111011",
  45613=>"010100010",
  45614=>"111010000",
  45615=>"000101011",
  45616=>"010111000",
  45617=>"000101000",
  45618=>"001001100",
  45619=>"111000011",
  45620=>"000000001",
  45621=>"010111011",
  45622=>"000011011",
  45623=>"000000000",
  45624=>"000010010",
  45625=>"001000011",
  45626=>"001001010",
  45627=>"011000000",
  45628=>"010110111",
  45629=>"111111111",
  45630=>"000000101",
  45631=>"110110110",
  45632=>"000101111",
  45633=>"101001000",
  45634=>"010010010",
  45635=>"001110000",
  45636=>"101111010",
  45637=>"111010000",
  45638=>"111001110",
  45639=>"111101101",
  45640=>"000001010",
  45641=>"110111010",
  45642=>"111010011",
  45643=>"110000111",
  45644=>"101100101",
  45645=>"010011010",
  45646=>"000001000",
  45647=>"111010011",
  45648=>"000010111",
  45649=>"111111111",
  45650=>"110011110",
  45651=>"011111010",
  45652=>"001000001",
  45653=>"000100000",
  45654=>"000111110",
  45655=>"111111011",
  45656=>"110011111",
  45657=>"000010001",
  45658=>"000010010",
  45659=>"000111010",
  45660=>"000001010",
  45661=>"000001111",
  45662=>"010010000",
  45663=>"000010010",
  45664=>"010110010",
  45665=>"010111111",
  45666=>"001000101",
  45667=>"000011010",
  45668=>"010010110",
  45669=>"010011000",
  45670=>"000000000",
  45671=>"000010111",
  45672=>"010011010",
  45673=>"011001000",
  45674=>"000010010",
  45675=>"000010110",
  45676=>"011011111",
  45677=>"001001010",
  45678=>"000000001",
  45679=>"000011110",
  45680=>"000111110",
  45681=>"000010010",
  45682=>"001100110",
  45683=>"000000010",
  45684=>"000010010",
  45685=>"101000101",
  45686=>"010111010",
  45687=>"010110110",
  45688=>"010010000",
  45689=>"010011010",
  45690=>"000001010",
  45691=>"010111010",
  45692=>"100100110",
  45693=>"110111000",
  45694=>"010111001",
  45695=>"100111111",
  45696=>"101101000",
  45697=>"110100000",
  45698=>"010010010",
  45699=>"010000001",
  45700=>"110010010",
  45701=>"000101011",
  45702=>"011100000",
  45703=>"011111011",
  45704=>"000111001",
  45705=>"011011010",
  45706=>"001010011",
  45707=>"000100101",
  45708=>"001010000",
  45709=>"000000010",
  45710=>"011111111",
  45711=>"101000101",
  45712=>"000001100",
  45713=>"110111001",
  45714=>"011000111",
  45715=>"000110011",
  45716=>"110111011",
  45717=>"000000010",
  45718=>"010111010",
  45719=>"110111011",
  45720=>"010111001",
  45721=>"111111000",
  45722=>"000010010",
  45723=>"000000000",
  45724=>"000000010",
  45725=>"111010010",
  45726=>"010111010",
  45727=>"101000101",
  45728=>"010010000",
  45729=>"000010010",
  45730=>"010110110",
  45731=>"110111111",
  45732=>"010000011",
  45733=>"010011010",
  45734=>"001011011",
  45735=>"000000101",
  45736=>"000111110",
  45737=>"000111110",
  45738=>"000000000",
  45739=>"000000100",
  45740=>"101000111",
  45741=>"000000101",
  45742=>"110110010",
  45743=>"011010010",
  45744=>"101101101",
  45745=>"010011110",
  45746=>"000101110",
  45747=>"000000110",
  45748=>"010111010",
  45749=>"010111111",
  45750=>"111111100",
  45751=>"000000001",
  45752=>"011010011",
  45753=>"011010011",
  45754=>"110000110",
  45755=>"011010110",
  45756=>"101001001",
  45757=>"111111100",
  45758=>"001011011",
  45759=>"010000010",
  45760=>"000011010",
  45761=>"000000110",
  45762=>"011111010",
  45763=>"111111100",
  45764=>"001001000",
  45765=>"110110110",
  45766=>"010010011",
  45767=>"000000000",
  45768=>"111111111",
  45769=>"011111000",
  45770=>"111001100",
  45771=>"000010000",
  45772=>"010011000",
  45773=>"000000001",
  45774=>"010000111",
  45775=>"110110000",
  45776=>"010100110",
  45777=>"010111010",
  45778=>"111011011",
  45779=>"010011010",
  45780=>"000001010",
  45781=>"100111111",
  45782=>"000000010",
  45783=>"110101010",
  45784=>"000011010",
  45785=>"010001010",
  45786=>"100000100",
  45787=>"001000000",
  45788=>"010110000",
  45789=>"111011010",
  45790=>"010010010",
  45791=>"010000010",
  45792=>"010000000",
  45793=>"101000010",
  45794=>"010111000",
  45795=>"010111000",
  45796=>"000000010",
  45797=>"000010010",
  45798=>"010000000",
  45799=>"000111110",
  45800=>"010010010",
  45801=>"010111010",
  45802=>"000000110",
  45803=>"000000110",
  45804=>"010010000",
  45805=>"001111111",
  45806=>"010101010",
  45807=>"010000011",
  45808=>"010010010",
  45809=>"011101100",
  45810=>"110111011",
  45811=>"010011000",
  45812=>"110010010",
  45813=>"001000010",
  45814=>"001000010",
  45815=>"000101100",
  45816=>"000010010",
  45817=>"000010011",
  45818=>"000000010",
  45819=>"000001000",
  45820=>"010111010",
  45821=>"000000000",
  45822=>"000101000",
  45823=>"000000010",
  45824=>"011010111",
  45825=>"100111011",
  45826=>"011100101",
  45827=>"010111010",
  45828=>"110110110",
  45829=>"000010100",
  45830=>"100101101",
  45831=>"111111101",
  45832=>"110010000",
  45833=>"111101101",
  45834=>"010001001",
  45835=>"101111110",
  45836=>"100000000",
  45837=>"000000000",
  45838=>"111110110",
  45839=>"111111111",
  45840=>"001101101",
  45841=>"111110000",
  45842=>"000011011",
  45843=>"001000000",
  45844=>"101101000",
  45845=>"111111010",
  45846=>"011111000",
  45847=>"001101101",
  45848=>"001001000",
  45849=>"000000110",
  45850=>"111111010",
  45851=>"111100100",
  45852=>"100100100",
  45853=>"000111010",
  45854=>"000111111",
  45855=>"111111000",
  45856=>"111101001",
  45857=>"110111100",
  45858=>"111111111",
  45859=>"011111010",
  45860=>"001111111",
  45861=>"000001111",
  45862=>"010011000",
  45863=>"111101111",
  45864=>"100101010",
  45865=>"111111000",
  45866=>"111111000",
  45867=>"000010111",
  45868=>"100110100",
  45869=>"010011010",
  45870=>"101111111",
  45871=>"101000001",
  45872=>"000100000",
  45873=>"100110100",
  45874=>"101010111",
  45875=>"011000000",
  45876=>"001101101",
  45877=>"010101000",
  45878=>"011011001",
  45879=>"110010110",
  45880=>"000000010",
  45881=>"111111000",
  45882=>"100001001",
  45883=>"101001100",
  45884=>"100111000",
  45885=>"000011111",
  45886=>"101000000",
  45887=>"001000001",
  45888=>"111111000",
  45889=>"000010111",
  45890=>"111110100",
  45891=>"111111110",
  45892=>"101000001",
  45893=>"100010000",
  45894=>"000000100",
  45895=>"010111000",
  45896=>"011111001",
  45897=>"110100000",
  45898=>"111111111",
  45899=>"111001000",
  45900=>"010111111",
  45901=>"000111010",
  45902=>"011011001",
  45903=>"000000000",
  45904=>"111000110",
  45905=>"000111111",
  45906=>"000111110",
  45907=>"100111010",
  45908=>"111101010",
  45909=>"011011011",
  45910=>"001011010",
  45911=>"111101001",
  45912=>"110111100",
  45913=>"000110000",
  45914=>"010011010",
  45915=>"001101000",
  45916=>"111111000",
  45917=>"100100000",
  45918=>"111101000",
  45919=>"111111111",
  45920=>"111111111",
  45921=>"111111110",
  45922=>"001000000",
  45923=>"010010000",
  45924=>"101111000",
  45925=>"111100000",
  45926=>"111111101",
  45927=>"111001101",
  45928=>"110101000",
  45929=>"001111111",
  45930=>"000010000",
  45931=>"000011000",
  45932=>"000010000",
  45933=>"111111000",
  45934=>"000011000",
  45935=>"101000100",
  45936=>"111111000",
  45937=>"111011111",
  45938=>"111111100",
  45939=>"111111000",
  45940=>"001111000",
  45941=>"111011110",
  45942=>"111001000",
  45943=>"000111011",
  45944=>"000000000",
  45945=>"011101000",
  45946=>"010000101",
  45947=>"000111000",
  45948=>"110010100",
  45949=>"100011000",
  45950=>"000000000",
  45951=>"001000000",
  45952=>"100000111",
  45953=>"000000100",
  45954=>"101111000",
  45955=>"000111110",
  45956=>"011111011",
  45957=>"001010000",
  45958=>"011110011",
  45959=>"111101000",
  45960=>"000111100",
  45961=>"111101110",
  45962=>"111101000",
  45963=>"100111111",
  45964=>"110111110",
  45965=>"000000001",
  45966=>"000101000",
  45967=>"000010000",
  45968=>"001011110",
  45969=>"100101000",
  45970=>"011011010",
  45971=>"111000000",
  45972=>"011111000",
  45973=>"000101000",
  45974=>"101101000",
  45975=>"011011000",
  45976=>"000000000",
  45977=>"000000111",
  45978=>"011001000",
  45979=>"000000000",
  45980=>"101111010",
  45981=>"100100000",
  45982=>"011011101",
  45983=>"110100000",
  45984=>"110110010",
  45985=>"111101000",
  45986=>"111001000",
  45987=>"011111111",
  45988=>"000110000",
  45989=>"000111000",
  45990=>"110111111",
  45991=>"001100101",
  45992=>"101000010",
  45993=>"101010010",
  45994=>"011011011",
  45995=>"000010000",
  45996=>"100000111",
  45997=>"010011010",
  45998=>"110011011",
  45999=>"000100000",
  46000=>"100100111",
  46001=>"111111101",
  46002=>"000010000",
  46003=>"010011000",
  46004=>"000100000",
  46005=>"111000000",
  46006=>"011001001",
  46007=>"010000001",
  46008=>"101110100",
  46009=>"110110100",
  46010=>"000000101",
  46011=>"010101000",
  46012=>"111011010",
  46013=>"011000101",
  46014=>"011110100",
  46015=>"111101111",
  46016=>"101111000",
  46017=>"011011010",
  46018=>"100111000",
  46019=>"000100110",
  46020=>"111101111",
  46021=>"010011111",
  46022=>"011111000",
  46023=>"111111101",
  46024=>"110111111",
  46025=>"101100111",
  46026=>"011010010",
  46027=>"111111010",
  46028=>"111110000",
  46029=>"010000001",
  46030=>"000000000",
  46031=>"000000100",
  46032=>"011001111",
  46033=>"000000000",
  46034=>"101000011",
  46035=>"111111011",
  46036=>"001111000",
  46037=>"110000000",
  46038=>"010110000",
  46039=>"100101000",
  46040=>"100100000",
  46041=>"000000000",
  46042=>"111001011",
  46043=>"111000101",
  46044=>"100111100",
  46045=>"000001101",
  46046=>"111011001",
  46047=>"010100001",
  46048=>"100100000",
  46049=>"111101101",
  46050=>"010011001",
  46051=>"111111000",
  46052=>"111101001",
  46053=>"000111000",
  46054=>"101000000",
  46055=>"111110010",
  46056=>"111010000",
  46057=>"111111001",
  46058=>"100100000",
  46059=>"111011100",
  46060=>"010000111",
  46061=>"110111111",
  46062=>"000111011",
  46063=>"011011000",
  46064=>"010111010",
  46065=>"110101011",
  46066=>"101111000",
  46067=>"101111000",
  46068=>"111111010",
  46069=>"001001101",
  46070=>"001010010",
  46071=>"111011111",
  46072=>"100100000",
  46073=>"000110000",
  46074=>"000111010",
  46075=>"010100000",
  46076=>"010010010",
  46077=>"010010000",
  46078=>"011011001",
  46079=>"101010000",
  46080=>"000000011",
  46081=>"010000111",
  46082=>"101101000",
  46083=>"111101101",
  46084=>"111111010",
  46085=>"001001000",
  46086=>"110010011",
  46087=>"010010111",
  46088=>"000000111",
  46089=>"000111111",
  46090=>"100011000",
  46091=>"100111011",
  46092=>"000111101",
  46093=>"011011111",
  46094=>"111010011",
  46095=>"000100101",
  46096=>"000010110",
  46097=>"001111010",
  46098=>"110111000",
  46099=>"100100111",
  46100=>"101010110",
  46101=>"111111010",
  46102=>"101100111",
  46103=>"000000101",
  46104=>"101101101",
  46105=>"110110111",
  46106=>"111000111",
  46107=>"111011111",
  46108=>"110101101",
  46109=>"101111101",
  46110=>"010100101",
  46111=>"001100000",
  46112=>"110010010",
  46113=>"111011111",
  46114=>"111001000",
  46115=>"111101001",
  46116=>"001011000",
  46117=>"000000100",
  46118=>"111000111",
  46119=>"001111001",
  46120=>"111000011",
  46121=>"111010010",
  46122=>"111001111",
  46123=>"011011111",
  46124=>"111001001",
  46125=>"101001101",
  46126=>"111111000",
  46127=>"000000000",
  46128=>"000000000",
  46129=>"111101101",
  46130=>"101100100",
  46131=>"111000000",
  46132=>"000000111",
  46133=>"101101111",
  46134=>"000100110",
  46135=>"000111111",
  46136=>"000111101",
  46137=>"011101100",
  46138=>"010110000",
  46139=>"110000000",
  46140=>"110001001",
  46141=>"000110011",
  46142=>"000101101",
  46143=>"011010001",
  46144=>"000000111",
  46145=>"010110111",
  46146=>"001010101",
  46147=>"000100101",
  46148=>"000000000",
  46149=>"000001101",
  46150=>"110010101",
  46151=>"001100011",
  46152=>"000000101",
  46153=>"111000000",
  46154=>"000010001",
  46155=>"000011111",
  46156=>"001111010",
  46157=>"101111010",
  46158=>"001010010",
  46159=>"001110000",
  46160=>"111010010",
  46161=>"101000011",
  46162=>"011000010",
  46163=>"000001011",
  46164=>"000111111",
  46165=>"000000101",
  46166=>"011001011",
  46167=>"101111111",
  46168=>"110110000",
  46169=>"110110110",
  46170=>"011000000",
  46171=>"110110000",
  46172=>"010110111",
  46173=>"011001001",
  46174=>"100000101",
  46175=>"000001101",
  46176=>"010010111",
  46177=>"100110010",
  46178=>"000011111",
  46179=>"110100000",
  46180=>"111111000",
  46181=>"111011111",
  46182=>"010000000",
  46183=>"111111100",
  46184=>"010111101",
  46185=>"101100000",
  46186=>"000010010",
  46187=>"010011111",
  46188=>"010111000",
  46189=>"111111000",
  46190=>"000001000",
  46191=>"000010101",
  46192=>"110110010",
  46193=>"000110000",
  46194=>"000000011",
  46195=>"111101101",
  46196=>"000000010",
  46197=>"000001011",
  46198=>"111001111",
  46199=>"000111111",
  46200=>"000001001",
  46201=>"010010101",
  46202=>"110000000",
  46203=>"101101000",
  46204=>"001111111",
  46205=>"110100100",
  46206=>"010111111",
  46207=>"111011000",
  46208=>"000000001",
  46209=>"000101100",
  46210=>"111100101",
  46211=>"111111000",
  46212=>"000010010",
  46213=>"010000100",
  46214=>"001000101",
  46215=>"011000001",
  46216=>"111010000",
  46217=>"111000000",
  46218=>"110110111",
  46219=>"000000001",
  46220=>"111001000",
  46221=>"000101100",
  46222=>"010000101",
  46223=>"010000110",
  46224=>"011011011",
  46225=>"000100010",
  46226=>"001001000",
  46227=>"000011111",
  46228=>"111000000",
  46229=>"101101101",
  46230=>"110000101",
  46231=>"100000011",
  46232=>"100011101",
  46233=>"101001110",
  46234=>"101100010",
  46235=>"010101100",
  46236=>"001101111",
  46237=>"110111010",
  46238=>"001100000",
  46239=>"100011111",
  46240=>"001000101",
  46241=>"001001111",
  46242=>"111011101",
  46243=>"111111000",
  46244=>"110110000",
  46245=>"010011001",
  46246=>"101001001",
  46247=>"000010111",
  46248=>"100111111",
  46249=>"001000010",
  46250=>"101000010",
  46251=>"001001010",
  46252=>"011000101",
  46253=>"011110010",
  46254=>"001111011",
  46255=>"111111101",
  46256=>"010001001",
  46257=>"111011001",
  46258=>"101111111",
  46259=>"001011101",
  46260=>"111111101",
  46261=>"111111101",
  46262=>"100000100",
  46263=>"101000011",
  46264=>"011100100",
  46265=>"110010110",
  46266=>"000000001",
  46267=>"000111100",
  46268=>"111100000",
  46269=>"110111111",
  46270=>"000111011",
  46271=>"111111101",
  46272=>"000010000",
  46273=>"000000001",
  46274=>"000001111",
  46275=>"111111001",
  46276=>"000000000",
  46277=>"001001000",
  46278=>"000100110",
  46279=>"001000100",
  46280=>"111000000",
  46281=>"001001111",
  46282=>"100011101",
  46283=>"101001111",
  46284=>"000100101",
  46285=>"100111111",
  46286=>"100111111",
  46287=>"000111000",
  46288=>"111111010",
  46289=>"011010000",
  46290=>"011111111",
  46291=>"000000000",
  46292=>"100000010",
  46293=>"110100100",
  46294=>"101111000",
  46295=>"011011111",
  46296=>"000100101",
  46297=>"000000110",
  46298=>"111010101",
  46299=>"111000000",
  46300=>"000000000",
  46301=>"001100000",
  46302=>"100110101",
  46303=>"001000111",
  46304=>"011111111",
  46305=>"101101000",
  46306=>"111000000",
  46307=>"111011100",
  46308=>"000001010",
  46309=>"000000000",
  46310=>"110011111",
  46311=>"010111111",
  46312=>"000010000",
  46313=>"111100000",
  46314=>"000010010",
  46315=>"010101111",
  46316=>"000010111",
  46317=>"000000000",
  46318=>"100010010",
  46319=>"000000000",
  46320=>"010100100",
  46321=>"100100001",
  46322=>"100111001",
  46323=>"110000001",
  46324=>"000000111",
  46325=>"111000000",
  46326=>"000100001",
  46327=>"111111001",
  46328=>"000001111",
  46329=>"000100100",
  46330=>"111110011",
  46331=>"011110101",
  46332=>"000010110",
  46333=>"110101001",
  46334=>"011000101",
  46335=>"011111111",
  46336=>"101000000",
  46337=>"000000111",
  46338=>"000000000",
  46339=>"001101111",
  46340=>"110001010",
  46341=>"001001000",
  46342=>"010100100",
  46343=>"000111111",
  46344=>"111001001",
  46345=>"111000000",
  46346=>"000000100",
  46347=>"010000101",
  46348=>"010010111",
  46349=>"111000111",
  46350=>"001010010",
  46351=>"000000000",
  46352=>"000001000",
  46353=>"101000101",
  46354=>"000110111",
  46355=>"111000100",
  46356=>"100000110",
  46357=>"000010010",
  46358=>"000101111",
  46359=>"010000000",
  46360=>"101000001",
  46361=>"000000000",
  46362=>"000000100",
  46363=>"110111110",
  46364=>"110111001",
  46365=>"111000001",
  46366=>"101110011",
  46367=>"111101111",
  46368=>"000000000",
  46369=>"000000111",
  46370=>"100101100",
  46371=>"000101111",
  46372=>"001001000",
  46373=>"010110001",
  46374=>"000111010",
  46375=>"010111111",
  46376=>"111000000",
  46377=>"000111111",
  46378=>"000011000",
  46379=>"100000000",
  46380=>"000111111",
  46381=>"011111000",
  46382=>"111010111",
  46383=>"101110001",
  46384=>"001111001",
  46385=>"111010000",
  46386=>"100100110",
  46387=>"111111101",
  46388=>"000000101",
  46389=>"101101001",
  46390=>"100100001",
  46391=>"101111001",
  46392=>"000110000",
  46393=>"101001111",
  46394=>"111101111",
  46395=>"101111010",
  46396=>"000111110",
  46397=>"010111111",
  46398=>"101100100",
  46399=>"011001111",
  46400=>"101000010",
  46401=>"110010111",
  46402=>"100111111",
  46403=>"000000000",
  46404=>"011000000",
  46405=>"110001000",
  46406=>"110000001",
  46407=>"100110101",
  46408=>"000111111",
  46409=>"010000110",
  46410=>"101101101",
  46411=>"111111011",
  46412=>"101110010",
  46413=>"110100000",
  46414=>"010011100",
  46415=>"111000000",
  46416=>"101101101",
  46417=>"010111111",
  46418=>"010010111",
  46419=>"110010110",
  46420=>"011000110",
  46421=>"001100100",
  46422=>"100111011",
  46423=>"001000100",
  46424=>"001101111",
  46425=>"110110000",
  46426=>"000110111",
  46427=>"111100100",
  46428=>"000100111",
  46429=>"010000000",
  46430=>"111111000",
  46431=>"100100000",
  46432=>"000110111",
  46433=>"010000000",
  46434=>"111111110",
  46435=>"001111101",
  46436=>"000100010",
  46437=>"010110000",
  46438=>"100000000",
  46439=>"100011000",
  46440=>"001000010",
  46441=>"011100000",
  46442=>"111111000",
  46443=>"000110110",
  46444=>"000110110",
  46445=>"000000010",
  46446=>"111110111",
  46447=>"111010000",
  46448=>"101111010",
  46449=>"010010010",
  46450=>"001001100",
  46451=>"101101001",
  46452=>"000011010",
  46453=>"111001000",
  46454=>"110100111",
  46455=>"000010000",
  46456=>"011111110",
  46457=>"110010000",
  46458=>"110001001",
  46459=>"000000000",
  46460=>"101000100",
  46461=>"111100100",
  46462=>"111000110",
  46463=>"111000000",
  46464=>"000000000",
  46465=>"000000010",
  46466=>"111101000",
  46467=>"110010101",
  46468=>"010000111",
  46469=>"111101001",
  46470=>"110111110",
  46471=>"000000000",
  46472=>"000110000",
  46473=>"000111010",
  46474=>"010000000",
  46475=>"111101000",
  46476=>"111001000",
  46477=>"000000001",
  46478=>"110010000",
  46479=>"001001000",
  46480=>"010111001",
  46481=>"000000010",
  46482=>"000101110",
  46483=>"110000110",
  46484=>"111111010",
  46485=>"001000000",
  46486=>"000111111",
  46487=>"010010010",
  46488=>"010111101",
  46489=>"101111111",
  46490=>"111000000",
  46491=>"000100010",
  46492=>"010101000",
  46493=>"001101000",
  46494=>"101101000",
  46495=>"000111110",
  46496=>"100001011",
  46497=>"110100001",
  46498=>"110000010",
  46499=>"000101110",
  46500=>"111011110",
  46501=>"001001000",
  46502=>"011111010",
  46503=>"011110111",
  46504=>"111000110",
  46505=>"000000111",
  46506=>"111000111",
  46507=>"111110101",
  46508=>"111111010",
  46509=>"111100000",
  46510=>"100101101",
  46511=>"010001000",
  46512=>"010110111",
  46513=>"011011000",
  46514=>"110000000",
  46515=>"100011000",
  46516=>"111000001",
  46517=>"100111111",
  46518=>"000000100",
  46519=>"111000000",
  46520=>"011111111",
  46521=>"000010100",
  46522=>"111011000",
  46523=>"011111000",
  46524=>"100110011",
  46525=>"100000110",
  46526=>"100000100",
  46527=>"000000010",
  46528=>"111000000",
  46529=>"111000000",
  46530=>"000110011",
  46531=>"100000000",
  46532=>"000110011",
  46533=>"011111100",
  46534=>"000000111",
  46535=>"000110100",
  46536=>"010010000",
  46537=>"000110010",
  46538=>"000001000",
  46539=>"100000000",
  46540=>"111101000",
  46541=>"000100000",
  46542=>"111100000",
  46543=>"011011000",
  46544=>"111000101",
  46545=>"001111111",
  46546=>"011111010",
  46547=>"111101110",
  46548=>"010010000",
  46549=>"100100101",
  46550=>"000000111",
  46551=>"000111111",
  46552=>"001111000",
  46553=>"001000000",
  46554=>"011100011",
  46555=>"111000000",
  46556=>"100111011",
  46557=>"000000000",
  46558=>"000001101",
  46559=>"101000010",
  46560=>"110011000",
  46561=>"011001000",
  46562=>"111111101",
  46563=>"000001100",
  46564=>"000001000",
  46565=>"010000000",
  46566=>"111000110",
  46567=>"001111101",
  46568=>"100111111",
  46569=>"100000111",
  46570=>"111001000",
  46571=>"111000010",
  46572=>"000111111",
  46573=>"101001000",
  46574=>"000000010",
  46575=>"010100100",
  46576=>"111101111",
  46577=>"100011000",
  46578=>"111111010",
  46579=>"111111111",
  46580=>"011110111",
  46581=>"100000101",
  46582=>"011001000",
  46583=>"000111100",
  46584=>"111000000",
  46585=>"000001000",
  46586=>"111101101",
  46587=>"111111100",
  46588=>"100111111",
  46589=>"001000000",
  46590=>"111000000",
  46591=>"000110110",
  46592=>"011011010",
  46593=>"000000110",
  46594=>"000000000",
  46595=>"111111000",
  46596=>"100000100",
  46597=>"010110000",
  46598=>"110010111",
  46599=>"000111111",
  46600=>"111101001",
  46601=>"101101111",
  46602=>"100000000",
  46603=>"111111011",
  46604=>"010010011",
  46605=>"101101111",
  46606=>"110101011",
  46607=>"000000011",
  46608=>"100000000",
  46609=>"111111100",
  46610=>"110110000",
  46611=>"010000101",
  46612=>"111111111",
  46613=>"000000000",
  46614=>"011011011",
  46615=>"111110111",
  46616=>"000110100",
  46617=>"000000001",
  46618=>"000000000",
  46619=>"111111100",
  46620=>"111111110",
  46621=>"011101000",
  46622=>"110100000",
  46623=>"111111011",
  46624=>"000010010",
  46625=>"010011110",
  46626=>"100110101",
  46627=>"010111010",
  46628=>"110111000",
  46629=>"110100000",
  46630=>"111110110",
  46631=>"111010000",
  46632=>"101000111",
  46633=>"111111000",
  46634=>"111011110",
  46635=>"111111110",
  46636=>"110111000",
  46637=>"110010000",
  46638=>"010110111",
  46639=>"001000000",
  46640=>"101000100",
  46641=>"110100111",
  46642=>"110100111",
  46643=>"111011011",
  46644=>"111110001",
  46645=>"111111111",
  46646=>"111111110",
  46647=>"110000011",
  46648=>"111110111",
  46649=>"111000000",
  46650=>"101000100",
  46651=>"111111010",
  46652=>"100100111",
  46653=>"110111111",
  46654=>"101000111",
  46655=>"111101110",
  46656=>"111011111",
  46657=>"111000000",
  46658=>"110110100",
  46659=>"100100100",
  46660=>"111010010",
  46661=>"010000000",
  46662=>"000100111",
  46663=>"110110101",
  46664=>"000110110",
  46665=>"001001110",
  46666=>"000000011",
  46667=>"000000000",
  46668=>"000000000",
  46669=>"000111111",
  46670=>"010000000",
  46671=>"110111011",
  46672=>"111111111",
  46673=>"000111111",
  46674=>"000000010",
  46675=>"011001000",
  46676=>"001000000",
  46677=>"100010000",
  46678=>"001001101",
  46679=>"000000000",
  46680=>"000101111",
  46681=>"111111011",
  46682=>"111111110",
  46683=>"001000000",
  46684=>"000000000",
  46685=>"011001111",
  46686=>"111111010",
  46687=>"001111010",
  46688=>"001001110",
  46689=>"001100110",
  46690=>"000000001",
  46691=>"100111111",
  46692=>"101110000",
  46693=>"000000101",
  46694=>"000100101",
  46695=>"011011000",
  46696=>"000110100",
  46697=>"110001000",
  46698=>"110000110",
  46699=>"111000000",
  46700=>"111000000",
  46701=>"100110111",
  46702=>"000000011",
  46703=>"000001111",
  46704=>"101100000",
  46705=>"111111000",
  46706=>"111111111",
  46707=>"000000000",
  46708=>"111000000",
  46709=>"000000000",
  46710=>"000000101",
  46711=>"111111110",
  46712=>"001000111",
  46713=>"110101100",
  46714=>"010010111",
  46715=>"000110111",
  46716=>"100110011",
  46717=>"100100000",
  46718=>"111101110",
  46719=>"000001101",
  46720=>"010000000",
  46721=>"100100100",
  46722=>"000000100",
  46723=>"010000100",
  46724=>"111111111",
  46725=>"100000001",
  46726=>"111011001",
  46727=>"001011011",
  46728=>"011011111",
  46729=>"000000000",
  46730=>"000000000",
  46731=>"111000000",
  46732=>"000000000",
  46733=>"000011111",
  46734=>"111111111",
  46735=>"001000001",
  46736=>"101111001",
  46737=>"111111000",
  46738=>"000000110",
  46739=>"000000000",
  46740=>"000101111",
  46741=>"111111010",
  46742=>"000000000",
  46743=>"000110000",
  46744=>"010010100",
  46745=>"111111111",
  46746=>"000111110",
  46747=>"000000000",
  46748=>"110110000",
  46749=>"000111111",
  46750=>"110010010",
  46751=>"001001101",
  46752=>"000111001",
  46753=>"111110010",
  46754=>"111110000",
  46755=>"111101101",
  46756=>"111111111",
  46757=>"110100000",
  46758=>"111110111",
  46759=>"111110000",
  46760=>"000111111",
  46761=>"110000000",
  46762=>"000000111",
  46763=>"111101110",
  46764=>"110100000",
  46765=>"000000000",
  46766=>"100000011",
  46767=>"010010010",
  46768=>"011010100",
  46769=>"010010110",
  46770=>"000000000",
  46771=>"101101110",
  46772=>"111011011",
  46773=>"000000111",
  46774=>"001000000",
  46775=>"000010101",
  46776=>"001011001",
  46777=>"000110110",
  46778=>"111110001",
  46779=>"000000000",
  46780=>"001001000",
  46781=>"100111111",
  46782=>"111100101",
  46783=>"111111010",
  46784=>"000000000",
  46785=>"111111111",
  46786=>"010111010",
  46787=>"011001000",
  46788=>"000000000",
  46789=>"111110110",
  46790=>"101100010",
  46791=>"000000110",
  46792=>"000000110",
  46793=>"000000000",
  46794=>"010000000",
  46795=>"010111000",
  46796=>"001001000",
  46797=>"001011011",
  46798=>"111011001",
  46799=>"111110110",
  46800=>"111111111",
  46801=>"111000000",
  46802=>"010110111",
  46803=>"000100110",
  46804=>"000000101",
  46805=>"100110111",
  46806=>"100000000",
  46807=>"000111000",
  46808=>"001000000",
  46809=>"011111110",
  46810=>"000111111",
  46811=>"000000110",
  46812=>"111011000",
  46813=>"010000111",
  46814=>"000000000",
  46815=>"011100001",
  46816=>"000000000",
  46817=>"000000011",
  46818=>"111100000",
  46819=>"000000000",
  46820=>"000000000",
  46821=>"001000000",
  46822=>"011101101",
  46823=>"011010111",
  46824=>"000000110",
  46825=>"100111011",
  46826=>"000000000",
  46827=>"000000000",
  46828=>"111110010",
  46829=>"011000000",
  46830=>"000001010",
  46831=>"110000000",
  46832=>"111100000",
  46833=>"111011011",
  46834=>"010011110",
  46835=>"111100000",
  46836=>"111010000",
  46837=>"000111110",
  46838=>"000000000",
  46839=>"111111001",
  46840=>"010111000",
  46841=>"110111111",
  46842=>"010110000",
  46843=>"010001001",
  46844=>"111110000",
  46845=>"100010000",
  46846=>"001011011",
  46847=>"011111011",
  46848=>"110111100",
  46849=>"010101101",
  46850=>"000000101",
  46851=>"000010010",
  46852=>"000000001",
  46853=>"111110000",
  46854=>"000010010",
  46855=>"111111100",
  46856=>"000000001",
  46857=>"000000000",
  46858=>"000001000",
  46859=>"000000000",
  46860=>"010010000",
  46861=>"010111111",
  46862=>"110001001",
  46863=>"111111000",
  46864=>"001011100",
  46865=>"100111111",
  46866=>"010010010",
  46867=>"000000000",
  46868=>"000000111",
  46869=>"110101100",
  46870=>"010110110",
  46871=>"101111011",
  46872=>"011111000",
  46873=>"011011001",
  46874=>"111111111",
  46875=>"000001000",
  46876=>"000000000",
  46877=>"011000000",
  46878=>"111010000",
  46879=>"111000000",
  46880=>"000010101",
  46881=>"010010101",
  46882=>"111000011",
  46883=>"001100010",
  46884=>"111110000",
  46885=>"010110010",
  46886=>"000011010",
  46887=>"000001000",
  46888=>"111111101",
  46889=>"001110101",
  46890=>"100000110",
  46891=>"010111101",
  46892=>"011011011",
  46893=>"111110010",
  46894=>"111111001",
  46895=>"011001111",
  46896=>"000000111",
  46897=>"110001001",
  46898=>"001010000",
  46899=>"111001101",
  46900=>"000110111",
  46901=>"000000111",
  46902=>"110110001",
  46903=>"101000000",
  46904=>"000001111",
  46905=>"011100000",
  46906=>"000100100",
  46907=>"000001111",
  46908=>"100110101",
  46909=>"000111011",
  46910=>"000001110",
  46911=>"000000110",
  46912=>"011000101",
  46913=>"111111101",
  46914=>"111111011",
  46915=>"111101111",
  46916=>"000000111",
  46917=>"101000010",
  46918=>"000000000",
  46919=>"111101000",
  46920=>"111001100",
  46921=>"111111000",
  46922=>"111000001",
  46923=>"101000000",
  46924=>"101100000",
  46925=>"011111000",
  46926=>"000100000",
  46927=>"111110111",
  46928=>"000010101",
  46929=>"010000000",
  46930=>"011010000",
  46931=>"001000100",
  46932=>"010000000",
  46933=>"011000111",
  46934=>"011001001",
  46935=>"111111011",
  46936=>"110111101",
  46937=>"111001000",
  46938=>"010000011",
  46939=>"110111000",
  46940=>"000000011",
  46941=>"000001001",
  46942=>"001000100",
  46943=>"101101101",
  46944=>"000111111",
  46945=>"111100110",
  46946=>"111010000",
  46947=>"000000100",
  46948=>"100100000",
  46949=>"111100000",
  46950=>"110110000",
  46951=>"101101111",
  46952=>"000100110",
  46953=>"111111101",
  46954=>"100011011",
  46955=>"001010000",
  46956=>"011111111",
  46957=>"000101000",
  46958=>"000000111",
  46959=>"010111111",
  46960=>"010111011",
  46961=>"111111111",
  46962=>"011101100",
  46963=>"101111010",
  46964=>"000111111",
  46965=>"000000101",
  46966=>"001111111",
  46967=>"011011001",
  46968=>"111111100",
  46969=>"010100000",
  46970=>"111001000",
  46971=>"000101101",
  46972=>"011110101",
  46973=>"000100000",
  46974=>"000001111",
  46975=>"010000110",
  46976=>"101111010",
  46977=>"010111000",
  46978=>"110000000",
  46979=>"111001001",
  46980=>"111111111",
  46981=>"101001000",
  46982=>"011111111",
  46983=>"111110110",
  46984=>"001111011",
  46985=>"101101101",
  46986=>"101111111",
  46987=>"100000000",
  46988=>"000101000",
  46989=>"110001111",
  46990=>"010001111",
  46991=>"000001010",
  46992=>"110110011",
  46993=>"001101111",
  46994=>"000101111",
  46995=>"011100100",
  46996=>"010000000",
  46997=>"111010000",
  46998=>"101000100",
  46999=>"110000111",
  47000=>"000101110",
  47001=>"000111111",
  47002=>"001101111",
  47003=>"000001101",
  47004=>"000011011",
  47005=>"011000100",
  47006=>"000100111",
  47007=>"000000001",
  47008=>"000100000",
  47009=>"110000000",
  47010=>"111100000",
  47011=>"010100111",
  47012=>"010000100",
  47013=>"010011011",
  47014=>"101001000",
  47015=>"101000011",
  47016=>"111111010",
  47017=>"000110111",
  47018=>"100110111",
  47019=>"110111110",
  47020=>"101000011",
  47021=>"111111110",
  47022=>"100100100",
  47023=>"111010000",
  47024=>"100000000",
  47025=>"110001001",
  47026=>"000000100",
  47027=>"111000100",
  47028=>"110110110",
  47029=>"101100100",
  47030=>"110100000",
  47031=>"001010000",
  47032=>"001010111",
  47033=>"110010001",
  47034=>"010000000",
  47035=>"000011111",
  47036=>"101100000",
  47037=>"111111110",
  47038=>"000000001",
  47039=>"101101111",
  47040=>"000110111",
  47041=>"000000000",
  47042=>"000111111",
  47043=>"110110111",
  47044=>"011000000",
  47045=>"101001000",
  47046=>"111010000",
  47047=>"000100010",
  47048=>"111010101",
  47049=>"100001110",
  47050=>"100101100",
  47051=>"001000100",
  47052=>"000000000",
  47053=>"000001111",
  47054=>"101101001",
  47055=>"000001011",
  47056=>"100111000",
  47057=>"000100110",
  47058=>"011000000",
  47059=>"001101011",
  47060=>"110011101",
  47061=>"111100100",
  47062=>"010010000",
  47063=>"001111101",
  47064=>"101101111",
  47065=>"000000111",
  47066=>"111100000",
  47067=>"000000000",
  47068=>"111011110",
  47069=>"000011111",
  47070=>"111111010",
  47071=>"011111000",
  47072=>"100111001",
  47073=>"100010100",
  47074=>"110000000",
  47075=>"001111111",
  47076=>"000000000",
  47077=>"011101111",
  47078=>"000000000",
  47079=>"010100000",
  47080=>"101100111",
  47081=>"100111111",
  47082=>"101100001",
  47083=>"000000111",
  47084=>"101100000",
  47085=>"010111101",
  47086=>"000000000",
  47087=>"000000000",
  47088=>"000000111",
  47089=>"100000100",
  47090=>"000010000",
  47091=>"011001000",
  47092=>"110111001",
  47093=>"010111111",
  47094=>"000000000",
  47095=>"110000000",
  47096=>"000000101",
  47097=>"000111111",
  47098=>"010011000",
  47099=>"110010000",
  47100=>"101000001",
  47101=>"000000100",
  47102=>"110111000",
  47103=>"000000000",
  47104=>"110111001",
  47105=>"100101010",
  47106=>"001001111",
  47107=>"101000000",
  47108=>"100000100",
  47109=>"010001100",
  47110=>"100000001",
  47111=>"101011011",
  47112=>"100101111",
  47113=>"000011011",
  47114=>"010010100",
  47115=>"000010111",
  47116=>"111000000",
  47117=>"010111111",
  47118=>"100100100",
  47119=>"000100110",
  47120=>"000110111",
  47121=>"111111000",
  47122=>"111010000",
  47123=>"001001001",
  47124=>"001111101",
  47125=>"111101101",
  47126=>"110010000",
  47127=>"001010010",
  47128=>"100000001",
  47129=>"101111111",
  47130=>"000111111",
  47131=>"000000000",
  47132=>"000000111",
  47133=>"111111011",
  47134=>"011010000",
  47135=>"011010111",
  47136=>"011001101",
  47137=>"111011000",
  47138=>"000010110",
  47139=>"011010000",
  47140=>"000110100",
  47141=>"100000100",
  47142=>"111001000",
  47143=>"100111101",
  47144=>"111101111",
  47145=>"001010010",
  47146=>"000000110",
  47147=>"010000001",
  47148=>"011111101",
  47149=>"010010111",
  47150=>"000001000",
  47151=>"001000111",
  47152=>"111101000",
  47153=>"101100110",
  47154=>"100010000",
  47155=>"010000101",
  47156=>"111111100",
  47157=>"111101100",
  47158=>"011011001",
  47159=>"000111110",
  47160=>"011000001",
  47161=>"101100101",
  47162=>"000010000",
  47163=>"100010010",
  47164=>"000000100",
  47165=>"111111110",
  47166=>"000110100",
  47167=>"100000011",
  47168=>"101000000",
  47169=>"010100110",
  47170=>"000000010",
  47171=>"000000100",
  47172=>"111111000",
  47173=>"000000110",
  47174=>"000000000",
  47175=>"101000000",
  47176=>"001111111",
  47177=>"100000000",
  47178=>"101100111",
  47179=>"000000001",
  47180=>"000010010",
  47181=>"111111111",
  47182=>"111111001",
  47183=>"010111111",
  47184=>"111011000",
  47185=>"101011111",
  47186=>"000001010",
  47187=>"111001011",
  47188=>"110000101",
  47189=>"100010110",
  47190=>"110010011",
  47191=>"010000001",
  47192=>"000101001",
  47193=>"101000000",
  47194=>"011001100",
  47195=>"000000001",
  47196=>"111010000",
  47197=>"010001100",
  47198=>"111111010",
  47199=>"001000001",
  47200=>"000010000",
  47201=>"001100000",
  47202=>"000111000",
  47203=>"000100001",
  47204=>"110010111",
  47205=>"001011001",
  47206=>"111000110",
  47207=>"011101111",
  47208=>"000000011",
  47209=>"100000000",
  47210=>"000010011",
  47211=>"111000000",
  47212=>"110011000",
  47213=>"010010111",
  47214=>"000010000",
  47215=>"000001111",
  47216=>"011011011",
  47217=>"100010111",
  47218=>"100100100",
  47219=>"010010010",
  47220=>"000010111",
  47221=>"000000101",
  47222=>"000100011",
  47223=>"111111000",
  47224=>"011000001",
  47225=>"000000000",
  47226=>"100010010",
  47227=>"101100101",
  47228=>"110101110",
  47229=>"011110001",
  47230=>"010000001",
  47231=>"000000101",
  47232=>"101010000",
  47233=>"111000000",
  47234=>"100000101",
  47235=>"111111000",
  47236=>"111000000",
  47237=>"000001000",
  47238=>"000000001",
  47239=>"000001011",
  47240=>"011110110",
  47241=>"110100101",
  47242=>"000011011",
  47243=>"101000000",
  47244=>"000000101",
  47245=>"101001101",
  47246=>"000000101",
  47247=>"000000100",
  47248=>"100101001",
  47249=>"100000000",
  47250=>"000000101",
  47251=>"100000001",
  47252=>"000000001",
  47253=>"000000000",
  47254=>"001010000",
  47255=>"111111000",
  47256=>"110111111",
  47257=>"101000001",
  47258=>"001011111",
  47259=>"000000101",
  47260=>"011111110",
  47261=>"000010000",
  47262=>"000101111",
  47263=>"011010000",
  47264=>"000011001",
  47265=>"101011101",
  47266=>"101000100",
  47267=>"111110010",
  47268=>"011000100",
  47269=>"000110110",
  47270=>"111111000",
  47271=>"000000111",
  47272=>"110010111",
  47273=>"001101000",
  47274=>"101101101",
  47275=>"010111000",
  47276=>"110001000",
  47277=>"111110010",
  47278=>"111111100",
  47279=>"111010110",
  47280=>"111001010",
  47281=>"010001101",
  47282=>"111101111",
  47283=>"100110010",
  47284=>"111111011",
  47285=>"110001000",
  47286=>"111011011",
  47287=>"000010111",
  47288=>"000000001",
  47289=>"100100100",
  47290=>"011000001",
  47291=>"111010010",
  47292=>"100011110",
  47293=>"001111010",
  47294=>"001001101",
  47295=>"010000010",
  47296=>"100000000",
  47297=>"111000000",
  47298=>"000001000",
  47299=>"111110110",
  47300=>"011000000",
  47301=>"101000000",
  47302=>"100110111",
  47303=>"110101111",
  47304=>"100011111",
  47305=>"011000001",
  47306=>"101111111",
  47307=>"111011111",
  47308=>"000100100",
  47309=>"011101000",
  47310=>"010000000",
  47311=>"010000000",
  47312=>"001100101",
  47313=>"110110110",
  47314=>"101011111",
  47315=>"000010010",
  47316=>"100100101",
  47317=>"011110011",
  47318=>"000001101",
  47319=>"101101111",
  47320=>"111000010",
  47321=>"010000101",
  47322=>"101110101",
  47323=>"110000000",
  47324=>"011011101",
  47325=>"010010100",
  47326=>"111111111",
  47327=>"010000000",
  47328=>"000001000",
  47329=>"000000000",
  47330=>"111000110",
  47331=>"000101111",
  47332=>"110100001",
  47333=>"000111001",
  47334=>"000111111",
  47335=>"100101001",
  47336=>"000111011",
  47337=>"111110000",
  47338=>"100011001",
  47339=>"111011010",
  47340=>"111000001",
  47341=>"000000000",
  47342=>"010011110",
  47343=>"010110001",
  47344=>"101101101",
  47345=>"011000000",
  47346=>"110100011",
  47347=>"100110111",
  47348=>"001111111",
  47349=>"000000000",
  47350=>"000101000",
  47351=>"010000000",
  47352=>"000000000",
  47353=>"001111010",
  47354=>"111111011",
  47355=>"001000000",
  47356=>"111111010",
  47357=>"111101110",
  47358=>"011010001",
  47359=>"100100001",
  47360=>"100100100",
  47361=>"011001100",
  47362=>"110111001",
  47363=>"000000000",
  47364=>"110111100",
  47365=>"000000000",
  47366=>"100000000",
  47367=>"100101111",
  47368=>"111110000",
  47369=>"111111010",
  47370=>"110111011",
  47371=>"000000000",
  47372=>"100000000",
  47373=>"110100111",
  47374=>"001011110",
  47375=>"011101111",
  47376=>"000110000",
  47377=>"011111001",
  47378=>"010111010",
  47379=>"001100000",
  47380=>"110111111",
  47381=>"000110000",
  47382=>"010101100",
  47383=>"110000111",
  47384=>"111000000",
  47385=>"111000101",
  47386=>"011001000",
  47387=>"000111011",
  47388=>"011001111",
  47389=>"100111111",
  47390=>"100111000",
  47391=>"111001000",
  47392=>"010111111",
  47393=>"000000000",
  47394=>"111100100",
  47395=>"010000000",
  47396=>"110111110",
  47397=>"000011011",
  47398=>"010011010",
  47399=>"000111111",
  47400=>"111111111",
  47401=>"111011111",
  47402=>"000000000",
  47403=>"000000000",
  47404=>"000001001",
  47405=>"001100010",
  47406=>"100000101",
  47407=>"011001111",
  47408=>"000000111",
  47409=>"110110111",
  47410=>"111110111",
  47411=>"000000011",
  47412=>"000000000",
  47413=>"000000000",
  47414=>"011111011",
  47415=>"100000010",
  47416=>"100100011",
  47417=>"101101000",
  47418=>"100100101",
  47419=>"000111110",
  47420=>"010000111",
  47421=>"111111011",
  47422=>"010101101",
  47423=>"000110110",
  47424=>"000011000",
  47425=>"000011101",
  47426=>"111110111",
  47427=>"010010010",
  47428=>"010010010",
  47429=>"101001000",
  47430=>"001111101",
  47431=>"011000011",
  47432=>"000000010",
  47433=>"000111111",
  47434=>"111101001",
  47435=>"000000000",
  47436=>"010110010",
  47437=>"001011011",
  47438=>"111010111",
  47439=>"111111111",
  47440=>"000010010",
  47441=>"111111111",
  47442=>"000000000",
  47443=>"001001011",
  47444=>"000011000",
  47445=>"000000000",
  47446=>"011001011",
  47447=>"111011111",
  47448=>"111101000",
  47449=>"111111111",
  47450=>"001011000",
  47451=>"000000010",
  47452=>"100000000",
  47453=>"101001001",
  47454=>"110111011",
  47455=>"110011111",
  47456=>"010111111",
  47457=>"110000010",
  47458=>"000100100",
  47459=>"010111110",
  47460=>"100000100",
  47461=>"110111111",
  47462=>"000111110",
  47463=>"011111100",
  47464=>"000000010",
  47465=>"000111111",
  47466=>"111111111",
  47467=>"001000110",
  47468=>"111111111",
  47469=>"000011111",
  47470=>"000000101",
  47471=>"010110100",
  47472=>"011011111",
  47473=>"000000101",
  47474=>"011111010",
  47475=>"100000000",
  47476=>"111101111",
  47477=>"100100100",
  47478=>"111001111",
  47479=>"010010010",
  47480=>"101001000",
  47481=>"000000000",
  47482=>"000000000",
  47483=>"101110010",
  47484=>"001000101",
  47485=>"110101110",
  47486=>"000101111",
  47487=>"111011010",
  47488=>"100111111",
  47489=>"111000000",
  47490=>"000100000",
  47491=>"011011111",
  47492=>"000000000",
  47493=>"111111111",
  47494=>"100110110",
  47495=>"100000100",
  47496=>"100111111",
  47497=>"100110110",
  47498=>"111111111",
  47499=>"000001111",
  47500=>"110000000",
  47501=>"000000100",
  47502=>"101000000",
  47503=>"000000000",
  47504=>"001001001",
  47505=>"001010000",
  47506=>"010111011",
  47507=>"011000000",
  47508=>"111000010",
  47509=>"011001001",
  47510=>"000111011",
  47511=>"110100110",
  47512=>"110111101",
  47513=>"101000000",
  47514=>"011010011",
  47515=>"000000000",
  47516=>"000000000",
  47517=>"000010000",
  47518=>"000001000",
  47519=>"001000000",
  47520=>"000000000",
  47521=>"011110000",
  47522=>"111101111",
  47523=>"111111000",
  47524=>"100100101",
  47525=>"011001010",
  47526=>"111001100",
  47527=>"000010000",
  47528=>"101111110",
  47529=>"100010111",
  47530=>"100000100",
  47531=>"110101001",
  47532=>"111101111",
  47533=>"011111011",
  47534=>"100001011",
  47535=>"100000100",
  47536=>"000000100",
  47537=>"000001011",
  47538=>"000000001",
  47539=>"111000000",
  47540=>"111110011",
  47541=>"111000100",
  47542=>"111111111",
  47543=>"000100111",
  47544=>"000000001",
  47545=>"011011010",
  47546=>"000111111",
  47547=>"000100110",
  47548=>"101111011",
  47549=>"111111111",
  47550=>"110000010",
  47551=>"000100001",
  47552=>"101000000",
  47553=>"000000000",
  47554=>"000000111",
  47555=>"100110110",
  47556=>"000000010",
  47557=>"001000100",
  47558=>"000010101",
  47559=>"000000000",
  47560=>"100100000",
  47561=>"111000000",
  47562=>"111111011",
  47563=>"011011010",
  47564=>"001111011",
  47565=>"100100000",
  47566=>"000000000",
  47567=>"111110000",
  47568=>"011011010",
  47569=>"110110110",
  47570=>"011000000",
  47571=>"101100100",
  47572=>"000000000",
  47573=>"000101100",
  47574=>"000010011",
  47575=>"001101111",
  47576=>"000000100",
  47577=>"001010010",
  47578=>"111110101",
  47579=>"100000100",
  47580=>"100000000",
  47581=>"000001101",
  47582=>"011000000",
  47583=>"001000000",
  47584=>"000110000",
  47585=>"100000000",
  47586=>"101000000",
  47587=>"000010001",
  47588=>"000010000",
  47589=>"000000001",
  47590=>"111000000",
  47591=>"000000100",
  47592=>"000101111",
  47593=>"000000101",
  47594=>"011111110",
  47595=>"001000101",
  47596=>"111101101",
  47597=>"000000000",
  47598=>"101001000",
  47599=>"111000000",
  47600=>"111111111",
  47601=>"110001101",
  47602=>"100100111",
  47603=>"111111110",
  47604=>"011010111",
  47605=>"000111010",
  47606=>"000000010",
  47607=>"000100111",
  47608=>"000000101",
  47609=>"100001011",
  47610=>"110000000",
  47611=>"000001101",
  47612=>"000010000",
  47613=>"000000100",
  47614=>"100111010",
  47615=>"000100100",
  47616=>"011011111",
  47617=>"000000000",
  47618=>"010010010",
  47619=>"111110000",
  47620=>"101001000",
  47621=>"000010001",
  47622=>"000101111",
  47623=>"110111111",
  47624=>"111000101",
  47625=>"001101111",
  47626=>"001000000",
  47627=>"000000000",
  47628=>"110010011",
  47629=>"111111111",
  47630=>"100000001",
  47631=>"010101011",
  47632=>"000111110",
  47633=>"101101000",
  47634=>"000100000",
  47635=>"000000000",
  47636=>"000000100",
  47637=>"110111100",
  47638=>"000011000",
  47639=>"101111111",
  47640=>"000000000",
  47641=>"000000000",
  47642=>"000000000",
  47643=>"101001111",
  47644=>"101101101",
  47645=>"101111001",
  47646=>"100010011",
  47647=>"111111101",
  47648=>"101000000",
  47649=>"000100000",
  47650=>"100110010",
  47651=>"000000101",
  47652=>"001000101",
  47653=>"100111001",
  47654=>"000010000",
  47655=>"001001111",
  47656=>"101111111",
  47657=>"101010101",
  47658=>"000000001",
  47659=>"000000000",
  47660=>"000000111",
  47661=>"100111011",
  47662=>"111100100",
  47663=>"100100011",
  47664=>"111001011",
  47665=>"111000111",
  47666=>"000101100",
  47667=>"100010010",
  47668=>"000101110",
  47669=>"110010010",
  47670=>"000001000",
  47671=>"111101101",
  47672=>"101110110",
  47673=>"111111111",
  47674=>"100101101",
  47675=>"000000001",
  47676=>"101111100",
  47677=>"000111111",
  47678=>"000001011",
  47679=>"111111111",
  47680=>"111010000",
  47681=>"000000110",
  47682=>"111101101",
  47683=>"001001101",
  47684=>"000010111",
  47685=>"110000000",
  47686=>"000011010",
  47687=>"000111010",
  47688=>"111111111",
  47689=>"000000101",
  47690=>"100101101",
  47691=>"110010111",
  47692=>"111111111",
  47693=>"000010111",
  47694=>"110100111",
  47695=>"001000010",
  47696=>"000001101",
  47697=>"001111000",
  47698=>"101001010",
  47699=>"001011111",
  47700=>"000010111",
  47701=>"000000010",
  47702=>"000100110",
  47703=>"001001010",
  47704=>"100110000",
  47705=>"001010110",
  47706=>"000100111",
  47707=>"011011110",
  47708=>"001000100",
  47709=>"001000001",
  47710=>"111011010",
  47711=>"100100101",
  47712=>"000000000",
  47713=>"000111111",
  47714=>"000010000",
  47715=>"101111111",
  47716=>"110001111",
  47717=>"111001100",
  47718=>"110000001",
  47719=>"111001000",
  47720=>"011111111",
  47721=>"101000000",
  47722=>"011100000",
  47723=>"111111011",
  47724=>"000111001",
  47725=>"000000000",
  47726=>"000011001",
  47727=>"111101010",
  47728=>"001101111",
  47729=>"101000100",
  47730=>"000110010",
  47731=>"100110110",
  47732=>"111111111",
  47733=>"001001101",
  47734=>"111111000",
  47735=>"000001110",
  47736=>"000000110",
  47737=>"000000000",
  47738=>"000110111",
  47739=>"000101111",
  47740=>"100000000",
  47741=>"100100101",
  47742=>"000110110",
  47743=>"010111101",
  47744=>"000000111",
  47745=>"010010010",
  47746=>"111000000",
  47747=>"110101100",
  47748=>"010000010",
  47749=>"110111000",
  47750=>"001010110",
  47751=>"000100001",
  47752=>"000111111",
  47753=>"000001011",
  47754=>"111111111",
  47755=>"011000110",
  47756=>"011010000",
  47757=>"000011011",
  47758=>"010110010",
  47759=>"000110101",
  47760=>"001000100",
  47761=>"010110101",
  47762=>"101111101",
  47763=>"111011010",
  47764=>"111111110",
  47765=>"000000000",
  47766=>"010010010",
  47767=>"111000101",
  47768=>"000000000",
  47769=>"011000001",
  47770=>"000110000",
  47771=>"000000000",
  47772=>"001001000",
  47773=>"000001101",
  47774=>"101101011",
  47775=>"000000000",
  47776=>"100001111",
  47777=>"111111011",
  47778=>"000111111",
  47779=>"000010010",
  47780=>"000000110",
  47781=>"000001001",
  47782=>"010000100",
  47783=>"000111111",
  47784=>"000000010",
  47785=>"110010000",
  47786=>"000000000",
  47787=>"000000000",
  47788=>"000001001",
  47789=>"101101111",
  47790=>"110100001",
  47791=>"011111110",
  47792=>"111111101",
  47793=>"001101101",
  47794=>"100000111",
  47795=>"000001000",
  47796=>"111000100",
  47797=>"111111001",
  47798=>"000011001",
  47799=>"101111111",
  47800=>"100101101",
  47801=>"110100000",
  47802=>"111111100",
  47803=>"101010001",
  47804=>"111000000",
  47805=>"011000000",
  47806=>"000000010",
  47807=>"000100100",
  47808=>"111111111",
  47809=>"010000000",
  47810=>"101111111",
  47811=>"001001100",
  47812=>"000100100",
  47813=>"001000110",
  47814=>"111000011",
  47815=>"101111010",
  47816=>"000101111",
  47817=>"111111110",
  47818=>"000000000",
  47819=>"011010000",
  47820=>"011001100",
  47821=>"001100000",
  47822=>"000000000",
  47823=>"111101100",
  47824=>"111111111",
  47825=>"100000011",
  47826=>"111010000",
  47827=>"101000000",
  47828=>"010000000",
  47829=>"000100000",
  47830=>"100100111",
  47831=>"101001111",
  47832=>"000000111",
  47833=>"010001011",
  47834=>"110100010",
  47835=>"101000000",
  47836=>"001010010",
  47837=>"000001100",
  47838=>"110010011",
  47839=>"111111110",
  47840=>"000010011",
  47841=>"100011011",
  47842=>"010011111",
  47843=>"000100100",
  47844=>"011010001",
  47845=>"010110111",
  47846=>"001011110",
  47847=>"101011100",
  47848=>"000001010",
  47849=>"000000010",
  47850=>"000000100",
  47851=>"000011000",
  47852=>"111000000",
  47853=>"000001100",
  47854=>"000000001",
  47855=>"101000101",
  47856=>"111110000",
  47857=>"100000110",
  47858=>"001100110",
  47859=>"101000011",
  47860=>"110101000",
  47861=>"000100101",
  47862=>"000000000",
  47863=>"100000011",
  47864=>"010011010",
  47865=>"100101100",
  47866=>"100110100",
  47867=>"111000000",
  47868=>"101101010",
  47869=>"000100101",
  47870=>"110100001",
  47871=>"000101000",
  47872=>"011011100",
  47873=>"000000000",
  47874=>"101000000",
  47875=>"010010011",
  47876=>"000100000",
  47877=>"010011000",
  47878=>"000001000",
  47879=>"011010010",
  47880=>"011110100",
  47881=>"010011110",
  47882=>"000000111",
  47883=>"000000010",
  47884=>"011000001",
  47885=>"000010011",
  47886=>"100100001",
  47887=>"110001000",
  47888=>"000011011",
  47889=>"100000111",
  47890=>"101100101",
  47891=>"100000010",
  47892=>"011010011",
  47893=>"000100111",
  47894=>"000000000",
  47895=>"111101111",
  47896=>"100000001",
  47897=>"011000101",
  47898=>"011111111",
  47899=>"000011011",
  47900=>"111100101",
  47901=>"101000000",
  47902=>"010010000",
  47903=>"111000101",
  47904=>"111111000",
  47905=>"011100100",
  47906=>"111111101",
  47907=>"000000111",
  47908=>"001111001",
  47909=>"011110000",
  47910=>"100110110",
  47911=>"101001000",
  47912=>"011001010",
  47913=>"111111000",
  47914=>"111011011",
  47915=>"111011000",
  47916=>"001011111",
  47917=>"101101110",
  47918=>"011011100",
  47919=>"000000000",
  47920=>"010011000",
  47921=>"101101101",
  47922=>"111101110",
  47923=>"101000000",
  47924=>"000111011",
  47925=>"101001110",
  47926=>"000000000",
  47927=>"010110000",
  47928=>"010101000",
  47929=>"000000111",
  47930=>"101100111",
  47931=>"000100000",
  47932=>"000100000",
  47933=>"111000000",
  47934=>"000011011",
  47935=>"010111111",
  47936=>"010001010",
  47937=>"111011000",
  47938=>"111111000",
  47939=>"000011010",
  47940=>"111000010",
  47941=>"010100010",
  47942=>"101010011",
  47943=>"101000101",
  47944=>"000001110",
  47945=>"010011100",
  47946=>"000000011",
  47947=>"100010010",
  47948=>"111111111",
  47949=>"000111111",
  47950=>"001111110",
  47951=>"101111110",
  47952=>"100010111",
  47953=>"111101111",
  47954=>"000110100",
  47955=>"001001010",
  47956=>"100111111",
  47957=>"001000110",
  47958=>"001100100",
  47959=>"000111111",
  47960=>"001000111",
  47961=>"010110001",
  47962=>"101101101",
  47963=>"011011010",
  47964=>"001000000",
  47965=>"100001000",
  47966=>"000000111",
  47967=>"000010010",
  47968=>"000010111",
  47969=>"111000011",
  47970=>"000010111",
  47971=>"011100100",
  47972=>"000111100",
  47973=>"111001000",
  47974=>"111110000",
  47975=>"111100100",
  47976=>"111010110",
  47977=>"111101101",
  47978=>"010011111",
  47979=>"111010101",
  47980=>"110000001",
  47981=>"000111111",
  47982=>"000011011",
  47983=>"011111100",
  47984=>"000111100",
  47985=>"011011000",
  47986=>"000000000",
  47987=>"111100100",
  47988=>"010110111",
  47989=>"001000100",
  47990=>"101010010",
  47991=>"010011101",
  47992=>"000000000",
  47993=>"111101001",
  47994=>"111101101",
  47995=>"011001000",
  47996=>"100000000",
  47997=>"010110000",
  47998=>"000101011",
  47999=>"000010010",
  48000=>"000000000",
  48001=>"100100110",
  48002=>"011010000",
  48003=>"111110111",
  48004=>"011101000",
  48005=>"101000000",
  48006=>"110111000",
  48007=>"000110110",
  48008=>"010111001",
  48009=>"100100111",
  48010=>"100011011",
  48011=>"000000100",
  48012=>"101001011",
  48013=>"001111010",
  48014=>"010001011",
  48015=>"000000001",
  48016=>"111101101",
  48017=>"111111000",
  48018=>"100100110",
  48019=>"000010100",
  48020=>"000010010",
  48021=>"000000010",
  48022=>"110111001",
  48023=>"001101000",
  48024=>"000010010",
  48025=>"101001111",
  48026=>"100100011",
  48027=>"100100111",
  48028=>"000010000",
  48029=>"001010000",
  48030=>"010000111",
  48031=>"100101100",
  48032=>"100100110",
  48033=>"001000000",
  48034=>"010000011",
  48035=>"100000001",
  48036=>"111100101",
  48037=>"100011011",
  48038=>"010101000",
  48039=>"000111111",
  48040=>"100000000",
  48041=>"001101011",
  48042=>"010101111",
  48043=>"000000000",
  48044=>"011110100",
  48045=>"010011110",
  48046=>"011110111",
  48047=>"111110010",
  48048=>"010111111",
  48049=>"100000001",
  48050=>"101111000",
  48051=>"101101000",
  48052=>"001111100",
  48053=>"101011100",
  48054=>"011010000",
  48055=>"111011000",
  48056=>"000001000",
  48057=>"000110101",
  48058=>"011011100",
  48059=>"000101100",
  48060=>"011000001",
  48061=>"111110111",
  48062=>"001111000",
  48063=>"001101111",
  48064=>"100010110",
  48065=>"010011111",
  48066=>"111001011",
  48067=>"000011101",
  48068=>"011101101",
  48069=>"000100001",
  48070=>"010000000",
  48071=>"111011110",
  48072=>"111011111",
  48073=>"000110000",
  48074=>"011000000",
  48075=>"011011010",
  48076=>"100010010",
  48077=>"000000000",
  48078=>"100011011",
  48079=>"011001000",
  48080=>"100100111",
  48081=>"011111000",
  48082=>"010000100",
  48083=>"111101110",
  48084=>"000001011",
  48085=>"000110110",
  48086=>"100001101",
  48087=>"010001000",
  48088=>"110101111",
  48089=>"000000111",
  48090=>"011011111",
  48091=>"101000001",
  48092=>"000100000",
  48093=>"111011111",
  48094=>"000000101",
  48095=>"011000000",
  48096=>"000011111",
  48097=>"111001101",
  48098=>"111101100",
  48099=>"000011110",
  48100=>"000000000",
  48101=>"110100100",
  48102=>"111011010",
  48103=>"000011111",
  48104=>"000011010",
  48105=>"000010000",
  48106=>"100000111",
  48107=>"011111111",
  48108=>"100000110",
  48109=>"010110110",
  48110=>"000000000",
  48111=>"000000000",
  48112=>"111000111",
  48113=>"000101111",
  48114=>"011011000",
  48115=>"001101101",
  48116=>"010110000",
  48117=>"101000111",
  48118=>"000000001",
  48119=>"011111000",
  48120=>"100000010",
  48121=>"101100111",
  48122=>"010000111",
  48123=>"000000111",
  48124=>"100011011",
  48125=>"111100101",
  48126=>"011110110",
  48127=>"101011000",
  48128=>"000100000",
  48129=>"000001010",
  48130=>"100000000",
  48131=>"000001000",
  48132=>"111111011",
  48133=>"000000001",
  48134=>"000000111",
  48135=>"000000001",
  48136=>"100010110",
  48137=>"111101111",
  48138=>"111111111",
  48139=>"110010000",
  48140=>"110010111",
  48141=>"111101111",
  48142=>"000101000",
  48143=>"110111111",
  48144=>"111110011",
  48145=>"000000100",
  48146=>"011010010",
  48147=>"000000110",
  48148=>"100001000",
  48149=>"111010000",
  48150=>"111111111",
  48151=>"110011111",
  48152=>"001001001",
  48153=>"101111001",
  48154=>"000010001",
  48155=>"100100101",
  48156=>"000001000",
  48157=>"000000001",
  48158=>"010011110",
  48159=>"000000001",
  48160=>"000001000",
  48161=>"000000001",
  48162=>"001000011",
  48163=>"111001001",
  48164=>"100000101",
  48165=>"100110000",
  48166=>"111011010",
  48167=>"111111111",
  48168=>"111000111",
  48169=>"001000100",
  48170=>"000000110",
  48171=>"110110011",
  48172=>"011111111",
  48173=>"011000000",
  48174=>"100100100",
  48175=>"100001001",
  48176=>"101100000",
  48177=>"000000000",
  48178=>"000000011",
  48179=>"000000011",
  48180=>"111111000",
  48181=>"000000000",
  48182=>"110100100",
  48183=>"000000000",
  48184=>"000000000",
  48185=>"001001001",
  48186=>"010010010",
  48187=>"110111111",
  48188=>"000000000",
  48189=>"111111111",
  48190=>"000101111",
  48191=>"110110111",
  48192=>"100110111",
  48193=>"111110010",
  48194=>"000011111",
  48195=>"110111011",
  48196=>"100101111",
  48197=>"011000100",
  48198=>"100110111",
  48199=>"111111111",
  48200=>"000000000",
  48201=>"111111111",
  48202=>"111000101",
  48203=>"010111111",
  48204=>"001000000",
  48205=>"011011011",
  48206=>"111111111",
  48207=>"111111111",
  48208=>"100000101",
  48209=>"111111011",
  48210=>"111101111",
  48211=>"000000000",
  48212=>"000111111",
  48213=>"000000010",
  48214=>"010100110",
  48215=>"101001111",
  48216=>"000001001",
  48217=>"111111111",
  48218=>"000100100",
  48219=>"111110111",
  48220=>"000000001",
  48221=>"000000000",
  48222=>"010000010",
  48223=>"111111110",
  48224=>"111001111",
  48225=>"110111111",
  48226=>"000000001",
  48227=>"001111011",
  48228=>"000001101",
  48229=>"011111000",
  48230=>"000110111",
  48231=>"010000000",
  48232=>"001111110",
  48233=>"101111010",
  48234=>"000000110",
  48235=>"000000100",
  48236=>"101000111",
  48237=>"101101001",
  48238=>"110111110",
  48239=>"100101001",
  48240=>"110110110",
  48241=>"000000100",
  48242=>"001001100",
  48243=>"110110111",
  48244=>"011011111",
  48245=>"000000111",
  48246=>"000000000",
  48247=>"010011111",
  48248=>"111111111",
  48249=>"011111111",
  48250=>"000000110",
  48251=>"100000100",
  48252=>"010110110",
  48253=>"000000000",
  48254=>"111011111",
  48255=>"101111101",
  48256=>"000101011",
  48257=>"111111111",
  48258=>"000000000",
  48259=>"001100111",
  48260=>"000000000",
  48261=>"000001111",
  48262=>"011011010",
  48263=>"010010000",
  48264=>"101001011",
  48265=>"101111111",
  48266=>"111111010",
  48267=>"000000110",
  48268=>"000111011",
  48269=>"111110110",
  48270=>"000110110",
  48271=>"000000101",
  48272=>"001001111",
  48273=>"000000000",
  48274=>"000000000",
  48275=>"011010111",
  48276=>"000110111",
  48277=>"000000110",
  48278=>"111110110",
  48279=>"000000011",
  48280=>"111100010",
  48281=>"111111111",
  48282=>"011110110",
  48283=>"110110110",
  48284=>"000111111",
  48285=>"111110000",
  48286=>"000000000",
  48287=>"000101101",
  48288=>"110110011",
  48289=>"111111111",
  48290=>"101000101",
  48291=>"011111011",
  48292=>"111000000",
  48293=>"110111111",
  48294=>"111111001",
  48295=>"001001001",
  48296=>"000001011",
  48297=>"000000000",
  48298=>"001000000",
  48299=>"101101111",
  48300=>"111111111",
  48301=>"000000000",
  48302=>"101101101",
  48303=>"111111110",
  48304=>"111111111",
  48305=>"000000100",
  48306=>"000110000",
  48307=>"011011100",
  48308=>"111001111",
  48309=>"001111010",
  48310=>"000011111",
  48311=>"000010000",
  48312=>"001001000",
  48313=>"000111110",
  48314=>"001110100",
  48315=>"100111110",
  48316=>"100000001",
  48317=>"111011100",
  48318=>"111110110",
  48319=>"001001110",
  48320=>"110110010",
  48321=>"111110000",
  48322=>"110101000",
  48323=>"010010110",
  48324=>"000000000",
  48325=>"100000000",
  48326=>"100000111",
  48327=>"010111110",
  48328=>"001000000",
  48329=>"111111110",
  48330=>"010011111",
  48331=>"110111000",
  48332=>"100100011",
  48333=>"000010010",
  48334=>"000000001",
  48335=>"000111001",
  48336=>"111111000",
  48337=>"110110110",
  48338=>"101000000",
  48339=>"000000000",
  48340=>"011011001",
  48341=>"001001000",
  48342=>"000000001",
  48343=>"111100000",
  48344=>"111001001",
  48345=>"111100000",
  48346=>"001011011",
  48347=>"111111110",
  48348=>"011111110",
  48349=>"001111111",
  48350=>"110111111",
  48351=>"000000000",
  48352=>"111110000",
  48353=>"010001111",
  48354=>"001000000",
  48355=>"111111111",
  48356=>"101001001",
  48357=>"111000111",
  48358=>"100000101",
  48359=>"111111111",
  48360=>"000000000",
  48361=>"000101111",
  48362=>"111111111",
  48363=>"111111111",
  48364=>"111101001",
  48365=>"000011000",
  48366=>"000000001",
  48367=>"000000000",
  48368=>"000000001",
  48369=>"001001000",
  48370=>"101110101",
  48371=>"110000000",
  48372=>"001111111",
  48373=>"110111001",
  48374=>"000001111",
  48375=>"110000000",
  48376=>"010000000",
  48377=>"000000000",
  48378=>"111111111",
  48379=>"000101000",
  48380=>"000010000",
  48381=>"000100111",
  48382=>"100100100",
  48383=>"000111111",
  48384=>"001001001",
  48385=>"000100111",
  48386=>"101100101",
  48387=>"011010011",
  48388=>"110100111",
  48389=>"010010010",
  48390=>"111100100",
  48391=>"000010011",
  48392=>"000100101",
  48393=>"000000001",
  48394=>"101100100",
  48395=>"111100000",
  48396=>"000011010",
  48397=>"000010000",
  48398=>"100111011",
  48399=>"001100111",
  48400=>"110000101",
  48401=>"000000111",
  48402=>"101000111",
  48403=>"111100100",
  48404=>"000000101",
  48405=>"000000010",
  48406=>"111111111",
  48407=>"111101100",
  48408=>"111100100",
  48409=>"110001101",
  48410=>"000000010",
  48411=>"111101111",
  48412=>"000100101",
  48413=>"100000000",
  48414=>"111111011",
  48415=>"101000000",
  48416=>"000000000",
  48417=>"010011011",
  48418=>"101101111",
  48419=>"000010010",
  48420=>"001011010",
  48421=>"010110100",
  48422=>"000010010",
  48423=>"000000111",
  48424=>"101010111",
  48425=>"001010000",
  48426=>"101000100",
  48427=>"110000000",
  48428=>"111001001",
  48429=>"111100111",
  48430=>"011000100",
  48431=>"111111110",
  48432=>"011011111",
  48433=>"011110101",
  48434=>"000111111",
  48435=>"111000000",
  48436=>"111000000",
  48437=>"000100000",
  48438=>"000010011",
  48439=>"010111100",
  48440=>"010010000",
  48441=>"000001001",
  48442=>"011100111",
  48443=>"100100000",
  48444=>"000111110",
  48445=>"110111010",
  48446=>"000000000",
  48447=>"100110110",
  48448=>"000000110",
  48449=>"101011001",
  48450=>"011111111",
  48451=>"011011000",
  48452=>"000000010",
  48453=>"011000100",
  48454=>"000000000",
  48455=>"000010000",
  48456=>"000001010",
  48457=>"000011111",
  48458=>"101000000",
  48459=>"111100100",
  48460=>"111011000",
  48461=>"100110011",
  48462=>"011011010",
  48463=>"101000111",
  48464=>"101110000",
  48465=>"111010000",
  48466=>"111101111",
  48467=>"010000000",
  48468=>"111101100",
  48469=>"010111111",
  48470=>"010011001",
  48471=>"111000000",
  48472=>"111000100",
  48473=>"100110100",
  48474=>"100010010",
  48475=>"000011001",
  48476=>"000011011",
  48477=>"111001001",
  48478=>"100011111",
  48479=>"000000010",
  48480=>"000011111",
  48481=>"000000111",
  48482=>"111000000",
  48483=>"111101101",
  48484=>"000100000",
  48485=>"111110010",
  48486=>"111100000",
  48487=>"001011000",
  48488=>"111011111",
  48489=>"010111000",
  48490=>"000010010",
  48491=>"001000000",
  48492=>"100100000",
  48493=>"011000101",
  48494=>"010000000",
  48495=>"111000010",
  48496=>"000000100",
  48497=>"010011000",
  48498=>"000010111",
  48499=>"111011011",
  48500=>"000111111",
  48501=>"100100100",
  48502=>"010011010",
  48503=>"000111010",
  48504=>"101111000",
  48505=>"011011011",
  48506=>"111000000",
  48507=>"000101100",
  48508=>"100110100",
  48509=>"010100000",
  48510=>"111100111",
  48511=>"100000000",
  48512=>"111011010",
  48513=>"000000000",
  48514=>"000111011",
  48515=>"000000011",
  48516=>"101001000",
  48517=>"111000000",
  48518=>"100111000",
  48519=>"110101100",
  48520=>"000000100",
  48521=>"101100000",
  48522=>"111100110",
  48523=>"111011000",
  48524=>"000000101",
  48525=>"101101111",
  48526=>"110111110",
  48527=>"001000000",
  48528=>"100100000",
  48529=>"100100101",
  48530=>"111100111",
  48531=>"111011100",
  48532=>"100110000",
  48533=>"110110000",
  48534=>"011111011",
  48535=>"000011011",
  48536=>"010100100",
  48537=>"011100111",
  48538=>"000111011",
  48539=>"100100110",
  48540=>"001111000",
  48541=>"110111100",
  48542=>"011010000",
  48543=>"111000000",
  48544=>"000100111",
  48545=>"110111010",
  48546=>"000011001",
  48547=>"011100011",
  48548=>"000000000",
  48549=>"000011100",
  48550=>"101111010",
  48551=>"000011011",
  48552=>"100111111",
  48553=>"000010111",
  48554=>"111000000",
  48555=>"110100100",
  48556=>"111010000",
  48557=>"000011011",
  48558=>"111110110",
  48559=>"111111011",
  48560=>"000100100",
  48561=>"011001001",
  48562=>"111111100",
  48563=>"000111100",
  48564=>"000011011",
  48565=>"111111111",
  48566=>"000100110",
  48567=>"000011001",
  48568=>"101111011",
  48569=>"001111000",
  48570=>"111010001",
  48571=>"111000010",
  48572=>"011000001",
  48573=>"000111111",
  48574=>"000011111",
  48575=>"111100011",
  48576=>"111000000",
  48577=>"001000000",
  48578=>"001101111",
  48579=>"011011010",
  48580=>"110101101",
  48581=>"001011101",
  48582=>"111110100",
  48583=>"111001101",
  48584=>"000000100",
  48585=>"000011010",
  48586=>"010111011",
  48587=>"000100111",
  48588=>"100100000",
  48589=>"000001111",
  48590=>"101001000",
  48591=>"001001000",
  48592=>"000000111",
  48593=>"000110110",
  48594=>"111000000",
  48595=>"000111011",
  48596=>"111100110",
  48597=>"110100110",
  48598=>"100000000",
  48599=>"000001111",
  48600=>"111000000",
  48601=>"000100000",
  48602=>"001111100",
  48603=>"111000000",
  48604=>"110011111",
  48605=>"100101111",
  48606=>"000100000",
  48607=>"111111000",
  48608=>"000111111",
  48609=>"011000010",
  48610=>"111000000",
  48611=>"000000110",
  48612=>"000100000",
  48613=>"111000100",
  48614=>"110000101",
  48615=>"000001011",
  48616=>"010011111",
  48617=>"001000001",
  48618=>"100100000",
  48619=>"111000100",
  48620=>"000111111",
  48621=>"000000000",
  48622=>"000100000",
  48623=>"000100100",
  48624=>"111000000",
  48625=>"000111101",
  48626=>"100011000",
  48627=>"000011110",
  48628=>"010110011",
  48629=>"111111111",
  48630=>"000000110",
  48631=>"000101011",
  48632=>"110000000",
  48633=>"101001111",
  48634=>"010100010",
  48635=>"101001001",
  48636=>"000111000",
  48637=>"011100100",
  48638=>"001001001",
  48639=>"101100000",
  48640=>"110101000",
  48641=>"100010101",
  48642=>"101000111",
  48643=>"000000010",
  48644=>"111101101",
  48645=>"101100111",
  48646=>"000111000",
  48647=>"111111010",
  48648=>"001000000",
  48649=>"111000100",
  48650=>"001000101",
  48651=>"011000110",
  48652=>"111000101",
  48653=>"000101101",
  48654=>"100100100",
  48655=>"111111011",
  48656=>"000010101",
  48657=>"000000000",
  48658=>"011001010",
  48659=>"111111000",
  48660=>"010011011",
  48661=>"000000000",
  48662=>"110111100",
  48663=>"111011101",
  48664=>"110000111",
  48665=>"000111000",
  48666=>"111101111",
  48667=>"000000111",
  48668=>"011000010",
  48669=>"000000000",
  48670=>"000000111",
  48671=>"111000000",
  48672=>"000111001",
  48673=>"111000111",
  48674=>"000100101",
  48675=>"001100111",
  48676=>"110011001",
  48677=>"000001111",
  48678=>"000010000",
  48679=>"111111110",
  48680=>"001001000",
  48681=>"011110101",
  48682=>"111111011",
  48683=>"010011000",
  48684=>"111010011",
  48685=>"111000000",
  48686=>"101110100",
  48687=>"100000011",
  48688=>"110000111",
  48689=>"111111101",
  48690=>"101000000",
  48691=>"000000001",
  48692=>"001000111",
  48693=>"000000000",
  48694=>"100111011",
  48695=>"110000110",
  48696=>"111111010",
  48697=>"010000111",
  48698=>"111010101",
  48699=>"111000111",
  48700=>"000000000",
  48701=>"111010001",
  48702=>"111000000",
  48703=>"111111001",
  48704=>"010000000",
  48705=>"111000001",
  48706=>"110111000",
  48707=>"111000110",
  48708=>"010000000",
  48709=>"000001000",
  48710=>"000111000",
  48711=>"100000000",
  48712=>"110000000",
  48713=>"111000111",
  48714=>"110110000",
  48715=>"101010100",
  48716=>"111000111",
  48717=>"001011100",
  48718=>"111111011",
  48719=>"000000111",
  48720=>"000000010",
  48721=>"111011101",
  48722=>"101010000",
  48723=>"001001010",
  48724=>"101000110",
  48725=>"101001100",
  48726=>"111110001",
  48727=>"110000101",
  48728=>"111010010",
  48729=>"111111000",
  48730=>"111110011",
  48731=>"011111100",
  48732=>"000111000",
  48733=>"010000010",
  48734=>"010111000",
  48735=>"110000111",
  48736=>"001001111",
  48737=>"000111110",
  48738=>"111000111",
  48739=>"110111111",
  48740=>"011000001",
  48741=>"000010100",
  48742=>"111001111",
  48743=>"000011001",
  48744=>"010000111",
  48745=>"111010111",
  48746=>"111111000",
  48747=>"000000000",
  48748=>"111101101",
  48749=>"000011000",
  48750=>"010111100",
  48751=>"010011101",
  48752=>"001000010",
  48753=>"101000100",
  48754=>"001111100",
  48755=>"110110000",
  48756=>"111011000",
  48757=>"000001011",
  48758=>"100010001",
  48759=>"110001000",
  48760=>"000111111",
  48761=>"000111110",
  48762=>"000000000",
  48763=>"111000000",
  48764=>"010000011",
  48765=>"001001010",
  48766=>"011111010",
  48767=>"111000111",
  48768=>"000100000",
  48769=>"111000000",
  48770=>"000000000",
  48771=>"000111110",
  48772=>"000100000",
  48773=>"001000000",
  48774=>"100101111",
  48775=>"110000100",
  48776=>"000000000",
  48777=>"111000100",
  48778=>"010111000",
  48779=>"100000000",
  48780=>"000111000",
  48781=>"100111000",
  48782=>"101000001",
  48783=>"100000000",
  48784=>"010000111",
  48785=>"010000010",
  48786=>"001111111",
  48787=>"010111010",
  48788=>"111100000",
  48789=>"100110101",
  48790=>"000000000",
  48791=>"110010000",
  48792=>"011101111",
  48793=>"111111000",
  48794=>"000000111",
  48795=>"000000001",
  48796=>"111111111",
  48797=>"000111110",
  48798=>"000111110",
  48799=>"111000111",
  48800=>"110000110",
  48801=>"011010110",
  48802=>"110111111",
  48803=>"100000000",
  48804=>"000111101",
  48805=>"000000011",
  48806=>"100000000",
  48807=>"111111111",
  48808=>"000000101",
  48809=>"111011111",
  48810=>"111000111",
  48811=>"110010111",
  48812=>"101111000",
  48813=>"010111010",
  48814=>"100000000",
  48815=>"000111011",
  48816=>"100100000",
  48817=>"011000001",
  48818=>"111111111",
  48819=>"010001011",
  48820=>"010000100",
  48821=>"000000110",
  48822=>"001000100",
  48823=>"000000000",
  48824=>"001000111",
  48825=>"111001011",
  48826=>"111111000",
  48827=>"010000111",
  48828=>"000111000",
  48829=>"111111111",
  48830=>"001111111",
  48831=>"000100000",
  48832=>"110010000",
  48833=>"010000110",
  48834=>"000100000",
  48835=>"011101000",
  48836=>"111000000",
  48837=>"001000000",
  48838=>"000110100",
  48839=>"111111111",
  48840=>"111111000",
  48841=>"110000111",
  48842=>"100111000",
  48843=>"000000000",
  48844=>"000010000",
  48845=>"111100100",
  48846=>"000000111",
  48847=>"000001111",
  48848=>"111011111",
  48849=>"010011111",
  48850=>"100101001",
  48851=>"111000000",
  48852=>"010010000",
  48853=>"000000110",
  48854=>"111000111",
  48855=>"011011111",
  48856=>"000000000",
  48857=>"111111100",
  48858=>"010111011",
  48859=>"010010110",
  48860=>"001110111",
  48861=>"100010111",
  48862=>"000000001",
  48863=>"101101100",
  48864=>"111110111",
  48865=>"110000111",
  48866=>"000000000",
  48867=>"001010000",
  48868=>"001101001",
  48869=>"010000111",
  48870=>"000011111",
  48871=>"110001110",
  48872=>"000100000",
  48873=>"111111110",
  48874=>"111000011",
  48875=>"000000111",
  48876=>"000000111",
  48877=>"111111111",
  48878=>"011011000",
  48879=>"111101100",
  48880=>"111111110",
  48881=>"110000000",
  48882=>"110110000",
  48883=>"010111111",
  48884=>"001111000",
  48885=>"110000110",
  48886=>"011000111",
  48887=>"101000001",
  48888=>"110110100",
  48889=>"111111000",
  48890=>"011000000",
  48891=>"000001000",
  48892=>"111111111",
  48893=>"000111000",
  48894=>"111101111",
  48895=>"000010011",
  48896=>"110110110",
  48897=>"111100000",
  48898=>"000000000",
  48899=>"111001000",
  48900=>"110110110",
  48901=>"000000100",
  48902=>"101111111",
  48903=>"100100101",
  48904=>"000000100",
  48905=>"010111111",
  48906=>"100010011",
  48907=>"000000000",
  48908=>"000000000",
  48909=>"010000111",
  48910=>"011110000",
  48911=>"010001000",
  48912=>"000000000",
  48913=>"100000101",
  48914=>"111100000",
  48915=>"000110011",
  48916=>"011000000",
  48917=>"110111111",
  48918=>"111011010",
  48919=>"100100110",
  48920=>"100000000",
  48921=>"111111111",
  48922=>"100100111",
  48923=>"011011100",
  48924=>"010100000",
  48925=>"011111100",
  48926=>"111001111",
  48927=>"000000000",
  48928=>"010111000",
  48929=>"100000000",
  48930=>"000000000",
  48931=>"100000110",
  48932=>"000000111",
  48933=>"111100000",
  48934=>"000000101",
  48935=>"000000000",
  48936=>"110111111",
  48937=>"100001001",
  48938=>"101111001",
  48939=>"100000000",
  48940=>"100100110",
  48941=>"000000000",
  48942=>"000111111",
  48943=>"000100110",
  48944=>"000000000",
  48945=>"000110111",
  48946=>"000110000",
  48947=>"110111111",
  48948=>"111001101",
  48949=>"111011101",
  48950=>"100000001",
  48951=>"011011100",
  48952=>"111100000",
  48953=>"101000000",
  48954=>"000000000",
  48955=>"111100100",
  48956=>"110111000",
  48957=>"111111100",
  48958=>"000000100",
  48959=>"010011101",
  48960=>"001001101",
  48961=>"101111111",
  48962=>"100101110",
  48963=>"100000100",
  48964=>"000010000",
  48965=>"101001000",
  48966=>"000111010",
  48967=>"000000111",
  48968=>"100100100",
  48969=>"001000011",
  48970=>"101100111",
  48971=>"101100110",
  48972=>"000100000",
  48973=>"000000000",
  48974=>"001001101",
  48975=>"000000011",
  48976=>"100000000",
  48977=>"111110111",
  48978=>"100110000",
  48979=>"001000100",
  48980=>"001000001",
  48981=>"010111101",
  48982=>"011011110",
  48983=>"000000100",
  48984=>"100000000",
  48985=>"100110111",
  48986=>"001011101",
  48987=>"100110011",
  48988=>"000100100",
  48989=>"000001000",
  48990=>"011111000",
  48991=>"001001001",
  48992=>"101100111",
  48993=>"001111010",
  48994=>"000000101",
  48995=>"000100001",
  48996=>"111111010",
  48997=>"111110111",
  48998=>"101111111",
  48999=>"010110111",
  49000=>"010011010",
  49001=>"000010011",
  49002=>"010011011",
  49003=>"011110100",
  49004=>"001000000",
  49005=>"011111010",
  49006=>"111100101",
  49007=>"100000010",
  49008=>"110110110",
  49009=>"111101101",
  49010=>"001100100",
  49011=>"000000000",
  49012=>"011111111",
  49013=>"100000111",
  49014=>"000000000",
  49015=>"111111111",
  49016=>"011011000",
  49017=>"111111000",
  49018=>"011111011",
  49019=>"011101110",
  49020=>"110110111",
  49021=>"000000000",
  49022=>"000110111",
  49023=>"000001111",
  49024=>"000101101",
  49025=>"111100111",
  49026=>"011010011",
  49027=>"011111000",
  49028=>"011111001",
  49029=>"010111000",
  49030=>"000011100",
  49031=>"101100100",
  49032=>"011011001",
  49033=>"001000000",
  49034=>"011011011",
  49035=>"000100000",
  49036=>"111111000",
  49037=>"000000000",
  49038=>"011011100",
  49039=>"001000000",
  49040=>"111111111",
  49041=>"111101000",
  49042=>"000000000",
  49043=>"101100101",
  49044=>"110010100",
  49045=>"000000101",
  49046=>"111011000",
  49047=>"000011110",
  49048=>"011010010",
  49049=>"010000110",
  49050=>"111111011",
  49051=>"000000011",
  49052=>"001000111",
  49053=>"011011000",
  49054=>"100100111",
  49055=>"100100111",
  49056=>"100100110",
  49057=>"011011000",
  49058=>"111101101",
  49059=>"001111000",
  49060=>"000101111",
  49061=>"000000111",
  49062=>"100010001",
  49063=>"000000100",
  49064=>"001111111",
  49065=>"100010000",
  49066=>"001100001",
  49067=>"000100000",
  49068=>"110100100",
  49069=>"000000000",
  49070=>"010001001",
  49071=>"111111010",
  49072=>"000101001",
  49073=>"000100110",
  49074=>"001101001",
  49075=>"100000001",
  49076=>"001011111",
  49077=>"100100000",
  49078=>"100100001",
  49079=>"011111101",
  49080=>"001001100",
  49081=>"111010101",
  49082=>"011001010",
  49083=>"111100100",
  49084=>"011111001",
  49085=>"010011010",
  49086=>"000100100",
  49087=>"100000000",
  49088=>"100000100",
  49089=>"000100111",
  49090=>"000111100",
  49091=>"001101111",
  49092=>"011110000",
  49093=>"010110000",
  49094=>"111011100",
  49095=>"111111000",
  49096=>"010100000",
  49097=>"100000111",
  49098=>"001101111",
  49099=>"111111111",
  49100=>"000100100",
  49101=>"011011010",
  49102=>"000001111",
  49103=>"111111100",
  49104=>"101100111",
  49105=>"010110010",
  49106=>"100001111",
  49107=>"011001000",
  49108=>"100100111",
  49109=>"100001001",
  49110=>"100000111",
  49111=>"111011110",
  49112=>"100000101",
  49113=>"001111010",
  49114=>"001001011",
  49115=>"000010111",
  49116=>"101000001",
  49117=>"110010011",
  49118=>"000100000",
  49119=>"111011010",
  49120=>"100000111",
  49121=>"101100100",
  49122=>"000000011",
  49123=>"001111011",
  49124=>"101000111",
  49125=>"000000111",
  49126=>"000100000",
  49127=>"010110100",
  49128=>"001100100",
  49129=>"001000000",
  49130=>"100100100",
  49131=>"101100100",
  49132=>"000000101",
  49133=>"000010111",
  49134=>"101100110",
  49135=>"000100111",
  49136=>"000000000",
  49137=>"000011110",
  49138=>"100100111",
  49139=>"001111110",
  49140=>"011011101",
  49141=>"101111101",
  49142=>"001000010",
  49143=>"001001011",
  49144=>"100000111",
  49145=>"001011011",
  49146=>"000000000",
  49147=>"001111011",
  49148=>"111111000",
  49149=>"111111110",
  49150=>"000000100",
  49151=>"100100111",
  49152=>"010000100",
  49153=>"001110110",
  49154=>"001001111",
  49155=>"111000001",
  49156=>"000000110",
  49157=>"001000111",
  49158=>"000000000",
  49159=>"000000110",
  49160=>"100101110",
  49161=>"000000000",
  49162=>"101000110",
  49163=>"001000000",
  49164=>"011001101",
  49165=>"001001000",
  49166=>"000110011",
  49167=>"100010001",
  49168=>"110110111",
  49169=>"000011111",
  49170=>"000000110",
  49171=>"001110000",
  49172=>"011001001",
  49173=>"001000000",
  49174=>"100000000",
  49175=>"010111111",
  49176=>"000000111",
  49177=>"110010000",
  49178=>"110110000",
  49179=>"001000000",
  49180=>"001000101",
  49181=>"000000000",
  49182=>"111000000",
  49183=>"110110000",
  49184=>"001111111",
  49185=>"101110100",
  49186=>"100101100",
  49187=>"110110110",
  49188=>"000000011",
  49189=>"011111011",
  49190=>"001000111",
  49191=>"111111000",
  49192=>"000001111",
  49193=>"111001010",
  49194=>"000100000",
  49195=>"110111000",
  49196=>"110111011",
  49197=>"000000111",
  49198=>"000101010",
  49199=>"001000110",
  49200=>"000000001",
  49201=>"000000110",
  49202=>"011111110",
  49203=>"000001111",
  49204=>"110000001",
  49205=>"000001001",
  49206=>"111111011",
  49207=>"001000110",
  49208=>"110000000",
  49209=>"001000000",
  49210=>"001000000",
  49211=>"010100111",
  49212=>"110011010",
  49213=>"110111010",
  49214=>"000000001",
  49215=>"010111001",
  49216=>"000110111",
  49217=>"001111000",
  49218=>"110111011",
  49219=>"001110110",
  49220=>"111010010",
  49221=>"001000001",
  49222=>"000000111",
  49223=>"110000001",
  49224=>"011111000",
  49225=>"110110111",
  49226=>"001000110",
  49227=>"111110100",
  49228=>"111000001",
  49229=>"000100010",
  49230=>"100010011",
  49231=>"110110000",
  49232=>"110000010",
  49233=>"010010000",
  49234=>"111111011",
  49235=>"011000000",
  49236=>"001001101",
  49237=>"010010110",
  49238=>"111010110",
  49239=>"110110000",
  49240=>"111000101",
  49241=>"110010111",
  49242=>"101101111",
  49243=>"111110010",
  49244=>"010110000",
  49245=>"001001010",
  49246=>"101101111",
  49247=>"010110111",
  49248=>"111000110",
  49249=>"110110000",
  49250=>"001001111",
  49251=>"011001111",
  49252=>"100000000",
  49253=>"111011011",
  49254=>"110110010",
  49255=>"010111000",
  49256=>"000010111",
  49257=>"000000110",
  49258=>"000100110",
  49259=>"111110011",
  49260=>"000000000",
  49261=>"000001111",
  49262=>"010010000",
  49263=>"000001110",
  49264=>"110111110",
  49265=>"110110110",
  49266=>"111110100",
  49267=>"000000111",
  49268=>"111111110",
  49269=>"000000010",
  49270=>"000010010",
  49271=>"111001011",
  49272=>"000001000",
  49273=>"101110111",
  49274=>"001110111",
  49275=>"100001000",
  49276=>"100110010",
  49277=>"100000001",
  49278=>"010110001",
  49279=>"110010100",
  49280=>"000000000",
  49281=>"000000000",
  49282=>"101000110",
  49283=>"001101000",
  49284=>"001000001",
  49285=>"110001001",
  49286=>"110110000",
  49287=>"010100100",
  49288=>"101101111",
  49289=>"110000010",
  49290=>"100101110",
  49291=>"000000111",
  49292=>"000010000",
  49293=>"001001111",
  49294=>"011001111",
  49295=>"000000110",
  49296=>"100000100",
  49297=>"111111010",
  49298=>"111110000",
  49299=>"110000110",
  49300=>"000110101",
  49301=>"001001011",
  49302=>"100100110",
  49303=>"000001000",
  49304=>"110111001",
  49305=>"110110000",
  49306=>"001001111",
  49307=>"000000000",
  49308=>"001000001",
  49309=>"001001101",
  49310=>"110000000",
  49311=>"000010110",
  49312=>"111001011",
  49313=>"001001011",
  49314=>"111110000",
  49315=>"110100111",
  49316=>"001000000",
  49317=>"110000010",
  49318=>"001010000",
  49319=>"110111110",
  49320=>"000000101",
  49321=>"001100110",
  49322=>"000000000",
  49323=>"001001011",
  49324=>"101110110",
  49325=>"111001001",
  49326=>"100010000",
  49327=>"111111111",
  49328=>"100111110",
  49329=>"011001001",
  49330=>"011001111",
  49331=>"000100000",
  49332=>"111111110",
  49333=>"101111111",
  49334=>"111111111",
  49335=>"000101001",
  49336=>"111110100",
  49337=>"110110010",
  49338=>"010111110",
  49339=>"111000101",
  49340=>"000000000",
  49341=>"011011111",
  49342=>"110000010",
  49343=>"111111000",
  49344=>"000000001",
  49345=>"111000000",
  49346=>"110010110",
  49347=>"001000010",
  49348=>"100001001",
  49349=>"100000000",
  49350=>"001111110",
  49351=>"001101111",
  49352=>"111001100",
  49353=>"110110000",
  49354=>"110001110",
  49355=>"110110000",
  49356=>"110110010",
  49357=>"011010100",
  49358=>"000000001",
  49359=>"000110110",
  49360=>"000000011",
  49361=>"110110110",
  49362=>"010010100",
  49363=>"110111110",
  49364=>"000000001",
  49365=>"100100110",
  49366=>"101001110",
  49367=>"001000000",
  49368=>"111000000",
  49369=>"000110000",
  49370=>"100100001",
  49371=>"000000111",
  49372=>"000000111",
  49373=>"111101100",
  49374=>"110000000",
  49375=>"110000000",
  49376=>"000110010",
  49377=>"001000111",
  49378=>"000000000",
  49379=>"101100111",
  49380=>"110110000",
  49381=>"101001001",
  49382=>"000001100",
  49383=>"010000000",
  49384=>"110110100",
  49385=>"001001101",
  49386=>"001011001",
  49387=>"000000011",
  49388=>"110110110",
  49389=>"110001100",
  49390=>"010011000",
  49391=>"000000000",
  49392=>"110110000",
  49393=>"011001000",
  49394=>"000000001",
  49395=>"100100000",
  49396=>"000001001",
  49397=>"101111111",
  49398=>"000000110",
  49399=>"000000000",
  49400=>"000000001",
  49401=>"000001011",
  49402=>"001001011",
  49403=>"000001111",
  49404=>"111001010",
  49405=>"110110000",
  49406=>"011011110",
  49407=>"000010110",
  49408=>"011001000",
  49409=>"000011010",
  49410=>"100000000",
  49411=>"100101011",
  49412=>"001111111",
  49413=>"011000000",
  49414=>"100110110",
  49415=>"000011111",
  49416=>"000100111",
  49417=>"000100000",
  49418=>"100000001",
  49419=>"101100111",
  49420=>"011011001",
  49421=>"111101101",
  49422=>"000010111",
  49423=>"000100111",
  49424=>"000111011",
  49425=>"100101111",
  49426=>"000110000",
  49427=>"110001011",
  49428=>"111111111",
  49429=>"110101100",
  49430=>"000001000",
  49431=>"101110010",
  49432=>"000000000",
  49433=>"111111101",
  49434=>"011101010",
  49435=>"000100101",
  49436=>"101011011",
  49437=>"101100000",
  49438=>"110000000",
  49439=>"000111000",
  49440=>"000101101",
  49441=>"000111001",
  49442=>"001011010",
  49443=>"011111000",
  49444=>"111111110",
  49445=>"011000000",
  49446=>"111100100",
  49447=>"000000000",
  49448=>"011111111",
  49449=>"001110010",
  49450=>"100000011",
  49451=>"010010000",
  49452=>"000001110",
  49453=>"111111111",
  49454=>"111110000",
  49455=>"000001000",
  49456=>"111000000",
  49457=>"110110011",
  49458=>"111101000",
  49459=>"000011011",
  49460=>"000000000",
  49461=>"010111010",
  49462=>"110000001",
  49463=>"100100100",
  49464=>"111000000",
  49465=>"000000101",
  49466=>"000000100",
  49467=>"010010011",
  49468=>"110110100",
  49469=>"111111000",
  49470=>"010000000",
  49471=>"100000000",
  49472=>"101100111",
  49473=>"011000011",
  49474=>"000100100",
  49475=>"001100100",
  49476=>"110011000",
  49477=>"101100011",
  49478=>"000010000",
  49479=>"111010010",
  49480=>"101101101",
  49481=>"000000000",
  49482=>"101000011",
  49483=>"011011011",
  49484=>"100000000",
  49485=>"010010011",
  49486=>"011011111",
  49487=>"001011101",
  49488=>"100101000",
  49489=>"111101111",
  49490=>"110100011",
  49491=>"011000001",
  49492=>"010100000",
  49493=>"100111101",
  49494=>"011000000",
  49495=>"000110010",
  49496=>"110100001",
  49497=>"000001001",
  49498=>"110110000",
  49499=>"010010011",
  49500=>"111010000",
  49501=>"001001001",
  49502=>"000011111",
  49503=>"000000000",
  49504=>"111011000",
  49505=>"101111111",
  49506=>"000000100",
  49507=>"100100000",
  49508=>"000000100",
  49509=>"100110000",
  49510=>"000001000",
  49511=>"011000100",
  49512=>"010000101",
  49513=>"000000111",
  49514=>"010111011",
  49515=>"100000010",
  49516=>"111010000",
  49517=>"000000000",
  49518=>"011100000",
  49519=>"011010100",
  49520=>"001110111",
  49521=>"000000101",
  49522=>"001010111",
  49523=>"000011011",
  49524=>"010010011",
  49525=>"100000000",
  49526=>"000111111",
  49527=>"011011000",
  49528=>"000010010",
  49529=>"001000011",
  49530=>"000111111",
  49531=>"000011001",
  49532=>"101110011",
  49533=>"100000000",
  49534=>"111000100",
  49535=>"000000100",
  49536=>"111001010",
  49537=>"111011000",
  49538=>"100100010",
  49539=>"111101000",
  49540=>"000000011",
  49541=>"111101111",
  49542=>"011000100",
  49543=>"000011001",
  49544=>"010001111",
  49545=>"111111111",
  49546=>"111000000",
  49547=>"110000010",
  49548=>"000100101",
  49549=>"100100111",
  49550=>"000000100",
  49551=>"000000001",
  49552=>"000000111",
  49553=>"000000000",
  49554=>"000000000",
  49555=>"000011111",
  49556=>"000011101",
  49557=>"000000111",
  49558=>"110000101",
  49559=>"100001111",
  49560=>"000011011",
  49561=>"000000111",
  49562=>"111100000",
  49563=>"000000111",
  49564=>"100000000",
  49565=>"010000101",
  49566=>"111111011",
  49567=>"111010000",
  49568=>"101011000",
  49569=>"100000010",
  49570=>"001000000",
  49571=>"011000000",
  49572=>"000000000",
  49573=>"100110110",
  49574=>"000110000",
  49575=>"110111011",
  49576=>"000010111",
  49577=>"000010011",
  49578=>"110000101",
  49579=>"000011000",
  49580=>"101111101",
  49581=>"100100011",
  49582=>"001001111",
  49583=>"011111101",
  49584=>"000000000",
  49585=>"001000110",
  49586=>"100001111",
  49587=>"000100001",
  49588=>"000000000",
  49589=>"111111111",
  49590=>"011011011",
  49591=>"011011000",
  49592=>"001010000",
  49593=>"001111111",
  49594=>"011111010",
  49595=>"111100000",
  49596=>"011001000",
  49597=>"111111000",
  49598=>"001000001",
  49599=>"000000001",
  49600=>"100000000",
  49601=>"111000111",
  49602=>"000000011",
  49603=>"000110000",
  49604=>"000011000",
  49605=>"110111101",
  49606=>"101000010",
  49607=>"010011000",
  49608=>"101111000",
  49609=>"111100110",
  49610=>"111111011",
  49611=>"001011011",
  49612=>"110000100",
  49613=>"101011010",
  49614=>"011111010",
  49615=>"100110001",
  49616=>"110101111",
  49617=>"001000110",
  49618=>"010000100",
  49619=>"100011011",
  49620=>"000000100",
  49621=>"110011001",
  49622=>"100000000",
  49623=>"000011000",
  49624=>"111111000",
  49625=>"011101111",
  49626=>"011011010",
  49627=>"000000110",
  49628=>"111100000",
  49629=>"011000011",
  49630=>"011100110",
  49631=>"000000000",
  49632=>"000011000",
  49633=>"100000100",
  49634=>"000100111",
  49635=>"010100111",
  49636=>"101000000",
  49637=>"110101000",
  49638=>"111101110",
  49639=>"010000010",
  49640=>"100101111",
  49641=>"101101000",
  49642=>"000100000",
  49643=>"100111001",
  49644=>"000100111",
  49645=>"001011111",
  49646=>"000100000",
  49647=>"010010000",
  49648=>"100110111",
  49649=>"001111100",
  49650=>"100100000",
  49651=>"100000110",
  49652=>"110111101",
  49653=>"100111100",
  49654=>"000111000",
  49655=>"001000000",
  49656=>"000001111",
  49657=>"101101110",
  49658=>"011011010",
  49659=>"100100011",
  49660=>"010001000",
  49661=>"101001001",
  49662=>"111111011",
  49663=>"000000000",
  49664=>"001001010",
  49665=>"000111011",
  49666=>"101001101",
  49667=>"001001010",
  49668=>"110100110",
  49669=>"000000101",
  49670=>"111101101",
  49671=>"111101000",
  49672=>"110000000",
  49673=>"000000100",
  49674=>"111111001",
  49675=>"011000000",
  49676=>"000000100",
  49677=>"010011110",
  49678=>"010011010",
  49679=>"111111111",
  49680=>"110000100",
  49681=>"100000101",
  49682=>"010111011",
  49683=>"001000001",
  49684=>"101101101",
  49685=>"001000011",
  49686=>"111111011",
  49687=>"001000010",
  49688=>"101100000",
  49689=>"111101100",
  49690=>"110000000",
  49691=>"000000000",
  49692=>"111111010",
  49693=>"001000100",
  49694=>"111111111",
  49695=>"011110010",
  49696=>"011111001",
  49697=>"000000001",
  49698=>"001010111",
  49699=>"000000000",
  49700=>"100100100",
  49701=>"000001111",
  49702=>"111010010",
  49703=>"000100100",
  49704=>"110111000",
  49705=>"101001101",
  49706=>"101101111",
  49707=>"000111111",
  49708=>"010101100",
  49709=>"111111001",
  49710=>"001000101",
  49711=>"111001000",
  49712=>"110011000",
  49713=>"111100000",
  49714=>"000110011",
  49715=>"111101101",
  49716=>"001001000",
  49717=>"011001001",
  49718=>"000000111",
  49719=>"100000100",
  49720=>"010101000",
  49721=>"000000100",
  49722=>"101101111",
  49723=>"011000000",
  49724=>"011011000",
  49725=>"011111011",
  49726=>"000000000",
  49727=>"110110100",
  49728=>"101000101",
  49729=>"000111110",
  49730=>"010000000",
  49731=>"011001000",
  49732=>"111111010",
  49733=>"100100000",
  49734=>"010111000",
  49735=>"010010001",
  49736=>"001011011",
  49737=>"111001001",
  49738=>"000101101",
  49739=>"110000110",
  49740=>"000000111",
  49741=>"001010000",
  49742=>"111011001",
  49743=>"111101100",
  49744=>"000010010",
  49745=>"000110110",
  49746=>"111111101",
  49747=>"111100000",
  49748=>"000000110",
  49749=>"100001011",
  49750=>"011011001",
  49751=>"000100101",
  49752=>"000111011",
  49753=>"100100101",
  49754=>"101001011",
  49755=>"100001111",
  49756=>"111001000",
  49757=>"101001101",
  49758=>"000111111",
  49759=>"001000000",
  49760=>"111111010",
  49761=>"010000000",
  49762=>"111111101",
  49763=>"001100000",
  49764=>"111111000",
  49765=>"100111110",
  49766=>"010011111",
  49767=>"111011011",
  49768=>"010111011",
  49769=>"101100100",
  49770=>"000010010",
  49771=>"111111000",
  49772=>"111101101",
  49773=>"100110111",
  49774=>"111010010",
  49775=>"000100101",
  49776=>"110110000",
  49777=>"000001000",
  49778=>"000100000",
  49779=>"111000100",
  49780=>"101111011",
  49781=>"000000111",
  49782=>"000001101",
  49783=>"110000000",
  49784=>"000001111",
  49785=>"011011001",
  49786=>"100110000",
  49787=>"000000000",
  49788=>"111000000",
  49789=>"110000000",
  49790=>"010010111",
  49791=>"101000001",
  49792=>"101101111",
  49793=>"100010000",
  49794=>"111100010",
  49795=>"111011000",
  49796=>"001000000",
  49797=>"010000000",
  49798=>"100110110",
  49799=>"000000111",
  49800=>"111001000",
  49801=>"000101101",
  49802=>"100111101",
  49803=>"111000100",
  49804=>"110111111",
  49805=>"001000100",
  49806=>"000011111",
  49807=>"001001101",
  49808=>"100110110",
  49809=>"010110011",
  49810=>"101000010",
  49811=>"110000000",
  49812=>"011011001",
  49813=>"100000100",
  49814=>"000000101",
  49815=>"001011001",
  49816=>"010110110",
  49817=>"000010111",
  49818=>"010000110",
  49819=>"000100000",
  49820=>"001101100",
  49821=>"110111101",
  49822=>"100000000",
  49823=>"000000101",
  49824=>"100100110",
  49825=>"101101000",
  49826=>"111000000",
  49827=>"000100111",
  49828=>"000000101",
  49829=>"111001011",
  49830=>"111010000",
  49831=>"000000110",
  49832=>"010000001",
  49833=>"110110111",
  49834=>"000100000",
  49835=>"000000000",
  49836=>"010000000",
  49837=>"111111000",
  49838=>"000011001",
  49839=>"111010000",
  49840=>"000010011",
  49841=>"010001001",
  49842=>"100100111",
  49843=>"000010110",
  49844=>"011011110",
  49845=>"110101111",
  49846=>"111100000",
  49847=>"010111000",
  49848=>"101100000",
  49849=>"011000000",
  49850=>"010010010",
  49851=>"000101111",
  49852=>"100000110",
  49853=>"010111011",
  49854=>"101001000",
  49855=>"000101000",
  49856=>"101001101",
  49857=>"101100100",
  49858=>"100110110",
  49859=>"110100100",
  49860=>"111101111",
  49861=>"111110000",
  49862=>"011011101",
  49863=>"000000111",
  49864=>"010000110",
  49865=>"001000010",
  49866=>"101111101",
  49867=>"111111110",
  49868=>"001000000",
  49869=>"110110000",
  49870=>"100000011",
  49871=>"000001111",
  49872=>"101001000",
  49873=>"110110100",
  49874=>"111101100",
  49875=>"011000100",
  49876=>"000000100",
  49877=>"000100110",
  49878=>"100100000",
  49879=>"101110011",
  49880=>"100101111",
  49881=>"001010000",
  49882=>"011000000",
  49883=>"000000111",
  49884=>"111011100",
  49885=>"111010010",
  49886=>"101001010",
  49887=>"111111000",
  49888=>"111000000",
  49889=>"111110110",
  49890=>"101111110",
  49891=>"110110000",
  49892=>"111111111",
  49893=>"101000000",
  49894=>"011000000",
  49895=>"000100100",
  49896=>"000000000",
  49897=>"101111000",
  49898=>"100100000",
  49899=>"100000010",
  49900=>"000000010",
  49901=>"111111110",
  49902=>"001000000",
  49903=>"111010001",
  49904=>"111000000",
  49905=>"011011101",
  49906=>"111000000",
  49907=>"110011010",
  49908=>"100011101",
  49909=>"100010010",
  49910=>"000000000",
  49911=>"100111111",
  49912=>"000000111",
  49913=>"100001111",
  49914=>"000000000",
  49915=>"111111100",
  49916=>"111111110",
  49917=>"011111010",
  49918=>"000000000",
  49919=>"000101101",
  49920=>"111111111",
  49921=>"111011100",
  49922=>"100100110",
  49923=>"010100001",
  49924=>"111110111",
  49925=>"110000101",
  49926=>"101000101",
  49927=>"000111111",
  49928=>"011001001",
  49929=>"000000001",
  49930=>"001010000",
  49931=>"000000000",
  49932=>"000100000",
  49933=>"000000100",
  49934=>"101100010",
  49935=>"100111110",
  49936=>"000000000",
  49937=>"110010011",
  49938=>"111111011",
  49939=>"000101010",
  49940=>"010111111",
  49941=>"100111010",
  49942=>"000001101",
  49943=>"101111010",
  49944=>"100000000",
  49945=>"111111111",
  49946=>"111100100",
  49947=>"000000100",
  49948=>"110100111",
  49949=>"010111000",
  49950=>"111100011",
  49951=>"001000000",
  49952=>"111000001",
  49953=>"010100010",
  49954=>"000000010",
  49955=>"111100000",
  49956=>"100110100",
  49957=>"011111111",
  49958=>"111110000",
  49959=>"000000101",
  49960=>"111101000",
  49961=>"000000000",
  49962=>"000000000",
  49963=>"111010111",
  49964=>"000110000",
  49965=>"111011010",
  49966=>"011011110",
  49967=>"111100011",
  49968=>"010010101",
  49969=>"011110111",
  49970=>"101101111",
  49971=>"010111011",
  49972=>"000111111",
  49973=>"001111111",
  49974=>"000011010",
  49975=>"000111111",
  49976=>"010101111",
  49977=>"101111111",
  49978=>"011101101",
  49979=>"000001111",
  49980=>"011111111",
  49981=>"111111010",
  49982=>"101000001",
  49983=>"101001011",
  49984=>"111111101",
  49985=>"101111101",
  49986=>"000000011",
  49987=>"100101110",
  49988=>"001000000",
  49989=>"000101111",
  49990=>"000100000",
  49991=>"000110001",
  49992=>"001111001",
  49993=>"010001100",
  49994=>"001100000",
  49995=>"011110111",
  49996=>"111111111",
  49997=>"000111111",
  49998=>"000001001",
  49999=>"000111111",
  50000=>"000100111",
  50001=>"111111110",
  50002=>"101100101",
  50003=>"001101100",
  50004=>"000000000",
  50005=>"001110110",
  50006=>"010001000",
  50007=>"101000101",
  50008=>"000000000",
  50009=>"101110001",
  50010=>"101000000",
  50011=>"111011111",
  50012=>"110110000",
  50013=>"010000001",
  50014=>"000000111",
  50015=>"101101101",
  50016=>"001000101",
  50017=>"111000000",
  50018=>"000000100",
  50019=>"000100000",
  50020=>"000101100",
  50021=>"111100000",
  50022=>"110101111",
  50023=>"100101111",
  50024=>"000100111",
  50025=>"111101111",
  50026=>"000000000",
  50027=>"111111100",
  50028=>"000111101",
  50029=>"000111000",
  50030=>"000100101",
  50031=>"100000010",
  50032=>"000001101",
  50033=>"111011000",
  50034=>"111011011",
  50035=>"111001010",
  50036=>"000101011",
  50037=>"000001111",
  50038=>"111000000",
  50039=>"001010001",
  50040=>"000001000",
  50041=>"010000001",
  50042=>"010000101",
  50043=>"000000000",
  50044=>"110000010",
  50045=>"111110011",
  50046=>"010101111",
  50047=>"101000000",
  50048=>"110110101",
  50049=>"000000010",
  50050=>"000010111",
  50051=>"000010010",
  50052=>"000011010",
  50053=>"011000010",
  50054=>"100111110",
  50055=>"111111011",
  50056=>"000100111",
  50057=>"000010011",
  50058=>"111001000",
  50059=>"010001010",
  50060=>"000101101",
  50061=>"000000101",
  50062=>"010111111",
  50063=>"011000000",
  50064=>"111111011",
  50065=>"011110001",
  50066=>"010000011",
  50067=>"111000000",
  50068=>"110111111",
  50069=>"100101101",
  50070=>"110111010",
  50071=>"010100100",
  50072=>"001010100",
  50073=>"101111101",
  50074=>"010010110",
  50075=>"100000000",
  50076=>"101000000",
  50077=>"000000101",
  50078=>"011011010",
  50079=>"111101111",
  50080=>"100111010",
  50081=>"110011111",
  50082=>"011000000",
  50083=>"111000000",
  50084=>"011000010",
  50085=>"111111010",
  50086=>"110001011",
  50087=>"000000010",
  50088=>"110010010",
  50089=>"000000011",
  50090=>"011111111",
  50091=>"100100111",
  50092=>"010011101",
  50093=>"111000100",
  50094=>"011111101",
  50095=>"100000010",
  50096=>"000000001",
  50097=>"100000100",
  50098=>"110111000",
  50099=>"111001000",
  50100=>"101111001",
  50101=>"111010010",
  50102=>"111111000",
  50103=>"110000011",
  50104=>"111011001",
  50105=>"101111011",
  50106=>"011011011",
  50107=>"010110000",
  50108=>"000100000",
  50109=>"000000000",
  50110=>"100000100",
  50111=>"000000101",
  50112=>"111000000",
  50113=>"010111011",
  50114=>"110110000",
  50115=>"000001000",
  50116=>"010010000",
  50117=>"000111100",
  50118=>"111111100",
  50119=>"111100011",
  50120=>"000000000",
  50121=>"000000000",
  50122=>"000000011",
  50123=>"000111111",
  50124=>"111000000",
  50125=>"001010110",
  50126=>"111010010",
  50127=>"011111111",
  50128=>"101000000",
  50129=>"001111111",
  50130=>"110110111",
  50131=>"001101111",
  50132=>"000101010",
  50133=>"111110110",
  50134=>"101000001",
  50135=>"000000011",
  50136=>"111111000",
  50137=>"000000000",
  50138=>"011100100",
  50139=>"111100101",
  50140=>"100101111",
  50141=>"100101100",
  50142=>"001010000",
  50143=>"100000101",
  50144=>"111000000",
  50145=>"111000001",
  50146=>"000000000",
  50147=>"101111111",
  50148=>"111000000",
  50149=>"111100101",
  50150=>"100000000",
  50151=>"111010110",
  50152=>"100100000",
  50153=>"001100100",
  50154=>"110011010",
  50155=>"111100101",
  50156=>"000000000",
  50157=>"111001101",
  50158=>"111101000",
  50159=>"000000000",
  50160=>"000000011",
  50161=>"001111000",
  50162=>"001001100",
  50163=>"100001111",
  50164=>"001110111",
  50165=>"100001011",
  50166=>"110000000",
  50167=>"111001011",
  50168=>"010000000",
  50169=>"010111010",
  50170=>"100000101",
  50171=>"011110111",
  50172=>"111111111",
  50173=>"111101111",
  50174=>"000011011",
  50175=>"110111111",
  50176=>"101101110",
  50177=>"111111111",
  50178=>"011010101",
  50179=>"000000011",
  50180=>"011011011",
  50181=>"010111000",
  50182=>"101000000",
  50183=>"100110000",
  50184=>"110111100",
  50185=>"000001001",
  50186=>"001111111",
  50187=>"010100000",
  50188=>"011110000",
  50189=>"000100111",
  50190=>"110100001",
  50191=>"000000001",
  50192=>"100000000",
  50193=>"101111111",
  50194=>"111110000",
  50195=>"001000000",
  50196=>"111111111",
  50197=>"000011011",
  50198=>"110101111",
  50199=>"010010011",
  50200=>"000000111",
  50201=>"001011000",
  50202=>"111111111",
  50203=>"011000000",
  50204=>"000100100",
  50205=>"011001100",
  50206=>"011011010",
  50207=>"001101111",
  50208=>"100110000",
  50209=>"100111111",
  50210=>"111101001",
  50211=>"011000000",
  50212=>"010000000",
  50213=>"000000011",
  50214=>"000011111",
  50215=>"000000000",
  50216=>"000011111",
  50217=>"000111111",
  50218=>"100001111",
  50219=>"000101000",
  50220=>"000001001",
  50221=>"101110111",
  50222=>"110011111",
  50223=>"000000000",
  50224=>"000110111",
  50225=>"001000000",
  50226=>"101110100",
  50227=>"010111000",
  50228=>"111011001",
  50229=>"100001111",
  50230=>"010111111",
  50231=>"001000000",
  50232=>"010111010",
  50233=>"111100000",
  50234=>"100000000",
  50235=>"111000001",
  50236=>"001011110",
  50237=>"110111111",
  50238=>"100000000",
  50239=>"111010110",
  50240=>"111111000",
  50241=>"000000000",
  50242=>"100011100",
  50243=>"101000000",
  50244=>"000111111",
  50245=>"000100100",
  50246=>"101000000",
  50247=>"001001101",
  50248=>"001110000",
  50249=>"000100100",
  50250=>"000000000",
  50251=>"000000100",
  50252=>"100000000",
  50253=>"000000000",
  50254=>"111110000",
  50255=>"111001111",
  50256=>"000010011",
  50257=>"111011101",
  50258=>"011001000",
  50259=>"100111000",
  50260=>"001000000",
  50261=>"011111111",
  50262=>"010011000",
  50263=>"001000000",
  50264=>"101000100",
  50265=>"001101001",
  50266=>"110111111",
  50267=>"010110110",
  50268=>"000010100",
  50269=>"111111010",
  50270=>"000011111",
  50271=>"001000011",
  50272=>"101000000",
  50273=>"000000000",
  50274=>"000000100",
  50275=>"011101001",
  50276=>"000111111",
  50277=>"111111100",
  50278=>"100000000",
  50279=>"111111111",
  50280=>"111111111",
  50281=>"001000111",
  50282=>"010111111",
  50283=>"001110000",
  50284=>"111110000",
  50285=>"000011111",
  50286=>"010000100",
  50287=>"110000000",
  50288=>"111110111",
  50289=>"111111011",
  50290=>"101111011",
  50291=>"111100000",
  50292=>"000011110",
  50293=>"000000100",
  50294=>"111111010",
  50295=>"000111010",
  50296=>"001111111",
  50297=>"000000000",
  50298=>"101010111",
  50299=>"011000101",
  50300=>"111011010",
  50301=>"011111001",
  50302=>"001111111",
  50303=>"000000000",
  50304=>"000000000",
  50305=>"011111111",
  50306=>"000000111",
  50307=>"000000000",
  50308=>"011000000",
  50309=>"111101001",
  50310=>"000000000",
  50311=>"001000000",
  50312=>"110011001",
  50313=>"111100100",
  50314=>"111100100",
  50315=>"001001000",
  50316=>"000000101",
  50317=>"010011111",
  50318=>"000000000",
  50319=>"100000000",
  50320=>"000000000",
  50321=>"011010000",
  50322=>"000011111",
  50323=>"111111000",
  50324=>"110010010",
  50325=>"110111000",
  50326=>"111100100",
  50327=>"011000000",
  50328=>"000110000",
  50329=>"000111001",
  50330=>"111000000",
  50331=>"111000000",
  50332=>"111101000",
  50333=>"111000000",
  50334=>"011010000",
  50335=>"111000000",
  50336=>"110100010",
  50337=>"111111000",
  50338=>"000000111",
  50339=>"001000000",
  50340=>"010111011",
  50341=>"000000010",
  50342=>"010011111",
  50343=>"111101100",
  50344=>"101011101",
  50345=>"100000011",
  50346=>"110000000",
  50347=>"000000110",
  50348=>"101000001",
  50349=>"000000110",
  50350=>"000010001",
  50351=>"100000001",
  50352=>"100000000",
  50353=>"100110000",
  50354=>"000000101",
  50355=>"111110110",
  50356=>"000111000",
  50357=>"101000111",
  50358=>"000010111",
  50359=>"000000000",
  50360=>"110101011",
  50361=>"111001000",
  50362=>"000000010",
  50363=>"000100110",
  50364=>"011001010",
  50365=>"011111011",
  50366=>"111111110",
  50367=>"101111101",
  50368=>"000000000",
  50369=>"100000100",
  50370=>"011011000",
  50371=>"110110110",
  50372=>"111000100",
  50373=>"101110111",
  50374=>"101000011",
  50375=>"010000000",
  50376=>"111111100",
  50377=>"111101101",
  50378=>"000111111",
  50379=>"110000111",
  50380=>"000000000",
  50381=>"111110101",
  50382=>"101101111",
  50383=>"010111000",
  50384=>"011010010",
  50385=>"000100000",
  50386=>"000000000",
  50387=>"000000000",
  50388=>"111000100",
  50389=>"001011011",
  50390=>"111000000",
  50391=>"000001011",
  50392=>"101000000",
  50393=>"111101111",
  50394=>"111011001",
  50395=>"000100100",
  50396=>"011011010",
  50397=>"000000111",
  50398=>"100000000",
  50399=>"001010001",
  50400=>"010110100",
  50401=>"001010100",
  50402=>"111111011",
  50403=>"111100000",
  50404=>"000000100",
  50405=>"111000000",
  50406=>"111000000",
  50407=>"000011100",
  50408=>"000111111",
  50409=>"000111110",
  50410=>"000110011",
  50411=>"100100000",
  50412=>"111010000",
  50413=>"111101000",
  50414=>"010010111",
  50415=>"011011000",
  50416=>"111101000",
  50417=>"001011111",
  50418=>"010000000",
  50419=>"110111111",
  50420=>"000111011",
  50421=>"111000101",
  50422=>"100000000",
  50423=>"001001001",
  50424=>"000111011",
  50425=>"101111110",
  50426=>"000011000",
  50427=>"010000000",
  50428=>"101000000",
  50429=>"001000000",
  50430=>"000100110",
  50431=>"111000000",
  50432=>"011000000",
  50433=>"010110011",
  50434=>"001000000",
  50435=>"110001111",
  50436=>"111111011",
  50437=>"111110000",
  50438=>"110111110",
  50439=>"111111111",
  50440=>"111001000",
  50441=>"111001101",
  50442=>"100100010",
  50443=>"000000000",
  50444=>"111111101",
  50445=>"011111001",
  50446=>"011000111",
  50447=>"000011100",
  50448=>"110111010",
  50449=>"000000100",
  50450=>"111000111",
  50451=>"111000000",
  50452=>"111101100",
  50453=>"111111000",
  50454=>"000000000",
  50455=>"111101111",
  50456=>"010110010",
  50457=>"111011000",
  50458=>"101111011",
  50459=>"000111111",
  50460=>"011010010",
  50461=>"101001001",
  50462=>"111000100",
  50463=>"000011111",
  50464=>"000000000",
  50465=>"111111111",
  50466=>"000001001",
  50467=>"000111101",
  50468=>"000000111",
  50469=>"111001000",
  50470=>"111100000",
  50471=>"000000000",
  50472=>"101111001",
  50473=>"101111111",
  50474=>"111000101",
  50475=>"000111110",
  50476=>"001111011",
  50477=>"111110111",
  50478=>"111111000",
  50479=>"100111111",
  50480=>"111111111",
  50481=>"001001000",
  50482=>"000000001",
  50483=>"110111110",
  50484=>"000000000",
  50485=>"010001100",
  50486=>"000000000",
  50487=>"111001000",
  50488=>"111000000",
  50489=>"101000111",
  50490=>"000110111",
  50491=>"000000010",
  50492=>"100001000",
  50493=>"111111011",
  50494=>"010000110",
  50495=>"000100100",
  50496=>"000000000",
  50497=>"110010000",
  50498=>"111111111",
  50499=>"100000000",
  50500=>"111111000",
  50501=>"111111101",
  50502=>"000000000",
  50503=>"010110000",
  50504=>"110001010",
  50505=>"111111000",
  50506=>"111111111",
  50507=>"000000010",
  50508=>"111111111",
  50509=>"100100000",
  50510=>"110110110",
  50511=>"011111111",
  50512=>"001101101",
  50513=>"000110101",
  50514=>"111110111",
  50515=>"111010000",
  50516=>"000000000",
  50517=>"000000000",
  50518=>"110110000",
  50519=>"111011111",
  50520=>"010011000",
  50521=>"010010111",
  50522=>"100101100",
  50523=>"000000011",
  50524=>"000110110",
  50525=>"010011011",
  50526=>"000000000",
  50527=>"001000000",
  50528=>"111001111",
  50529=>"001011110",
  50530=>"101101101",
  50531=>"000111110",
  50532=>"111111111",
  50533=>"100100110",
  50534=>"111111011",
  50535=>"111000000",
  50536=>"011010010",
  50537=>"110111110",
  50538=>"110110100",
  50539=>"000110010",
  50540=>"100101101",
  50541=>"111111111",
  50542=>"111010000",
  50543=>"010010010",
  50544=>"000000101",
  50545=>"110010010",
  50546=>"000000000",
  50547=>"111111111",
  50548=>"011000111",
  50549=>"101000000",
  50550=>"111111010",
  50551=>"000111111",
  50552=>"001100111",
  50553=>"100000101",
  50554=>"000001111",
  50555=>"111101111",
  50556=>"000000000",
  50557=>"111101100",
  50558=>"000000111",
  50559=>"101111101",
  50560=>"001001001",
  50561=>"000000000",
  50562=>"110000101",
  50563=>"010110100",
  50564=>"010011000",
  50565=>"000000011",
  50566=>"111010010",
  50567=>"011011011",
  50568=>"001111000",
  50569=>"000100000",
  50570=>"011010010",
  50571=>"000111001",
  50572=>"111001000",
  50573=>"001000110",
  50574=>"111011101",
  50575=>"110100000",
  50576=>"011101111",
  50577=>"000000000",
  50578=>"010000010",
  50579=>"010000010",
  50580=>"000110110",
  50581=>"111110111",
  50582=>"111000000",
  50583=>"101101100",
  50584=>"111111001",
  50585=>"111111110",
  50586=>"101110111",
  50587=>"101111111",
  50588=>"111000010",
  50589=>"000000000",
  50590=>"011011000",
  50591=>"000110100",
  50592=>"001000011",
  50593=>"010000111",
  50594=>"111111111",
  50595=>"111000000",
  50596=>"110100000",
  50597=>"101111111",
  50598=>"111111101",
  50599=>"111001001",
  50600=>"110000111",
  50601=>"011001011",
  50602=>"000000101",
  50603=>"001110111",
  50604=>"000000101",
  50605=>"111111000",
  50606=>"000000000",
  50607=>"100111111",
  50608=>"000000001",
  50609=>"100101111",
  50610=>"111111111",
  50611=>"100000000",
  50612=>"100101110",
  50613=>"111111010",
  50614=>"001000100",
  50615=>"101111100",
  50616=>"001000000",
  50617=>"000111111",
  50618=>"111111111",
  50619=>"010111111",
  50620=>"111111010",
  50621=>"001100101",
  50622=>"011000101",
  50623=>"000111000",
  50624=>"000000000",
  50625=>"011111110",
  50626=>"111110001",
  50627=>"101111011",
  50628=>"111111111",
  50629=>"000000100",
  50630=>"010111011",
  50631=>"101100111",
  50632=>"111000101",
  50633=>"000011001",
  50634=>"110111100",
  50635=>"111001000",
  50636=>"101000011",
  50637=>"000000000",
  50638=>"000000000",
  50639=>"000001101",
  50640=>"100110110",
  50641=>"010100010",
  50642=>"010101001",
  50643=>"110011111",
  50644=>"000000000",
  50645=>"010110000",
  50646=>"000000000",
  50647=>"111001111",
  50648=>"000000000",
  50649=>"000000000",
  50650=>"100000000",
  50651=>"111111110",
  50652=>"000000000",
  50653=>"111111011",
  50654=>"000011010",
  50655=>"111101111",
  50656=>"111111010",
  50657=>"101111111",
  50658=>"000000101",
  50659=>"100100000",
  50660=>"000111111",
  50661=>"101011111",
  50662=>"111111111",
  50663=>"000000001",
  50664=>"111001000",
  50665=>"010010111",
  50666=>"000010001",
  50667=>"000111001",
  50668=>"101001111",
  50669=>"000101101",
  50670=>"001001001",
  50671=>"110111001",
  50672=>"000000001",
  50673=>"010000010",
  50674=>"111001110",
  50675=>"110110110",
  50676=>"010001000",
  50677=>"000111001",
  50678=>"111000011",
  50679=>"000000010",
  50680=>"111000000",
  50681=>"010111111",
  50682=>"111000010",
  50683=>"000000001",
  50684=>"111000000",
  50685=>"111000000",
  50686=>"111111101",
  50687=>"100000000",
  50688=>"000111011",
  50689=>"010000101",
  50690=>"000011110",
  50691=>"110000000",
  50692=>"011100100",
  50693=>"010000110",
  50694=>"101000000",
  50695=>"111010111",
  50696=>"000000001",
  50697=>"010000000",
  50698=>"000000000",
  50699=>"101111100",
  50700=>"111000000",
  50701=>"011000000",
  50702=>"011100100",
  50703=>"011000000",
  50704=>"101110000",
  50705=>"110000000",
  50706=>"001101100",
  50707=>"000000101",
  50708=>"000011111",
  50709=>"010000010",
  50710=>"100111011",
  50711=>"100000000",
  50712=>"111101000",
  50713=>"010111111",
  50714=>"001000000",
  50715=>"011110110",
  50716=>"100111011",
  50717=>"111111011",
  50718=>"010000001",
  50719=>"010111111",
  50720=>"100010110",
  50721=>"111111111",
  50722=>"111000100",
  50723=>"000000010",
  50724=>"001001101",
  50725=>"000100100",
  50726=>"010010010",
  50727=>"010000000",
  50728=>"011010010",
  50729=>"101000001",
  50730=>"010000000",
  50731=>"110111100",
  50732=>"111101101",
  50733=>"111110000",
  50734=>"110111001",
  50735=>"111110011",
  50736=>"101000000",
  50737=>"101101100",
  50738=>"000001111",
  50739=>"100110110",
  50740=>"000000000",
  50741=>"011110110",
  50742=>"001000100",
  50743=>"000001111",
  50744=>"111000000",
  50745=>"100100000",
  50746=>"000101001",
  50747=>"000010101",
  50748=>"001011111",
  50749=>"111111111",
  50750=>"000000000",
  50751=>"001100111",
  50752=>"000001100",
  50753=>"010000110",
  50754=>"101101001",
  50755=>"001000100",
  50756=>"111000100",
  50757=>"010011101",
  50758=>"000000000",
  50759=>"010000100",
  50760=>"101100000",
  50761=>"111110111",
  50762=>"101100000",
  50763=>"111001010",
  50764=>"010000000",
  50765=>"001100000",
  50766=>"011011001",
  50767=>"100110000",
  50768=>"000000101",
  50769=>"000000000",
  50770=>"110000111",
  50771=>"110110001",
  50772=>"011010000",
  50773=>"100001001",
  50774=>"000000101",
  50775=>"000000000",
  50776=>"101001001",
  50777=>"100101100",
  50778=>"000001111",
  50779=>"111001000",
  50780=>"010100000",
  50781=>"001101001",
  50782=>"000000110",
  50783=>"101001000",
  50784=>"101111111",
  50785=>"010001100",
  50786=>"101000101",
  50787=>"000001101",
  50788=>"110111000",
  50789=>"011111111",
  50790=>"110111111",
  50791=>"010101110",
  50792=>"111010111",
  50793=>"010000000",
  50794=>"110100101",
  50795=>"000000000",
  50796=>"101001001",
  50797=>"111111000",
  50798=>"010000000",
  50799=>"000111101",
  50800=>"111111100",
  50801=>"111000000",
  50802=>"100100001",
  50803=>"010101000",
  50804=>"000001101",
  50805=>"000001000",
  50806=>"111010000",
  50807=>"000110111",
  50808=>"000000111",
  50809=>"100011111",
  50810=>"111101111",
  50811=>"101111010",
  50812=>"110011000",
  50813=>"001001100",
  50814=>"010110111",
  50815=>"000111101",
  50816=>"010100000",
  50817=>"001111101",
  50818=>"110011000",
  50819=>"110111011",
  50820=>"000101111",
  50821=>"100000010",
  50822=>"000101001",
  50823=>"000100001",
  50824=>"101111100",
  50825=>"111000000",
  50826=>"111111111",
  50827=>"000000110",
  50828=>"000010010",
  50829=>"100111101",
  50830=>"111110010",
  50831=>"001100010",
  50832=>"111111100",
  50833=>"111110101",
  50834=>"010000001",
  50835=>"011010010",
  50836=>"101111010",
  50837=>"011000000",
  50838=>"000011000",
  50839=>"101101100",
  50840=>"010110110",
  50841=>"010110110",
  50842=>"000111001",
  50843=>"000010110",
  50844=>"111010000",
  50845=>"000010010",
  50846=>"000000111",
  50847=>"111101000",
  50848=>"111100100",
  50849=>"010000111",
  50850=>"000001000",
  50851=>"000000000",
  50852=>"001100000",
  50853=>"110001101",
  50854=>"000001000",
  50855=>"000010111",
  50856=>"010000000",
  50857=>"111011110",
  50858=>"111111101",
  50859=>"001001000",
  50860=>"011111011",
  50861=>"000000000",
  50862=>"011100100",
  50863=>"000010010",
  50864=>"111010010",
  50865=>"101001010",
  50866=>"111101100",
  50867=>"100001000",
  50868=>"101111111",
  50869=>"111110101",
  50870=>"010000100",
  50871=>"010111011",
  50872=>"110110100",
  50873=>"100110000",
  50874=>"000111111",
  50875=>"111000111",
  50876=>"111111011",
  50877=>"110111111",
  50878=>"100000100",
  50879=>"010000011",
  50880=>"000100000",
  50881=>"111110010",
  50882=>"111010111",
  50883=>"101001001",
  50884=>"011000000",
  50885=>"110100100",
  50886=>"010000000",
  50887=>"010111011",
  50888=>"110111001",
  50889=>"010010110",
  50890=>"110111101",
  50891=>"010000010",
  50892=>"000001111",
  50893=>"011001000",
  50894=>"000001011",
  50895=>"000101111",
  50896=>"001000001",
  50897=>"100111011",
  50898=>"110000000",
  50899=>"111000101",
  50900=>"001001011",
  50901=>"101101111",
  50902=>"101101101",
  50903=>"111001110",
  50904=>"000011000",
  50905=>"001111101",
  50906=>"111101001",
  50907=>"010000000",
  50908=>"001101110",
  50909=>"011111000",
  50910=>"110101101",
  50911=>"111110110",
  50912=>"111010111",
  50913=>"101000000",
  50914=>"000000111",
  50915=>"110011100",
  50916=>"000101111",
  50917=>"101111111",
  50918=>"010000000",
  50919=>"100000011",
  50920=>"111000100",
  50921=>"000000111",
  50922=>"100000001",
  50923=>"001010100",
  50924=>"111000000",
  50925=>"000101000",
  50926=>"011010000",
  50927=>"000101010",
  50928=>"000110101",
  50929=>"011001001",
  50930=>"110000000",
  50931=>"001111101",
  50932=>"001011110",
  50933=>"000001111",
  50934=>"000000101",
  50935=>"110110011",
  50936=>"000000000",
  50937=>"111111111",
  50938=>"111101101",
  50939=>"111001111",
  50940=>"101111101",
  50941=>"010111011",
  50942=>"001000011",
  50943=>"111011010",
  50944=>"011111010",
  50945=>"111110000",
  50946=>"101000000",
  50947=>"001000010",
  50948=>"000100001",
  50949=>"111000001",
  50950=>"000101111",
  50951=>"000110010",
  50952=>"001001111",
  50953=>"110000000",
  50954=>"110110111",
  50955=>"110100011",
  50956=>"100000100",
  50957=>"001001000",
  50958=>"100100011",
  50959=>"101111100",
  50960=>"001000010",
  50961=>"011000100",
  50962=>"001000000",
  50963=>"111010010",
  50964=>"000010000",
  50965=>"101000001",
  50966=>"101000001",
  50967=>"100111011",
  50968=>"101101110",
  50969=>"110110101",
  50970=>"111111001",
  50971=>"011100101",
  50972=>"111101111",
  50973=>"101001111",
  50974=>"000010010",
  50975=>"001101100",
  50976=>"110001101",
  50977=>"000010000",
  50978=>"000000000",
  50979=>"000000000",
  50980=>"000111111",
  50981=>"000110100",
  50982=>"010000010",
  50983=>"000010011",
  50984=>"110111111",
  50985=>"110000000",
  50986=>"100100000",
  50987=>"101101101",
  50988=>"100111111",
  50989=>"101100000",
  50990=>"000000011",
  50991=>"011101111",
  50992=>"010110000",
  50993=>"011101001",
  50994=>"000111111",
  50995=>"000000111",
  50996=>"000100110",
  50997=>"111000001",
  50998=>"110100001",
  50999=>"000000010",
  51000=>"010111000",
  51001=>"101000000",
  51002=>"111101101",
  51003=>"011000111",
  51004=>"001110110",
  51005=>"111111111",
  51006=>"000010011",
  51007=>"110111001",
  51008=>"011000100",
  51009=>"101110000",
  51010=>"001000000",
  51011=>"011001001",
  51012=>"111001101",
  51013=>"010000000",
  51014=>"010111111",
  51015=>"111000010",
  51016=>"011000000",
  51017=>"001111101",
  51018=>"000001101",
  51019=>"111110111",
  51020=>"110101101",
  51021=>"101110000",
  51022=>"101111111",
  51023=>"100101111",
  51024=>"001001000",
  51025=>"111000000",
  51026=>"000010011",
  51027=>"001001001",
  51028=>"010010000",
  51029=>"001111111",
  51030=>"001111111",
  51031=>"001010010",
  51032=>"101111001",
  51033=>"101101011",
  51034=>"000100100",
  51035=>"000011111",
  51036=>"000110010",
  51037=>"111001001",
  51038=>"011111000",
  51039=>"100100000",
  51040=>"111100000",
  51041=>"101011011",
  51042=>"111000000",
  51043=>"000000101",
  51044=>"000111101",
  51045=>"101011100",
  51046=>"100110111",
  51047=>"101001101",
  51048=>"101001001",
  51049=>"000101111",
  51050=>"010010011",
  51051=>"111111101",
  51052=>"101001001",
  51053=>"001011000",
  51054=>"000000000",
  51055=>"000011011",
  51056=>"010110111",
  51057=>"111010111",
  51058=>"011001110",
  51059=>"100000111",
  51060=>"101011010",
  51061=>"101001000",
  51062=>"111111110",
  51063=>"100100000",
  51064=>"011000000",
  51065=>"000010010",
  51066=>"000110110",
  51067=>"011101101",
  51068=>"000111110",
  51069=>"011101101",
  51070=>"111101111",
  51071=>"000001101",
  51072=>"010000000",
  51073=>"110000000",
  51074=>"000000010",
  51075=>"000001000",
  51076=>"111010010",
  51077=>"010101001",
  51078=>"110001111",
  51079=>"000011011",
  51080=>"000000100",
  51081=>"000000000",
  51082=>"000011010",
  51083=>"010000000",
  51084=>"100100010",
  51085=>"110100000",
  51086=>"111001001",
  51087=>"000000000",
  51088=>"111001101",
  51089=>"111011101",
  51090=>"110110000",
  51091=>"000000000",
  51092=>"001110010",
  51093=>"111000000",
  51094=>"000000000",
  51095=>"010100000",
  51096=>"010111111",
  51097=>"000000000",
  51098=>"110111011",
  51099=>"000100000",
  51100=>"111101111",
  51101=>"111011011",
  51102=>"111011110",
  51103=>"000000101",
  51104=>"111000000",
  51105=>"111000000",
  51106=>"010101101",
  51107=>"110000101",
  51108=>"010100111",
  51109=>"110110010",
  51110=>"110000111",
  51111=>"010000000",
  51112=>"010101001",
  51113=>"000110110",
  51114=>"010000001",
  51115=>"000000000",
  51116=>"110111000",
  51117=>"000100101",
  51118=>"110100011",
  51119=>"000100110",
  51120=>"100110011",
  51121=>"000100110",
  51122=>"111100100",
  51123=>"001000101",
  51124=>"111001001",
  51125=>"100000100",
  51126=>"001100000",
  51127=>"111111001",
  51128=>"010111011",
  51129=>"000110111",
  51130=>"110101101",
  51131=>"111101010",
  51132=>"110000010",
  51133=>"111111011",
  51134=>"011001000",
  51135=>"000000111",
  51136=>"001000001",
  51137=>"000000101",
  51138=>"111001111",
  51139=>"011110111",
  51140=>"010010001",
  51141=>"100100110",
  51142=>"111111111",
  51143=>"101111111",
  51144=>"010101111",
  51145=>"010100101",
  51146=>"110001111",
  51147=>"101101000",
  51148=>"110011010",
  51149=>"000111010",
  51150=>"100111111",
  51151=>"111101111",
  51152=>"100101000",
  51153=>"101101100",
  51154=>"000011000",
  51155=>"011111100",
  51156=>"000010000",
  51157=>"000011011",
  51158=>"111000000",
  51159=>"111111111",
  51160=>"110101111",
  51161=>"000010010",
  51162=>"100000001",
  51163=>"000001101",
  51164=>"000100111",
  51165=>"000110101",
  51166=>"010011001",
  51167=>"010110010",
  51168=>"000010000",
  51169=>"101001001",
  51170=>"111101111",
  51171=>"000001101",
  51172=>"000010000",
  51173=>"110101110",
  51174=>"001001000",
  51175=>"110011000",
  51176=>"000010010",
  51177=>"000000000",
  51178=>"001011111",
  51179=>"111100111",
  51180=>"100110111",
  51181=>"000000010",
  51182=>"000000000",
  51183=>"000010011",
  51184=>"100100010",
  51185=>"000001000",
  51186=>"000001011",
  51187=>"110100101",
  51188=>"110010001",
  51189=>"000101100",
  51190=>"000000110",
  51191=>"111101101",
  51192=>"010000000",
  51193=>"101101011",
  51194=>"111101001",
  51195=>"000111010",
  51196=>"010111111",
  51197=>"000010010",
  51198=>"011011001",
  51199=>"001110010",
  51200=>"010010000",
  51201=>"111101111",
  51202=>"111010101",
  51203=>"000000111",
  51204=>"011001000",
  51205=>"000000000",
  51206=>"110100000",
  51207=>"000110111",
  51208=>"001001111",
  51209=>"010010000",
  51210=>"011001000",
  51211=>"010110110",
  51212=>"000000000",
  51213=>"000000000",
  51214=>"001011011",
  51215=>"001000010",
  51216=>"000000010",
  51217=>"111001000",
  51218=>"001001001",
  51219=>"101010111",
  51220=>"111101111",
  51221=>"111000101",
  51222=>"101011100",
  51223=>"000000000",
  51224=>"111000110",
  51225=>"010111111",
  51226=>"011111111",
  51227=>"110010000",
  51228=>"111100100",
  51229=>"110101011",
  51230=>"001000001",
  51231=>"001001111",
  51232=>"010000000",
  51233=>"011101111",
  51234=>"100011111",
  51235=>"010000000",
  51236=>"111100000",
  51237=>"000000100",
  51238=>"000101111",
  51239=>"101101101",
  51240=>"101000001",
  51241=>"000001000",
  51242=>"010011001",
  51243=>"110000010",
  51244=>"011011001",
  51245=>"010000111",
  51246=>"000101101",
  51247=>"000000100",
  51248=>"010101111",
  51249=>"101001001",
  51250=>"001100111",
  51251=>"010111111",
  51252=>"111110000",
  51253=>"001101111",
  51254=>"111000000",
  51255=>"000111010",
  51256=>"000111110",
  51257=>"000000100",
  51258=>"100100111",
  51259=>"011111110",
  51260=>"000100100",
  51261=>"111111001",
  51262=>"000000010",
  51263=>"000000101",
  51264=>"111010000",
  51265=>"000000000",
  51266=>"101010110",
  51267=>"001001011",
  51268=>"000000110",
  51269=>"001101001",
  51270=>"011010010",
  51271=>"010000000",
  51272=>"001101111",
  51273=>"000001011",
  51274=>"000000010",
  51275=>"010000000",
  51276=>"000111110",
  51277=>"111011001",
  51278=>"111000000",
  51279=>"001011110",
  51280=>"111111000",
  51281=>"111010001",
  51282=>"011000011",
  51283=>"011111110",
  51284=>"001001010",
  51285=>"000000100",
  51286=>"111111100",
  51287=>"010010000",
  51288=>"000000100",
  51289=>"100100011",
  51290=>"100101111",
  51291=>"110110001",
  51292=>"001001101",
  51293=>"001001011",
  51294=>"011101101",
  51295=>"111100100",
  51296=>"111000110",
  51297=>"000001111",
  51298=>"110111110",
  51299=>"001111110",
  51300=>"100111100",
  51301=>"011111111",
  51302=>"000000110",
  51303=>"111111100",
  51304=>"001001111",
  51305=>"001101001",
  51306=>"110101011",
  51307=>"000001001",
  51308=>"000101101",
  51309=>"111111000",
  51310=>"111110100",
  51311=>"000000111",
  51312=>"011011001",
  51313=>"001000110",
  51314=>"111000000",
  51315=>"000000100",
  51316=>"000000010",
  51317=>"101101111",
  51318=>"110110110",
  51319=>"101000010",
  51320=>"010100010",
  51321=>"110110000",
  51322=>"101101101",
  51323=>"000001111",
  51324=>"110110110",
  51325=>"110100000",
  51326=>"111010010",
  51327=>"000000010",
  51328=>"111111011",
  51329=>"101000111",
  51330=>"000101101",
  51331=>"111010111",
  51332=>"001101001",
  51333=>"100100111",
  51334=>"000000001",
  51335=>"111000011",
  51336=>"101101001",
  51337=>"110110110",
  51338=>"000101011",
  51339=>"111100000",
  51340=>"101000001",
  51341=>"001001000",
  51342=>"110010000",
  51343=>"001000001",
  51344=>"110100101",
  51345=>"000000000",
  51346=>"111100101",
  51347=>"010000101",
  51348=>"111010011",
  51349=>"000000000",
  51350=>"000111000",
  51351=>"100110001",
  51352=>"111110100",
  51353=>"000001110",
  51354=>"111110010",
  51355=>"000000110",
  51356=>"010010011",
  51357=>"011111010",
  51358=>"111111110",
  51359=>"000001010",
  51360=>"010100001",
  51361=>"000001111",
  51362=>"101001000",
  51363=>"000011011",
  51364=>"000001111",
  51365=>"011011010",
  51366=>"101001001",
  51367=>"001111110",
  51368=>"110011111",
  51369=>"000010111",
  51370=>"101101111",
  51371=>"111001000",
  51372=>"001100101",
  51373=>"000011111",
  51374=>"111111011",
  51375=>"110111111",
  51376=>"000000110",
  51377=>"001111100",
  51378=>"111111000",
  51379=>"001100110",
  51380=>"100110101",
  51381=>"000110111",
  51382=>"100000100",
  51383=>"000100001",
  51384=>"000011011",
  51385=>"110010110",
  51386=>"010000010",
  51387=>"011001000",
  51388=>"001001000",
  51389=>"111111010",
  51390=>"000001011",
  51391=>"000000100",
  51392=>"000001101",
  51393=>"110111000",
  51394=>"000000111",
  51395=>"101011000",
  51396=>"010001000",
  51397=>"000011001",
  51398=>"010100111",
  51399=>"010110110",
  51400=>"100111110",
  51401=>"000000000",
  51402=>"000010001",
  51403=>"010110110",
  51404=>"001000000",
  51405=>"011011111",
  51406=>"111011000",
  51407=>"100101000",
  51408=>"000111110",
  51409=>"111101000",
  51410=>"000110111",
  51411=>"101101100",
  51412=>"101101100",
  51413=>"111100000",
  51414=>"000000110",
  51415=>"111101001",
  51416=>"101001011",
  51417=>"011000111",
  51418=>"100100100",
  51419=>"000100000",
  51420=>"110100011",
  51421=>"000000000",
  51422=>"111110001",
  51423=>"001101111",
  51424=>"000000000",
  51425=>"001111011",
  51426=>"001001110",
  51427=>"100110110",
  51428=>"101000100",
  51429=>"110100101",
  51430=>"111110000",
  51431=>"111100100",
  51432=>"001111111",
  51433=>"110100110",
  51434=>"110010001",
  51435=>"111110111",
  51436=>"111010000",
  51437=>"101101101",
  51438=>"110010000",
  51439=>"000101111",
  51440=>"001010010",
  51441=>"010000100",
  51442=>"000000101",
  51443=>"000000110",
  51444=>"000100011",
  51445=>"101111010",
  51446=>"101000000",
  51447=>"100110110",
  51448=>"101000101",
  51449=>"111111111",
  51450=>"111111000",
  51451=>"001011111",
  51452=>"000001101",
  51453=>"010001000",
  51454=>"100100100",
  51455=>"000111111",
  51456=>"000001100",
  51457=>"010000000",
  51458=>"000000000",
  51459=>"000000000",
  51460=>"100011111",
  51461=>"111010001",
  51462=>"011111110",
  51463=>"000011011",
  51464=>"000110000",
  51465=>"101000000",
  51466=>"000000000",
  51467=>"101100010",
  51468=>"010100000",
  51469=>"000111110",
  51470=>"000001011",
  51471=>"000000000",
  51472=>"010011111",
  51473=>"110000110",
  51474=>"111000000",
  51475=>"000000101",
  51476=>"111110110",
  51477=>"010011111",
  51478=>"011101001",
  51479=>"000010111",
  51480=>"100000000",
  51481=>"111111111",
  51482=>"111111111",
  51483=>"101001000",
  51484=>"101000010",
  51485=>"000101000",
  51486=>"001010000",
  51487=>"000111111",
  51488=>"110000000",
  51489=>"001010010",
  51490=>"000000010",
  51491=>"101111111",
  51492=>"100110111",
  51493=>"001111111",
  51494=>"101000000",
  51495=>"011000000",
  51496=>"000111000",
  51497=>"001000110",
  51498=>"000000000",
  51499=>"000000010",
  51500=>"111110001",
  51501=>"111010100",
  51502=>"110110100",
  51503=>"111111110",
  51504=>"100000111",
  51505=>"001011100",
  51506=>"000111111",
  51507=>"111001110",
  51508=>"001000000",
  51509=>"001000000",
  51510=>"110000001",
  51511=>"000000000",
  51512=>"111010000",
  51513=>"000111111",
  51514=>"000000100",
  51515=>"000011111",
  51516=>"011110110",
  51517=>"111111111",
  51518=>"000000001",
  51519=>"000111100",
  51520=>"110000000",
  51521=>"001111001",
  51522=>"111010000",
  51523=>"101010000",
  51524=>"101000001",
  51525=>"000000010",
  51526=>"001101011",
  51527=>"111111111",
  51528=>"110111111",
  51529=>"101000001",
  51530=>"101000000",
  51531=>"101000110",
  51532=>"111010000",
  51533=>"001111000",
  51534=>"000011010",
  51535=>"010111101",
  51536=>"001101100",
  51537=>"110110110",
  51538=>"110110111",
  51539=>"011001100",
  51540=>"000000000",
  51541=>"111111001",
  51542=>"011111111",
  51543=>"110110111",
  51544=>"000100000",
  51545=>"000000001",
  51546=>"100111111",
  51547=>"011111111",
  51548=>"111011000",
  51549=>"001001001",
  51550=>"000111010",
  51551=>"110110001",
  51552=>"000000000",
  51553=>"101101100",
  51554=>"000000000",
  51555=>"001011100",
  51556=>"000000100",
  51557=>"000100000",
  51558=>"000000010",
  51559=>"111010000",
  51560=>"000010010",
  51561=>"000000000",
  51562=>"010000000",
  51563=>"111101111",
  51564=>"100001001",
  51565=>"000000000",
  51566=>"000000000",
  51567=>"000000000",
  51568=>"100100101",
  51569=>"110000000",
  51570=>"001001100",
  51571=>"100000101",
  51572=>"111001111",
  51573=>"011000000",
  51574=>"000110110",
  51575=>"010111010",
  51576=>"000010110",
  51577=>"001001111",
  51578=>"001000101",
  51579=>"000111011",
  51580=>"000100000",
  51581=>"000100001",
  51582=>"000000000",
  51583=>"101101100",
  51584=>"101111111",
  51585=>"111111001",
  51586=>"000011000",
  51587=>"000000010",
  51588=>"110000000",
  51589=>"011001001",
  51590=>"100111111",
  51591=>"100101100",
  51592=>"101011011",
  51593=>"111010111",
  51594=>"110000110",
  51595=>"111000001",
  51596=>"000111111",
  51597=>"101110101",
  51598=>"000001001",
  51599=>"101001001",
  51600=>"101111101",
  51601=>"111111111",
  51602=>"000000110",
  51603=>"111000100",
  51604=>"111000101",
  51605=>"110010000",
  51606=>"111000101",
  51607=>"001001000",
  51608=>"111111111",
  51609=>"000010010",
  51610=>"111001101",
  51611=>"111010000",
  51612=>"111111010",
  51613=>"111111111",
  51614=>"010000000",
  51615=>"111000001",
  51616=>"011111111",
  51617=>"110010111",
  51618=>"011111111",
  51619=>"110000000",
  51620=>"010000001",
  51621=>"110111011",
  51622=>"011100001",
  51623=>"010001100",
  51624=>"111110010",
  51625=>"000000000",
  51626=>"000000000",
  51627=>"011001111",
  51628=>"000011000",
  51629=>"000010000",
  51630=>"010101101",
  51631=>"010110010",
  51632=>"000111110",
  51633=>"000111100",
  51634=>"000100000",
  51635=>"000000000",
  51636=>"001101001",
  51637=>"000000000",
  51638=>"000010001",
  51639=>"000000000",
  51640=>"011000011",
  51641=>"111000111",
  51642=>"010110100",
  51643=>"010010111",
  51644=>"101101111",
  51645=>"111011000",
  51646=>"000011000",
  51647=>"110111111",
  51648=>"010111011",
  51649=>"000111101",
  51650=>"111001100",
  51651=>"001111001",
  51652=>"000000000",
  51653=>"100010110",
  51654=>"111111001",
  51655=>"010111110",
  51656=>"001000000",
  51657=>"011111101",
  51658=>"000000000",
  51659=>"000111011",
  51660=>"000011010",
  51661=>"000000000",
  51662=>"010100101",
  51663=>"000000011",
  51664=>"101111110",
  51665=>"000001010",
  51666=>"000111110",
  51667=>"100001001",
  51668=>"010111010",
  51669=>"000000110",
  51670=>"111000000",
  51671=>"100000000",
  51672=>"010111111",
  51673=>"000000101",
  51674=>"110111110",
  51675=>"111000001",
  51676=>"110000011",
  51677=>"000111000",
  51678=>"110110111",
  51679=>"000010111",
  51680=>"010111111",
  51681=>"111010110",
  51682=>"000111000",
  51683=>"100100101",
  51684=>"000110110",
  51685=>"010001000",
  51686=>"101001101",
  51687=>"000100100",
  51688=>"111111001",
  51689=>"111100000",
  51690=>"001000000",
  51691=>"001000001",
  51692=>"111111111",
  51693=>"110111111",
  51694=>"000000000",
  51695=>"010110111",
  51696=>"101101101",
  51697=>"111001100",
  51698=>"111010000",
  51699=>"000000000",
  51700=>"000000000",
  51701=>"101101101",
  51702=>"101001111",
  51703=>"100101111",
  51704=>"000111111",
  51705=>"011000000",
  51706=>"111101111",
  51707=>"111000001",
  51708=>"000000101",
  51709=>"001000010",
  51710=>"110110010",
  51711=>"010000110",
  51712=>"001001100",
  51713=>"111000001",
  51714=>"111110101",
  51715=>"000010110",
  51716=>"000100100",
  51717=>"100000000",
  51718=>"001101000",
  51719=>"000000110",
  51720=>"000110110",
  51721=>"111010010",
  51722=>"000000000",
  51723=>"111110111",
  51724=>"101111101",
  51725=>"101011111",
  51726=>"100001001",
  51727=>"111110000",
  51728=>"000000010",
  51729=>"110000011",
  51730=>"010111011",
  51731=>"110000000",
  51732=>"000111001",
  51733=>"110010000",
  51734=>"111011111",
  51735=>"111111111",
  51736=>"101101111",
  51737=>"111101001",
  51738=>"011000000",
  51739=>"100101111",
  51740=>"100000111",
  51741=>"000110111",
  51742=>"110000011",
  51743=>"000010000",
  51744=>"101111111",
  51745=>"001110101",
  51746=>"110010000",
  51747=>"010010000",
  51748=>"101100100",
  51749=>"101101100",
  51750=>"110111000",
  51751=>"000000000",
  51752=>"010111000",
  51753=>"101101101",
  51754=>"101101100",
  51755=>"010000111",
  51756=>"101100101",
  51757=>"101010000",
  51758=>"110100101",
  51759=>"111110111",
  51760=>"010000010",
  51761=>"001001001",
  51762=>"000010111",
  51763=>"101001010",
  51764=>"000000101",
  51765=>"010010100",
  51766=>"000000100",
  51767=>"000000111",
  51768=>"010111011",
  51769=>"000100000",
  51770=>"000000011",
  51771=>"101111011",
  51772=>"000100011",
  51773=>"111111111",
  51774=>"111010001",
  51775=>"100110000",
  51776=>"011111000",
  51777=>"010000000",
  51778=>"010110111",
  51779=>"001001100",
  51780=>"010111000",
  51781=>"000000110",
  51782=>"111111101",
  51783=>"110010011",
  51784=>"100100000",
  51785=>"100110011",
  51786=>"111111111",
  51787=>"000101001",
  51788=>"000000111",
  51789=>"001001000",
  51790=>"100100100",
  51791=>"111011000",
  51792=>"010000100",
  51793=>"111001111",
  51794=>"010011010",
  51795=>"011011000",
  51796=>"010111101",
  51797=>"001011101",
  51798=>"001011000",
  51799=>"001000111",
  51800=>"111111000",
  51801=>"001111011",
  51802=>"011110100",
  51803=>"011101100",
  51804=>"110111111",
  51805=>"000010001",
  51806=>"000010110",
  51807=>"100000001",
  51808=>"101000000",
  51809=>"010000000",
  51810=>"111001001",
  51811=>"110011111",
  51812=>"000101010",
  51813=>"111001110",
  51814=>"000101000",
  51815=>"010100000",
  51816=>"111110000",
  51817=>"110000001",
  51818=>"111000111",
  51819=>"000000000",
  51820=>"001100101",
  51821=>"000000000",
  51822=>"111011101",
  51823=>"010111111",
  51824=>"001101000",
  51825=>"110000001",
  51826=>"000000101",
  51827=>"000000000",
  51828=>"111111111",
  51829=>"000000100",
  51830=>"000000000",
  51831=>"000000111",
  51832=>"110111111",
  51833=>"010110111",
  51834=>"101010110",
  51835=>"000000000",
  51836=>"000110110",
  51837=>"100110000",
  51838=>"010110111",
  51839=>"000101000",
  51840=>"101100010",
  51841=>"110000100",
  51842=>"000111111",
  51843=>"000111110",
  51844=>"001000000",
  51845=>"010010000",
  51846=>"011001001",
  51847=>"101000001",
  51848=>"000101000",
  51849=>"100000000",
  51850=>"110100010",
  51851=>"000011100",
  51852=>"000110000",
  51853=>"000000010",
  51854=>"010111101",
  51855=>"101001001",
  51856=>"001101100",
  51857=>"111100000",
  51858=>"011101010",
  51859=>"111110111",
  51860=>"011111011",
  51861=>"000000111",
  51862=>"111111101",
  51863=>"001111011",
  51864=>"010010111",
  51865=>"000111111",
  51866=>"110010000",
  51867=>"010010010",
  51868=>"000011000",
  51869=>"010111011",
  51870=>"010010011",
  51871=>"111000000",
  51872=>"111011000",
  51873=>"111111110",
  51874=>"000010010",
  51875=>"111010111",
  51876=>"110011011",
  51877=>"111001011",
  51878=>"000101011",
  51879=>"000110000",
  51880=>"011000001",
  51881=>"011111111",
  51882=>"000010100",
  51883=>"001000000",
  51884=>"101111011",
  51885=>"000101100",
  51886=>"111010110",
  51887=>"111010000",
  51888=>"111111010",
  51889=>"001101000",
  51890=>"000000000",
  51891=>"001000100",
  51892=>"000011000",
  51893=>"110011111",
  51894=>"111011000",
  51895=>"000001000",
  51896=>"000001100",
  51897=>"100110110",
  51898=>"001101010",
  51899=>"111110111",
  51900=>"110111100",
  51901=>"011001111",
  51902=>"001011011",
  51903=>"011000010",
  51904=>"010110100",
  51905=>"100001000",
  51906=>"010000001",
  51907=>"101111111",
  51908=>"000000001",
  51909=>"110111011",
  51910=>"100100011",
  51911=>"000001111",
  51912=>"000101110",
  51913=>"111101101",
  51914=>"111011111",
  51915=>"010010000",
  51916=>"000010011",
  51917=>"000001011",
  51918=>"000100111",
  51919=>"000001111",
  51920=>"000110010",
  51921=>"011100110",
  51922=>"001101111",
  51923=>"010010110",
  51924=>"000011101",
  51925=>"110101001",
  51926=>"110111111",
  51927=>"110101011",
  51928=>"000111000",
  51929=>"000000010",
  51930=>"111110100",
  51931=>"000000000",
  51932=>"011110111",
  51933=>"010111110",
  51934=>"111111000",
  51935=>"011000011",
  51936=>"010111111",
  51937=>"100000111",
  51938=>"000011101",
  51939=>"100000000",
  51940=>"110000010",
  51941=>"011001011",
  51942=>"111111010",
  51943=>"101101111",
  51944=>"111100100",
  51945=>"011010110",
  51946=>"001000000",
  51947=>"001011111",
  51948=>"111110111",
  51949=>"001101101",
  51950=>"110010010",
  51951=>"000000110",
  51952=>"111111100",
  51953=>"011101110",
  51954=>"000000010",
  51955=>"100110000",
  51956=>"100111001",
  51957=>"100101000",
  51958=>"000000011",
  51959=>"111010001",
  51960=>"000010110",
  51961=>"110110101",
  51962=>"111111101",
  51963=>"000111111",
  51964=>"000000110",
  51965=>"101001100",
  51966=>"101011010",
  51967=>"111100111",
  51968=>"011001001",
  51969=>"000000001",
  51970=>"110110100",
  51971=>"101111110",
  51972=>"001001010",
  51973=>"000100110",
  51974=>"101111101",
  51975=>"100110111",
  51976=>"011001011",
  51977=>"001000111",
  51978=>"000000001",
  51979=>"000001000",
  51980=>"111001001",
  51981=>"000010001",
  51982=>"100100100",
  51983=>"101011000",
  51984=>"101000100",
  51985=>"000000011",
  51986=>"000000000",
  51987=>"000000111",
  51988=>"100111111",
  51989=>"110110110",
  51990=>"011001010",
  51991=>"000000000",
  51992=>"001000000",
  51993=>"110100000",
  51994=>"101111111",
  51995=>"000000001",
  51996=>"000000001",
  51997=>"000000000",
  51998=>"000000000",
  51999=>"111110010",
  52000=>"000000000",
  52001=>"010110110",
  52002=>"000001010",
  52003=>"001001001",
  52004=>"100100000",
  52005=>"000011010",
  52006=>"010010010",
  52007=>"011000111",
  52008=>"011110010",
  52009=>"010001101",
  52010=>"111110000",
  52011=>"110100000",
  52012=>"110110110",
  52013=>"000110111",
  52014=>"010011000",
  52015=>"101101010",
  52016=>"001000000",
  52017=>"001100111",
  52018=>"001001101",
  52019=>"001001111",
  52020=>"000000001",
  52021=>"000111110",
  52022=>"011000000",
  52023=>"011010000",
  52024=>"000100111",
  52025=>"000100000",
  52026=>"000000101",
  52027=>"000000001",
  52028=>"110011011",
  52029=>"110111010",
  52030=>"000101001",
  52031=>"000110110",
  52032=>"111111111",
  52033=>"001001111",
  52034=>"111111000",
  52035=>"011111011",
  52036=>"000010111",
  52037=>"000000100",
  52038=>"100101111",
  52039=>"000110110",
  52040=>"111111111",
  52041=>"001110010",
  52042=>"010000001",
  52043=>"111010111",
  52044=>"000110111",
  52045=>"011001110",
  52046=>"000000001",
  52047=>"011101111",
  52048=>"111111110",
  52049=>"110111000",
  52050=>"111101111",
  52051=>"001100000",
  52052=>"001101000",
  52053=>"011011111",
  52054=>"011001001",
  52055=>"001001111",
  52056=>"110111000",
  52057=>"011011110",
  52058=>"111011010",
  52059=>"100100000",
  52060=>"000000000",
  52061=>"001001001",
  52062=>"010010000",
  52063=>"110111101",
  52064=>"101101000",
  52065=>"010010000",
  52066=>"001001101",
  52067=>"111111110",
  52068=>"000000110",
  52069=>"100000110",
  52070=>"010111110",
  52071=>"111111000",
  52072=>"011101111",
  52073=>"000001101",
  52074=>"111101011",
  52075=>"000000000",
  52076=>"010000000",
  52077=>"101101001",
  52078=>"111111100",
  52079=>"111000110",
  52080=>"001001100",
  52081=>"010000000",
  52082=>"110000000",
  52083=>"001000001",
  52084=>"111110010",
  52085=>"000000000",
  52086=>"010000100",
  52087=>"001010000",
  52088=>"110110000",
  52089=>"000101000",
  52090=>"000111110",
  52091=>"000001001",
  52092=>"101010000",
  52093=>"100000000",
  52094=>"010100000",
  52095=>"001001111",
  52096=>"100001001",
  52097=>"100100100",
  52098=>"111000000",
  52099=>"111000000",
  52100=>"111001000",
  52101=>"111111111",
  52102=>"100100110",
  52103=>"000000100",
  52104=>"100110111",
  52105=>"000111101",
  52106=>"101100111",
  52107=>"000000000",
  52108=>"011000000",
  52109=>"111101111",
  52110=>"000000000",
  52111=>"000001000",
  52112=>"011001010",
  52113=>"111110000",
  52114=>"111001111",
  52115=>"000000010",
  52116=>"000000111",
  52117=>"000000111",
  52118=>"110111111",
  52119=>"110110000",
  52120=>"000000000",
  52121=>"001111100",
  52122=>"000010111",
  52123=>"000000011",
  52124=>"000000011",
  52125=>"000000100",
  52126=>"111111111",
  52127=>"000100101",
  52128=>"110111111",
  52129=>"001000101",
  52130=>"010001101",
  52131=>"111111111",
  52132=>"010111000",
  52133=>"111111111",
  52134=>"111111000",
  52135=>"100101000",
  52136=>"000000000",
  52137=>"000001001",
  52138=>"001001001",
  52139=>"000000110",
  52140=>"001101111",
  52141=>"011111111",
  52142=>"100101111",
  52143=>"111111011",
  52144=>"000000000",
  52145=>"011101001",
  52146=>"001001001",
  52147=>"011001000",
  52148=>"111111011",
  52149=>"111111110",
  52150=>"111010000",
  52151=>"110110000",
  52152=>"111111110",
  52153=>"110010000",
  52154=>"111010000",
  52155=>"110000010",
  52156=>"000001001",
  52157=>"111111101",
  52158=>"101011111",
  52159=>"000000111",
  52160=>"111110111",
  52161=>"001111100",
  52162=>"111110110",
  52163=>"000000110",
  52164=>"000000111",
  52165=>"000111011",
  52166=>"111000111",
  52167=>"111100101",
  52168=>"100000000",
  52169=>"110110111",
  52170=>"000000010",
  52171=>"001000011",
  52172=>"110110000",
  52173=>"011101001",
  52174=>"101001000",
  52175=>"111001000",
  52176=>"111110111",
  52177=>"111101111",
  52178=>"000000110",
  52179=>"101101000",
  52180=>"001000000",
  52181=>"001001001",
  52182=>"000001001",
  52183=>"001111111",
  52184=>"000000000",
  52185=>"111111111",
  52186=>"110110111",
  52187=>"001000101",
  52188=>"110100001",
  52189=>"000110010",
  52190=>"111110110",
  52191=>"010000010",
  52192=>"011110000",
  52193=>"000011011",
  52194=>"000000000",
  52195=>"001101110",
  52196=>"101101001",
  52197=>"000001001",
  52198=>"000000000",
  52199=>"011101110",
  52200=>"111101100",
  52201=>"011001000",
  52202=>"001101001",
  52203=>"001001001",
  52204=>"010010000",
  52205=>"000000001",
  52206=>"110100000",
  52207=>"001100110",
  52208=>"000000010",
  52209=>"010100100",
  52210=>"110111000",
  52211=>"111111110",
  52212=>"110100111",
  52213=>"101010010",
  52214=>"001000010",
  52215=>"111000010",
  52216=>"000000111",
  52217=>"000110111",
  52218=>"111111110",
  52219=>"000010110",
  52220=>"011111000",
  52221=>"111101111",
  52222=>"100100110",
  52223=>"000001000",
  52224=>"110000111",
  52225=>"110111110",
  52226=>"101001100",
  52227=>"000000001",
  52228=>"111111111",
  52229=>"111001101",
  52230=>"000110000",
  52231=>"100111111",
  52232=>"000000111",
  52233=>"100001000",
  52234=>"011011010",
  52235=>"000000001",
  52236=>"001001111",
  52237=>"101101001",
  52238=>"100000000",
  52239=>"111111011",
  52240=>"111001001",
  52241=>"111001111",
  52242=>"111101000",
  52243=>"000011001",
  52244=>"000110110",
  52245=>"011010011",
  52246=>"111111010",
  52247=>"010110001",
  52248=>"111000000",
  52249=>"000001111",
  52250=>"111111111",
  52251=>"000000110",
  52252=>"101000010",
  52253=>"111111111",
  52254=>"111010000",
  52255=>"000000000",
  52256=>"001001001",
  52257=>"100111010",
  52258=>"000000000",
  52259=>"110001101",
  52260=>"100110000",
  52261=>"000001111",
  52262=>"000000100",
  52263=>"010000000",
  52264=>"111111111",
  52265=>"000001000",
  52266=>"101001000",
  52267=>"110011110",
  52268=>"000010100",
  52269=>"111111111",
  52270=>"111001011",
  52271=>"011000001",
  52272=>"111111011",
  52273=>"000110100",
  52274=>"001111000",
  52275=>"110111000",
  52276=>"010001111",
  52277=>"100100000",
  52278=>"001000000",
  52279=>"000110010",
  52280=>"110000001",
  52281=>"000010000",
  52282=>"010001111",
  52283=>"010110000",
  52284=>"000001110",
  52285=>"111110100",
  52286=>"000001001",
  52287=>"000001001",
  52288=>"000000111",
  52289=>"111100001",
  52290=>"000101000",
  52291=>"001001000",
  52292=>"000010000",
  52293=>"000111110",
  52294=>"101010000",
  52295=>"110110101",
  52296=>"101111111",
  52297=>"000000000",
  52298=>"001100101",
  52299=>"000010110",
  52300=>"001001111",
  52301=>"011011001",
  52302=>"000110011",
  52303=>"000110000",
  52304=>"110000001",
  52305=>"111111101",
  52306=>"011010000",
  52307=>"010010001",
  52308=>"000000011",
  52309=>"110110000",
  52310=>"000100110",
  52311=>"111100110",
  52312=>"110011001",
  52313=>"001111000",
  52314=>"000100111",
  52315=>"000010110",
  52316=>"000000000",
  52317=>"000000110",
  52318=>"011111000",
  52319=>"000000101",
  52320=>"111000000",
  52321=>"000001111",
  52322=>"101001111",
  52323=>"111001001",
  52324=>"000000000",
  52325=>"000010011",
  52326=>"000101101",
  52327=>"000000110",
  52328=>"000000000",
  52329=>"001001000",
  52330=>"100001001",
  52331=>"010000000",
  52332=>"001000110",
  52333=>"001101111",
  52334=>"101111000",
  52335=>"110111011",
  52336=>"001010011",
  52337=>"111110000",
  52338=>"100000001",
  52339=>"000111000",
  52340=>"110101111",
  52341=>"100111011",
  52342=>"000000000",
  52343=>"000000000",
  52344=>"101111111",
  52345=>"000010010",
  52346=>"110101001",
  52347=>"001111001",
  52348=>"010000001",
  52349=>"100101100",
  52350=>"010011000",
  52351=>"000000111",
  52352=>"110011011",
  52353=>"111001000",
  52354=>"000010010",
  52355=>"000110100",
  52356=>"011000000",
  52357=>"000000000",
  52358=>"100000110",
  52359=>"000001011",
  52360=>"100111110",
  52361=>"000000000",
  52362=>"101101100",
  52363=>"001000001",
  52364=>"000001011",
  52365=>"101111111",
  52366=>"000010000",
  52367=>"001001100",
  52368=>"000001000",
  52369=>"001111110",
  52370=>"000001000",
  52371=>"110110000",
  52372=>"000110110",
  52373=>"101001000",
  52374=>"111111011",
  52375=>"100100000",
  52376=>"000101110",
  52377=>"111110111",
  52378=>"000101010",
  52379=>"111001000",
  52380=>"000001101",
  52381=>"001000010",
  52382=>"000000011",
  52383=>"010100110",
  52384=>"011011110",
  52385=>"110010111",
  52386=>"000001110",
  52387=>"000010111",
  52388=>"111000011",
  52389=>"100100010",
  52390=>"000000010",
  52391=>"000011000",
  52392=>"111110110",
  52393=>"000000000",
  52394=>"111001111",
  52395=>"110011111",
  52396=>"001111111",
  52397=>"100000110",
  52398=>"101010110",
  52399=>"000000111",
  52400=>"111111110",
  52401=>"000010001",
  52402=>"111111111",
  52403=>"010001000",
  52404=>"101100000",
  52405=>"110110000",
  52406=>"111101101",
  52407=>"000000110",
  52408=>"000100110",
  52409=>"001111010",
  52410=>"000000000",
  52411=>"000000011",
  52412=>"101000110",
  52413=>"111001111",
  52414=>"111010010",
  52415=>"000001001",
  52416=>"110110010",
  52417=>"000001110",
  52418=>"111110001",
  52419=>"100100010",
  52420=>"000000111",
  52421=>"110110111",
  52422=>"000001110",
  52423=>"001000111",
  52424=>"101111000",
  52425=>"101001111",
  52426=>"111001011",
  52427=>"000100001",
  52428=>"000000000",
  52429=>"100000001",
  52430=>"110100111",
  52431=>"010001111",
  52432=>"101101001",
  52433=>"010111111",
  52434=>"000000111",
  52435=>"001010111",
  52436=>"111101111",
  52437=>"100100111",
  52438=>"001000000",
  52439=>"111110000",
  52440=>"000110111",
  52441=>"111111101",
  52442=>"100110110",
  52443=>"101001111",
  52444=>"110111001",
  52445=>"001001001",
  52446=>"010111111",
  52447=>"000001111",
  52448=>"001001111",
  52449=>"111000011",
  52450=>"011111111",
  52451=>"100110111",
  52452=>"000000001",
  52453=>"000100010",
  52454=>"101111000",
  52455=>"000100110",
  52456=>"011001111",
  52457=>"000110111",
  52458=>"101110111",
  52459=>"111001001",
  52460=>"001001101",
  52461=>"000001011",
  52462=>"111101110",
  52463=>"111110100",
  52464=>"000111110",
  52465=>"011111110",
  52466=>"001011010",
  52467=>"000000000",
  52468=>"000010010",
  52469=>"101001000",
  52470=>"001001111",
  52471=>"010000111",
  52472=>"110000000",
  52473=>"000000000",
  52474=>"010111111",
  52475=>"100110100",
  52476=>"111111001",
  52477=>"101111111",
  52478=>"100111111",
  52479=>"000000000",
  52480=>"000010110",
  52481=>"111111001",
  52482=>"000000111",
  52483=>"111010000",
  52484=>"010000011",
  52485=>"101101111",
  52486=>"111000000",
  52487=>"011110000",
  52488=>"000000011",
  52489=>"000111000",
  52490=>"111101000",
  52491=>"111111111",
  52492=>"000000111",
  52493=>"000000111",
  52494=>"100000100",
  52495=>"010111111",
  52496=>"111101000",
  52497=>"000000111",
  52498=>"000010111",
  52499=>"101100000",
  52500=>"000000011",
  52501=>"111101100",
  52502=>"111110001",
  52503=>"010111110",
  52504=>"000100110",
  52505=>"111111101",
  52506=>"010001010",
  52507=>"111000000",
  52508=>"001100000",
  52509=>"101111101",
  52510=>"000011000",
  52511=>"000000101",
  52512=>"110000111",
  52513=>"111000000",
  52514=>"000000111",
  52515=>"000010000",
  52516=>"011010110",
  52517=>"000000000",
  52518=>"111100010",
  52519=>"010010111",
  52520=>"011011100",
  52521=>"010000001",
  52522=>"111011000",
  52523=>"111111010",
  52524=>"011000000",
  52525=>"111110010",
  52526=>"111111101",
  52527=>"000000100",
  52528=>"111011111",
  52529=>"110110011",
  52530=>"010111111",
  52531=>"111001110",
  52532=>"101000000",
  52533=>"000000000",
  52534=>"101100000",
  52535=>"100100000",
  52536=>"110000000",
  52537=>"000101101",
  52538=>"000000111",
  52539=>"001010010",
  52540=>"011001100",
  52541=>"011000000",
  52542=>"001001111",
  52543=>"101000000",
  52544=>"010111111",
  52545=>"000111000",
  52546=>"110010101",
  52547=>"000000000",
  52548=>"111111000",
  52549=>"001101001",
  52550=>"110110000",
  52551=>"001000111",
  52552=>"110111110",
  52553=>"111110010",
  52554=>"001101000",
  52555=>"111100000",
  52556=>"000000111",
  52557=>"110000111",
  52558=>"110001100",
  52559=>"110000100",
  52560=>"000101101",
  52561=>"111000000",
  52562=>"010101111",
  52563=>"001010010",
  52564=>"000000000",
  52565=>"111100001",
  52566=>"110010000",
  52567=>"111000000",
  52568=>"011001111",
  52569=>"011010111",
  52570=>"100100111",
  52571=>"111110111",
  52572=>"111000000",
  52573=>"001110110",
  52574=>"000111111",
  52575=>"001010000",
  52576=>"110010111",
  52577=>"111111000",
  52578=>"000111111",
  52579=>"011011001",
  52580=>"110001011",
  52581=>"000000100",
  52582=>"000010101",
  52583=>"100001001",
  52584=>"110000010",
  52585=>"000000011",
  52586=>"000111111",
  52587=>"000101111",
  52588=>"111000000",
  52589=>"000000111",
  52590=>"111000000",
  52591=>"010000000",
  52592=>"111110110",
  52593=>"111010000",
  52594=>"000010000",
  52595=>"001000111",
  52596=>"100000000",
  52597=>"000111101",
  52598=>"111010011",
  52599=>"000001000",
  52600=>"101010010",
  52601=>"011111111",
  52602=>"001110000",
  52603=>"000011111",
  52604=>"010001000",
  52605=>"000010011",
  52606=>"100000000",
  52607=>"000101100",
  52608=>"111000000",
  52609=>"101001010",
  52610=>"111110000",
  52611=>"111111100",
  52612=>"000101101",
  52613=>"000111001",
  52614=>"010000000",
  52615=>"111010000",
  52616=>"011010000",
  52617=>"000111001",
  52618=>"011011110",
  52619=>"000011111",
  52620=>"100101001",
  52621=>"111000100",
  52622=>"100000000",
  52623=>"001001001",
  52624=>"000011110",
  52625=>"000000000",
  52626=>"000000000",
  52627=>"101001011",
  52628=>"111100000",
  52629=>"101011011",
  52630=>"110100101",
  52631=>"111110110",
  52632=>"010111100",
  52633=>"111001000",
  52634=>"100000111",
  52635=>"100000000",
  52636=>"011000000",
  52637=>"100000000",
  52638=>"111010000",
  52639=>"110000110",
  52640=>"001010110",
  52641=>"010011111",
  52642=>"111010111",
  52643=>"111111000",
  52644=>"000011111",
  52645=>"110011000",
  52646=>"001011111",
  52647=>"101000000",
  52648=>"111101000",
  52649=>"111000000",
  52650=>"100010110",
  52651=>"000000000",
  52652=>"000000111",
  52653=>"111110010",
  52654=>"000000011",
  52655=>"111111000",
  52656=>"101111011",
  52657=>"110110111",
  52658=>"100110000",
  52659=>"110000010",
  52660=>"110110111",
  52661=>"111010011",
  52662=>"101011101",
  52663=>"010111111",
  52664=>"110000100",
  52665=>"111011000",
  52666=>"011100000",
  52667=>"011010000",
  52668=>"000101111",
  52669=>"000100111",
  52670=>"110000000",
  52671=>"000000000",
  52672=>"011011000",
  52673=>"010000000",
  52674=>"000000000",
  52675=>"000000000",
  52676=>"001101111",
  52677=>"100100100",
  52678=>"111011011",
  52679=>"000111111",
  52680=>"101110111",
  52681=>"001101111",
  52682=>"111100000",
  52683=>"100100111",
  52684=>"101010100",
  52685=>"111100000",
  52686=>"010001100",
  52687=>"000000111",
  52688=>"001100111",
  52689=>"001000000",
  52690=>"111111001",
  52691=>"011010110",
  52692=>"100110000",
  52693=>"111001001",
  52694=>"111000110",
  52695=>"111000000",
  52696=>"111111011",
  52697=>"100000000",
  52698=>"110010110",
  52699=>"000101111",
  52700=>"111111000",
  52701=>"000000111",
  52702=>"111001101",
  52703=>"111111000",
  52704=>"000000010",
  52705=>"001011001",
  52706=>"000111111",
  52707=>"000100011",
  52708=>"101000000",
  52709=>"100001100",
  52710=>"110000010",
  52711=>"110100100",
  52712=>"010011010",
  52713=>"101101111",
  52714=>"000000000",
  52715=>"000011011",
  52716=>"000001011",
  52717=>"000100100",
  52718=>"101000000",
  52719=>"111000000",
  52720=>"000000100",
  52721=>"001000011",
  52722=>"110010101",
  52723=>"010011110",
  52724=>"011011011",
  52725=>"100111101",
  52726=>"000000111",
  52727=>"111111111",
  52728=>"010010000",
  52729=>"010000111",
  52730=>"011001100",
  52731=>"111110110",
  52732=>"111100000",
  52733=>"111111011",
  52734=>"000000110",
  52735=>"110110000",
  52736=>"100111011",
  52737=>"110011101",
  52738=>"001000111",
  52739=>"010010001",
  52740=>"100010000",
  52741=>"000000101",
  52742=>"001110000",
  52743=>"000101101",
  52744=>"100001111",
  52745=>"111100111",
  52746=>"000000001",
  52747=>"101101101",
  52748=>"110110010",
  52749=>"000100110",
  52750=>"010110000",
  52751=>"000000111",
  52752=>"001110101",
  52753=>"100000000",
  52754=>"111111010",
  52755=>"011111001",
  52756=>"111111111",
  52757=>"011001101",
  52758=>"010111011",
  52759=>"000000001",
  52760=>"000100111",
  52761=>"111100110",
  52762=>"000000111",
  52763=>"000000010",
  52764=>"100111001",
  52765=>"101101010",
  52766=>"110111101",
  52767=>"100000000",
  52768=>"100000111",
  52769=>"000000011",
  52770=>"111011000",
  52771=>"101000100",
  52772=>"110110100",
  52773=>"011000000",
  52774=>"100000010",
  52775=>"000000000",
  52776=>"000111011",
  52777=>"101000000",
  52778=>"111100111",
  52779=>"101111100",
  52780=>"111011110",
  52781=>"011111011",
  52782=>"100111101",
  52783=>"000000101",
  52784=>"000000000",
  52785=>"110110111",
  52786=>"011101110",
  52787=>"111100000",
  52788=>"000000000",
  52789=>"111010000",
  52790=>"000000010",
  52791=>"000110010",
  52792=>"000111111",
  52793=>"000110000",
  52794=>"110101101",
  52795=>"000000000",
  52796=>"000110000",
  52797=>"111010101",
  52798=>"100000010",
  52799=>"000011111",
  52800=>"111111000",
  52801=>"000110000",
  52802=>"101101101",
  52803=>"000110111",
  52804=>"111111011",
  52805=>"001010101",
  52806=>"000011111",
  52807=>"111111011",
  52808=>"011111111",
  52809=>"111111000",
  52810=>"000100101",
  52811=>"110111101",
  52812=>"011100111",
  52813=>"111111010",
  52814=>"100010001",
  52815=>"111111111",
  52816=>"100010010",
  52817=>"111111110",
  52818=>"111111100",
  52819=>"111011001",
  52820=>"111111010",
  52821=>"010011001",
  52822=>"100111111",
  52823=>"111101111",
  52824=>"001000110",
  52825=>"010010000",
  52826=>"011000000",
  52827=>"100110011",
  52828=>"000010000",
  52829=>"010011000",
  52830=>"010111110",
  52831=>"011011010",
  52832=>"010000001",
  52833=>"010110000",
  52834=>"011100111",
  52835=>"011011000",
  52836=>"101110000",
  52837=>"011001001",
  52838=>"000110111",
  52839=>"100101111",
  52840=>"111000010",
  52841=>"001100000",
  52842=>"100111111",
  52843=>"101011000",
  52844=>"100111101",
  52845=>"111000111",
  52846=>"000000000",
  52847=>"000000111",
  52848=>"011011011",
  52849=>"000000101",
  52850=>"000000000",
  52851=>"111101111",
  52852=>"100100110",
  52853=>"000000101",
  52854=>"000000000",
  52855=>"010000111",
  52856=>"110000111",
  52857=>"110000111",
  52858=>"111011101",
  52859=>"000000000",
  52860=>"110011001",
  52861=>"111110100",
  52862=>"000000111",
  52863=>"110000000",
  52864=>"000101111",
  52865=>"011111100",
  52866=>"000010111",
  52867=>"001100000",
  52868=>"111011010",
  52869=>"001001111",
  52870=>"100100101",
  52871=>"100100100",
  52872=>"111111000",
  52873=>"000000001",
  52874=>"000000010",
  52875=>"010101111",
  52876=>"001000010",
  52877=>"000101011",
  52878=>"000011000",
  52879=>"001001111",
  52880=>"111011111",
  52881=>"000000000",
  52882=>"000000000",
  52883=>"100110000",
  52884=>"000011100",
  52885=>"000101110",
  52886=>"111111100",
  52887=>"001110100",
  52888=>"100000011",
  52889=>"011000001",
  52890=>"001100111",
  52891=>"111100101",
  52892=>"011011111",
  52893=>"000100000",
  52894=>"111010010",
  52895=>"111110110",
  52896=>"001010011",
  52897=>"011011111",
  52898=>"000000101",
  52899=>"111111111",
  52900=>"111110000",
  52901=>"001000010",
  52902=>"011011000",
  52903=>"110111001",
  52904=>"000111101",
  52905=>"010011000",
  52906=>"101101111",
  52907=>"110111011",
  52908=>"111101100",
  52909=>"010110011",
  52910=>"011111000",
  52911=>"111000001",
  52912=>"110100101",
  52913=>"100111000",
  52914=>"111011000",
  52915=>"110001001",
  52916=>"000110000",
  52917=>"111111111",
  52918=>"111110000",
  52919=>"110000111",
  52920=>"010011010",
  52921=>"100011001",
  52922=>"000010011",
  52923=>"101111010",
  52924=>"000011010",
  52925=>"111101111",
  52926=>"111111111",
  52927=>"100000000",
  52928=>"010111010",
  52929=>"110011001",
  52930=>"111111000",
  52931=>"100110011",
  52932=>"111001111",
  52933=>"111111111",
  52934=>"000100111",
  52935=>"011000100",
  52936=>"100000100",
  52937=>"010100010",
  52938=>"101000111",
  52939=>"000000111",
  52940=>"000000000",
  52941=>"011110110",
  52942=>"010000011",
  52943=>"111111110",
  52944=>"010111111",
  52945=>"110110111",
  52946=>"100011101",
  52947=>"000010010",
  52948=>"000111011",
  52949=>"100000000",
  52950=>"010111010",
  52951=>"011110000",
  52952=>"001000000",
  52953=>"000011001",
  52954=>"111110100",
  52955=>"111100101",
  52956=>"110110110",
  52957=>"010100111",
  52958=>"110000010",
  52959=>"000010111",
  52960=>"000100111",
  52961=>"111010010",
  52962=>"010000001",
  52963=>"111011001",
  52964=>"000000000",
  52965=>"101100111",
  52966=>"000000101",
  52967=>"100110010",
  52968=>"101100111",
  52969=>"101100011",
  52970=>"001000000",
  52971=>"000000101",
  52972=>"000000111",
  52973=>"111000000",
  52974=>"110111111",
  52975=>"000101111",
  52976=>"101001111",
  52977=>"111111011",
  52978=>"010111001",
  52979=>"010001000",
  52980=>"001011110",
  52981=>"100100001",
  52982=>"111100001",
  52983=>"110100001",
  52984=>"010011000",
  52985=>"000000111",
  52986=>"100011110",
  52987=>"100110010",
  52988=>"011011111",
  52989=>"101000111",
  52990=>"110110010",
  52991=>"000111100",
  52992=>"011001010",
  52993=>"000000010",
  52994=>"000010000",
  52995=>"111000110",
  52996=>"000000111",
  52997=>"110101100",
  52998=>"000000100",
  52999=>"111101110",
  53000=>"011011000",
  53001=>"000000101",
  53002=>"000111110",
  53003=>"000011010",
  53004=>"000111010",
  53005=>"111111100",
  53006=>"000011011",
  53007=>"001101100",
  53008=>"111101111",
  53009=>"000111111",
  53010=>"111000000",
  53011=>"000000111",
  53012=>"110010100",
  53013=>"010010000",
  53014=>"011001100",
  53015=>"011010010",
  53016=>"000000011",
  53017=>"000101110",
  53018=>"010000000",
  53019=>"000111111",
  53020=>"111001111",
  53021=>"110100111",
  53022=>"111101000",
  53023=>"100101001",
  53024=>"000101111",
  53025=>"000111000",
  53026=>"000010110",
  53027=>"001001011",
  53028=>"111101100",
  53029=>"001001011",
  53030=>"111000001",
  53031=>"000000100",
  53032=>"110110000",
  53033=>"100000001",
  53034=>"101000100",
  53035=>"000000000",
  53036=>"100001011",
  53037=>"111010000",
  53038=>"111111001",
  53039=>"111111001",
  53040=>"000000000",
  53041=>"001001011",
  53042=>"101001101",
  53043=>"111000000",
  53044=>"000111111",
  53045=>"000010001",
  53046=>"111111111",
  53047=>"111001001",
  53048=>"111101011",
  53049=>"110110000",
  53050=>"000101000",
  53051=>"000111100",
  53052=>"101011011",
  53053=>"111111111",
  53054=>"110000000",
  53055=>"110011111",
  53056=>"010110111",
  53057=>"000000111",
  53058=>"001001000",
  53059=>"011011001",
  53060=>"111000011",
  53061=>"110010000",
  53062=>"000111110",
  53063=>"111111000",
  53064=>"110111100",
  53065=>"111111111",
  53066=>"111001101",
  53067=>"100111111",
  53068=>"001000011",
  53069=>"000011011",
  53070=>"111111100",
  53071=>"000010111",
  53072=>"100100111",
  53073=>"111000000",
  53074=>"111111000",
  53075=>"111000111",
  53076=>"111111111",
  53077=>"111010111",
  53078=>"000001001",
  53079=>"111111111",
  53080=>"000010110",
  53081=>"111001001",
  53082=>"000100011",
  53083=>"000111011",
  53084=>"110110111",
  53085=>"001001001",
  53086=>"000010111",
  53087=>"111100100",
  53088=>"001010011",
  53089=>"010100111",
  53090=>"010011110",
  53091=>"101001111",
  53092=>"110101110",
  53093=>"000001001",
  53094=>"000111110",
  53095=>"111000000",
  53096=>"000110111",
  53097=>"000000000",
  53098=>"111011000",
  53099=>"111000010",
  53100=>"111000000",
  53101=>"000001110",
  53102=>"111111110",
  53103=>"000000110",
  53104=>"100100000",
  53105=>"000001001",
  53106=>"011111110",
  53107=>"000000011",
  53108=>"111000000",
  53109=>"101000000",
  53110=>"000000100",
  53111=>"100110110",
  53112=>"111010110",
  53113=>"010000110",
  53114=>"000000000",
  53115=>"010111111",
  53116=>"011001101",
  53117=>"110100000",
  53118=>"110111101",
  53119=>"110111101",
  53120=>"110110001",
  53121=>"111101100",
  53122=>"001111001",
  53123=>"000000010",
  53124=>"111111000",
  53125=>"001111010",
  53126=>"000000111",
  53127=>"100100100",
  53128=>"111011011",
  53129=>"100111111",
  53130=>"110111111",
  53131=>"010000010",
  53132=>"000111111",
  53133=>"000111111",
  53134=>"110101111",
  53135=>"000001001",
  53136=>"101100100",
  53137=>"000000110",
  53138=>"111111101",
  53139=>"111000000",
  53140=>"111101001",
  53141=>"111101101",
  53142=>"000010010",
  53143=>"110100000",
  53144=>"000000010",
  53145=>"011000010",
  53146=>"000010111",
  53147=>"111111111",
  53148=>"000001111",
  53149=>"000000111",
  53150=>"000000111",
  53151=>"111000000",
  53152=>"000111100",
  53153=>"111111000",
  53154=>"111101100",
  53155=>"000000111",
  53156=>"111000000",
  53157=>"000010000",
  53158=>"111111001",
  53159=>"000000111",
  53160=>"111111111",
  53161=>"100100000",
  53162=>"111011000",
  53163=>"000000010",
  53164=>"101111100",
  53165=>"111001000",
  53166=>"100101011",
  53167=>"110110110",
  53168=>"001000010",
  53169=>"011011001",
  53170=>"101001101",
  53171=>"000001100",
  53172=>"010110110",
  53173=>"111111101",
  53174=>"000111111",
  53175=>"000000100",
  53176=>"100100100",
  53177=>"111001101",
  53178=>"000000010",
  53179=>"001001111",
  53180=>"000110110",
  53181=>"110000011",
  53182=>"111111110",
  53183=>"111101101",
  53184=>"010110111",
  53185=>"000110111",
  53186=>"101111111",
  53187=>"111111000",
  53188=>"100111000",
  53189=>"110110010",
  53190=>"111110000",
  53191=>"011011000",
  53192=>"000011010",
  53193=>"100110000",
  53194=>"111101100",
  53195=>"000111111",
  53196=>"000000111",
  53197=>"110100001",
  53198=>"000010000",
  53199=>"010001000",
  53200=>"000010010",
  53201=>"001011011",
  53202=>"010111000",
  53203=>"101100000",
  53204=>"110111110",
  53205=>"000000100",
  53206=>"111111110",
  53207=>"111111010",
  53208=>"000000110",
  53209=>"110010011",
  53210=>"001100100",
  53211=>"000000010",
  53212=>"111111011",
  53213=>"011110111",
  53214=>"010111111",
  53215=>"111110010",
  53216=>"001110111",
  53217=>"000000000",
  53218=>"010011010",
  53219=>"100100111",
  53220=>"010111111",
  53221=>"000111000",
  53222=>"110000000",
  53223=>"110101101",
  53224=>"010010000",
  53225=>"101000110",
  53226=>"010110111",
  53227=>"001111111",
  53228=>"000000101",
  53229=>"101001000",
  53230=>"011010000",
  53231=>"011000000",
  53232=>"111111010",
  53233=>"011011010",
  53234=>"111001001",
  53235=>"110101101",
  53236=>"110110101",
  53237=>"000000000",
  53238=>"000000111",
  53239=>"000000111",
  53240=>"010010000",
  53241=>"111101000",
  53242=>"111111111",
  53243=>"111111010",
  53244=>"111111111",
  53245=>"010110111",
  53246=>"110100111",
  53247=>"101001000",
  53248=>"110100100",
  53249=>"000111111",
  53250=>"011000111",
  53251=>"000111111",
  53252=>"000111000",
  53253=>"000000011",
  53254=>"111111100",
  53255=>"011011111",
  53256=>"000100001",
  53257=>"010000111",
  53258=>"111000100",
  53259=>"000000000",
  53260=>"101111010",
  53261=>"000000011",
  53262=>"001011100",
  53263=>"101000001",
  53264=>"000100000",
  53265=>"111000000",
  53266=>"110000010",
  53267=>"111100001",
  53268=>"000001111",
  53269=>"111111000",
  53270=>"000111001",
  53271=>"000111110",
  53272=>"000000101",
  53273=>"000111111",
  53274=>"100100000",
  53275=>"110000111",
  53276=>"000100000",
  53277=>"001000000",
  53278=>"101001011",
  53279=>"111000000",
  53280=>"000000000",
  53281=>"000100110",
  53282=>"111000100",
  53283=>"100111000",
  53284=>"010010000",
  53285=>"011011011",
  53286=>"100110000",
  53287=>"101000000",
  53288=>"110111111",
  53289=>"000010000",
  53290=>"000000000",
  53291=>"111000000",
  53292=>"111111011",
  53293=>"111111000",
  53294=>"101100111",
  53295=>"000000011",
  53296=>"100001000",
  53297=>"110011010",
  53298=>"000000101",
  53299=>"000000111",
  53300=>"111000101",
  53301=>"111001000",
  53302=>"011011111",
  53303=>"010011000",
  53304=>"101010111",
  53305=>"000000111",
  53306=>"000101010",
  53307=>"000101111",
  53308=>"011011011",
  53309=>"010011011",
  53310=>"010000101",
  53311=>"011011001",
  53312=>"101000111",
  53313=>"001001011",
  53314=>"101001111",
  53315=>"011100010",
  53316=>"001000010",
  53317=>"101101101",
  53318=>"111111000",
  53319=>"000000011",
  53320=>"010111111",
  53321=>"101000110",
  53322=>"000000000",
  53323=>"111000000",
  53324=>"101000111",
  53325=>"011111111",
  53326=>"000110111",
  53327=>"111000000",
  53328=>"000001000",
  53329=>"011111111",
  53330=>"101111001",
  53331=>"001100000",
  53332=>"000000000",
  53333=>"100110100",
  53334=>"111010000",
  53335=>"000000100",
  53336=>"000111111",
  53337=>"000011110",
  53338=>"011000000",
  53339=>"000100011",
  53340=>"001000101",
  53341=>"000100110",
  53342=>"111111000",
  53343=>"000001011",
  53344=>"000001111",
  53345=>"111101100",
  53346=>"001000111",
  53347=>"100101110",
  53348=>"100000011",
  53349=>"000000100",
  53350=>"001001110",
  53351=>"110110001",
  53352=>"001110111",
  53353=>"111011111",
  53354=>"110011000",
  53355=>"000101001",
  53356=>"001000111",
  53357=>"111110010",
  53358=>"001001001",
  53359=>"010111111",
  53360=>"001011010",
  53361=>"000110110",
  53362=>"100100100",
  53363=>"010111001",
  53364=>"000011000",
  53365=>"100100101",
  53366=>"101010111",
  53367=>"111001001",
  53368=>"010000111",
  53369=>"111011010",
  53370=>"110111101",
  53371=>"100111110",
  53372=>"111011001",
  53373=>"100011010",
  53374=>"111011101",
  53375=>"110010001",
  53376=>"001001000",
  53377=>"000110101",
  53378=>"000000111",
  53379=>"011110000",
  53380=>"111111000",
  53381=>"110000000",
  53382=>"100101111",
  53383=>"000011001",
  53384=>"010110000",
  53385=>"000001000",
  53386=>"111111000",
  53387=>"001000111",
  53388=>"010110101",
  53389=>"001000001",
  53390=>"000000000",
  53391=>"101000000",
  53392=>"000111011",
  53393=>"111110000",
  53394=>"010000111",
  53395=>"000010111",
  53396=>"100111000",
  53397=>"001000111",
  53398=>"101101111",
  53399=>"001110110",
  53400=>"110010000",
  53401=>"000000110",
  53402=>"000111000",
  53403=>"111000011",
  53404=>"111110011",
  53405=>"001000111",
  53406=>"001111000",
  53407=>"111001111",
  53408=>"011111011",
  53409=>"111010111",
  53410=>"111111110",
  53411=>"000000000",
  53412=>"111110001",
  53413=>"110011001",
  53414=>"111111111",
  53415=>"001111111",
  53416=>"011111000",
  53417=>"000100001",
  53418=>"000000000",
  53419=>"000000100",
  53420=>"011000011",
  53421=>"000000000",
  53422=>"110100100",
  53423=>"111111000",
  53424=>"101000000",
  53425=>"000100100",
  53426=>"101001111",
  53427=>"100111011",
  53428=>"111010010",
  53429=>"101100111",
  53430=>"111010100",
  53431=>"001101001",
  53432=>"110110100",
  53433=>"111111100",
  53434=>"100101000",
  53435=>"100000000",
  53436=>"111000000",
  53437=>"000011001",
  53438=>"001010100",
  53439=>"000101000",
  53440=>"101000000",
  53441=>"010000000",
  53442=>"000000000",
  53443=>"111110100",
  53444=>"110000000",
  53445=>"010000001",
  53446=>"111110000",
  53447=>"110111000",
  53448=>"110000111",
  53449=>"110000001",
  53450=>"000000100",
  53451=>"111001111",
  53452=>"001001010",
  53453=>"000111101",
  53454=>"111000101",
  53455=>"110000000",
  53456=>"011011000",
  53457=>"111011000",
  53458=>"111010111",
  53459=>"111000000",
  53460=>"000000000",
  53461=>"000000001",
  53462=>"001000000",
  53463=>"000001000",
  53464=>"111111000",
  53465=>"111011100",
  53466=>"100001111",
  53467=>"011000000",
  53468=>"001011111",
  53469=>"111111111",
  53470=>"101101101",
  53471=>"001101010",
  53472=>"010000001",
  53473=>"001000111",
  53474=>"111110000",
  53475=>"100100000",
  53476=>"101001000",
  53477=>"011000000",
  53478=>"001011111",
  53479=>"111111011",
  53480=>"000000110",
  53481=>"001000111",
  53482=>"011001001",
  53483=>"101000001",
  53484=>"000000000",
  53485=>"000111101",
  53486=>"000100000",
  53487=>"000010000",
  53488=>"111000000",
  53489=>"100000110",
  53490=>"111101001",
  53491=>"100001010",
  53492=>"100001011",
  53493=>"010000000",
  53494=>"000101000",
  53495=>"111111100",
  53496=>"000111111",
  53497=>"111011100",
  53498=>"000011000",
  53499=>"001000001",
  53500=>"110001000",
  53501=>"001000000",
  53502=>"110000000",
  53503=>"000000110",
  53504=>"010000000",
  53505=>"000000001",
  53506=>"000000101",
  53507=>"001000000",
  53508=>"101001111",
  53509=>"000100010",
  53510=>"101000011",
  53511=>"100001111",
  53512=>"101100111",
  53513=>"101001001",
  53514=>"001001011",
  53515=>"010010111",
  53516=>"000000010",
  53517=>"010000000",
  53518=>"001111110",
  53519=>"111011010",
  53520=>"010110111",
  53521=>"000111101",
  53522=>"101001010",
  53523=>"000011011",
  53524=>"111111010",
  53525=>"000000010",
  53526=>"010110110",
  53527=>"001111111",
  53528=>"101000000",
  53529=>"101100111",
  53530=>"001011111",
  53531=>"000010110",
  53532=>"010100000",
  53533=>"000000000",
  53534=>"001000000",
  53535=>"111111000",
  53536=>"010000101",
  53537=>"000000111",
  53538=>"101100100",
  53539=>"101011010",
  53540=>"010110011",
  53541=>"000000001",
  53542=>"001000000",
  53543=>"100101100",
  53544=>"110110110",
  53545=>"110111111",
  53546=>"010000000",
  53547=>"010000000",
  53548=>"001011011",
  53549=>"000000000",
  53550=>"000100001",
  53551=>"110110111",
  53552=>"001000000",
  53553=>"100110111",
  53554=>"000111111",
  53555=>"111010111",
  53556=>"000000000",
  53557=>"111111111",
  53558=>"011000000",
  53559=>"100000000",
  53560=>"000010111",
  53561=>"001011001",
  53562=>"111101000",
  53563=>"000101111",
  53564=>"000111111",
  53565=>"111110110",
  53566=>"000000001",
  53567=>"110110110",
  53568=>"001001101",
  53569=>"101011001",
  53570=>"111110000",
  53571=>"110111100",
  53572=>"111101010",
  53573=>"101101010",
  53574=>"011101111",
  53575=>"001011010",
  53576=>"001111111",
  53577=>"001000000",
  53578=>"101000000",
  53579=>"111111111",
  53580=>"000000000",
  53581=>"001001111",
  53582=>"011010111",
  53583=>"111011111",
  53584=>"110000000",
  53585=>"100111110",
  53586=>"001000000",
  53587=>"001001000",
  53588=>"000000000",
  53589=>"000111011",
  53590=>"011011011",
  53591=>"000000001",
  53592=>"010110000",
  53593=>"110011000",
  53594=>"111111000",
  53595=>"110100010",
  53596=>"000000111",
  53597=>"011001100",
  53598=>"101110100",
  53599=>"011000001",
  53600=>"111111000",
  53601=>"010011011",
  53602=>"100000100",
  53603=>"110110000",
  53604=>"000111111",
  53605=>"111100010",
  53606=>"110111110",
  53607=>"111100000",
  53608=>"011111000",
  53609=>"000111010",
  53610=>"000010111",
  53611=>"010011111",
  53612=>"101001111",
  53613=>"000010111",
  53614=>"101000101",
  53615=>"000001111",
  53616=>"011011011",
  53617=>"000010111",
  53618=>"110000000",
  53619=>"001000000",
  53620=>"111111111",
  53621=>"100001000",
  53622=>"011111010",
  53623=>"101111111",
  53624=>"001111100",
  53625=>"010111111",
  53626=>"110010000",
  53627=>"000001111",
  53628=>"101100111",
  53629=>"101101001",
  53630=>"111101101",
  53631=>"111100101",
  53632=>"001001001",
  53633=>"100000010",
  53634=>"110000111",
  53635=>"111111111",
  53636=>"100100000",
  53637=>"001000000",
  53638=>"001100100",
  53639=>"100011110",
  53640=>"111111110",
  53641=>"000000001",
  53642=>"111111000",
  53643=>"000000001",
  53644=>"001101000",
  53645=>"111100111",
  53646=>"000101100",
  53647=>"101001001",
  53648=>"100111000",
  53649=>"110111110",
  53650=>"000001101",
  53651=>"111010111",
  53652=>"001111111",
  53653=>"000101111",
  53654=>"111010110",
  53655=>"101100101",
  53656=>"110111000",
  53657=>"100100000",
  53658=>"010110010",
  53659=>"100011111",
  53660=>"011000000",
  53661=>"010000001",
  53662=>"001000101",
  53663=>"000000110",
  53664=>"000111110",
  53665=>"111111101",
  53666=>"101001000",
  53667=>"010111010",
  53668=>"000101010",
  53669=>"111001010",
  53670=>"000001101",
  53671=>"001111111",
  53672=>"000000000",
  53673=>"001011011",
  53674=>"000000000",
  53675=>"010001101",
  53676=>"001010111",
  53677=>"000000000",
  53678=>"011011001",
  53679=>"111010000",
  53680=>"000010111",
  53681=>"001110111",
  53682=>"101101111",
  53683=>"110110111",
  53684=>"111110010",
  53685=>"111101111",
  53686=>"000000000",
  53687=>"010110001",
  53688=>"000011011",
  53689=>"001011011",
  53690=>"000010000",
  53691=>"111111011",
  53692=>"001111000",
  53693=>"000110111",
  53694=>"011011011",
  53695=>"001000000",
  53696=>"000000101",
  53697=>"010110000",
  53698=>"010011000",
  53699=>"110010000",
  53700=>"000001101",
  53701=>"000000001",
  53702=>"011000100",
  53703=>"101000000",
  53704=>"000000010",
  53705=>"000100000",
  53706=>"001000001",
  53707=>"000000001",
  53708=>"111101000",
  53709=>"101011110",
  53710=>"111011001",
  53711=>"111111100",
  53712=>"110010000",
  53713=>"111100110",
  53714=>"101111111",
  53715=>"011110000",
  53716=>"000000011",
  53717=>"000111001",
  53718=>"011111000",
  53719=>"000001111",
  53720=>"000000011",
  53721=>"101011011",
  53722=>"100111110",
  53723=>"110000000",
  53724=>"111101111",
  53725=>"111010111",
  53726=>"111101010",
  53727=>"000000000",
  53728=>"101101011",
  53729=>"100000010",
  53730=>"110101000",
  53731=>"110111111",
  53732=>"000000001",
  53733=>"000000011",
  53734=>"111010111",
  53735=>"111111001",
  53736=>"111000000",
  53737=>"011111111",
  53738=>"110110100",
  53739=>"111111110",
  53740=>"000011011",
  53741=>"000000000",
  53742=>"001111010",
  53743=>"000101000",
  53744=>"000010010",
  53745=>"001000000",
  53746=>"000000000",
  53747=>"111011000",
  53748=>"000110010",
  53749=>"111000000",
  53750=>"111011000",
  53751=>"111111100",
  53752=>"000000111",
  53753=>"011000111",
  53754=>"111111110",
  53755=>"000111110",
  53756=>"110111110",
  53757=>"111111111",
  53758=>"101011011",
  53759=>"010010000",
  53760=>"011001110",
  53761=>"010010010",
  53762=>"000000111",
  53763=>"101101000",
  53764=>"111011001",
  53765=>"000001011",
  53766=>"111110000",
  53767=>"111111101",
  53768=>"001101110",
  53769=>"000010111",
  53770=>"111100001",
  53771=>"100101101",
  53772=>"101101000",
  53773=>"010111000",
  53774=>"011111100",
  53775=>"111111011",
  53776=>"111111011",
  53777=>"111111000",
  53778=>"000111111",
  53779=>"000010000",
  53780=>"000111010",
  53781=>"011111100",
  53782=>"111111011",
  53783=>"000111001",
  53784=>"001110111",
  53785=>"011001001",
  53786=>"001111011",
  53787=>"000000000",
  53788=>"110000000",
  53789=>"000000000",
  53790=>"000110011",
  53791=>"110110000",
  53792=>"010000000",
  53793=>"101101010",
  53794=>"101010111",
  53795=>"000000111",
  53796=>"111111011",
  53797=>"000001000",
  53798=>"000101101",
  53799=>"111011111",
  53800=>"100001000",
  53801=>"000000111",
  53802=>"000100000",
  53803=>"101010001",
  53804=>"000111000",
  53805=>"111000000",
  53806=>"100010101",
  53807=>"111110000",
  53808=>"111101000",
  53809=>"111001011",
  53810=>"011010111",
  53811=>"010011000",
  53812=>"000000000",
  53813=>"001000000",
  53814=>"010010000",
  53815=>"111000000",
  53816=>"001100111",
  53817=>"110100000",
  53818=>"101101010",
  53819=>"100101101",
  53820=>"010000000",
  53821=>"011010111",
  53822=>"101001000",
  53823=>"101110000",
  53824=>"000000111",
  53825=>"010000110",
  53826=>"000010000",
  53827=>"011011100",
  53828=>"001101111",
  53829=>"001000000",
  53830=>"100110000",
  53831=>"111111111",
  53832=>"101100011",
  53833=>"001000000",
  53834=>"111111000",
  53835=>"010111001",
  53836=>"001001011",
  53837=>"001011010",
  53838=>"000100100",
  53839=>"100000101",
  53840=>"000000000",
  53841=>"000111111",
  53842=>"101001111",
  53843=>"111100010",
  53844=>"000010001",
  53845=>"000100011",
  53846=>"011111000",
  53847=>"000001011",
  53848=>"000000101",
  53849=>"111111110",
  53850=>"111000000",
  53851=>"111111010",
  53852=>"000111111",
  53853=>"001100000",
  53854=>"010010111",
  53855=>"110011000",
  53856=>"000011110",
  53857=>"010000010",
  53858=>"000000111",
  53859=>"111001000",
  53860=>"111101000",
  53861=>"011111000",
  53862=>"010001000",
  53863=>"000000010",
  53864=>"111111010",
  53865=>"000000111",
  53866=>"011010111",
  53867=>"010000001",
  53868=>"000000111",
  53869=>"001101000",
  53870=>"110000000",
  53871=>"001011010",
  53872=>"111111000",
  53873=>"111100110",
  53874=>"010010000",
  53875=>"000000001",
  53876=>"011010000",
  53877=>"000100000",
  53878=>"010100000",
  53879=>"000000111",
  53880=>"000010111",
  53881=>"010111111",
  53882=>"111010000",
  53883=>"000111111",
  53884=>"111011110",
  53885=>"100001001",
  53886=>"111111111",
  53887=>"000000010",
  53888=>"001001111",
  53889=>"111000111",
  53890=>"000101111",
  53891=>"100100111",
  53892=>"000000010",
  53893=>"111111111",
  53894=>"000000000",
  53895=>"100001000",
  53896=>"100100000",
  53897=>"111000111",
  53898=>"101000111",
  53899=>"000000111",
  53900=>"000000011",
  53901=>"101000111",
  53902=>"111101000",
  53903=>"100100000",
  53904=>"101101000",
  53905=>"111111001",
  53906=>"000101000",
  53907=>"010011101",
  53908=>"001010000",
  53909=>"000000010",
  53910=>"010000000",
  53911=>"011000000",
  53912=>"110010000",
  53913=>"000110111",
  53914=>"000101101",
  53915=>"010000101",
  53916=>"110011111",
  53917=>"000101111",
  53918=>"000010000",
  53919=>"111011000",
  53920=>"101001111",
  53921=>"111111111",
  53922=>"011110100",
  53923=>"101100111",
  53924=>"000111000",
  53925=>"011001010",
  53926=>"000000000",
  53927=>"000111010",
  53928=>"001100101",
  53929=>"111010000",
  53930=>"111000000",
  53931=>"000110011",
  53932=>"101110110",
  53933=>"101101111",
  53934=>"111111001",
  53935=>"111000001",
  53936=>"000110000",
  53937=>"011001000",
  53938=>"110000000",
  53939=>"000001111",
  53940=>"000111000",
  53941=>"111111000",
  53942=>"000000000",
  53943=>"000000111",
  53944=>"110000000",
  53945=>"101001001",
  53946=>"000000111",
  53947=>"110101111",
  53948=>"000000000",
  53949=>"001000101",
  53950=>"000000111",
  53951=>"111000000",
  53952=>"111101000",
  53953=>"010000000",
  53954=>"111111000",
  53955=>"001100000",
  53956=>"100111111",
  53957=>"111101001",
  53958=>"100011011",
  53959=>"000111111",
  53960=>"000110110",
  53961=>"110010011",
  53962=>"111101100",
  53963=>"110000000",
  53964=>"010011000",
  53965=>"111110111",
  53966=>"000110000",
  53967=>"011001110",
  53968=>"111000000",
  53969=>"111111100",
  53970=>"111000101",
  53971=>"111111011",
  53972=>"111001001",
  53973=>"100011000",
  53974=>"111111000",
  53975=>"010011000",
  53976=>"111111000",
  53977=>"101011110",
  53978=>"101100111",
  53979=>"001000111",
  53980=>"111110100",
  53981=>"000000000",
  53982=>"111010011",
  53983=>"001000001",
  53984=>"000001111",
  53985=>"000000000",
  53986=>"111110000",
  53987=>"111111001",
  53988=>"000001000",
  53989=>"111111001",
  53990=>"000110110",
  53991=>"111111111",
  53992=>"111000110",
  53993=>"000000000",
  53994=>"110001100",
  53995=>"000000000",
  53996=>"000111000",
  53997=>"000000101",
  53998=>"000111000",
  53999=>"101111110",
  54000=>"001100000",
  54001=>"011001100",
  54002=>"111111000",
  54003=>"001011000",
  54004=>"111111011",
  54005=>"000000000",
  54006=>"100000111",
  54007=>"010000100",
  54008=>"101110111",
  54009=>"111111001",
  54010=>"101001011",
  54011=>"001000000",
  54012=>"111111000",
  54013=>"111110000",
  54014=>"000011110",
  54015=>"111111000",
  54016=>"011000000",
  54017=>"000001000",
  54018=>"000000000",
  54019=>"000000000",
  54020=>"000000001",
  54021=>"101100110",
  54022=>"010000000",
  54023=>"001000010",
  54024=>"000001111",
  54025=>"101101111",
  54026=>"001000000",
  54027=>"000000111",
  54028=>"111010110",
  54029=>"111000110",
  54030=>"000001011",
  54031=>"000000000",
  54032=>"111111111",
  54033=>"010000111",
  54034=>"000110010",
  54035=>"000011111",
  54036=>"000010110",
  54037=>"111111111",
  54038=>"000000000",
  54039=>"000000000",
  54040=>"010011001",
  54041=>"111111111",
  54042=>"111111111",
  54043=>"111111010",
  54044=>"111111111",
  54045=>"000001001",
  54046=>"000000010",
  54047=>"111111111",
  54048=>"100001000",
  54049=>"000010000",
  54050=>"000010000",
  54051=>"111111111",
  54052=>"000000000",
  54053=>"111111110",
  54054=>"111101100",
  54055=>"111001101",
  54056=>"111011001",
  54057=>"010000000",
  54058=>"001010101",
  54059=>"111111111",
  54060=>"010010000",
  54061=>"000000000",
  54062=>"001010000",
  54063=>"000000001",
  54064=>"000000000",
  54065=>"100000000",
  54066=>"001000001",
  54067=>"000001111",
  54068=>"010001000",
  54069=>"000001000",
  54070=>"111111001",
  54071=>"000000111",
  54072=>"000000000",
  54073=>"000010000",
  54074=>"011011001",
  54075=>"000000111",
  54076=>"000001111",
  54077=>"111111110",
  54078=>"000000110",
  54079=>"000000011",
  54080=>"100110110",
  54081=>"111111010",
  54082=>"111000000",
  54083=>"101101110",
  54084=>"110110110",
  54085=>"000010010",
  54086=>"010111100",
  54087=>"000000111",
  54088=>"001101100",
  54089=>"111110100",
  54090=>"000010010",
  54091=>"000000011",
  54092=>"111111111",
  54093=>"001000001",
  54094=>"001000000",
  54095=>"100000000",
  54096=>"111101101",
  54097=>"110000011",
  54098=>"001000111",
  54099=>"000000000",
  54100=>"010110010",
  54101=>"001011100",
  54102=>"000000000",
  54103=>"111111111",
  54104=>"000100000",
  54105=>"000000000",
  54106=>"101101100",
  54107=>"101101011",
  54108=>"001000000",
  54109=>"000001001",
  54110=>"111111111",
  54111=>"100011011",
  54112=>"101101111",
  54113=>"101100101",
  54114=>"111111110",
  54115=>"010111010",
  54116=>"101001100",
  54117=>"110011011",
  54118=>"011101100",
  54119=>"011111111",
  54120=>"000100110",
  54121=>"000000010",
  54122=>"111111111",
  54123=>"110111111",
  54124=>"111110111",
  54125=>"000000010",
  54126=>"111111111",
  54127=>"000100011",
  54128=>"001011011",
  54129=>"000000000",
  54130=>"111111110",
  54131=>"000110111",
  54132=>"111000000",
  54133=>"000100100",
  54134=>"000000100",
  54135=>"110100100",
  54136=>"111111111",
  54137=>"000100111",
  54138=>"000000000",
  54139=>"000000000",
  54140=>"000111111",
  54141=>"000000001",
  54142=>"001000000",
  54143=>"101111111",
  54144=>"111011000",
  54145=>"100100000",
  54146=>"111000000",
  54147=>"000000000",
  54148=>"000100000",
  54149=>"000110010",
  54150=>"111111011",
  54151=>"111111111",
  54152=>"111100011",
  54153=>"011010000",
  54154=>"000000000",
  54155=>"000000011",
  54156=>"111111010",
  54157=>"011011001",
  54158=>"000010111",
  54159=>"000001111",
  54160=>"001001001",
  54161=>"001010000",
  54162=>"111111111",
  54163=>"111110101",
  54164=>"011111111",
  54165=>"000000101",
  54166=>"110111011",
  54167=>"100000000",
  54168=>"111000100",
  54169=>"111111111",
  54170=>"111110111",
  54171=>"000001100",
  54172=>"011010000",
  54173=>"000000000",
  54174=>"111000000",
  54175=>"000000000",
  54176=>"011101000",
  54177=>"101101000",
  54178=>"111100000",
  54179=>"101000110",
  54180=>"111000001",
  54181=>"110111111",
  54182=>"000001011",
  54183=>"100000011",
  54184=>"010000110",
  54185=>"000000000",
  54186=>"101101101",
  54187=>"001010110",
  54188=>"001111011",
  54189=>"111110111",
  54190=>"000000011",
  54191=>"111111111",
  54192=>"101100010",
  54193=>"000000011",
  54194=>"000000011",
  54195=>"000000000",
  54196=>"000000100",
  54197=>"000000011",
  54198=>"011110110",
  54199=>"010111001",
  54200=>"011110111",
  54201=>"110111111",
  54202=>"111111001",
  54203=>"111100111",
  54204=>"000110111",
  54205=>"111111111",
  54206=>"001001111",
  54207=>"000000110",
  54208=>"111111111",
  54209=>"111111011",
  54210=>"000000111",
  54211=>"100100100",
  54212=>"111111000",
  54213=>"000000111",
  54214=>"100000001",
  54215=>"100001010",
  54216=>"111011011",
  54217=>"111111111",
  54218=>"110011001",
  54219=>"111110110",
  54220=>"000100011",
  54221=>"010011111",
  54222=>"100110111",
  54223=>"000000000",
  54224=>"000010000",
  54225=>"001001011",
  54226=>"111111110",
  54227=>"000000000",
  54228=>"011100010",
  54229=>"000000001",
  54230=>"110110010",
  54231=>"111000011",
  54232=>"111010000",
  54233=>"000000111",
  54234=>"000000010",
  54235=>"010000000",
  54236=>"011010101",
  54237=>"000001100",
  54238=>"110111111",
  54239=>"010000000",
  54240=>"010111111",
  54241=>"010000000",
  54242=>"111111111",
  54243=>"100000100",
  54244=>"110111110",
  54245=>"110111111",
  54246=>"111111111",
  54247=>"001000100",
  54248=>"100000000",
  54249=>"100000000",
  54250=>"000000000",
  54251=>"101000111",
  54252=>"111111111",
  54253=>"000010010",
  54254=>"000000000",
  54255=>"100000000",
  54256=>"101111111",
  54257=>"000000011",
  54258=>"001000111",
  54259=>"000000000",
  54260=>"100000000",
  54261=>"011011000",
  54262=>"010010111",
  54263=>"101000100",
  54264=>"111110110",
  54265=>"000000000",
  54266=>"000000000",
  54267=>"000000111",
  54268=>"000000000",
  54269=>"110000110",
  54270=>"000011111",
  54271=>"010000000",
  54272=>"110000000",
  54273=>"000111111",
  54274=>"101000000",
  54275=>"111000010",
  54276=>"100000111",
  54277=>"000000000",
  54278=>"101010100",
  54279=>"101110110",
  54280=>"101100111",
  54281=>"000000100",
  54282=>"000011000",
  54283=>"111010110",
  54284=>"111111011",
  54285=>"000000000",
  54286=>"000100110",
  54287=>"111111010",
  54288=>"110010000",
  54289=>"111011111",
  54290=>"111101111",
  54291=>"000000100",
  54292=>"101101111",
  54293=>"101101101",
  54294=>"110011011",
  54295=>"101111011",
  54296=>"010111001",
  54297=>"101111100",
  54298=>"000110000",
  54299=>"001000111",
  54300=>"101101101",
  54301=>"001111111",
  54302=>"011110000",
  54303=>"111000000",
  54304=>"111101111",
  54305=>"111111111",
  54306=>"000010111",
  54307=>"000111111",
  54308=>"101111111",
  54309=>"000000011",
  54310=>"000000001",
  54311=>"110111111",
  54312=>"111001111",
  54313=>"011111111",
  54314=>"000111000",
  54315=>"110111011",
  54316=>"000000100",
  54317=>"000111111",
  54318=>"101100000",
  54319=>"110110111",
  54320=>"111000111",
  54321=>"000000111",
  54322=>"111111010",
  54323=>"010110101",
  54324=>"000010000",
  54325=>"111111110",
  54326=>"001011110",
  54327=>"000100111",
  54328=>"110000000",
  54329=>"000000011",
  54330=>"110000011",
  54331=>"000000000",
  54332=>"001101001",
  54333=>"010110110",
  54334=>"000000000",
  54335=>"110001110",
  54336=>"100000111",
  54337=>"000000111",
  54338=>"001000000",
  54339=>"110110001",
  54340=>"111001000",
  54341=>"101001001",
  54342=>"001000000",
  54343=>"011101000",
  54344=>"110101011",
  54345=>"001101001",
  54346=>"111110110",
  54347=>"101001100",
  54348=>"100000001",
  54349=>"101100100",
  54350=>"011000111",
  54351=>"100100000",
  54352=>"101111111",
  54353=>"111010000",
  54354=>"111011110",
  54355=>"111001001",
  54356=>"011000101",
  54357=>"111111100",
  54358=>"111111110",
  54359=>"000000000",
  54360=>"111000001",
  54361=>"100101011",
  54362=>"000000011",
  54363=>"101111110",
  54364=>"001001010",
  54365=>"010000110",
  54366=>"111101111",
  54367=>"011010100",
  54368=>"000110000",
  54369=>"101011000",
  54370=>"101000000",
  54371=>"110111111",
  54372=>"101000111",
  54373=>"111111111",
  54374=>"111011010",
  54375=>"000000010",
  54376=>"101111101",
  54377=>"111000000",
  54378=>"111100111",
  54379=>"111000000",
  54380=>"100010111",
  54381=>"000000000",
  54382=>"000000000",
  54383=>"000111000",
  54384=>"010001000",
  54385=>"000000110",
  54386=>"100010001",
  54387=>"000000000",
  54388=>"011000000",
  54389=>"001000100",
  54390=>"000000000",
  54391=>"000000000",
  54392=>"111000010",
  54393=>"110001000",
  54394=>"001001000",
  54395=>"110101110",
  54396=>"111010101",
  54397=>"111100100",
  54398=>"001111111",
  54399=>"101000001",
  54400=>"101001000",
  54401=>"111110010",
  54402=>"101100011",
  54403=>"101000111",
  54404=>"100001111",
  54405=>"111101101",
  54406=>"001000010",
  54407=>"000001001",
  54408=>"001100000",
  54409=>"001000101",
  54410=>"111100111",
  54411=>"111001000",
  54412=>"100101100",
  54413=>"000000100",
  54414=>"010001101",
  54415=>"000100000",
  54416=>"011111011",
  54417=>"001000000",
  54418=>"000000000",
  54419=>"110111000",
  54420=>"011010000",
  54421=>"101111000",
  54422=>"111010110",
  54423=>"110101111",
  54424=>"111111111",
  54425=>"000010101",
  54426=>"111000101",
  54427=>"100000000",
  54428=>"010100111",
  54429=>"000001001",
  54430=>"111010010",
  54431=>"000010001",
  54432=>"001001000",
  54433=>"001111110",
  54434=>"000110000",
  54435=>"000111111",
  54436=>"010010100",
  54437=>"001101110",
  54438=>"001001000",
  54439=>"000011001",
  54440=>"000111111",
  54441=>"000101111",
  54442=>"111000001",
  54443=>"010000011",
  54444=>"100000111",
  54445=>"101000101",
  54446=>"011001111",
  54447=>"000101101",
  54448=>"110111111",
  54449=>"110010100",
  54450=>"110000010",
  54451=>"000100010",
  54452=>"110111111",
  54453=>"100111111",
  54454=>"110011101",
  54455=>"001000000",
  54456=>"000101101",
  54457=>"110011000",
  54458=>"101001010",
  54459=>"111111000",
  54460=>"000000111",
  54461=>"001010100",
  54462=>"001000001",
  54463=>"111010000",
  54464=>"111001000",
  54465=>"000000000",
  54466=>"101001011",
  54467=>"010000111",
  54468=>"001001000",
  54469=>"111100000",
  54470=>"000000010",
  54471=>"111101100",
  54472=>"000110111",
  54473=>"000000001",
  54474=>"111111110",
  54475=>"111000001",
  54476=>"000100111",
  54477=>"010010100",
  54478=>"000001001",
  54479=>"110100100",
  54480=>"000000110",
  54481=>"011101111",
  54482=>"100110111",
  54483=>"110111101",
  54484=>"101001000",
  54485=>"011110010",
  54486=>"000010000",
  54487=>"000000111",
  54488=>"000111111",
  54489=>"000001001",
  54490=>"110101000",
  54491=>"111000100",
  54492=>"111100110",
  54493=>"101010010",
  54494=>"011010000",
  54495=>"111101011",
  54496=>"001000110",
  54497=>"011100010",
  54498=>"111000011",
  54499=>"111001111",
  54500=>"001101101",
  54501=>"111000000",
  54502=>"000000000",
  54503=>"100000101",
  54504=>"001001011",
  54505=>"000111000",
  54506=>"011010000",
  54507=>"001000000",
  54508=>"000010111",
  54509=>"111111000",
  54510=>"000000000",
  54511=>"001000000",
  54512=>"000000110",
  54513=>"001001101",
  54514=>"101001110",
  54515=>"011011111",
  54516=>"001100000",
  54517=>"000100101",
  54518=>"101000000",
  54519=>"000000010",
  54520=>"000100000",
  54521=>"010110110",
  54522=>"111110000",
  54523=>"010100010",
  54524=>"011000101",
  54525=>"111000111",
  54526=>"011011111",
  54527=>"000000100",
  54528=>"011001001",
  54529=>"110100100",
  54530=>"110000110",
  54531=>"100000000",
  54532=>"100111011",
  54533=>"000000010",
  54534=>"000000000",
  54535=>"110111111",
  54536=>"000110100",
  54537=>"000011011",
  54538=>"010001011",
  54539=>"000011011",
  54540=>"000100100",
  54541=>"100100111",
  54542=>"010111001",
  54543=>"001000100",
  54544=>"011011000",
  54545=>"100100010",
  54546=>"100000011",
  54547=>"000101111",
  54548=>"111111010",
  54549=>"011000100",
  54550=>"011100100",
  54551=>"000111111",
  54552=>"000011010",
  54553=>"111011011",
  54554=>"111011010",
  54555=>"100000000",
  54556=>"000100100",
  54557=>"110011111",
  54558=>"010011010",
  54559=>"100000000",
  54560=>"111101000",
  54561=>"110100100",
  54562=>"111101111",
  54563=>"000100101",
  54564=>"100011001",
  54565=>"011010010",
  54566=>"111011010",
  54567=>"000000000",
  54568=>"111000000",
  54569=>"111111100",
  54570=>"000100100",
  54571=>"000000000",
  54572=>"111110111",
  54573=>"111111111",
  54574=>"011011110",
  54575=>"000000111",
  54576=>"111000000",
  54577=>"111011100",
  54578=>"011100000",
  54579=>"111110000",
  54580=>"101000000",
  54581=>"011000111",
  54582=>"000110101",
  54583=>"000000011",
  54584=>"000100001",
  54585=>"000100100",
  54586=>"011100110",
  54587=>"000000000",
  54588=>"100111001",
  54589=>"011100000",
  54590=>"100000000",
  54591=>"000011011",
  54592=>"111111000",
  54593=>"111011000",
  54594=>"111110101",
  54595=>"000011011",
  54596=>"011000100",
  54597=>"011000000",
  54598=>"000100000",
  54599=>"111100111",
  54600=>"011111110",
  54601=>"001011011",
  54602=>"111011000",
  54603=>"111100100",
  54604=>"011011011",
  54605=>"001011000",
  54606=>"000110110",
  54607=>"011111100",
  54608=>"001100000",
  54609=>"011101001",
  54610=>"111110111",
  54611=>"010101100",
  54612=>"000111011",
  54613=>"000011011",
  54614=>"000110010",
  54615=>"000011011",
  54616=>"111010100",
  54617=>"010110110",
  54618=>"000001000",
  54619=>"011011011",
  54620=>"000000000",
  54621=>"011100010",
  54622=>"111100100",
  54623=>"110011011",
  54624=>"100100100",
  54625=>"001111111",
  54626=>"111000100",
  54627=>"001110111",
  54628=>"000010000",
  54629=>"110110000",
  54630=>"100011000",
  54631=>"001011011",
  54632=>"000111111",
  54633=>"101110011",
  54634=>"011011001",
  54635=>"111111101",
  54636=>"100000110",
  54637=>"101100011",
  54638=>"000110000",
  54639=>"111100000",
  54640=>"101001001",
  54641=>"001010111",
  54642=>"001001000",
  54643=>"111000100",
  54644=>"011010000",
  54645=>"001000000",
  54646=>"000000011",
  54647=>"011011011",
  54648=>"111000000",
  54649=>"100100011",
  54650=>"111100100",
  54651=>"000000101",
  54652=>"000110010",
  54653=>"011110000",
  54654=>"010000000",
  54655=>"000111011",
  54656=>"111000101",
  54657=>"000011011",
  54658=>"011011000",
  54659=>"110100001",
  54660=>"011011100",
  54661=>"110111111",
  54662=>"011111001",
  54663=>"000010011",
  54664=>"110110011",
  54665=>"110111100",
  54666=>"011000000",
  54667=>"100000110",
  54668=>"000011010",
  54669=>"000000101",
  54670=>"000001111",
  54671=>"000000000",
  54672=>"011101110",
  54673=>"000010010",
  54674=>"000011000",
  54675=>"110100000",
  54676=>"010111111",
  54677=>"000000000",
  54678=>"111111111",
  54679=>"010000100",
  54680=>"000100000",
  54681=>"011111011",
  54682=>"001001000",
  54683=>"010000100",
  54684=>"110100100",
  54685=>"001011010",
  54686=>"101101110",
  54687=>"011000000",
  54688=>"100010111",
  54689=>"100111111",
  54690=>"110000000",
  54691=>"000101000",
  54692=>"011101000",
  54693=>"001111111",
  54694=>"101100111",
  54695=>"001100100",
  54696=>"010000110",
  54697=>"000100000",
  54698=>"100100110",
  54699=>"010000100",
  54700=>"111000111",
  54701=>"001011000",
  54702=>"001100000",
  54703=>"000000100",
  54704=>"100111110",
  54705=>"101000100",
  54706=>"001111111",
  54707=>"001100000",
  54708=>"000111111",
  54709=>"110100111",
  54710=>"011111101",
  54711=>"011100000",
  54712=>"011011010",
  54713=>"000111011",
  54714=>"000011001",
  54715=>"011011001",
  54716=>"111111100",
  54717=>"011000000",
  54718=>"010010111",
  54719=>"001000010",
  54720=>"010011010",
  54721=>"100011011",
  54722=>"011000011",
  54723=>"100010110",
  54724=>"000000000",
  54725=>"110000000",
  54726=>"000000011",
  54727=>"101111011",
  54728=>"100111110",
  54729=>"000011011",
  54730=>"111101111",
  54731=>"000011000",
  54732=>"000011001",
  54733=>"000001011",
  54734=>"000000011",
  54735=>"100111011",
  54736=>"000000111",
  54737=>"011001001",
  54738=>"110111011",
  54739=>"000000100",
  54740=>"111000100",
  54741=>"110100100",
  54742=>"000100010",
  54743=>"110000000",
  54744=>"110100011",
  54745=>"100100100",
  54746=>"100000100",
  54747=>"111100111",
  54748=>"110111111",
  54749=>"110101011",
  54750=>"010000000",
  54751=>"010011000",
  54752=>"000000000",
  54753=>"010100100",
  54754=>"000111011",
  54755=>"101111111",
  54756=>"100011000",
  54757=>"111100101",
  54758=>"000000000",
  54759=>"000110001",
  54760=>"001000111",
  54761=>"110000000",
  54762=>"000010000",
  54763=>"010101111",
  54764=>"000000100",
  54765=>"000000111",
  54766=>"000000000",
  54767=>"000001001",
  54768=>"111111011",
  54769=>"001001101",
  54770=>"000000011",
  54771=>"001001101",
  54772=>"101101010",
  54773=>"000000100",
  54774=>"000000001",
  54775=>"000000101",
  54776=>"000100000",
  54777=>"100110011",
  54778=>"010000110",
  54779=>"000001111",
  54780=>"111100100",
  54781=>"010011011",
  54782=>"010110000",
  54783=>"110000000",
  54784=>"000011100",
  54785=>"000000010",
  54786=>"010010010",
  54787=>"001101111",
  54788=>"000000011",
  54789=>"000000001",
  54790=>"011111111",
  54791=>"110111011",
  54792=>"000000100",
  54793=>"111010101",
  54794=>"111111111",
  54795=>"110111010",
  54796=>"000111111",
  54797=>"000101000",
  54798=>"111111110",
  54799=>"111111111",
  54800=>"000000111",
  54801=>"111110111",
  54802=>"111110110",
  54803=>"111000111",
  54804=>"011111101",
  54805=>"000000101",
  54806=>"011111101",
  54807=>"111111111",
  54808=>"000001100",
  54809=>"000000111",
  54810=>"000000000",
  54811=>"010100100",
  54812=>"000000000",
  54813=>"111101000",
  54814=>"001111111",
  54815=>"101100000",
  54816=>"000111101",
  54817=>"110111000",
  54818=>"001101100",
  54819=>"000010011",
  54820=>"001011111",
  54821=>"000001001",
  54822=>"000111110",
  54823=>"110111111",
  54824=>"111011110",
  54825=>"000000000",
  54826=>"111111101",
  54827=>"000000100",
  54828=>"000001011",
  54829=>"000000010",
  54830=>"000000110",
  54831=>"110011000",
  54832=>"000101001",
  54833=>"110110111",
  54834=>"000101001",
  54835=>"001101000",
  54836=>"110111111",
  54837=>"000110001",
  54838=>"111111111",
  54839=>"101111100",
  54840=>"000101111",
  54841=>"111101000",
  54842=>"111101000",
  54843=>"000101111",
  54844=>"000000000",
  54845=>"111111111",
  54846=>"000101111",
  54847=>"100100100",
  54848=>"000001111",
  54849=>"000000000",
  54850=>"101001101",
  54851=>"111111111",
  54852=>"111111111",
  54853=>"000000111",
  54854=>"111110111",
  54855=>"000001011",
  54856=>"000000000",
  54857=>"111101000",
  54858=>"111101101",
  54859=>"110000010",
  54860=>"000000000",
  54861=>"110100111",
  54862=>"001010110",
  54863=>"000000111",
  54864=>"111111111",
  54865=>"100011101",
  54866=>"001011001",
  54867=>"000001000",
  54868=>"000010010",
  54869=>"000001000",
  54870=>"111011010",
  54871=>"110111111",
  54872=>"001000101",
  54873=>"110100101",
  54874=>"111101011",
  54875=>"111000111",
  54876=>"000000000",
  54877=>"100100111",
  54878=>"000000111",
  54879=>"110111111",
  54880=>"000011000",
  54881=>"010010000",
  54882=>"110111111",
  54883=>"111011000",
  54884=>"001000101",
  54885=>"011100000",
  54886=>"000000000",
  54887=>"111111100",
  54888=>"111111110",
  54889=>"111101000",
  54890=>"000100000",
  54891=>"001000000",
  54892=>"000111111",
  54893=>"111011011",
  54894=>"111111101",
  54895=>"111011000",
  54896=>"011011011",
  54897=>"010101000",
  54898=>"111111111",
  54899=>"000000000",
  54900=>"011110000",
  54901=>"000000000",
  54902=>"000111100",
  54903=>"000111111",
  54904=>"010110110",
  54905=>"111111000",
  54906=>"111110000",
  54907=>"001101111",
  54908=>"111111111",
  54909=>"011000001",
  54910=>"111101111",
  54911=>"010010011",
  54912=>"001001010",
  54913=>"011000101",
  54914=>"000000000",
  54915=>"101111101",
  54916=>"010110010",
  54917=>"000000000",
  54918=>"000000100",
  54919=>"101000110",
  54920=>"000100111",
  54921=>"111011010",
  54922=>"000000000",
  54923=>"101000010",
  54924=>"001000010",
  54925=>"000010000",
  54926=>"000000000",
  54927=>"010110011",
  54928=>"111101100",
  54929=>"100000000",
  54930=>"100011011",
  54931=>"111110000",
  54932=>"000000000",
  54933=>"111111111",
  54934=>"000000010",
  54935=>"000100000",
  54936=>"000010010",
  54937=>"101001000",
  54938=>"110110010",
  54939=>"000010011",
  54940=>"000110111",
  54941=>"000000111",
  54942=>"010001001",
  54943=>"011011000",
  54944=>"000000100",
  54945=>"000111000",
  54946=>"000000100",
  54947=>"111111111",
  54948=>"110111111",
  54949=>"001010011",
  54950=>"001000000",
  54951=>"000000111",
  54952=>"111100000",
  54953=>"000000000",
  54954=>"110100100",
  54955=>"011111111",
  54956=>"001011000",
  54957=>"111010000",
  54958=>"111101111",
  54959=>"001000000",
  54960=>"000000001",
  54961=>"111011001",
  54962=>"000110010",
  54963=>"011111111",
  54964=>"111100100",
  54965=>"111111010",
  54966=>"000111011",
  54967=>"000000101",
  54968=>"000000000",
  54969=>"000010001",
  54970=>"000000000",
  54971=>"000111111",
  54972=>"000000000",
  54973=>"111111111",
  54974=>"000001000",
  54975=>"111011000",
  54976=>"000000111",
  54977=>"111000111",
  54978=>"001000011",
  54979=>"110110010",
  54980=>"000001111",
  54981=>"100001000",
  54982=>"111111111",
  54983=>"000001000",
  54984=>"111101101",
  54985=>"000011010",
  54986=>"010101111",
  54987=>"010010111",
  54988=>"100100000",
  54989=>"111111011",
  54990=>"111111111",
  54991=>"111111111",
  54992=>"111111111",
  54993=>"000010000",
  54994=>"101000001",
  54995=>"111111010",
  54996=>"000000011",
  54997=>"011111101",
  54998=>"000011000",
  54999=>"011101000",
  55000=>"000000000",
  55001=>"111010000",
  55002=>"001001000",
  55003=>"111111111",
  55004=>"101111000",
  55005=>"111000000",
  55006=>"111100110",
  55007=>"001000000",
  55008=>"111111110",
  55009=>"011101000",
  55010=>"101000001",
  55011=>"011011011",
  55012=>"111000000",
  55013=>"000000000",
  55014=>"000000000",
  55015=>"111111111",
  55016=>"000100110",
  55017=>"101111110",
  55018=>"111111111",
  55019=>"000111111",
  55020=>"000111111",
  55021=>"010111010",
  55022=>"111110000",
  55023=>"100000000",
  55024=>"000000010",
  55025=>"000000000",
  55026=>"000011000",
  55027=>"011001000",
  55028=>"001100101",
  55029=>"111111111",
  55030=>"000011111",
  55031=>"101101111",
  55032=>"011111111",
  55033=>"111111111",
  55034=>"000000001",
  55035=>"001000000",
  55036=>"000100110",
  55037=>"111010110",
  55038=>"110001110",
  55039=>"000111111",
  55040=>"011001100",
  55041=>"111100100",
  55042=>"111100100",
  55043=>"000101111",
  55044=>"111110111",
  55045=>"111110101",
  55046=>"000011011",
  55047=>"001100010",
  55048=>"000000110",
  55049=>"000000000",
  55050=>"010110011",
  55051=>"101011111",
  55052=>"000100010",
  55053=>"000010000",
  55054=>"110110110",
  55055=>"000110010",
  55056=>"100111101",
  55057=>"000011010",
  55058=>"111001010",
  55059=>"010000000",
  55060=>"001100100",
  55061=>"111101101",
  55062=>"111101101",
  55063=>"101111111",
  55064=>"111101000",
  55065=>"111111010",
  55066=>"011111111",
  55067=>"001101110",
  55068=>"011111111",
  55069=>"000011111",
  55070=>"010101101",
  55071=>"011111110",
  55072=>"111101101",
  55073=>"111100100",
  55074=>"101100110",
  55075=>"111100001",
  55076=>"011110110",
  55077=>"001100111",
  55078=>"110100100",
  55079=>"000001010",
  55080=>"111101111",
  55081=>"101100111",
  55082=>"100010011",
  55083=>"111011110",
  55084=>"000110111",
  55085=>"011011000",
  55086=>"101111100",
  55087=>"110110100",
  55088=>"010111101",
  55089=>"111111001",
  55090=>"001111111",
  55091=>"110111111",
  55092=>"000000100",
  55093=>"110010100",
  55094=>"101100000",
  55095=>"000000000",
  55096=>"011111110",
  55097=>"000000000",
  55098=>"100100010",
  55099=>"110011000",
  55100=>"011000110",
  55101=>"111111000",
  55102=>"111100100",
  55103=>"000111011",
  55104=>"000101001",
  55105=>"000110100",
  55106=>"010100100",
  55107=>"111111000",
  55108=>"000010010",
  55109=>"000000000",
  55110=>"000000000",
  55111=>"001101011",
  55112=>"011101000",
  55113=>"100101111",
  55114=>"110110101",
  55115=>"100111011",
  55116=>"111101011",
  55117=>"100101111",
  55118=>"101100110",
  55119=>"110110100",
  55120=>"111111000",
  55121=>"111100100",
  55122=>"000010111",
  55123=>"000011011",
  55124=>"010000101",
  55125=>"011000100",
  55126=>"000010010",
  55127=>"111000100",
  55128=>"100111110",
  55129=>"000000001",
  55130=>"011101011",
  55131=>"000000110",
  55132=>"000010010",
  55133=>"011011000",
  55134=>"111111101",
  55135=>"111100000",
  55136=>"111111111",
  55137=>"000000000",
  55138=>"100000100",
  55139=>"011110000",
  55140=>"111000100",
  55141=>"111000100",
  55142=>"000000000",
  55143=>"101001011",
  55144=>"011000111",
  55145=>"010100111",
  55146=>"111111011",
  55147=>"100101111",
  55148=>"010000100",
  55149=>"010010010",
  55150=>"000000000",
  55151=>"000001010",
  55152=>"100111111",
  55153=>"000101100",
  55154=>"110001000",
  55155=>"001111111",
  55156=>"000000000",
  55157=>"010000100",
  55158=>"010111111",
  55159=>"100100000",
  55160=>"111111000",
  55161=>"100110010",
  55162=>"000101000",
  55163=>"000111100",
  55164=>"111111011",
  55165=>"011000000",
  55166=>"111100101",
  55167=>"111111101",
  55168=>"100011000",
  55169=>"111000000",
  55170=>"110110100",
  55171=>"000100111",
  55172=>"111111111",
  55173=>"111000010",
  55174=>"100100100",
  55175=>"010100000",
  55176=>"010111111",
  55177=>"010000000",
  55178=>"100000000",
  55179=>"100000011",
  55180=>"011100000",
  55181=>"000100000",
  55182=>"111111110",
  55183=>"010000000",
  55184=>"101100001",
  55185=>"011001101",
  55186=>"000000000",
  55187=>"111101101",
  55188=>"010111101",
  55189=>"001101101",
  55190=>"100111111",
  55191=>"101011100",
  55192=>"000000101",
  55193=>"010111110",
  55194=>"000001110",
  55195=>"101100000",
  55196=>"111100100",
  55197=>"110101101",
  55198=>"000000110",
  55199=>"001111110",
  55200=>"110111010",
  55201=>"111011100",
  55202=>"000111010",
  55203=>"110111111",
  55204=>"111101111",
  55205=>"000110010",
  55206=>"100100101",
  55207=>"000000111",
  55208=>"000111011",
  55209=>"000001000",
  55210=>"111100000",
  55211=>"111100000",
  55212=>"101010011",
  55213=>"010011010",
  55214=>"011000000",
  55215=>"000010000",
  55216=>"100011011",
  55217=>"111111111",
  55218=>"000010000",
  55219=>"110011000",
  55220=>"000001011",
  55221=>"100111000",
  55222=>"000011010",
  55223=>"011100000",
  55224=>"110110000",
  55225=>"000110101",
  55226=>"010000000",
  55227=>"010110111",
  55228=>"010000011",
  55229=>"011111111",
  55230=>"000011011",
  55231=>"010111101",
  55232=>"110010000",
  55233=>"111111111",
  55234=>"111010000",
  55235=>"100001011",
  55236=>"011010010",
  55237=>"110001101",
  55238=>"000000011",
  55239=>"011100101",
  55240=>"011101000",
  55241=>"111000100",
  55242=>"111111011",
  55243=>"111000100",
  55244=>"001011000",
  55245=>"111100111",
  55246=>"101010010",
  55247=>"011101100",
  55248=>"100000000",
  55249=>"010111011",
  55250=>"000100111",
  55251=>"000011011",
  55252=>"000000000",
  55253=>"111100001",
  55254=>"111101100",
  55255=>"100000101",
  55256=>"000011001",
  55257=>"010111000",
  55258=>"011111110",
  55259=>"101110000",
  55260=>"111100001",
  55261=>"001111000",
  55262=>"000011011",
  55263=>"000010000",
  55264=>"001100000",
  55265=>"110100000",
  55266=>"110111111",
  55267=>"000100110",
  55268=>"111100111",
  55269=>"100100101",
  55270=>"000111010",
  55271=>"100100000",
  55272=>"011011011",
  55273=>"000010010",
  55274=>"100100010",
  55275=>"100000100",
  55276=>"011010101",
  55277=>"100111111",
  55278=>"111000000",
  55279=>"000111111",
  55280=>"010011011",
  55281=>"011100100",
  55282=>"000101100",
  55283=>"100110110",
  55284=>"101000100",
  55285=>"111101000",
  55286=>"100000010",
  55287=>"001010011",
  55288=>"111111100",
  55289=>"111111011",
  55290=>"111111111",
  55291=>"000110111",
  55292=>"000101011",
  55293=>"011011111",
  55294=>"011011111",
  55295=>"111101001",
  55296=>"100001000",
  55297=>"101100100",
  55298=>"000000000",
  55299=>"001000111",
  55300=>"000000110",
  55301=>"000110010",
  55302=>"111011111",
  55303=>"110101000",
  55304=>"110010000",
  55305=>"110010010",
  55306=>"000110010",
  55307=>"000001011",
  55308=>"111101001",
  55309=>"100001001",
  55310=>"000100101",
  55311=>"111101000",
  55312=>"111110111",
  55313=>"111010010",
  55314=>"010000000",
  55315=>"001010010",
  55316=>"000101111",
  55317=>"101001001",
  55318=>"100100000",
  55319=>"110111110",
  55320=>"111000010",
  55321=>"110111111",
  55322=>"111111111",
  55323=>"101000110",
  55324=>"111100100",
  55325=>"110000000",
  55326=>"111111001",
  55327=>"010000000",
  55328=>"111010000",
  55329=>"000010110",
  55330=>"010000001",
  55331=>"111011010",
  55332=>"000110110",
  55333=>"000100001",
  55334=>"111110010",
  55335=>"000110110",
  55336=>"000011111",
  55337=>"111111110",
  55338=>"101111010",
  55339=>"010010001",
  55340=>"100111100",
  55341=>"101111011",
  55342=>"010000100",
  55343=>"000000100",
  55344=>"010010000",
  55345=>"010001100",
  55346=>"010010111",
  55347=>"000000101",
  55348=>"100110010",
  55349=>"000111111",
  55350=>"011011011",
  55351=>"000100000",
  55352=>"111010001",
  55353=>"111001000",
  55354=>"000000101",
  55355=>"100010010",
  55356=>"110000100",
  55357=>"111001000",
  55358=>"110010000",
  55359=>"000001111",
  55360=>"111110000",
  55361=>"111110010",
  55362=>"111000000",
  55363=>"110000000",
  55364=>"111111000",
  55365=>"000101111",
  55366=>"000101011",
  55367=>"011010111",
  55368=>"111110011",
  55369=>"111110000",
  55370=>"111000000",
  55371=>"000011110",
  55372=>"000000000",
  55373=>"010011000",
  55374=>"000101000",
  55375=>"000000101",
  55376=>"000010010",
  55377=>"111111111",
  55378=>"101111001",
  55379=>"000011000",
  55380=>"111000010",
  55381=>"100100100",
  55382=>"000011111",
  55383=>"111010110",
  55384=>"010000001",
  55385=>"011010011",
  55386=>"000100110",
  55387=>"010001011",
  55388=>"000111101",
  55389=>"010000000",
  55390=>"111111111",
  55391=>"001000000",
  55392=>"111111000",
  55393=>"000000000",
  55394=>"111010000",
  55395=>"000010001",
  55396=>"100000001",
  55397=>"000001011",
  55398=>"101000000",
  55399=>"000001101",
  55400=>"111000111",
  55401=>"111101101",
  55402=>"000010111",
  55403=>"000100000",
  55404=>"111000100",
  55405=>"000110110",
  55406=>"000001001",
  55407=>"000000000",
  55408=>"000100100",
  55409=>"000000000",
  55410=>"110110110",
  55411=>"000000000",
  55412=>"001001001",
  55413=>"101000000",
  55414=>"111001101",
  55415=>"111000000",
  55416=>"111001010",
  55417=>"000000000",
  55418=>"001010111",
  55419=>"000001001",
  55420=>"110100000",
  55421=>"000100000",
  55422=>"000010010",
  55423=>"000000000",
  55424=>"101111111",
  55425=>"111111000",
  55426=>"000101000",
  55427=>"010000010",
  55428=>"110011100",
  55429=>"000110111",
  55430=>"001001100",
  55431=>"000101001",
  55432=>"001001001",
  55433=>"001000011",
  55434=>"000101111",
  55435=>"010000101",
  55436=>"000100000",
  55437=>"000001000",
  55438=>"101101101",
  55439=>"001000100",
  55440=>"011000000",
  55441=>"111000011",
  55442=>"000111110",
  55443=>"011011001",
  55444=>"101100011",
  55445=>"111010000",
  55446=>"011111100",
  55447=>"000100100",
  55448=>"000101110",
  55449=>"101101111",
  55450=>"111101110",
  55451=>"111010000",
  55452=>"111000111",
  55453=>"111000000",
  55454=>"101111011",
  55455=>"111000000",
  55456=>"000011011",
  55457=>"101010000",
  55458=>"001000010",
  55459=>"101011010",
  55460=>"000000010",
  55461=>"000100100",
  55462=>"000000000",
  55463=>"000110110",
  55464=>"001100010",
  55465=>"000000000",
  55466=>"011101000",
  55467=>"111010000",
  55468=>"110100110",
  55469=>"000000000",
  55470=>"000000000",
  55471=>"000000000",
  55472=>"111101000",
  55473=>"000111111",
  55474=>"010000000",
  55475=>"110110110",
  55476=>"100110111",
  55477=>"111011111",
  55478=>"010100101",
  55479=>"000110111",
  55480=>"111001011",
  55481=>"111001100",
  55482=>"000101110",
  55483=>"111001010",
  55484=>"101101101",
  55485=>"010111011",
  55486=>"110010000",
  55487=>"010111000",
  55488=>"001000101",
  55489=>"000101100",
  55490=>"101111011",
  55491=>"110100100",
  55492=>"001000111",
  55493=>"000100000",
  55494=>"111101001",
  55495=>"111000000",
  55496=>"000100101",
  55497=>"101101000",
  55498=>"000111111",
  55499=>"001111111",
  55500=>"000000000",
  55501=>"111011000",
  55502=>"010111000",
  55503=>"000001111",
  55504=>"000000000",
  55505=>"000001001",
  55506=>"000100110",
  55507=>"111111000",
  55508=>"111101001",
  55509=>"000011011",
  55510=>"101110000",
  55511=>"000110111",
  55512=>"001101111",
  55513=>"001000110",
  55514=>"010100100",
  55515=>"010110111",
  55516=>"110101001",
  55517=>"000001100",
  55518=>"000001001",
  55519=>"010011010",
  55520=>"010000001",
  55521=>"111000101",
  55522=>"000101111",
  55523=>"011111111",
  55524=>"101011000",
  55525=>"010100111",
  55526=>"001001001",
  55527=>"000001000",
  55528=>"111001001",
  55529=>"000011010",
  55530=>"000010111",
  55531=>"111111000",
  55532=>"101101111",
  55533=>"000111000",
  55534=>"010111000",
  55535=>"000000000",
  55536=>"000010000",
  55537=>"000001001",
  55538=>"101000000",
  55539=>"000111111",
  55540=>"000100100",
  55541=>"000001001",
  55542=>"000100000",
  55543=>"111000111",
  55544=>"101010111",
  55545=>"010111101",
  55546=>"011111111",
  55547=>"000000001",
  55548=>"111111001",
  55549=>"000101111",
  55550=>"000000011",
  55551=>"000000000",
  55552=>"001011011",
  55553=>"000000000",
  55554=>"111000000",
  55555=>"100100111",
  55556=>"001011011",
  55557=>"111101001",
  55558=>"100000100",
  55559=>"111001010",
  55560=>"000100100",
  55561=>"000000100",
  55562=>"101001111",
  55563=>"010000111",
  55564=>"110000101",
  55565=>"111111100",
  55566=>"010011110",
  55567=>"101000110",
  55568=>"000000010",
  55569=>"101011111",
  55570=>"111100111",
  55571=>"011000000",
  55572=>"111011000",
  55573=>"100111011",
  55574=>"111000011",
  55575=>"111001011",
  55576=>"111000000",
  55577=>"000000000",
  55578=>"000100000",
  55579=>"110100100",
  55580=>"101100000",
  55581=>"100100000",
  55582=>"010110110",
  55583=>"000110110",
  55584=>"000000000",
  55585=>"000111111",
  55586=>"000111111",
  55587=>"000011010",
  55588=>"011111001",
  55589=>"111011000",
  55590=>"000010000",
  55591=>"100010000",
  55592=>"111001111",
  55593=>"101001001",
  55594=>"000000101",
  55595=>"000011010",
  55596=>"110100100",
  55597=>"000000001",
  55598=>"011111100",
  55599=>"000111010",
  55600=>"111110100",
  55601=>"001101011",
  55602=>"111011001",
  55603=>"111110010",
  55604=>"111101111",
  55605=>"010111011",
  55606=>"110111000",
  55607=>"000100110",
  55608=>"111110111",
  55609=>"111000001",
  55610=>"111111000",
  55611=>"001001011",
  55612=>"111010100",
  55613=>"110111011",
  55614=>"000000100",
  55615=>"011011001",
  55616=>"010011001",
  55617=>"000010010",
  55618=>"111110000",
  55619=>"011000100",
  55620=>"000011011",
  55621=>"101000100",
  55622=>"101000011",
  55623=>"000000000",
  55624=>"100111111",
  55625=>"111000000",
  55626=>"111000100",
  55627=>"101100101",
  55628=>"111011010",
  55629=>"110111110",
  55630=>"001001011",
  55631=>"100000011",
  55632=>"000000000",
  55633=>"110111000",
  55634=>"000000001",
  55635=>"000011100",
  55636=>"111101000",
  55637=>"111101100",
  55638=>"111111111",
  55639=>"100000001",
  55640=>"010111111",
  55641=>"011001000",
  55642=>"101011011",
  55643=>"011011000",
  55644=>"000010110",
  55645=>"101000111",
  55646=>"111110111",
  55647=>"000001000",
  55648=>"011011000",
  55649=>"000000010",
  55650=>"111000001",
  55651=>"111111111",
  55652=>"001000011",
  55653=>"011111011",
  55654=>"010001000",
  55655=>"000011011",
  55656=>"100000111",
  55657=>"101011010",
  55658=>"001100000",
  55659=>"000111000",
  55660=>"000111111",
  55661=>"100000011",
  55662=>"111111000",
  55663=>"101000101",
  55664=>"010111110",
  55665=>"000011100",
  55666=>"001000010",
  55667=>"000010001",
  55668=>"111100001",
  55669=>"101100010",
  55670=>"111001000",
  55671=>"001011011",
  55672=>"111011111",
  55673=>"110001111",
  55674=>"100101111",
  55675=>"000101111",
  55676=>"110100000",
  55677=>"010100100",
  55678=>"110111100",
  55679=>"111000000",
  55680=>"000010011",
  55681=>"111000000",
  55682=>"111111101",
  55683=>"000001011",
  55684=>"100100000",
  55685=>"011001001",
  55686=>"001010000",
  55687=>"101100000",
  55688=>"010000001",
  55689=>"100111010",
  55690=>"000000000",
  55691=>"010010000",
  55692=>"100110000",
  55693=>"101100001",
  55694=>"111000101",
  55695=>"110000100",
  55696=>"111111110",
  55697=>"111011011",
  55698=>"101000000",
  55699=>"100111100",
  55700=>"000100000",
  55701=>"010000100",
  55702=>"011000001",
  55703=>"000010001",
  55704=>"111011111",
  55705=>"111111100",
  55706=>"011011000",
  55707=>"000100100",
  55708=>"111100100",
  55709=>"001001111",
  55710=>"011110100",
  55711=>"010011001",
  55712=>"010010001",
  55713=>"001000000",
  55714=>"110000001",
  55715=>"110111110",
  55716=>"000111101",
  55717=>"110011011",
  55718=>"000110110",
  55719=>"010011111",
  55720=>"101110000",
  55721=>"100100000",
  55722=>"101100000",
  55723=>"101010110",
  55724=>"100000011",
  55725=>"101100100",
  55726=>"001000110",
  55727=>"000100111",
  55728=>"011101101",
  55729=>"010000000",
  55730=>"111101010",
  55731=>"111010010",
  55732=>"000001001",
  55733=>"011000000",
  55734=>"000011011",
  55735=>"000011011",
  55736=>"000000100",
  55737=>"100101001",
  55738=>"010001100",
  55739=>"111101101",
  55740=>"011010000",
  55741=>"111111111",
  55742=>"001001000",
  55743=>"110111101",
  55744=>"100011001",
  55745=>"000000010",
  55746=>"101111100",
  55747=>"001010110",
  55748=>"100101110",
  55749=>"001001011",
  55750=>"000110101",
  55751=>"111111101",
  55752=>"111000011",
  55753=>"000011011",
  55754=>"110111111",
  55755=>"100100111",
  55756=>"011000000",
  55757=>"001001100",
  55758=>"001000000",
  55759=>"100001101",
  55760=>"000010111",
  55761=>"000000011",
  55762=>"111100100",
  55763=>"100001111",
  55764=>"001010000",
  55765=>"101000000",
  55766=>"111100100",
  55767=>"011111111",
  55768=>"000000001",
  55769=>"010000011",
  55770=>"011001111",
  55771=>"111000101",
  55772=>"001101001",
  55773=>"101111111",
  55774=>"011111011",
  55775=>"111100101",
  55776=>"100010010",
  55777=>"111111111",
  55778=>"010000011",
  55779=>"001000110",
  55780=>"010000100",
  55781=>"111111100",
  55782=>"000111000",
  55783=>"100001110",
  55784=>"010011000",
  55785=>"100110101",
  55786=>"100000100",
  55787=>"100000101",
  55788=>"010011111",
  55789=>"010011001",
  55790=>"110000000",
  55791=>"000011011",
  55792=>"010101000",
  55793=>"100100110",
  55794=>"011010101",
  55795=>"100100110",
  55796=>"100110110",
  55797=>"111000001",
  55798=>"000000000",
  55799=>"111100000",
  55800=>"000101101",
  55801=>"111101011",
  55802=>"000100111",
  55803=>"000000101",
  55804=>"000000011",
  55805=>"011000011",
  55806=>"010110010",
  55807=>"110000000",
  55808=>"110110110",
  55809=>"111111100",
  55810=>"111100000",
  55811=>"000011110",
  55812=>"111111111",
  55813=>"111011111",
  55814=>"001000010",
  55815=>"100111111",
  55816=>"000001001",
  55817=>"010000000",
  55818=>"111111110",
  55819=>"100101010",
  55820=>"000000000",
  55821=>"000000111",
  55822=>"001110001",
  55823=>"000000000",
  55824=>"000100000",
  55825=>"111111000",
  55826=>"110000000",
  55827=>"000011000",
  55828=>"011111111",
  55829=>"101100000",
  55830=>"111111110",
  55831=>"111111001",
  55832=>"100100001",
  55833=>"010001001",
  55834=>"101101111",
  55835=>"111111111",
  55836=>"111111111",
  55837=>"011111111",
  55838=>"000101011",
  55839=>"000101111",
  55840=>"111111110",
  55841=>"000111111",
  55842=>"000000000",
  55843=>"011111010",
  55844=>"100110100",
  55845=>"000000001",
  55846=>"111111111",
  55847=>"010111010",
  55848=>"111111100",
  55849=>"111111111",
  55850=>"000000000",
  55851=>"000000000",
  55852=>"100110101",
  55853=>"000000000",
  55854=>"111111000",
  55855=>"001010111",
  55856=>"111101111",
  55857=>"111111101",
  55858=>"100000000",
  55859=>"111111111",
  55860=>"111111110",
  55861=>"000101000",
  55862=>"000000110",
  55863=>"000000101",
  55864=>"010110000",
  55865=>"000000000",
  55866=>"000100111",
  55867=>"111111111",
  55868=>"100000000",
  55869=>"111011001",
  55870=>"111000000",
  55871=>"000001100",
  55872=>"111111111",
  55873=>"000000000",
  55874=>"000011110",
  55875=>"100111111",
  55876=>"000000100",
  55877=>"000001011",
  55878=>"111111111",
  55879=>"000000000",
  55880=>"000000000",
  55881=>"010110000",
  55882=>"001000001",
  55883=>"000000001",
  55884=>"000000000",
  55885=>"011111111",
  55886=>"110111111",
  55887=>"111111111",
  55888=>"000101111",
  55889=>"111010111",
  55890=>"000011001",
  55891=>"110000100",
  55892=>"111111110",
  55893=>"000001000",
  55894=>"111111110",
  55895=>"110110010",
  55896=>"111101101",
  55897=>"001001011",
  55898=>"010011011",
  55899=>"000000000",
  55900=>"000010000",
  55901=>"111000100",
  55902=>"111111100",
  55903=>"111011010",
  55904=>"000111111",
  55905=>"100001000",
  55906=>"110111110",
  55907=>"110111110",
  55908=>"000000000",
  55909=>"111001100",
  55910=>"000000010",
  55911=>"111111111",
  55912=>"110000000",
  55913=>"000000111",
  55914=>"010001000",
  55915=>"000000001",
  55916=>"111111110",
  55917=>"000000000",
  55918=>"000000111",
  55919=>"111000110",
  55920=>"010010111",
  55921=>"000000000",
  55922=>"000000111",
  55923=>"010000001",
  55924=>"000010000",
  55925=>"100001111",
  55926=>"000110000",
  55927=>"000001011",
  55928=>"111111101",
  55929=>"101100000",
  55930=>"000011110",
  55931=>"000000001",
  55932=>"111011011",
  55933=>"001000011",
  55934=>"111011101",
  55935=>"000000000",
  55936=>"011001000",
  55937=>"111000000",
  55938=>"000011110",
  55939=>"010111111",
  55940=>"000000000",
  55941=>"111101100",
  55942=>"000000001",
  55943=>"000000000",
  55944=>"000101011",
  55945=>"111000111",
  55946=>"111111111",
  55947=>"001011111",
  55948=>"001000000",
  55949=>"000011001",
  55950=>"011011011",
  55951=>"000001001",
  55952=>"000110110",
  55953=>"111000000",
  55954=>"000000000",
  55955=>"111101101",
  55956=>"000001011",
  55957=>"000000000",
  55958=>"000111001",
  55959=>"110010110",
  55960=>"000101110",
  55961=>"000000110",
  55962=>"111101010",
  55963=>"111010001",
  55964=>"011011001",
  55965=>"100100000",
  55966=>"010010010",
  55967=>"111111010",
  55968=>"000000000",
  55969=>"111010111",
  55970=>"111011001",
  55971=>"000000000",
  55972=>"010011111",
  55973=>"000010011",
  55974=>"111011111",
  55975=>"000000100",
  55976=>"111111100",
  55977=>"000100111",
  55978=>"000000100",
  55979=>"101111101",
  55980=>"001000111",
  55981=>"000000010",
  55982=>"011001011",
  55983=>"000000001",
  55984=>"000110100",
  55985=>"000000000",
  55986=>"010011001",
  55987=>"100100000",
  55988=>"110111110",
  55989=>"110011011",
  55990=>"111111111",
  55991=>"111111000",
  55992=>"000000000",
  55993=>"000100100",
  55994=>"000000011",
  55995=>"101101111",
  55996=>"111111000",
  55997=>"000000000",
  55998=>"000001111",
  55999=>"111100111",
  56000=>"000000000",
  56001=>"011000001",
  56002=>"000011010",
  56003=>"000101100",
  56004=>"000000000",
  56005=>"000011000",
  56006=>"000000000",
  56007=>"111101000",
  56008=>"111101111",
  56009=>"111111111",
  56010=>"111111111",
  56011=>"010111000",
  56012=>"000000000",
  56013=>"001011100",
  56014=>"011011111",
  56015=>"110111011",
  56016=>"110000000",
  56017=>"010011111",
  56018=>"010000001",
  56019=>"100111100",
  56020=>"000000000",
  56021=>"111110011",
  56022=>"111111010",
  56023=>"110111111",
  56024=>"111111000",
  56025=>"001111111",
  56026=>"000000001",
  56027=>"110000110",
  56028=>"110101001",
  56029=>"000101111",
  56030=>"111111111",
  56031=>"000000100",
  56032=>"010110000",
  56033=>"101111110",
  56034=>"000000000",
  56035=>"111110100",
  56036=>"000010000",
  56037=>"000001000",
  56038=>"110101011",
  56039=>"110000000",
  56040=>"000111111",
  56041=>"111111111",
  56042=>"101111000",
  56043=>"000001001",
  56044=>"001111111",
  56045=>"110001000",
  56046=>"111000000",
  56047=>"111111000",
  56048=>"111101001",
  56049=>"100000000",
  56050=>"111011011",
  56051=>"110000000",
  56052=>"000001001",
  56053=>"111111111",
  56054=>"100000000",
  56055=>"000000010",
  56056=>"000000000",
  56057=>"111110000",
  56058=>"000000000",
  56059=>"111110100",
  56060=>"111000000",
  56061=>"110000000",
  56062=>"000001000",
  56063=>"111111110",
  56064=>"001100011",
  56065=>"111111101",
  56066=>"000110111",
  56067=>"100111111",
  56068=>"000111011",
  56069=>"000000000",
  56070=>"011101111",
  56071=>"010111011",
  56072=>"100111111",
  56073=>"111111100",
  56074=>"111100000",
  56075=>"000000000",
  56076=>"000000111",
  56077=>"010010000",
  56078=>"000001101",
  56079=>"111111000",
  56080=>"111000000",
  56081=>"111111111",
  56082=>"001010111",
  56083=>"001010001",
  56084=>"111100111",
  56085=>"000101000",
  56086=>"110011011",
  56087=>"111111101",
  56088=>"101000000",
  56089=>"111100100",
  56090=>"111111101",
  56091=>"000111010",
  56092=>"111111000",
  56093=>"101111000",
  56094=>"000000000",
  56095=>"000000111",
  56096=>"101000000",
  56097=>"010000001",
  56098=>"011101101",
  56099=>"111111000",
  56100=>"111110000",
  56101=>"100100100",
  56102=>"111001000",
  56103=>"110111111",
  56104=>"111001101",
  56105=>"010000000",
  56106=>"110000000",
  56107=>"101000110",
  56108=>"101110101",
  56109=>"001010111",
  56110=>"101000110",
  56111=>"000000011",
  56112=>"111000000",
  56113=>"001111110",
  56114=>"000101101",
  56115=>"000001000",
  56116=>"010000000",
  56117=>"011010110",
  56118=>"111100100",
  56119=>"000010110",
  56120=>"100001000",
  56121=>"000100111",
  56122=>"001011111",
  56123=>"111000001",
  56124=>"000100110",
  56125=>"111001000",
  56126=>"000000010",
  56127=>"111011110",
  56128=>"001000111",
  56129=>"101101001",
  56130=>"111100111",
  56131=>"000000011",
  56132=>"000001111",
  56133=>"000111111",
  56134=>"111101111",
  56135=>"110000111",
  56136=>"100111001",
  56137=>"010101000",
  56138=>"111010111",
  56139=>"111111010",
  56140=>"000111111",
  56141=>"100011010",
  56142=>"100111111",
  56143=>"000000011",
  56144=>"000100111",
  56145=>"111101000",
  56146=>"101111101",
  56147=>"001001001",
  56148=>"000000101",
  56149=>"100110010",
  56150=>"111100011",
  56151=>"111101000",
  56152=>"000000011",
  56153=>"011111100",
  56154=>"000110110",
  56155=>"111100000",
  56156=>"111001000",
  56157=>"001110110",
  56158=>"111010011",
  56159=>"000001100",
  56160=>"111101111",
  56161=>"000010111",
  56162=>"000101111",
  56163=>"000001111",
  56164=>"000000010",
  56165=>"011111001",
  56166=>"010001010",
  56167=>"000111101",
  56168=>"110100111",
  56169=>"011000000",
  56170=>"111110101",
  56171=>"010000101",
  56172=>"110111111",
  56173=>"101000000",
  56174=>"011100000",
  56175=>"001111010",
  56176=>"110011011",
  56177=>"010000101",
  56178=>"111001001",
  56179=>"000000111",
  56180=>"111110111",
  56181=>"101111111",
  56182=>"111101000",
  56183=>"000000110",
  56184=>"000000011",
  56185=>"000000000",
  56186=>"111111000",
  56187=>"000000011",
  56188=>"000000001",
  56189=>"100001110",
  56190=>"111000000",
  56191=>"000000001",
  56192=>"111000000",
  56193=>"000001010",
  56194=>"111111010",
  56195=>"111001011",
  56196=>"101111111",
  56197=>"100000000",
  56198=>"101101111",
  56199=>"001000010",
  56200=>"011110110",
  56201=>"000111011",
  56202=>"011000111",
  56203=>"000000101",
  56204=>"000000111",
  56205=>"001010111",
  56206=>"101101010",
  56207=>"001001101",
  56208=>"011111110",
  56209=>"111000000",
  56210=>"111010000",
  56211=>"000000000",
  56212=>"000101000",
  56213=>"100001000",
  56214=>"000111111",
  56215=>"101111000",
  56216=>"111000000",
  56217=>"011001101",
  56218=>"111000000",
  56219=>"001000000",
  56220=>"000000001",
  56221=>"000000111",
  56222=>"111001101",
  56223=>"000001001",
  56224=>"001111000",
  56225=>"000000111",
  56226=>"001000000",
  56227=>"011001101",
  56228=>"000010000",
  56229=>"101001011",
  56230=>"110110110",
  56231=>"010101000",
  56232=>"111110111",
  56233=>"000110001",
  56234=>"000000000",
  56235=>"111110100",
  56236=>"010000110",
  56237=>"000000111",
  56238=>"110100101",
  56239=>"000000101",
  56240=>"111000111",
  56241=>"001001010",
  56242=>"000110111",
  56243=>"000001001",
  56244=>"000100101",
  56245=>"111001000",
  56246=>"111100100",
  56247=>"000000000",
  56248=>"000011010",
  56249=>"000001100",
  56250=>"101000010",
  56251=>"000000001",
  56252=>"010001001",
  56253=>"000101111",
  56254=>"101100010",
  56255=>"010000110",
  56256=>"000000101",
  56257=>"111000000",
  56258=>"010100101",
  56259=>"001011010",
  56260=>"000010111",
  56261=>"100110011",
  56262=>"111101000",
  56263=>"010000000",
  56264=>"000101000",
  56265=>"111100110",
  56266=>"111001000",
  56267=>"111110111",
  56268=>"000100111",
  56269=>"011110000",
  56270=>"000101000",
  56271=>"110000001",
  56272=>"000111111",
  56273=>"001110111",
  56274=>"100000000",
  56275=>"110111001",
  56276=>"000000100",
  56277=>"100001010",
  56278=>"000011111",
  56279=>"111111101",
  56280=>"001000000",
  56281=>"000110001",
  56282=>"110110010",
  56283=>"010101111",
  56284=>"001110110",
  56285=>"101100111",
  56286=>"111101101",
  56287=>"000000101",
  56288=>"000100111",
  56289=>"000101011",
  56290=>"001001001",
  56291=>"111011011",
  56292=>"000000000",
  56293=>"101101111",
  56294=>"001111111",
  56295=>"111101110",
  56296=>"000011001",
  56297=>"010010000",
  56298=>"011011100",
  56299=>"110001000",
  56300=>"111111100",
  56301=>"100010000",
  56302=>"010000000",
  56303=>"101000000",
  56304=>"100000000",
  56305=>"011011111",
  56306=>"000010101",
  56307=>"100011111",
  56308=>"111011111",
  56309=>"001101000",
  56310=>"000000000",
  56311=>"011101111",
  56312=>"111000000",
  56313=>"111000001",
  56314=>"111000010",
  56315=>"000110111",
  56316=>"110110010",
  56317=>"001000100",
  56318=>"001110110",
  56319=>"001110011",
  56320=>"111011100",
  56321=>"000100111",
  56322=>"100000100",
  56323=>"000000010",
  56324=>"000011011",
  56325=>"111000111",
  56326=>"011011010",
  56327=>"000110111",
  56328=>"010010000",
  56329=>"010111000",
  56330=>"110011111",
  56331=>"000000110",
  56332=>"100100101",
  56333=>"011011010",
  56334=>"101011001",
  56335=>"000000000",
  56336=>"110101111",
  56337=>"110011110",
  56338=>"000010100",
  56339=>"000111111",
  56340=>"111011101",
  56341=>"010100100",
  56342=>"000100011",
  56343=>"000010000",
  56344=>"000011000",
  56345=>"010010000",
  56346=>"000100101",
  56347=>"111111110",
  56348=>"111111000",
  56349=>"111011000",
  56350=>"101111010",
  56351=>"000110100",
  56352=>"000000111",
  56353=>"000010000",
  56354=>"001110101",
  56355=>"000101010",
  56356=>"000001000",
  56357=>"110010000",
  56358=>"000100100",
  56359=>"000000010",
  56360=>"101100111",
  56361=>"010011011",
  56362=>"111111011",
  56363=>"111100100",
  56364=>"111111011",
  56365=>"001000111",
  56366=>"111100111",
  56367=>"010011110",
  56368=>"001010111",
  56369=>"001001001",
  56370=>"101001110",
  56371=>"011110111",
  56372=>"011111010",
  56373=>"111111110",
  56374=>"111111111",
  56375=>"111111110",
  56376=>"011111111",
  56377=>"000011000",
  56378=>"010110111",
  56379=>"000111000",
  56380=>"100100001",
  56381=>"111111001",
  56382=>"000000010",
  56383=>"101111111",
  56384=>"000000000",
  56385=>"010000010",
  56386=>"101100111",
  56387=>"001100110",
  56388=>"010011000",
  56389=>"000000101",
  56390=>"001011000",
  56391=>"101001000",
  56392=>"000001111",
  56393=>"100100111",
  56394=>"101100101",
  56395=>"100100000",
  56396=>"000111010",
  56397=>"001101101",
  56398=>"100110110",
  56399=>"011010010",
  56400=>"010011011",
  56401=>"000101111",
  56402=>"101111000",
  56403=>"011000011",
  56404=>"111101101",
  56405=>"001111011",
  56406=>"100110110",
  56407=>"001000000",
  56408=>"100110111",
  56409=>"000001001",
  56410=>"001111011",
  56411=>"110110100",
  56412=>"100000111",
  56413=>"001001001",
  56414=>"111111000",
  56415=>"110100101",
  56416=>"000100100",
  56417=>"100000101",
  56418=>"100100000",
  56419=>"110110110",
  56420=>"010011001",
  56421=>"011011111",
  56422=>"111111111",
  56423=>"010011000",
  56424=>"010010010",
  56425=>"000000000",
  56426=>"110101100",
  56427=>"111000000",
  56428=>"000000011",
  56429=>"011000000",
  56430=>"100100000",
  56431=>"111000011",
  56432=>"011001001",
  56433=>"000000111",
  56434=>"111111111",
  56435=>"100000000",
  56436=>"111000000",
  56437=>"100101110",
  56438=>"111111111",
  56439=>"111000000",
  56440=>"000000011",
  56441=>"010000000",
  56442=>"111101000",
  56443=>"010011110",
  56444=>"100110001",
  56445=>"010000100",
  56446=>"111100111",
  56447=>"110111111",
  56448=>"101000000",
  56449=>"111100110",
  56450=>"011011010",
  56451=>"111011010",
  56452=>"011100000",
  56453=>"111011010",
  56454=>"011001000",
  56455=>"100001000",
  56456=>"000111110",
  56457=>"000000000",
  56458=>"000000100",
  56459=>"111000100",
  56460=>"000000000",
  56461=>"000100111",
  56462=>"101001001",
  56463=>"101000001",
  56464=>"111111101",
  56465=>"010011101",
  56466=>"011010000",
  56467=>"000100011",
  56468=>"000010011",
  56469=>"111000001",
  56470=>"101001000",
  56471=>"000000001",
  56472=>"000010010",
  56473=>"000100111",
  56474=>"100100100",
  56475=>"001100000",
  56476=>"000100011",
  56477=>"001100000",
  56478=>"000000111",
  56479=>"101111111",
  56480=>"000100000",
  56481=>"000000011",
  56482=>"110000101",
  56483=>"111011010",
  56484=>"010010111",
  56485=>"000000010",
  56486=>"001000011",
  56487=>"001011000",
  56488=>"111000111",
  56489=>"000100000",
  56490=>"000000110",
  56491=>"111000000",
  56492=>"111111001",
  56493=>"011111000",
  56494=>"110110110",
  56495=>"111000111",
  56496=>"010000111",
  56497=>"001100100",
  56498=>"110110000",
  56499=>"000110010",
  56500=>"101111110",
  56501=>"010000000",
  56502=>"011000100",
  56503=>"111000011",
  56504=>"001000100",
  56505=>"000110110",
  56506=>"111011000",
  56507=>"111011010",
  56508=>"010000000",
  56509=>"110111001",
  56510=>"110110100",
  56511=>"000000011",
  56512=>"000000000",
  56513=>"100101100",
  56514=>"111000000",
  56515=>"001011001",
  56516=>"111000001",
  56517=>"100111101",
  56518=>"000011011",
  56519=>"110100100",
  56520=>"010100011",
  56521=>"000100000",
  56522=>"000000000",
  56523=>"100100111",
  56524=>"010011011",
  56525=>"001011010",
  56526=>"111111011",
  56527=>"101000110",
  56528=>"110011010",
  56529=>"101000110",
  56530=>"000000000",
  56531=>"100100101",
  56532=>"111101101",
  56533=>"000000000",
  56534=>"000011011",
  56535=>"111010000",
  56536=>"100100101",
  56537=>"011000100",
  56538=>"010000100",
  56539=>"101100100",
  56540=>"011111111",
  56541=>"001010011",
  56542=>"100000000",
  56543=>"000001111",
  56544=>"110000000",
  56545=>"101100111",
  56546=>"111100100",
  56547=>"000000000",
  56548=>"000000000",
  56549=>"011111000",
  56550=>"010000010",
  56551=>"010100110",
  56552=>"110000111",
  56553=>"000000000",
  56554=>"111011011",
  56555=>"100111000",
  56556=>"100100101",
  56557=>"101000100",
  56558=>"110100000",
  56559=>"010101010",
  56560=>"000000000",
  56561=>"011001110",
  56562=>"101100000",
  56563=>"011111000",
  56564=>"010000011",
  56565=>"000011000",
  56566=>"000010010",
  56567=>"011101100",
  56568=>"111100111",
  56569=>"000011111",
  56570=>"000000000",
  56571=>"110100000",
  56572=>"000000000",
  56573=>"100100000",
  56574=>"110110100",
  56575=>"100000100",
  56576=>"010001000",
  56577=>"000101111",
  56578=>"111000000",
  56579=>"000110110",
  56580=>"100110100",
  56581=>"101011010",
  56582=>"111100000",
  56583=>"101010101",
  56584=>"010011001",
  56585=>"010111010",
  56586=>"011111101",
  56587=>"000000000",
  56588=>"011101101",
  56589=>"000000001",
  56590=>"000000101",
  56591=>"000000000",
  56592=>"111111000",
  56593=>"101000000",
  56594=>"010111010",
  56595=>"000111000",
  56596=>"111111111",
  56597=>"010000100",
  56598=>"000000011",
  56599=>"111111010",
  56600=>"111101001",
  56601=>"011000000",
  56602=>"100000000",
  56603=>"100100101",
  56604=>"110000000",
  56605=>"111111111",
  56606=>"010000000",
  56607=>"000000000",
  56608=>"111100000",
  56609=>"000000101",
  56610=>"000000000",
  56611=>"000010011",
  56612=>"111110110",
  56613=>"010010001",
  56614=>"000110000",
  56615=>"100101001",
  56616=>"101001110",
  56617=>"111101001",
  56618=>"110101100",
  56619=>"010111111",
  56620=>"111111011",
  56621=>"010000101",
  56622=>"100010011",
  56623=>"010010111",
  56624=>"101011000",
  56625=>"001010010",
  56626=>"111100000",
  56627=>"100000101",
  56628=>"111000000",
  56629=>"010110001",
  56630=>"000010011",
  56631=>"010110100",
  56632=>"101111100",
  56633=>"101101111",
  56634=>"000010010",
  56635=>"111010010",
  56636=>"000111001",
  56637=>"111111111",
  56638=>"100000000",
  56639=>"011011011",
  56640=>"000000111",
  56641=>"000110011",
  56642=>"010010100",
  56643=>"000111011",
  56644=>"110101010",
  56645=>"010000000",
  56646=>"110010110",
  56647=>"111111110",
  56648=>"101000000",
  56649=>"000010010",
  56650=>"111101111",
  56651=>"100011011",
  56652=>"111100100",
  56653=>"111110011",
  56654=>"100110001",
  56655=>"111111111",
  56656=>"111111011",
  56657=>"111110111",
  56658=>"101010011",
  56659=>"110001001",
  56660=>"000000000",
  56661=>"100100111",
  56662=>"101111011",
  56663=>"101111000",
  56664=>"001000101",
  56665=>"001011111",
  56666=>"000100100",
  56667=>"011011001",
  56668=>"000000111",
  56669=>"100000000",
  56670=>"101000000",
  56671=>"001111110",
  56672=>"000000001",
  56673=>"000011011",
  56674=>"000000110",
  56675=>"110111001",
  56676=>"000100101",
  56677=>"110100100",
  56678=>"101111111",
  56679=>"000111001",
  56680=>"110011000",
  56681=>"111110111",
  56682=>"111111111",
  56683=>"100011010",
  56684=>"101110111",
  56685=>"111000000",
  56686=>"000011000",
  56687=>"111000000",
  56688=>"100111110",
  56689=>"100110111",
  56690=>"000011011",
  56691=>"101000000",
  56692=>"111111000",
  56693=>"110000000",
  56694=>"000000100",
  56695=>"111111011",
  56696=>"000110000",
  56697=>"100100010",
  56698=>"111101001",
  56699=>"001011111",
  56700=>"001110011",
  56701=>"100100110",
  56702=>"100110000",
  56703=>"010011011",
  56704=>"001100000",
  56705=>"111111111",
  56706=>"101011010",
  56707=>"000111111",
  56708=>"010110101",
  56709=>"111111010",
  56710=>"000010100",
  56711=>"000001000",
  56712=>"001011011",
  56713=>"101001000",
  56714=>"001100000",
  56715=>"100000000",
  56716=>"111000100",
  56717=>"100111001",
  56718=>"000010110",
  56719=>"100000100",
  56720=>"011011001",
  56721=>"000001011",
  56722=>"011011010",
  56723=>"001000010",
  56724=>"100001110",
  56725=>"011111101",
  56726=>"111100100",
  56727=>"010110100",
  56728=>"111111111",
  56729=>"100011010",
  56730=>"011111111",
  56731=>"111011000",
  56732=>"111100000",
  56733=>"000000000",
  56734=>"110110000",
  56735=>"111100101",
  56736=>"011011011",
  56737=>"011010000",
  56738=>"110110000",
  56739=>"100000100",
  56740=>"100111110",
  56741=>"011110110",
  56742=>"010000110",
  56743=>"000010001",
  56744=>"001000000",
  56745=>"001100000",
  56746=>"101101111",
  56747=>"100100101",
  56748=>"000000111",
  56749=>"000100111",
  56750=>"100111000",
  56751=>"001111111",
  56752=>"100111011",
  56753=>"100100000",
  56754=>"111010011",
  56755=>"000000001",
  56756=>"010010111",
  56757=>"000000000",
  56758=>"011100100",
  56759=>"000000000",
  56760=>"011111010",
  56761=>"001100000",
  56762=>"100101111",
  56763=>"111001000",
  56764=>"001100001",
  56765=>"111000000",
  56766=>"110110110",
  56767=>"000111111",
  56768=>"011011010",
  56769=>"000111110",
  56770=>"011000000",
  56771=>"110111101",
  56772=>"101100010",
  56773=>"111100000",
  56774=>"000111111",
  56775=>"100000100",
  56776=>"001000000",
  56777=>"010111010",
  56778=>"100000010",
  56779=>"000111110",
  56780=>"000011000",
  56781=>"100100001",
  56782=>"011111000",
  56783=>"000110111",
  56784=>"011111010",
  56785=>"011000001",
  56786=>"100100000",
  56787=>"100111111",
  56788=>"110010111",
  56789=>"101001000",
  56790=>"101100101",
  56791=>"000100011",
  56792=>"111111111",
  56793=>"111011011",
  56794=>"110011011",
  56795=>"111000100",
  56796=>"000000011",
  56797=>"001111110",
  56798=>"100100110",
  56799=>"101101111",
  56800=>"010011011",
  56801=>"101100001",
  56802=>"001111011",
  56803=>"000100001",
  56804=>"000000000",
  56805=>"000000000",
  56806=>"111110010",
  56807=>"001111101",
  56808=>"110111111",
  56809=>"101111001",
  56810=>"101101010",
  56811=>"111000001",
  56812=>"111100100",
  56813=>"000100011",
  56814=>"111001010",
  56815=>"010000010",
  56816=>"101111000",
  56817=>"110100100",
  56818=>"001011011",
  56819=>"010110110",
  56820=>"100001100",
  56821=>"000000011",
  56822=>"111100010",
  56823=>"000011110",
  56824=>"110111000",
  56825=>"111111100",
  56826=>"011011110",
  56827=>"110000010",
  56828=>"111111111",
  56829=>"000110010",
  56830=>"001011001",
  56831=>"000000101",
  56832=>"010000000",
  56833=>"000010010",
  56834=>"000000001",
  56835=>"001001111",
  56836=>"000000000",
  56837=>"001001101",
  56838=>"000000000",
  56839=>"101010111",
  56840=>"000000000",
  56841=>"000000000",
  56842=>"111111011",
  56843=>"101001101",
  56844=>"000000000",
  56845=>"101001000",
  56846=>"010000001",
  56847=>"001111111",
  56848=>"000010011",
  56849=>"010010010",
  56850=>"110110110",
  56851=>"000110111",
  56852=>"010101111",
  56853=>"000011010",
  56854=>"111100000",
  56855=>"110110010",
  56856=>"010000000",
  56857=>"011111111",
  56858=>"000001111",
  56859=>"000000100",
  56860=>"000101110",
  56861=>"101000010",
  56862=>"010011100",
  56863=>"000101001",
  56864=>"001001111",
  56865=>"111100001",
  56866=>"011100000",
  56867=>"001101111",
  56868=>"111101110",
  56869=>"001001011",
  56870=>"000111010",
  56871=>"000000000",
  56872=>"010111111",
  56873=>"010011011",
  56874=>"111110111",
  56875=>"011111010",
  56876=>"111111111",
  56877=>"011001111",
  56878=>"111111011",
  56879=>"001000000",
  56880=>"111101001",
  56881=>"100101011",
  56882=>"010111110",
  56883=>"111111111",
  56884=>"011010000",
  56885=>"010001000",
  56886=>"111110011",
  56887=>"000000000",
  56888=>"011111111",
  56889=>"000000011",
  56890=>"000000000",
  56891=>"110000111",
  56892=>"111100111",
  56893=>"111111010",
  56894=>"000000001",
  56895=>"001000100",
  56896=>"111111111",
  56897=>"110010010",
  56898=>"111111111",
  56899=>"000000000",
  56900=>"110111111",
  56901=>"000000000",
  56902=>"000001101",
  56903=>"110110111",
  56904=>"000100011",
  56905=>"101000101",
  56906=>"111111111",
  56907=>"100110010",
  56908=>"101000000",
  56909=>"111011011",
  56910=>"111101110",
  56911=>"010111111",
  56912=>"000001000",
  56913=>"111010000",
  56914=>"101101111",
  56915=>"011000000",
  56916=>"000000000",
  56917=>"000000100",
  56918=>"001001000",
  56919=>"000010110",
  56920=>"000000000",
  56921=>"000100111",
  56922=>"100100000",
  56923=>"001011001",
  56924=>"111001101",
  56925=>"100100101",
  56926=>"010110111",
  56927=>"000000001",
  56928=>"111000000",
  56929=>"001000101",
  56930=>"000000001",
  56931=>"111111101",
  56932=>"101101000",
  56933=>"101000000",
  56934=>"111101010",
  56935=>"000110011",
  56936=>"111001000",
  56937=>"111111111",
  56938=>"000000000",
  56939=>"010111001",
  56940=>"111110111",
  56941=>"010110111",
  56942=>"000000000",
  56943=>"000100010",
  56944=>"100100000",
  56945=>"110111010",
  56946=>"111010110",
  56947=>"000110010",
  56948=>"000000111",
  56949=>"000101101",
  56950=>"011011110",
  56951=>"000000001",
  56952=>"010011101",
  56953=>"000001111",
  56954=>"111000010",
  56955=>"111101100",
  56956=>"111000011",
  56957=>"111001101",
  56958=>"110000000",
  56959=>"000000000",
  56960=>"111000000",
  56961=>"000110110",
  56962=>"010001011",
  56963=>"101101100",
  56964=>"010000101",
  56965=>"101000000",
  56966=>"010111010",
  56967=>"110001111",
  56968=>"011011111",
  56969=>"111101000",
  56970=>"000000000",
  56971=>"010110111",
  56972=>"000000000",
  56973=>"000101111",
  56974=>"010000000",
  56975=>"000110100",
  56976=>"011011011",
  56977=>"000000001",
  56978=>"000000010",
  56979=>"111001111",
  56980=>"100100010",
  56981=>"000000111",
  56982=>"010110010",
  56983=>"100111111",
  56984=>"101001000",
  56985=>"110110101",
  56986=>"000111010",
  56987=>"001000000",
  56988=>"100100000",
  56989=>"101001000",
  56990=>"000111110",
  56991=>"100000000",
  56992=>"010000010",
  56993=>"101000111",
  56994=>"000111111",
  56995=>"111110100",
  56996=>"011000000",
  56997=>"100110110",
  56998=>"000010101",
  56999=>"111111111",
  57000=>"010000110",
  57001=>"111110111",
  57002=>"001000000",
  57003=>"000000000",
  57004=>"110001000",
  57005=>"000001011",
  57006=>"000001001",
  57007=>"111111111",
  57008=>"000000010",
  57009=>"010110100",
  57010=>"000000000",
  57011=>"001100100",
  57012=>"001111111",
  57013=>"111101101",
  57014=>"000011111",
  57015=>"010111111",
  57016=>"110101111",
  57017=>"111101011",
  57018=>"101001001",
  57019=>"110111010",
  57020=>"110111111",
  57021=>"000010000",
  57022=>"000000001",
  57023=>"000001101",
  57024=>"010110000",
  57025=>"000000000",
  57026=>"101010010",
  57027=>"111100100",
  57028=>"100110011",
  57029=>"010001010",
  57030=>"110000101",
  57031=>"101000100",
  57032=>"111101111",
  57033=>"110111100",
  57034=>"010111000",
  57035=>"011001000",
  57036=>"111010010",
  57037=>"111100100",
  57038=>"000000100",
  57039=>"111100001",
  57040=>"000000111",
  57041=>"111100110",
  57042=>"000111100",
  57043=>"000001111",
  57044=>"000000000",
  57045=>"000010010",
  57046=>"000000000",
  57047=>"000000010",
  57048=>"011111111",
  57049=>"010111101",
  57050=>"111000111",
  57051=>"001001000",
  57052=>"100011011",
  57053=>"101110111",
  57054=>"001111111",
  57055=>"000000110",
  57056=>"111000101",
  57057=>"001011111",
  57058=>"000010010",
  57059=>"101110110",
  57060=>"000000000",
  57061=>"001000000",
  57062=>"111001111",
  57063=>"011000100",
  57064=>"011001111",
  57065=>"000101111",
  57066=>"111110110",
  57067=>"000110000",
  57068=>"100101101",
  57069=>"000111111",
  57070=>"000110110",
  57071=>"101001110",
  57072=>"111101111",
  57073=>"001110101",
  57074=>"000000000",
  57075=>"001000011",
  57076=>"111100011",
  57077=>"001111000",
  57078=>"001101010",
  57079=>"111111111",
  57080=>"000010111",
  57081=>"000111111",
  57082=>"010111111",
  57083=>"111111001",
  57084=>"000010000",
  57085=>"001001101",
  57086=>"000100100",
  57087=>"001011001",
  57088=>"101000110",
  57089=>"000010111",
  57090=>"000011010",
  57091=>"111010111",
  57092=>"001001000",
  57093=>"110110111",
  57094=>"101101001",
  57095=>"111010111",
  57096=>"001101101",
  57097=>"011000000",
  57098=>"100000000",
  57099=>"000000010",
  57100=>"000011000",
  57101=>"010110000",
  57102=>"100011100",
  57103=>"111110101",
  57104=>"011100000",
  57105=>"010010010",
  57106=>"100100110",
  57107=>"100110001",
  57108=>"100011000",
  57109=>"000010111",
  57110=>"110111111",
  57111=>"110100111",
  57112=>"010110000",
  57113=>"101111111",
  57114=>"111011101",
  57115=>"111000111",
  57116=>"111111111",
  57117=>"110000011",
  57118=>"111010011",
  57119=>"101101111",
  57120=>"101111100",
  57121=>"000000111",
  57122=>"000000001",
  57123=>"111111000",
  57124=>"000101101",
  57125=>"100000011",
  57126=>"111111101",
  57127=>"111111100",
  57128=>"001111111",
  57129=>"000010001",
  57130=>"010000000",
  57131=>"100111111",
  57132=>"001001101",
  57133=>"000000001",
  57134=>"111111000",
  57135=>"000100000",
  57136=>"000000011",
  57137=>"000001000",
  57138=>"000010111",
  57139=>"111000010",
  57140=>"101011010",
  57141=>"000000000",
  57142=>"000000100",
  57143=>"011001000",
  57144=>"110010100",
  57145=>"000000000",
  57146=>"111101111",
  57147=>"101011000",
  57148=>"101111011",
  57149=>"101111101",
  57150=>"000000000",
  57151=>"011000000",
  57152=>"001000111",
  57153=>"010110100",
  57154=>"010111101",
  57155=>"010011001",
  57156=>"110000010",
  57157=>"000000011",
  57158=>"010111000",
  57159=>"111111000",
  57160=>"000000111",
  57161=>"111110000",
  57162=>"000100000",
  57163=>"111101010",
  57164=>"100100101",
  57165=>"010101100",
  57166=>"100100001",
  57167=>"101111000",
  57168=>"000111101",
  57169=>"000000000",
  57170=>"110011010",
  57171=>"101001001",
  57172=>"000010110",
  57173=>"001000101",
  57174=>"100001000",
  57175=>"011010010",
  57176=>"011001001",
  57177=>"111001000",
  57178=>"000110101",
  57179=>"010100000",
  57180=>"110010000",
  57181=>"001001101",
  57182=>"110000111",
  57183=>"001000100",
  57184=>"001111111",
  57185=>"111101110",
  57186=>"110100100",
  57187=>"100101101",
  57188=>"111101000",
  57189=>"111101101",
  57190=>"110111100",
  57191=>"110111000",
  57192=>"101000111",
  57193=>"111010010",
  57194=>"111010110",
  57195=>"101111111",
  57196=>"001010000",
  57197=>"111000000",
  57198=>"110100000",
  57199=>"001000010",
  57200=>"100001000",
  57201=>"111010000",
  57202=>"000000011",
  57203=>"111111011",
  57204=>"111010110",
  57205=>"000100011",
  57206=>"010111111",
  57207=>"000110000",
  57208=>"110111010",
  57209=>"111000011",
  57210=>"000000111",
  57211=>"111001000",
  57212=>"000000011",
  57213=>"111100000",
  57214=>"111111111",
  57215=>"101101101",
  57216=>"000010000",
  57217=>"100000111",
  57218=>"111111000",
  57219=>"101001000",
  57220=>"111000000",
  57221=>"111111110",
  57222=>"001001000",
  57223=>"101100100",
  57224=>"000100000",
  57225=>"111111111",
  57226=>"111111100",
  57227=>"101111010",
  57228=>"000101101",
  57229=>"110110111",
  57230=>"010000100",
  57231=>"011011110",
  57232=>"001101001",
  57233=>"000011111",
  57234=>"111000000",
  57235=>"011010010",
  57236=>"011001100",
  57237=>"111010000",
  57238=>"111101111",
  57239=>"100100100",
  57240=>"111000000",
  57241=>"000111111",
  57242=>"100000100",
  57243=>"000000111",
  57244=>"000010111",
  57245=>"111011111",
  57246=>"111010011",
  57247=>"001000000",
  57248=>"000000001",
  57249=>"011000111",
  57250=>"011000000",
  57251=>"100000111",
  57252=>"111110000",
  57253=>"100100000",
  57254=>"001111000",
  57255=>"010011101",
  57256=>"111010000",
  57257=>"000111111",
  57258=>"000100011",
  57259=>"010000000",
  57260=>"011110011",
  57261=>"111111000",
  57262=>"110000110",
  57263=>"111111000",
  57264=>"111000001",
  57265=>"000001001",
  57266=>"000100111",
  57267=>"000000011",
  57268=>"110111101",
  57269=>"000010101",
  57270=>"001000000",
  57271=>"000000101",
  57272=>"101111110",
  57273=>"110111001",
  57274=>"111000010",
  57275=>"111010001",
  57276=>"000011011",
  57277=>"000111111",
  57278=>"111111001",
  57279=>"000010000",
  57280=>"000000010",
  57281=>"000000000",
  57282=>"111111111",
  57283=>"000101001",
  57284=>"010010111",
  57285=>"110110110",
  57286=>"000011000",
  57287=>"111001111",
  57288=>"100000101",
  57289=>"000001101",
  57290=>"001110000",
  57291=>"010110110",
  57292=>"111100000",
  57293=>"000110110",
  57294=>"000011111",
  57295=>"001110111",
  57296=>"000111000",
  57297=>"100100111",
  57298=>"101101010",
  57299=>"111011011",
  57300=>"100111111",
  57301=>"100100111",
  57302=>"000000101",
  57303=>"111000111",
  57304=>"001010010",
  57305=>"101000010",
  57306=>"000100000",
  57307=>"111100101",
  57308=>"000110110",
  57309=>"100111111",
  57310=>"000000010",
  57311=>"111010000",
  57312=>"000101000",
  57313=>"010111111",
  57314=>"111101000",
  57315=>"111101001",
  57316=>"111111011",
  57317=>"000000101",
  57318=>"000011111",
  57319=>"011001000",
  57320=>"111010111",
  57321=>"101111111",
  57322=>"011001011",
  57323=>"000111111",
  57324=>"000000001",
  57325=>"000000000",
  57326=>"000000000",
  57327=>"101101100",
  57328=>"100000010",
  57329=>"011011001",
  57330=>"110111100",
  57331=>"111101001",
  57332=>"101100000",
  57333=>"100101111",
  57334=>"000010111",
  57335=>"101111111",
  57336=>"000000110",
  57337=>"000000010",
  57338=>"101111111",
  57339=>"101111011",
  57340=>"111101100",
  57341=>"000000000",
  57342=>"011000000",
  57343=>"111111000",
  57344=>"100101011",
  57345=>"001000100",
  57346=>"000000111",
  57347=>"000110110",
  57348=>"001000000",
  57349=>"111101001",
  57350=>"011000000",
  57351=>"111111101",
  57352=>"001101111",
  57353=>"000001101",
  57354=>"000000011",
  57355=>"010000111",
  57356=>"111111010",
  57357=>"001111111",
  57358=>"000000000",
  57359=>"011111111",
  57360=>"001101101",
  57361=>"000000000",
  57362=>"111110111",
  57363=>"010000000",
  57364=>"101100110",
  57365=>"000000101",
  57366=>"000000000",
  57367=>"011111111",
  57368=>"111100111",
  57369=>"111111111",
  57370=>"101101111",
  57371=>"010000100",
  57372=>"111000010",
  57373=>"001011000",
  57374=>"000100100",
  57375=>"000000001",
  57376=>"111011111",
  57377=>"001110111",
  57378=>"001011111",
  57379=>"001000000",
  57380=>"000010000",
  57381=>"001001111",
  57382=>"100000001",
  57383=>"000110111",
  57384=>"011010111",
  57385=>"010111111",
  57386=>"001111000",
  57387=>"000000100",
  57388=>"001011110",
  57389=>"011010111",
  57390=>"111101101",
  57391=>"011010000",
  57392=>"001111110",
  57393=>"111101100",
  57394=>"000000000",
  57395=>"000001100",
  57396=>"001000101",
  57397=>"000000000",
  57398=>"000000000",
  57399=>"000100101",
  57400=>"111000000",
  57401=>"000101101",
  57402=>"111010111",
  57403=>"000000000",
  57404=>"011001011",
  57405=>"011011111",
  57406=>"000000101",
  57407=>"000001001",
  57408=>"101111111",
  57409=>"011111010",
  57410=>"101111111",
  57411=>"001000001",
  57412=>"000010000",
  57413=>"101111010",
  57414=>"010101100",
  57415=>"001001110",
  57416=>"111011111",
  57417=>"111111111",
  57418=>"000010111",
  57419=>"101101101",
  57420=>"111111111",
  57421=>"000000110",
  57422=>"110100010",
  57423=>"000000110",
  57424=>"000000000",
  57425=>"110111110",
  57426=>"000000111",
  57427=>"111110001",
  57428=>"001000001",
  57429=>"101101101",
  57430=>"010010000",
  57431=>"000010111",
  57432=>"001101000",
  57433=>"111111111",
  57434=>"000000000",
  57435=>"000100100",
  57436=>"000000011",
  57437=>"100110000",
  57438=>"111111111",
  57439=>"101000000",
  57440=>"100110111",
  57441=>"010000000",
  57442=>"111111111",
  57443=>"001010000",
  57444=>"001000011",
  57445=>"010111000",
  57446=>"111111100",
  57447=>"001101001",
  57448=>"000000010",
  57449=>"111000001",
  57450=>"111001101",
  57451=>"111111010",
  57452=>"011111001",
  57453=>"011000000",
  57454=>"010111000",
  57455=>"001110111",
  57456=>"111100111",
  57457=>"101110111",
  57458=>"000000001",
  57459=>"111111011",
  57460=>"111101000",
  57461=>"101101000",
  57462=>"100000001",
  57463=>"001111100",
  57464=>"000000000",
  57465=>"111001100",
  57466=>"000001101",
  57467=>"111111110",
  57468=>"001001001",
  57469=>"111011010",
  57470=>"111111111",
  57471=>"000100111",
  57472=>"001000000",
  57473=>"000100000",
  57474=>"000111000",
  57475=>"101011000",
  57476=>"000101111",
  57477=>"010001000",
  57478=>"000100010",
  57479=>"010100111",
  57480=>"111000110",
  57481=>"000000001",
  57482=>"101001111",
  57483=>"111011000",
  57484=>"001101111",
  57485=>"000000100",
  57486=>"011111111",
  57487=>"000000000",
  57488=>"110100010",
  57489=>"100001000",
  57490=>"110101001",
  57491=>"011001101",
  57492=>"110100000",
  57493=>"000000000",
  57494=>"111111110",
  57495=>"100111011",
  57496=>"101101010",
  57497=>"000000001",
  57498=>"111111111",
  57499=>"000010011",
  57500=>"010101000",
  57501=>"010111111",
  57502=>"000001111",
  57503=>"010111001",
  57504=>"011110111",
  57505=>"000000001",
  57506=>"111111111",
  57507=>"100111101",
  57508=>"000100101",
  57509=>"000000100",
  57510=>"111110110",
  57511=>"111101000",
  57512=>"000000000",
  57513=>"000000001",
  57514=>"111110000",
  57515=>"000000000",
  57516=>"010111110",
  57517=>"000000111",
  57518=>"000000000",
  57519=>"111111111",
  57520=>"000101111",
  57521=>"100101001",
  57522=>"111000100",
  57523=>"111111011",
  57524=>"111011011",
  57525=>"111110000",
  57526=>"010111110",
  57527=>"111101101",
  57528=>"100100111",
  57529=>"110101111",
  57530=>"101000001",
  57531=>"111111111",
  57532=>"111000011",
  57533=>"111111110",
  57534=>"000101100",
  57535=>"000111111",
  57536=>"000000111",
  57537=>"010000000",
  57538=>"001011010",
  57539=>"011000001",
  57540=>"111111111",
  57541=>"001001001",
  57542=>"000101000",
  57543=>"000100100",
  57544=>"010111111",
  57545=>"000001000",
  57546=>"000000101",
  57547=>"100111111",
  57548=>"000101101",
  57549=>"110000100",
  57550=>"101101001",
  57551=>"101111111",
  57552=>"000000000",
  57553=>"111111000",
  57554=>"111111111",
  57555=>"111111111",
  57556=>"000000000",
  57557=>"001001111",
  57558=>"000111110",
  57559=>"101011000",
  57560=>"111111001",
  57561=>"111111111",
  57562=>"011011010",
  57563=>"000010011",
  57564=>"000000001",
  57565=>"010110101",
  57566=>"111111010",
  57567=>"001101111",
  57568=>"100000001",
  57569=>"001011111",
  57570=>"111011011",
  57571=>"011001001",
  57572=>"000000001",
  57573=>"111111101",
  57574=>"111101001",
  57575=>"000001001",
  57576=>"000000100",
  57577=>"111101111",
  57578=>"000000001",
  57579=>"010010111",
  57580=>"111111010",
  57581=>"000101111",
  57582=>"111111111",
  57583=>"000010100",
  57584=>"110000111",
  57585=>"000000000",
  57586=>"110111111",
  57587=>"000110111",
  57588=>"101101111",
  57589=>"000000000",
  57590=>"101000110",
  57591=>"110111011",
  57592=>"000100100",
  57593=>"000001100",
  57594=>"000110000",
  57595=>"001001001",
  57596=>"000000011",
  57597=>"100011001",
  57598=>"010100111",
  57599=>"000000010",
  57600=>"000101111",
  57601=>"000000100",
  57602=>"010010010",
  57603=>"000001111",
  57604=>"100000000",
  57605=>"000001111",
  57606=>"111111100",
  57607=>"101101000",
  57608=>"110101101",
  57609=>"101101101",
  57610=>"100000000",
  57611=>"000101111",
  57612=>"000001101",
  57613=>"101100101",
  57614=>"000000110",
  57615=>"101111110",
  57616=>"011000101",
  57617=>"111111010",
  57618=>"111111110",
  57619=>"000100000",
  57620=>"111000000",
  57621=>"111000000",
  57622=>"100000000",
  57623=>"000010111",
  57624=>"010010000",
  57625=>"111111010",
  57626=>"011000101",
  57627=>"111000101",
  57628=>"111111111",
  57629=>"000000001",
  57630=>"000101001",
  57631=>"101000010",
  57632=>"000011111",
  57633=>"011000010",
  57634=>"111010010",
  57635=>"111000000",
  57636=>"011000001",
  57637=>"000011011",
  57638=>"010010011",
  57639=>"001000101",
  57640=>"111010000",
  57641=>"110111101",
  57642=>"001001111",
  57643=>"001000000",
  57644=>"010100111",
  57645=>"110010000",
  57646=>"000101101",
  57647=>"001000011",
  57648=>"011111110",
  57649=>"101110110",
  57650=>"111111110",
  57651=>"110000111",
  57652=>"000010000",
  57653=>"000001010",
  57654=>"111001000",
  57655=>"111111111",
  57656=>"000101000",
  57657=>"101000100",
  57658=>"110000010",
  57659=>"111111101",
  57660=>"001001011",
  57661=>"111111011",
  57662=>"000000000",
  57663=>"000001001",
  57664=>"101001000",
  57665=>"000101110",
  57666=>"100001111",
  57667=>"000100100",
  57668=>"110000010",
  57669=>"101100000",
  57670=>"111111111",
  57671=>"101011000",
  57672=>"000000010",
  57673=>"000001101",
  57674=>"000010000",
  57675=>"101101100",
  57676=>"111111111",
  57677=>"111011000",
  57678=>"110000001",
  57679=>"010111001",
  57680=>"000000010",
  57681=>"111000000",
  57682=>"000101111",
  57683=>"111110110",
  57684=>"010000100",
  57685=>"001000000",
  57686=>"000101110",
  57687=>"111001101",
  57688=>"111000010",
  57689=>"000000100",
  57690=>"001101101",
  57691=>"111000101",
  57692=>"000001000",
  57693=>"000000100",
  57694=>"111111011",
  57695=>"000001000",
  57696=>"111111111",
  57697=>"000000010",
  57698=>"000000010",
  57699=>"000111101",
  57700=>"001000111",
  57701=>"000101000",
  57702=>"000101111",
  57703=>"100100111",
  57704=>"111000110",
  57705=>"000000000",
  57706=>"111000011",
  57707=>"000111111",
  57708=>"001011111",
  57709=>"111000110",
  57710=>"000000100",
  57711=>"101111111",
  57712=>"000011011",
  57713=>"001000000",
  57714=>"111001000",
  57715=>"101111111",
  57716=>"100001000",
  57717=>"000000001",
  57718=>"000000101",
  57719=>"110111111",
  57720=>"011110100",
  57721=>"111101010",
  57722=>"011000110",
  57723=>"000000010",
  57724=>"011001001",
  57725=>"001011011",
  57726=>"111001111",
  57727=>"100000111",
  57728=>"111101101",
  57729=>"111011111",
  57730=>"101111101",
  57731=>"000010000",
  57732=>"111000000",
  57733=>"001111111",
  57734=>"100100111",
  57735=>"110110110",
  57736=>"010110000",
  57737=>"101000010",
  57738=>"100010011",
  57739=>"111111110",
  57740=>"000001000",
  57741=>"000000110",
  57742=>"001001101",
  57743=>"000000000",
  57744=>"110101100",
  57745=>"000111111",
  57746=>"111000101",
  57747=>"000000001",
  57748=>"101010011",
  57749=>"000000101",
  57750=>"000000111",
  57751=>"111101111",
  57752=>"011111111",
  57753=>"001000101",
  57754=>"010000110",
  57755=>"001000001",
  57756=>"110001011",
  57757=>"111001000",
  57758=>"111001000",
  57759=>"111001110",
  57760=>"100100100",
  57761=>"010110100",
  57762=>"001100111",
  57763=>"110010000",
  57764=>"001001101",
  57765=>"011011111",
  57766=>"111110101",
  57767=>"000101101",
  57768=>"111111000",
  57769=>"000000000",
  57770=>"000111100",
  57771=>"110111111",
  57772=>"111110111",
  57773=>"100000000",
  57774=>"000001011",
  57775=>"111111110",
  57776=>"011111101",
  57777=>"011001011",
  57778=>"101011111",
  57779=>"000000000",
  57780=>"001111100",
  57781=>"001010111",
  57782=>"111111011",
  57783=>"111001111",
  57784=>"100100100",
  57785=>"011000000",
  57786=>"000111111",
  57787=>"100101000",
  57788=>"100100010",
  57789=>"000000010",
  57790=>"000100100",
  57791=>"000100101",
  57792=>"111010110",
  57793=>"111110111",
  57794=>"011111111",
  57795=>"100100100",
  57796=>"000001111",
  57797=>"001000100",
  57798=>"000100100",
  57799=>"101000010",
  57800=>"111101001",
  57801=>"111110110",
  57802=>"111011001",
  57803=>"111010111",
  57804=>"000000100",
  57805=>"110100000",
  57806=>"000000000",
  57807=>"110001111",
  57808=>"110110110",
  57809=>"001011011",
  57810=>"111101000",
  57811=>"001110110",
  57812=>"001111101",
  57813=>"111100000",
  57814=>"000100110",
  57815=>"000001000",
  57816=>"001001000",
  57817=>"000000010",
  57818=>"110010011",
  57819=>"111110000",
  57820=>"000000001",
  57821=>"000111111",
  57822=>"111001110",
  57823=>"110000101",
  57824=>"010010010",
  57825=>"010000011",
  57826=>"111000101",
  57827=>"001010011",
  57828=>"111110101",
  57829=>"100101000",
  57830=>"101001101",
  57831=>"000000101",
  57832=>"000100100",
  57833=>"000000000",
  57834=>"001001000",
  57835=>"000100000",
  57836=>"010110111",
  57837=>"111000100",
  57838=>"101100100",
  57839=>"111000000",
  57840=>"111101111",
  57841=>"110110001",
  57842=>"000101111",
  57843=>"000011011",
  57844=>"011011101",
  57845=>"111111001",
  57846=>"101111111",
  57847=>"111111100",
  57848=>"111010000",
  57849=>"000000000",
  57850=>"111110110",
  57851=>"011010000",
  57852=>"001001000",
  57853=>"000111111",
  57854=>"111100111",
  57855=>"010011011",
  57856=>"000010000",
  57857=>"000000000",
  57858=>"100000101",
  57859=>"000000111",
  57860=>"111101101",
  57861=>"000000100",
  57862=>"001000000",
  57863=>"000101011",
  57864=>"111011011",
  57865=>"000000011",
  57866=>"011001111",
  57867=>"101000111",
  57868=>"000101111",
  57869=>"000000000",
  57870=>"010111000",
  57871=>"111111011",
  57872=>"010000001",
  57873=>"111111110",
  57874=>"110000000",
  57875=>"000111111",
  57876=>"010111111",
  57877=>"000001000",
  57878=>"001111000",
  57879=>"111111000",
  57880=>"000000010",
  57881=>"000000111",
  57882=>"001000000",
  57883=>"110110100",
  57884=>"010101011",
  57885=>"111001101",
  57886=>"111100000",
  57887=>"011000110",
  57888=>"111111000",
  57889=>"011001010",
  57890=>"001111111",
  57891=>"000000000",
  57892=>"000111110",
  57893=>"111001000",
  57894=>"101000100",
  57895=>"011001001",
  57896=>"001001111",
  57897=>"111101000",
  57898=>"010000000",
  57899=>"010110110",
  57900=>"000100110",
  57901=>"000000010",
  57902=>"111000111",
  57903=>"100111110",
  57904=>"110001000",
  57905=>"110110100",
  57906=>"111111000",
  57907=>"011111111",
  57908=>"110110111",
  57909=>"111111111",
  57910=>"011111111",
  57911=>"011110000",
  57912=>"000011111",
  57913=>"110000100",
  57914=>"000000100",
  57915=>"000111110",
  57916=>"001001111",
  57917=>"000111111",
  57918=>"010000000",
  57919=>"001000000",
  57920=>"000111111",
  57921=>"110110000",
  57922=>"011111010",
  57923=>"010100000",
  57924=>"111111111",
  57925=>"000010010",
  57926=>"011001010",
  57927=>"111000100",
  57928=>"000000001",
  57929=>"000000001",
  57930=>"100111000",
  57931=>"010001000",
  57932=>"001000111",
  57933=>"011011011",
  57934=>"011011001",
  57935=>"101000001",
  57936=>"001010111",
  57937=>"110111111",
  57938=>"111100000",
  57939=>"001110100",
  57940=>"000101111",
  57941=>"001111101",
  57942=>"000110100",
  57943=>"000001000",
  57944=>"000000111",
  57945=>"110110000",
  57946=>"000000011",
  57947=>"011110111",
  57948=>"001001000",
  57949=>"000101111",
  57950=>"011000100",
  57951=>"110000101",
  57952=>"111001001",
  57953=>"000000110",
  57954=>"111111111",
  57955=>"000000110",
  57956=>"000011010",
  57957=>"000011000",
  57958=>"011001000",
  57959=>"001101111",
  57960=>"000000100",
  57961=>"111111000",
  57962=>"000000101",
  57963=>"111100111",
  57964=>"111001001",
  57965=>"110000000",
  57966=>"000010000",
  57967=>"111111111",
  57968=>"001001000",
  57969=>"110111000",
  57970=>"110111111",
  57971=>"111110011",
  57972=>"111001111",
  57973=>"000110110",
  57974=>"000001000",
  57975=>"000100100",
  57976=>"010000000",
  57977=>"000000000",
  57978=>"000010011",
  57979=>"001111111",
  57980=>"110011001",
  57981=>"000001001",
  57982=>"010011000",
  57983=>"000000000",
  57984=>"000111000",
  57985=>"000010110",
  57986=>"000111111",
  57987=>"001011101",
  57988=>"111000000",
  57989=>"000001111",
  57990=>"110010000",
  57991=>"100100100",
  57992=>"100100110",
  57993=>"011000100",
  57994=>"001000000",
  57995=>"111111111",
  57996=>"000000000",
  57997=>"000000000",
  57998=>"111000000",
  57999=>"000001000",
  58000=>"100100110",
  58001=>"000001101",
  58002=>"000001000",
  58003=>"000000001",
  58004=>"001010000",
  58005=>"000101001",
  58006=>"111111000",
  58007=>"010110110",
  58008=>"000001010",
  58009=>"000000101",
  58010=>"101000101",
  58011=>"111111111",
  58012=>"011011000",
  58013=>"111111111",
  58014=>"111000000",
  58015=>"010000010",
  58016=>"000001001",
  58017=>"110111100",
  58018=>"000000000",
  58019=>"001001111",
  58020=>"000011111",
  58021=>"001011110",
  58022=>"000000000",
  58023=>"100000011",
  58024=>"000010000",
  58025=>"000001000",
  58026=>"111000001",
  58027=>"100010000",
  58028=>"111000010",
  58029=>"101101111",
  58030=>"011101101",
  58031=>"111000000",
  58032=>"001000111",
  58033=>"000000110",
  58034=>"000000000",
  58035=>"011011011",
  58036=>"110111111",
  58037=>"111111101",
  58038=>"000101111",
  58039=>"001000111",
  58040=>"100100110",
  58041=>"001001001",
  58042=>"000000110",
  58043=>"111101000",
  58044=>"100111110",
  58045=>"001001111",
  58046=>"110110000",
  58047=>"111111000",
  58048=>"000000111",
  58049=>"010111010",
  58050=>"110001111",
  58051=>"011011001",
  58052=>"011000000",
  58053=>"111100100",
  58054=>"111010111",
  58055=>"111010000",
  58056=>"001000111",
  58057=>"110110010",
  58058=>"100101110",
  58059=>"000001111",
  58060=>"000100100",
  58061=>"000100100",
  58062=>"111111001",
  58063=>"000011100",
  58064=>"111111111",
  58065=>"110011011",
  58066=>"001000100",
  58067=>"000001001",
  58068=>"000000001",
  58069=>"011000001",
  58070=>"000000010",
  58071=>"111110000",
  58072=>"000000000",
  58073=>"101110000",
  58074=>"000100111",
  58075=>"111111000",
  58076=>"010111010",
  58077=>"111101000",
  58078=>"010111011",
  58079=>"000001111",
  58080=>"010000000",
  58081=>"011000001",
  58082=>"111000100",
  58083=>"011011000",
  58084=>"111001000",
  58085=>"110001111",
  58086=>"111000100",
  58087=>"110111011",
  58088=>"111101001",
  58089=>"100000000",
  58090=>"110100100",
  58091=>"000100000",
  58092=>"100101100",
  58093=>"111000001",
  58094=>"010111010",
  58095=>"111000101",
  58096=>"101001001",
  58097=>"111010000",
  58098=>"001100000",
  58099=>"000011010",
  58100=>"000000000",
  58101=>"100000010",
  58102=>"000000000",
  58103=>"010111000",
  58104=>"111111000",
  58105=>"100000111",
  58106=>"000111010",
  58107=>"111110000",
  58108=>"111100000",
  58109=>"001000000",
  58110=>"100110010",
  58111=>"000110000",
  58112=>"110011001",
  58113=>"001000000",
  58114=>"111000000",
  58115=>"100000000",
  58116=>"010000000",
  58117=>"111101101",
  58118=>"111101010",
  58119=>"000000111",
  58120=>"001111111",
  58121=>"000000001",
  58122=>"110100001",
  58123=>"010100000",
  58124=>"100000000",
  58125=>"100101010",
  58126=>"111100000",
  58127=>"101001000",
  58128=>"000000011",
  58129=>"011000111",
  58130=>"011000000",
  58131=>"000001000",
  58132=>"111111001",
  58133=>"111110000",
  58134=>"110111000",
  58135=>"111001111",
  58136=>"111000000",
  58137=>"001001010",
  58138=>"010110101",
  58139=>"110000000",
  58140=>"000000000",
  58141=>"111000100",
  58142=>"111110100",
  58143=>"000100110",
  58144=>"001001000",
  58145=>"011111111",
  58146=>"110001000",
  58147=>"000111010",
  58148=>"001001100",
  58149=>"110100000",
  58150=>"010111111",
  58151=>"111001101",
  58152=>"101000110",
  58153=>"010110000",
  58154=>"001011011",
  58155=>"010000000",
  58156=>"001110101",
  58157=>"100100010",
  58158=>"111101101",
  58159=>"110001000",
  58160=>"000001111",
  58161=>"010101110",
  58162=>"000001111",
  58163=>"110111111",
  58164=>"001000000",
  58165=>"001011000",
  58166=>"011110010",
  58167=>"000011000",
  58168=>"110011111",
  58169=>"001000000",
  58170=>"111000100",
  58171=>"000000010",
  58172=>"001000111",
  58173=>"011111111",
  58174=>"000000100",
  58175=>"000100011",
  58176=>"000000000",
  58177=>"110101111",
  58178=>"101110110",
  58179=>"001011001",
  58180=>"000111110",
  58181=>"000000000",
  58182=>"110000000",
  58183=>"101001010",
  58184=>"100100110",
  58185=>"000001000",
  58186=>"000000000",
  58187=>"000000011",
  58188=>"111111000",
  58189=>"100101001",
  58190=>"000101011",
  58191=>"001000101",
  58192=>"001110111",
  58193=>"111011111",
  58194=>"101000010",
  58195=>"111001000",
  58196=>"111110000",
  58197=>"001000110",
  58198=>"100000000",
  58199=>"110000000",
  58200=>"111100100",
  58201=>"110100100",
  58202=>"000000001",
  58203=>"100110011",
  58204=>"000111111",
  58205=>"000001001",
  58206=>"111111011",
  58207=>"110100000",
  58208=>"000111111",
  58209=>"010000101",
  58210=>"001011010",
  58211=>"011011001",
  58212=>"000101000",
  58213=>"100100100",
  58214=>"011011101",
  58215=>"101000000",
  58216=>"100110000",
  58217=>"111101000",
  58218=>"100000110",
  58219=>"101010111",
  58220=>"010111111",
  58221=>"111000111",
  58222=>"111111101",
  58223=>"111101111",
  58224=>"011001000",
  58225=>"111110111",
  58226=>"010010000",
  58227=>"000000011",
  58228=>"111001000",
  58229=>"000000101",
  58230=>"100000000",
  58231=>"000110011",
  58232=>"000010110",
  58233=>"111111101",
  58234=>"111111010",
  58235=>"000000010",
  58236=>"110000011",
  58237=>"110100000",
  58238=>"000111011",
  58239=>"001001000",
  58240=>"000010000",
  58241=>"010001100",
  58242=>"100110111",
  58243=>"011000111",
  58244=>"111001000",
  58245=>"000001011",
  58246=>"011001000",
  58247=>"000000100",
  58248=>"110101001",
  58249=>"110000000",
  58250=>"000000101",
  58251=>"000000010",
  58252=>"101000010",
  58253=>"111111100",
  58254=>"110000111",
  58255=>"000000000",
  58256=>"010011100",
  58257=>"011000100",
  58258=>"001001000",
  58259=>"111001111",
  58260=>"011010000",
  58261=>"111000000",
  58262=>"100111111",
  58263=>"000011101",
  58264=>"111111111",
  58265=>"100010101",
  58266=>"101101111",
  58267=>"000101101",
  58268=>"000111111",
  58269=>"000110110",
  58270=>"010100010",
  58271=>"010011000",
  58272=>"100000011",
  58273=>"110110111",
  58274=>"111000111",
  58275=>"111001001",
  58276=>"010010000",
  58277=>"000001001",
  58278=>"111110000",
  58279=>"001011111",
  58280=>"111111111",
  58281=>"000110110",
  58282=>"001000000",
  58283=>"010001000",
  58284=>"001000000",
  58285=>"000000000",
  58286=>"110100110",
  58287=>"000111100",
  58288=>"001000000",
  58289=>"000011111",
  58290=>"000000000",
  58291=>"001001111",
  58292=>"011000001",
  58293=>"000111000",
  58294=>"000111111",
  58295=>"000000000",
  58296=>"000000111",
  58297=>"100110101",
  58298=>"000001000",
  58299=>"111111001",
  58300=>"001101111",
  58301=>"111110111",
  58302=>"000111001",
  58303=>"000011111",
  58304=>"100000000",
  58305=>"000000010",
  58306=>"111111111",
  58307=>"011111101",
  58308=>"111111100",
  58309=>"111110111",
  58310=>"111111000",
  58311=>"000001111",
  58312=>"000111111",
  58313=>"000110111",
  58314=>"011111111",
  58315=>"001000001",
  58316=>"111000111",
  58317=>"011100100",
  58318=>"001011011",
  58319=>"000000111",
  58320=>"001111101",
  58321=>"000100110",
  58322=>"110000000",
  58323=>"001000000",
  58324=>"000101110",
  58325=>"010100010",
  58326=>"010111111",
  58327=>"001001001",
  58328=>"101101111",
  58329=>"000100000",
  58330=>"011110111",
  58331=>"111000000",
  58332=>"110110100",
  58333=>"100010000",
  58334=>"000111011",
  58335=>"101000000",
  58336=>"101000011",
  58337=>"111000000",
  58338=>"111101001",
  58339=>"010110001",
  58340=>"110111111",
  58341=>"110111001",
  58342=>"000111111",
  58343=>"100011111",
  58344=>"000010111",
  58345=>"000000000",
  58346=>"000000100",
  58347=>"000000111",
  58348=>"000010111",
  58349=>"000111111",
  58350=>"000000000",
  58351=>"000110110",
  58352=>"000001000",
  58353=>"111011111",
  58354=>"111111001",
  58355=>"111001001",
  58356=>"011110101",
  58357=>"111011111",
  58358=>"000000010",
  58359=>"111111111",
  58360=>"000000111",
  58361=>"101111110",
  58362=>"000000010",
  58363=>"000111111",
  58364=>"001000000",
  58365=>"000000000",
  58366=>"000111111",
  58367=>"111000000",
  58368=>"001001000",
  58369=>"101100111",
  58370=>"110011101",
  58371=>"000110011",
  58372=>"101101011",
  58373=>"110101011",
  58374=>"011011011",
  58375=>"111100010",
  58376=>"000000101",
  58377=>"000000010",
  58378=>"100100110",
  58379=>"000101000",
  58380=>"111010001",
  58381=>"010111001",
  58382=>"011000111",
  58383=>"001101110",
  58384=>"101111011",
  58385=>"000000000",
  58386=>"000000100",
  58387=>"101010011",
  58388=>"000101111",
  58389=>"011110000",
  58390=>"001001101",
  58391=>"001101100",
  58392=>"000010000",
  58393=>"000111000",
  58394=>"011010000",
  58395=>"111100111",
  58396=>"110111111",
  58397=>"010111101",
  58398=>"001001101",
  58399=>"000000101",
  58400=>"111111111",
  58401=>"000000000",
  58402=>"100101111",
  58403=>"000100010",
  58404=>"111101101",
  58405=>"111100000",
  58406=>"010000001",
  58407=>"011001001",
  58408=>"110011101",
  58409=>"000100011",
  58410=>"101100111",
  58411=>"001111010",
  58412=>"111101110",
  58413=>"011100011",
  58414=>"111000001",
  58415=>"011100101",
  58416=>"000000111",
  58417=>"001001001",
  58418=>"011010110",
  58419=>"111110000",
  58420=>"000101101",
  58421=>"010000000",
  58422=>"001100110",
  58423=>"001001111",
  58424=>"010010010",
  58425=>"000100101",
  58426=>"100010111",
  58427=>"011000000",
  58428=>"110110110",
  58429=>"101101101",
  58430=>"000000100",
  58431=>"001001000",
  58432=>"011000000",
  58433=>"101101111",
  58434=>"010001001",
  58435=>"100001001",
  58436=>"000000010",
  58437=>"010000000",
  58438=>"000110010",
  58439=>"000000111",
  58440=>"111111011",
  58441=>"000101010",
  58442=>"101100111",
  58443=>"101000001",
  58444=>"010010010",
  58445=>"101101100",
  58446=>"100101101",
  58447=>"010111110",
  58448=>"000000111",
  58449=>"000001101",
  58450=>"101111111",
  58451=>"000000001",
  58452=>"111110111",
  58453=>"011111111",
  58454=>"011001100",
  58455=>"101011000",
  58456=>"110010000",
  58457=>"100000101",
  58458=>"110000010",
  58459=>"111100100",
  58460=>"010111011",
  58461=>"001000001",
  58462=>"111111000",
  58463=>"001100100",
  58464=>"110010011",
  58465=>"111111111",
  58466=>"011001101",
  58467=>"000000110",
  58468=>"110000100",
  58469=>"000100101",
  58470=>"011111110",
  58471=>"100001100",
  58472=>"000010000",
  58473=>"000111000",
  58474=>"000000110",
  58475=>"000111010",
  58476=>"111111111",
  58477=>"010010110",
  58478=>"100111111",
  58479=>"000101111",
  58480=>"101101100",
  58481=>"010000111",
  58482=>"100001001",
  58483=>"010000000",
  58484=>"101000111",
  58485=>"000001000",
  58486=>"110000000",
  58487=>"111111011",
  58488=>"000000001",
  58489=>"000000010",
  58490=>"000000101",
  58491=>"101001000",
  58492=>"110010011",
  58493=>"100100100",
  58494=>"000111101",
  58495=>"001000111",
  58496=>"101000000",
  58497=>"000000011",
  58498=>"111111111",
  58499=>"001111111",
  58500=>"000000111",
  58501=>"110000101",
  58502=>"001001101",
  58503=>"010000000",
  58504=>"111001001",
  58505=>"111000000",
  58506=>"111101111",
  58507=>"010000010",
  58508=>"111110000",
  58509=>"110101001",
  58510=>"111111111",
  58511=>"000000000",
  58512=>"111101001",
  58513=>"111001000",
  58514=>"100111010",
  58515=>"100000000",
  58516=>"101011111",
  58517=>"000001001",
  58518=>"111101001",
  58519=>"001000000",
  58520=>"000111000",
  58521=>"000010000",
  58522=>"110111100",
  58523=>"100111110",
  58524=>"011010110",
  58525=>"110101100",
  58526=>"000110010",
  58527=>"000000101",
  58528=>"110110100",
  58529=>"000101101",
  58530=>"111001000",
  58531=>"011100101",
  58532=>"010000110",
  58533=>"001000100",
  58534=>"110110000",
  58535=>"110111011",
  58536=>"011111101",
  58537=>"111011000",
  58538=>"101000001",
  58539=>"100000011",
  58540=>"001111000",
  58541=>"011010111",
  58542=>"001100110",
  58543=>"011000000",
  58544=>"110010000",
  58545=>"011000000",
  58546=>"101100100",
  58547=>"100000111",
  58548=>"111100000",
  58549=>"000000011",
  58550=>"000000000",
  58551=>"011100000",
  58552=>"011011111",
  58553=>"110010101",
  58554=>"100111010",
  58555=>"000000001",
  58556=>"111111000",
  58557=>"010011000",
  58558=>"000101001",
  58559=>"010010110",
  58560=>"011000000",
  58561=>"000000000",
  58562=>"001110111",
  58563=>"111101100",
  58564=>"010110110",
  58565=>"001011011",
  58566=>"000000111",
  58567=>"101100010",
  58568=>"011110000",
  58569=>"101001000",
  58570=>"010110111",
  58571=>"011011101",
  58572=>"000000001",
  58573=>"011011110",
  58574=>"000000000",
  58575=>"000000111",
  58576=>"000100000",
  58577=>"101001101",
  58578=>"000101111",
  58579=>"101001011",
  58580=>"111001001",
  58581=>"100100110",
  58582=>"000111011",
  58583=>"101010011",
  58584=>"011011000",
  58585=>"000110111",
  58586=>"011001000",
  58587=>"000000000",
  58588=>"100100101",
  58589=>"010010111",
  58590=>"001111101",
  58591=>"010010111",
  58592=>"001111000",
  58593=>"101100101",
  58594=>"011110000",
  58595=>"111110100",
  58596=>"010010100",
  58597=>"111101101",
  58598=>"011010010",
  58599=>"100000111",
  58600=>"000010011",
  58601=>"000000110",
  58602=>"001000001",
  58603=>"110101111",
  58604=>"000111011",
  58605=>"000100000",
  58606=>"000000001",
  58607=>"101100111",
  58608=>"101111011",
  58609=>"000110110",
  58610=>"010000111",
  58611=>"100100100",
  58612=>"100000101",
  58613=>"001000111",
  58614=>"000000000",
  58615=>"000111101",
  58616=>"001001011",
  58617=>"000011110",
  58618=>"101101101",
  58619=>"101111111",
  58620=>"001101111",
  58621=>"111011111",
  58622=>"111001000",
  58623=>"111000111",
  58624=>"011011000",
  58625=>"010000000",
  58626=>"001000001",
  58627=>"010000110",
  58628=>"000100001",
  58629=>"000000000",
  58630=>"011111011",
  58631=>"100100011",
  58632=>"000110010",
  58633=>"000000100",
  58634=>"000100111",
  58635=>"100000000",
  58636=>"111000000",
  58637=>"010011110",
  58638=>"000011111",
  58639=>"100000000",
  58640=>"000100100",
  58641=>"001001011",
  58642=>"100001000",
  58643=>"110100000",
  58644=>"011110010",
  58645=>"000101111",
  58646=>"110111111",
  58647=>"111101101",
  58648=>"000000000",
  58649=>"111101001",
  58650=>"110101000",
  58651=>"111001110",
  58652=>"111000110",
  58653=>"100000000",
  58654=>"100100000",
  58655=>"000110000",
  58656=>"000100011",
  58657=>"001011111",
  58658=>"000011111",
  58659=>"110110111",
  58660=>"101101001",
  58661=>"000000000",
  58662=>"000100010",
  58663=>"101000100",
  58664=>"001111011",
  58665=>"011001111",
  58666=>"001001100",
  58667=>"110000110",
  58668=>"100100111",
  58669=>"000100000",
  58670=>"111010000",
  58671=>"010000111",
  58672=>"000000001",
  58673=>"110111111",
  58674=>"001100100",
  58675=>"001001000",
  58676=>"010110000",
  58677=>"010100000",
  58678=>"000100011",
  58679=>"100110000",
  58680=>"000100110",
  58681=>"100010010",
  58682=>"000001101",
  58683=>"011111111",
  58684=>"000000000",
  58685=>"010011000",
  58686=>"100100100",
  58687=>"000110000",
  58688=>"111101111",
  58689=>"011011001",
  58690=>"111011011",
  58691=>"110110000",
  58692=>"001111011",
  58693=>"001100001",
  58694=>"111001111",
  58695=>"100110111",
  58696=>"110100000",
  58697=>"010110110",
  58698=>"001000100",
  58699=>"000111011",
  58700=>"110000000",
  58701=>"110101101",
  58702=>"011011000",
  58703=>"000000100",
  58704=>"010111001",
  58705=>"111001101",
  58706=>"100000000",
  58707=>"011101000",
  58708=>"111010010",
  58709=>"111101111",
  58710=>"111111001",
  58711=>"111100100",
  58712=>"001011101",
  58713=>"001101111",
  58714=>"001001100",
  58715=>"110111100",
  58716=>"011110011",
  58717=>"100101000",
  58718=>"111111111",
  58719=>"000000011",
  58720=>"110010010",
  58721=>"000010000",
  58722=>"111010000",
  58723=>"000010001",
  58724=>"010001000",
  58725=>"010011000",
  58726=>"010011000",
  58727=>"000111111",
  58728=>"110000010",
  58729=>"111100100",
  58730=>"010010111",
  58731=>"100100110",
  58732=>"000000110",
  58733=>"001101101",
  58734=>"100100100",
  58735=>"001000000",
  58736=>"010010001",
  58737=>"110100110",
  58738=>"011000000",
  58739=>"001011011",
  58740=>"110100111",
  58741=>"001101110",
  58742=>"110010010",
  58743=>"110010000",
  58744=>"110111110",
  58745=>"000101011",
  58746=>"001101011",
  58747=>"000100111",
  58748=>"000000000",
  58749=>"000000111",
  58750=>"000001010",
  58751=>"010011010",
  58752=>"111000100",
  58753=>"011000101",
  58754=>"110100110",
  58755=>"000000110",
  58756=>"000010110",
  58757=>"000010000",
  58758=>"010110000",
  58759=>"101111000",
  58760=>"010011001",
  58761=>"001001011",
  58762=>"001100110",
  58763=>"010100101",
  58764=>"100100101",
  58765=>"110110110",
  58766=>"111101011",
  58767=>"001000000",
  58768=>"111101111",
  58769=>"011111000",
  58770=>"011010110",
  58771=>"100100011",
  58772=>"000100110",
  58773=>"100000100",
  58774=>"110010110",
  58775=>"100010011",
  58776=>"110000010",
  58777=>"101010100",
  58778=>"110110111",
  58779=>"100100000",
  58780=>"000100001",
  58781=>"100111110",
  58782=>"011000010",
  58783=>"011100100",
  58784=>"110100110",
  58785=>"011111101",
  58786=>"000100110",
  58787=>"000000010",
  58788=>"010000010",
  58789=>"000000010",
  58790=>"001111001",
  58791=>"010110100",
  58792=>"000000011",
  58793=>"100111011",
  58794=>"100000111",
  58795=>"011101101",
  58796=>"101011011",
  58797=>"110010010",
  58798=>"000000011",
  58799=>"100110110",
  58800=>"000010110",
  58801=>"000100000",
  58802=>"100100000",
  58803=>"010100000",
  58804=>"110111110",
  58805=>"001011001",
  58806=>"101100101",
  58807=>"000000011",
  58808=>"111111101",
  58809=>"000001011",
  58810=>"111001101",
  58811=>"010100110",
  58812=>"100000001",
  58813=>"110111111",
  58814=>"111000111",
  58815=>"001101111",
  58816=>"000100100",
  58817=>"110110100",
  58818=>"111100110",
  58819=>"011111001",
  58820=>"000100111",
  58821=>"011111011",
  58822=>"000000110",
  58823=>"110111111",
  58824=>"111110011",
  58825=>"011011001",
  58826=>"000000000",
  58827=>"001000110",
  58828=>"100010010",
  58829=>"100110110",
  58830=>"101100000",
  58831=>"001100000",
  58832=>"000001011",
  58833=>"011101100",
  58834=>"001000101",
  58835=>"110100100",
  58836=>"110110110",
  58837=>"110001111",
  58838=>"000000010",
  58839=>"000000000",
  58840=>"011011010",
  58841=>"101111110",
  58842=>"001100000",
  58843=>"000100101",
  58844=>"100000000",
  58845=>"100110001",
  58846=>"011001011",
  58847=>"100100000",
  58848=>"000110010",
  58849=>"011101001",
  58850=>"000000001",
  58851=>"011001000",
  58852=>"001000010",
  58853=>"011111111",
  58854=>"101001001",
  58855=>"011111100",
  58856=>"000110111",
  58857=>"100001111",
  58858=>"011100100",
  58859=>"011100111",
  58860=>"101100000",
  58861=>"111100110",
  58862=>"111000011",
  58863=>"010000100",
  58864=>"000000101",
  58865=>"000000100",
  58866=>"010010000",
  58867=>"000000110",
  58868=>"000100011",
  58869=>"100011101",
  58870=>"000100110",
  58871=>"000100110",
  58872=>"111100110",
  58873=>"100110111",
  58874=>"000100110",
  58875=>"100111011",
  58876=>"111110110",
  58877=>"001000101",
  58878=>"100100111",
  58879=>"110010000",
  58880=>"011011000",
  58881=>"011100001",
  58882=>"101000000",
  58883=>"111100111",
  58884=>"110111111",
  58885=>"111101000",
  58886=>"010010000",
  58887=>"111111110",
  58888=>"011010000",
  58889=>"110010011",
  58890=>"100111111",
  58891=>"111000100",
  58892=>"100000011",
  58893=>"110110100",
  58894=>"000001111",
  58895=>"011101001",
  58896=>"111111000",
  58897=>"101111111",
  58898=>"010110011",
  58899=>"110010101",
  58900=>"011111111",
  58901=>"111010111",
  58902=>"100101000",
  58903=>"111100111",
  58904=>"101000010",
  58905=>"001110000",
  58906=>"111000000",
  58907=>"000010111",
  58908=>"010000101",
  58909=>"101001101",
  58910=>"010011111",
  58911=>"000101100",
  58912=>"111001001",
  58913=>"000000010",
  58914=>"000000000",
  58915=>"110111011",
  58916=>"000011000",
  58917=>"110110000",
  58918=>"101000000",
  58919=>"000000111",
  58920=>"011011000",
  58921=>"011000000",
  58922=>"001100110",
  58923=>"010000000",
  58924=>"100001011",
  58925=>"101000100",
  58926=>"000001011",
  58927=>"000000000",
  58928=>"011000111",
  58929=>"010110110",
  58930=>"000000001",
  58931=>"010010111",
  58932=>"010111000",
  58933=>"000000010",
  58934=>"110111110",
  58935=>"010000101",
  58936=>"111111000",
  58937=>"101000101",
  58938=>"000110000",
  58939=>"111101101",
  58940=>"100110100",
  58941=>"111101110",
  58942=>"000000100",
  58943=>"100111111",
  58944=>"111111011",
  58945=>"111111000",
  58946=>"000000111",
  58947=>"111011111",
  58948=>"001001111",
  58949=>"100000101",
  58950=>"000000000",
  58951=>"111111000",
  58952=>"100000000",
  58953=>"101000000",
  58954=>"101100101",
  58955=>"000111111",
  58956=>"111010111",
  58957=>"100100110",
  58958=>"011011011",
  58959=>"000000011",
  58960=>"010111111",
  58961=>"111010011",
  58962=>"110111111",
  58963=>"011100100",
  58964=>"010010000",
  58965=>"001111110",
  58966=>"011011001",
  58967=>"101000000",
  58968=>"100100110",
  58969=>"100100100",
  58970=>"011111110",
  58971=>"000100111",
  58972=>"010111010",
  58973=>"000001000",
  58974=>"000000100",
  58975=>"001001111",
  58976=>"001000100",
  58977=>"000100011",
  58978=>"000000000",
  58979=>"100111001",
  58980=>"000110000",
  58981=>"001100100",
  58982=>"010010000",
  58983=>"010100000",
  58984=>"000110111",
  58985=>"000010001",
  58986=>"010000010",
  58987=>"111000000",
  58988=>"100100000",
  58989=>"000101000",
  58990=>"000000101",
  58991=>"000000110",
  58992=>"000100100",
  58993=>"001010101",
  58994=>"011111011",
  58995=>"000000000",
  58996=>"000100111",
  58997=>"101100101",
  58998=>"100100101",
  58999=>"111000101",
  59000=>"000111010",
  59001=>"010000111",
  59002=>"000111111",
  59003=>"111100011",
  59004=>"100110010",
  59005=>"110001001",
  59006=>"111110110",
  59007=>"000100000",
  59008=>"000000001",
  59009=>"111000000",
  59010=>"010011010",
  59011=>"111000111",
  59012=>"000011111",
  59013=>"111100101",
  59014=>"011011000",
  59015=>"000000100",
  59016=>"000011011",
  59017=>"000000000",
  59018=>"010111110",
  59019=>"100111110",
  59020=>"001000000",
  59021=>"101000111",
  59022=>"101001010",
  59023=>"101000000",
  59024=>"001011001",
  59025=>"111111000",
  59026=>"011100000",
  59027=>"000010011",
  59028=>"000010010",
  59029=>"111000001",
  59030=>"000010111",
  59031=>"110100100",
  59032=>"000000000",
  59033=>"100111111",
  59034=>"010011011",
  59035=>"111110010",
  59036=>"010000000",
  59037=>"001000010",
  59038=>"010110001",
  59039=>"000000000",
  59040=>"000100100",
  59041=>"111010000",
  59042=>"101000100",
  59043=>"000000111",
  59044=>"000100111",
  59045=>"001001011",
  59046=>"111001001",
  59047=>"010111011",
  59048=>"000000111",
  59049=>"011000000",
  59050=>"000000011",
  59051=>"011011011",
  59052=>"111111000",
  59053=>"111100000",
  59054=>"110100011",
  59055=>"100100010",
  59056=>"111101100",
  59057=>"000101000",
  59058=>"000111000",
  59059=>"000000011",
  59060=>"111111111",
  59061=>"111111100",
  59062=>"111011011",
  59063=>"001011000",
  59064=>"001011001",
  59065=>"000100011",
  59066=>"110000000",
  59067=>"001111110",
  59068=>"010001101",
  59069=>"111111111",
  59070=>"000111111",
  59071=>"011000000",
  59072=>"110010000",
  59073=>"000000000",
  59074=>"011111101",
  59075=>"001111110",
  59076=>"000001101",
  59077=>"101100010",
  59078=>"101110111",
  59079=>"111110000",
  59080=>"000011000",
  59081=>"101111000",
  59082=>"111010000",
  59083=>"001001001",
  59084=>"000000010",
  59085=>"001011010",
  59086=>"111111000",
  59087=>"111010000",
  59088=>"010000110",
  59089=>"101111000",
  59090=>"000000010",
  59091=>"010111100",
  59092=>"101101111",
  59093=>"000100000",
  59094=>"101101101",
  59095=>"010101011",
  59096=>"101100100",
  59097=>"000000010",
  59098=>"000000001",
  59099=>"000100100",
  59100=>"111101110",
  59101=>"001111000",
  59102=>"101101000",
  59103=>"010011101",
  59104=>"000111010",
  59105=>"000001000",
  59106=>"000000000",
  59107=>"001001111",
  59108=>"000100011",
  59109=>"111101111",
  59110=>"111101110",
  59111=>"000101101",
  59112=>"111000000",
  59113=>"000000111",
  59114=>"011111000",
  59115=>"111111111",
  59116=>"000000000",
  59117=>"000000000",
  59118=>"000000000",
  59119=>"111000001",
  59120=>"010000101",
  59121=>"001111111",
  59122=>"000000010",
  59123=>"111111011",
  59124=>"110111111",
  59125=>"000101101",
  59126=>"100000000",
  59127=>"010000100",
  59128=>"000000010",
  59129=>"100000010",
  59130=>"111000101",
  59131=>"000111110",
  59132=>"011011000",
  59133=>"111000000",
  59134=>"010101101",
  59135=>"101000101",
  59136=>"101011001",
  59137=>"101111101",
  59138=>"000000101",
  59139=>"111101111",
  59140=>"000101000",
  59141=>"110000000",
  59142=>"000000010",
  59143=>"111101101",
  59144=>"100000011",
  59145=>"111000000",
  59146=>"100110111",
  59147=>"111100111",
  59148=>"000011001",
  59149=>"000000000",
  59150=>"000101001",
  59151=>"000101111",
  59152=>"010000111",
  59153=>"110110111",
  59154=>"000001000",
  59155=>"111000000",
  59156=>"010011101",
  59157=>"000000000",
  59158=>"111110011",
  59159=>"000000111",
  59160=>"111111000",
  59161=>"011111111",
  59162=>"011010101",
  59163=>"000000111",
  59164=>"101001100",
  59165=>"110000100",
  59166=>"010010001",
  59167=>"111100000",
  59168=>"111101000",
  59169=>"100000000",
  59170=>"000001000",
  59171=>"110001101",
  59172=>"111000100",
  59173=>"100110111",
  59174=>"111111010",
  59175=>"000101111",
  59176=>"111111010",
  59177=>"000110010",
  59178=>"000000000",
  59179=>"110000000",
  59180=>"101000000",
  59181=>"111100110",
  59182=>"100000001",
  59183=>"010001111",
  59184=>"000110111",
  59185=>"000000000",
  59186=>"000011111",
  59187=>"000111101",
  59188=>"100000111",
  59189=>"111110000",
  59190=>"110010000",
  59191=>"101000000",
  59192=>"011001111",
  59193=>"111100101",
  59194=>"000000111",
  59195=>"100101101",
  59196=>"100100100",
  59197=>"000101101",
  59198=>"000000000",
  59199=>"111111010",
  59200=>"100011111",
  59201=>"101100001",
  59202=>"111111111",
  59203=>"011111010",
  59204=>"000010010",
  59205=>"000000000",
  59206=>"010000000",
  59207=>"011111011",
  59208=>"000000101",
  59209=>"000100011",
  59210=>"101101111",
  59211=>"000010111",
  59212=>"101001011",
  59213=>"010011000",
  59214=>"000111101",
  59215=>"000001111",
  59216=>"101111000",
  59217=>"010010000",
  59218=>"000000100",
  59219=>"011101000",
  59220=>"101101111",
  59221=>"001110000",
  59222=>"001011010",
  59223=>"001001101",
  59224=>"000100011",
  59225=>"111101000",
  59226=>"111100100",
  59227=>"000100111",
  59228=>"000000111",
  59229=>"100001010",
  59230=>"010010011",
  59231=>"100011010",
  59232=>"111111111",
  59233=>"000111111",
  59234=>"101000111",
  59235=>"001001001",
  59236=>"000100001",
  59237=>"100111011",
  59238=>"000110000",
  59239=>"111000000",
  59240=>"010110000",
  59241=>"010111111",
  59242=>"111010010",
  59243=>"111000101",
  59244=>"000000100",
  59245=>"010111110",
  59246=>"111111111",
  59247=>"100010111",
  59248=>"100000111",
  59249=>"100000111",
  59250=>"010000000",
  59251=>"000000011",
  59252=>"000100111",
  59253=>"101000000",
  59254=>"000010111",
  59255=>"001111010",
  59256=>"001000101",
  59257=>"000101101",
  59258=>"000000110",
  59259=>"101000000",
  59260=>"101110000",
  59261=>"110110000",
  59262=>"111100101",
  59263=>"101000111",
  59264=>"010010000",
  59265=>"101000101",
  59266=>"000011111",
  59267=>"000010111",
  59268=>"000101111",
  59269=>"111111101",
  59270=>"011001001",
  59271=>"000000011",
  59272=>"111110000",
  59273=>"101100100",
  59274=>"010111111",
  59275=>"101000000",
  59276=>"010111000",
  59277=>"101101111",
  59278=>"000101101",
  59279=>"000000100",
  59280=>"011100000",
  59281=>"100100000",
  59282=>"010000101",
  59283=>"000000011",
  59284=>"001001100",
  59285=>"000000000",
  59286=>"010011000",
  59287=>"100011011",
  59288=>"011111111",
  59289=>"111000000",
  59290=>"001010011",
  59291=>"000000000",
  59292=>"100100101",
  59293=>"111111000",
  59294=>"101101000",
  59295=>"000100000",
  59296=>"100101011",
  59297=>"010111010",
  59298=>"001101111",
  59299=>"101111110",
  59300=>"110010100",
  59301=>"010110110",
  59302=>"100110011",
  59303=>"000000110",
  59304=>"111111000",
  59305=>"000010101",
  59306=>"001111111",
  59307=>"000000000",
  59308=>"000111101",
  59309=>"001101111",
  59310=>"100100100",
  59311=>"111110000",
  59312=>"010111111",
  59313=>"000101100",
  59314=>"000000010",
  59315=>"000000100",
  59316=>"101011011",
  59317=>"111010000",
  59318=>"000011011",
  59319=>"001101111",
  59320=>"000000001",
  59321=>"100110100",
  59322=>"111000001",
  59323=>"010111111",
  59324=>"000000100",
  59325=>"001011111",
  59326=>"001011011",
  59327=>"111000001",
  59328=>"001000101",
  59329=>"010110111",
  59330=>"010111011",
  59331=>"000100011",
  59332=>"000000111",
  59333=>"100000001",
  59334=>"110001000",
  59335=>"000010000",
  59336=>"000010101",
  59337=>"010010000",
  59338=>"111111000",
  59339=>"101000101",
  59340=>"010000000",
  59341=>"111000001",
  59342=>"101111100",
  59343=>"000000000",
  59344=>"111100111",
  59345=>"100110110",
  59346=>"000000110",
  59347=>"000111111",
  59348=>"100000001",
  59349=>"010100001",
  59350=>"101101101",
  59351=>"010110101",
  59352=>"100000101",
  59353=>"100000000",
  59354=>"000011000",
  59355=>"000110010",
  59356=>"001011110",
  59357=>"101011111",
  59358=>"010111000",
  59359=>"010100000",
  59360=>"010000001",
  59361=>"001100101",
  59362=>"111000111",
  59363=>"110001001",
  59364=>"000111101",
  59365=>"110010010",
  59366=>"111000010",
  59367=>"101011001",
  59368=>"010000011",
  59369=>"101000101",
  59370=>"000001011",
  59371=>"000011000",
  59372=>"010010111",
  59373=>"010111000",
  59374=>"000000000",
  59375=>"000000010",
  59376=>"101000000",
  59377=>"001000100",
  59378=>"110110001",
  59379=>"101000001",
  59380=>"111110100",
  59381=>"001000101",
  59382=>"000000000",
  59383=>"001000011",
  59384=>"101000111",
  59385=>"000000111",
  59386=>"110110000",
  59387=>"111000001",
  59388=>"101000111",
  59389=>"011000101",
  59390=>"101110001",
  59391=>"000000010",
  59392=>"010011011",
  59393=>"001000110",
  59394=>"111000000",
  59395=>"100000001",
  59396=>"010000011",
  59397=>"110110000",
  59398=>"000000000",
  59399=>"111011110",
  59400=>"010001011",
  59401=>"000000000",
  59402=>"110100000",
  59403=>"000000001",
  59404=>"111000000",
  59405=>"000111111",
  59406=>"001001011",
  59407=>"111101000",
  59408=>"010111101",
  59409=>"000001001",
  59410=>"110001000",
  59411=>"110010000",
  59412=>"111111001",
  59413=>"101100000",
  59414=>"000011111",
  59415=>"111000000",
  59416=>"010001001",
  59417=>"111111111",
  59418=>"000111010",
  59419=>"000111011",
  59420=>"010101001",
  59421=>"110000100",
  59422=>"100010000",
  59423=>"111000000",
  59424=>"000000000",
  59425=>"000010000",
  59426=>"001101111",
  59427=>"000100110",
  59428=>"000100001",
  59429=>"010010001",
  59430=>"000000110",
  59431=>"000011010",
  59432=>"000110010",
  59433=>"110111111",
  59434=>"111000100",
  59435=>"000001000",
  59436=>"010111110",
  59437=>"000011001",
  59438=>"000000000",
  59439=>"110001000",
  59440=>"000000111",
  59441=>"000111101",
  59442=>"001000100",
  59443=>"110111001",
  59444=>"001000000",
  59445=>"000000000",
  59446=>"000111101",
  59447=>"011000000",
  59448=>"110011000",
  59449=>"111000000",
  59450=>"111101000",
  59451=>"000110101",
  59452=>"000110111",
  59453=>"000001000",
  59454=>"001000001",
  59455=>"011111111",
  59456=>"101110110",
  59457=>"100110011",
  59458=>"000000000",
  59459=>"000011000",
  59460=>"111111111",
  59461=>"010000101",
  59462=>"000111000",
  59463=>"111111101",
  59464=>"110111111",
  59465=>"011001011",
  59466=>"111101111",
  59467=>"111000001",
  59468=>"000110110",
  59469=>"111011000",
  59470=>"000011011",
  59471=>"010110110",
  59472=>"000000010",
  59473=>"000111100",
  59474=>"111011111",
  59475=>"010011100",
  59476=>"110000000",
  59477=>"110111110",
  59478=>"010011001",
  59479=>"010010011",
  59480=>"000111110",
  59481=>"000101111",
  59482=>"000011111",
  59483=>"000000000",
  59484=>"001000111",
  59485=>"111000001",
  59486=>"011011010",
  59487=>"010100000",
  59488=>"000110110",
  59489=>"010110111",
  59490=>"001000111",
  59491=>"000100110",
  59492=>"011011001",
  59493=>"111000000",
  59494=>"100111111",
  59495=>"110000000",
  59496=>"010111110",
  59497=>"111000000",
  59498=>"000111010",
  59499=>"111011111",
  59500=>"111001000",
  59501=>"000000000",
  59502=>"011101111",
  59503=>"110100001",
  59504=>"000110111",
  59505=>"111001111",
  59506=>"000010111",
  59507=>"001100011",
  59508=>"000111111",
  59509=>"000000001",
  59510=>"110000000",
  59511=>"000111000",
  59512=>"111010000",
  59513=>"111011011",
  59514=>"000000010",
  59515=>"110000001",
  59516=>"111000110",
  59517=>"000100000",
  59518=>"111111000",
  59519=>"111000100",
  59520=>"111010000",
  59521=>"111000010",
  59522=>"011111110",
  59523=>"111001001",
  59524=>"000110000",
  59525=>"111001001",
  59526=>"100110111",
  59527=>"100100110",
  59528=>"011111111",
  59529=>"111100000",
  59530=>"000000101",
  59531=>"101010000",
  59532=>"111000010",
  59533=>"111100000",
  59534=>"111000000",
  59535=>"000000000",
  59536=>"000110111",
  59537=>"110110111",
  59538=>"101111111",
  59539=>"111000110",
  59540=>"110110111",
  59541=>"111000000",
  59542=>"001000011",
  59543=>"000011001",
  59544=>"000000000",
  59545=>"111011110",
  59546=>"010111111",
  59547=>"010001000",
  59548=>"101000101",
  59549=>"111000000",
  59550=>"000000000",
  59551=>"111000000",
  59552=>"011100011",
  59553=>"000111101",
  59554=>"111001001",
  59555=>"000000001",
  59556=>"111010000",
  59557=>"011111111",
  59558=>"000111100",
  59559=>"010000010",
  59560=>"000111100",
  59561=>"000111111",
  59562=>"010011111",
  59563=>"000110001",
  59564=>"101110000",
  59565=>"000000001",
  59566=>"010100001",
  59567=>"111100000",
  59568=>"000000000",
  59569=>"001001001",
  59570=>"101010000",
  59571=>"010000100",
  59572=>"010111110",
  59573=>"001000100",
  59574=>"000110111",
  59575=>"000111111",
  59576=>"000110111",
  59577=>"101011101",
  59578=>"011111011",
  59579=>"111110010",
  59580=>"100000000",
  59581=>"111111111",
  59582=>"000110111",
  59583=>"000000001",
  59584=>"111101001",
  59585=>"000000000",
  59586=>"000000111",
  59587=>"010110000",
  59588=>"101000000",
  59589=>"101101100",
  59590=>"110100100",
  59591=>"000110000",
  59592=>"010001101",
  59593=>"101110110",
  59594=>"101101111",
  59595=>"101000000",
  59596=>"111000000",
  59597=>"110001000",
  59598=>"101010010",
  59599=>"000010111",
  59600=>"010000000",
  59601=>"000110110",
  59602=>"110110110",
  59603=>"111110001",
  59604=>"111000000",
  59605=>"111000110",
  59606=>"111000011",
  59607=>"010011000",
  59608=>"111001000",
  59609=>"000000101",
  59610=>"001001000",
  59611=>"111000000",
  59612=>"010111101",
  59613=>"010111011",
  59614=>"001110010",
  59615=>"111111100",
  59616=>"001001110",
  59617=>"000000001",
  59618=>"111001000",
  59619=>"000001111",
  59620=>"111000000",
  59621=>"111001111",
  59622=>"100001001",
  59623=>"111111001",
  59624=>"111111111",
  59625=>"010010111",
  59626=>"011001000",
  59627=>"000000110",
  59628=>"000110111",
  59629=>"000000111",
  59630=>"000000000",
  59631=>"010001110",
  59632=>"011110100",
  59633=>"101001111",
  59634=>"111000000",
  59635=>"111001001",
  59636=>"000111111",
  59637=>"010011011",
  59638=>"101000000",
  59639=>"010000101",
  59640=>"110010000",
  59641=>"111000000",
  59642=>"111000001",
  59643=>"000110110",
  59644=>"111110100",
  59645=>"111101001",
  59646=>"000100100",
  59647=>"110000000",
  59648=>"001101111",
  59649=>"011000110",
  59650=>"000101111",
  59651=>"010011000",
  59652=>"000100111",
  59653=>"110101100",
  59654=>"111011111",
  59655=>"011010110",
  59656=>"111001111",
  59657=>"000000000",
  59658=>"000110110",
  59659=>"000000000",
  59660=>"000011000",
  59661=>"111100111",
  59662=>"101101110",
  59663=>"110000011",
  59664=>"111111001",
  59665=>"000110100",
  59666=>"110101100",
  59667=>"000010111",
  59668=>"111110111",
  59669=>"101100100",
  59670=>"001110110",
  59671=>"111111101",
  59672=>"000100110",
  59673=>"001100100",
  59674=>"111101111",
  59675=>"000000111",
  59676=>"001000101",
  59677=>"111111101",
  59678=>"111100000",
  59679=>"101001001",
  59680=>"000010010",
  59681=>"101100000",
  59682=>"000101111",
  59683=>"000101000",
  59684=>"101100000",
  59685=>"100000100",
  59686=>"000000100",
  59687=>"001111111",
  59688=>"000111000",
  59689=>"001101110",
  59690=>"011000111",
  59691=>"111010000",
  59692=>"011011000",
  59693=>"010100101",
  59694=>"011100110",
  59695=>"000111011",
  59696=>"000000000",
  59697=>"101111111",
  59698=>"100100101",
  59699=>"111100111",
  59700=>"000010000",
  59701=>"111111110",
  59702=>"110000010",
  59703=>"011001101",
  59704=>"111101101",
  59705=>"111101101",
  59706=>"100000000",
  59707=>"100011101",
  59708=>"001011000",
  59709=>"111111111",
  59710=>"011010011",
  59711=>"111001001",
  59712=>"100001000",
  59713=>"100101100",
  59714=>"111101011",
  59715=>"101100110",
  59716=>"000100111",
  59717=>"111000010",
  59718=>"010000101",
  59719=>"000010000",
  59720=>"110001000",
  59721=>"000111101",
  59722=>"010100011",
  59723=>"101000100",
  59724=>"111101111",
  59725=>"101101100",
  59726=>"000110011",
  59727=>"111001001",
  59728=>"001000100",
  59729=>"111110010",
  59730=>"111011111",
  59731=>"001001001",
  59732=>"010011111",
  59733=>"101100000",
  59734=>"100000001",
  59735=>"111100111",
  59736=>"111100101",
  59737=>"101011011",
  59738=>"101001001",
  59739=>"101100000",
  59740=>"100101111",
  59741=>"010001011",
  59742=>"101101111",
  59743=>"101001100",
  59744=>"011000000",
  59745=>"111010000",
  59746=>"001000100",
  59747=>"111100000",
  59748=>"000000111",
  59749=>"100011001",
  59750=>"111100100",
  59751=>"000010010",
  59752=>"100010111",
  59753=>"101000100",
  59754=>"100101010",
  59755=>"001100111",
  59756=>"110000100",
  59757=>"000011111",
  59758=>"100111111",
  59759=>"100100111",
  59760=>"001110000",
  59761=>"100110110",
  59762=>"011000110",
  59763=>"000000000",
  59764=>"000011111",
  59765=>"101000000",
  59766=>"100000111",
  59767=>"000011010",
  59768=>"000000000",
  59769=>"101110111",
  59770=>"100000111",
  59771=>"001000101",
  59772=>"111111111",
  59773=>"000000000",
  59774=>"001000110",
  59775=>"101000110",
  59776=>"010000000",
  59777=>"111001001",
  59778=>"000000000",
  59779=>"011111110",
  59780=>"111110111",
  59781=>"010110110",
  59782=>"011001000",
  59783=>"001001000",
  59784=>"000101100",
  59785=>"101100111",
  59786=>"010111011",
  59787=>"000000000",
  59788=>"100100100",
  59789=>"000010000",
  59790=>"000011010",
  59791=>"000000000",
  59792=>"000001000",
  59793=>"101001101",
  59794=>"101100111",
  59795=>"100000000",
  59796=>"000111001",
  59797=>"100100101",
  59798=>"101111100",
  59799=>"110100100",
  59800=>"001010000",
  59801=>"101000000",
  59802=>"000010000",
  59803=>"000010100",
  59804=>"111100100",
  59805=>"000000000",
  59806=>"111111100",
  59807=>"111101111",
  59808=>"000000000",
  59809=>"111111111",
  59810=>"000110111",
  59811=>"000100100",
  59812=>"000001111",
  59813=>"100110000",
  59814=>"001101011",
  59815=>"100111011",
  59816=>"001011111",
  59817=>"001101000",
  59818=>"100000101",
  59819=>"100100100",
  59820=>"100100100",
  59821=>"111101111",
  59822=>"110110101",
  59823=>"010010000",
  59824=>"101000000",
  59825=>"011100111",
  59826=>"101101110",
  59827=>"000001110",
  59828=>"010011101",
  59829=>"010010000",
  59830=>"000011011",
  59831=>"000011000",
  59832=>"010100000",
  59833=>"110110100",
  59834=>"011011011",
  59835=>"001000111",
  59836=>"000010110",
  59837=>"011111111",
  59838=>"011100110",
  59839=>"000111000",
  59840=>"111101101",
  59841=>"000000000",
  59842=>"110010100",
  59843=>"000011011",
  59844=>"101110010",
  59845=>"101100100",
  59846=>"011011100",
  59847=>"101100111",
  59848=>"100101111",
  59849=>"111000111",
  59850=>"010111001",
  59851=>"001101000",
  59852=>"110011010",
  59853=>"000111110",
  59854=>"000011000",
  59855=>"101000100",
  59856=>"111101110",
  59857=>"011001111",
  59858=>"000000111",
  59859=>"110111001",
  59860=>"101100000",
  59861=>"011001000",
  59862=>"111101111",
  59863=>"010010000",
  59864=>"000000001",
  59865=>"000000111",
  59866=>"000010000",
  59867=>"000011000",
  59868=>"101011101",
  59869=>"011001111",
  59870=>"010111111",
  59871=>"000000011",
  59872=>"101100101",
  59873=>"111001100",
  59874=>"010011010",
  59875=>"101001001",
  59876=>"101000001",
  59877=>"101011011",
  59878=>"111111111",
  59879=>"000010000",
  59880=>"000000010",
  59881=>"111010000",
  59882=>"110011011",
  59883=>"100111011",
  59884=>"000000011",
  59885=>"100000000",
  59886=>"110000001",
  59887=>"100000010",
  59888=>"000000001",
  59889=>"001000001",
  59890=>"000000000",
  59891=>"111110011",
  59892=>"110000001",
  59893=>"101001011",
  59894=>"000000000",
  59895=>"000011000",
  59896=>"110001000",
  59897=>"111110001",
  59898=>"101100111",
  59899=>"011111100",
  59900=>"101100001",
  59901=>"000001011",
  59902=>"001011001",
  59903=>"001000000",
  59904=>"001101100",
  59905=>"100001111",
  59906=>"101000101",
  59907=>"000101011",
  59908=>"001001011",
  59909=>"111110100",
  59910=>"100000100",
  59911=>"111111111",
  59912=>"000000000",
  59913=>"100000000",
  59914=>"101000000",
  59915=>"111101111",
  59916=>"000001111",
  59917=>"010111001",
  59918=>"001001011",
  59919=>"111111010",
  59920=>"011000010",
  59921=>"101000111",
  59922=>"111100001",
  59923=>"011011000",
  59924=>"001010000",
  59925=>"101000000",
  59926=>"111001000",
  59927=>"101101110",
  59928=>"101000110",
  59929=>"111111101",
  59930=>"000000100",
  59931=>"100000000",
  59932=>"010010010",
  59933=>"000000000",
  59934=>"110110000",
  59935=>"000010010",
  59936=>"010011100",
  59937=>"010111111",
  59938=>"100011010",
  59939=>"000000000",
  59940=>"000011011",
  59941=>"110110011",
  59942=>"000010010",
  59943=>"011010001",
  59944=>"011111001",
  59945=>"000110110",
  59946=>"101001001",
  59947=>"101111100",
  59948=>"001011011",
  59949=>"101000011",
  59950=>"111100000",
  59951=>"010111111",
  59952=>"010110110",
  59953=>"001011011",
  59954=>"111000010",
  59955=>"100101101",
  59956=>"010000000",
  59957=>"001001000",
  59958=>"100000000",
  59959=>"000100101",
  59960=>"001101101",
  59961=>"001000000",
  59962=>"111101000",
  59963=>"000100111",
  59964=>"001110000",
  59965=>"111111010",
  59966=>"100000000",
  59967=>"111010000",
  59968=>"111011011",
  59969=>"000000101",
  59970=>"100000011",
  59971=>"111000100",
  59972=>"110000011",
  59973=>"111010111",
  59974=>"101000000",
  59975=>"000001000",
  59976=>"010010011",
  59977=>"001111001",
  59978=>"111100001",
  59979=>"011111011",
  59980=>"000100000",
  59981=>"000100100",
  59982=>"000110110",
  59983=>"100110111",
  59984=>"000101111",
  59985=>"010110111",
  59986=>"011011000",
  59987=>"111101000",
  59988=>"111000110",
  59989=>"111110110",
  59990=>"011100101",
  59991=>"001000111",
  59992=>"111111100",
  59993=>"000111000",
  59994=>"110110111",
  59995=>"010100111",
  59996=>"000100000",
  59997=>"001001001",
  59998=>"100010000",
  59999=>"111000000",
  60000=>"010111110",
  60001=>"000000000",
  60002=>"110111000",
  60003=>"111101000",
  60004=>"010001101",
  60005=>"001001101",
  60006=>"010010000",
  60007=>"001001000",
  60008=>"000000101",
  60009=>"110000101",
  60010=>"111111101",
  60011=>"010011110",
  60012=>"001000110",
  60013=>"001101000",
  60014=>"111101111",
  60015=>"100000001",
  60016=>"110110001",
  60017=>"000100101",
  60018=>"011000110",
  60019=>"011111000",
  60020=>"111010010",
  60021=>"000000010",
  60022=>"100000101",
  60023=>"011010000",
  60024=>"111000001",
  60025=>"111010000",
  60026=>"111010010",
  60027=>"101111111",
  60028=>"000110110",
  60029=>"010100000",
  60030=>"011000011",
  60031=>"101100000",
  60032=>"000101110",
  60033=>"010111111",
  60034=>"111000010",
  60035=>"110001001",
  60036=>"010000000",
  60037=>"111111111",
  60038=>"111101110",
  60039=>"011000000",
  60040=>"000100000",
  60041=>"000000000",
  60042=>"100100010",
  60043=>"011001000",
  60044=>"001010000",
  60045=>"000010110",
  60046=>"101001001",
  60047=>"001001000",
  60048=>"000100100",
  60049=>"000100111",
  60050=>"000100000",
  60051=>"111001101",
  60052=>"000000000",
  60053=>"111000101",
  60054=>"111101001",
  60055=>"010011011",
  60056=>"000110111",
  60057=>"000111111",
  60058=>"111101101",
  60059=>"111101011",
  60060=>"111101101",
  60061=>"111101101",
  60062=>"101101001",
  60063=>"000000101",
  60064=>"000010000",
  60065=>"101100000",
  60066=>"011001001",
  60067=>"101001010",
  60068=>"000000010",
  60069=>"000000010",
  60070=>"010110100",
  60071=>"101000100",
  60072=>"101100000",
  60073=>"010010111",
  60074=>"111100000",
  60075=>"010101000",
  60076=>"010101001",
  60077=>"111101111",
  60078=>"001001001",
  60079=>"101000111",
  60080=>"011101000",
  60081=>"111010011",
  60082=>"000010010",
  60083=>"000001000",
  60084=>"101000001",
  60085=>"000100000",
  60086=>"111111111",
  60087=>"000111101",
  60088=>"100011011",
  60089=>"110000110",
  60090=>"011000001",
  60091=>"111111001",
  60092=>"000000000",
  60093=>"111111111",
  60094=>"000100100",
  60095=>"001101010",
  60096=>"101001001",
  60097=>"111100111",
  60098=>"111100110",
  60099=>"011101001",
  60100=>"000101010",
  60101=>"000101111",
  60102=>"000000011",
  60103=>"000010000",
  60104=>"101001101",
  60105=>"010000000",
  60106=>"101101101",
  60107=>"111001101",
  60108=>"111000100",
  60109=>"000010011",
  60110=>"010111101",
  60111=>"010111100",
  60112=>"111111000",
  60113=>"111101110",
  60114=>"010011101",
  60115=>"111101010",
  60116=>"000010110",
  60117=>"001101111",
  60118=>"000111111",
  60119=>"111100101",
  60120=>"000110000",
  60121=>"001001100",
  60122=>"000000000",
  60123=>"100000101",
  60124=>"111001000",
  60125=>"111011000",
  60126=>"010111110",
  60127=>"010111011",
  60128=>"000011010",
  60129=>"111100100",
  60130=>"011010000",
  60131=>"011101000",
  60132=>"111000101",
  60133=>"000010110",
  60134=>"011111111",
  60135=>"001111000",
  60136=>"000000011",
  60137=>"001000000",
  60138=>"100000000",
  60139=>"000000000",
  60140=>"000000011",
  60141=>"010001111",
  60142=>"000000100",
  60143=>"001011010",
  60144=>"010111000",
  60145=>"001000110",
  60146=>"111000000",
  60147=>"010000000",
  60148=>"110101110",
  60149=>"111101101",
  60150=>"000000000",
  60151=>"101101001",
  60152=>"111001001",
  60153=>"111001010",
  60154=>"110000000",
  60155=>"101101000",
  60156=>"001101101",
  60157=>"101000000",
  60158=>"110110111",
  60159=>"101000000",
  60160=>"010100100",
  60161=>"010000001",
  60162=>"111001001",
  60163=>"101001110",
  60164=>"011011010",
  60165=>"111110000",
  60166=>"000110111",
  60167=>"101000010",
  60168=>"100101100",
  60169=>"001001111",
  60170=>"010111001",
  60171=>"000001111",
  60172=>"101000001",
  60173=>"111001001",
  60174=>"100110111",
  60175=>"001000001",
  60176=>"100000100",
  60177=>"111110110",
  60178=>"111111100",
  60179=>"011000000",
  60180=>"011110000",
  60181=>"111110010",
  60182=>"010101101",
  60183=>"100000110",
  60184=>"111110000",
  60185=>"010111011",
  60186=>"010011100",
  60187=>"000000111",
  60188=>"001010111",
  60189=>"000000000",
  60190=>"111010100",
  60191=>"000011101",
  60192=>"101101111",
  60193=>"010000001",
  60194=>"000000011",
  60195=>"111111111",
  60196=>"000101100",
  60197=>"000010011",
  60198=>"111110010",
  60199=>"010001001",
  60200=>"000111111",
  60201=>"001111111",
  60202=>"110000000",
  60203=>"001101111",
  60204=>"111111100",
  60205=>"101111010",
  60206=>"010000110",
  60207=>"000010000",
  60208=>"010010000",
  60209=>"000100100",
  60210=>"110111001",
  60211=>"000111111",
  60212=>"111111111",
  60213=>"001001000",
  60214=>"110100011",
  60215=>"001101110",
  60216=>"110100010",
  60217=>"000010011",
  60218=>"000111100",
  60219=>"100111111",
  60220=>"100000011",
  60221=>"011111101",
  60222=>"000000101",
  60223=>"110010001",
  60224=>"110111111",
  60225=>"000000100",
  60226=>"000000111",
  60227=>"001100000",
  60228=>"111001011",
  60229=>"111100101",
  60230=>"000110010",
  60231=>"010111111",
  60232=>"011000111",
  60233=>"011110111",
  60234=>"100100111",
  60235=>"110000100",
  60236=>"111001000",
  60237=>"001011111",
  60238=>"100110100",
  60239=>"010111111",
  60240=>"001111000",
  60241=>"110111000",
  60242=>"011010100",
  60243=>"000000100",
  60244=>"000100000",
  60245=>"100100110",
  60246=>"000101101",
  60247=>"000110101",
  60248=>"000011010",
  60249=>"001001000",
  60250=>"001111000",
  60251=>"010011010",
  60252=>"010000100",
  60253=>"000000000",
  60254=>"111111000",
  60255=>"100000000",
  60256=>"111001101",
  60257=>"000111110",
  60258=>"101000111",
  60259=>"101100000",
  60260=>"001000000",
  60261=>"001100100",
  60262=>"111111000",
  60263=>"000000100",
  60264=>"111000110",
  60265=>"000111111",
  60266=>"111000000",
  60267=>"111010010",
  60268=>"000101111",
  60269=>"010111011",
  60270=>"010111010",
  60271=>"010010010",
  60272=>"001001111",
  60273=>"000000111",
  60274=>"011001110",
  60275=>"000111000",
  60276=>"111000011",
  60277=>"101000011",
  60278=>"000000101",
  60279=>"011000101",
  60280=>"111000101",
  60281=>"111000111",
  60282=>"101000001",
  60283=>"000000001",
  60284=>"000101001",
  60285=>"010000001",
  60286=>"000100000",
  60287=>"100111101",
  60288=>"010011010",
  60289=>"100010010",
  60290=>"111000010",
  60291=>"011000010",
  60292=>"111101101",
  60293=>"000000010",
  60294=>"011011110",
  60295=>"000001011",
  60296=>"100100100",
  60297=>"000000111",
  60298=>"000010101",
  60299=>"000000111",
  60300=>"000000000",
  60301=>"111111010",
  60302=>"001100110",
  60303=>"001000011",
  60304=>"011011001",
  60305=>"000010111",
  60306=>"010000010",
  60307=>"000010111",
  60308=>"000000001",
  60309=>"111000111",
  60310=>"000111000",
  60311=>"100110000",
  60312=>"111000101",
  60313=>"110010010",
  60314=>"110010010",
  60315=>"000000000",
  60316=>"000111010",
  60317=>"111100000",
  60318=>"010000000",
  60319=>"000101111",
  60320=>"011011011",
  60321=>"001000011",
  60322=>"000000001",
  60323=>"001110111",
  60324=>"010000011",
  60325=>"110110100",
  60326=>"101111000",
  60327=>"101000000",
  60328=>"110111110",
  60329=>"111000000",
  60330=>"111001111",
  60331=>"111111111",
  60332=>"000010111",
  60333=>"100000100",
  60334=>"001011011",
  60335=>"001101111",
  60336=>"101000000",
  60337=>"000110110",
  60338=>"000100100",
  60339=>"000010110",
  60340=>"000000000",
  60341=>"101100000",
  60342=>"111100100",
  60343=>"000000101",
  60344=>"001000111",
  60345=>"000000110",
  60346=>"110010000",
  60347=>"111011011",
  60348=>"000000011",
  60349=>"011011011",
  60350=>"001001011",
  60351=>"100100000",
  60352=>"000111110",
  60353=>"010111010",
  60354=>"111010010",
  60355=>"000001000",
  60356=>"000000001",
  60357=>"110110001",
  60358=>"000000111",
  60359=>"000111000",
  60360=>"110000000",
  60361=>"011111010",
  60362=>"111110000",
  60363=>"010110111",
  60364=>"011000001",
  60365=>"000101111",
  60366=>"001111000",
  60367=>"111011110",
  60368=>"111011000",
  60369=>"001100010",
  60370=>"010010011",
  60371=>"111101011",
  60372=>"111000000",
  60373=>"001011000",
  60374=>"111111111",
  60375=>"110001001",
  60376=>"000010010",
  60377=>"101000001",
  60378=>"100110110",
  60379=>"000101001",
  60380=>"000001001",
  60381=>"111101001",
  60382=>"111101101",
  60383=>"010000010",
  60384=>"010111111",
  60385=>"110111111",
  60386=>"101001101",
  60387=>"001011001",
  60388=>"000010000",
  60389=>"000000000",
  60390=>"111101111",
  60391=>"001101100",
  60392=>"110000100",
  60393=>"000000111",
  60394=>"111111110",
  60395=>"001101111",
  60396=>"000110111",
  60397=>"101000001",
  60398=>"000000000",
  60399=>"000000010",
  60400=>"111101001",
  60401=>"011011100",
  60402=>"000000010",
  60403=>"000000001",
  60404=>"000001001",
  60405=>"010111000",
  60406=>"000100000",
  60407=>"111100111",
  60408=>"111000001",
  60409=>"000000111",
  60410=>"111010111",
  60411=>"111010010",
  60412=>"010010000",
  60413=>"111111111",
  60414=>"000100000",
  60415=>"111001000",
  60416=>"111110110",
  60417=>"000000000",
  60418=>"000000100",
  60419=>"111111111",
  60420=>"110111101",
  60421=>"001001111",
  60422=>"111110000",
  60423=>"111111111",
  60424=>"000001001",
  60425=>"000100010",
  60426=>"110110110",
  60427=>"010000000",
  60428=>"000000000",
  60429=>"000000111",
  60430=>"111110111",
  60431=>"000000111",
  60432=>"111011000",
  60433=>"110111111",
  60434=>"111110111",
  60435=>"000000000",
  60436=>"100110111",
  60437=>"000000000",
  60438=>"111111010",
  60439=>"010111011",
  60440=>"101001111",
  60441=>"000000000",
  60442=>"100000111",
  60443=>"000001011",
  60444=>"111111000",
  60445=>"110010101",
  60446=>"101111111",
  60447=>"010010000",
  60448=>"011111111",
  60449=>"110000000",
  60450=>"111111111",
  60451=>"000000000",
  60452=>"000000000",
  60453=>"100110000",
  60454=>"000000001",
  60455=>"100100100",
  60456=>"100100001",
  60457=>"001001100",
  60458=>"011011001",
  60459=>"011101000",
  60460=>"111110100",
  60461=>"110000000",
  60462=>"111111111",
  60463=>"111011111",
  60464=>"000010111",
  60465=>"000000111",
  60466=>"101001000",
  60467=>"110110110",
  60468=>"111111011",
  60469=>"000001000",
  60470=>"111000100",
  60471=>"000001101",
  60472=>"111111111",
  60473=>"000000111",
  60474=>"011001101",
  60475=>"000000000",
  60476=>"101101001",
  60477=>"111111111",
  60478=>"000000000",
  60479=>"000010001",
  60480=>"101111011",
  60481=>"101111000",
  60482=>"001000001",
  60483=>"001000110",
  60484=>"110111111",
  60485=>"111111101",
  60486=>"000000001",
  60487=>"001111111",
  60488=>"010000100",
  60489=>"110110000",
  60490=>"101000000",
  60491=>"111101110",
  60492=>"000000000",
  60493=>"000000011",
  60494=>"000110110",
  60495=>"010111111",
  60496=>"111110111",
  60497=>"110110000",
  60498=>"000000000",
  60499=>"011011111",
  60500=>"000000000",
  60501=>"100100100",
  60502=>"110110110",
  60503=>"011111111",
  60504=>"100000000",
  60505=>"100100010",
  60506=>"011001000",
  60507=>"100000000",
  60508=>"001111011",
  60509=>"001011110",
  60510=>"000000111",
  60511=>"000000110",
  60512=>"101000101",
  60513=>"010110110",
  60514=>"101111111",
  60515=>"110110000",
  60516=>"100010010",
  60517=>"111111111",
  60518=>"011000001",
  60519=>"100000001",
  60520=>"110111111",
  60521=>"011110010",
  60522=>"001001000",
  60523=>"110000000",
  60524=>"100111111",
  60525=>"000011001",
  60526=>"010000000",
  60527=>"000000000",
  60528=>"110110110",
  60529=>"111111000",
  60530=>"110011011",
  60531=>"000000000",
  60532=>"000000100",
  60533=>"000000100",
  60534=>"111111101",
  60535=>"100000011",
  60536=>"000000000",
  60537=>"000001000",
  60538=>"000000000",
  60539=>"011111111",
  60540=>"100111111",
  60541=>"001000001",
  60542=>"000000000",
  60543=>"000010111",
  60544=>"000111101",
  60545=>"111111000",
  60546=>"000000100",
  60547=>"111101111",
  60548=>"001000000",
  60549=>"000000111",
  60550=>"011111110",
  60551=>"010010011",
  60552=>"011011111",
  60553=>"110110100",
  60554=>"010111010",
  60555=>"000000111",
  60556=>"000000000",
  60557=>"000000000",
  60558=>"111011011",
  60559=>"101100100",
  60560=>"001011001",
  60561=>"011011000",
  60562=>"000000000",
  60563=>"000000001",
  60564=>"010010010",
  60565=>"000000000",
  60566=>"111011111",
  60567=>"110100100",
  60568=>"010000000",
  60569=>"111000000",
  60570=>"000000000",
  60571=>"111111111",
  60572=>"001100100",
  60573=>"000001111",
  60574=>"000111000",
  60575=>"101000100",
  60576=>"011101010",
  60577=>"111111001",
  60578=>"111111111",
  60579=>"010000010",
  60580=>"010111100",
  60581=>"111111101",
  60582=>"100000010",
  60583=>"101000001",
  60584=>"000000100",
  60585=>"011001101",
  60586=>"001000101",
  60587=>"111000100",
  60588=>"001001111",
  60589=>"111101111",
  60590=>"111111111",
  60591=>"010111001",
  60592=>"000000001",
  60593=>"011111100",
  60594=>"011111011",
  60595=>"000011001",
  60596=>"111001000",
  60597=>"011111110",
  60598=>"000000100",
  60599=>"001111111",
  60600=>"111111000",
  60601=>"010000100",
  60602=>"010000000",
  60603=>"000000000",
  60604=>"000000000",
  60605=>"110111001",
  60606=>"000000100",
  60607=>"111111010",
  60608=>"010010000",
  60609=>"000000111",
  60610=>"100111110",
  60611=>"111001101",
  60612=>"000000111",
  60613=>"111111100",
  60614=>"010111111",
  60615=>"001101111",
  60616=>"000000101",
  60617=>"111001001",
  60618=>"101001000",
  60619=>"110000000",
  60620=>"010000000",
  60621=>"000110111",
  60622=>"111111110",
  60623=>"111111001",
  60624=>"000000000",
  60625=>"111011111",
  60626=>"010010101",
  60627=>"111110101",
  60628=>"000000111",
  60629=>"111111001",
  60630=>"110000111",
  60631=>"010111111",
  60632=>"000110110",
  60633=>"000000001",
  60634=>"000101000",
  60635=>"001001111",
  60636=>"111110110",
  60637=>"011011000",
  60638=>"000000001",
  60639=>"011101111",
  60640=>"111000000",
  60641=>"111111000",
  60642=>"000111100",
  60643=>"101111011",
  60644=>"000000000",
  60645=>"000010000",
  60646=>"000101101",
  60647=>"110110111",
  60648=>"000000000",
  60649=>"111001000",
  60650=>"110111000",
  60651=>"111111111",
  60652=>"011000001",
  60653=>"000000000",
  60654=>"000000000",
  60655=>"001101111",
  60656=>"000000100",
  60657=>"010111010",
  60658=>"000111111",
  60659=>"110010001",
  60660=>"001111111",
  60661=>"111111101",
  60662=>"111000000",
  60663=>"100000000",
  60664=>"001001000",
  60665=>"111110000",
  60666=>"111111110",
  60667=>"110101000",
  60668=>"000000100",
  60669=>"111111000",
  60670=>"000000110",
  60671=>"111111111",
  60672=>"100000100",
  60673=>"111111111",
  60674=>"010010101",
  60675=>"000000000",
  60676=>"001110010",
  60677=>"000000001",
  60678=>"100101100",
  60679=>"101010111",
  60680=>"000001011",
  60681=>"011010111",
  60682=>"110111001",
  60683=>"000000000",
  60684=>"000000110",
  60685=>"101000100",
  60686=>"011010010",
  60687=>"111000000",
  60688=>"111111111",
  60689=>"111111000",
  60690=>"101111111",
  60691=>"111110111",
  60692=>"000111010",
  60693=>"000000111",
  60694=>"111111111",
  60695=>"010111111",
  60696=>"111000000",
  60697=>"111111111",
  60698=>"111000111",
  60699=>"010010000",
  60700=>"110000010",
  60701=>"000000000",
  60702=>"000110111",
  60703=>"111111111",
  60704=>"111001001",
  60705=>"011000010",
  60706=>"100111100",
  60707=>"011000000",
  60708=>"110110100",
  60709=>"000000000",
  60710=>"000000111",
  60711=>"111111110",
  60712=>"000111000",
  60713=>"000100111",
  60714=>"000110110",
  60715=>"000000100",
  60716=>"000110111",
  60717=>"111100000",
  60718=>"111000000",
  60719=>"000011011",
  60720=>"111110001",
  60721=>"000100101",
  60722=>"111001000",
  60723=>"111111001",
  60724=>"010110010",
  60725=>"000011111",
  60726=>"111111110",
  60727=>"101001101",
  60728=>"001101110",
  60729=>"000000000",
  60730=>"000000111",
  60731=>"111111111",
  60732=>"000000001",
  60733=>"000010111",
  60734=>"001000111",
  60735=>"100000011",
  60736=>"111111101",
  60737=>"000000000",
  60738=>"101101101",
  60739=>"110100010",
  60740=>"101101111",
  60741=>"100100000",
  60742=>"000000000",
  60743=>"101001101",
  60744=>"001000000",
  60745=>"000000110",
  60746=>"101100000",
  60747=>"000000000",
  60748=>"000000110",
  60749=>"001111001",
  60750=>"000000000",
  60751=>"111111000",
  60752=>"000110000",
  60753=>"111110000",
  60754=>"111111111",
  60755=>"001110110",
  60756=>"001010000",
  60757=>"000000010",
  60758=>"011111011",
  60759=>"000001000",
  60760=>"101101111",
  60761=>"011110111",
  60762=>"010100100",
  60763=>"000100110",
  60764=>"111111101",
  60765=>"111100100",
  60766=>"000111111",
  60767=>"011001011",
  60768=>"000000111",
  60769=>"000100000",
  60770=>"001000111",
  60771=>"010011001",
  60772=>"101001001",
  60773=>"001111100",
  60774=>"111111111",
  60775=>"111111111",
  60776=>"000000001",
  60777=>"011111111",
  60778=>"111010111",
  60779=>"010101100",
  60780=>"000000000",
  60781=>"000000000",
  60782=>"001000000",
  60783=>"000101111",
  60784=>"001011011",
  60785=>"001000000",
  60786=>"111111011",
  60787=>"000000010",
  60788=>"111111100",
  60789=>"111000010",
  60790=>"000000011",
  60791=>"001001100",
  60792=>"110000000",
  60793=>"111111101",
  60794=>"010010000",
  60795=>"111100111",
  60796=>"000000001",
  60797=>"100001011",
  60798=>"000000010",
  60799=>"001000111",
  60800=>"000111111",
  60801=>"000000000",
  60802=>"000000000",
  60803=>"100000111",
  60804=>"100110111",
  60805=>"111111010",
  60806=>"000000000",
  60807=>"001000000",
  60808=>"111100010",
  60809=>"111111111",
  60810=>"111111100",
  60811=>"101111111",
  60812=>"001000111",
  60813=>"111111111",
  60814=>"000011011",
  60815=>"001000111",
  60816=>"001011100",
  60817=>"111001000",
  60818=>"000000010",
  60819=>"001000000",
  60820=>"001000000",
  60821=>"010111000",
  60822=>"110000110",
  60823=>"000000001",
  60824=>"001101000",
  60825=>"101101111",
  60826=>"111000110",
  60827=>"110010000",
  60828=>"000000000",
  60829=>"000000000",
  60830=>"000100000",
  60831=>"000000110",
  60832=>"000000000",
  60833=>"001000000",
  60834=>"101100010",
  60835=>"111001100",
  60836=>"000001111",
  60837=>"001011011",
  60838=>"110111111",
  60839=>"000000111",
  60840=>"010111111",
  60841=>"000000110",
  60842=>"100100111",
  60843=>"000110000",
  60844=>"110111111",
  60845=>"101101111",
  60846=>"000000000",
  60847=>"110000110",
  60848=>"111100000",
  60849=>"001000100",
  60850=>"110111100",
  60851=>"100110111",
  60852=>"110100100",
  60853=>"111000111",
  60854=>"110111111",
  60855=>"100010011",
  60856=>"000000000",
  60857=>"000000000",
  60858=>"111111000",
  60859=>"111000000",
  60860=>"001000010",
  60861=>"011111001",
  60862=>"111001110",
  60863=>"000100100",
  60864=>"001000111",
  60865=>"111000000",
  60866=>"010010000",
  60867=>"000000110",
  60868=>"000000101",
  60869=>"100110111",
  60870=>"000111101",
  60871=>"001010011",
  60872=>"101101111",
  60873=>"000000000",
  60874=>"110111111",
  60875=>"011000111",
  60876=>"111000000",
  60877=>"000010110",
  60878=>"000010101",
  60879=>"111100111",
  60880=>"000000110",
  60881=>"000000000",
  60882=>"000000111",
  60883=>"110110010",
  60884=>"101101111",
  60885=>"001000000",
  60886=>"011101111",
  60887=>"111101001",
  60888=>"001001111",
  60889=>"000000000",
  60890=>"000000010",
  60891=>"000000111",
  60892=>"100111111",
  60893=>"000000000",
  60894=>"000111000",
  60895=>"101111111",
  60896=>"000000000",
  60897=>"111111111",
  60898=>"100101000",
  60899=>"011001010",
  60900=>"101000000",
  60901=>"111110101",
  60902=>"000000010",
  60903=>"000000001",
  60904=>"011000011",
  60905=>"111011101",
  60906=>"011110000",
  60907=>"111111111",
  60908=>"001001111",
  60909=>"000000111",
  60910=>"110000000",
  60911=>"100000111",
  60912=>"000000111",
  60913=>"010001001",
  60914=>"000110101",
  60915=>"011011010",
  60916=>"000000010",
  60917=>"101101000",
  60918=>"101000010",
  60919=>"110111111",
  60920=>"110010011",
  60921=>"001000011",
  60922=>"111111111",
  60923=>"001000000",
  60924=>"111111000",
  60925=>"111000000",
  60926=>"101010101",
  60927=>"000000010",
  60928=>"111011111",
  60929=>"110000000",
  60930=>"000111111",
  60931=>"000111000",
  60932=>"011000101",
  60933=>"100111100",
  60934=>"000000111",
  60935=>"111010100",
  60936=>"000000111",
  60937=>"000101000",
  60938=>"011011001",
  60939=>"101101111",
  60940=>"000000111",
  60941=>"000000000",
  60942=>"110010000",
  60943=>"100111101",
  60944=>"111010000",
  60945=>"111000000",
  60946=>"111000000",
  60947=>"000000000",
  60948=>"101011111",
  60949=>"111101000",
  60950=>"000000000",
  60951=>"111001101",
  60952=>"010000000",
  60953=>"111011000",
  60954=>"000000000",
  60955=>"011111000",
  60956=>"111110000",
  60957=>"010111000",
  60958=>"000011111",
  60959=>"000111111",
  60960=>"111000000",
  60961=>"111010000",
  60962=>"100110111",
  60963=>"000000111",
  60964=>"100000100",
  60965=>"111111000",
  60966=>"111000000",
  60967=>"000000011",
  60968=>"000000000",
  60969=>"111000111",
  60970=>"010000000",
  60971=>"000100111",
  60972=>"111011000",
  60973=>"010000000",
  60974=>"111000100",
  60975=>"001000100",
  60976=>"000001000",
  60977=>"111110100",
  60978=>"111011111",
  60979=>"111010000",
  60980=>"001000100",
  60981=>"000000000",
  60982=>"000101111",
  60983=>"111101000",
  60984=>"000010011",
  60985=>"111000000",
  60986=>"100000000",
  60987=>"000000000",
  60988=>"010110001",
  60989=>"010100100",
  60990=>"000000000",
  60991=>"011011000",
  60992=>"011110111",
  60993=>"111010001",
  60994=>"000100000",
  60995=>"001001111",
  60996=>"000111010",
  60997=>"111101101",
  60998=>"000000000",
  60999=>"000111111",
  61000=>"111100000",
  61001=>"111000000",
  61002=>"101000000",
  61003=>"111000000",
  61004=>"101000000",
  61005=>"011001001",
  61006=>"111001100",
  61007=>"111101010",
  61008=>"100000000",
  61009=>"111000111",
  61010=>"010111111",
  61011=>"001101000",
  61012=>"110001000",
  61013=>"101000000",
  61014=>"000000000",
  61015=>"100111000",
  61016=>"011110111",
  61017=>"111000011",
  61018=>"011100100",
  61019=>"111010000",
  61020=>"111010000",
  61021=>"010000000",
  61022=>"000000111",
  61023=>"100100111",
  61024=>"000000010",
  61025=>"011000000",
  61026=>"000111111",
  61027=>"110001001",
  61028=>"111001001",
  61029=>"000011000",
  61030=>"010000000",
  61031=>"111000000",
  61032=>"000111110",
  61033=>"111010000",
  61034=>"010011000",
  61035=>"111110111",
  61036=>"111111111",
  61037=>"111000100",
  61038=>"000000000",
  61039=>"111010000",
  61040=>"011000100",
  61041=>"111000010",
  61042=>"000111110",
  61043=>"010000000",
  61044=>"111001000",
  61045=>"101000000",
  61046=>"100111100",
  61047=>"000000001",
  61048=>"000000011",
  61049=>"010010000",
  61050=>"101101000",
  61051=>"101100110",
  61052=>"101011110",
  61053=>"110001000",
  61054=>"000110010",
  61055=>"001111111",
  61056=>"000010000",
  61057=>"000001111",
  61058=>"000000111",
  61059=>"111000000",
  61060=>"111000000",
  61061=>"011000100",
  61062=>"110011001",
  61063=>"111000000",
  61064=>"110100000",
  61065=>"100110110",
  61066=>"111000000",
  61067=>"010011000",
  61068=>"000000010",
  61069=>"100110110",
  61070=>"000000000",
  61071=>"111001000",
  61072=>"011000001",
  61073=>"010111111",
  61074=>"001000000",
  61075=>"111101101",
  61076=>"111100011",
  61077=>"100000000",
  61078=>"111011111",
  61079=>"100100101",
  61080=>"100000000",
  61081=>"000000111",
  61082=>"010100000",
  61083=>"000001111",
  61084=>"000000011",
  61085=>"100000000",
  61086=>"010101100",
  61087=>"101101111",
  61088=>"000001011",
  61089=>"011000111",
  61090=>"011011000",
  61091=>"111001111",
  61092=>"000000100",
  61093=>"111000000",
  61094=>"000101111",
  61095=>"111001100",
  61096=>"101101000",
  61097=>"000000000",
  61098=>"101111111",
  61099=>"000101010",
  61100=>"100001000",
  61101=>"001100010",
  61102=>"111001011",
  61103=>"001010001",
  61104=>"100001111",
  61105=>"111001101",
  61106=>"000011111",
  61107=>"000000011",
  61108=>"111000000",
  61109=>"010110001",
  61110=>"101000000",
  61111=>"111110100",
  61112=>"110011010",
  61113=>"111111010",
  61114=>"010001000",
  61115=>"000101111",
  61116=>"111000000",
  61117=>"000111111",
  61118=>"100101101",
  61119=>"111000000",
  61120=>"010001011",
  61121=>"110000000",
  61122=>"110111000",
  61123=>"111000000",
  61124=>"000000000",
  61125=>"011001000",
  61126=>"111010111",
  61127=>"100111111",
  61128=>"000000000",
  61129=>"100000000",
  61130=>"111100000",
  61131=>"001001111",
  61132=>"011000000",
  61133=>"001000001",
  61134=>"010100100",
  61135=>"000110010",
  61136=>"010000110",
  61137=>"110001011",
  61138=>"001100000",
  61139=>"000001000",
  61140=>"101000111",
  61141=>"011001000",
  61142=>"001001011",
  61143=>"111111001",
  61144=>"011000111",
  61145=>"000010000",
  61146=>"000010111",
  61147=>"100000010",
  61148=>"010000000",
  61149=>"111111100",
  61150=>"111000100",
  61151=>"111111001",
  61152=>"000000000",
  61153=>"101101010",
  61154=>"000101111",
  61155=>"011011111",
  61156=>"010000000",
  61157=>"010111111",
  61158=>"000000111",
  61159=>"010011110",
  61160=>"010111101",
  61161=>"000000000",
  61162=>"111110100",
  61163=>"100101010",
  61164=>"100111111",
  61165=>"111111000",
  61166=>"001000000",
  61167=>"100000000",
  61168=>"001111111",
  61169=>"101101000",
  61170=>"111000010",
  61171=>"111000000",
  61172=>"111000010",
  61173=>"011001100",
  61174=>"111100000",
  61175=>"111000000",
  61176=>"000010111",
  61177=>"010111111",
  61178=>"111000100",
  61179=>"111111000",
  61180=>"011000100",
  61181=>"100000000",
  61182=>"011001000",
  61183=>"111011011",
  61184=>"001101010",
  61185=>"110000000",
  61186=>"111010010",
  61187=>"101101111",
  61188=>"000111110",
  61189=>"001001100",
  61190=>"111110000",
  61191=>"110001111",
  61192=>"110011000",
  61193=>"110110011",
  61194=>"001101010",
  61195=>"000001000",
  61196=>"101000000",
  61197=>"100111000",
  61198=>"011000010",
  61199=>"010110111",
  61200=>"000001101",
  61201=>"000010111",
  61202=>"000000001",
  61203=>"001001000",
  61204=>"100000000",
  61205=>"110110000",
  61206=>"111011001",
  61207=>"000000110",
  61208=>"111101101",
  61209=>"001011011",
  61210=>"111111000",
  61211=>"111111000",
  61212=>"000000111",
  61213=>"111111000",
  61214=>"111111111",
  61215=>"111010000",
  61216=>"111101111",
  61217=>"100100000",
  61218=>"000111111",
  61219=>"010010111",
  61220=>"010110000",
  61221=>"000000010",
  61222=>"111111000",
  61223=>"000010111",
  61224=>"001000000",
  61225=>"000111100",
  61226=>"000000111",
  61227=>"011111001",
  61228=>"111100110",
  61229=>"101001101",
  61230=>"000010111",
  61231=>"111010000",
  61232=>"000111010",
  61233=>"111111000",
  61234=>"000010111",
  61235=>"001111111",
  61236=>"111111010",
  61237=>"000000000",
  61238=>"111000000",
  61239=>"010011010",
  61240=>"000000111",
  61241=>"111100000",
  61242=>"100100101",
  61243=>"000001000",
  61244=>"100000000",
  61245=>"101111111",
  61246=>"110000000",
  61247=>"000000000",
  61248=>"111111111",
  61249=>"110111111",
  61250=>"100100110",
  61251=>"001000000",
  61252=>"010100010",
  61253=>"001011101",
  61254=>"000000000",
  61255=>"111111101",
  61256=>"000000000",
  61257=>"111111000",
  61258=>"111111111",
  61259=>"000000100",
  61260=>"011110010",
  61261=>"111000000",
  61262=>"110101100",
  61263=>"011010000",
  61264=>"111111010",
  61265=>"000111111",
  61266=>"111111111",
  61267=>"111010010",
  61268=>"111000000",
  61269=>"000000001",
  61270=>"011111000",
  61271=>"000010010",
  61272=>"111111111",
  61273=>"001011001",
  61274=>"111111000",
  61275=>"011111111",
  61276=>"111000111",
  61277=>"001001001",
  61278=>"010010000",
  61279=>"111000000",
  61280=>"111111011",
  61281=>"000111000",
  61282=>"001000000",
  61283=>"111111000",
  61284=>"110100000",
  61285=>"111000001",
  61286=>"111101111",
  61287=>"111111000",
  61288=>"101000001",
  61289=>"000000111",
  61290=>"101111111",
  61291=>"000010000",
  61292=>"110101000",
  61293=>"000000000",
  61294=>"000010010",
  61295=>"111111000",
  61296=>"111111000",
  61297=>"000101111",
  61298=>"111001000",
  61299=>"000010010",
  61300=>"001000111",
  61301=>"001000111",
  61302=>"111101000",
  61303=>"000111011",
  61304=>"000010000",
  61305=>"100000110",
  61306=>"000111000",
  61307=>"111111111",
  61308=>"000000000",
  61309=>"100100000",
  61310=>"001000010",
  61311=>"110001000",
  61312=>"111111010",
  61313=>"011111110",
  61314=>"010001000",
  61315=>"011101111",
  61316=>"010111110",
  61317=>"000000100",
  61318=>"001000000",
  61319=>"110000000",
  61320=>"111011001",
  61321=>"000111000",
  61322=>"000000000",
  61323=>"100111011",
  61324=>"111011110",
  61325=>"010000000",
  61326=>"111001101",
  61327=>"011001011",
  61328=>"110111101",
  61329=>"111011000",
  61330=>"000000111",
  61331=>"110000000",
  61332=>"111111000",
  61333=>"000000010",
  61334=>"111001000",
  61335=>"001111001",
  61336=>"111111111",
  61337=>"000000111",
  61338=>"110110000",
  61339=>"111111001",
  61340=>"010111111",
  61341=>"001000111",
  61342=>"100111111",
  61343=>"001100110",
  61344=>"001000000",
  61345=>"110111111",
  61346=>"111001000",
  61347=>"111111110",
  61348=>"001000000",
  61349=>"111011000",
  61350=>"000111011",
  61351=>"001000000",
  61352=>"000000111",
  61353=>"110111101",
  61354=>"111111000",
  61355=>"001000000",
  61356=>"110000000",
  61357=>"010111110",
  61358=>"110100100",
  61359=>"110010000",
  61360=>"111111100",
  61361=>"011000000",
  61362=>"101001100",
  61363=>"101101110",
  61364=>"110100100",
  61365=>"001000000",
  61366=>"011000001",
  61367=>"001111111",
  61368=>"011000000",
  61369=>"010001000",
  61370=>"110111111",
  61371=>"010011010",
  61372=>"001101110",
  61373=>"100000000",
  61374=>"011101000",
  61375=>"001011111",
  61376=>"111010010",
  61377=>"101111010",
  61378=>"111000001",
  61379=>"110000100",
  61380=>"000000111",
  61381=>"100101001",
  61382=>"110110111",
  61383=>"111111000",
  61384=>"000000000",
  61385=>"111111000",
  61386=>"111111001",
  61387=>"111001111",
  61388=>"111010000",
  61389=>"111000000",
  61390=>"111000000",
  61391=>"111011000",
  61392=>"111111111",
  61393=>"100011001",
  61394=>"111111001",
  61395=>"111111000",
  61396=>"111110000",
  61397=>"111000000",
  61398=>"010111000",
  61399=>"000000000",
  61400=>"011000000",
  61401=>"110111010",
  61402=>"110111110",
  61403=>"000000111",
  61404=>"111100000",
  61405=>"010110111",
  61406=>"010011111",
  61407=>"000000000",
  61408=>"010010000",
  61409=>"111111111",
  61410=>"100000000",
  61411=>"100111000",
  61412=>"000000000",
  61413=>"001001000",
  61414=>"000000001",
  61415=>"011111010",
  61416=>"111111111",
  61417=>"011000100",
  61418=>"101100000",
  61419=>"111111000",
  61420=>"110111111",
  61421=>"000000000",
  61422=>"000111111",
  61423=>"011001011",
  61424=>"000000000",
  61425=>"001110100",
  61426=>"000010010",
  61427=>"111111100",
  61428=>"101111001",
  61429=>"111111001",
  61430=>"110000000",
  61431=>"100111000",
  61432=>"000000110",
  61433=>"001000000",
  61434=>"101111000",
  61435=>"111010000",
  61436=>"001000000",
  61437=>"000000000",
  61438=>"111110000",
  61439=>"000000000",
  61440=>"011011011",
  61441=>"000011110",
  61442=>"010000111",
  61443=>"000001000",
  61444=>"000000100",
  61445=>"110011000",
  61446=>"000100000",
  61447=>"100110110",
  61448=>"111111000",
  61449=>"110000000",
  61450=>"100000000",
  61451=>"111010011",
  61452=>"000000000",
  61453=>"000101111",
  61454=>"111001000",
  61455=>"000001101",
  61456=>"000110010",
  61457=>"110000000",
  61458=>"000001101",
  61459=>"010110111",
  61460=>"110110100",
  61461=>"111010110",
  61462=>"001100100",
  61463=>"000011011",
  61464=>"010000000",
  61465=>"110001000",
  61466=>"111110000",
  61467=>"101010000",
  61468=>"110111010",
  61469=>"000111111",
  61470=>"010101000",
  61471=>"001000111",
  61472=>"011001001",
  61473=>"110111000",
  61474=>"000010111",
  61475=>"111111001",
  61476=>"000000000",
  61477=>"111110110",
  61478=>"101010000",
  61479=>"111111101",
  61480=>"011010111",
  61481=>"110111111",
  61482=>"010110000",
  61483=>"010000111",
  61484=>"111011110",
  61485=>"000111111",
  61486=>"000011101",
  61487=>"000100110",
  61488=>"000010010",
  61489=>"100011111",
  61490=>"101000001",
  61491=>"111111000",
  61492=>"000000010",
  61493=>"111010000",
  61494=>"110010000",
  61495=>"001011000",
  61496=>"000111101",
  61497=>"101001000",
  61498=>"000101101",
  61499=>"000000110",
  61500=>"000011111",
  61501=>"101111111",
  61502=>"000000000",
  61503=>"000100111",
  61504=>"111001000",
  61505=>"111000100",
  61506=>"111111111",
  61507=>"001000011",
  61508=>"010011011",
  61509=>"000010010",
  61510=>"110110001",
  61511=>"110000111",
  61512=>"000011111",
  61513=>"010011000",
  61514=>"000110111",
  61515=>"011101000",
  61516=>"000000000",
  61517=>"011000000",
  61518=>"001111111",
  61519=>"110111000",
  61520=>"111000110",
  61521=>"010010011",
  61522=>"111111110",
  61523=>"001100001",
  61524=>"110110110",
  61525=>"001101100",
  61526=>"000000011",
  61527=>"111010001",
  61528=>"000111110",
  61529=>"000111111",
  61530=>"101000011",
  61531=>"100100101",
  61532=>"010101000",
  61533=>"000001111",
  61534=>"000010011",
  61535=>"000100100",
  61536=>"111110000",
  61537=>"101101011",
  61538=>"110000001",
  61539=>"000110110",
  61540=>"101000001",
  61541=>"001001101",
  61542=>"110100000",
  61543=>"111110110",
  61544=>"000111110",
  61545=>"000101101",
  61546=>"010110111",
  61547=>"110000000",
  61548=>"000111110",
  61549=>"110010000",
  61550=>"010110000",
  61551=>"010111000",
  61552=>"001010101",
  61553=>"000101001",
  61554=>"011000000",
  61555=>"010010001",
  61556=>"111111000",
  61557=>"000010111",
  61558=>"111111101",
  61559=>"111000001",
  61560=>"010110001",
  61561=>"010000111",
  61562=>"101110000",
  61563=>"000111111",
  61564=>"001001010",
  61565=>"100000100",
  61566=>"100000000",
  61567=>"101000111",
  61568=>"000111000",
  61569=>"001000011",
  61570=>"110000101",
  61571=>"000100111",
  61572=>"111110010",
  61573=>"101001000",
  61574=>"011000111",
  61575=>"011001001",
  61576=>"000001110",
  61577=>"111111110",
  61578=>"000010010",
  61579=>"010000100",
  61580=>"111000111",
  61581=>"100001001",
  61582=>"000000000",
  61583=>"000000001",
  61584=>"000000100",
  61585=>"101101001",
  61586=>"100001110",
  61587=>"001000000",
  61588=>"000101100",
  61589=>"111111000",
  61590=>"111111000",
  61591=>"100001000",
  61592=>"011000111",
  61593=>"010110000",
  61594=>"110000111",
  61595=>"000000000",
  61596=>"110010000",
  61597=>"000011010",
  61598=>"111101001",
  61599=>"010000001",
  61600=>"001101011",
  61601=>"111111000",
  61602=>"000000001",
  61603=>"111110101",
  61604=>"010011000",
  61605=>"000001110",
  61606=>"100111011",
  61607=>"111111000",
  61608=>"000110110",
  61609=>"000111110",
  61610=>"000000111",
  61611=>"110010110",
  61612=>"110110110",
  61613=>"111000101",
  61614=>"111100110",
  61615=>"110111001",
  61616=>"000000001",
  61617=>"100100010",
  61618=>"001101111",
  61619=>"011100101",
  61620=>"100101011",
  61621=>"010110011",
  61622=>"010010111",
  61623=>"011111101",
  61624=>"001100111",
  61625=>"000100001",
  61626=>"010000011",
  61627=>"010111111",
  61628=>"010010111",
  61629=>"100000111",
  61630=>"001001110",
  61631=>"000000010",
  61632=>"010000000",
  61633=>"111001000",
  61634=>"110111110",
  61635=>"001100111",
  61636=>"101000000",
  61637=>"011001111",
  61638=>"111111010",
  61639=>"111001000",
  61640=>"000000100",
  61641=>"000000010",
  61642=>"000010111",
  61643=>"000000000",
  61644=>"111111000",
  61645=>"101101000",
  61646=>"111000111",
  61647=>"000111000",
  61648=>"010010111",
  61649=>"001001110",
  61650=>"010101011",
  61651=>"000000001",
  61652=>"001100000",
  61653=>"000000110",
  61654=>"000110110",
  61655=>"111111110",
  61656=>"000000000",
  61657=>"011111110",
  61658=>"000101101",
  61659=>"000000001",
  61660=>"000111110",
  61661=>"110111110",
  61662=>"000110111",
  61663=>"010101000",
  61664=>"111000000",
  61665=>"111111010",
  61666=>"000000010",
  61667=>"100101011",
  61668=>"000000001",
  61669=>"000000010",
  61670=>"111001000",
  61671=>"111110111",
  61672=>"111111000",
  61673=>"000110101",
  61674=>"000000000",
  61675=>"000000011",
  61676=>"000001001",
  61677=>"001000111",
  61678=>"000000001",
  61679=>"000000000",
  61680=>"010010111",
  61681=>"110000100",
  61682=>"100011011",
  61683=>"001011110",
  61684=>"100101001",
  61685=>"001000110",
  61686=>"000000111",
  61687=>"000000110",
  61688=>"110001001",
  61689=>"111111000",
  61690=>"000111111",
  61691=>"111001110",
  61692=>"001001101",
  61693=>"000010111",
  61694=>"000001010",
  61695=>"011110111",
  61696=>"001001100",
  61697=>"000000000",
  61698=>"001001001",
  61699=>"001000001",
  61700=>"100000100",
  61701=>"111111111",
  61702=>"101001101",
  61703=>"001101000",
  61704=>"000100000",
  61705=>"000110110",
  61706=>"100110010",
  61707=>"110011000",
  61708=>"001001111",
  61709=>"011111100",
  61710=>"101111010",
  61711=>"101111000",
  61712=>"110010000",
  61713=>"000010000",
  61714=>"000110110",
  61715=>"101001011",
  61716=>"000011111",
  61717=>"000111110",
  61718=>"001001111",
  61719=>"001001111",
  61720=>"000000001",
  61721=>"110001010",
  61722=>"110100111",
  61723=>"110110010",
  61724=>"001000000",
  61725=>"001001111",
  61726=>"111001010",
  61727=>"000000111",
  61728=>"011110111",
  61729=>"001001111",
  61730=>"111101001",
  61731=>"001101111",
  61732=>"011001000",
  61733=>"111111011",
  61734=>"000011010",
  61735=>"001111001",
  61736=>"110011011",
  61737=>"100110000",
  61738=>"110111000",
  61739=>"001000110",
  61740=>"110111110",
  61741=>"000000111",
  61742=>"111111111",
  61743=>"010000000",
  61744=>"000000111",
  61745=>"101000000",
  61746=>"110001000",
  61747=>"101110111",
  61748=>"110110001",
  61749=>"011110000",
  61750=>"010110001",
  61751=>"110000000",
  61752=>"110001111",
  61753=>"100000000",
  61754=>"000000000",
  61755=>"000101111",
  61756=>"111111100",
  61757=>"001001011",
  61758=>"000001111",
  61759=>"110110000",
  61760=>"100100101",
  61761=>"001000000",
  61762=>"000111011",
  61763=>"110110000",
  61764=>"001001111",
  61765=>"100110000",
  61766=>"000111000",
  61767=>"001001111",
  61768=>"110111111",
  61769=>"110010111",
  61770=>"101000000",
  61771=>"000000110",
  61772=>"111111000",
  61773=>"111000000",
  61774=>"011001000",
  61775=>"111000001",
  61776=>"001001000",
  61777=>"110111111",
  61778=>"001110110",
  61779=>"111001000",
  61780=>"001001000",
  61781=>"111111110",
  61782=>"001001110",
  61783=>"110111111",
  61784=>"000000010",
  61785=>"100101000",
  61786=>"001110011",
  61787=>"101101100",
  61788=>"110000111",
  61789=>"100000100",
  61790=>"110110000",
  61791=>"110110000",
  61792=>"010000000",
  61793=>"110110111",
  61794=>"000000111",
  61795=>"010100110",
  61796=>"111001011",
  61797=>"111101110",
  61798=>"110110011",
  61799=>"110010000",
  61800=>"000110100",
  61801=>"111111010",
  61802=>"110110000",
  61803=>"100100010",
  61804=>"010010011",
  61805=>"110110000",
  61806=>"000011011",
  61807=>"111011111",
  61808=>"100000000",
  61809=>"110110111",
  61810=>"101011000",
  61811=>"001000111",
  61812=>"111000010",
  61813=>"000000000",
  61814=>"100010110",
  61815=>"110111001",
  61816=>"001111000",
  61817=>"001001110",
  61818=>"000001111",
  61819=>"111111111",
  61820=>"000110011",
  61821=>"000000000",
  61822=>"000000101",
  61823=>"110000000",
  61824=>"101010000",
  61825=>"111000001",
  61826=>"110011000",
  61827=>"001000111",
  61828=>"111000000",
  61829=>"000110111",
  61830=>"110111010",
  61831=>"100110100",
  61832=>"000001000",
  61833=>"001000100",
  61834=>"110010011",
  61835=>"000110111",
  61836=>"110110000",
  61837=>"001111011",
  61838=>"000111110",
  61839=>"000000000",
  61840=>"011001001",
  61841=>"001101010",
  61842=>"000001111",
  61843=>"010000000",
  61844=>"001111111",
  61845=>"110110001",
  61846=>"110111111",
  61847=>"000011100",
  61848=>"110111001",
  61849=>"110110111",
  61850=>"000000110",
  61851=>"000000001",
  61852=>"000000101",
  61853=>"010110000",
  61854=>"000110111",
  61855=>"000000111",
  61856=>"111100110",
  61857=>"110110100",
  61858=>"111111111",
  61859=>"011001100",
  61860=>"111011010",
  61861=>"000011001",
  61862=>"001111110",
  61863=>"001111000",
  61864=>"110100010",
  61865=>"100111111",
  61866=>"001001001",
  61867=>"000000000",
  61868=>"101000111",
  61869=>"000000000",
  61870=>"011001101",
  61871=>"000011111",
  61872=>"000000000",
  61873=>"111001111",
  61874=>"111000001",
  61875=>"100100000",
  61876=>"111111000",
  61877=>"000100110",
  61878=>"100001001",
  61879=>"101111100",
  61880=>"111110111",
  61881=>"010110111",
  61882=>"110110101",
  61883=>"110010010",
  61884=>"111010010",
  61885=>"110111111",
  61886=>"011001000",
  61887=>"001000000",
  61888=>"000000111",
  61889=>"001000000",
  61890=>"000111111",
  61891=>"011001000",
  61892=>"001100000",
  61893=>"111000111",
  61894=>"110111111",
  61895=>"010010110",
  61896=>"010111101",
  61897=>"010011000",
  61898=>"000000001",
  61899=>"010011001",
  61900=>"010111000",
  61901=>"100111011",
  61902=>"000000001",
  61903=>"111011110",
  61904=>"101101111",
  61905=>"100100011",
  61906=>"000011000",
  61907=>"000000000",
  61908=>"001000001",
  61909=>"000000111",
  61910=>"000100010",
  61911=>"001000111",
  61912=>"001111111",
  61913=>"000000110",
  61914=>"111001011",
  61915=>"001000111",
  61916=>"001001110",
  61917=>"111111100",
  61918=>"000000011",
  61919=>"110111001",
  61920=>"111001010",
  61921=>"001000111",
  61922=>"101111000",
  61923=>"111100011",
  61924=>"000000111",
  61925=>"111001111",
  61926=>"111011111",
  61927=>"001001111",
  61928=>"100110111",
  61929=>"101111111",
  61930=>"011110000",
  61931=>"001001111",
  61932=>"000000010",
  61933=>"010110000",
  61934=>"000000001",
  61935=>"111010110",
  61936=>"001111111",
  61937=>"100000110",
  61938=>"111011010",
  61939=>"011011000",
  61940=>"101001111",
  61941=>"001001111",
  61942=>"100000001",
  61943=>"001001111",
  61944=>"000001000",
  61945=>"001000111",
  61946=>"110000101",
  61947=>"000111111",
  61948=>"000110000",
  61949=>"111000010",
  61950=>"000000000",
  61951=>"000000001",
  61952=>"110111011",
  61953=>"011010001",
  61954=>"001000111",
  61955=>"000000000",
  61956=>"110100100",
  61957=>"111111101",
  61958=>"111101111",
  61959=>"000111111",
  61960=>"000010000",
  61961=>"101101010",
  61962=>"001001101",
  61963=>"000000101",
  61964=>"010000111",
  61965=>"000000010",
  61966=>"110100000",
  61967=>"001111111",
  61968=>"111100110",
  61969=>"000000010",
  61970=>"111010101",
  61971=>"111101000",
  61972=>"001101010",
  61973=>"000111111",
  61974=>"111111100",
  61975=>"111101100",
  61976=>"000001000",
  61977=>"001000111",
  61978=>"101101110",
  61979=>"000000110",
  61980=>"100110111",
  61981=>"000001010",
  61982=>"111111100",
  61983=>"011000100",
  61984=>"111111010",
  61985=>"111111010",
  61986=>"011111001",
  61987=>"010111100",
  61988=>"011101100",
  61989=>"000010111",
  61990=>"010000110",
  61991=>"111001110",
  61992=>"000000110",
  61993=>"000100010",
  61994=>"000000100",
  61995=>"001000000",
  61996=>"010010001",
  61997=>"100101000",
  61998=>"001111111",
  61999=>"011001000",
  62000=>"110101000",
  62001=>"100110110",
  62002=>"000111111",
  62003=>"111111011",
  62004=>"000000111",
  62005=>"000001010",
  62006=>"001000101",
  62007=>"000111111",
  62008=>"000001100",
  62009=>"000000101",
  62010=>"001101111",
  62011=>"001001011",
  62012=>"100001011",
  62013=>"110111000",
  62014=>"111111111",
  62015=>"000100100",
  62016=>"000111111",
  62017=>"001111111",
  62018=>"111111111",
  62019=>"101101100",
  62020=>"010110111",
  62021=>"101000101",
  62022=>"000111111",
  62023=>"110100111",
  62024=>"100110101",
  62025=>"111001110",
  62026=>"111001000",
  62027=>"010100000",
  62028=>"110111111",
  62029=>"010000110",
  62030=>"111011011",
  62031=>"100010000",
  62032=>"111111000",
  62033=>"010110010",
  62034=>"001111111",
  62035=>"000001100",
  62036=>"101001111",
  62037=>"011111111",
  62038=>"111011011",
  62039=>"100100111",
  62040=>"000000000",
  62041=>"100110100",
  62042=>"011000000",
  62043=>"100100100",
  62044=>"000001001",
  62045=>"000000000",
  62046=>"110111111",
  62047=>"001000001",
  62048=>"010111000",
  62049=>"111001000",
  62050=>"111101100",
  62051=>"011001000",
  62052=>"000000000",
  62053=>"110110010",
  62054=>"111001111",
  62055=>"110100111",
  62056=>"000101111",
  62057=>"111101001",
  62058=>"000000000",
  62059=>"111111111",
  62060=>"010001000",
  62061=>"000111111",
  62062=>"000000001",
  62063=>"000000111",
  62064=>"111011001",
  62065=>"000000100",
  62066=>"100000011",
  62067=>"000001000",
  62068=>"101010110",
  62069=>"001001111",
  62070=>"000000001",
  62071=>"100010000",
  62072=>"000000111",
  62073=>"111111000",
  62074=>"000000000",
  62075=>"101101111",
  62076=>"000001001",
  62077=>"110100010",
  62078=>"000000110",
  62079=>"111000000",
  62080=>"000111111",
  62081=>"011011010",
  62082=>"101101101",
  62083=>"000010111",
  62084=>"101101000",
  62085=>"000000001",
  62086=>"000000111",
  62087=>"111100100",
  62088=>"110100100",
  62089=>"111111111",
  62090=>"101101011",
  62091=>"011000000",
  62092=>"000000000",
  62093=>"010110010",
  62094=>"000000000",
  62095=>"000000000",
  62096=>"110100000",
  62097=>"111111000",
  62098=>"110011000",
  62099=>"111100100",
  62100=>"000000000",
  62101=>"000001000",
  62102=>"010111111",
  62103=>"001011011",
  62104=>"000110111",
  62105=>"111111001",
  62106=>"100111111",
  62107=>"101100010",
  62108=>"000010110",
  62109=>"110111111",
  62110=>"000000000",
  62111=>"000000010",
  62112=>"010110101",
  62113=>"001110110",
  62114=>"010000100",
  62115=>"000001001",
  62116=>"000000001",
  62117=>"011111011",
  62118=>"000110000",
  62119=>"000000000",
  62120=>"000001011",
  62121=>"000010000",
  62122=>"001101010",
  62123=>"010000000",
  62124=>"111000110",
  62125=>"101111111",
  62126=>"110110000",
  62127=>"111111011",
  62128=>"001100000",
  62129=>"000000001",
  62130=>"111000101",
  62131=>"110000000",
  62132=>"011100000",
  62133=>"000000000",
  62134=>"100000000",
  62135=>"000000000",
  62136=>"000000100",
  62137=>"000011011",
  62138=>"000100111",
  62139=>"110111000",
  62140=>"010111111",
  62141=>"010110010",
  62142=>"001011001",
  62143=>"001111111",
  62144=>"101000001",
  62145=>"101000111",
  62146=>"000111111",
  62147=>"010000110",
  62148=>"011101011",
  62149=>"111000100",
  62150=>"110111100",
  62151=>"001000110",
  62152=>"111011110",
  62153=>"010000000",
  62154=>"001000000",
  62155=>"011111000",
  62156=>"101101000",
  62157=>"000100101",
  62158=>"000000001",
  62159=>"111111110",
  62160=>"001000111",
  62161=>"110110010",
  62162=>"001000000",
  62163=>"011111111",
  62164=>"011010110",
  62165=>"110110000",
  62166=>"000000111",
  62167=>"000000101",
  62168=>"111000000",
  62169=>"010101000",
  62170=>"000011111",
  62171=>"001001111",
  62172=>"111011001",
  62173=>"110010000",
  62174=>"000000001",
  62175=>"000000101",
  62176=>"000000101",
  62177=>"001000000",
  62178=>"101000000",
  62179=>"011011000",
  62180=>"000000000",
  62181=>"101000000",
  62182=>"000000111",
  62183=>"010111010",
  62184=>"001100101",
  62185=>"010011111",
  62186=>"101101110",
  62187=>"000000000",
  62188=>"000001000",
  62189=>"111010010",
  62190=>"000000100",
  62191=>"111111001",
  62192=>"111000011",
  62193=>"110100011",
  62194=>"001111110",
  62195=>"010111001",
  62196=>"000110010",
  62197=>"101000000",
  62198=>"101111111",
  62199=>"110100110",
  62200=>"000000010",
  62201=>"001010110",
  62202=>"010000101",
  62203=>"000000000",
  62204=>"111111010",
  62205=>"010101101",
  62206=>"000011011",
  62207=>"000010000",
  62208=>"100111100",
  62209=>"111000000",
  62210=>"101101100",
  62211=>"000001000",
  62212=>"100111111",
  62213=>"001000101",
  62214=>"000111011",
  62215=>"000000000",
  62216=>"010111000",
  62217=>"101101000",
  62218=>"101000000",
  62219=>"000000000",
  62220=>"111100000",
  62221=>"110111111",
  62222=>"000100000",
  62223=>"011000111",
  62224=>"101000000",
  62225=>"100101101",
  62226=>"100001101",
  62227=>"111100000",
  62228=>"110010000",
  62229=>"111101111",
  62230=>"100111110",
  62231=>"101101101",
  62232=>"111001100",
  62233=>"111010100",
  62234=>"111101000",
  62235=>"101101001",
  62236=>"101100111",
  62237=>"100000111",
  62238=>"101101111",
  62239=>"000111111",
  62240=>"010100000",
  62241=>"010010000",
  62242=>"100101011",
  62243=>"000000010",
  62244=>"000001111",
  62245=>"001100111",
  62246=>"101101000",
  62247=>"001000101",
  62248=>"001001100",
  62249=>"011010000",
  62250=>"111000001",
  62251=>"100100101",
  62252=>"110110111",
  62253=>"000100011",
  62254=>"111110101",
  62255=>"101001001",
  62256=>"111111110",
  62257=>"001000111",
  62258=>"101100110",
  62259=>"101001010",
  62260=>"111000101",
  62261=>"000111111",
  62262=>"111100001",
  62263=>"001111111",
  62264=>"010010111",
  62265=>"000010011",
  62266=>"001101101",
  62267=>"101101011",
  62268=>"000011111",
  62269=>"111111000",
  62270=>"000000000",
  62271=>"000100110",
  62272=>"001000000",
  62273=>"000000110",
  62274=>"011111111",
  62275=>"000000100",
  62276=>"101100010",
  62277=>"111010100",
  62278=>"101101111",
  62279=>"000010000",
  62280=>"000011101",
  62281=>"111101111",
  62282=>"000000101",
  62283=>"000111101",
  62284=>"110100111",
  62285=>"000100101",
  62286=>"000000101",
  62287=>"000101110",
  62288=>"000100100",
  62289=>"111111111",
  62290=>"010111010",
  62291=>"000101101",
  62292=>"111110000",
  62293=>"000110100",
  62294=>"000001111",
  62295=>"000101000",
  62296=>"001001110",
  62297=>"000001000",
  62298=>"000100011",
  62299=>"000001100",
  62300=>"101000010",
  62301=>"100110101",
  62302=>"010010110",
  62303=>"000000001",
  62304=>"001000100",
  62305=>"100101000",
  62306=>"101000000",
  62307=>"001011101",
  62308=>"000000001",
  62309=>"000111001",
  62310=>"110011010",
  62311=>"000010010",
  62312=>"000000010",
  62313=>"111100101",
  62314=>"001001011",
  62315=>"110111001",
  62316=>"000000000",
  62317=>"111001010",
  62318=>"000000000",
  62319=>"010110100",
  62320=>"000001111",
  62321=>"000000000",
  62322=>"101001100",
  62323=>"000101110",
  62324=>"110000000",
  62325=>"101001101",
  62326=>"001010101",
  62327=>"010010111",
  62328=>"101000000",
  62329=>"011000100",
  62330=>"000001101",
  62331=>"110110111",
  62332=>"001001000",
  62333=>"000101011",
  62334=>"001100110",
  62335=>"100000000",
  62336=>"111000000",
  62337=>"010010010",
  62338=>"100000100",
  62339=>"000110000",
  62340=>"000000011",
  62341=>"011110010",
  62342=>"000000111",
  62343=>"100100000",
  62344=>"100110101",
  62345=>"101011010",
  62346=>"000100111",
  62347=>"110111001",
  62348=>"000011010",
  62349=>"001100101",
  62350=>"000010101",
  62351=>"001001101",
  62352=>"010111110",
  62353=>"001010101",
  62354=>"111101110",
  62355=>"000000111",
  62356=>"001100010",
  62357=>"101000010",
  62358=>"110010110",
  62359=>"100100101",
  62360=>"110000000",
  62361=>"000000110",
  62362=>"101100001",
  62363=>"101101111",
  62364=>"111101010",
  62365=>"111000111",
  62366=>"001000010",
  62367=>"010000111",
  62368=>"000000111",
  62369=>"101111111",
  62370=>"111111111",
  62371=>"101100000",
  62372=>"100001000",
  62373=>"010101111",
  62374=>"011111000",
  62375=>"111011111",
  62376=>"111001110",
  62377=>"000001010",
  62378=>"111001001",
  62379=>"101000000",
  62380=>"001000000",
  62381=>"000000010",
  62382=>"001110110",
  62383=>"101110110",
  62384=>"000000000",
  62385=>"100000010",
  62386=>"000110101",
  62387=>"001001001",
  62388=>"111111000",
  62389=>"000000001",
  62390=>"100000100",
  62391=>"011000000",
  62392=>"100110111",
  62393=>"001000000",
  62394=>"111110101",
  62395=>"101101111",
  62396=>"010010000",
  62397=>"001010000",
  62398=>"000000010",
  62399=>"001111011",
  62400=>"000000011",
  62401=>"101100100",
  62402=>"111101101",
  62403=>"100001011",
  62404=>"010010000",
  62405=>"100000100",
  62406=>"000100110",
  62407=>"000100100",
  62408=>"011010111",
  62409=>"000011110",
  62410=>"011110000",
  62411=>"000010010",
  62412=>"100111111",
  62413=>"110100000",
  62414=>"111111000",
  62415=>"010010001",
  62416=>"100101011",
  62417=>"011111111",
  62418=>"101110001",
  62419=>"010111111",
  62420=>"001000000",
  62421=>"010011001",
  62422=>"110000010",
  62423=>"010000000",
  62424=>"000101111",
  62425=>"111000010",
  62426=>"011010001",
  62427=>"111101101",
  62428=>"100010000",
  62429=>"011000110",
  62430=>"111111101",
  62431=>"111111010",
  62432=>"000010110",
  62433=>"101101111",
  62434=>"101110110",
  62435=>"100001111",
  62436=>"111101100",
  62437=>"111111111",
  62438=>"110111111",
  62439=>"000011011",
  62440=>"110111101",
  62441=>"110111101",
  62442=>"111000000",
  62443=>"011011000",
  62444=>"010010000",
  62445=>"000000010",
  62446=>"000000100",
  62447=>"100101101",
  62448=>"010110000",
  62449=>"001001000",
  62450=>"000000111",
  62451=>"110110100",
  62452=>"010010001",
  62453=>"111100010",
  62454=>"100101000",
  62455=>"101100101",
  62456=>"000000000",
  62457=>"010101101",
  62458=>"111110100",
  62459=>"000011000",
  62460=>"001111111",
  62461=>"000000011",
  62462=>"001001011",
  62463=>"111001000",
  62464=>"011011001",
  62465=>"010001001",
  62466=>"001000001",
  62467=>"000000001",
  62468=>"011011011",
  62469=>"110110101",
  62470=>"000000000",
  62471=>"011000001",
  62472=>"011011110",
  62473=>"000000000",
  62474=>"100000000",
  62475=>"000111011",
  62476=>"101000111",
  62477=>"000000110",
  62478=>"001111001",
  62479=>"000111110",
  62480=>"000000111",
  62481=>"011000011",
  62482=>"000010110",
  62483=>"000100110",
  62484=>"111110011",
  62485=>"100000000",
  62486=>"110100100",
  62487=>"111000111",
  62488=>"001101100",
  62489=>"100000000",
  62490=>"101000100",
  62491=>"111111000",
  62492=>"101000000",
  62493=>"000100111",
  62494=>"111111100",
  62495=>"000000011",
  62496=>"000000000",
  62497=>"110111100",
  62498=>"001001000",
  62499=>"000000000",
  62500=>"011001100",
  62501=>"110110010",
  62502=>"011010010",
  62503=>"010011000",
  62504=>"111011000",
  62505=>"001111111",
  62506=>"101000011",
  62507=>"110110000",
  62508=>"001011011",
  62509=>"100111111",
  62510=>"000100111",
  62511=>"000000111",
  62512=>"000000111",
  62513=>"000001111",
  62514=>"101101011",
  62515=>"111000000",
  62516=>"000000000",
  62517=>"010110111",
  62518=>"110000001",
  62519=>"000000000",
  62520=>"011111111",
  62521=>"001000000",
  62522=>"100000101",
  62523=>"000000100",
  62524=>"110111011",
  62525=>"111111100",
  62526=>"000000000",
  62527=>"001111000",
  62528=>"000000001",
  62529=>"111110111",
  62530=>"000111101",
  62531=>"011010000",
  62532=>"011111100",
  62533=>"000001101",
  62534=>"111000110",
  62535=>"101111010",
  62536=>"000011010",
  62537=>"111111010",
  62538=>"111001101",
  62539=>"111000101",
  62540=>"000000000",
  62541=>"111011001",
  62542=>"010011110",
  62543=>"101000111",
  62544=>"000101111",
  62545=>"110010001",
  62546=>"111111101",
  62547=>"111001100",
  62548=>"000111000",
  62549=>"010011110",
  62550=>"111001101",
  62551=>"101101111",
  62552=>"001001110",
  62553=>"100110111",
  62554=>"110001101",
  62555=>"111110111",
  62556=>"100110001",
  62557=>"010000000",
  62558=>"101010111",
  62559=>"000001001",
  62560=>"010111010",
  62561=>"000101100",
  62562=>"110010000",
  62563=>"001000101",
  62564=>"110010011",
  62565=>"000000001",
  62566=>"111111000",
  62567=>"111000000",
  62568=>"111111100",
  62569=>"111111010",
  62570=>"110111111",
  62571=>"100000000",
  62572=>"000000011",
  62573=>"000000111",
  62574=>"001000101",
  62575=>"111101111",
  62576=>"100110011",
  62577=>"000111111",
  62578=>"010000100",
  62579=>"101111111",
  62580=>"011001011",
  62581=>"000000000",
  62582=>"111110111",
  62583=>"111111000",
  62584=>"011001101",
  62585=>"111111101",
  62586=>"001001000",
  62587=>"000000110",
  62588=>"000111011",
  62589=>"011100000",
  62590=>"010000010",
  62591=>"111010000",
  62592=>"111110101",
  62593=>"010000000",
  62594=>"110111011",
  62595=>"100000000",
  62596=>"111111101",
  62597=>"001000010",
  62598=>"011111110",
  62599=>"000100000",
  62600=>"010111100",
  62601=>"101000010",
  62602=>"100000111",
  62603=>"000000000",
  62604=>"000000000",
  62605=>"111001000",
  62606=>"000000101",
  62607=>"000000000",
  62608=>"001111110",
  62609=>"000110000",
  62610=>"111000111",
  62611=>"111101000",
  62612=>"111111000",
  62613=>"111010000",
  62614=>"000101001",
  62615=>"011111101",
  62616=>"011110100",
  62617=>"000010001",
  62618=>"000010010",
  62619=>"000000000",
  62620=>"000001010",
  62621=>"010111000",
  62622=>"111110110",
  62623=>"000000100",
  62624=>"000100000",
  62625=>"111111111",
  62626=>"110110001",
  62627=>"010000101",
  62628=>"111011100",
  62629=>"111001001",
  62630=>"000001000",
  62631=>"000110111",
  62632=>"111111000",
  62633=>"001101101",
  62634=>"000000100",
  62635=>"111101111",
  62636=>"001001100",
  62637=>"111111000",
  62638=>"100111111",
  62639=>"001100111",
  62640=>"000000000",
  62641=>"100101001",
  62642=>"010000000",
  62643=>"011000000",
  62644=>"010100100",
  62645=>"101000111",
  62646=>"000000000",
  62647=>"101110010",
  62648=>"011111110",
  62649=>"101101001",
  62650=>"010011111",
  62651=>"111111010",
  62652=>"000111100",
  62653=>"111111111",
  62654=>"100111011",
  62655=>"000101111",
  62656=>"101000000",
  62657=>"101000000",
  62658=>"111110111",
  62659=>"010000011",
  62660=>"111111010",
  62661=>"000000000",
  62662=>"111000000",
  62663=>"011110000",
  62664=>"000001000",
  62665=>"000000000",
  62666=>"010011100",
  62667=>"000000001",
  62668=>"000010010",
  62669=>"001101010",
  62670=>"000001001",
  62671=>"000101000",
  62672=>"001111110",
  62673=>"100100011",
  62674=>"011101000",
  62675=>"010111111",
  62676=>"101000101",
  62677=>"011000111",
  62678=>"001111011",
  62679=>"000111111",
  62680=>"100000001",
  62681=>"111000000",
  62682=>"000000101",
  62683=>"000000111",
  62684=>"000001011",
  62685=>"000111110",
  62686=>"100000010",
  62687=>"011010001",
  62688=>"000000001",
  62689=>"111101101",
  62690=>"101111001",
  62691=>"101101111",
  62692=>"101000111",
  62693=>"000011011",
  62694=>"000101111",
  62695=>"011001111",
  62696=>"010010011",
  62697=>"110101111",
  62698=>"001000001",
  62699=>"000000001",
  62700=>"110111000",
  62701=>"100101001",
  62702=>"010000000",
  62703=>"000001000",
  62704=>"000000111",
  62705=>"000000100",
  62706=>"100000000",
  62707=>"011001001",
  62708=>"010110100",
  62709=>"001000000",
  62710=>"000000001",
  62711=>"110000000",
  62712=>"111111111",
  62713=>"000001011",
  62714=>"111001111",
  62715=>"001001010",
  62716=>"110000111",
  62717=>"100101111",
  62718=>"111110000",
  62719=>"001000100",
  62720=>"000001000",
  62721=>"000100000",
  62722=>"100010011",
  62723=>"101111111",
  62724=>"110111010",
  62725=>"000001011",
  62726=>"000011111",
  62727=>"000111110",
  62728=>"011011010",
  62729=>"011010100",
  62730=>"110110010",
  62731=>"100111111",
  62732=>"110100100",
  62733=>"010000001",
  62734=>"000000000",
  62735=>"100001000",
  62736=>"110111101",
  62737=>"111111001",
  62738=>"111100110",
  62739=>"100000110",
  62740=>"100000011",
  62741=>"011011101",
  62742=>"110100100",
  62743=>"110111111",
  62744=>"100000111",
  62745=>"100111101",
  62746=>"000000111",
  62747=>"011011011",
  62748=>"111011101",
  62749=>"000000100",
  62750=>"110111011",
  62751=>"000100001",
  62752=>"110100000",
  62753=>"000101111",
  62754=>"000001010",
  62755=>"011101000",
  62756=>"100110011",
  62757=>"111111111",
  62758=>"100010100",
  62759=>"111010000",
  62760=>"000001001",
  62761=>"111111011",
  62762=>"110110000",
  62763=>"100100100",
  62764=>"000100100",
  62765=>"101100000",
  62766=>"111110111",
  62767=>"000000110",
  62768=>"111110010",
  62769=>"110100100",
  62770=>"011111000",
  62771=>"000011001",
  62772=>"100100100",
  62773=>"110110000",
  62774=>"011000001",
  62775=>"000000001",
  62776=>"101111010",
  62777=>"000000011",
  62778=>"000000001",
  62779=>"111110110",
  62780=>"010000111",
  62781=>"000100001",
  62782=>"010000000",
  62783=>"100000000",
  62784=>"100111110",
  62785=>"110000000",
  62786=>"100100001",
  62787=>"000110100",
  62788=>"111000001",
  62789=>"100111011",
  62790=>"001001010",
  62791=>"100000000",
  62792=>"011011000",
  62793=>"011101111",
  62794=>"100000111",
  62795=>"111101111",
  62796=>"000001101",
  62797=>"010110111",
  62798=>"000100100",
  62799=>"111111101",
  62800=>"100000101",
  62801=>"100110111",
  62802=>"111011011",
  62803=>"101100100",
  62804=>"100110010",
  62805=>"110110111",
  62806=>"000100100",
  62807=>"101011011",
  62808=>"001001111",
  62809=>"000100100",
  62810=>"001001000",
  62811=>"000111100",
  62812=>"111111000",
  62813=>"001000000",
  62814=>"011111111",
  62815=>"100100001",
  62816=>"111000000",
  62817=>"111011000",
  62818=>"111011111",
  62819=>"111110101",
  62820=>"000100011",
  62821=>"001101000",
  62822=>"000000000",
  62823=>"000000100",
  62824=>"000001001",
  62825=>"000110010",
  62826=>"011111111",
  62827=>"001011111",
  62828=>"011110010",
  62829=>"011011011",
  62830=>"001100000",
  62831=>"011111011",
  62832=>"100100111",
  62833=>"100100010",
  62834=>"101110000",
  62835=>"001000000",
  62836=>"100111011",
  62837=>"001111111",
  62838=>"111011100",
  62839=>"111011011",
  62840=>"000010000",
  62841=>"001111011",
  62842=>"111000111",
  62843=>"011100110",
  62844=>"001100100",
  62845=>"111000011",
  62846=>"111011101",
  62847=>"100100000",
  62848=>"100011011",
  62849=>"011000100",
  62850=>"110011001",
  62851=>"011000000",
  62852=>"010000100",
  62853=>"010101000",
  62854=>"000000000",
  62855=>"010100000",
  62856=>"000100100",
  62857=>"110110010",
  62858=>"001001000",
  62859=>"001000011",
  62860=>"011011001",
  62861=>"110001010",
  62862=>"011001000",
  62863=>"000001100",
  62864=>"110110100",
  62865=>"111001100",
  62866=>"111000001",
  62867=>"100100100",
  62868=>"000101100",
  62869=>"100111011",
  62870=>"100100000",
  62871=>"000000000",
  62872=>"000001011",
  62873=>"011011010",
  62874=>"000101000",
  62875=>"001100000",
  62876=>"010010111",
  62877=>"110000111",
  62878=>"010010000",
  62879=>"111100100",
  62880=>"100100000",
  62881=>"111011001",
  62882=>"111100010",
  62883=>"110010101",
  62884=>"011011011",
  62885=>"001001000",
  62886=>"011111000",
  62887=>"111100000",
  62888=>"111111011",
  62889=>"000111111",
  62890=>"111000000",
  62891=>"111100110",
  62892=>"001111110",
  62893=>"100000111",
  62894=>"001000010",
  62895=>"111001100",
  62896=>"011100101",
  62897=>"001001000",
  62898=>"111100011",
  62899=>"011100110",
  62900=>"101101000",
  62901=>"011001000",
  62902=>"111011110",
  62903=>"000000100",
  62904=>"001011000",
  62905=>"101111011",
  62906=>"111001011",
  62907=>"110110000",
  62908=>"001101011",
  62909=>"110111111",
  62910=>"010000001",
  62911=>"001000101",
  62912=>"111011001",
  62913=>"110100000",
  62914=>"111101010",
  62915=>"100100101",
  62916=>"000000000",
  62917=>"000101111",
  62918=>"100111011",
  62919=>"111000000",
  62920=>"101000100",
  62921=>"000011011",
  62922=>"100010011",
  62923=>"010111010",
  62924=>"000111000",
  62925=>"000000001",
  62926=>"000011001",
  62927=>"110010000",
  62928=>"100001000",
  62929=>"000111110",
  62930=>"011000001",
  62931=>"110100000",
  62932=>"110111001",
  62933=>"110111111",
  62934=>"000100000",
  62935=>"000100010",
  62936=>"110100100",
  62937=>"111100000",
  62938=>"010100110",
  62939=>"011011001",
  62940=>"000100110",
  62941=>"111001010",
  62942=>"001110000",
  62943=>"111111011",
  62944=>"000111000",
  62945=>"010010000",
  62946=>"011001000",
  62947=>"100111110",
  62948=>"101001000",
  62949=>"100001111",
  62950=>"100110010",
  62951=>"001111110",
  62952=>"011101101",
  62953=>"111000000",
  62954=>"111001000",
  62955=>"111111101",
  62956=>"000011000",
  62957=>"000100011",
  62958=>"000011011",
  62959=>"111000000",
  62960=>"000111001",
  62961=>"000100110",
  62962=>"110000011",
  62963=>"110000001",
  62964=>"000110100",
  62965=>"001000000",
  62966=>"001011110",
  62967=>"010001100",
  62968=>"000111111",
  62969=>"001001001",
  62970=>"111111100",
  62971=>"000100101",
  62972=>"000101101",
  62973=>"010111110",
  62974=>"000111000",
  62975=>"000010111",
  62976=>"001001000",
  62977=>"010100011",
  62978=>"001001111",
  62979=>"001001111",
  62980=>"000000110",
  62981=>"111001001",
  62982=>"001001001",
  62983=>"010000000",
  62984=>"001001111",
  62985=>"000000110",
  62986=>"100101101",
  62987=>"111011011",
  62988=>"001001011",
  62989=>"011111110",
  62990=>"011001011",
  62991=>"010111111",
  62992=>"011011110",
  62993=>"011001011",
  62994=>"001000111",
  62995=>"110100000",
  62996=>"011001110",
  62997=>"110110100",
  62998=>"101111011",
  62999=>"001110101",
  63000=>"011001111",
  63001=>"100100100",
  63002=>"110011111",
  63003=>"011001111",
  63004=>"100100110",
  63005=>"100010110",
  63006=>"111111111",
  63007=>"100011000",
  63008=>"100111101",
  63009=>"001011111",
  63010=>"000110000",
  63011=>"110000000",
  63012=>"000100000",
  63013=>"111011000",
  63014=>"000000110",
  63015=>"001101111",
  63016=>"110110110",
  63017=>"111011111",
  63018=>"001100000",
  63019=>"000000000",
  63020=>"010000100",
  63021=>"111010011",
  63022=>"110110110",
  63023=>"111001110",
  63024=>"110111000",
  63025=>"000000000",
  63026=>"000110111",
  63027=>"100000100",
  63028=>"100110110",
  63029=>"010000001",
  63030=>"111001000",
  63031=>"100100110",
  63032=>"101000000",
  63033=>"001001111",
  63034=>"000000101",
  63035=>"000100000",
  63036=>"100110000",
  63037=>"001100001",
  63038=>"000000011",
  63039=>"000000001",
  63040=>"111011001",
  63041=>"111111000",
  63042=>"011001001",
  63043=>"011011001",
  63044=>"011011000",
  63045=>"001001011",
  63046=>"100110000",
  63047=>"101000101",
  63048=>"111011100",
  63049=>"010000100",
  63050=>"011011011",
  63051=>"100100000",
  63052=>"100001000",
  63053=>"100010110",
  63054=>"000001001",
  63055=>"000000100",
  63056=>"011000111",
  63057=>"100111110",
  63058=>"101011111",
  63059=>"100111100",
  63060=>"011000010",
  63061=>"111110111",
  63062=>"110110100",
  63063=>"001001011",
  63064=>"010000000",
  63065=>"110100100",
  63066=>"110111100",
  63067=>"100110000",
  63068=>"110110100",
  63069=>"100100100",
  63070=>"111111011",
  63071=>"001010011",
  63072=>"000100001",
  63073=>"001001111",
  63074=>"001001011",
  63075=>"100100100",
  63076=>"011011001",
  63077=>"000110110",
  63078=>"111110100",
  63079=>"111110110",
  63080=>"101101001",
  63081=>"100001001",
  63082=>"000111111",
  63083=>"001111111",
  63084=>"110010110",
  63085=>"010011001",
  63086=>"110110000",
  63087=>"111101001",
  63088=>"000100000",
  63089=>"111100100",
  63090=>"001000000",
  63091=>"001001000",
  63092=>"001001000",
  63093=>"000001100",
  63094=>"100001110",
  63095=>"110110111",
  63096=>"110111111",
  63097=>"010100000",
  63098=>"001100100",
  63099=>"001001001",
  63100=>"100100101",
  63101=>"111001000",
  63102=>"101111110",
  63103=>"011001111",
  63104=>"110111000",
  63105=>"000000001",
  63106=>"100100100",
  63107=>"100100111",
  63108=>"111011111",
  63109=>"101111000",
  63110=>"100100000",
  63111=>"000001000",
  63112=>"110010000",
  63113=>"111000010",
  63114=>"111111000",
  63115=>"011000110",
  63116=>"001111001",
  63117=>"001000001",
  63118=>"001001110",
  63119=>"100000100",
  63120=>"111100101",
  63121=>"110011001",
  63122=>"100111000",
  63123=>"011001001",
  63124=>"100000110",
  63125=>"001001111",
  63126=>"000100100",
  63127=>"001001000",
  63128=>"101101010",
  63129=>"000001110",
  63130=>"100110100",
  63131=>"100001000",
  63132=>"111000000",
  63133=>"111100000",
  63134=>"011100000",
  63135=>"010011111",
  63136=>"100001011",
  63137=>"111010001",
  63138=>"001001110",
  63139=>"111111011",
  63140=>"001011000",
  63141=>"110000100",
  63142=>"001000111",
  63143=>"000100100",
  63144=>"110000100",
  63145=>"011001010",
  63146=>"110010110",
  63147=>"011001111",
  63148=>"110111001",
  63149=>"001001111",
  63150=>"010011110",
  63151=>"001000111",
  63152=>"001111010",
  63153=>"001001010",
  63154=>"111001111",
  63155=>"111001001",
  63156=>"111111100",
  63157=>"110110000",
  63158=>"111110110",
  63159=>"000111000",
  63160=>"110100111",
  63161=>"001100000",
  63162=>"110010000",
  63163=>"111111000",
  63164=>"100010010",
  63165=>"101001000",
  63166=>"011011111",
  63167=>"101000000",
  63168=>"111100111",
  63169=>"110110100",
  63170=>"100101101",
  63171=>"001110100",
  63172=>"000110000",
  63173=>"110011001",
  63174=>"111001001",
  63175=>"000110110",
  63176=>"110100111",
  63177=>"100001001",
  63178=>"110110110",
  63179=>"000100100",
  63180=>"110100000",
  63181=>"001100101",
  63182=>"100110100",
  63183=>"100100111",
  63184=>"001011011",
  63185=>"001110010",
  63186=>"101000001",
  63187=>"011110101",
  63188=>"111100110",
  63189=>"100111100",
  63190=>"011001011",
  63191=>"110110110",
  63192=>"100110000",
  63193=>"011011010",
  63194=>"000000001",
  63195=>"110001011",
  63196=>"000101001",
  63197=>"111011010",
  63198=>"110110000",
  63199=>"111111000",
  63200=>"011001011",
  63201=>"011001011",
  63202=>"111011001",
  63203=>"001001101",
  63204=>"111001001",
  63205=>"011001011",
  63206=>"001001001",
  63207=>"100110000",
  63208=>"111011011",
  63209=>"010110100",
  63210=>"111111100",
  63211=>"001000000",
  63212=>"011001001",
  63213=>"110111111",
  63214=>"110100110",
  63215=>"110110010",
  63216=>"100000000",
  63217=>"001000011",
  63218=>"010001110",
  63219=>"100100110",
  63220=>"100111111",
  63221=>"000111110",
  63222=>"000100100",
  63223=>"100000100",
  63224=>"001110100",
  63225=>"000111100",
  63226=>"110001011",
  63227=>"001011100",
  63228=>"110110100",
  63229=>"010000000",
  63230=>"100111101",
  63231=>"111101101",
  63232=>"000000110",
  63233=>"101000000",
  63234=>"001000000",
  63235=>"000111010",
  63236=>"000000000",
  63237=>"110000111",
  63238=>"000011010",
  63239=>"000000000",
  63240=>"110010111",
  63241=>"000000001",
  63242=>"001011110",
  63243=>"000000000",
  63244=>"000111110",
  63245=>"101000110",
  63246=>"000010010",
  63247=>"011111001",
  63248=>"000000101",
  63249=>"111010011",
  63250=>"111111011",
  63251=>"000100111",
  63252=>"000000000",
  63253=>"000000000",
  63254=>"111111100",
  63255=>"110110010",
  63256=>"011000010",
  63257=>"100111111",
  63258=>"011000111",
  63259=>"000000000",
  63260=>"000000101",
  63261=>"001101001",
  63262=>"000000000",
  63263=>"111111111",
  63264=>"111000111",
  63265=>"000101000",
  63266=>"001100000",
  63267=>"101001111",
  63268=>"000100110",
  63269=>"001000111",
  63270=>"000010010",
  63271=>"111001010",
  63272=>"000000001",
  63273=>"111001001",
  63274=>"010111110",
  63275=>"111111111",
  63276=>"010101011",
  63277=>"101010000",
  63278=>"111111010",
  63279=>"000001001",
  63280=>"110111111",
  63281=>"110110110",
  63282=>"000101101",
  63283=>"010000010",
  63284=>"101000000",
  63285=>"001010011",
  63286=>"001110010",
  63287=>"000000000",
  63288=>"010111001",
  63289=>"000000000",
  63290=>"100111000",
  63291=>"010010000",
  63292=>"011000010",
  63293=>"111111101",
  63294=>"101001101",
  63295=>"100111001",
  63296=>"111010111",
  63297=>"000000001",
  63298=>"000111000",
  63299=>"001000100",
  63300=>"110110000",
  63301=>"111110010",
  63302=>"000000000",
  63303=>"000000111",
  63304=>"110010101",
  63305=>"010000000",
  63306=>"100001011",
  63307=>"111110110",
  63308=>"100101101",
  63309=>"011011011",
  63310=>"000001011",
  63311=>"111111111",
  63312=>"000000000",
  63313=>"111110110",
  63314=>"101000010",
  63315=>"101110000",
  63316=>"000000001",
  63317=>"110000000",
  63318=>"000001001",
  63319=>"000000000",
  63320=>"111111011",
  63321=>"101111111",
  63322=>"000010100",
  63323=>"011111100",
  63324=>"111111010",
  63325=>"000100100",
  63326=>"111000000",
  63327=>"000000001",
  63328=>"010000001",
  63329=>"110110000",
  63330=>"000000100",
  63331=>"000001001",
  63332=>"000111110",
  63333=>"111001111",
  63334=>"110010000",
  63335=>"000000000",
  63336=>"000011000",
  63337=>"000010010",
  63338=>"111000000",
  63339=>"101000110",
  63340=>"100100000",
  63341=>"010010011",
  63342=>"000000000",
  63343=>"000000000",
  63344=>"101111111",
  63345=>"111111000",
  63346=>"011110011",
  63347=>"000101000",
  63348=>"000000000",
  63349=>"000110000",
  63350=>"000111000",
  63351=>"111010111",
  63352=>"011111101",
  63353=>"111111000",
  63354=>"111100100",
  63355=>"111111011",
  63356=>"100010100",
  63357=>"000110111",
  63358=>"000000010",
  63359=>"111000000",
  63360=>"110111001",
  63361=>"111100000",
  63362=>"011011010",
  63363=>"011110110",
  63364=>"001101001",
  63365=>"000111111",
  63366=>"010010110",
  63367=>"100110011",
  63368=>"111111101",
  63369=>"101101000",
  63370=>"001111001",
  63371=>"001000000",
  63372=>"000000000",
  63373=>"011111101",
  63374=>"110110110",
  63375=>"001001000",
  63376=>"111111111",
  63377=>"100011111",
  63378=>"111001101",
  63379=>"101000110",
  63380=>"000110010",
  63381=>"111101100",
  63382=>"100010000",
  63383=>"110110010",
  63384=>"100101101",
  63385=>"110110111",
  63386=>"000110110",
  63387=>"000000111",
  63388=>"111000110",
  63389=>"010111000",
  63390=>"111000000",
  63391=>"000000000",
  63392=>"001011011",
  63393=>"111111011",
  63394=>"000000111",
  63395=>"101011111",
  63396=>"000110110",
  63397=>"110111010",
  63398=>"111001000",
  63399=>"000000001",
  63400=>"011010010",
  63401=>"000000000",
  63402=>"111111111",
  63403=>"001101000",
  63404=>"111111110",
  63405=>"101101111",
  63406=>"000101011",
  63407=>"001111110",
  63408=>"000000010",
  63409=>"001110110",
  63410=>"111111010",
  63411=>"000001011",
  63412=>"111111111",
  63413=>"010011001",
  63414=>"101011111",
  63415=>"101000110",
  63416=>"010010000",
  63417=>"001011011",
  63418=>"101000010",
  63419=>"110111111",
  63420=>"000100000",
  63421=>"000000111",
  63422=>"110110101",
  63423=>"010000101",
  63424=>"111111010",
  63425=>"011011010",
  63426=>"111111000",
  63427=>"110110100",
  63428=>"000001111",
  63429=>"110110001",
  63430=>"000000100",
  63431=>"000000111",
  63432=>"000000111",
  63433=>"101111111",
  63434=>"101000111",
  63435=>"010110000",
  63436=>"111010010",
  63437=>"000000010",
  63438=>"001101110",
  63439=>"111011000",
  63440=>"001000000",
  63441=>"101111110",
  63442=>"000001100",
  63443=>"111101101",
  63444=>"001111111",
  63445=>"001100001",
  63446=>"000000000",
  63447=>"110000111",
  63448=>"000000000",
  63449=>"000001101",
  63450=>"100110111",
  63451=>"000111111",
  63452=>"111001111",
  63453=>"111111111",
  63454=>"000000000",
  63455=>"000000101",
  63456=>"111111001",
  63457=>"111000000",
  63458=>"111010000",
  63459=>"001011011",
  63460=>"000000000",
  63461=>"000000010",
  63462=>"000000010",
  63463=>"010111100",
  63464=>"111000111",
  63465=>"000100100",
  63466=>"110010000",
  63467=>"010000111",
  63468=>"000001101",
  63469=>"000000001",
  63470=>"000111010",
  63471=>"000000010",
  63472=>"101101111",
  63473=>"011010110",
  63474=>"101111000",
  63475=>"010111011",
  63476=>"000001011",
  63477=>"000101001",
  63478=>"000100110",
  63479=>"000001000",
  63480=>"000110100",
  63481=>"000000000",
  63482=>"111111110",
  63483=>"111111001",
  63484=>"000010010",
  63485=>"000000010",
  63486=>"100111011",
  63487=>"000111111",
  63488=>"111110111",
  63489=>"010010000",
  63490=>"100000000",
  63491=>"000010111",
  63492=>"011111011",
  63493=>"111111010",
  63494=>"011110100",
  63495=>"010000000",
  63496=>"000111010",
  63497=>"100111000",
  63498=>"101111011",
  63499=>"000000100",
  63500=>"100000101",
  63501=>"111111111",
  63502=>"111101000",
  63503=>"101001010",
  63504=>"001001100",
  63505=>"110000110",
  63506=>"001000000",
  63507=>"011100000",
  63508=>"000100100",
  63509=>"000010000",
  63510=>"010110011",
  63511=>"110110001",
  63512=>"000001111",
  63513=>"000000100",
  63514=>"011011000",
  63515=>"000111100",
  63516=>"101100010",
  63517=>"000000111",
  63518=>"111010001",
  63519=>"000000010",
  63520=>"111111111",
  63521=>"111111111",
  63522=>"101000110",
  63523=>"011111111",
  63524=>"001011010",
  63525=>"101001010",
  63526=>"110110000",
  63527=>"000000000",
  63528=>"011111010",
  63529=>"000010000",
  63530=>"101111000",
  63531=>"010010000",
  63532=>"000011011",
  63533=>"101111001",
  63534=>"111111011",
  63535=>"011000010",
  63536=>"000000110",
  63537=>"001011011",
  63538=>"111011110",
  63539=>"111111111",
  63540=>"101110111",
  63541=>"100000000",
  63542=>"100000000",
  63543=>"000000000",
  63544=>"111010000",
  63545=>"100000100",
  63546=>"111111111",
  63547=>"010111110",
  63548=>"100000001",
  63549=>"111111111",
  63550=>"000000001",
  63551=>"001111110",
  63552=>"111000101",
  63553=>"000110111",
  63554=>"111111000",
  63555=>"110111011",
  63556=>"100111111",
  63557=>"001100110",
  63558=>"011000011",
  63559=>"111101011",
  63560=>"110001000",
  63561=>"000000000",
  63562=>"100000101",
  63563=>"000000100",
  63564=>"011111110",
  63565=>"101110011",
  63566=>"100111111",
  63567=>"010000010",
  63568=>"010000000",
  63569=>"111111111",
  63570=>"000000011",
  63571=>"001001001",
  63572=>"111000001",
  63573=>"111111111",
  63574=>"011011011",
  63575=>"011000100",
  63576=>"111111101",
  63577=>"101111111",
  63578=>"000001001",
  63579=>"110110010",
  63580=>"111111100",
  63581=>"000011000",
  63582=>"000000000",
  63583=>"001101111",
  63584=>"000011010",
  63585=>"110100010",
  63586=>"100100100",
  63587=>"000110111",
  63588=>"100110000",
  63589=>"110110111",
  63590=>"011110000",
  63591=>"111111000",
  63592=>"111111111",
  63593=>"111111000",
  63594=>"110010111",
  63595=>"101111000",
  63596=>"000000111",
  63597=>"011111000",
  63598=>"100000000",
  63599=>"011001111",
  63600=>"100110111",
  63601=>"000010111",
  63602=>"101000100",
  63603=>"000000001",
  63604=>"000111000",
  63605=>"000000000",
  63606=>"001110110",
  63607=>"110000000",
  63608=>"100101111",
  63609=>"111100000",
  63610=>"000001000",
  63611=>"000111011",
  63612=>"011011001",
  63613=>"010110100",
  63614=>"110111010",
  63615=>"000100000",
  63616=>"000111011",
  63617=>"111101100",
  63618=>"010010110",
  63619=>"011010011",
  63620=>"000111000",
  63621=>"000000000",
  63622=>"001101111",
  63623=>"011000100",
  63624=>"001001011",
  63625=>"000000111",
  63626=>"111000000",
  63627=>"101000110",
  63628=>"000111000",
  63629=>"110011000",
  63630=>"100000000",
  63631=>"001000001",
  63632=>"001001100",
  63633=>"011011111",
  63634=>"111111011",
  63635=>"011000001",
  63636=>"011000000",
  63637=>"101111110",
  63638=>"001000000",
  63639=>"000001011",
  63640=>"011101110",
  63641=>"101000101",
  63642=>"111111110",
  63643=>"010100000",
  63644=>"000011111",
  63645=>"111111110",
  63646=>"010100111",
  63647=>"000000100",
  63648=>"010001111",
  63649=>"000000111",
  63650=>"000000000",
  63651=>"111001000",
  63652=>"011110010",
  63653=>"000000010",
  63654=>"001000001",
  63655=>"100011010",
  63656=>"111111000",
  63657=>"000011010",
  63658=>"111110111",
  63659=>"000111111",
  63660=>"011001111",
  63661=>"111111111",
  63662=>"111011010",
  63663=>"000001000",
  63664=>"000000010",
  63665=>"010000000",
  63666=>"000100100",
  63667=>"011111011",
  63668=>"100110000",
  63669=>"000100110",
  63670=>"011001010",
  63671=>"000000100",
  63672=>"001001110",
  63673=>"111001000",
  63674=>"000000010",
  63675=>"100111111",
  63676=>"011010000",
  63677=>"101101101",
  63678=>"010111111",
  63679=>"111010001",
  63680=>"100000000",
  63681=>"000000101",
  63682=>"010010010",
  63683=>"111010101",
  63684=>"111000100",
  63685=>"010011111",
  63686=>"010010111",
  63687=>"101110111",
  63688=>"110001100",
  63689=>"111110100",
  63690=>"010101111",
  63691=>"101000100",
  63692=>"000011111",
  63693=>"010110100",
  63694=>"000000100",
  63695=>"000111111",
  63696=>"000111111",
  63697=>"000110110",
  63698=>"000000100",
  63699=>"000111111",
  63700=>"000000000",
  63701=>"010000001",
  63702=>"010011000",
  63703=>"101011111",
  63704=>"000000100",
  63705=>"101001010",
  63706=>"000010111",
  63707=>"000000000",
  63708=>"100111110",
  63709=>"111111111",
  63710=>"001000001",
  63711=>"011110000",
  63712=>"111111010",
  63713=>"000000000",
  63714=>"000000000",
  63715=>"101111100",
  63716=>"000000100",
  63717=>"111110000",
  63718=>"000100111",
  63719=>"111101010",
  63720=>"000111111",
  63721=>"000000100",
  63722=>"111011011",
  63723=>"101111110",
  63724=>"100000000",
  63725=>"110000111",
  63726=>"010111010",
  63727=>"010011001",
  63728=>"000100000",
  63729=>"010111101",
  63730=>"000000010",
  63731=>"000111110",
  63732=>"101001111",
  63733=>"010101010",
  63734=>"001000000",
  63735=>"001111010",
  63736=>"000000100",
  63737=>"010111111",
  63738=>"000000000",
  63739=>"001010010",
  63740=>"101000000",
  63741=>"111000010",
  63742=>"110110110",
  63743=>"111100001",
  63744=>"011010010",
  63745=>"010010010",
  63746=>"000011110",
  63747=>"111110010",
  63748=>"001011001",
  63749=>"010000010",
  63750=>"111111111",
  63751=>"111111100",
  63752=>"000000000",
  63753=>"001001101",
  63754=>"110110010",
  63755=>"101001101",
  63756=>"101000000",
  63757=>"111111000",
  63758=>"111111011",
  63759=>"001001101",
  63760=>"000101110",
  63761=>"010111000",
  63762=>"001001001",
  63763=>"000111111",
  63764=>"010010010",
  63765=>"001101100",
  63766=>"000001000",
  63767=>"010110111",
  63768=>"000000000",
  63769=>"111111111",
  63770=>"100100111",
  63771=>"111000000",
  63772=>"000001111",
  63773=>"101000111",
  63774=>"010010111",
  63775=>"001001001",
  63776=>"000011011",
  63777=>"000000001",
  63778=>"001000000",
  63779=>"000000000",
  63780=>"011001011",
  63781=>"110111100",
  63782=>"000000000",
  63783=>"000000000",
  63784=>"000001101",
  63785=>"000001000",
  63786=>"110110010",
  63787=>"111111101",
  63788=>"011111111",
  63789=>"101110110",
  63790=>"111110100",
  63791=>"000100000",
  63792=>"010011110",
  63793=>"101101101",
  63794=>"000000001",
  63795=>"110110111",
  63796=>"111111111",
  63797=>"111111110",
  63798=>"001111010",
  63799=>"110111010",
  63800=>"010000010",
  63801=>"111110010",
  63802=>"000000001",
  63803=>"000000100",
  63804=>"000000000",
  63805=>"111111111",
  63806=>"111101010",
  63807=>"100110010",
  63808=>"010000100",
  63809=>"111100110",
  63810=>"101000000",
  63811=>"011001101",
  63812=>"000000000",
  63813=>"010000101",
  63814=>"110110110",
  63815=>"001001011",
  63816=>"101011000",
  63817=>"001001111",
  63818=>"111111000",
  63819=>"010111111",
  63820=>"001001010",
  63821=>"111111111",
  63822=>"100111111",
  63823=>"110100000",
  63824=>"111000100",
  63825=>"110111010",
  63826=>"000010010",
  63827=>"001001011",
  63828=>"001000000",
  63829=>"100111001",
  63830=>"100100100",
  63831=>"000000111",
  63832=>"000000111",
  63833=>"110100000",
  63834=>"111100100",
  63835=>"110110110",
  63836=>"000001111",
  63837=>"001011011",
  63838=>"110111111",
  63839=>"100000111",
  63840=>"111001101",
  63841=>"000000000",
  63842=>"001000001",
  63843=>"001011111",
  63844=>"100110100",
  63845=>"000001001",
  63846=>"100110111",
  63847=>"111101101",
  63848=>"000010001",
  63849=>"000011111",
  63850=>"111000100",
  63851=>"001101010",
  63852=>"000000101",
  63853=>"110111010",
  63854=>"010010000",
  63855=>"100011111",
  63856=>"001011001",
  63857=>"110110000",
  63858=>"110110011",
  63859=>"001110110",
  63860=>"111001000",
  63861=>"000001000",
  63862=>"000001000",
  63863=>"100000100",
  63864=>"010000000",
  63865=>"110000000",
  63866=>"011001010",
  63867=>"001010111",
  63868=>"100110110",
  63869=>"100000100",
  63870=>"111111100",
  63871=>"000001111",
  63872=>"000000000",
  63873=>"111001111",
  63874=>"010010000",
  63875=>"001000101",
  63876=>"000101111",
  63877=>"101000000",
  63878=>"110101011",
  63879=>"111111010",
  63880=>"101111111",
  63881=>"100110000",
  63882=>"100100000",
  63883=>"000011101",
  63884=>"011101101",
  63885=>"000000101",
  63886=>"111111110",
  63887=>"100001000",
  63888=>"101101100",
  63889=>"111001001",
  63890=>"110111111",
  63891=>"011000000",
  63892=>"000111101",
  63893=>"000000000",
  63894=>"001000000",
  63895=>"100000000",
  63896=>"000000000",
  63897=>"111101100",
  63898=>"101000001",
  63899=>"000000100",
  63900=>"000011110",
  63901=>"111111001",
  63902=>"111111000",
  63903=>"111001001",
  63904=>"111001000",
  63905=>"000000001",
  63906=>"110011110",
  63907=>"101111110",
  63908=>"000000111",
  63909=>"110010110",
  63910=>"000010111",
  63911=>"000110011",
  63912=>"010110110",
  63913=>"000000000",
  63914=>"111000000",
  63915=>"000110000",
  63916=>"011011111",
  63917=>"001000101",
  63918=>"100011000",
  63919=>"110111101",
  63920=>"011111101",
  63921=>"101110100",
  63922=>"101000101",
  63923=>"000000000",
  63924=>"111111111",
  63925=>"010010101",
  63926=>"100000110",
  63927=>"000010000",
  63928=>"001000100",
  63929=>"110111111",
  63930=>"110100111",
  63931=>"010110001",
  63932=>"000010100",
  63933=>"000000000",
  63934=>"000000001",
  63935=>"111000110",
  63936=>"010110010",
  63937=>"111111010",
  63938=>"010000000",
  63939=>"111011011",
  63940=>"111000000",
  63941=>"100100100",
  63942=>"010000010",
  63943=>"110111111",
  63944=>"111001100",
  63945=>"111100110",
  63946=>"111110000",
  63947=>"111111111",
  63948=>"010000000",
  63949=>"011001110",
  63950=>"111000010",
  63951=>"111101000",
  63952=>"000000000",
  63953=>"111011111",
  63954=>"111001011",
  63955=>"001001000",
  63956=>"101111111",
  63957=>"110110000",
  63958=>"100110010",
  63959=>"111000000",
  63960=>"110010010",
  63961=>"000010111",
  63962=>"100000000",
  63963=>"000111111",
  63964=>"111000100",
  63965=>"000001111",
  63966=>"000100011",
  63967=>"111011010",
  63968=>"000101001",
  63969=>"111111111",
  63970=>"111111101",
  63971=>"110111110",
  63972=>"100100110",
  63973=>"010110001",
  63974=>"010000000",
  63975=>"111010000",
  63976=>"001000000",
  63977=>"010000010",
  63978=>"010111010",
  63979=>"001010000",
  63980=>"000000000",
  63981=>"001001111",
  63982=>"001011000",
  63983=>"101011000",
  63984=>"000000000",
  63985=>"011011001",
  63986=>"111000111",
  63987=>"010000000",
  63988=>"110110000",
  63989=>"000111110",
  63990=>"000000110",
  63991=>"000001001",
  63992=>"000000000",
  63993=>"110111101",
  63994=>"111101111",
  63995=>"110111111",
  63996=>"000000111",
  63997=>"000100000",
  63998=>"100100001",
  63999=>"110111010",
  64000=>"001001111",
  64001=>"000111111",
  64002=>"110000000",
  64003=>"111111111",
  64004=>"000010011",
  64005=>"000000001",
  64006=>"111000000",
  64007=>"000011001",
  64008=>"000000000",
  64009=>"111100001",
  64010=>"110000000",
  64011=>"111001010",
  64012=>"000000101",
  64013=>"001101111",
  64014=>"010011011",
  64015=>"111111111",
  64016=>"000000000",
  64017=>"001010010",
  64018=>"010000000",
  64019=>"000010011",
  64020=>"101011111",
  64021=>"111111011",
  64022=>"011111111",
  64023=>"111011111",
  64024=>"111000000",
  64025=>"101111011",
  64026=>"000010110",
  64027=>"011110111",
  64028=>"010000101",
  64029=>"110100000",
  64030=>"111110111",
  64031=>"111111111",
  64032=>"100101000",
  64033=>"111000011",
  64034=>"100111011",
  64035=>"111111101",
  64036=>"011001011",
  64037=>"111110111",
  64038=>"100000010",
  64039=>"001000000",
  64040=>"111000000",
  64041=>"111111011",
  64042=>"000000000",
  64043=>"000101101",
  64044=>"001111111",
  64045=>"111000000",
  64046=>"111111101",
  64047=>"111111000",
  64048=>"111011000",
  64049=>"001001001",
  64050=>"100101111",
  64051=>"101110000",
  64052=>"111011000",
  64053=>"110111111",
  64054=>"000111111",
  64055=>"000110111",
  64056=>"111010110",
  64057=>"000000111",
  64058=>"001100000",
  64059=>"101101111",
  64060=>"011111011",
  64061=>"111010111",
  64062=>"000000111",
  64063=>"000000000",
  64064=>"111101000",
  64065=>"111010011",
  64066=>"111111101",
  64067=>"001010000",
  64068=>"111101111",
  64069=>"000100000",
  64070=>"000000000",
  64071=>"111010010",
  64072=>"100100111",
  64073=>"000000000",
  64074=>"000100101",
  64075=>"101001111",
  64076=>"100000000",
  64077=>"000000000",
  64078=>"000100110",
  64079=>"000011000",
  64080=>"000101011",
  64081=>"111010000",
  64082=>"011000000",
  64083=>"111011001",
  64084=>"000100111",
  64085=>"111111100",
  64086=>"011001001",
  64087=>"101001000",
  64088=>"101110000",
  64089=>"001111111",
  64090=>"000001001",
  64091=>"101111111",
  64092=>"110111111",
  64093=>"110001001",
  64094=>"101000000",
  64095=>"000001100",
  64096=>"000000111",
  64097=>"000000000",
  64098=>"100101111",
  64099=>"000110110",
  64100=>"001111111",
  64101=>"100110100",
  64102=>"000000000",
  64103=>"111111110",
  64104=>"000000000",
  64105=>"111000000",
  64106=>"011000000",
  64107=>"111011111",
  64108=>"000010000",
  64109=>"111100000",
  64110=>"011000111",
  64111=>"000001000",
  64112=>"000001110",
  64113=>"111010101",
  64114=>"000111011",
  64115=>"111011000",
  64116=>"111111111",
  64117=>"101101101",
  64118=>"111111111",
  64119=>"101111111",
  64120=>"000010000",
  64121=>"111111111",
  64122=>"000000001",
  64123=>"011000000",
  64124=>"000111110",
  64125=>"111100100",
  64126=>"100000000",
  64127=>"111101100",
  64128=>"111111111",
  64129=>"111011000",
  64130=>"011011011",
  64131=>"010111001",
  64132=>"000000000",
  64133=>"001111111",
  64134=>"111011010",
  64135=>"000100111",
  64136=>"000111011",
  64137=>"000000000",
  64138=>"000000000",
  64139=>"111100000",
  64140=>"000000000",
  64141=>"011010010",
  64142=>"111011111",
  64143=>"000000000",
  64144=>"011011111",
  64145=>"000010111",
  64146=>"101001111",
  64147=>"110111000",
  64148=>"000100101",
  64149=>"111000000",
  64150=>"001011011",
  64151=>"000111111",
  64152=>"001001000",
  64153=>"111011000",
  64154=>"111010000",
  64155=>"000000111",
  64156=>"100100100",
  64157=>"000011011",
  64158=>"111111110",
  64159=>"111111111",
  64160=>"000000010",
  64161=>"101000000",
  64162=>"111111111",
  64163=>"111010001",
  64164=>"111010000",
  64165=>"000111111",
  64166=>"111111111",
  64167=>"000111111",
  64168=>"111011000",
  64169=>"011010111",
  64170=>"000000000",
  64171=>"101000000",
  64172=>"111011001",
  64173=>"110000000",
  64174=>"001010110",
  64175=>"000111011",
  64176=>"000000010",
  64177=>"000001111",
  64178=>"111101100",
  64179=>"000000000",
  64180=>"000110110",
  64181=>"101111011",
  64182=>"000101111",
  64183=>"101111000",
  64184=>"110111111",
  64185=>"000101101",
  64186=>"101001010",
  64187=>"010010111",
  64188=>"001000010",
  64189=>"111100000",
  64190=>"010000110",
  64191=>"101111111",
  64192=>"111000100",
  64193=>"000111111",
  64194=>"011010111",
  64195=>"110111111",
  64196=>"101001000",
  64197=>"001000000",
  64198=>"010100000",
  64199=>"101001101",
  64200=>"010000000",
  64201=>"000111111",
  64202=>"110001111",
  64203=>"000000111",
  64204=>"000000000",
  64205=>"110111111",
  64206=>"000111111",
  64207=>"111000100",
  64208=>"111000000",
  64209=>"000110111",
  64210=>"001101001",
  64211=>"111000110",
  64212=>"111101110",
  64213=>"001000110",
  64214=>"111000111",
  64215=>"101110000",
  64216=>"111111111",
  64217=>"000000111",
  64218=>"100100100",
  64219=>"111000000",
  64220=>"111110101",
  64221=>"111000000",
  64222=>"101111111",
  64223=>"100000010",
  64224=>"101000101",
  64225=>"111000100",
  64226=>"111000000",
  64227=>"000011111",
  64228=>"000000010",
  64229=>"010111111",
  64230=>"000111111",
  64231=>"000000000",
  64232=>"000000000",
  64233=>"000000000",
  64234=>"001000000",
  64235=>"000011011",
  64236=>"000100101",
  64237=>"001111101",
  64238=>"111000000",
  64239=>"111111111",
  64240=>"111111101",
  64241=>"011000000",
  64242=>"111111111",
  64243=>"000111111",
  64244=>"011110111",
  64245=>"000000000",
  64246=>"111101011",
  64247=>"101000100",
  64248=>"101101111",
  64249=>"101000000",
  64250=>"111111000",
  64251=>"000101111",
  64252=>"101000101",
  64253=>"000000000",
  64254=>"101100110",
  64255=>"000111011",
  64256=>"100100110",
  64257=>"010110000",
  64258=>"100000001",
  64259=>"010010000",
  64260=>"011001000",
  64261=>"000001110",
  64262=>"100000000",
  64263=>"111010100",
  64264=>"011101001",
  64265=>"100000000",
  64266=>"111111010",
  64267=>"111101001",
  64268=>"000010010",
  64269=>"011000101",
  64270=>"100100100",
  64271=>"000000000",
  64272=>"100000000",
  64273=>"111000001",
  64274=>"010111111",
  64275=>"100000000",
  64276=>"110111111",
  64277=>"010111111",
  64278=>"001111010",
  64279=>"110100000",
  64280=>"001000000",
  64281=>"111011000",
  64282=>"000000110",
  64283=>"111000100",
  64284=>"100000000",
  64285=>"000101101",
  64286=>"000001111",
  64287=>"100000100",
  64288=>"011011000",
  64289=>"111111110",
  64290=>"100000000",
  64291=>"011010000",
  64292=>"011001011",
  64293=>"000001011",
  64294=>"111111111",
  64295=>"010000111",
  64296=>"010011000",
  64297=>"000000000",
  64298=>"000100110",
  64299=>"000000000",
  64300=>"111011011",
  64301=>"001010100",
  64302=>"000111111",
  64303=>"011011011",
  64304=>"011111111",
  64305=>"111111111",
  64306=>"001111010",
  64307=>"000010000",
  64308=>"000010111",
  64309=>"111111111",
  64310=>"100101011",
  64311=>"100000000",
  64312=>"101000111",
  64313=>"000000001",
  64314=>"010011010",
  64315=>"100000000",
  64316=>"010111001",
  64317=>"111111111",
  64318=>"000000000",
  64319=>"111001100",
  64320=>"000010010",
  64321=>"000000110",
  64322=>"010011011",
  64323=>"110001101",
  64324=>"011011011",
  64325=>"101111111",
  64326=>"100000001",
  64327=>"110000111",
  64328=>"111111010",
  64329=>"111101000",
  64330=>"000100110",
  64331=>"101001000",
  64332=>"101000000",
  64333=>"101110110",
  64334=>"110011011",
  64335=>"011100000",
  64336=>"000001000",
  64337=>"111000000",
  64338=>"100100111",
  64339=>"001101011",
  64340=>"101111100",
  64341=>"001000001",
  64342=>"000010000",
  64343=>"010000000",
  64344=>"111111011",
  64345=>"011000100",
  64346=>"000110100",
  64347=>"011100110",
  64348=>"101000000",
  64349=>"110110110",
  64350=>"010111110",
  64351=>"011101101",
  64352=>"001001101",
  64353=>"000001101",
  64354=>"000111111",
  64355=>"011011011",
  64356=>"011111111",
  64357=>"010110111",
  64358=>"010000110",
  64359=>"111101101",
  64360=>"101110000",
  64361=>"111101111",
  64362=>"000011100",
  64363=>"000000011",
  64364=>"011000000",
  64365=>"011111111",
  64366=>"000101101",
  64367=>"000010011",
  64368=>"110110110",
  64369=>"110010001",
  64370=>"001101111",
  64371=>"000100001",
  64372=>"000000000",
  64373=>"100111111",
  64374=>"000000000",
  64375=>"000111111",
  64376=>"000010111",
  64377=>"111010110",
  64378=>"001000101",
  64379=>"010100111",
  64380=>"011001001",
  64381=>"000011111",
  64382=>"000101000",
  64383=>"111100100",
  64384=>"000000010",
  64385=>"101100111",
  64386=>"111001110",
  64387=>"111000000",
  64388=>"101000000",
  64389=>"111000001",
  64390=>"000000100",
  64391=>"000010000",
  64392=>"111001011",
  64393=>"001001111",
  64394=>"110000101",
  64395=>"000100010",
  64396=>"110101000",
  64397=>"000100001",
  64398=>"110000001",
  64399=>"000000000",
  64400=>"011111111",
  64401=>"001000000",
  64402=>"000101100",
  64403=>"011111110",
  64404=>"100000000",
  64405=>"011000000",
  64406=>"111111111",
  64407=>"011000100",
  64408=>"000100001",
  64409=>"000010001",
  64410=>"111110100",
  64411=>"000000000",
  64412=>"110100101",
  64413=>"011001000",
  64414=>"001100111",
  64415=>"101001000",
  64416=>"111111111",
  64417=>"010010100",
  64418=>"011011000",
  64419=>"101000000",
  64420=>"011111011",
  64421=>"101100100",
  64422=>"110000000",
  64423=>"010010010",
  64424=>"111111010",
  64425=>"000000000",
  64426=>"111000000",
  64427=>"000110111",
  64428=>"010101101",
  64429=>"000000101",
  64430=>"111011111",
  64431=>"011000000",
  64432=>"001011001",
  64433=>"011110110",
  64434=>"010111011",
  64435=>"010011001",
  64436=>"011000000",
  64437=>"001111111",
  64438=>"011011010",
  64439=>"000000000",
  64440=>"011111100",
  64441=>"111001001",
  64442=>"000000000",
  64443=>"100110110",
  64444=>"000010100",
  64445=>"111111111",
  64446=>"010100100",
  64447=>"000000000",
  64448=>"000010111",
  64449=>"101000100",
  64450=>"000100100",
  64451=>"100110110",
  64452=>"010000101",
  64453=>"001001000",
  64454=>"000000000",
  64455=>"000000111",
  64456=>"110111111",
  64457=>"000000000",
  64458=>"100000000",
  64459=>"111000111",
  64460=>"100100100",
  64461=>"110100101",
  64462=>"011101100",
  64463=>"001111111",
  64464=>"111000000",
  64465=>"010100110",
  64466=>"111111100",
  64467=>"010100000",
  64468=>"000000001",
  64469=>"001011011",
  64470=>"011001011",
  64471=>"000111111",
  64472=>"110100100",
  64473=>"101101000",
  64474=>"111111011",
  64475=>"011111111",
  64476=>"110010110",
  64477=>"011100000",
  64478=>"111000000",
  64479=>"000000000",
  64480=>"000000000",
  64481=>"000010111",
  64482=>"110100101",
  64483=>"000111011",
  64484=>"000000000",
  64485=>"000000100",
  64486=>"101101000",
  64487=>"010110111",
  64488=>"000111010",
  64489=>"001111000",
  64490=>"111010110",
  64491=>"000000000",
  64492=>"001000000",
  64493=>"010000000",
  64494=>"101000011",
  64495=>"111000100",
  64496=>"100111111",
  64497=>"001100100",
  64498=>"111001110",
  64499=>"111011010",
  64500=>"001001001",
  64501=>"110100000",
  64502=>"000000010",
  64503=>"111101101",
  64504=>"111111110",
  64505=>"000100101",
  64506=>"100000010",
  64507=>"000000100",
  64508=>"000010111",
  64509=>"111101101",
  64510=>"100100010",
  64511=>"000001101",
  64512=>"101110100",
  64513=>"100110000",
  64514=>"011001001",
  64515=>"100110000",
  64516=>"011111000",
  64517=>"000100100",
  64518=>"001001111",
  64519=>"111111011",
  64520=>"001011011",
  64521=>"011011010",
  64522=>"111000001",
  64523=>"000000000",
  64524=>"000000111",
  64525=>"100100000",
  64526=>"100001011",
  64527=>"011101111",
  64528=>"110101000",
  64529=>"100000100",
  64530=>"111110101",
  64531=>"110111001",
  64532=>"000100111",
  64533=>"000110100",
  64534=>"101000101",
  64535=>"101000000",
  64536=>"100100000",
  64537=>"000100100",
  64538=>"100110000",
  64539=>"111001111",
  64540=>"101100110",
  64541=>"010011011",
  64542=>"000110100",
  64543=>"001001011",
  64544=>"001011000",
  64545=>"100100100",
  64546=>"001110110",
  64547=>"111011011",
  64548=>"001011011",
  64549=>"000100000",
  64550=>"011001001",
  64551=>"110111110",
  64552=>"000011000",
  64553=>"100100000",
  64554=>"000000011",
  64555=>"011010000",
  64556=>"111111101",
  64557=>"110000100",
  64558=>"000100110",
  64559=>"000100000",
  64560=>"000100100",
  64561=>"001001001",
  64562=>"100110100",
  64563=>"100101100",
  64564=>"100110011",
  64565=>"101000000",
  64566=>"001011110",
  64567=>"111111011",
  64568=>"100100100",
  64569=>"100100110",
  64570=>"110110100",
  64571=>"110110110",
  64572=>"000001001",
  64573=>"011011011",
  64574=>"000100100",
  64575=>"011011111",
  64576=>"111111111",
  64577=>"110100011",
  64578=>"101111111",
  64579=>"011011110",
  64580=>"100110111",
  64581=>"100110100",
  64582=>"001001110",
  64583=>"000011111",
  64584=>"100010000",
  64585=>"011011000",
  64586=>"100100000",
  64587=>"101100100",
  64588=>"010001001",
  64589=>"011000101",
  64590=>"000111111",
  64591=>"011100000",
  64592=>"011011010",
  64593=>"011011100",
  64594=>"111111110",
  64595=>"000100010",
  64596=>"011100100",
  64597=>"100110001",
  64598=>"111111101",
  64599=>"111100110",
  64600=>"110110110",
  64601=>"110110000",
  64602=>"001000001",
  64603=>"100110110",
  64604=>"100100100",
  64605=>"000100001",
  64606=>"100100100",
  64607=>"101011111",
  64608=>"011001011",
  64609=>"111110000",
  64610=>"011001111",
  64611=>"110101111",
  64612=>"010111111",
  64613=>"001011000",
  64614=>"111001111",
  64615=>"011011011",
  64616=>"000110011",
  64617=>"110110000",
  64618=>"001000110",
  64619=>"000110111",
  64620=>"100110001",
  64621=>"110001010",
  64622=>"000001111",
  64623=>"000100101",
  64624=>"110111001",
  64625=>"100110100",
  64626=>"011001001",
  64627=>"100110011",
  64628=>"111110111",
  64629=>"100100100",
  64630=>"110100000",
  64631=>"011001001",
  64632=>"001010001",
  64633=>"111000000",
  64634=>"000100100",
  64635=>"100110011",
  64636=>"010011001",
  64637=>"010110100",
  64638=>"011011011",
  64639=>"011001011",
  64640=>"000101111",
  64641=>"010010001",
  64642=>"111000110",
  64643=>"111110011",
  64644=>"010100100",
  64645=>"111000111",
  64646=>"011110100",
  64647=>"111111110",
  64648=>"000001011",
  64649=>"111011111",
  64650=>"111101100",
  64651=>"000110111",
  64652=>"011001001",
  64653=>"101001110",
  64654=>"001111001",
  64655=>"000100100",
  64656=>"000011001",
  64657=>"001010011",
  64658=>"000011011",
  64659=>"011110110",
  64660=>"000000010",
  64661=>"100100110",
  64662=>"101100001",
  64663=>"000100100",
  64664=>"000001000",
  64665=>"001100100",
  64666=>"111011000",
  64667=>"100001001",
  64668=>"100111110",
  64669=>"011011011",
  64670=>"100100110",
  64671=>"000000000",
  64672=>"100111011",
  64673=>"110100100",
  64674=>"011000010",
  64675=>"100101001",
  64676=>"110000110",
  64677=>"001001011",
  64678=>"101100100",
  64679=>"010001011",
  64680=>"100100100",
  64681=>"110010000",
  64682=>"110111100",
  64683=>"110110011",
  64684=>"111111011",
  64685=>"001000000",
  64686=>"011110001",
  64687=>"000001011",
  64688=>"100000010",
  64689=>"001001000",
  64690=>"100100110",
  64691=>"111110011",
  64692=>"011011011",
  64693=>"000000011",
  64694=>"100110110",
  64695=>"000100000",
  64696=>"000100110",
  64697=>"000000000",
  64698=>"001011000",
  64699=>"001011111",
  64700=>"000100000",
  64701=>"011011011",
  64702=>"011001001",
  64703=>"000000100",
  64704=>"001011111",
  64705=>"111011011",
  64706=>"110111001",
  64707=>"001001001",
  64708=>"100100000",
  64709=>"000100100",
  64710=>"000000100",
  64711=>"010011000",
  64712=>"011001011",
  64713=>"010000000",
  64714=>"100110001",
  64715=>"101011111",
  64716=>"001001010",
  64717=>"001011011",
  64718=>"011011000",
  64719=>"001001111",
  64720=>"100011111",
  64721=>"011101011",
  64722=>"001100000",
  64723=>"001001110",
  64724=>"011011011",
  64725=>"111111000",
  64726=>"100010000",
  64727=>"000110100",
  64728=>"001011111",
  64729=>"100000000",
  64730=>"010100101",
  64731=>"100100100",
  64732=>"111110100",
  64733=>"110110101",
  64734=>"110100110",
  64735=>"000100100",
  64736=>"001000001",
  64737=>"000101100",
  64738=>"011011111",
  64739=>"111011010",
  64740=>"101001001",
  64741=>"110010100",
  64742=>"011011011",
  64743=>"011011111",
  64744=>"010110100",
  64745=>"001000010",
  64746=>"000000000",
  64747=>"111001000",
  64748=>"100000000",
  64749=>"111111110",
  64750=>"000000000",
  64751=>"100000000",
  64752=>"001110110",
  64753=>"101111100",
  64754=>"100100100",
  64755=>"111111101",
  64756=>"000111110",
  64757=>"110111111",
  64758=>"100101101",
  64759=>"101000000",
  64760=>"100100110",
  64761=>"110010110",
  64762=>"100100100",
  64763=>"011111001",
  64764=>"111010011",
  64765=>"110001101",
  64766=>"100010111",
  64767=>"111010010",
  64768=>"100000000",
  64769=>"111110101",
  64770=>"110000100",
  64771=>"011011011",
  64772=>"100000000",
  64773=>"111000000",
  64774=>"110110110",
  64775=>"011110011",
  64776=>"000110111",
  64777=>"011110100",
  64778=>"100100000",
  64779=>"100010011",
  64780=>"001011111",
  64781=>"000011111",
  64782=>"000001001",
  64783=>"110011011",
  64784=>"100100110",
  64785=>"000100110",
  64786=>"000001011",
  64787=>"100110011",
  64788=>"100110011",
  64789=>"011001000",
  64790=>"111010000",
  64791=>"100100100",
  64792=>"110110110",
  64793=>"111111111",
  64794=>"000001101",
  64795=>"000011001",
  64796=>"010011011",
  64797=>"000100100",
  64798=>"000100110",
  64799=>"000000100",
  64800=>"111100100",
  64801=>"000011001",
  64802=>"101100100",
  64803=>"110000100",
  64804=>"100110000",
  64805=>"000111111",
  64806=>"100100100",
  64807=>"000111000",
  64808=>"111010110",
  64809=>"000000100",
  64810=>"001100100",
  64811=>"011000011",
  64812=>"001100011",
  64813=>"000110111",
  64814=>"001000100",
  64815=>"011111011",
  64816=>"100100011",
  64817=>"000001000",
  64818=>"000000001",
  64819=>"100111111",
  64820=>"100000000",
  64821=>"100111011",
  64822=>"100100110",
  64823=>"010111100",
  64824=>"011000000",
  64825=>"000000100",
  64826=>"000000010",
  64827=>"100111111",
  64828=>"001100110",
  64829=>"111111110",
  64830=>"000101101",
  64831=>"110111110",
  64832=>"110110110",
  64833=>"100110010",
  64834=>"011001000",
  64835=>"001001100",
  64836=>"110100110",
  64837=>"100000100",
  64838=>"111110110",
  64839=>"011001000",
  64840=>"001110110",
  64841=>"101011111",
  64842=>"100100110",
  64843=>"000100101",
  64844=>"111110100",
  64845=>"000100110",
  64846=>"100111110",
  64847=>"111100001",
  64848=>"000000000",
  64849=>"111111001",
  64850=>"111110111",
  64851=>"000010010",
  64852=>"000011011",
  64853=>"001000000",
  64854=>"001100110",
  64855=>"000011011",
  64856=>"001011101",
  64857=>"010010100",
  64858=>"101001100",
  64859=>"001001100",
  64860=>"010111011",
  64861=>"001000101",
  64862=>"111111110",
  64863=>"110100000",
  64864=>"110110110",
  64865=>"000000100",
  64866=>"110110100",
  64867=>"011001011",
  64868=>"100000010",
  64869=>"000010100",
  64870=>"000001011",
  64871=>"111001011",
  64872=>"101110110",
  64873=>"010100100",
  64874=>"011011011",
  64875=>"111100110",
  64876=>"111000111",
  64877=>"000000011",
  64878=>"011011000",
  64879=>"010000111",
  64880=>"100110110",
  64881=>"001111011",
  64882=>"100100100",
  64883=>"101000100",
  64884=>"011011011",
  64885=>"100100100",
  64886=>"011011010",
  64887=>"000111011",
  64888=>"011000011",
  64889=>"000100110",
  64890=>"100100100",
  64891=>"001011111",
  64892=>"100110110",
  64893=>"100000000",
  64894=>"011011100",
  64895=>"000011000",
  64896=>"110110010",
  64897=>"111100000",
  64898=>"000111110",
  64899=>"000101000",
  64900=>"000100011",
  64901=>"001101111",
  64902=>"110010001",
  64903=>"100000001",
  64904=>"100100101",
  64905=>"100110111",
  64906=>"110110100",
  64907=>"011111110",
  64908=>"101011100",
  64909=>"000111111",
  64910=>"001111111",
  64911=>"100100100",
  64912=>"100111110",
  64913=>"111111000",
  64914=>"000010000",
  64915=>"000100110",
  64916=>"000000100",
  64917=>"000000000",
  64918=>"101100111",
  64919=>"110000000",
  64920=>"111111011",
  64921=>"000000011",
  64922=>"111000000",
  64923=>"001000011",
  64924=>"110011001",
  64925=>"000100100",
  64926=>"000001111",
  64927=>"110100111",
  64928=>"111110110",
  64929=>"100111110",
  64930=>"101000000",
  64931=>"100110111",
  64932=>"000000111",
  64933=>"100111110",
  64934=>"100100101",
  64935=>"111111111",
  64936=>"000100000",
  64937=>"001011011",
  64938=>"111011011",
  64939=>"111000000",
  64940=>"000011101",
  64941=>"000011000",
  64942=>"001100111",
  64943=>"011001011",
  64944=>"111011000",
  64945=>"010011010",
  64946=>"111101000",
  64947=>"001000000",
  64948=>"010011011",
  64949=>"101101000",
  64950=>"000011011",
  64951=>"100010111",
  64952=>"110000001",
  64953=>"000110100",
  64954=>"011001000",
  64955=>"100000011",
  64956=>"111101000",
  64957=>"011011011",
  64958=>"000001001",
  64959=>"111011000",
  64960=>"010100100",
  64961=>"000001000",
  64962=>"001011011",
  64963=>"101001000",
  64964=>"000000110",
  64965=>"100100111",
  64966=>"111110000",
  64967=>"001000100",
  64968=>"000100010",
  64969=>"010111111",
  64970=>"110010010",
  64971=>"100100111",
  64972=>"110011000",
  64973=>"000000110",
  64974=>"110000100",
  64975=>"100011011",
  64976=>"011011000",
  64977=>"000000000",
  64978=>"100010011",
  64979=>"101111000",
  64980=>"111111111",
  64981=>"100000101",
  64982=>"111100111",
  64983=>"111100000",
  64984=>"011111111",
  64985=>"000000111",
  64986=>"101111111",
  64987=>"111100111",
  64988=>"100110110",
  64989=>"000001011",
  64990=>"001011111",
  64991=>"000000001",
  64992=>"010010000",
  64993=>"101011011",
  64994=>"001011011",
  64995=>"100110110",
  64996=>"100110000",
  64997=>"001000010",
  64998=>"011101101",
  64999=>"110110001",
  65000=>"011011101",
  65001=>"100111001",
  65002=>"000100110",
  65003=>"101000100",
  65004=>"011011011",
  65005=>"111111110",
  65006=>"110000000",
  65007=>"000100000",
  65008=>"000100100",
  65009=>"100000111",
  65010=>"011000000",
  65011=>"011011010",
  65012=>"000110100",
  65013=>"111101111",
  65014=>"011011111",
  65015=>"001001001",
  65016=>"100100000",
  65017=>"011001001",
  65018=>"111100100",
  65019=>"000000111",
  65020=>"111000000",
  65021=>"001011100",
  65022=>"100110101",
  65023=>"000000111",
  65024=>"011001101",
  65025=>"110101100",
  65026=>"000000110",
  65027=>"000000110",
  65028=>"001010110",
  65029=>"000010010",
  65030=>"110110000",
  65031=>"011111111",
  65032=>"001000111",
  65033=>"001000000",
  65034=>"000111111",
  65035=>"000011110",
  65036=>"001001101",
  65037=>"000000000",
  65038=>"010001011",
  65039=>"111100011",
  65040=>"111110010",
  65041=>"111000000",
  65042=>"110101100",
  65043=>"011110000",
  65044=>"101101101",
  65045=>"111111101",
  65046=>"110010010",
  65047=>"010111000",
  65048=>"000111000",
  65049=>"111000000",
  65050=>"011011000",
  65051=>"000010010",
  65052=>"101001000",
  65053=>"000000000",
  65054=>"110111011",
  65055=>"000000101",
  65056=>"000000111",
  65057=>"000000000",
  65058=>"000101100",
  65059=>"000011010",
  65060=>"011000100",
  65061=>"110001011",
  65062=>"010111111",
  65063=>"101001000",
  65064=>"111010111",
  65065=>"000011000",
  65066=>"100111111",
  65067=>"111011000",
  65068=>"111100001",
  65069=>"101101000",
  65070=>"111000101",
  65071=>"010001000",
  65072=>"111000000",
  65073=>"001011011",
  65074=>"010000000",
  65075=>"001000000",
  65076=>"110011111",
  65077=>"011101101",
  65078=>"111110101",
  65079=>"111101000",
  65080=>"111000000",
  65081=>"000000000",
  65082=>"000000100",
  65083=>"010000001",
  65084=>"100000000",
  65085=>"010001000",
  65086=>"000101100",
  65087=>"011111111",
  65088=>"110011000",
  65089=>"111000101",
  65090=>"101000101",
  65091=>"001010011",
  65092=>"000010000",
  65093=>"001101111",
  65094=>"001000000",
  65095=>"111101000",
  65096=>"111001100",
  65097=>"000011111",
  65098=>"000100101",
  65099=>"111111101",
  65100=>"111000001",
  65101=>"000001011",
  65102=>"000000111",
  65103=>"111111111",
  65104=>"000000000",
  65105=>"110000000",
  65106=>"111111001",
  65107=>"011001110",
  65108=>"110111001",
  65109=>"111111000",
  65110=>"011001001",
  65111=>"101010011",
  65112=>"000000000",
  65113=>"000000101",
  65114=>"000111111",
  65115=>"110000100",
  65116=>"111111000",
  65117=>"000001111",
  65118=>"011000111",
  65119=>"000000110",
  65120=>"111111111",
  65121=>"000000110",
  65122=>"001110111",
  65123=>"011000101",
  65124=>"000001110",
  65125=>"000010001",
  65126=>"011111111",
  65127=>"001111010",
  65128=>"001000110",
  65129=>"101000000",
  65130=>"101001011",
  65131=>"111111000",
  65132=>"111000000",
  65133=>"000111111",
  65134=>"111000000",
  65135=>"111011001",
  65136=>"101111111",
  65137=>"110001100",
  65138=>"011111011",
  65139=>"101000001",
  65140=>"111000001",
  65141=>"111000000",
  65142=>"000000001",
  65143=>"000000101",
  65144=>"000111111",
  65145=>"111101100",
  65146=>"000000000",
  65147=>"000000010",
  65148=>"000000010",
  65149=>"100000110",
  65150=>"000010111",
  65151=>"000111111",
  65152=>"010000000",
  65153=>"000000000",
  65154=>"111010000",
  65155=>"100010010",
  65156=>"101101101",
  65157=>"110101111",
  65158=>"111001101",
  65159=>"100000100",
  65160=>"000011111",
  65161=>"100011111",
  65162=>"000111111",
  65163=>"100110110",
  65164=>"000110111",
  65165=>"111111101",
  65166=>"010001000",
  65167=>"000000001",
  65168=>"111001101",
  65169=>"000000111",
  65170=>"000010000",
  65171=>"000000001",
  65172=>"010010010",
  65173=>"111010010",
  65174=>"100011111",
  65175=>"000000001",
  65176=>"111011000",
  65177=>"111110100",
  65178=>"000000010",
  65179=>"000001111",
  65180=>"110001010",
  65181=>"000000111",
  65182=>"101000000",
  65183=>"111000000",
  65184=>"000000111",
  65185=>"000100000",
  65186=>"000111111",
  65187=>"100010101",
  65188=>"111111000",
  65189=>"110000011",
  65190=>"011110110",
  65191=>"000100111",
  65192=>"111010000",
  65193=>"000001000",
  65194=>"110110111",
  65195=>"000000000",
  65196=>"111111111",
  65197=>"011000010",
  65198=>"100101110",
  65199=>"001111100",
  65200=>"101111110",
  65201=>"001001001",
  65202=>"000001111",
  65203=>"000001100",
  65204=>"011111110",
  65205=>"000111101",
  65206=>"111111100",
  65207=>"000011111",
  65208=>"001000010",
  65209=>"000011010",
  65210=>"100010000",
  65211=>"101000011",
  65212=>"000000101",
  65213=>"000001111",
  65214=>"000111111",
  65215=>"111000000",
  65216=>"111101101",
  65217=>"110111000",
  65218=>"101010000",
  65219=>"001001101",
  65220=>"111000000",
  65221=>"110110100",
  65222=>"111111100",
  65223=>"000000000",
  65224=>"011001111",
  65225=>"111010010",
  65226=>"111010000",
  65227=>"011010010",
  65228=>"000110111",
  65229=>"000011100",
  65230=>"000111100",
  65231=>"000110000",
  65232=>"000010111",
  65233=>"011001110",
  65234=>"010000000",
  65235=>"001000010",
  65236=>"000011001",
  65237=>"100101111",
  65238=>"100010010",
  65239=>"011000000",
  65240=>"111100000",
  65241=>"011011000",
  65242=>"000001111",
  65243=>"010000101",
  65244=>"111000000",
  65245=>"101100111",
  65246=>"010110000",
  65247=>"000111100",
  65248=>"101000010",
  65249=>"111000111",
  65250=>"000000010",
  65251=>"111100110",
  65252=>"001100000",
  65253=>"010101101",
  65254=>"011000111",
  65255=>"111101101",
  65256=>"100011000",
  65257=>"111111101",
  65258=>"001010111",
  65259=>"111010000",
  65260=>"000011111",
  65261=>"110000100",
  65262=>"000000000",
  65263=>"100011100",
  65264=>"111111010",
  65265=>"111011111",
  65266=>"111000010",
  65267=>"111111001",
  65268=>"110100101",
  65269=>"000101111",
  65270=>"000001001",
  65271=>"110000001",
  65272=>"111000000",
  65273=>"000111111",
  65274=>"111000100",
  65275=>"001111101",
  65276=>"000111110",
  65277=>"111111000",
  65278=>"110010111",
  65279=>"100100000",
  65280=>"000001001",
  65281=>"001000111",
  65282=>"000000000",
  65283=>"000000110",
  65284=>"111000101",
  65285=>"000000111",
  65286=>"000101110",
  65287=>"000000010",
  65288=>"101000000",
  65289=>"000110111",
  65290=>"000010110",
  65291=>"111000010",
  65292=>"000000000",
  65293=>"110010001",
  65294=>"000000000",
  65295=>"110111111",
  65296=>"000001001",
  65297=>"111111111",
  65298=>"010000101",
  65299=>"000111110",
  65300=>"001100110",
  65301=>"001000000",
  65302=>"011101100",
  65303=>"010010111",
  65304=>"000000000",
  65305=>"111000111",
  65306=>"100100001",
  65307=>"000111100",
  65308=>"000101110",
  65309=>"101100100",
  65310=>"101000000",
  65311=>"101101101",
  65312=>"100001100",
  65313=>"110111011",
  65314=>"000000010",
  65315=>"000111111",
  65316=>"000000011",
  65317=>"000000111",
  65318=>"011001000",
  65319=>"000101111",
  65320=>"111111010",
  65321=>"110100111",
  65322=>"000111111",
  65323=>"001011110",
  65324=>"111011111",
  65325=>"000000000",
  65326=>"000000000",
  65327=>"010101110",
  65328=>"001001000",
  65329=>"000100000",
  65330=>"000000011",
  65331=>"000101100",
  65332=>"010111111",
  65333=>"111111111",
  65334=>"110111011",
  65335=>"100010011",
  65336=>"101000111",
  65337=>"000101101",
  65338=>"000110000",
  65339=>"101000000",
  65340=>"100001000",
  65341=>"111111000",
  65342=>"101010110",
  65343=>"010111001",
  65344=>"111111111",
  65345=>"010101011",
  65346=>"011000111",
  65347=>"000001111",
  65348=>"010111010",
  65349=>"001000111",
  65350=>"000111111",
  65351=>"110001010",
  65352=>"000100111",
  65353=>"110111111",
  65354=>"000001000",
  65355=>"000010001",
  65356=>"000000010",
  65357=>"000011111",
  65358=>"111100110",
  65359=>"010010111",
  65360=>"111111111",
  65361=>"111111000",
  65362=>"000100110",
  65363=>"001100110",
  65364=>"110100000",
  65365=>"100000110",
  65366=>"000101111",
  65367=>"000000000",
  65368=>"000001101",
  65369=>"111001011",
  65370=>"000111111",
  65371=>"011011110",
  65372=>"111111111",
  65373=>"000000000",
  65374=>"010110101",
  65375=>"000010111",
  65376=>"110101111",
  65377=>"000111110",
  65378=>"000101111",
  65379=>"010110100",
  65380=>"000100100",
  65381=>"111111100",
  65382=>"010111110",
  65383=>"000011111",
  65384=>"000101011",
  65385=>"000000000",
  65386=>"000000110",
  65387=>"010001110",
  65388=>"010000100",
  65389=>"000000010",
  65390=>"000001001",
  65391=>"111111001",
  65392=>"100000010",
  65393=>"111110111",
  65394=>"011111110",
  65395=>"000001011",
  65396=>"000000011",
  65397=>"000000000",
  65398=>"000110011",
  65399=>"111111111",
  65400=>"011010111",
  65401=>"110111101",
  65402=>"000001000",
  65403=>"111000111",
  65404=>"001011010",
  65405=>"110000010",
  65406=>"111100001",
  65407=>"000001000",
  65408=>"110110100",
  65409=>"111101000",
  65410=>"111001000",
  65411=>"111111010",
  65412=>"001101000",
  65413=>"111101100",
  65414=>"110100110",
  65415=>"001000000",
  65416=>"001000100",
  65417=>"000001101",
  65418=>"010011010",
  65419=>"101110111",
  65420=>"101101011",
  65421=>"111100101",
  65422=>"111000000",
  65423=>"000000000",
  65424=>"001001011",
  65425=>"010101111",
  65426=>"000000010",
  65427=>"000000000",
  65428=>"101000100",
  65429=>"000000010",
  65430=>"100111001",
  65431=>"010011011",
  65432=>"010000111",
  65433=>"001000011",
  65434=>"011110111",
  65435=>"101000000",
  65436=>"000100101",
  65437=>"111111010",
  65438=>"000000111",
  65439=>"100111011",
  65440=>"011000000",
  65441=>"110000000",
  65442=>"111100010",
  65443=>"000010000",
  65444=>"111001010",
  65445=>"110000000",
  65446=>"001111000",
  65447=>"010110110",
  65448=>"000000000",
  65449=>"110111000",
  65450=>"111010000",
  65451=>"000110110",
  65452=>"100000101",
  65453=>"000101010",
  65454=>"000010011",
  65455=>"111011110",
  65456=>"011000000",
  65457=>"000001100",
  65458=>"010100000",
  65459=>"001000100",
  65460=>"111000001",
  65461=>"111010100",
  65462=>"111111101",
  65463=>"001101111",
  65464=>"001100000",
  65465=>"100000001",
  65466=>"001000000",
  65467=>"000000010",
  65468=>"000010000",
  65469=>"000100111",
  65470=>"001000000",
  65471=>"010010111",
  65472=>"000000000",
  65473=>"000000000",
  65474=>"010000111",
  65475=>"000101001",
  65476=>"000001000",
  65477=>"100000011",
  65478=>"000000001",
  65479=>"010011000",
  65480=>"101000101",
  65481=>"110010000",
  65482=>"111010010",
  65483=>"110000000",
  65484=>"000000000",
  65485=>"100110110",
  65486=>"011010010",
  65487=>"111111011",
  65488=>"100000010",
  65489=>"110100111",
  65490=>"111000011",
  65491=>"110000010",
  65492=>"101101111",
  65493=>"000100100",
  65494=>"010101111",
  65495=>"001111001",
  65496=>"000000111",
  65497=>"111000000",
  65498=>"111110000",
  65499=>"000000111",
  65500=>"110001001",
  65501=>"111110010",
  65502=>"111111000",
  65503=>"111011001",
  65504=>"000111111",
  65505=>"001001000",
  65506=>"000000110",
  65507=>"000000010",
  65508=>"010000000",
  65509=>"111001000",
  65510=>"111000110",
  65511=>"111101100",
  65512=>"111000111",
  65513=>"111111110",
  65514=>"000100010",
  65515=>"000000111",
  65516=>"001001000",
  65517=>"111011111",
  65518=>"000000000",
  65519=>"001111001",
  65520=>"111000000",
  65521=>"001000010",
  65522=>"010000010",
  65523=>"111001101",
  65524=>"100101111",
  65525=>"000001000",
  65526=>"000010010",
  65527=>"001001101",
  65528=>"000000111",
  65529=>"000000101",
  65530=>"111011110",
  65531=>"101001000",
  65532=>"000011001",
  65533=>"111100110",
  65534=>"000111111",
  65535=>"000000000");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;