LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L2_2_BNROM IS
    PORT (
        coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); -- Instruction bus
        address : IN unsigned(3 DOWNTO 0));
END L2_2_BNROM;

ARCHITECTURE RTL OF L2_2_BNROM IS

    TYPE ROM_mem IS ARRAY (0 TO 15) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem :=
    (0=>"0000111000100000"&"0010001110111010",
    1=>"0011000000100111"&"0001010001101011",
    2=>"0000100100010100"&"0001100010001000",
    3=>"0001010101001000"&"0001011010100010",
    4=>"0000010110010101"&"0001000010110011",
    5=>"0010001010101110"&"0001101000001001",
    6=>"0001000100001001"&"0001100000000001",
    7=>"0001000101010001"&"0001001011101100",
    8=>"0000110101010010"&"0010001000101001",
    9=>"0001000011110100"&"0001110010011100",
    10=>"0010010111101011"&"0001101111101001",
    11=>"0000111111011110"&"0010000000000100",
    12=>"0001001100110000"&"0001011010101100",
    13=>"0001111011100110"&"0001011001111010",
    14=>"1111100000011011"&"0001110000011000",
    15=>"0000110101010101"&"0001011100010110");
BEGIN
    coefs <= ROM_content(to_integer(address));
END RTL;