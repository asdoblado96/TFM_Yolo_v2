LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_12_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_12_WROM;

ARCHITECTURE RTL OF L8_12_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"000010111",
  1=>"100110001",
  2=>"001010001",
  3=>"001000110",
  4=>"000010101",
  5=>"100111100",
  6=>"101000011",
  7=>"100000001",
  8=>"110111010",
  9=>"100010001",
  10=>"000101100",
  11=>"111100010",
  12=>"110001111",
  13=>"110001111",
  14=>"000100001",
  15=>"100000111",
  16=>"101100110",
  17=>"000010010",
  18=>"101100100",
  19=>"011111000",
  20=>"101010011",
  21=>"101001010",
  22=>"010110011",
  23=>"001011111",
  24=>"011101111",
  25=>"100110100",
  26=>"110110111",
  27=>"011111011",
  28=>"100101111",
  29=>"000101110",
  30=>"100110000",
  31=>"111110010",
  32=>"001110101",
  33=>"100100011",
  34=>"000001010",
  35=>"011110111",
  36=>"010100100",
  37=>"001110010",
  38=>"111001001",
  39=>"010011000",
  40=>"000001000",
  41=>"000000000",
  42=>"001111011",
  43=>"010010111",
  44=>"000000010",
  45=>"110001110",
  46=>"010010000",
  47=>"110000011",
  48=>"101000101",
  49=>"100010010",
  50=>"000010110",
  51=>"000101000",
  52=>"101001101",
  53=>"111011000",
  54=>"100001101",
  55=>"110001111",
  56=>"100100100",
  57=>"011111001",
  58=>"110111010",
  59=>"110000101",
  60=>"100010110",
  61=>"000000000",
  62=>"001000011",
  63=>"101000100",
  64=>"110111000",
  65=>"001100010",
  66=>"101011001",
  67=>"101110010",
  68=>"010111011",
  69=>"001011101",
  70=>"101001111",
  71=>"010111101",
  72=>"000011010",
  73=>"110000001",
  74=>"000100010",
  75=>"110000011",
  76=>"001100000",
  77=>"111010111",
  78=>"111010001",
  79=>"011000110",
  80=>"011010100",
  81=>"010011111",
  82=>"110011001",
  83=>"011000100",
  84=>"000010100",
  85=>"010000000",
  86=>"111001111",
  87=>"000111001",
  88=>"101111111",
  89=>"000000010",
  90=>"101100110",
  91=>"010100000",
  92=>"110101011",
  93=>"010111101",
  94=>"001010111",
  95=>"010111001",
  96=>"110000010",
  97=>"100100010",
  98=>"111110110",
  99=>"011001101",
  100=>"111011101",
  101=>"000011001",
  102=>"011100111",
  103=>"000101000",
  104=>"011100011",
  105=>"010000101",
  106=>"010000000",
  107=>"101010011",
  108=>"010000000",
  109=>"111111111",
  110=>"100010100",
  111=>"001101001",
  112=>"001111001",
  113=>"101101101",
  114=>"011110010",
  115=>"011001111",
  116=>"000000110",
  117=>"011001011",
  118=>"000100010",
  119=>"101110100",
  120=>"010101100",
  121=>"000111000",
  122=>"000111101",
  123=>"100100010",
  124=>"000010110",
  125=>"001010111",
  126=>"110000100",
  127=>"000101100",
  128=>"000100000",
  129=>"001010010",
  130=>"011111001",
  131=>"111111001",
  132=>"100011111",
  133=>"000001011",
  134=>"111100001",
  135=>"001001100",
  136=>"000100111",
  137=>"111010000",
  138=>"011010111",
  139=>"101001010",
  140=>"111111010",
  141=>"111101101",
  142=>"101001100",
  143=>"110110111",
  144=>"010000001",
  145=>"111000110",
  146=>"111001101",
  147=>"110101101",
  148=>"111100110",
  149=>"111000111",
  150=>"001100001",
  151=>"111111100",
  152=>"000001000",
  153=>"100111111",
  154=>"010111100",
  155=>"101000010",
  156=>"001101000",
  157=>"011001011",
  158=>"110000000",
  159=>"010100110",
  160=>"010100110",
  161=>"010010111",
  162=>"111001101",
  163=>"011001100",
  164=>"011101010",
  165=>"111111111",
  166=>"010001110",
  167=>"110110110",
  168=>"010000011",
  169=>"101101001",
  170=>"100110001",
  171=>"001000111",
  172=>"010011110",
  173=>"011011111",
  174=>"010101001",
  175=>"000010010",
  176=>"111001100",
  177=>"001111111",
  178=>"010001110",
  179=>"111100101",
  180=>"000010000",
  181=>"110100100",
  182=>"011000110",
  183=>"010000011",
  184=>"011001101",
  185=>"111010110",
  186=>"110001000",
  187=>"101011000",
  188=>"100101000",
  189=>"101010100",
  190=>"011100100",
  191=>"010110100",
  192=>"111111011",
  193=>"000111110",
  194=>"100110010",
  195=>"010100111",
  196=>"110101001",
  197=>"000001100",
  198=>"011010111",
  199=>"111111101",
  200=>"100000000",
  201=>"001011011",
  202=>"111101111",
  203=>"011000110",
  204=>"101100000",
  205=>"110100010",
  206=>"010001010",
  207=>"001001010",
  208=>"011110000",
  209=>"000011000",
  210=>"001011001",
  211=>"011110111",
  212=>"110100100",
  213=>"000111000",
  214=>"000001111",
  215=>"111101111",
  216=>"100011110",
  217=>"111011110",
  218=>"110110000",
  219=>"100011011",
  220=>"010100000",
  221=>"001111100",
  222=>"001000101",
  223=>"101000001",
  224=>"100110100",
  225=>"000101111",
  226=>"110000011",
  227=>"111010111",
  228=>"101110010",
  229=>"100111000",
  230=>"100111100",
  231=>"111000000",
  232=>"001101001",
  233=>"000011101",
  234=>"101000011",
  235=>"001000001",
  236=>"111111101",
  237=>"011110110",
  238=>"110101000",
  239=>"101000000",
  240=>"010100101",
  241=>"111010111",
  242=>"001010100",
  243=>"010000111",
  244=>"110010111",
  245=>"010111010",
  246=>"001110000",
  247=>"000000110",
  248=>"110100010",
  249=>"101110101",
  250=>"001100000",
  251=>"000101010",
  252=>"101011010",
  253=>"011010001",
  254=>"101101101",
  255=>"101011100",
  256=>"110011100",
  257=>"101101010",
  258=>"110110010",
  259=>"011100010",
  260=>"110010101",
  261=>"111110100",
  262=>"001011010",
  263=>"010110111",
  264=>"010100100",
  265=>"110001100",
  266=>"011100110",
  267=>"111110111",
  268=>"001001001",
  269=>"000110100",
  270=>"000001010",
  271=>"110101101",
  272=>"000000000",
  273=>"111101100",
  274=>"111101111",
  275=>"111110100",
  276=>"001010011",
  277=>"101010111",
  278=>"010000000",
  279=>"000001110",
  280=>"011010001",
  281=>"110001101",
  282=>"011011110",
  283=>"010110100",
  284=>"110000111",
  285=>"111010011",
  286=>"001000100",
  287=>"000000000",
  288=>"111000000",
  289=>"101110101",
  290=>"111011100",
  291=>"110000101",
  292=>"011100111",
  293=>"101001100",
  294=>"111110011",
  295=>"010000000",
  296=>"011001100",
  297=>"011100010",
  298=>"110110100",
  299=>"000100011",
  300=>"100111101",
  301=>"000000110",
  302=>"110000011",
  303=>"101011110",
  304=>"010111110",
  305=>"110010010",
  306=>"110001110",
  307=>"000001111",
  308=>"110110111",
  309=>"110000010",
  310=>"111100110",
  311=>"101111110",
  312=>"111011010",
  313=>"011011001",
  314=>"101101101",
  315=>"000101110",
  316=>"011010000",
  317=>"111000111",
  318=>"110101101",
  319=>"101100101",
  320=>"000001101",
  321=>"101100011",
  322=>"100110010",
  323=>"000011011",
  324=>"010111111",
  325=>"111001111",
  326=>"111100001",
  327=>"011010011",
  328=>"011000110",
  329=>"000010110",
  330=>"100100001",
  331=>"110101000",
  332=>"111000010",
  333=>"111100001",
  334=>"000000100",
  335=>"110000100",
  336=>"010000011",
  337=>"011000011",
  338=>"101100000",
  339=>"101001001",
  340=>"000000110",
  341=>"001000011",
  342=>"101001101",
  343=>"000001101",
  344=>"101000000",
  345=>"000110010",
  346=>"011000110",
  347=>"001000110",
  348=>"101111101",
  349=>"011111111",
  350=>"101001010",
  351=>"000100101",
  352=>"000110000",
  353=>"111110011",
  354=>"000011110",
  355=>"110101100",
  356=>"000100010",
  357=>"111010101",
  358=>"110100000",
  359=>"010000110",
  360=>"010101000",
  361=>"001110001",
  362=>"111111110",
  363=>"110010000",
  364=>"100011000",
  365=>"010001000",
  366=>"011000100",
  367=>"110111001",
  368=>"000110000",
  369=>"111101110",
  370=>"001111110",
  371=>"111100101",
  372=>"100001101",
  373=>"001001111",
  374=>"010101000",
  375=>"010011101",
  376=>"111110100",
  377=>"010001000",
  378=>"110100010",
  379=>"110100110",
  380=>"110001001",
  381=>"000010110",
  382=>"111110011",
  383=>"000101001",
  384=>"110110101",
  385=>"101001111",
  386=>"000111001",
  387=>"000111011",
  388=>"001001100",
  389=>"000110101",
  390=>"011001000",
  391=>"001110110",
  392=>"000101010",
  393=>"011010011",
  394=>"100100100",
  395=>"111111011",
  396=>"110110110",
  397=>"010100101",
  398=>"010010000",
  399=>"111000100",
  400=>"000000001",
  401=>"011001111",
  402=>"110111110",
  403=>"011101101",
  404=>"010101110",
  405=>"000000001",
  406=>"010000100",
  407=>"001001001",
  408=>"011000110",
  409=>"100111010",
  410=>"111010001",
  411=>"001110011",
  412=>"010100011",
  413=>"100010011",
  414=>"010010100",
  415=>"000110110",
  416=>"010010111",
  417=>"001111110",
  418=>"000001001",
  419=>"001011010",
  420=>"110010111",
  421=>"000101000",
  422=>"001101010",
  423=>"101001010",
  424=>"010001101",
  425=>"101001100",
  426=>"011110111",
  427=>"010110100",
  428=>"110101101",
  429=>"100110101",
  430=>"110001111",
  431=>"111010011",
  432=>"110110001",
  433=>"100101000",
  434=>"001011010",
  435=>"000100111",
  436=>"000100100",
  437=>"101101100",
  438=>"110100110",
  439=>"100000100",
  440=>"100001110",
  441=>"010001100",
  442=>"111110101",
  443=>"100111101",
  444=>"111100001",
  445=>"001011111",
  446=>"000100110",
  447=>"110010110",
  448=>"011111101",
  449=>"101001100",
  450=>"101110010",
  451=>"001001111",
  452=>"101101110",
  453=>"000000011",
  454=>"000111011",
  455=>"100011000",
  456=>"010010000",
  457=>"111101001",
  458=>"000010111",
  459=>"101100010",
  460=>"110101100",
  461=>"000011110",
  462=>"000000001",
  463=>"101010011",
  464=>"011010111",
  465=>"100010010",
  466=>"000000110",
  467=>"100000001",
  468=>"110011011",
  469=>"110000110",
  470=>"001101110",
  471=>"000010000",
  472=>"000000111",
  473=>"110100001",
  474=>"001001101",
  475=>"111011000",
  476=>"101001110",
  477=>"000110110",
  478=>"001010101",
  479=>"111010000",
  480=>"010010011",
  481=>"100010110",
  482=>"110110100",
  483=>"101001011",
  484=>"010001001",
  485=>"101011011",
  486=>"100000000",
  487=>"000011110",
  488=>"110010000",
  489=>"111100110",
  490=>"110001100",
  491=>"011011000",
  492=>"001001010",
  493=>"010010000",
  494=>"010000000",
  495=>"000011110",
  496=>"100101010",
  497=>"111010100",
  498=>"011010111",
  499=>"010110101",
  500=>"111000101",
  501=>"111001001",
  502=>"000110011",
  503=>"110011110",
  504=>"000100111",
  505=>"011111001",
  506=>"111001111",
  507=>"000000101",
  508=>"000101000",
  509=>"011000100",
  510=>"011100001",
  511=>"001001010",
  512=>"001110110",
  513=>"000000100",
  514=>"011100101",
  515=>"110111010",
  516=>"010010101",
  517=>"010100010",
  518=>"001110001",
  519=>"100000010",
  520=>"110010110",
  521=>"001110011",
  522=>"011110111",
  523=>"101110000",
  524=>"001101110",
  525=>"101001000",
  526=>"000000100",
  527=>"001111000",
  528=>"010110111",
  529=>"001100111",
  530=>"000000111",
  531=>"100101100",
  532=>"010111101",
  533=>"001001010",
  534=>"111001000",
  535=>"000101001",
  536=>"010000001",
  537=>"000100111",
  538=>"000000101",
  539=>"100010001",
  540=>"000000101",
  541=>"001011000",
  542=>"011000011",
  543=>"010101000",
  544=>"000010111",
  545=>"100010111",
  546=>"100101001",
  547=>"110010011",
  548=>"110101000",
  549=>"001100111",
  550=>"101010000",
  551=>"011110000",
  552=>"101011001",
  553=>"001111111",
  554=>"011001000",
  555=>"101000100",
  556=>"100101110",
  557=>"000000110",
  558=>"100111111",
  559=>"111110100",
  560=>"010101101",
  561=>"001011110",
  562=>"000100100",
  563=>"110000111",
  564=>"110010100",
  565=>"111010110",
  566=>"010010100",
  567=>"010111101",
  568=>"010011011",
  569=>"101101111",
  570=>"001001010",
  571=>"010010001",
  572=>"010111010",
  573=>"000000011",
  574=>"111100100",
  575=>"111110110",
  576=>"111110010",
  577=>"010000100",
  578=>"101000111",
  579=>"110101001",
  580=>"000110011",
  581=>"000100001",
  582=>"111110101",
  583=>"111111110",
  584=>"010110100",
  585=>"000110011",
  586=>"001010100",
  587=>"100101101",
  588=>"110011111",
  589=>"010100100",
  590=>"011101110",
  591=>"100010011",
  592=>"000010010",
  593=>"110110001",
  594=>"000100100",
  595=>"110101011",
  596=>"100011111",
  597=>"111110000",
  598=>"101011111",
  599=>"000110100",
  600=>"111110101",
  601=>"000000000",
  602=>"111101000",
  603=>"000100100",
  604=>"110010101",
  605=>"001001110",
  606=>"111000110",
  607=>"110110000",
  608=>"100101001",
  609=>"000000000",
  610=>"000110011",
  611=>"001000111",
  612=>"001011111",
  613=>"010101100",
  614=>"100000011",
  615=>"100010011",
  616=>"010010101",
  617=>"101101010",
  618=>"101000001",
  619=>"101000100",
  620=>"001011010",
  621=>"011110110",
  622=>"101110001",
  623=>"101010101",
  624=>"000110101",
  625=>"101011111",
  626=>"110011010",
  627=>"001110000",
  628=>"100110010",
  629=>"000000001",
  630=>"011110000",
  631=>"110010100",
  632=>"010100100",
  633=>"110110111",
  634=>"110110111",
  635=>"010110011",
  636=>"001001001",
  637=>"011101100",
  638=>"110111011",
  639=>"101100101",
  640=>"100110101",
  641=>"100001001",
  642=>"100110111",
  643=>"001010111",
  644=>"001110010",
  645=>"100010111",
  646=>"010001100",
  647=>"101001000",
  648=>"000101111",
  649=>"000010011",
  650=>"010000111",
  651=>"101100110",
  652=>"011010000",
  653=>"010110110",
  654=>"011101111",
  655=>"011000000",
  656=>"010011100",
  657=>"100101101",
  658=>"101001001",
  659=>"100111111",
  660=>"110011011",
  661=>"011001010",
  662=>"110101111",
  663=>"110001010",
  664=>"111010000",
  665=>"001010111",
  666=>"011000111",
  667=>"110101101",
  668=>"111010011",
  669=>"111000100",
  670=>"000110110",
  671=>"001000000",
  672=>"110001011",
  673=>"000000100",
  674=>"111011100",
  675=>"001011100",
  676=>"110110100",
  677=>"111010111",
  678=>"110011000",
  679=>"111000010",
  680=>"111010000",
  681=>"101100100",
  682=>"100100110",
  683=>"010111011",
  684=>"101100110",
  685=>"110000000",
  686=>"001100000",
  687=>"101100110",
  688=>"101101000",
  689=>"110110110",
  690=>"110111111",
  691=>"100110110",
  692=>"100110010",
  693=>"111000000",
  694=>"111111011",
  695=>"111111011",
  696=>"110111010",
  697=>"100100111",
  698=>"011010110",
  699=>"101001101",
  700=>"100111111",
  701=>"100100000",
  702=>"101111100",
  703=>"001111011",
  704=>"100100001",
  705=>"110010110",
  706=>"100000100",
  707=>"000011010",
  708=>"110110111",
  709=>"010001100",
  710=>"000110110",
  711=>"011111010",
  712=>"010011100",
  713=>"011110100",
  714=>"011010100",
  715=>"001000010",
  716=>"000011001",
  717=>"100111111",
  718=>"110000100",
  719=>"001010100",
  720=>"011001010",
  721=>"100101100",
  722=>"000001011",
  723=>"001000110",
  724=>"100010011",
  725=>"001010111",
  726=>"100001111",
  727=>"100000111",
  728=>"100111010",
  729=>"110110010",
  730=>"110001011",
  731=>"101001000",
  732=>"110000000",
  733=>"011100011",
  734=>"001011101",
  735=>"111110111",
  736=>"011110001",
  737=>"001100001",
  738=>"111101001",
  739=>"010101101",
  740=>"000110111",
  741=>"111000001",
  742=>"011011110",
  743=>"110111110",
  744=>"001111011",
  745=>"110001011",
  746=>"001010000",
  747=>"100000110",
  748=>"100001001",
  749=>"110110010",
  750=>"011101111",
  751=>"000000100",
  752=>"000100101",
  753=>"001110101",
  754=>"000001111",
  755=>"110011100",
  756=>"100111101",
  757=>"011101010",
  758=>"101100000",
  759=>"100111110",
  760=>"111010111",
  761=>"001000010",
  762=>"001111011",
  763=>"011001000",
  764=>"100110100",
  765=>"000110010",
  766=>"001000110",
  767=>"010111000",
  768=>"000000110",
  769=>"000000101",
  770=>"011110011",
  771=>"010000110",
  772=>"110011101",
  773=>"001111011",
  774=>"101000111",
  775=>"110001111",
  776=>"001110000",
  777=>"010100001",
  778=>"111011111",
  779=>"001001001",
  780=>"011011110",
  781=>"000011100",
  782=>"010001100",
  783=>"111110101",
  784=>"101000010",
  785=>"000100000",
  786=>"101001100",
  787=>"011011110",
  788=>"000111011",
  789=>"110010110",
  790=>"011111010",
  791=>"010001011",
  792=>"000010011",
  793=>"011000110",
  794=>"110111101",
  795=>"011000010",
  796=>"111101001",
  797=>"101111010",
  798=>"101111110",
  799=>"101111100",
  800=>"101100011",
  801=>"111010011",
  802=>"111111000",
  803=>"100101001",
  804=>"101111110",
  805=>"111110001",
  806=>"101011010",
  807=>"110101110",
  808=>"101001011",
  809=>"010011101",
  810=>"111100000",
  811=>"111100110",
  812=>"111001101",
  813=>"101010011",
  814=>"001010011",
  815=>"001010001",
  816=>"110011100",
  817=>"100000110",
  818=>"011000101",
  819=>"000000001",
  820=>"101111110",
  821=>"111111001",
  822=>"001110010",
  823=>"010011100",
  824=>"110111101",
  825=>"001101110",
  826=>"001011011",
  827=>"111011000",
  828=>"000000001",
  829=>"000100110",
  830=>"011111100",
  831=>"011101010",
  832=>"001100111",
  833=>"011111011",
  834=>"001001001",
  835=>"010011010",
  836=>"100010000",
  837=>"110011011",
  838=>"100000101",
  839=>"110101100",
  840=>"001100100",
  841=>"111001101",
  842=>"100111010",
  843=>"000111011",
  844=>"000101001",
  845=>"100001100",
  846=>"100001111",
  847=>"001000101",
  848=>"001000111",
  849=>"001111110",
  850=>"110110100",
  851=>"000111100",
  852=>"011101111",
  853=>"111101101",
  854=>"100000000",
  855=>"110000010",
  856=>"010111011",
  857=>"001001000",
  858=>"111001011",
  859=>"011111111",
  860=>"001001010",
  861=>"011011011",
  862=>"100010000",
  863=>"000110101",
  864=>"000100000",
  865=>"000101001",
  866=>"110011111",
  867=>"101111110",
  868=>"110110010",
  869=>"000101000",
  870=>"110011100",
  871=>"111111001",
  872=>"000000000",
  873=>"111001000",
  874=>"100000101",
  875=>"110001010",
  876=>"111001001",
  877=>"110110011",
  878=>"110101100",
  879=>"000000101",
  880=>"111000101",
  881=>"011100011",
  882=>"000111101",
  883=>"010101100",
  884=>"111100001",
  885=>"101100011",
  886=>"001111010",
  887=>"000100100",
  888=>"111111010",
  889=>"100011000",
  890=>"111010000",
  891=>"100011110",
  892=>"000110000",
  893=>"100001101",
  894=>"111001101",
  895=>"010000100",
  896=>"100110011",
  897=>"110111001",
  898=>"110011100",
  899=>"110111010",
  900=>"000100000",
  901=>"010011001",
  902=>"010110111",
  903=>"110001110",
  904=>"101100100",
  905=>"110011100",
  906=>"110001111",
  907=>"011111001",
  908=>"000111100",
  909=>"100000011",
  910=>"000110111",
  911=>"110100100",
  912=>"100111101",
  913=>"111111011",
  914=>"000010000",
  915=>"110101110",
  916=>"000001101",
  917=>"100111010",
  918=>"000110000",
  919=>"101010111",
  920=>"111011011",
  921=>"110110110",
  922=>"010110011",
  923=>"101001000",
  924=>"011101111",
  925=>"010010101",
  926=>"010101110",
  927=>"000000000",
  928=>"100000010",
  929=>"100010100",
  930=>"100100011",
  931=>"001100011",
  932=>"010000111",
  933=>"110100001",
  934=>"110101101",
  935=>"001110100",
  936=>"000010010",
  937=>"110000000",
  938=>"001010110",
  939=>"000010100",
  940=>"001000001",
  941=>"110101100",
  942=>"101101011",
  943=>"100101101",
  944=>"000111001",
  945=>"010100101",
  946=>"010000111",
  947=>"110110100",
  948=>"011010011",
  949=>"110010000",
  950=>"100111001",
  951=>"001000010",
  952=>"001010100",
  953=>"101101001",
  954=>"100000011",
  955=>"001101011",
  956=>"001000101",
  957=>"100000101",
  958=>"101111000",
  959=>"110110001",
  960=>"001100000",
  961=>"100100110",
  962=>"111011001",
  963=>"111010000",
  964=>"011111010",
  965=>"011101001",
  966=>"100001010",
  967=>"110110111",
  968=>"010101110",
  969=>"010011011",
  970=>"101111111",
  971=>"101111011",
  972=>"101000010",
  973=>"010010100",
  974=>"101110000",
  975=>"001000100",
  976=>"010000000",
  977=>"000110100",
  978=>"000010011",
  979=>"001111001",
  980=>"001100011",
  981=>"010111001",
  982=>"111000010",
  983=>"000100111",
  984=>"110100100",
  985=>"100000110",
  986=>"000000011",
  987=>"101000101",
  988=>"010001111",
  989=>"001011111",
  990=>"110011101",
  991=>"010011000",
  992=>"001000111",
  993=>"010100011",
  994=>"011111001",
  995=>"001000110",
  996=>"100100100",
  997=>"010011011",
  998=>"111110101",
  999=>"100100011",
  1000=>"100101111",
  1001=>"110011001",
  1002=>"010000010",
  1003=>"101010011",
  1004=>"111011011",
  1005=>"000011001",
  1006=>"001001011",
  1007=>"001010111",
  1008=>"011101101",
  1009=>"101010000",
  1010=>"000110100",
  1011=>"111111111",
  1012=>"111000010",
  1013=>"000101000",
  1014=>"110110010",
  1015=>"100011000",
  1016=>"001110010",
  1017=>"110000100",
  1018=>"001000110",
  1019=>"000001010",
  1020=>"100110111",
  1021=>"111010101",
  1022=>"011010100",
  1023=>"111001010",
  1024=>"000101101",
  1025=>"101100000",
  1026=>"100011100",
  1027=>"101000011",
  1028=>"101011101",
  1029=>"110110010",
  1030=>"001000000",
  1031=>"001101100",
  1032=>"000010111",
  1033=>"000001001",
  1034=>"110111111",
  1035=>"000000011",
  1036=>"001001111",
  1037=>"000011000",
  1038=>"111000000",
  1039=>"000010011",
  1040=>"110110011",
  1041=>"110111111",
  1042=>"000111110",
  1043=>"010111111",
  1044=>"110110101",
  1045=>"000001100",
  1046=>"001101110",
  1047=>"110110101",
  1048=>"010101110",
  1049=>"000010100",
  1050=>"100001000",
  1051=>"101010011",
  1052=>"101001001",
  1053=>"101110000",
  1054=>"111010101",
  1055=>"100100000",
  1056=>"011110101",
  1057=>"101100110",
  1058=>"100001110",
  1059=>"011110010",
  1060=>"111000001",
  1061=>"110011111",
  1062=>"011110000",
  1063=>"110011001",
  1064=>"000000001",
  1065=>"111000111",
  1066=>"000101100",
  1067=>"111111110",
  1068=>"100001010",
  1069=>"010010100",
  1070=>"001100011",
  1071=>"001011010",
  1072=>"010000010",
  1073=>"001011101",
  1074=>"000001101",
  1075=>"100111110",
  1076=>"110101100",
  1077=>"100100010",
  1078=>"101100101",
  1079=>"110111100",
  1080=>"010011110",
  1081=>"011110001",
  1082=>"000000001",
  1083=>"010101010",
  1084=>"101001011",
  1085=>"000110101",
  1086=>"111111001",
  1087=>"010111111",
  1088=>"001000101",
  1089=>"001110100",
  1090=>"101001100",
  1091=>"010000111",
  1092=>"110110110",
  1093=>"001111100",
  1094=>"000100001",
  1095=>"110011101",
  1096=>"100111101",
  1097=>"001011110",
  1098=>"101010101",
  1099=>"110000001",
  1100=>"100000011",
  1101=>"101000000",
  1102=>"110101100",
  1103=>"011101100",
  1104=>"001100110",
  1105=>"110000011",
  1106=>"001101000",
  1107=>"000001011",
  1108=>"000001101",
  1109=>"101011100",
  1110=>"111111101",
  1111=>"100100110",
  1112=>"111110011",
  1113=>"110001111",
  1114=>"111011010",
  1115=>"000011100",
  1116=>"100000101",
  1117=>"101011110",
  1118=>"101001001",
  1119=>"011001101",
  1120=>"010010011",
  1121=>"101111101",
  1122=>"100011101",
  1123=>"000001000",
  1124=>"011000100",
  1125=>"110001101",
  1126=>"111101110",
  1127=>"111100101",
  1128=>"010011101",
  1129=>"010110001",
  1130=>"010001101",
  1131=>"001001000",
  1132=>"111100010",
  1133=>"000101010",
  1134=>"100110011",
  1135=>"010111010",
  1136=>"111100111",
  1137=>"110110000",
  1138=>"111100010",
  1139=>"001010000",
  1140=>"100000010",
  1141=>"100110001",
  1142=>"111001110",
  1143=>"011101011",
  1144=>"010001100",
  1145=>"111010111",
  1146=>"010111100",
  1147=>"011010101",
  1148=>"010111100",
  1149=>"101110100",
  1150=>"101011110",
  1151=>"011011001",
  1152=>"000000011",
  1153=>"111001000",
  1154=>"101011001",
  1155=>"100000010",
  1156=>"111100000",
  1157=>"010011010",
  1158=>"110001111",
  1159=>"100000001",
  1160=>"111010101",
  1161=>"100100010",
  1162=>"100001101",
  1163=>"111001100",
  1164=>"110100010",
  1165=>"010111011",
  1166=>"011000000",
  1167=>"111011000",
  1168=>"011010011",
  1169=>"110110010",
  1170=>"110011001",
  1171=>"101100011",
  1172=>"010011101",
  1173=>"110101011",
  1174=>"011101101",
  1175=>"100100001",
  1176=>"100011010",
  1177=>"001101000",
  1178=>"000111011",
  1179=>"010010010",
  1180=>"000011001",
  1181=>"110010010",
  1182=>"111101110",
  1183=>"010010100",
  1184=>"000000101",
  1185=>"100000001",
  1186=>"111111001",
  1187=>"101110110",
  1188=>"001100011",
  1189=>"111001001",
  1190=>"000110101",
  1191=>"001100101",
  1192=>"111101011",
  1193=>"111110111",
  1194=>"111111100",
  1195=>"110011010",
  1196=>"001000010",
  1197=>"000101101",
  1198=>"111100101",
  1199=>"100111001",
  1200=>"101001000",
  1201=>"011110000",
  1202=>"101110000",
  1203=>"100100001",
  1204=>"011101010",
  1205=>"100000111",
  1206=>"000010011",
  1207=>"100110000",
  1208=>"010001100",
  1209=>"101100101",
  1210=>"001010001",
  1211=>"110101000",
  1212=>"110011000",
  1213=>"000010110",
  1214=>"101111101",
  1215=>"111001100",
  1216=>"101001000",
  1217=>"000100011",
  1218=>"111100000",
  1219=>"001100001",
  1220=>"011110110",
  1221=>"011111001",
  1222=>"110101111",
  1223=>"101010000",
  1224=>"001010000",
  1225=>"101101110",
  1226=>"001010111",
  1227=>"110101110",
  1228=>"000100110",
  1229=>"010000001",
  1230=>"101011111",
  1231=>"111011001",
  1232=>"010100111",
  1233=>"000010110",
  1234=>"001001000",
  1235=>"011101111",
  1236=>"011111110",
  1237=>"110001010",
  1238=>"101100101",
  1239=>"010000111",
  1240=>"111010011",
  1241=>"011101010",
  1242=>"110000010",
  1243=>"110100001",
  1244=>"011010101",
  1245=>"100001000",
  1246=>"111010101",
  1247=>"101111000",
  1248=>"011010011",
  1249=>"001001011",
  1250=>"001001011",
  1251=>"010100000",
  1252=>"110111001",
  1253=>"101110110",
  1254=>"010110010",
  1255=>"111011101",
  1256=>"111101011",
  1257=>"010110111",
  1258=>"100000001",
  1259=>"010101001",
  1260=>"011100010",
  1261=>"111010100",
  1262=>"111010101",
  1263=>"000100000",
  1264=>"110000111",
  1265=>"000011101",
  1266=>"011110011",
  1267=>"000001110",
  1268=>"111110111",
  1269=>"000101001",
  1270=>"111110111",
  1271=>"110101001",
  1272=>"010001000",
  1273=>"011011011",
  1274=>"110000111",
  1275=>"001000011",
  1276=>"001110100",
  1277=>"011010000",
  1278=>"011110101",
  1279=>"011100010",
  1280=>"111010100",
  1281=>"101100101",
  1282=>"000000001",
  1283=>"011110100",
  1284=>"110010110",
  1285=>"011011111",
  1286=>"011101001",
  1287=>"011011100",
  1288=>"011000100",
  1289=>"111111110",
  1290=>"110100010",
  1291=>"000001001",
  1292=>"010001001",
  1293=>"000010110",
  1294=>"111101101",
  1295=>"100111110",
  1296=>"101001101",
  1297=>"110010100",
  1298=>"100001000",
  1299=>"110111001",
  1300=>"000100111",
  1301=>"100011100",
  1302=>"100011101",
  1303=>"001011110",
  1304=>"100011110",
  1305=>"011000001",
  1306=>"001100111",
  1307=>"111101000",
  1308=>"110001000",
  1309=>"001111101",
  1310=>"100110000",
  1311=>"110101010",
  1312=>"110011110",
  1313=>"001101001",
  1314=>"110001010",
  1315=>"011010010",
  1316=>"010011000",
  1317=>"010100010",
  1318=>"010011001",
  1319=>"111010001",
  1320=>"100100000",
  1321=>"000001111",
  1322=>"111101000",
  1323=>"100000101",
  1324=>"011110111",
  1325=>"100010001",
  1326=>"100100010",
  1327=>"111110000",
  1328=>"100011000",
  1329=>"111100100",
  1330=>"010001111",
  1331=>"000100000",
  1332=>"000101010",
  1333=>"001010011",
  1334=>"101010010",
  1335=>"110101000",
  1336=>"011100011",
  1337=>"111000010",
  1338=>"001001101",
  1339=>"100110101",
  1340=>"000000101",
  1341=>"100010110",
  1342=>"011001111",
  1343=>"011110010",
  1344=>"111011100",
  1345=>"101010001",
  1346=>"110100111",
  1347=>"100011110",
  1348=>"011111001",
  1349=>"111001101",
  1350=>"111100111",
  1351=>"101010100",
  1352=>"101001111",
  1353=>"110001010",
  1354=>"011000011",
  1355=>"000010001",
  1356=>"010001000",
  1357=>"010111000",
  1358=>"110110110",
  1359=>"000000010",
  1360=>"001000010",
  1361=>"001110101",
  1362=>"000011110",
  1363=>"001001001",
  1364=>"001000001",
  1365=>"010011100",
  1366=>"001011010",
  1367=>"101100100",
  1368=>"100100000",
  1369=>"000110000",
  1370=>"001100011",
  1371=>"101101010",
  1372=>"110100000",
  1373=>"110111111",
  1374=>"101111011",
  1375=>"101110001",
  1376=>"111110100",
  1377=>"110010001",
  1378=>"101001110",
  1379=>"101000010",
  1380=>"111000000",
  1381=>"010010010",
  1382=>"110001110",
  1383=>"000111001",
  1384=>"100011010",
  1385=>"101101100",
  1386=>"001000010",
  1387=>"000010001",
  1388=>"101001111",
  1389=>"100110100",
  1390=>"101111111",
  1391=>"000010101",
  1392=>"010001000",
  1393=>"111111101",
  1394=>"101101110",
  1395=>"011101011",
  1396=>"000001110",
  1397=>"111100011",
  1398=>"110010101",
  1399=>"011010000",
  1400=>"000001011",
  1401=>"011110011",
  1402=>"010011101",
  1403=>"100100111",
  1404=>"010011010",
  1405=>"011100001",
  1406=>"111100110",
  1407=>"010110000",
  1408=>"101100100",
  1409=>"000100100",
  1410=>"110011011",
  1411=>"110110011",
  1412=>"110001110",
  1413=>"110101001",
  1414=>"000100010",
  1415=>"101011111",
  1416=>"111110110",
  1417=>"010011011",
  1418=>"111101111",
  1419=>"000110100",
  1420=>"011101100",
  1421=>"010010011",
  1422=>"100010011",
  1423=>"111100001",
  1424=>"000110101",
  1425=>"010101110",
  1426=>"011001000",
  1427=>"110011100",
  1428=>"110010100",
  1429=>"001101000",
  1430=>"000011100",
  1431=>"000010001",
  1432=>"010100101",
  1433=>"011000010",
  1434=>"010011000",
  1435=>"010010101",
  1436=>"111000001",
  1437=>"010010010",
  1438=>"101010001",
  1439=>"110110000",
  1440=>"110010001",
  1441=>"001100001",
  1442=>"010011100",
  1443=>"111100011",
  1444=>"010100110",
  1445=>"101110101",
  1446=>"110111001",
  1447=>"010010010",
  1448=>"100001110",
  1449=>"111111110",
  1450=>"000001101",
  1451=>"000001101",
  1452=>"111110000",
  1453=>"110100001",
  1454=>"000000011",
  1455=>"011101010",
  1456=>"101000110",
  1457=>"001010010",
  1458=>"110101001",
  1459=>"111100000",
  1460=>"110100001",
  1461=>"100110100",
  1462=>"111100000",
  1463=>"010100000",
  1464=>"100110010",
  1465=>"011100011",
  1466=>"000111111",
  1467=>"111100100",
  1468=>"000001001",
  1469=>"011011000",
  1470=>"010001100",
  1471=>"000000111",
  1472=>"011001011",
  1473=>"111001000",
  1474=>"001001110",
  1475=>"111001110",
  1476=>"011101011",
  1477=>"011111000",
  1478=>"010001011",
  1479=>"000000010",
  1480=>"110100010",
  1481=>"000101110",
  1482=>"100101111",
  1483=>"111010101",
  1484=>"111100001",
  1485=>"010000111",
  1486=>"010010101",
  1487=>"111001100",
  1488=>"000100011",
  1489=>"001111011",
  1490=>"011111100",
  1491=>"110101010",
  1492=>"111100001",
  1493=>"001111100",
  1494=>"000010010",
  1495=>"100110100",
  1496=>"010011100",
  1497=>"111101011",
  1498=>"010111010",
  1499=>"011010110",
  1500=>"110100001",
  1501=>"111111110",
  1502=>"000111001",
  1503=>"100010110",
  1504=>"001111100",
  1505=>"011010111",
  1506=>"101001010",
  1507=>"100000101",
  1508=>"010110000",
  1509=>"011101100",
  1510=>"111001001",
  1511=>"101111100",
  1512=>"010011111",
  1513=>"101110110",
  1514=>"000101110",
  1515=>"011010111",
  1516=>"111001000",
  1517=>"110010010",
  1518=>"100111100",
  1519=>"110111010",
  1520=>"101011000",
  1521=>"100100100",
  1522=>"100000001",
  1523=>"101100101",
  1524=>"110100101",
  1525=>"000110000",
  1526=>"101111011",
  1527=>"000010001",
  1528=>"110101011",
  1529=>"001110111",
  1530=>"011000111",
  1531=>"101100110",
  1532=>"000100000",
  1533=>"011001110",
  1534=>"101100001",
  1535=>"111111111",
  1536=>"000010010",
  1537=>"101100100",
  1538=>"001110000",
  1539=>"101100010",
  1540=>"001010010",
  1541=>"010101110",
  1542=>"101000100",
  1543=>"000000010",
  1544=>"010100100",
  1545=>"110101100",
  1546=>"110011001",
  1547=>"101111001",
  1548=>"011100101",
  1549=>"100111110",
  1550=>"101110011",
  1551=>"101111101",
  1552=>"100110110",
  1553=>"111100100",
  1554=>"110000011",
  1555=>"101100110",
  1556=>"001010010",
  1557=>"111101110",
  1558=>"010100100",
  1559=>"000001110",
  1560=>"101111100",
  1561=>"001001000",
  1562=>"100001000",
  1563=>"101011100",
  1564=>"011001000",
  1565=>"010010110",
  1566=>"001101000",
  1567=>"011100010",
  1568=>"101001010",
  1569=>"110001111",
  1570=>"101001110",
  1571=>"011110010",
  1572=>"100111010",
  1573=>"110110111",
  1574=>"001110110",
  1575=>"110010111",
  1576=>"001001011",
  1577=>"101111001",
  1578=>"100111101",
  1579=>"011011111",
  1580=>"001000011",
  1581=>"010000101",
  1582=>"100000001",
  1583=>"100110000",
  1584=>"100001110",
  1585=>"111111100",
  1586=>"001000010",
  1587=>"100111100",
  1588=>"110011101",
  1589=>"111001000",
  1590=>"010000100",
  1591=>"001010001",
  1592=>"000101000",
  1593=>"111110100",
  1594=>"111000100",
  1595=>"011001011",
  1596=>"001010100",
  1597=>"110010010",
  1598=>"111001101",
  1599=>"010011100",
  1600=>"100010001",
  1601=>"101001000",
  1602=>"110100110",
  1603=>"111101001",
  1604=>"111110011",
  1605=>"011001111",
  1606=>"010001000",
  1607=>"110010000",
  1608=>"101001110",
  1609=>"001001111",
  1610=>"110110101",
  1611=>"011000001",
  1612=>"101110110",
  1613=>"010010111",
  1614=>"110001111",
  1615=>"010000101",
  1616=>"101000011",
  1617=>"100110110",
  1618=>"000110111",
  1619=>"011101110",
  1620=>"101111100",
  1621=>"010101000",
  1622=>"001101111",
  1623=>"001101100",
  1624=>"101001011",
  1625=>"111111100",
  1626=>"001010011",
  1627=>"101001100",
  1628=>"010000100",
  1629=>"100101111",
  1630=>"000000000",
  1631=>"111011110",
  1632=>"010011111",
  1633=>"100011111",
  1634=>"110011011",
  1635=>"110110110",
  1636=>"111100010",
  1637=>"100101001",
  1638=>"011101000",
  1639=>"111100100",
  1640=>"100001001",
  1641=>"110111100",
  1642=>"011111111",
  1643=>"000101100",
  1644=>"001100011",
  1645=>"010011000",
  1646=>"100100111",
  1647=>"001110010",
  1648=>"010011101",
  1649=>"000010101",
  1650=>"000110001",
  1651=>"111010101",
  1652=>"110010101",
  1653=>"000100110",
  1654=>"100011101",
  1655=>"110100001",
  1656=>"110100110",
  1657=>"100010110",
  1658=>"101110101",
  1659=>"011001111",
  1660=>"011101111",
  1661=>"000111110",
  1662=>"000110101",
  1663=>"010100111",
  1664=>"000010001",
  1665=>"001010101",
  1666=>"011111011",
  1667=>"001000000",
  1668=>"110111000",
  1669=>"101100100",
  1670=>"010001111",
  1671=>"011001100",
  1672=>"111110001",
  1673=>"111000001",
  1674=>"100000001",
  1675=>"101010111",
  1676=>"100001001",
  1677=>"101010110",
  1678=>"011010011",
  1679=>"110101110",
  1680=>"001111110",
  1681=>"000110011",
  1682=>"000001010",
  1683=>"000110011",
  1684=>"101000101",
  1685=>"101110110",
  1686=>"101000011",
  1687=>"100001111",
  1688=>"001010101",
  1689=>"101010000",
  1690=>"000000101",
  1691=>"101110110",
  1692=>"000001011",
  1693=>"011010110",
  1694=>"000010010",
  1695=>"101110000",
  1696=>"000101010",
  1697=>"100101001",
  1698=>"100100010",
  1699=>"101001010",
  1700=>"010101011",
  1701=>"111001001",
  1702=>"111001000",
  1703=>"010010000",
  1704=>"000000000",
  1705=>"100011111",
  1706=>"100110100",
  1707=>"001000000",
  1708=>"000010001",
  1709=>"111110000",
  1710=>"101101100",
  1711=>"101011001",
  1712=>"001001000",
  1713=>"110101110",
  1714=>"101101001",
  1715=>"111000010",
  1716=>"110011111",
  1717=>"001110010",
  1718=>"011010101",
  1719=>"110010011",
  1720=>"000100000",
  1721=>"101111110",
  1722=>"111010111",
  1723=>"101100110",
  1724=>"001101111",
  1725=>"000101010",
  1726=>"001000110",
  1727=>"110000111",
  1728=>"100001000",
  1729=>"010100001",
  1730=>"101101111",
  1731=>"000100010",
  1732=>"010011011",
  1733=>"000000111",
  1734=>"110001000",
  1735=>"001010000",
  1736=>"101100110",
  1737=>"010000000",
  1738=>"010011010",
  1739=>"101000110",
  1740=>"011001101",
  1741=>"110100010",
  1742=>"110100010",
  1743=>"110110111",
  1744=>"001101110",
  1745=>"010011001",
  1746=>"110001010",
  1747=>"110111001",
  1748=>"000110110",
  1749=>"001011111",
  1750=>"011000011",
  1751=>"010100011",
  1752=>"101011110",
  1753=>"000001110",
  1754=>"011001011",
  1755=>"101010111",
  1756=>"000100101",
  1757=>"110101000",
  1758=>"001011101",
  1759=>"100011101",
  1760=>"001111110",
  1761=>"110101101",
  1762=>"110010111",
  1763=>"110110111",
  1764=>"110100101",
  1765=>"111111110",
  1766=>"010000000",
  1767=>"111100111",
  1768=>"001001100",
  1769=>"110000000",
  1770=>"011000010",
  1771=>"111000001",
  1772=>"101011110",
  1773=>"101011101",
  1774=>"011001001",
  1775=>"000000010",
  1776=>"010000010",
  1777=>"111100000",
  1778=>"110101010",
  1779=>"100111000",
  1780=>"100110010",
  1781=>"111110111",
  1782=>"110010001",
  1783=>"111001001",
  1784=>"000010000",
  1785=>"010111110",
  1786=>"001110001",
  1787=>"011000011",
  1788=>"111001011",
  1789=>"010010000",
  1790=>"110110010",
  1791=>"101001001",
  1792=>"100000111",
  1793=>"000001011",
  1794=>"001010101",
  1795=>"001111000",
  1796=>"100000110",
  1797=>"111011000",
  1798=>"110001100",
  1799=>"101000000",
  1800=>"100010001",
  1801=>"010110010",
  1802=>"111010000",
  1803=>"001010110",
  1804=>"101101100",
  1805=>"100010101",
  1806=>"101000110",
  1807=>"000010110",
  1808=>"000011111",
  1809=>"111101100",
  1810=>"000001000",
  1811=>"101101011",
  1812=>"111010010",
  1813=>"001001010",
  1814=>"100001011",
  1815=>"001111101",
  1816=>"101000100",
  1817=>"101000100",
  1818=>"111001001",
  1819=>"101010000",
  1820=>"100111101",
  1821=>"011000001",
  1822=>"010000100",
  1823=>"100010010",
  1824=>"010100010",
  1825=>"101000000",
  1826=>"101100110",
  1827=>"001010101",
  1828=>"110000011",
  1829=>"010111100",
  1830=>"110011110",
  1831=>"111100111",
  1832=>"010110011",
  1833=>"000001100",
  1834=>"010010100",
  1835=>"001100100",
  1836=>"101100110",
  1837=>"111000110",
  1838=>"001011000",
  1839=>"100101111",
  1840=>"111000110",
  1841=>"011010000",
  1842=>"110101101",
  1843=>"001000101",
  1844=>"101001011",
  1845=>"110111000",
  1846=>"000010110",
  1847=>"011101110",
  1848=>"101011110",
  1849=>"001100110",
  1850=>"101100000",
  1851=>"110000111",
  1852=>"100010101",
  1853=>"001000000",
  1854=>"001000001",
  1855=>"000111111",
  1856=>"111011010",
  1857=>"011101000",
  1858=>"010010100",
  1859=>"111111110",
  1860=>"001001100",
  1861=>"101111011",
  1862=>"001011010",
  1863=>"110100101",
  1864=>"100110111",
  1865=>"110001000",
  1866=>"101101011",
  1867=>"110000110",
  1868=>"011101011",
  1869=>"000101000",
  1870=>"000011101",
  1871=>"111010010",
  1872=>"101011011",
  1873=>"101011101",
  1874=>"010110111",
  1875=>"111001110",
  1876=>"101000001",
  1877=>"000111010",
  1878=>"010011100",
  1879=>"100100010",
  1880=>"001000011",
  1881=>"111000000",
  1882=>"000100111",
  1883=>"011111111",
  1884=>"110010010",
  1885=>"101110100",
  1886=>"000011001",
  1887=>"101111100",
  1888=>"100110110",
  1889=>"100011010",
  1890=>"001011111",
  1891=>"111000000",
  1892=>"111110010",
  1893=>"000000000",
  1894=>"111110010",
  1895=>"001110001",
  1896=>"011011101",
  1897=>"111110000",
  1898=>"100010101",
  1899=>"010000101",
  1900=>"000001000",
  1901=>"010111101",
  1902=>"001000010",
  1903=>"011001110",
  1904=>"001101100",
  1905=>"101101110",
  1906=>"101011001",
  1907=>"111011000",
  1908=>"000110011",
  1909=>"000000000",
  1910=>"100101010",
  1911=>"001010001",
  1912=>"010101001",
  1913=>"010001011",
  1914=>"011110101",
  1915=>"110110010",
  1916=>"110100011",
  1917=>"111101111",
  1918=>"101101111",
  1919=>"110110110",
  1920=>"111001000",
  1921=>"010101011",
  1922=>"101001101",
  1923=>"100011100",
  1924=>"000000000",
  1925=>"011010101",
  1926=>"111010001",
  1927=>"110001100",
  1928=>"111000001",
  1929=>"111011011",
  1930=>"001100001",
  1931=>"110000100",
  1932=>"110100111",
  1933=>"000101000",
  1934=>"011111010",
  1935=>"001001110",
  1936=>"001100001",
  1937=>"010110011",
  1938=>"011000010",
  1939=>"010011010",
  1940=>"110011101",
  1941=>"100010101",
  1942=>"000001111",
  1943=>"000111111",
  1944=>"101000110",
  1945=>"010111110",
  1946=>"110100111",
  1947=>"111010010",
  1948=>"111110001",
  1949=>"101101111",
  1950=>"011000111",
  1951=>"101011011",
  1952=>"001010110",
  1953=>"110011010",
  1954=>"111001011",
  1955=>"111001001",
  1956=>"001110001",
  1957=>"001010011",
  1958=>"000010010",
  1959=>"011100001",
  1960=>"001110111",
  1961=>"111111111",
  1962=>"010110100",
  1963=>"111110111",
  1964=>"101101000",
  1965=>"111011110",
  1966=>"101001100",
  1967=>"111110011",
  1968=>"000011011",
  1969=>"100010101",
  1970=>"011011010",
  1971=>"110011000",
  1972=>"001010111",
  1973=>"111101011",
  1974=>"110010111",
  1975=>"000010010",
  1976=>"011011001",
  1977=>"100100010",
  1978=>"000000011",
  1979=>"111000001",
  1980=>"101100000",
  1981=>"001110001",
  1982=>"110100010",
  1983=>"101000000",
  1984=>"011001001",
  1985=>"101000110",
  1986=>"100010001",
  1987=>"010111001",
  1988=>"001111101",
  1989=>"101001011",
  1990=>"110000011",
  1991=>"001011101",
  1992=>"110110010",
  1993=>"001011001",
  1994=>"011111100",
  1995=>"110100101",
  1996=>"001001000",
  1997=>"100100101",
  1998=>"000100011",
  1999=>"111111000",
  2000=>"010000110",
  2001=>"100101100",
  2002=>"010101111",
  2003=>"001000100",
  2004=>"000001101",
  2005=>"100101110",
  2006=>"000010111",
  2007=>"000101111",
  2008=>"000010010",
  2009=>"110101101",
  2010=>"000101010",
  2011=>"001010000",
  2012=>"111010001",
  2013=>"000110001",
  2014=>"100011011",
  2015=>"001011010",
  2016=>"101111110",
  2017=>"110011011",
  2018=>"000101110",
  2019=>"010100110",
  2020=>"001010110",
  2021=>"000000000",
  2022=>"000111110",
  2023=>"100110000",
  2024=>"110000010",
  2025=>"111101101",
  2026=>"111001011",
  2027=>"101001001",
  2028=>"001011111",
  2029=>"110111011",
  2030=>"011111011",
  2031=>"100100100",
  2032=>"001100010",
  2033=>"000000100",
  2034=>"100100101",
  2035=>"001000011",
  2036=>"110110110",
  2037=>"000000101",
  2038=>"100011010",
  2039=>"001011110",
  2040=>"000000011",
  2041=>"010001000",
  2042=>"001000000",
  2043=>"101010111",
  2044=>"001010111",
  2045=>"001000001",
  2046=>"001100111",
  2047=>"100110000",
  2048=>"111100111",
  2049=>"101110000",
  2050=>"111010110",
  2051=>"011000001",
  2052=>"000011111",
  2053=>"111001011",
  2054=>"001001110",
  2055=>"011101001",
  2056=>"101001100",
  2057=>"100011010",
  2058=>"101011110",
  2059=>"001101101",
  2060=>"000110010",
  2061=>"110111101",
  2062=>"111011100",
  2063=>"000010000",
  2064=>"111101001",
  2065=>"101110110",
  2066=>"011000101",
  2067=>"011010110",
  2068=>"100000000",
  2069=>"110101101",
  2070=>"100100001",
  2071=>"000110000",
  2072=>"111000000",
  2073=>"100110110",
  2074=>"100011101",
  2075=>"110001010",
  2076=>"110000000",
  2077=>"110000110",
  2078=>"000000111",
  2079=>"010110111",
  2080=>"011101100",
  2081=>"000111000",
  2082=>"111001100",
  2083=>"010101110",
  2084=>"111011001",
  2085=>"000110100",
  2086=>"001101001",
  2087=>"111110110",
  2088=>"111001011",
  2089=>"101011111",
  2090=>"010010111",
  2091=>"100010100",
  2092=>"110001111",
  2093=>"000110111",
  2094=>"100100101",
  2095=>"001101111",
  2096=>"000001110",
  2097=>"100010100",
  2098=>"110101111",
  2099=>"011010110",
  2100=>"111001011",
  2101=>"000001110",
  2102=>"001001010",
  2103=>"000001100",
  2104=>"100101111",
  2105=>"001000011",
  2106=>"010101101",
  2107=>"100110100",
  2108=>"100111001",
  2109=>"011100010",
  2110=>"101011001",
  2111=>"011100011",
  2112=>"110110010",
  2113=>"101010000",
  2114=>"011100100",
  2115=>"001001111",
  2116=>"101010101",
  2117=>"000001101",
  2118=>"010000010",
  2119=>"010100000",
  2120=>"000001011",
  2121=>"011100111",
  2122=>"000101100",
  2123=>"100011001",
  2124=>"000101000",
  2125=>"100001101",
  2126=>"111100010",
  2127=>"100101011",
  2128=>"000110001",
  2129=>"101111111",
  2130=>"101011011",
  2131=>"101011110",
  2132=>"011111101",
  2133=>"000000100",
  2134=>"100010010",
  2135=>"101001101",
  2136=>"100100010",
  2137=>"100001111",
  2138=>"100100100",
  2139=>"111100101",
  2140=>"101000100",
  2141=>"001001001",
  2142=>"001101010",
  2143=>"100100010",
  2144=>"110010100",
  2145=>"100011000",
  2146=>"100011110",
  2147=>"110001001",
  2148=>"101101011",
  2149=>"010011111",
  2150=>"000100011",
  2151=>"010110111",
  2152=>"111100010",
  2153=>"011001001",
  2154=>"100000101",
  2155=>"110100001",
  2156=>"100110110",
  2157=>"000000000",
  2158=>"101100011",
  2159=>"001110110",
  2160=>"100111001",
  2161=>"010111101",
  2162=>"100011010",
  2163=>"101110101",
  2164=>"110111110",
  2165=>"001100001",
  2166=>"110010001",
  2167=>"110011001",
  2168=>"000111001",
  2169=>"110010111",
  2170=>"001010011",
  2171=>"011110011",
  2172=>"100111101",
  2173=>"100100001",
  2174=>"111100110",
  2175=>"100000010",
  2176=>"001101000",
  2177=>"100100000",
  2178=>"010101111",
  2179=>"001001000",
  2180=>"111101000",
  2181=>"101010101",
  2182=>"001011111",
  2183=>"010111010",
  2184=>"010010110",
  2185=>"000011110",
  2186=>"100000001",
  2187=>"110010011",
  2188=>"110101000",
  2189=>"001011010",
  2190=>"000001000",
  2191=>"010100000",
  2192=>"101100110",
  2193=>"110100001",
  2194=>"111011011",
  2195=>"011010011",
  2196=>"100010000",
  2197=>"100001000",
  2198=>"110100110",
  2199=>"111110110",
  2200=>"111000110",
  2201=>"001000010",
  2202=>"100000001",
  2203=>"011111000",
  2204=>"010100100",
  2205=>"001100111",
  2206=>"111101011",
  2207=>"111100100",
  2208=>"001101011",
  2209=>"101001011",
  2210=>"110110000",
  2211=>"101001101",
  2212=>"010011100",
  2213=>"001001010",
  2214=>"111011110",
  2215=>"111101000",
  2216=>"000011011",
  2217=>"000010011",
  2218=>"011000001",
  2219=>"001111110",
  2220=>"000000010",
  2221=>"111101110",
  2222=>"110010000",
  2223=>"111000000",
  2224=>"011011000",
  2225=>"011010000",
  2226=>"110010111",
  2227=>"010001010",
  2228=>"011010101",
  2229=>"010001000",
  2230=>"100010010",
  2231=>"001101011",
  2232=>"110111100",
  2233=>"111010101",
  2234=>"011101111",
  2235=>"010010000",
  2236=>"101011100",
  2237=>"101000111",
  2238=>"101010110",
  2239=>"101001001",
  2240=>"000010001",
  2241=>"101000101",
  2242=>"101000000",
  2243=>"011010011",
  2244=>"100100010",
  2245=>"110000010",
  2246=>"010101100",
  2247=>"000000000",
  2248=>"011100110",
  2249=>"110010000",
  2250=>"001111000",
  2251=>"110101010",
  2252=>"011110110",
  2253=>"111011011",
  2254=>"011001111",
  2255=>"101100000",
  2256=>"101111101",
  2257=>"100111110",
  2258=>"000100000",
  2259=>"111111101",
  2260=>"011000101",
  2261=>"111100100",
  2262=>"110001011",
  2263=>"011101111",
  2264=>"100111010",
  2265=>"100000010",
  2266=>"000101110",
  2267=>"010011000",
  2268=>"010011010",
  2269=>"101100100",
  2270=>"110011010",
  2271=>"111000001",
  2272=>"001011000",
  2273=>"000000001",
  2274=>"010010110",
  2275=>"100001010",
  2276=>"110001000",
  2277=>"011001110",
  2278=>"000100100",
  2279=>"011011011",
  2280=>"000010110",
  2281=>"001000110",
  2282=>"011000100",
  2283=>"101100001",
  2284=>"011111101",
  2285=>"111110011",
  2286=>"000001001",
  2287=>"000001000",
  2288=>"011111100",
  2289=>"010011000",
  2290=>"100010100",
  2291=>"100100001",
  2292=>"010001001",
  2293=>"000100110",
  2294=>"010011111",
  2295=>"110000100",
  2296=>"001001110",
  2297=>"110111011",
  2298=>"100100110",
  2299=>"101011100",
  2300=>"111000000",
  2301=>"100001111",
  2302=>"001101111",
  2303=>"001000001",
  2304=>"110101011",
  2305=>"101100110",
  2306=>"101000000",
  2307=>"111100101",
  2308=>"100111110",
  2309=>"100100110",
  2310=>"001111101",
  2311=>"000101010",
  2312=>"000011010",
  2313=>"110000001",
  2314=>"010000010",
  2315=>"100101001",
  2316=>"010110111",
  2317=>"001111111",
  2318=>"011111111",
  2319=>"010010101",
  2320=>"001001000",
  2321=>"010111001",
  2322=>"000111000",
  2323=>"001010110",
  2324=>"101000000",
  2325=>"001110110",
  2326=>"110010110",
  2327=>"111010110",
  2328=>"010101110",
  2329=>"111001000",
  2330=>"100110101",
  2331=>"111101011",
  2332=>"100010010",
  2333=>"101111101",
  2334=>"001001101",
  2335=>"100001010",
  2336=>"000110101",
  2337=>"000001101",
  2338=>"010010111",
  2339=>"000100010",
  2340=>"001011101",
  2341=>"011001100",
  2342=>"010100000",
  2343=>"100101111",
  2344=>"001111101",
  2345=>"000100110",
  2346=>"011111000",
  2347=>"111000001",
  2348=>"110101111",
  2349=>"000010011",
  2350=>"100000010",
  2351=>"110010100",
  2352=>"101001110",
  2353=>"111110111",
  2354=>"000100010",
  2355=>"000001011",
  2356=>"101000000",
  2357=>"011000100",
  2358=>"000001100",
  2359=>"011000000",
  2360=>"001001000",
  2361=>"000100001",
  2362=>"100111110",
  2363=>"011110010",
  2364=>"101111010",
  2365=>"111110111",
  2366=>"111111010",
  2367=>"101010110",
  2368=>"111101100",
  2369=>"111000001",
  2370=>"111101111",
  2371=>"000000000",
  2372=>"100010111",
  2373=>"011111110",
  2374=>"101010011",
  2375=>"010110000",
  2376=>"001100000",
  2377=>"001010100",
  2378=>"000110111",
  2379=>"110010111",
  2380=>"001001001",
  2381=>"000000110",
  2382=>"110111011",
  2383=>"100110011",
  2384=>"001001001",
  2385=>"111000010",
  2386=>"011100011",
  2387=>"101011110",
  2388=>"000010000",
  2389=>"100110011",
  2390=>"101111011",
  2391=>"010001111",
  2392=>"000100001",
  2393=>"001101011",
  2394=>"010110000",
  2395=>"100001000",
  2396=>"000001001",
  2397=>"100110100",
  2398=>"011011000",
  2399=>"000111101",
  2400=>"100101010",
  2401=>"111101010",
  2402=>"101101101",
  2403=>"000010001",
  2404=>"111111000",
  2405=>"100010101",
  2406=>"110100110",
  2407=>"000100001",
  2408=>"011100111",
  2409=>"001111000",
  2410=>"011110110",
  2411=>"100001110",
  2412=>"111010011",
  2413=>"100110110",
  2414=>"001111100",
  2415=>"110011100",
  2416=>"111101001",
  2417=>"000010000",
  2418=>"001001000",
  2419=>"001101011",
  2420=>"000101110",
  2421=>"010111001",
  2422=>"101010010",
  2423=>"110110100",
  2424=>"011101000",
  2425=>"100001010",
  2426=>"010101110",
  2427=>"110010000",
  2428=>"100001000",
  2429=>"011010100",
  2430=>"010000010",
  2431=>"111100010",
  2432=>"111000101",
  2433=>"100000010",
  2434=>"100011000",
  2435=>"001001100",
  2436=>"111111000",
  2437=>"001101110",
  2438=>"111011100",
  2439=>"111011101",
  2440=>"100101100",
  2441=>"100001111",
  2442=>"111001100",
  2443=>"101000001",
  2444=>"011110110",
  2445=>"111000000",
  2446=>"001110010",
  2447=>"111110100",
  2448=>"100011101",
  2449=>"011001000",
  2450=>"010101010",
  2451=>"011111111",
  2452=>"010010000",
  2453=>"010001111",
  2454=>"011101010",
  2455=>"011000000",
  2456=>"010010000",
  2457=>"100110100",
  2458=>"110010111",
  2459=>"100100000",
  2460=>"101101101",
  2461=>"010011011",
  2462=>"101100100",
  2463=>"010010111",
  2464=>"111111100",
  2465=>"001010100",
  2466=>"100101001",
  2467=>"000111001",
  2468=>"001010110",
  2469=>"000001101",
  2470=>"000010000",
  2471=>"101001100",
  2472=>"000001111",
  2473=>"010000000",
  2474=>"011101100",
  2475=>"111001000",
  2476=>"000000111",
  2477=>"010000000",
  2478=>"010010100",
  2479=>"011100111",
  2480=>"000000111",
  2481=>"101101000",
  2482=>"010100110",
  2483=>"000111010",
  2484=>"100000010",
  2485=>"110100110",
  2486=>"110010011",
  2487=>"111110110",
  2488=>"001011111",
  2489=>"001001000",
  2490=>"001001100",
  2491=>"000000000",
  2492=>"111110010",
  2493=>"001000010",
  2494=>"110011001",
  2495=>"101111110",
  2496=>"000110011",
  2497=>"000100000",
  2498=>"110100010",
  2499=>"101100111",
  2500=>"101100010",
  2501=>"010110000",
  2502=>"110101111",
  2503=>"111001100",
  2504=>"001001101",
  2505=>"111001011",
  2506=>"111010001",
  2507=>"001001001",
  2508=>"001110100",
  2509=>"000111101",
  2510=>"101010010",
  2511=>"000101011",
  2512=>"100111110",
  2513=>"100111100",
  2514=>"100111001",
  2515=>"101010011",
  2516=>"100001110",
  2517=>"010100001",
  2518=>"001110110",
  2519=>"101100110",
  2520=>"000001010",
  2521=>"100000000",
  2522=>"110111001",
  2523=>"101011101",
  2524=>"010010000",
  2525=>"100001101",
  2526=>"111100101",
  2527=>"010100111",
  2528=>"001001101",
  2529=>"001000001",
  2530=>"110001010",
  2531=>"111001011",
  2532=>"101010011",
  2533=>"110001010",
  2534=>"011011111",
  2535=>"100010001",
  2536=>"001001100",
  2537=>"000110111",
  2538=>"111101101",
  2539=>"001100111",
  2540=>"011110001",
  2541=>"101111101",
  2542=>"111010011",
  2543=>"111101110",
  2544=>"101111011",
  2545=>"100010010",
  2546=>"001011011",
  2547=>"101101010",
  2548=>"000010101",
  2549=>"101110101",
  2550=>"001011111",
  2551=>"100000000",
  2552=>"000111010",
  2553=>"110110110",
  2554=>"101011101",
  2555=>"100110000",
  2556=>"011001000",
  2557=>"111100000",
  2558=>"010001010",
  2559=>"111110110",
  2560=>"001000000",
  2561=>"111001101",
  2562=>"000110000",
  2563=>"010001011",
  2564=>"000101001",
  2565=>"100001101",
  2566=>"101011101",
  2567=>"100111101",
  2568=>"010000111",
  2569=>"011100111",
  2570=>"001000111",
  2571=>"101010110",
  2572=>"100001001",
  2573=>"011000010",
  2574=>"011101010",
  2575=>"011110110",
  2576=>"010101001",
  2577=>"101000101",
  2578=>"100110100",
  2579=>"111001110",
  2580=>"000000000",
  2581=>"001000100",
  2582=>"110000000",
  2583=>"110011111",
  2584=>"110001011",
  2585=>"001000100",
  2586=>"101000001",
  2587=>"011111010",
  2588=>"111100001",
  2589=>"101100101",
  2590=>"100100101",
  2591=>"101101011",
  2592=>"100010111",
  2593=>"000110110",
  2594=>"101100000",
  2595=>"010000000",
  2596=>"101110100",
  2597=>"001101000",
  2598=>"001110010",
  2599=>"111111100",
  2600=>"100101000",
  2601=>"010110000",
  2602=>"001001110",
  2603=>"101111000",
  2604=>"011011100",
  2605=>"001010000",
  2606=>"011100001",
  2607=>"001000010",
  2608=>"000011100",
  2609=>"000000011",
  2610=>"001101100",
  2611=>"100100000",
  2612=>"011000101",
  2613=>"010111010",
  2614=>"010100111",
  2615=>"101100011",
  2616=>"010111010",
  2617=>"000101100",
  2618=>"111100010",
  2619=>"001000000",
  2620=>"111011010",
  2621=>"010011001",
  2622=>"011111010",
  2623=>"100111010",
  2624=>"100100001",
  2625=>"101100010",
  2626=>"110000100",
  2627=>"110010100",
  2628=>"101000100",
  2629=>"110100011",
  2630=>"100001100",
  2631=>"110000000",
  2632=>"001100001",
  2633=>"000011010",
  2634=>"101110001",
  2635=>"110000110",
  2636=>"111001100",
  2637=>"101100001",
  2638=>"101110100",
  2639=>"011001011",
  2640=>"000010001",
  2641=>"010010110",
  2642=>"100000101",
  2643=>"100010100",
  2644=>"011001011",
  2645=>"111111111",
  2646=>"001100010",
  2647=>"111110000",
  2648=>"000101011",
  2649=>"111110011",
  2650=>"010001101",
  2651=>"001110100",
  2652=>"111111101",
  2653=>"001110101",
  2654=>"101100011",
  2655=>"100110111",
  2656=>"011010100",
  2657=>"000010001",
  2658=>"110001111",
  2659=>"000100111",
  2660=>"000000010",
  2661=>"111010100",
  2662=>"101001100",
  2663=>"000100101",
  2664=>"000010011",
  2665=>"110101011",
  2666=>"010110110",
  2667=>"010110110",
  2668=>"000010100",
  2669=>"000101011",
  2670=>"011010101",
  2671=>"011110000",
  2672=>"011111011",
  2673=>"011100011",
  2674=>"000010101",
  2675=>"101100000",
  2676=>"000010100",
  2677=>"010111010",
  2678=>"000000001",
  2679=>"100010011",
  2680=>"110011111",
  2681=>"010000111",
  2682=>"011001010",
  2683=>"100101110",
  2684=>"001000001",
  2685=>"000010111",
  2686=>"000101101",
  2687=>"000110011",
  2688=>"100111010",
  2689=>"010101010",
  2690=>"110110110",
  2691=>"001010011",
  2692=>"111000000",
  2693=>"000001001",
  2694=>"100101101",
  2695=>"100110101",
  2696=>"001111010",
  2697=>"001100111",
  2698=>"011110100",
  2699=>"110011100",
  2700=>"111101101",
  2701=>"111101011",
  2702=>"100101001",
  2703=>"100001100",
  2704=>"110100111",
  2705=>"000011001",
  2706=>"000100111",
  2707=>"001100001",
  2708=>"000011000",
  2709=>"100011110",
  2710=>"101010100",
  2711=>"000010100",
  2712=>"010111010",
  2713=>"001000101",
  2714=>"101000100",
  2715=>"100001000",
  2716=>"010110011",
  2717=>"111010010",
  2718=>"010010011",
  2719=>"001000001",
  2720=>"011100001",
  2721=>"101000010",
  2722=>"111000011",
  2723=>"001000010",
  2724=>"111000000",
  2725=>"110101010",
  2726=>"101110110",
  2727=>"000001010",
  2728=>"011111100",
  2729=>"110100111",
  2730=>"100010100",
  2731=>"111101011",
  2732=>"011011010",
  2733=>"001000100",
  2734=>"001010010",
  2735=>"000000001",
  2736=>"000000001",
  2737=>"110110000",
  2738=>"110000110",
  2739=>"001100011",
  2740=>"111110110",
  2741=>"011111101",
  2742=>"010011011",
  2743=>"001110010",
  2744=>"100010011",
  2745=>"101001111",
  2746=>"001011101",
  2747=>"010011110",
  2748=>"111100111",
  2749=>"101010111",
  2750=>"001010011",
  2751=>"110100100",
  2752=>"010100010",
  2753=>"011000100",
  2754=>"101011111",
  2755=>"111011110",
  2756=>"011010011",
  2757=>"001100100",
  2758=>"110001011",
  2759=>"100000011",
  2760=>"111010010",
  2761=>"111101100",
  2762=>"101001001",
  2763=>"001111000",
  2764=>"000101011",
  2765=>"011100110",
  2766=>"110001101",
  2767=>"001110100",
  2768=>"110101001",
  2769=>"000110100",
  2770=>"110111110",
  2771=>"111001011",
  2772=>"000011000",
  2773=>"111101001",
  2774=>"010011110",
  2775=>"011011010",
  2776=>"001011011",
  2777=>"010111010",
  2778=>"111101101",
  2779=>"111011101",
  2780=>"101101111",
  2781=>"111111000",
  2782=>"000110010",
  2783=>"100010100",
  2784=>"111100111",
  2785=>"110110111",
  2786=>"100101111",
  2787=>"101111111",
  2788=>"101100000",
  2789=>"111110110",
  2790=>"101010011",
  2791=>"001010110",
  2792=>"101001110",
  2793=>"111001100",
  2794=>"100110010",
  2795=>"001101101",
  2796=>"011010011",
  2797=>"111010111",
  2798=>"101110110",
  2799=>"001010100",
  2800=>"000011100",
  2801=>"110110100",
  2802=>"101011111",
  2803=>"011111011",
  2804=>"010111000",
  2805=>"111100111",
  2806=>"000000111",
  2807=>"111001010",
  2808=>"001110001",
  2809=>"001001100",
  2810=>"001011011",
  2811=>"001000101",
  2812=>"010100001",
  2813=>"000011110",
  2814=>"110001010",
  2815=>"111011111",
  2816=>"010000101",
  2817=>"000110101",
  2818=>"110111100",
  2819=>"101111101",
  2820=>"011100011",
  2821=>"101000010",
  2822=>"000011001",
  2823=>"010100110",
  2824=>"100011001",
  2825=>"111010000",
  2826=>"010010011",
  2827=>"100111100",
  2828=>"111000000",
  2829=>"111001100",
  2830=>"101010110",
  2831=>"010101111",
  2832=>"010111011",
  2833=>"100001000",
  2834=>"000011101",
  2835=>"100100111",
  2836=>"111110100",
  2837=>"011110101",
  2838=>"110001101",
  2839=>"110100100",
  2840=>"111101101",
  2841=>"001011110",
  2842=>"000000101",
  2843=>"011110111",
  2844=>"101111110",
  2845=>"000111000",
  2846=>"110010001",
  2847=>"110001110",
  2848=>"100110010",
  2849=>"000011101",
  2850=>"101111010",
  2851=>"011000001",
  2852=>"011011011",
  2853=>"111100101",
  2854=>"001111000",
  2855=>"011010100",
  2856=>"100011000",
  2857=>"001011001",
  2858=>"101000110",
  2859=>"010011011",
  2860=>"001000011",
  2861=>"110011110",
  2862=>"100101000",
  2863=>"010100110",
  2864=>"101100001",
  2865=>"100110110",
  2866=>"111000111",
  2867=>"000001101",
  2868=>"010100110",
  2869=>"010000110",
  2870=>"001111010",
  2871=>"110111110",
  2872=>"101111101",
  2873=>"000000111",
  2874=>"011011101",
  2875=>"100111100",
  2876=>"000000010",
  2877=>"110101111",
  2878=>"000000000",
  2879=>"011010111",
  2880=>"100001011",
  2881=>"001110100",
  2882=>"010010100",
  2883=>"101010100",
  2884=>"000011010",
  2885=>"010110010",
  2886=>"111111111",
  2887=>"111100000",
  2888=>"111110111",
  2889=>"111101010",
  2890=>"000001101",
  2891=>"000011110",
  2892=>"101111110",
  2893=>"000000001",
  2894=>"010111111",
  2895=>"110001000",
  2896=>"111011001",
  2897=>"101100000",
  2898=>"000111110",
  2899=>"010101010",
  2900=>"110001100",
  2901=>"011011101",
  2902=>"001001000",
  2903=>"011011010",
  2904=>"110010101",
  2905=>"110110001",
  2906=>"111010101",
  2907=>"100101001",
  2908=>"101101111",
  2909=>"101001100",
  2910=>"100010110",
  2911=>"001000010",
  2912=>"100111011",
  2913=>"111101111",
  2914=>"000001000",
  2915=>"011000101",
  2916=>"011100101",
  2917=>"100101010",
  2918=>"101100110",
  2919=>"100111110",
  2920=>"011101001",
  2921=>"011011111",
  2922=>"001000001",
  2923=>"011010111",
  2924=>"011100101",
  2925=>"000001100",
  2926=>"011100100",
  2927=>"100000100",
  2928=>"100100111",
  2929=>"000100000",
  2930=>"100011011",
  2931=>"000000111",
  2932=>"000010011",
  2933=>"101110011",
  2934=>"100000110",
  2935=>"000001000",
  2936=>"110010000",
  2937=>"000010101",
  2938=>"010100100",
  2939=>"110010011",
  2940=>"010100100",
  2941=>"111101111",
  2942=>"100110110",
  2943=>"100110010",
  2944=>"101001111",
  2945=>"000001101",
  2946=>"111010001",
  2947=>"100001100",
  2948=>"000001101",
  2949=>"101011010",
  2950=>"000111010",
  2951=>"011000110",
  2952=>"101111101",
  2953=>"000011001",
  2954=>"111110111",
  2955=>"010101000",
  2956=>"111010101",
  2957=>"010101001",
  2958=>"111100111",
  2959=>"101011110",
  2960=>"000110001",
  2961=>"101111001",
  2962=>"101011001",
  2963=>"000100101",
  2964=>"010100100",
  2965=>"001000110",
  2966=>"110010001",
  2967=>"101001010",
  2968=>"110111001",
  2969=>"111100111",
  2970=>"111011110",
  2971=>"100101001",
  2972=>"111101000",
  2973=>"011011010",
  2974=>"100100101",
  2975=>"101001011",
  2976=>"101111010",
  2977=>"111011011",
  2978=>"111100110",
  2979=>"011000111",
  2980=>"001101100",
  2981=>"010111100",
  2982=>"111111111",
  2983=>"110111101",
  2984=>"000111111",
  2985=>"101111111",
  2986=>"010110001",
  2987=>"111110101",
  2988=>"000010110",
  2989=>"001110001",
  2990=>"000111101",
  2991=>"000111111",
  2992=>"011010011",
  2993=>"111110110",
  2994=>"100011100",
  2995=>"100001111",
  2996=>"111100110",
  2997=>"010001101",
  2998=>"000010001",
  2999=>"101011010",
  3000=>"110101000",
  3001=>"011101111",
  3002=>"011001111",
  3003=>"010001010",
  3004=>"001001111",
  3005=>"111100000",
  3006=>"010111101",
  3007=>"111111101",
  3008=>"000111110",
  3009=>"000101110",
  3010=>"011000101",
  3011=>"000100000",
  3012=>"100001000",
  3013=>"101000111",
  3014=>"100100001",
  3015=>"000100001",
  3016=>"010010011",
  3017=>"010000001",
  3018=>"001011000",
  3019=>"111110110",
  3020=>"101001010",
  3021=>"111100001",
  3022=>"000000111",
  3023=>"001011010",
  3024=>"001110001",
  3025=>"001000100",
  3026=>"101101111",
  3027=>"110101111",
  3028=>"000110111",
  3029=>"110000101",
  3030=>"110011101",
  3031=>"011001000",
  3032=>"010011010",
  3033=>"111101101",
  3034=>"011001100",
  3035=>"010100001",
  3036=>"100011110",
  3037=>"000010000",
  3038=>"111011101",
  3039=>"101001010",
  3040=>"001010110",
  3041=>"110010011",
  3042=>"111000110",
  3043=>"110111110",
  3044=>"101111001",
  3045=>"001110010",
  3046=>"001110110",
  3047=>"111100100",
  3048=>"000100111",
  3049=>"100111011",
  3050=>"100001110",
  3051=>"000000001",
  3052=>"010101000",
  3053=>"100001111",
  3054=>"110110011",
  3055=>"010001100",
  3056=>"100000011",
  3057=>"110011100",
  3058=>"011100000",
  3059=>"001010101",
  3060=>"100000100",
  3061=>"000000000",
  3062=>"111011101",
  3063=>"000100010",
  3064=>"111100001",
  3065=>"010101011",
  3066=>"001010000",
  3067=>"001110000",
  3068=>"111100111",
  3069=>"110111100",
  3070=>"100011001",
  3071=>"000100110",
  3072=>"100010111",
  3073=>"001100001",
  3074=>"101011111",
  3075=>"101100000",
  3076=>"001111101",
  3077=>"100100111",
  3078=>"100010010",
  3079=>"100110010",
  3080=>"001011000",
  3081=>"101011001",
  3082=>"110111110",
  3083=>"001111010",
  3084=>"100011111",
  3085=>"010001101",
  3086=>"000100000",
  3087=>"001100001",
  3088=>"010100011",
  3089=>"100010111",
  3090=>"011000010",
  3091=>"010010111",
  3092=>"010111111",
  3093=>"010110100",
  3094=>"101111011",
  3095=>"001011100",
  3096=>"001000000",
  3097=>"100110110",
  3098=>"011100101",
  3099=>"110101001",
  3100=>"100110010",
  3101=>"111101110",
  3102=>"100010100",
  3103=>"000001001",
  3104=>"111001011",
  3105=>"111011100",
  3106=>"101000100",
  3107=>"110011111",
  3108=>"111011110",
  3109=>"000100010",
  3110=>"000111101",
  3111=>"110000011",
  3112=>"100111000",
  3113=>"100010000",
  3114=>"000110001",
  3115=>"000101010",
  3116=>"111000001",
  3117=>"010010010",
  3118=>"111010100",
  3119=>"000111010",
  3120=>"001010010",
  3121=>"100011100",
  3122=>"011000001",
  3123=>"001011000",
  3124=>"110110110",
  3125=>"110010100",
  3126=>"011110001",
  3127=>"011111111",
  3128=>"111110000",
  3129=>"000011101",
  3130=>"100101111",
  3131=>"001100101",
  3132=>"100110011",
  3133=>"000110011",
  3134=>"110011111",
  3135=>"001100101",
  3136=>"011011111",
  3137=>"000100010",
  3138=>"110111100",
  3139=>"101100001",
  3140=>"000000110",
  3141=>"000001111",
  3142=>"111010100",
  3143=>"010100000",
  3144=>"000101111",
  3145=>"101101110",
  3146=>"100000000",
  3147=>"111111001",
  3148=>"101010010",
  3149=>"111101001",
  3150=>"111100100",
  3151=>"111100010",
  3152=>"001101011",
  3153=>"000110110",
  3154=>"001010001",
  3155=>"011011001",
  3156=>"111111010",
  3157=>"010101111",
  3158=>"110001111",
  3159=>"110011111",
  3160=>"110000000",
  3161=>"111011111",
  3162=>"010100011",
  3163=>"111101111",
  3164=>"011011100",
  3165=>"011101000",
  3166=>"001010111",
  3167=>"000100010",
  3168=>"001011011",
  3169=>"111101101",
  3170=>"010011111",
  3171=>"000001001",
  3172=>"101001001",
  3173=>"011110110",
  3174=>"011111101",
  3175=>"010011001",
  3176=>"101011000",
  3177=>"110111011",
  3178=>"000010000",
  3179=>"101110101",
  3180=>"101110000",
  3181=>"001110000",
  3182=>"010110110",
  3183=>"001001101",
  3184=>"100010010",
  3185=>"011010010",
  3186=>"101001100",
  3187=>"101010101",
  3188=>"100001101",
  3189=>"010010011",
  3190=>"110010010",
  3191=>"101001111",
  3192=>"000110100",
  3193=>"000001010",
  3194=>"110000111",
  3195=>"010001101",
  3196=>"101000011",
  3197=>"101010100",
  3198=>"001111101",
  3199=>"111010010",
  3200=>"110110000",
  3201=>"100101000",
  3202=>"011010001",
  3203=>"011110101",
  3204=>"110110101",
  3205=>"110001101",
  3206=>"001011100",
  3207=>"011010010",
  3208=>"110100110",
  3209=>"100001010",
  3210=>"111111100",
  3211=>"001000000",
  3212=>"111001111",
  3213=>"111000100",
  3214=>"000000000",
  3215=>"110011001",
  3216=>"100101110",
  3217=>"100111011",
  3218=>"001011001",
  3219=>"110101100",
  3220=>"111000111",
  3221=>"010110110",
  3222=>"010101010",
  3223=>"110001101",
  3224=>"011101011",
  3225=>"000100000",
  3226=>"100101111",
  3227=>"010110000",
  3228=>"110110010",
  3229=>"011110101",
  3230=>"000001101",
  3231=>"110001000",
  3232=>"101011101",
  3233=>"100010110",
  3234=>"101101100",
  3235=>"000010011",
  3236=>"111111100",
  3237=>"001010100",
  3238=>"100100111",
  3239=>"101111110",
  3240=>"100010010",
  3241=>"001101110",
  3242=>"011101101",
  3243=>"000000100",
  3244=>"100011111",
  3245=>"110110110",
  3246=>"110100110",
  3247=>"001000000",
  3248=>"101111110",
  3249=>"010111101",
  3250=>"100000011",
  3251=>"000000010",
  3252=>"110111001",
  3253=>"111110111",
  3254=>"000110010",
  3255=>"101111010",
  3256=>"011100110",
  3257=>"101010001",
  3258=>"101111110",
  3259=>"010011100",
  3260=>"001110000",
  3261=>"011001101",
  3262=>"010100101",
  3263=>"100100000",
  3264=>"000110010",
  3265=>"000110000",
  3266=>"000101010",
  3267=>"000001100",
  3268=>"010111101",
  3269=>"000110000",
  3270=>"100011000",
  3271=>"110011000",
  3272=>"001100110",
  3273=>"111111100",
  3274=>"001101101",
  3275=>"100011111",
  3276=>"101001111",
  3277=>"101011000",
  3278=>"000101101",
  3279=>"000010000",
  3280=>"100001001",
  3281=>"100000010",
  3282=>"011111111",
  3283=>"010110100",
  3284=>"000011000",
  3285=>"101010100",
  3286=>"000000101",
  3287=>"111001101",
  3288=>"101100101",
  3289=>"000110101",
  3290=>"111111000",
  3291=>"000100100",
  3292=>"110101101",
  3293=>"010010001",
  3294=>"110100010",
  3295=>"010110011",
  3296=>"101110000",
  3297=>"111111110",
  3298=>"010100111",
  3299=>"000010000",
  3300=>"100111000",
  3301=>"111000001",
  3302=>"010010100",
  3303=>"011000100",
  3304=>"111101001",
  3305=>"011001011",
  3306=>"100001110",
  3307=>"010001000",
  3308=>"111001001",
  3309=>"110101100",
  3310=>"100010101",
  3311=>"001010110",
  3312=>"001110011",
  3313=>"111011111",
  3314=>"100011000",
  3315=>"101001111",
  3316=>"000101001",
  3317=>"110011110",
  3318=>"101011110",
  3319=>"110110000",
  3320=>"010110000",
  3321=>"100010001",
  3322=>"000001001",
  3323=>"000000101",
  3324=>"001001000",
  3325=>"111111100",
  3326=>"110100111",
  3327=>"111110000",
  3328=>"011000110",
  3329=>"111010100",
  3330=>"101000000",
  3331=>"011010001",
  3332=>"010111110",
  3333=>"101101100",
  3334=>"110111001",
  3335=>"011111111",
  3336=>"100011110",
  3337=>"111000000",
  3338=>"001110110",
  3339=>"111011111",
  3340=>"010001001",
  3341=>"010110110",
  3342=>"110100001",
  3343=>"011110001",
  3344=>"100110111",
  3345=>"001010101",
  3346=>"111101101",
  3347=>"001001010",
  3348=>"001011001",
  3349=>"101101011",
  3350=>"111010110",
  3351=>"100111011",
  3352=>"101011001",
  3353=>"111111001",
  3354=>"011111111",
  3355=>"000011001",
  3356=>"000000111",
  3357=>"101011010",
  3358=>"100010010",
  3359=>"111010111",
  3360=>"110001010",
  3361=>"110010001",
  3362=>"101100001",
  3363=>"011100011",
  3364=>"001010000",
  3365=>"100111011",
  3366=>"000011110",
  3367=>"010100100",
  3368=>"100101001",
  3369=>"010011001",
  3370=>"110000000",
  3371=>"101000101",
  3372=>"001100001",
  3373=>"110111110",
  3374=>"000111011",
  3375=>"001100100",
  3376=>"101110101",
  3377=>"101101111",
  3378=>"101001100",
  3379=>"000011011",
  3380=>"100100001",
  3381=>"011111010",
  3382=>"000100000",
  3383=>"010111001",
  3384=>"011001000",
  3385=>"111010111",
  3386=>"011001111",
  3387=>"000100111",
  3388=>"000000001",
  3389=>"111010000",
  3390=>"100010100",
  3391=>"000000110",
  3392=>"100111111",
  3393=>"100110001",
  3394=>"100100100",
  3395=>"101101000",
  3396=>"100011101",
  3397=>"101011100",
  3398=>"101110010",
  3399=>"010111010",
  3400=>"111001010",
  3401=>"001011101",
  3402=>"110010111",
  3403=>"101111111",
  3404=>"001001101",
  3405=>"101110001",
  3406=>"001111001",
  3407=>"101111010",
  3408=>"010100100",
  3409=>"111110011",
  3410=>"000111110",
  3411=>"110111110",
  3412=>"001100001",
  3413=>"111111101",
  3414=>"010000110",
  3415=>"111110111",
  3416=>"001011000",
  3417=>"001100011",
  3418=>"000001101",
  3419=>"011101011",
  3420=>"011110010",
  3421=>"101101101",
  3422=>"111111101",
  3423=>"010010111",
  3424=>"000110011",
  3425=>"011100000",
  3426=>"010100001",
  3427=>"111010000",
  3428=>"111000001",
  3429=>"010011100",
  3430=>"111110010",
  3431=>"010000011",
  3432=>"111100110",
  3433=>"111110010",
  3434=>"111111000",
  3435=>"110101010",
  3436=>"110101001",
  3437=>"000010100",
  3438=>"100111100",
  3439=>"100001000",
  3440=>"011111001",
  3441=>"001111111",
  3442=>"011110111",
  3443=>"110101101",
  3444=>"101011111",
  3445=>"000010100",
  3446=>"110010010",
  3447=>"000010110",
  3448=>"110101101",
  3449=>"000010010",
  3450=>"100100010",
  3451=>"100101110",
  3452=>"010111111",
  3453=>"001011110",
  3454=>"110101000",
  3455=>"011001111",
  3456=>"110110101",
  3457=>"000000000",
  3458=>"001001001",
  3459=>"000010000",
  3460=>"011010110",
  3461=>"000111000",
  3462=>"111011110",
  3463=>"000010110",
  3464=>"111010100",
  3465=>"010001101",
  3466=>"011011000",
  3467=>"100110101",
  3468=>"100111110",
  3469=>"110100010",
  3470=>"111001101",
  3471=>"111000101",
  3472=>"101100010",
  3473=>"100101001",
  3474=>"010100011",
  3475=>"110101010",
  3476=>"110000100",
  3477=>"111101111",
  3478=>"010100111",
  3479=>"100110101",
  3480=>"111001111",
  3481=>"001110001",
  3482=>"100011111",
  3483=>"101001000",
  3484=>"110110110",
  3485=>"101110110",
  3486=>"111011011",
  3487=>"110111101",
  3488=>"101111000",
  3489=>"100101000",
  3490=>"001101110",
  3491=>"111101001",
  3492=>"110011101",
  3493=>"001000000",
  3494=>"000000011",
  3495=>"000000001",
  3496=>"111110101",
  3497=>"111110000",
  3498=>"000101111",
  3499=>"011111010",
  3500=>"100110111",
  3501=>"111000001",
  3502=>"100000010",
  3503=>"100011101",
  3504=>"110111111",
  3505=>"101111001",
  3506=>"111101001",
  3507=>"000101111",
  3508=>"000100110",
  3509=>"101110011",
  3510=>"110110111",
  3511=>"100011101",
  3512=>"101111101",
  3513=>"101111101",
  3514=>"010111101",
  3515=>"110010100",
  3516=>"100001111",
  3517=>"110010000",
  3518=>"100110011",
  3519=>"111110000",
  3520=>"011100001",
  3521=>"000010010",
  3522=>"001110110",
  3523=>"110100011",
  3524=>"010011111",
  3525=>"110001100",
  3526=>"011111111",
  3527=>"101111011",
  3528=>"100100100",
  3529=>"000100111",
  3530=>"001100001",
  3531=>"000100111",
  3532=>"011101101",
  3533=>"101111110",
  3534=>"101000111",
  3535=>"011001111",
  3536=>"101001011",
  3537=>"000010100",
  3538=>"001111111",
  3539=>"000001011",
  3540=>"101010101",
  3541=>"110000110",
  3542=>"001010010",
  3543=>"111110010",
  3544=>"000000110",
  3545=>"010001100",
  3546=>"010000010",
  3547=>"111111000",
  3548=>"010010100",
  3549=>"000101110",
  3550=>"110101010",
  3551=>"111000110",
  3552=>"001111110",
  3553=>"101000001",
  3554=>"100000101",
  3555=>"011110000",
  3556=>"001000101",
  3557=>"011100000",
  3558=>"101100110",
  3559=>"101100100",
  3560=>"001101101",
  3561=>"100110101",
  3562=>"011111000",
  3563=>"010001001",
  3564=>"110011000",
  3565=>"110000100",
  3566=>"011001011",
  3567=>"111110110",
  3568=>"011001111",
  3569=>"100010100",
  3570=>"001101100",
  3571=>"010101111",
  3572=>"000101001",
  3573=>"000111011",
  3574=>"101001011",
  3575=>"101011001",
  3576=>"110100111",
  3577=>"010010011",
  3578=>"011111110",
  3579=>"010000000",
  3580=>"111001110",
  3581=>"110011111",
  3582=>"000111010",
  3583=>"100110100",
  3584=>"001001001",
  3585=>"000111000",
  3586=>"110110000",
  3587=>"011111101",
  3588=>"000010110",
  3589=>"011111101",
  3590=>"000010000",
  3591=>"111100101",
  3592=>"011010111",
  3593=>"110111000",
  3594=>"000100010",
  3595=>"111111001",
  3596=>"001000111",
  3597=>"010000101",
  3598=>"010111101",
  3599=>"110110000",
  3600=>"010010001",
  3601=>"111000110",
  3602=>"000001011",
  3603=>"111001000",
  3604=>"100010110",
  3605=>"101110010",
  3606=>"000111110",
  3607=>"100101000",
  3608=>"110011110",
  3609=>"010110111",
  3610=>"111100001",
  3611=>"111001100",
  3612=>"001111100",
  3613=>"111100001",
  3614=>"100011101",
  3615=>"010111000",
  3616=>"010011100",
  3617=>"010111111",
  3618=>"111001110",
  3619=>"001001110",
  3620=>"011110011",
  3621=>"111000010",
  3622=>"000100011",
  3623=>"100110000",
  3624=>"101101010",
  3625=>"101010000",
  3626=>"110100000",
  3627=>"111111000",
  3628=>"000000001",
  3629=>"000110011",
  3630=>"000011110",
  3631=>"100111111",
  3632=>"011100101",
  3633=>"111011010",
  3634=>"010001010",
  3635=>"111000011",
  3636=>"111111011",
  3637=>"101000000",
  3638=>"000001101",
  3639=>"011001010",
  3640=>"111011000",
  3641=>"010011010",
  3642=>"010011000",
  3643=>"101110100",
  3644=>"111111111",
  3645=>"111110110",
  3646=>"110100100",
  3647=>"011010001",
  3648=>"011100011",
  3649=>"011011011",
  3650=>"100000111",
  3651=>"111111011",
  3652=>"111001111",
  3653=>"001011100",
  3654=>"110111100",
  3655=>"000011011",
  3656=>"110111111",
  3657=>"101010010",
  3658=>"000111111",
  3659=>"010011000",
  3660=>"100010010",
  3661=>"100100111",
  3662=>"111011111",
  3663=>"001101011",
  3664=>"111011000",
  3665=>"000011101",
  3666=>"000111111",
  3667=>"110000101",
  3668=>"110101101",
  3669=>"101110111",
  3670=>"000101000",
  3671=>"100110110",
  3672=>"010001100",
  3673=>"111110110",
  3674=>"001010100",
  3675=>"100111010",
  3676=>"111100111",
  3677=>"000100110",
  3678=>"111100001",
  3679=>"101000101",
  3680=>"110101010",
  3681=>"100001100",
  3682=>"101100110",
  3683=>"010100000",
  3684=>"100001101",
  3685=>"101100110",
  3686=>"111110011",
  3687=>"010110100",
  3688=>"010000011",
  3689=>"011000011",
  3690=>"001110000",
  3691=>"110111111",
  3692=>"000000100",
  3693=>"100110011",
  3694=>"100110100",
  3695=>"001010110",
  3696=>"111100101",
  3697=>"000101110",
  3698=>"001011011",
  3699=>"010000101",
  3700=>"101100000",
  3701=>"110011110",
  3702=>"110000000",
  3703=>"001111110",
  3704=>"000010001",
  3705=>"001111111",
  3706=>"111111011",
  3707=>"001001111",
  3708=>"111111000",
  3709=>"100101110",
  3710=>"111101011",
  3711=>"100010010",
  3712=>"011111000",
  3713=>"101011101",
  3714=>"000000000",
  3715=>"111110110",
  3716=>"011111100",
  3717=>"111101111",
  3718=>"010110000",
  3719=>"100111111",
  3720=>"101111010",
  3721=>"001001010",
  3722=>"101010011",
  3723=>"011011111",
  3724=>"000100101",
  3725=>"000111000",
  3726=>"010011111",
  3727=>"011001000",
  3728=>"011000000",
  3729=>"011100001",
  3730=>"011010101",
  3731=>"100110001",
  3732=>"111001101",
  3733=>"001101111",
  3734=>"101111001",
  3735=>"001111011",
  3736=>"001100100",
  3737=>"100000111",
  3738=>"010000011",
  3739=>"101100001",
  3740=>"100010010",
  3741=>"010000000",
  3742=>"110000001",
  3743=>"011000001",
  3744=>"101010000",
  3745=>"101011000",
  3746=>"111101000",
  3747=>"010001101",
  3748=>"011111101",
  3749=>"010001011",
  3750=>"010101100",
  3751=>"000010001",
  3752=>"110110101",
  3753=>"110000100",
  3754=>"000011110",
  3755=>"111100010",
  3756=>"100011001",
  3757=>"110110010",
  3758=>"101000101",
  3759=>"110101011",
  3760=>"100011100",
  3761=>"010000011",
  3762=>"101010010",
  3763=>"011110101",
  3764=>"100011100",
  3765=>"011100001",
  3766=>"111000010",
  3767=>"011100010",
  3768=>"011110011",
  3769=>"000010000",
  3770=>"100000001",
  3771=>"011111001",
  3772=>"111000111",
  3773=>"010010111",
  3774=>"000101111",
  3775=>"000011000",
  3776=>"011011010",
  3777=>"100110110",
  3778=>"111111000",
  3779=>"000000010",
  3780=>"011110001",
  3781=>"101111000",
  3782=>"110101011",
  3783=>"100010111",
  3784=>"000010110",
  3785=>"110110011",
  3786=>"110111110",
  3787=>"001010101",
  3788=>"111101100",
  3789=>"001111010",
  3790=>"111010010",
  3791=>"100110011",
  3792=>"101111111",
  3793=>"000011110",
  3794=>"010100111",
  3795=>"010100001",
  3796=>"111011001",
  3797=>"111000001",
  3798=>"000101110",
  3799=>"011111111",
  3800=>"101101000",
  3801=>"100000001",
  3802=>"001101000",
  3803=>"000110000",
  3804=>"110010101",
  3805=>"000100111",
  3806=>"001110101",
  3807=>"010111100",
  3808=>"011101100",
  3809=>"110000001",
  3810=>"100001010",
  3811=>"011101011",
  3812=>"001001111",
  3813=>"100110111",
  3814=>"000001011",
  3815=>"111100100",
  3816=>"101001101",
  3817=>"100001010",
  3818=>"001001111",
  3819=>"111011101",
  3820=>"111000001",
  3821=>"111110110",
  3822=>"011111111",
  3823=>"110010001",
  3824=>"000001100",
  3825=>"010011010",
  3826=>"010111011",
  3827=>"001000001",
  3828=>"101100111",
  3829=>"111000001",
  3830=>"001101001",
  3831=>"110000111",
  3832=>"010010011",
  3833=>"010011111",
  3834=>"100011111",
  3835=>"011101110",
  3836=>"011111011",
  3837=>"110010110",
  3838=>"010010100",
  3839=>"100101101",
  3840=>"000110101",
  3841=>"010000001",
  3842=>"100010001",
  3843=>"001001000",
  3844=>"111001101",
  3845=>"001110001",
  3846=>"001010100",
  3847=>"101010101",
  3848=>"010111110",
  3849=>"111001000",
  3850=>"101101001",
  3851=>"101011101",
  3852=>"000110001",
  3853=>"100000010",
  3854=>"111001010",
  3855=>"101101000",
  3856=>"100101110",
  3857=>"100100011",
  3858=>"101101010",
  3859=>"010100110",
  3860=>"001000100",
  3861=>"010101011",
  3862=>"001000011",
  3863=>"100000001",
  3864=>"001101001",
  3865=>"010110001",
  3866=>"111111110",
  3867=>"011000001",
  3868=>"110110010",
  3869=>"100111000",
  3870=>"111011111",
  3871=>"011001011",
  3872=>"010110100",
  3873=>"011001000",
  3874=>"100101001",
  3875=>"011000000",
  3876=>"000100010",
  3877=>"100111111",
  3878=>"000101001",
  3879=>"101001110",
  3880=>"110000100",
  3881=>"011001011",
  3882=>"100100001",
  3883=>"001001000",
  3884=>"101100000",
  3885=>"000010111",
  3886=>"011001101",
  3887=>"110010101",
  3888=>"100111111",
  3889=>"011001001",
  3890=>"000010101",
  3891=>"101011110",
  3892=>"011111111",
  3893=>"101010110",
  3894=>"000100110",
  3895=>"000111100",
  3896=>"100011011",
  3897=>"000011001",
  3898=>"111101111",
  3899=>"011111100",
  3900=>"000111011",
  3901=>"100001110",
  3902=>"101010100",
  3903=>"110001000",
  3904=>"011000000",
  3905=>"100111110",
  3906=>"111101011",
  3907=>"101000011",
  3908=>"011110111",
  3909=>"000110111",
  3910=>"000000001",
  3911=>"101000101",
  3912=>"111100000",
  3913=>"011100000",
  3914=>"111001000",
  3915=>"000010111",
  3916=>"110100100",
  3917=>"000001111",
  3918=>"111001001",
  3919=>"101101101",
  3920=>"000100111",
  3921=>"110001100",
  3922=>"111110000",
  3923=>"101101100",
  3924=>"011100001",
  3925=>"001001110",
  3926=>"101001010",
  3927=>"011010000",
  3928=>"110101111",
  3929=>"101001110",
  3930=>"111010100",
  3931=>"011101111",
  3932=>"111010110",
  3933=>"110101111",
  3934=>"100100001",
  3935=>"000111110",
  3936=>"010101100",
  3937=>"111110111",
  3938=>"100111110",
  3939=>"011101100",
  3940=>"110100111",
  3941=>"001110100",
  3942=>"011010111",
  3943=>"101010001",
  3944=>"011000001",
  3945=>"011000000",
  3946=>"001100001",
  3947=>"100111000",
  3948=>"101111001",
  3949=>"101000000",
  3950=>"010101101",
  3951=>"111010101",
  3952=>"111110110",
  3953=>"010010010",
  3954=>"011110111",
  3955=>"100101100",
  3956=>"110010100",
  3957=>"111011001",
  3958=>"000110000",
  3959=>"100010100",
  3960=>"010011010",
  3961=>"110110110",
  3962=>"011010100",
  3963=>"100101111",
  3964=>"110000011",
  3965=>"101111100",
  3966=>"111111000",
  3967=>"101010101",
  3968=>"100101001",
  3969=>"111010111",
  3970=>"111111101",
  3971=>"111100010",
  3972=>"100001101",
  3973=>"010100000",
  3974=>"001101101",
  3975=>"100101101",
  3976=>"110111000",
  3977=>"011000100",
  3978=>"111011101",
  3979=>"000011000",
  3980=>"011110100",
  3981=>"101010111",
  3982=>"101111001",
  3983=>"100011110",
  3984=>"011111010",
  3985=>"111010001",
  3986=>"110001000",
  3987=>"000111000",
  3988=>"011001010",
  3989=>"011001000",
  3990=>"111011001",
  3991=>"001010010",
  3992=>"111001101",
  3993=>"110001110",
  3994=>"110011100",
  3995=>"101001111",
  3996=>"000001010",
  3997=>"001000100",
  3998=>"011011010",
  3999=>"010001010",
  4000=>"011010100",
  4001=>"010100011",
  4002=>"110010000",
  4003=>"010010110",
  4004=>"100100010",
  4005=>"011111001",
  4006=>"111010011",
  4007=>"010001100",
  4008=>"110010111",
  4009=>"100011001",
  4010=>"011110001",
  4011=>"110110010",
  4012=>"011000010",
  4013=>"010110010",
  4014=>"010010110",
  4015=>"110111110",
  4016=>"100000000",
  4017=>"111001100",
  4018=>"001011010",
  4019=>"000101110",
  4020=>"011010110",
  4021=>"001101111",
  4022=>"101111101",
  4023=>"010000000",
  4024=>"001111011",
  4025=>"101111010",
  4026=>"100100010",
  4027=>"111101110",
  4028=>"011001101",
  4029=>"110100111",
  4030=>"000110111",
  4031=>"001100000",
  4032=>"011100001",
  4033=>"000000110",
  4034=>"010101011",
  4035=>"101101010",
  4036=>"101001110",
  4037=>"000010111",
  4038=>"001011101",
  4039=>"111001110",
  4040=>"110111111",
  4041=>"110000100",
  4042=>"101110111",
  4043=>"011111000",
  4044=>"100111101",
  4045=>"001010101",
  4046=>"011000100",
  4047=>"111101111",
  4048=>"111110101",
  4049=>"000001001",
  4050=>"100110001",
  4051=>"111011111",
  4052=>"001111100",
  4053=>"111111100",
  4054=>"010000001",
  4055=>"101000000",
  4056=>"001110101",
  4057=>"111101100",
  4058=>"100111100",
  4059=>"010000110",
  4060=>"010000000",
  4061=>"110010110",
  4062=>"001001111",
  4063=>"011011011",
  4064=>"010011111",
  4065=>"000011001",
  4066=>"001000110",
  4067=>"000010000",
  4068=>"010111111",
  4069=>"010010011",
  4070=>"011001101",
  4071=>"111110010",
  4072=>"100010000",
  4073=>"100111100",
  4074=>"000010111",
  4075=>"011001110",
  4076=>"001000010",
  4077=>"000000000",
  4078=>"000000001",
  4079=>"010111011",
  4080=>"110110010",
  4081=>"000110100",
  4082=>"100001100",
  4083=>"100010111",
  4084=>"111100010",
  4085=>"111001010",
  4086=>"110001011",
  4087=>"010010010",
  4088=>"111110111",
  4089=>"011111010",
  4090=>"101111010",
  4091=>"000010001",
  4092=>"100001001",
  4093=>"101001110",
  4094=>"111011001",
  4095=>"110000010",
  4096=>"101101001",
  4097=>"101110100",
  4098=>"101000101",
  4099=>"101011000",
  4100=>"110111001",
  4101=>"101010000",
  4102=>"111001111",
  4103=>"111111011",
  4104=>"000110000",
  4105=>"100011011",
  4106=>"011111110",
  4107=>"001101111",
  4108=>"100000000",
  4109=>"101100010",
  4110=>"101001100",
  4111=>"001000000",
  4112=>"101101110",
  4113=>"000000000",
  4114=>"011011011",
  4115=>"001101100",
  4116=>"011100000",
  4117=>"101111010",
  4118=>"100010011",
  4119=>"101101101",
  4120=>"000001010",
  4121=>"100100100",
  4122=>"001101100",
  4123=>"101000110",
  4124=>"010110100",
  4125=>"001010110",
  4126=>"001011100",
  4127=>"111000001",
  4128=>"001101000",
  4129=>"111000000",
  4130=>"111000110",
  4131=>"011111100",
  4132=>"010110111",
  4133=>"010011110",
  4134=>"011001000",
  4135=>"011101000",
  4136=>"100001111",
  4137=>"001000011",
  4138=>"100101010",
  4139=>"110010011",
  4140=>"000111110",
  4141=>"110110101",
  4142=>"111111010",
  4143=>"001100001",
  4144=>"011111110",
  4145=>"011011000",
  4146=>"100110111",
  4147=>"011011111",
  4148=>"100100010",
  4149=>"111000001",
  4150=>"101000000",
  4151=>"111001110",
  4152=>"111000011",
  4153=>"011011111",
  4154=>"010001010",
  4155=>"011001110",
  4156=>"010100001",
  4157=>"110010001",
  4158=>"100100111",
  4159=>"000000001",
  4160=>"001110000",
  4161=>"000111000",
  4162=>"001010001",
  4163=>"101011001",
  4164=>"110010000",
  4165=>"011101001",
  4166=>"001100111",
  4167=>"010111010",
  4168=>"111111011",
  4169=>"011010000",
  4170=>"010111011",
  4171=>"111000010",
  4172=>"101000001",
  4173=>"000110011",
  4174=>"010111110",
  4175=>"111000100",
  4176=>"000110010",
  4177=>"010011011",
  4178=>"001100101",
  4179=>"110001011",
  4180=>"100000000",
  4181=>"110000110",
  4182=>"001111011",
  4183=>"100011110",
  4184=>"011011001",
  4185=>"111101101",
  4186=>"001011100",
  4187=>"110110000",
  4188=>"100100000",
  4189=>"110100000",
  4190=>"110111101",
  4191=>"011000010",
  4192=>"101101010",
  4193=>"000110101",
  4194=>"111111011",
  4195=>"001001001",
  4196=>"001011111",
  4197=>"110000010",
  4198=>"101101010",
  4199=>"000101110",
  4200=>"000111000",
  4201=>"110100011",
  4202=>"001001100",
  4203=>"111000111",
  4204=>"100111001",
  4205=>"111011100",
  4206=>"100010000",
  4207=>"000000001",
  4208=>"111100110",
  4209=>"101101100",
  4210=>"101001011",
  4211=>"011010110",
  4212=>"101110000",
  4213=>"101001110",
  4214=>"111011110",
  4215=>"011000111",
  4216=>"010001111",
  4217=>"110101000",
  4218=>"000010010",
  4219=>"011011100",
  4220=>"101111110",
  4221=>"001000111",
  4222=>"111101111",
  4223=>"100100100",
  4224=>"001001000",
  4225=>"111100101",
  4226=>"101110110",
  4227=>"101010100",
  4228=>"110111000",
  4229=>"111100011",
  4230=>"001000000",
  4231=>"001110011",
  4232=>"010011110",
  4233=>"111110100",
  4234=>"111100111",
  4235=>"100100110",
  4236=>"101100100",
  4237=>"110011010",
  4238=>"000001101",
  4239=>"011000100",
  4240=>"011001110",
  4241=>"111110100",
  4242=>"010010100",
  4243=>"101000111",
  4244=>"000010001",
  4245=>"000101101",
  4246=>"001111000",
  4247=>"000001110",
  4248=>"101111110",
  4249=>"000100110",
  4250=>"010001101",
  4251=>"011100111",
  4252=>"000111101",
  4253=>"101101111",
  4254=>"000010111",
  4255=>"010001011",
  4256=>"100100000",
  4257=>"011011110",
  4258=>"110011111",
  4259=>"101000000",
  4260=>"000111111",
  4261=>"000111001",
  4262=>"111111000",
  4263=>"100011010",
  4264=>"011110011",
  4265=>"111001001",
  4266=>"111000010",
  4267=>"111101101",
  4268=>"100101110",
  4269=>"111011110",
  4270=>"011011010",
  4271=>"110011000",
  4272=>"001011011",
  4273=>"111111000",
  4274=>"000011110",
  4275=>"011011101",
  4276=>"011000100",
  4277=>"110110001",
  4278=>"111111001",
  4279=>"111000101",
  4280=>"101010010",
  4281=>"110111011",
  4282=>"110011000",
  4283=>"011111111",
  4284=>"110010001",
  4285=>"011101111",
  4286=>"110010111",
  4287=>"100000000",
  4288=>"010001110",
  4289=>"011110010",
  4290=>"110001101",
  4291=>"110100000",
  4292=>"100110011",
  4293=>"101010011",
  4294=>"001000000",
  4295=>"100101000",
  4296=>"010010011",
  4297=>"011000100",
  4298=>"001110010",
  4299=>"110011001",
  4300=>"101010011",
  4301=>"011101010",
  4302=>"010011001",
  4303=>"011100011",
  4304=>"101111001",
  4305=>"110000000",
  4306=>"000101101",
  4307=>"111111010",
  4308=>"001110000",
  4309=>"110111110",
  4310=>"000100100",
  4311=>"111111001",
  4312=>"011000100",
  4313=>"010000100",
  4314=>"000011001",
  4315=>"110111101",
  4316=>"011101010",
  4317=>"000011100",
  4318=>"101000010",
  4319=>"010110100",
  4320=>"111110001",
  4321=>"110000011",
  4322=>"000100101",
  4323=>"100011011",
  4324=>"000000001",
  4325=>"110011111",
  4326=>"001001001",
  4327=>"011011001",
  4328=>"000111011",
  4329=>"100110001",
  4330=>"000000110",
  4331=>"010000011",
  4332=>"001110000",
  4333=>"000010011",
  4334=>"001010000",
  4335=>"010010010",
  4336=>"111110111",
  4337=>"011000111",
  4338=>"011000100",
  4339=>"100110101",
  4340=>"010010010",
  4341=>"001001001",
  4342=>"001110001",
  4343=>"011100010",
  4344=>"000101100",
  4345=>"110000011",
  4346=>"011001001",
  4347=>"101011010",
  4348=>"111000000",
  4349=>"010100100",
  4350=>"000001001",
  4351=>"011111111",
  4352=>"110001001",
  4353=>"110000100",
  4354=>"111011100",
  4355=>"111111011",
  4356=>"001001001",
  4357=>"101010001",
  4358=>"100001010",
  4359=>"000000001",
  4360=>"000000000",
  4361=>"100101101",
  4362=>"111001010",
  4363=>"100001011",
  4364=>"101111010",
  4365=>"100001000",
  4366=>"101100011",
  4367=>"100110000",
  4368=>"011000110",
  4369=>"000100100",
  4370=>"000100100",
  4371=>"011110101",
  4372=>"100011111",
  4373=>"000000101",
  4374=>"010101011",
  4375=>"110000010",
  4376=>"111110101",
  4377=>"001101110",
  4378=>"111000111",
  4379=>"111101110",
  4380=>"101001001",
  4381=>"010010010",
  4382=>"100101000",
  4383=>"111000110",
  4384=>"001010111",
  4385=>"111010000",
  4386=>"011000111",
  4387=>"001010111",
  4388=>"000000000",
  4389=>"010001100",
  4390=>"001100111",
  4391=>"101011011",
  4392=>"100110010",
  4393=>"100001000",
  4394=>"011011100",
  4395=>"100110001",
  4396=>"000001100",
  4397=>"100010111",
  4398=>"011001101",
  4399=>"101100110",
  4400=>"111110100",
  4401=>"000111100",
  4402=>"110011100",
  4403=>"001011000",
  4404=>"111110010",
  4405=>"101010110",
  4406=>"011011001",
  4407=>"100001101",
  4408=>"000000100",
  4409=>"101101011",
  4410=>"001000101",
  4411=>"101011010",
  4412=>"011001010",
  4413=>"001110010",
  4414=>"100011011",
  4415=>"011001111",
  4416=>"100100010",
  4417=>"111100011",
  4418=>"101111111",
  4419=>"111101111",
  4420=>"001100101",
  4421=>"101111000",
  4422=>"010101000",
  4423=>"000101101",
  4424=>"110000010",
  4425=>"101000001",
  4426=>"010010011",
  4427=>"001110111",
  4428=>"001000000",
  4429=>"111111111",
  4430=>"000100100",
  4431=>"001000010",
  4432=>"001101010",
  4433=>"011101100",
  4434=>"000000011",
  4435=>"011101111",
  4436=>"011111000",
  4437=>"010000000",
  4438=>"111111110",
  4439=>"000001100",
  4440=>"100100010",
  4441=>"011010110",
  4442=>"111001000",
  4443=>"001010111",
  4444=>"010100000",
  4445=>"111011101",
  4446=>"111010111",
  4447=>"111110001",
  4448=>"011011001",
  4449=>"100111000",
  4450=>"111010101",
  4451=>"010111100",
  4452=>"101101111",
  4453=>"001111111",
  4454=>"110101101",
  4455=>"101000110",
  4456=>"101011011",
  4457=>"100000000",
  4458=>"001110100",
  4459=>"101110100",
  4460=>"100011101",
  4461=>"100001000",
  4462=>"111001001",
  4463=>"011101001",
  4464=>"110010110",
  4465=>"010101010",
  4466=>"100010110",
  4467=>"111111111",
  4468=>"000010100",
  4469=>"111101011",
  4470=>"011100001",
  4471=>"111111100",
  4472=>"111001111",
  4473=>"001000111",
  4474=>"011110100",
  4475=>"010110110",
  4476=>"010000110",
  4477=>"101111010",
  4478=>"000000101",
  4479=>"111110011",
  4480=>"010101110",
  4481=>"011101111",
  4482=>"001100001",
  4483=>"100111100",
  4484=>"001101011",
  4485=>"010111011",
  4486=>"001010101",
  4487=>"000010001",
  4488=>"110100010",
  4489=>"111101100",
  4490=>"111100101",
  4491=>"010011001",
  4492=>"011010011",
  4493=>"101001010",
  4494=>"110011000",
  4495=>"001110111",
  4496=>"101101011",
  4497=>"111110101",
  4498=>"010100001",
  4499=>"001001111",
  4500=>"001111001",
  4501=>"010000010",
  4502=>"110111011",
  4503=>"101111101",
  4504=>"000010000",
  4505=>"100100100",
  4506=>"010111010",
  4507=>"100101111",
  4508=>"000000010",
  4509=>"010001010",
  4510=>"101111010",
  4511=>"000000010",
  4512=>"000010000",
  4513=>"100001100",
  4514=>"110011010",
  4515=>"111000000",
  4516=>"100001101",
  4517=>"000111100",
  4518=>"001011011",
  4519=>"000011110",
  4520=>"110111101",
  4521=>"011101101",
  4522=>"110010100",
  4523=>"001011100",
  4524=>"001111001",
  4525=>"011100110",
  4526=>"000011011",
  4527=>"100011100",
  4528=>"010100101",
  4529=>"001001111",
  4530=>"010000100",
  4531=>"001011101",
  4532=>"000111010",
  4533=>"011011001",
  4534=>"111011000",
  4535=>"101111001",
  4536=>"111010111",
  4537=>"001001111",
  4538=>"110110001",
  4539=>"011111010",
  4540=>"100011010",
  4541=>"111101111",
  4542=>"100101010",
  4543=>"010100010",
  4544=>"000011001",
  4545=>"101001010",
  4546=>"000001110",
  4547=>"000100110",
  4548=>"111100000",
  4549=>"011011000",
  4550=>"010100101",
  4551=>"100010000",
  4552=>"110001100",
  4553=>"111001010",
  4554=>"110000100",
  4555=>"001101101",
  4556=>"110010010",
  4557=>"101010001",
  4558=>"110011111",
  4559=>"111000110",
  4560=>"110100110",
  4561=>"000010010",
  4562=>"011101011",
  4563=>"110000111",
  4564=>"010010110",
  4565=>"100000011",
  4566=>"101100010",
  4567=>"000101011",
  4568=>"100000011",
  4569=>"111111101",
  4570=>"100010011",
  4571=>"010111010",
  4572=>"001011010",
  4573=>"011010001",
  4574=>"110110111",
  4575=>"110101100",
  4576=>"010000001",
  4577=>"011100110",
  4578=>"001100010",
  4579=>"101000110",
  4580=>"011011010",
  4581=>"111110000",
  4582=>"010000110",
  4583=>"110011111",
  4584=>"110101100",
  4585=>"001110101",
  4586=>"110010000",
  4587=>"010101100",
  4588=>"100101101",
  4589=>"111110100",
  4590=>"000110100",
  4591=>"101110011",
  4592=>"000100011",
  4593=>"111111000",
  4594=>"010101100",
  4595=>"110000000",
  4596=>"110101101",
  4597=>"001011101",
  4598=>"011101101",
  4599=>"010000100",
  4600=>"011111100",
  4601=>"111100101",
  4602=>"111011111",
  4603=>"101011101",
  4604=>"101010111",
  4605=>"001011101",
  4606=>"010110001",
  4607=>"100100001",
  4608=>"000001011",
  4609=>"101101101",
  4610=>"001000010",
  4611=>"011000101",
  4612=>"100000010",
  4613=>"010001100",
  4614=>"000010100",
  4615=>"000111101",
  4616=>"111111111",
  4617=>"111010101",
  4618=>"110110011",
  4619=>"000000110",
  4620=>"010011111",
  4621=>"101101001",
  4622=>"011010110",
  4623=>"110001101",
  4624=>"101011010",
  4625=>"110101100",
  4626=>"110011001",
  4627=>"010000000",
  4628=>"011011011",
  4629=>"110101101",
  4630=>"111010101",
  4631=>"110010010",
  4632=>"111100001",
  4633=>"100111001",
  4634=>"110011000",
  4635=>"101001110",
  4636=>"111011111",
  4637=>"011001011",
  4638=>"000001001",
  4639=>"011011011",
  4640=>"100111110",
  4641=>"111010000",
  4642=>"000110101",
  4643=>"001010001",
  4644=>"100010110",
  4645=>"010011010",
  4646=>"111111011",
  4647=>"010111010",
  4648=>"010001111",
  4649=>"110001101",
  4650=>"110100100",
  4651=>"000110100",
  4652=>"111101101",
  4653=>"110001111",
  4654=>"010110100",
  4655=>"000001010",
  4656=>"111000110",
  4657=>"011010010",
  4658=>"101101110",
  4659=>"101110101",
  4660=>"100111001",
  4661=>"010001100",
  4662=>"110010100",
  4663=>"000111011",
  4664=>"001100010",
  4665=>"001001000",
  4666=>"101100100",
  4667=>"101000110",
  4668=>"011110100",
  4669=>"011001000",
  4670=>"010001111",
  4671=>"010110011",
  4672=>"000000100",
  4673=>"111110000",
  4674=>"101001011",
  4675=>"110000100",
  4676=>"100011101",
  4677=>"001001001",
  4678=>"100010001",
  4679=>"010110101",
  4680=>"100011110",
  4681=>"101101000",
  4682=>"101011000",
  4683=>"000000111",
  4684=>"101110000",
  4685=>"000110011",
  4686=>"101111000",
  4687=>"101010101",
  4688=>"111111011",
  4689=>"011000101",
  4690=>"101011010",
  4691=>"011011111",
  4692=>"011011010",
  4693=>"010010100",
  4694=>"101110011",
  4695=>"100011001",
  4696=>"111011010",
  4697=>"110101100",
  4698=>"001100000",
  4699=>"011110110",
  4700=>"000101011",
  4701=>"100010010",
  4702=>"111111010",
  4703=>"000001101",
  4704=>"001100110",
  4705=>"111000100",
  4706=>"110101010",
  4707=>"100011110",
  4708=>"001000100",
  4709=>"000101010",
  4710=>"111010101",
  4711=>"011111000",
  4712=>"110100000",
  4713=>"001011011",
  4714=>"101111010",
  4715=>"100010010",
  4716=>"110110000",
  4717=>"000110001",
  4718=>"101101000",
  4719=>"000111011",
  4720=>"101101111",
  4721=>"001111001",
  4722=>"101000000",
  4723=>"011110010",
  4724=>"011111111",
  4725=>"010010110",
  4726=>"000001011",
  4727=>"000110010",
  4728=>"101100101",
  4729=>"111011101",
  4730=>"111010111",
  4731=>"010001100",
  4732=>"001000001",
  4733=>"111100100",
  4734=>"101101110",
  4735=>"000111000",
  4736=>"000001110",
  4737=>"000000111",
  4738=>"001010100",
  4739=>"010110111",
  4740=>"111101000",
  4741=>"101010001",
  4742=>"010100111",
  4743=>"011101001",
  4744=>"000011101",
  4745=>"100110100",
  4746=>"000000010",
  4747=>"101101011",
  4748=>"000001001",
  4749=>"010110000",
  4750=>"110000100",
  4751=>"001110000",
  4752=>"011100100",
  4753=>"001101001",
  4754=>"111010111",
  4755=>"010111011",
  4756=>"011000110",
  4757=>"110000000",
  4758=>"001100110",
  4759=>"110100010",
  4760=>"101001110",
  4761=>"110111110",
  4762=>"010110010",
  4763=>"001000001",
  4764=>"111110110",
  4765=>"000011001",
  4766=>"100111111",
  4767=>"010110011",
  4768=>"101100111",
  4769=>"110010110",
  4770=>"111011010",
  4771=>"101010011",
  4772=>"011011001",
  4773=>"011000001",
  4774=>"111001011",
  4775=>"010110110",
  4776=>"100011000",
  4777=>"011010110",
  4778=>"010111011",
  4779=>"111101110",
  4780=>"111111010",
  4781=>"111111111",
  4782=>"000010001",
  4783=>"100001011",
  4784=>"100111111",
  4785=>"010111010",
  4786=>"111010000",
  4787=>"000111111",
  4788=>"100010110",
  4789=>"110100100",
  4790=>"010111101",
  4791=>"100000000",
  4792=>"001011011",
  4793=>"110010011",
  4794=>"110000000",
  4795=>"111000000",
  4796=>"111110011",
  4797=>"011011011",
  4798=>"000101000",
  4799=>"101100110",
  4800=>"100001100",
  4801=>"001010010",
  4802=>"011000110",
  4803=>"000010001",
  4804=>"000011011",
  4805=>"010101110",
  4806=>"110100010",
  4807=>"100101110",
  4808=>"111101111",
  4809=>"001110110",
  4810=>"011010100",
  4811=>"001001111",
  4812=>"100010000",
  4813=>"101101101",
  4814=>"101010010",
  4815=>"010100010",
  4816=>"111011000",
  4817=>"101101110",
  4818=>"110011000",
  4819=>"111101000",
  4820=>"101101110",
  4821=>"111110010",
  4822=>"101110100",
  4823=>"001100001",
  4824=>"011000101",
  4825=>"011001100",
  4826=>"111110000",
  4827=>"100010101",
  4828=>"111000101",
  4829=>"001001110",
  4830=>"100011110",
  4831=>"110100100",
  4832=>"101101101",
  4833=>"100100111",
  4834=>"001000010",
  4835=>"101101011",
  4836=>"111101110",
  4837=>"001010010",
  4838=>"011100000",
  4839=>"000100010",
  4840=>"010101111",
  4841=>"011111101",
  4842=>"100000011",
  4843=>"011101111",
  4844=>"000111111",
  4845=>"010011010",
  4846=>"101111100",
  4847=>"000100000",
  4848=>"011111010",
  4849=>"101010011",
  4850=>"000000101",
  4851=>"001001100",
  4852=>"100100110",
  4853=>"111100110",
  4854=>"000111110",
  4855=>"011100001",
  4856=>"010010000",
  4857=>"001110001",
  4858=>"100010000",
  4859=>"001111000",
  4860=>"001010001",
  4861=>"000101010",
  4862=>"110011110",
  4863=>"010111000",
  4864=>"001010110",
  4865=>"000011111",
  4866=>"010001011",
  4867=>"011000110",
  4868=>"111010001",
  4869=>"011111001",
  4870=>"010110110",
  4871=>"010011011",
  4872=>"001100100",
  4873=>"000101011",
  4874=>"010110101",
  4875=>"101110001",
  4876=>"111001000",
  4877=>"000111000",
  4878=>"001001011",
  4879=>"110010110",
  4880=>"101100100",
  4881=>"111001101",
  4882=>"111100000",
  4883=>"000110111",
  4884=>"010001011",
  4885=>"010101001",
  4886=>"110100100",
  4887=>"010000000",
  4888=>"110111111",
  4889=>"110110101",
  4890=>"001001101",
  4891=>"111000100",
  4892=>"111100111",
  4893=>"000110101",
  4894=>"010010000",
  4895=>"111100011",
  4896=>"110111100",
  4897=>"001010110",
  4898=>"101110111",
  4899=>"010101101",
  4900=>"110101010",
  4901=>"100101010",
  4902=>"001110001",
  4903=>"000110011",
  4904=>"100010011",
  4905=>"110100100",
  4906=>"100101000",
  4907=>"011111111",
  4908=>"000110101",
  4909=>"111111010",
  4910=>"011110100",
  4911=>"100101000",
  4912=>"101011100",
  4913=>"100100100",
  4914=>"100011110",
  4915=>"010000101",
  4916=>"100011011",
  4917=>"000000010",
  4918=>"101110011",
  4919=>"011000101",
  4920=>"010001011",
  4921=>"010000000",
  4922=>"100010011",
  4923=>"010011000",
  4924=>"011110101",
  4925=>"111100010",
  4926=>"111001000",
  4927=>"011010000",
  4928=>"001010011",
  4929=>"000010111",
  4930=>"111001000",
  4931=>"001110010",
  4932=>"011100011",
  4933=>"000110000",
  4934=>"001010001",
  4935=>"001011010",
  4936=>"011111011",
  4937=>"000101010",
  4938=>"000011000",
  4939=>"010011111",
  4940=>"110100110",
  4941=>"011100010",
  4942=>"101000000",
  4943=>"000110000",
  4944=>"100000100",
  4945=>"000100001",
  4946=>"111001101",
  4947=>"100000001",
  4948=>"000100000",
  4949=>"111011000",
  4950=>"111100000",
  4951=>"000010011",
  4952=>"110101011",
  4953=>"111110001",
  4954=>"001110101",
  4955=>"100010111",
  4956=>"100101010",
  4957=>"001000111",
  4958=>"011100111",
  4959=>"110000101",
  4960=>"010101100",
  4961=>"110011011",
  4962=>"101100100",
  4963=>"011101001",
  4964=>"111001011",
  4965=>"100011001",
  4966=>"110110110",
  4967=>"110010110",
  4968=>"011111011",
  4969=>"000111011",
  4970=>"010110100",
  4971=>"111001000",
  4972=>"010111110",
  4973=>"111110000",
  4974=>"000000000",
  4975=>"011110100",
  4976=>"011100000",
  4977=>"101101010",
  4978=>"011111011",
  4979=>"111101011",
  4980=>"100011110",
  4981=>"111101010",
  4982=>"000111011",
  4983=>"100110110",
  4984=>"011001001",
  4985=>"111010000",
  4986=>"111101101",
  4987=>"000000010",
  4988=>"001110000",
  4989=>"111111001",
  4990=>"001100010",
  4991=>"111111011",
  4992=>"001111000",
  4993=>"111000010",
  4994=>"010100011",
  4995=>"111001000",
  4996=>"101011001",
  4997=>"011100111",
  4998=>"000010100",
  4999=>"111111111",
  5000=>"110101011",
  5001=>"111000000",
  5002=>"011101000",
  5003=>"001011001",
  5004=>"001011011",
  5005=>"010001100",
  5006=>"000101010",
  5007=>"010011010",
  5008=>"010010000",
  5009=>"010011000",
  5010=>"110000011",
  5011=>"001000000",
  5012=>"111111100",
  5013=>"000100001",
  5014=>"000010000",
  5015=>"101110110",
  5016=>"000001011",
  5017=>"000001000",
  5018=>"101010010",
  5019=>"001100000",
  5020=>"110100001",
  5021=>"011111111",
  5022=>"110000101",
  5023=>"000001000",
  5024=>"111001100",
  5025=>"110010111",
  5026=>"011111000",
  5027=>"110101000",
  5028=>"001000101",
  5029=>"101000100",
  5030=>"100011111",
  5031=>"000001111",
  5032=>"100110000",
  5033=>"001101101",
  5034=>"111111000",
  5035=>"111100101",
  5036=>"000010010",
  5037=>"001000110",
  5038=>"100001010",
  5039=>"010011000",
  5040=>"010011001",
  5041=>"001001000",
  5042=>"011110011",
  5043=>"010111101",
  5044=>"010010110",
  5045=>"111100110",
  5046=>"101101111",
  5047=>"110011010",
  5048=>"010011111",
  5049=>"001001110",
  5050=>"000101100",
  5051=>"010100101",
  5052=>"101011101",
  5053=>"111000010",
  5054=>"010100100",
  5055=>"010011110",
  5056=>"010110001",
  5057=>"101100001",
  5058=>"111101000",
  5059=>"110000110",
  5060=>"000100000",
  5061=>"010010000",
  5062=>"110111111",
  5063=>"001011010",
  5064=>"101100000",
  5065=>"000001010",
  5066=>"100111110",
  5067=>"001101100",
  5068=>"001001000",
  5069=>"010101000",
  5070=>"111100110",
  5071=>"100110111",
  5072=>"111100101",
  5073=>"001111110",
  5074=>"000110111",
  5075=>"101010011",
  5076=>"010110110",
  5077=>"111100111",
  5078=>"001000110",
  5079=>"011010010",
  5080=>"010000001",
  5081=>"011001000",
  5082=>"001000101",
  5083=>"000010110",
  5084=>"001101001",
  5085=>"100010110",
  5086=>"011011100",
  5087=>"110011011",
  5088=>"111111111",
  5089=>"111111100",
  5090=>"010100010",
  5091=>"111010100",
  5092=>"011000100",
  5093=>"110101010",
  5094=>"110101111",
  5095=>"101110101",
  5096=>"010001000",
  5097=>"011101100",
  5098=>"010001101",
  5099=>"001101111",
  5100=>"110111100",
  5101=>"010000101",
  5102=>"111001110",
  5103=>"011011101",
  5104=>"011100011",
  5105=>"001001111",
  5106=>"111001011",
  5107=>"100000010",
  5108=>"100001010",
  5109=>"011001101",
  5110=>"000000001",
  5111=>"011000001",
  5112=>"010000000",
  5113=>"111111111",
  5114=>"000101010",
  5115=>"111111001",
  5116=>"001101011",
  5117=>"011001000",
  5118=>"000101010",
  5119=>"000111110",
  5120=>"001000100",
  5121=>"010101010",
  5122=>"000111011",
  5123=>"100110110",
  5124=>"111000111",
  5125=>"100101100",
  5126=>"001101101",
  5127=>"011010100",
  5128=>"010110011",
  5129=>"110110110",
  5130=>"000010100",
  5131=>"000000001",
  5132=>"101110111",
  5133=>"001110010",
  5134=>"110010001",
  5135=>"110100000",
  5136=>"011001111",
  5137=>"000000101",
  5138=>"011000011",
  5139=>"111110111",
  5140=>"000110001",
  5141=>"000001011",
  5142=>"111111000",
  5143=>"100000000",
  5144=>"010000011",
  5145=>"101111100",
  5146=>"010001110",
  5147=>"001001110",
  5148=>"110110010",
  5149=>"011010000",
  5150=>"011111000",
  5151=>"110110100",
  5152=>"010011111",
  5153=>"010000000",
  5154=>"000101000",
  5155=>"001101110",
  5156=>"011111000",
  5157=>"000100100",
  5158=>"000100011",
  5159=>"000111111",
  5160=>"000111000",
  5161=>"110100111",
  5162=>"111001111",
  5163=>"001111100",
  5164=>"011110110",
  5165=>"111001111",
  5166=>"001011110",
  5167=>"101000101",
  5168=>"110010011",
  5169=>"110110100",
  5170=>"001001011",
  5171=>"100101010",
  5172=>"010110110",
  5173=>"011111001",
  5174=>"000011110",
  5175=>"111001011",
  5176=>"110101011",
  5177=>"000100000",
  5178=>"100011010",
  5179=>"101111101",
  5180=>"101111001",
  5181=>"100101100",
  5182=>"100100110",
  5183=>"100000011",
  5184=>"111100100",
  5185=>"000111010",
  5186=>"001000111",
  5187=>"010010111",
  5188=>"000010110",
  5189=>"111100010",
  5190=>"000001101",
  5191=>"101010111",
  5192=>"001101011",
  5193=>"100010001",
  5194=>"010111110",
  5195=>"011000011",
  5196=>"100100000",
  5197=>"100001011",
  5198=>"110100110",
  5199=>"000111111",
  5200=>"001010000",
  5201=>"011101001",
  5202=>"001111101",
  5203=>"000000011",
  5204=>"000101101",
  5205=>"001000011",
  5206=>"110101010",
  5207=>"000100110",
  5208=>"100011011",
  5209=>"010111111",
  5210=>"010100100",
  5211=>"000001100",
  5212=>"111100010",
  5213=>"111101010",
  5214=>"000101111",
  5215=>"010100001",
  5216=>"101101101",
  5217=>"010101000",
  5218=>"100111000",
  5219=>"010001001",
  5220=>"001000011",
  5221=>"111110101",
  5222=>"110101010",
  5223=>"110000000",
  5224=>"100001001",
  5225=>"010111001",
  5226=>"000000110",
  5227=>"001111110",
  5228=>"000000001",
  5229=>"110111000",
  5230=>"101000111",
  5231=>"100111010",
  5232=>"001010011",
  5233=>"011111110",
  5234=>"111100110",
  5235=>"100100101",
  5236=>"000011000",
  5237=>"000111101",
  5238=>"101111010",
  5239=>"000011101",
  5240=>"011011000",
  5241=>"010011111",
  5242=>"110011000",
  5243=>"001010100",
  5244=>"001010110",
  5245=>"000010110",
  5246=>"000011000",
  5247=>"111011100",
  5248=>"001011010",
  5249=>"000000110",
  5250=>"100001001",
  5251=>"000000011",
  5252=>"010101111",
  5253=>"001000000",
  5254=>"110110111",
  5255=>"100000110",
  5256=>"111111000",
  5257=>"010100110",
  5258=>"001110000",
  5259=>"100100110",
  5260=>"000010001",
  5261=>"001001001",
  5262=>"110101011",
  5263=>"000000100",
  5264=>"001110111",
  5265=>"001010010",
  5266=>"100101111",
  5267=>"110110111",
  5268=>"001000010",
  5269=>"001100111",
  5270=>"100101101",
  5271=>"110101101",
  5272=>"001011001",
  5273=>"000101010",
  5274=>"010111100",
  5275=>"001000111",
  5276=>"000011110",
  5277=>"010011110",
  5278=>"101110101",
  5279=>"100111111",
  5280=>"100110010",
  5281=>"111000001",
  5282=>"011100111",
  5283=>"110001101",
  5284=>"000001011",
  5285=>"010011000",
  5286=>"000101110",
  5287=>"010111000",
  5288=>"101000110",
  5289=>"111010000",
  5290=>"111010111",
  5291=>"110100110",
  5292=>"011100010",
  5293=>"111011111",
  5294=>"111100001",
  5295=>"001100010",
  5296=>"101000100",
  5297=>"110111010",
  5298=>"111001111",
  5299=>"000011011",
  5300=>"010111001",
  5301=>"010000101",
  5302=>"000110100",
  5303=>"000010011",
  5304=>"010111001",
  5305=>"101011011",
  5306=>"111001001",
  5307=>"010000010",
  5308=>"001111010",
  5309=>"100000000",
  5310=>"011101011",
  5311=>"101000100",
  5312=>"100100011",
  5313=>"011111110",
  5314=>"101001000",
  5315=>"100111101",
  5316=>"110110110",
  5317=>"111100010",
  5318=>"001011100",
  5319=>"011111000",
  5320=>"010101111",
  5321=>"101000111",
  5322=>"100101101",
  5323=>"011011001",
  5324=>"001101000",
  5325=>"000011110",
  5326=>"000101101",
  5327=>"100100010",
  5328=>"101011111",
  5329=>"101111001",
  5330=>"100010011",
  5331=>"100000101",
  5332=>"011111000",
  5333=>"111110000",
  5334=>"011100011",
  5335=>"110100111",
  5336=>"010110110",
  5337=>"010010011",
  5338=>"000101011",
  5339=>"001011110",
  5340=>"110011001",
  5341=>"101001101",
  5342=>"111101001",
  5343=>"110011010",
  5344=>"101111110",
  5345=>"000000110",
  5346=>"110010000",
  5347=>"010101000",
  5348=>"110101101",
  5349=>"000110010",
  5350=>"001100110",
  5351=>"011110110",
  5352=>"000011100",
  5353=>"011101010",
  5354=>"111001011",
  5355=>"111101001",
  5356=>"100010100",
  5357=>"010000010",
  5358=>"011000110",
  5359=>"011010000",
  5360=>"000110001",
  5361=>"010000000",
  5362=>"010100101",
  5363=>"000010111",
  5364=>"011111001",
  5365=>"101010111",
  5366=>"101000010",
  5367=>"001011011",
  5368=>"111111010",
  5369=>"101010101",
  5370=>"011000110",
  5371=>"011111000",
  5372=>"010101111",
  5373=>"011111110",
  5374=>"011001101",
  5375=>"111111001",
  5376=>"001100100",
  5377=>"110111010",
  5378=>"110111011",
  5379=>"010110010",
  5380=>"111010000",
  5381=>"010011000",
  5382=>"001100111",
  5383=>"000101001",
  5384=>"100101101",
  5385=>"011010111",
  5386=>"010111011",
  5387=>"111101110",
  5388=>"101000000",
  5389=>"000101000",
  5390=>"101100010",
  5391=>"000000001",
  5392=>"100010011",
  5393=>"100000011",
  5394=>"101110000",
  5395=>"101110011",
  5396=>"001010000",
  5397=>"101111010",
  5398=>"010011111",
  5399=>"101111110",
  5400=>"011001110",
  5401=>"000000110",
  5402=>"011100100",
  5403=>"001101110",
  5404=>"100110011",
  5405=>"000101111",
  5406=>"000001000",
  5407=>"001001000",
  5408=>"011000000",
  5409=>"000100011",
  5410=>"011110111",
  5411=>"010101100",
  5412=>"110010011",
  5413=>"110001100",
  5414=>"110011110",
  5415=>"000011101",
  5416=>"110000101",
  5417=>"101010010",
  5418=>"111101011",
  5419=>"011100001",
  5420=>"011101001",
  5421=>"100100000",
  5422=>"101001110",
  5423=>"000100000",
  5424=>"011101011",
  5425=>"011000010",
  5426=>"110011111",
  5427=>"001101101",
  5428=>"110111110",
  5429=>"010110000",
  5430=>"101101111",
  5431=>"110101111",
  5432=>"000010110",
  5433=>"010011001",
  5434=>"000100110",
  5435=>"100001110",
  5436=>"101000010",
  5437=>"100111100",
  5438=>"111000001",
  5439=>"100110111",
  5440=>"001011000",
  5441=>"010010111",
  5442=>"000110101",
  5443=>"110101001",
  5444=>"011011011",
  5445=>"010110101",
  5446=>"000100010",
  5447=>"101110011",
  5448=>"000110000",
  5449=>"001010100",
  5450=>"110011100",
  5451=>"100100001",
  5452=>"100011000",
  5453=>"111111010",
  5454=>"100001010",
  5455=>"001000111",
  5456=>"001101101",
  5457=>"000100010",
  5458=>"010001010",
  5459=>"001111100",
  5460=>"111000101",
  5461=>"010000110",
  5462=>"010010011",
  5463=>"111001110",
  5464=>"110011100",
  5465=>"111001001",
  5466=>"000000101",
  5467=>"111110000",
  5468=>"110111110",
  5469=>"010101010",
  5470=>"000100000",
  5471=>"001111110",
  5472=>"101101001",
  5473=>"010011110",
  5474=>"111100100",
  5475=>"111001100",
  5476=>"000001011",
  5477=>"010010011",
  5478=>"001010011",
  5479=>"111000101",
  5480=>"010111011",
  5481=>"000110100",
  5482=>"000110110",
  5483=>"000111110",
  5484=>"110010110",
  5485=>"111111010",
  5486=>"001011000",
  5487=>"111011011",
  5488=>"110101101",
  5489=>"000001000",
  5490=>"111011000",
  5491=>"100001110",
  5492=>"101001111",
  5493=>"110000110",
  5494=>"000110101",
  5495=>"110010001",
  5496=>"110101100",
  5497=>"000010110",
  5498=>"100001111",
  5499=>"000101110",
  5500=>"010101101",
  5501=>"010010101",
  5502=>"000001011",
  5503=>"011010100",
  5504=>"101101111",
  5505=>"001111001",
  5506=>"111110000",
  5507=>"111010111",
  5508=>"011110111",
  5509=>"001000011",
  5510=>"000010111",
  5511=>"011100100",
  5512=>"110101111",
  5513=>"011101011",
  5514=>"101000101",
  5515=>"000000010",
  5516=>"010001111",
  5517=>"100111111",
  5518=>"100000101",
  5519=>"111000100",
  5520=>"010010101",
  5521=>"000000010",
  5522=>"111101011",
  5523=>"100110101",
  5524=>"011000001",
  5525=>"000110100",
  5526=>"010010010",
  5527=>"110010000",
  5528=>"100010000",
  5529=>"100101011",
  5530=>"000011110",
  5531=>"111010101",
  5532=>"110101000",
  5533=>"101111101",
  5534=>"100100001",
  5535=>"010010111",
  5536=>"000110000",
  5537=>"101111011",
  5538=>"000100011",
  5539=>"110001000",
  5540=>"100101001",
  5541=>"000111001",
  5542=>"111100111",
  5543=>"001111010",
  5544=>"100001111",
  5545=>"001010101",
  5546=>"000011011",
  5547=>"010100110",
  5548=>"101011110",
  5549=>"110111101",
  5550=>"110111011",
  5551=>"010011100",
  5552=>"010110110",
  5553=>"010000001",
  5554=>"100100111",
  5555=>"101000111",
  5556=>"101110111",
  5557=>"001011100",
  5558=>"101111100",
  5559=>"111110000",
  5560=>"000000111",
  5561=>"111010000",
  5562=>"010001011",
  5563=>"111100111",
  5564=>"101010000",
  5565=>"111110011",
  5566=>"111001010",
  5567=>"111001100",
  5568=>"011000111",
  5569=>"000000111",
  5570=>"011100001",
  5571=>"101001010",
  5572=>"011010011",
  5573=>"110100010",
  5574=>"011001010",
  5575=>"010101000",
  5576=>"111010100",
  5577=>"010111010",
  5578=>"000110010",
  5579=>"001110000",
  5580=>"100000011",
  5581=>"001110100",
  5582=>"011100001",
  5583=>"110000111",
  5584=>"011010101",
  5585=>"000101001",
  5586=>"001001111",
  5587=>"001010001",
  5588=>"000001001",
  5589=>"001110101",
  5590=>"010001111",
  5591=>"111101100",
  5592=>"010011011",
  5593=>"111001101",
  5594=>"010011100",
  5595=>"101000000",
  5596=>"010101001",
  5597=>"011001110",
  5598=>"111101000",
  5599=>"001010100",
  5600=>"010010000",
  5601=>"111001011",
  5602=>"111001010",
  5603=>"100110010",
  5604=>"010011010",
  5605=>"101111000",
  5606=>"111010110",
  5607=>"111111110",
  5608=>"000100010",
  5609=>"001000010",
  5610=>"010000000",
  5611=>"111011010",
  5612=>"011100000",
  5613=>"101111011",
  5614=>"000011011",
  5615=>"100110110",
  5616=>"010111000",
  5617=>"110101100",
  5618=>"100010110",
  5619=>"111010100",
  5620=>"111001010",
  5621=>"111101111",
  5622=>"001000100",
  5623=>"000000011",
  5624=>"010010101",
  5625=>"111111010",
  5626=>"010010000",
  5627=>"111001110",
  5628=>"011010010",
  5629=>"101100110",
  5630=>"011000001",
  5631=>"100100101",
  5632=>"011011100",
  5633=>"000100010",
  5634=>"111011110",
  5635=>"101101010",
  5636=>"110010000",
  5637=>"010100001",
  5638=>"010100001",
  5639=>"100000001",
  5640=>"100000100",
  5641=>"111000010",
  5642=>"100101101",
  5643=>"000001100",
  5644=>"101010100",
  5645=>"100100111",
  5646=>"001110000",
  5647=>"001001001",
  5648=>"111101011",
  5649=>"000111100",
  5650=>"111011011",
  5651=>"011100000",
  5652=>"100001000",
  5653=>"000100100",
  5654=>"101001001",
  5655=>"111110001",
  5656=>"110101111",
  5657=>"100100111",
  5658=>"110001000",
  5659=>"000000001",
  5660=>"010111111",
  5661=>"010111100",
  5662=>"100011101",
  5663=>"011010101",
  5664=>"000000101",
  5665=>"000010110",
  5666=>"000010010",
  5667=>"101111000",
  5668=>"000010000",
  5669=>"010101011",
  5670=>"111110110",
  5671=>"101101101",
  5672=>"100000011",
  5673=>"010110110",
  5674=>"101101000",
  5675=>"111010110",
  5676=>"001101100",
  5677=>"011001010",
  5678=>"001000010",
  5679=>"110010010",
  5680=>"101011111",
  5681=>"100011100",
  5682=>"000111110",
  5683=>"001010001",
  5684=>"110011011",
  5685=>"011101110",
  5686=>"110000101",
  5687=>"000101011",
  5688=>"100010000",
  5689=>"100100100",
  5690=>"100001000",
  5691=>"110001101",
  5692=>"100110011",
  5693=>"000011110",
  5694=>"111000111",
  5695=>"101000000",
  5696=>"000100101",
  5697=>"111111101",
  5698=>"101011010",
  5699=>"000001010",
  5700=>"100010110",
  5701=>"000000110",
  5702=>"110100111",
  5703=>"010100001",
  5704=>"001001100",
  5705=>"101111111",
  5706=>"111010011",
  5707=>"110100011",
  5708=>"010000001",
  5709=>"110111000",
  5710=>"110110101",
  5711=>"010100110",
  5712=>"110010101",
  5713=>"100011000",
  5714=>"001000001",
  5715=>"000100000",
  5716=>"001001011",
  5717=>"001110101",
  5718=>"010100001",
  5719=>"101111100",
  5720=>"111111011",
  5721=>"001001001",
  5722=>"101000111",
  5723=>"111110110",
  5724=>"001011101",
  5725=>"000011110",
  5726=>"010100101",
  5727=>"011000110",
  5728=>"100110111",
  5729=>"011010010",
  5730=>"011010100",
  5731=>"011010000",
  5732=>"011011000",
  5733=>"100011111",
  5734=>"011111010",
  5735=>"010111111",
  5736=>"001100011",
  5737=>"010111101",
  5738=>"010000111",
  5739=>"001111101",
  5740=>"111110010",
  5741=>"001100110",
  5742=>"000110111",
  5743=>"110001110",
  5744=>"010010111",
  5745=>"100001010",
  5746=>"101010110",
  5747=>"010110101",
  5748=>"110001110",
  5749=>"010100011",
  5750=>"101011000",
  5751=>"101010101",
  5752=>"101011010",
  5753=>"010010010",
  5754=>"100000010",
  5755=>"111100011",
  5756=>"110010000",
  5757=>"101101001",
  5758=>"110011000",
  5759=>"011011111",
  5760=>"110000101",
  5761=>"101001101",
  5762=>"101111001",
  5763=>"110100111",
  5764=>"001100110",
  5765=>"100011001",
  5766=>"101000000",
  5767=>"010100101",
  5768=>"110001000",
  5769=>"010000101",
  5770=>"011011010",
  5771=>"010000011",
  5772=>"000011110",
  5773=>"011101111",
  5774=>"011100101",
  5775=>"110010111",
  5776=>"001101101",
  5777=>"111100010",
  5778=>"011010010",
  5779=>"110100011",
  5780=>"110111000",
  5781=>"110001110",
  5782=>"011000010",
  5783=>"111110100",
  5784=>"110000101",
  5785=>"101100000",
  5786=>"011110000",
  5787=>"101011000",
  5788=>"011111011",
  5789=>"101100000",
  5790=>"010011011",
  5791=>"001000100",
  5792=>"111001111",
  5793=>"000000111",
  5794=>"001000111",
  5795=>"100101110",
  5796=>"011110001",
  5797=>"000011011",
  5798=>"000100111",
  5799=>"101111111",
  5800=>"111001111",
  5801=>"010010111",
  5802=>"100101010",
  5803=>"101010101",
  5804=>"110000001",
  5805=>"110011011",
  5806=>"001011001",
  5807=>"010001011",
  5808=>"110000010",
  5809=>"101000010",
  5810=>"010010011",
  5811=>"100110001",
  5812=>"111101110",
  5813=>"100001000",
  5814=>"001100000",
  5815=>"111000101",
  5816=>"100101000",
  5817=>"101010011",
  5818=>"010001010",
  5819=>"010100001",
  5820=>"101000101",
  5821=>"000100110",
  5822=>"110001010",
  5823=>"000101001",
  5824=>"111100111",
  5825=>"010100110",
  5826=>"000000110",
  5827=>"111000010",
  5828=>"010110001",
  5829=>"000011111",
  5830=>"101110000",
  5831=>"110000010",
  5832=>"011000101",
  5833=>"110001100",
  5834=>"111001111",
  5835=>"110000110",
  5836=>"101111001",
  5837=>"110001001",
  5838=>"110010111",
  5839=>"011011011",
  5840=>"010010110",
  5841=>"011111111",
  5842=>"110111001",
  5843=>"100010101",
  5844=>"000010111",
  5845=>"011110000",
  5846=>"110110110",
  5847=>"100101100",
  5848=>"111101101",
  5849=>"000000111",
  5850=>"010001001",
  5851=>"011111100",
  5852=>"100000110",
  5853=>"111101101",
  5854=>"001010011",
  5855=>"100011000",
  5856=>"101011001",
  5857=>"010100010",
  5858=>"011010011",
  5859=>"110010010",
  5860=>"011101011",
  5861=>"101111100",
  5862=>"111101101",
  5863=>"000010100",
  5864=>"000010010",
  5865=>"111110111",
  5866=>"100101110",
  5867=>"111011010",
  5868=>"101001000",
  5869=>"010001000",
  5870=>"100001100",
  5871=>"000110011",
  5872=>"010000100",
  5873=>"101111011",
  5874=>"110101010",
  5875=>"101001111",
  5876=>"001100101",
  5877=>"101111111",
  5878=>"010000010",
  5879=>"001110110",
  5880=>"101011000",
  5881=>"111010011",
  5882=>"110110111",
  5883=>"000100101",
  5884=>"111101111",
  5885=>"110001001",
  5886=>"101001001",
  5887=>"100110000",
  5888=>"010110001",
  5889=>"111101001",
  5890=>"001011111",
  5891=>"100000101",
  5892=>"101000001",
  5893=>"110110000",
  5894=>"010100000",
  5895=>"010011010",
  5896=>"110010111",
  5897=>"100101011",
  5898=>"101100000",
  5899=>"000010101",
  5900=>"111101101",
  5901=>"001001100",
  5902=>"000001011",
  5903=>"111001011",
  5904=>"100100101",
  5905=>"000101011",
  5906=>"100011000",
  5907=>"110101101",
  5908=>"010111001",
  5909=>"001100110",
  5910=>"110110101",
  5911=>"101101100",
  5912=>"000101001",
  5913=>"000000101",
  5914=>"100011000",
  5915=>"100101010",
  5916=>"100101111",
  5917=>"011011101",
  5918=>"000000100",
  5919=>"000100000",
  5920=>"010001001",
  5921=>"011110100",
  5922=>"010000110",
  5923=>"100110000",
  5924=>"000101100",
  5925=>"111100011",
  5926=>"100100010",
  5927=>"011000100",
  5928=>"011000101",
  5929=>"000100100",
  5930=>"001101111",
  5931=>"100011100",
  5932=>"011100011",
  5933=>"111101101",
  5934=>"001001001",
  5935=>"010111010",
  5936=>"011100001",
  5937=>"111100001",
  5938=>"000011111",
  5939=>"010000011",
  5940=>"001001011",
  5941=>"101011110",
  5942=>"101010110",
  5943=>"010100111",
  5944=>"010111100",
  5945=>"010000001",
  5946=>"011110111",
  5947=>"001100100",
  5948=>"110101110",
  5949=>"000100110",
  5950=>"011111100",
  5951=>"100000000",
  5952=>"110110111",
  5953=>"000000000",
  5954=>"110010011",
  5955=>"001111010",
  5956=>"010011110",
  5957=>"010110111",
  5958=>"001011110",
  5959=>"001001100",
  5960=>"000000010",
  5961=>"011100001",
  5962=>"000011100",
  5963=>"001001000",
  5964=>"110110110",
  5965=>"000101011",
  5966=>"011010110",
  5967=>"100101001",
  5968=>"000001100",
  5969=>"111000100",
  5970=>"011000001",
  5971=>"000100010",
  5972=>"011001110",
  5973=>"001001111",
  5974=>"000101000",
  5975=>"111011011",
  5976=>"111011111",
  5977=>"111010111",
  5978=>"011010011",
  5979=>"100101001",
  5980=>"000111101",
  5981=>"010100010",
  5982=>"101000100",
  5983=>"000101001",
  5984=>"011111000",
  5985=>"101110110",
  5986=>"000110101",
  5987=>"110110111",
  5988=>"000011011",
  5989=>"000011000",
  5990=>"101101011",
  5991=>"000000110",
  5992=>"111111101",
  5993=>"110001001",
  5994=>"101001110",
  5995=>"011011110",
  5996=>"001000001",
  5997=>"001001000",
  5998=>"011111100",
  5999=>"010100010",
  6000=>"010101111",
  6001=>"101101101",
  6002=>"011111110",
  6003=>"101011011",
  6004=>"001110111",
  6005=>"111011001",
  6006=>"110110110",
  6007=>"001011011",
  6008=>"000101111",
  6009=>"111001101",
  6010=>"100101010",
  6011=>"110001111",
  6012=>"100011010",
  6013=>"000100111",
  6014=>"101100000",
  6015=>"000010001",
  6016=>"000001111",
  6017=>"011110100",
  6018=>"101001111",
  6019=>"111000110",
  6020=>"000100000",
  6021=>"011100100",
  6022=>"110000011",
  6023=>"000000101",
  6024=>"110011010",
  6025=>"001111101",
  6026=>"001110111",
  6027=>"000001111",
  6028=>"010100011",
  6029=>"010110101",
  6030=>"110000011",
  6031=>"000100101",
  6032=>"100110111",
  6033=>"001101100",
  6034=>"011010111",
  6035=>"000001101",
  6036=>"001101110",
  6037=>"100100110",
  6038=>"101010010",
  6039=>"010011111",
  6040=>"111101110",
  6041=>"000000101",
  6042=>"110001000",
  6043=>"110101011",
  6044=>"000001101",
  6045=>"000100000",
  6046=>"100000000",
  6047=>"001100001",
  6048=>"011011110",
  6049=>"011110011",
  6050=>"001100101",
  6051=>"100101111",
  6052=>"000111000",
  6053=>"111101111",
  6054=>"000000100",
  6055=>"111000111",
  6056=>"000000011",
  6057=>"111001010",
  6058=>"000100010",
  6059=>"110001100",
  6060=>"010101001",
  6061=>"001010101",
  6062=>"110110010",
  6063=>"110001011",
  6064=>"100101000",
  6065=>"001001110",
  6066=>"100100000",
  6067=>"001000000",
  6068=>"111111110",
  6069=>"001000100",
  6070=>"100001101",
  6071=>"101011000",
  6072=>"000001010",
  6073=>"010001100",
  6074=>"111011000",
  6075=>"011111000",
  6076=>"100101010",
  6077=>"111110000",
  6078=>"010011001",
  6079=>"001000101",
  6080=>"001000001",
  6081=>"001110101",
  6082=>"110011001",
  6083=>"011110001",
  6084=>"001110100",
  6085=>"001000011",
  6086=>"100111101",
  6087=>"111110011",
  6088=>"101101000",
  6089=>"110111100",
  6090=>"001001110",
  6091=>"110111000",
  6092=>"111111101",
  6093=>"011101111",
  6094=>"101100111",
  6095=>"100110111",
  6096=>"001101111",
  6097=>"000100111",
  6098=>"101001011",
  6099=>"010110101",
  6100=>"111010111",
  6101=>"010100010",
  6102=>"110101101",
  6103=>"110000001",
  6104=>"011111101",
  6105=>"110000110",
  6106=>"110000110",
  6107=>"110010000",
  6108=>"101111101",
  6109=>"010000011",
  6110=>"000101010",
  6111=>"101111111",
  6112=>"010111010",
  6113=>"100010011",
  6114=>"011111001",
  6115=>"010011010",
  6116=>"000111101",
  6117=>"000111000",
  6118=>"000010011",
  6119=>"010100111",
  6120=>"101010111",
  6121=>"001101001",
  6122=>"101000011",
  6123=>"011111110",
  6124=>"001010000",
  6125=>"010011010",
  6126=>"101111110",
  6127=>"000110011",
  6128=>"010101010",
  6129=>"010010010",
  6130=>"101000010",
  6131=>"100101100",
  6132=>"111110010",
  6133=>"010111000",
  6134=>"110010011",
  6135=>"010000111",
  6136=>"000010110",
  6137=>"111110110",
  6138=>"011000101",
  6139=>"001000110",
  6140=>"000010111",
  6141=>"010110000",
  6142=>"100101101",
  6143=>"100101001",
  6144=>"111010000",
  6145=>"010011101",
  6146=>"010000001",
  6147=>"000001100",
  6148=>"011000111",
  6149=>"001011010",
  6150=>"000011011",
  6151=>"010010010",
  6152=>"001010011",
  6153=>"101100011",
  6154=>"001001010",
  6155=>"010101000",
  6156=>"110000001",
  6157=>"000010011",
  6158=>"100111011",
  6159=>"010101110",
  6160=>"000010001",
  6161=>"101110111",
  6162=>"110100110",
  6163=>"010000000",
  6164=>"010000100",
  6165=>"011110000",
  6166=>"010100010",
  6167=>"111000101",
  6168=>"001001000",
  6169=>"001010111",
  6170=>"111111010",
  6171=>"111111010",
  6172=>"111110110",
  6173=>"101111110",
  6174=>"000001100",
  6175=>"110100101",
  6176=>"111010000",
  6177=>"111000010",
  6178=>"111001100",
  6179=>"110011010",
  6180=>"011000001",
  6181=>"011110100",
  6182=>"100101100",
  6183=>"101110001",
  6184=>"111001000",
  6185=>"010011001",
  6186=>"110110000",
  6187=>"100101011",
  6188=>"111111000",
  6189=>"110100111",
  6190=>"001011111",
  6191=>"001010110",
  6192=>"110110000",
  6193=>"110111100",
  6194=>"110100001",
  6195=>"100010100",
  6196=>"111011001",
  6197=>"111011011",
  6198=>"011011111",
  6199=>"101101001",
  6200=>"001011101",
  6201=>"001010110",
  6202=>"101101110",
  6203=>"001011111",
  6204=>"111000001",
  6205=>"111001010",
  6206=>"101110010",
  6207=>"010101000",
  6208=>"111010011",
  6209=>"100110110",
  6210=>"001010001",
  6211=>"010100110",
  6212=>"110010110",
  6213=>"001000011",
  6214=>"100111001",
  6215=>"110110111",
  6216=>"010011000",
  6217=>"110110100",
  6218=>"010000101",
  6219=>"101000100",
  6220=>"000010011",
  6221=>"101101011",
  6222=>"100100010",
  6223=>"100100011",
  6224=>"000111110",
  6225=>"111100111",
  6226=>"101100100",
  6227=>"000110011",
  6228=>"010000010",
  6229=>"000001011",
  6230=>"011110110",
  6231=>"101001100",
  6232=>"111011001",
  6233=>"100111001",
  6234=>"110101110",
  6235=>"101100100",
  6236=>"001110101",
  6237=>"101101001",
  6238=>"101111110",
  6239=>"000101001",
  6240=>"000010000",
  6241=>"111111111",
  6242=>"101101110",
  6243=>"000000010",
  6244=>"111111010",
  6245=>"000010111",
  6246=>"001101100",
  6247=>"010110001",
  6248=>"011100100",
  6249=>"101110001",
  6250=>"100010001",
  6251=>"000010100",
  6252=>"011011100",
  6253=>"001100001",
  6254=>"100000001",
  6255=>"001100000",
  6256=>"000101001",
  6257=>"010100001",
  6258=>"101110111",
  6259=>"110011000",
  6260=>"001001001",
  6261=>"000110100",
  6262=>"000000000",
  6263=>"011100100",
  6264=>"001111011",
  6265=>"111110000",
  6266=>"101101000",
  6267=>"110111010",
  6268=>"110011110",
  6269=>"110001001",
  6270=>"010000100",
  6271=>"010100101",
  6272=>"000100111",
  6273=>"011010001",
  6274=>"011100100",
  6275=>"111101010",
  6276=>"111111111",
  6277=>"111011001",
  6278=>"110111100",
  6279=>"110110001",
  6280=>"111010101",
  6281=>"000011011",
  6282=>"001110001",
  6283=>"010000100",
  6284=>"000001010",
  6285=>"000110100",
  6286=>"100111000",
  6287=>"110100001",
  6288=>"011111000",
  6289=>"111110110",
  6290=>"110110000",
  6291=>"111000111",
  6292=>"010100100",
  6293=>"001011010",
  6294=>"001101101",
  6295=>"101011110",
  6296=>"000110110",
  6297=>"101011011",
  6298=>"100100100",
  6299=>"001010011",
  6300=>"100110000",
  6301=>"101000010",
  6302=>"101101011",
  6303=>"000110010",
  6304=>"100000011",
  6305=>"010001101",
  6306=>"010011011",
  6307=>"100100110",
  6308=>"101010101",
  6309=>"001010110",
  6310=>"011101111",
  6311=>"011001101",
  6312=>"011001000",
  6313=>"110010011",
  6314=>"100110111",
  6315=>"111001101",
  6316=>"000111101",
  6317=>"100101100",
  6318=>"110100000",
  6319=>"111100110",
  6320=>"010011100",
  6321=>"010111011",
  6322=>"000110000",
  6323=>"110100111",
  6324=>"001001100",
  6325=>"100011101",
  6326=>"011101001",
  6327=>"010101100",
  6328=>"101110010",
  6329=>"001110001",
  6330=>"111111011",
  6331=>"011111110",
  6332=>"110101011",
  6333=>"100101101",
  6334=>"011010100",
  6335=>"101101011",
  6336=>"101010111",
  6337=>"101101010",
  6338=>"100111100",
  6339=>"001000011",
  6340=>"100011111",
  6341=>"010001001",
  6342=>"110001011",
  6343=>"000011101",
  6344=>"010010111",
  6345=>"101011101",
  6346=>"111011100",
  6347=>"100110111",
  6348=>"110011100",
  6349=>"011000100",
  6350=>"101001110",
  6351=>"101111111",
  6352=>"111001001",
  6353=>"111110010",
  6354=>"100000010",
  6355=>"100001111",
  6356=>"111101111",
  6357=>"011010110",
  6358=>"111011000",
  6359=>"011000101",
  6360=>"100000010",
  6361=>"101101101",
  6362=>"011011010",
  6363=>"111001100",
  6364=>"110111111",
  6365=>"101000010",
  6366=>"111000011",
  6367=>"000101101",
  6368=>"000111000",
  6369=>"101101111",
  6370=>"000111100",
  6371=>"101001111",
  6372=>"001010010",
  6373=>"101000101",
  6374=>"010000011",
  6375=>"110010110",
  6376=>"111010010",
  6377=>"001010000",
  6378=>"001000001",
  6379=>"101101100",
  6380=>"111001101",
  6381=>"010001111",
  6382=>"000010110",
  6383=>"111101111",
  6384=>"010001000",
  6385=>"101101101",
  6386=>"100010010",
  6387=>"001110110",
  6388=>"111011000",
  6389=>"011110110",
  6390=>"100111000",
  6391=>"101001100",
  6392=>"100010011",
  6393=>"000111100",
  6394=>"110101111",
  6395=>"100101001",
  6396=>"000010011",
  6397=>"100101011",
  6398=>"110101001",
  6399=>"000111011",
  6400=>"010111111",
  6401=>"111010110",
  6402=>"100101100",
  6403=>"100001101",
  6404=>"000110000",
  6405=>"111010010",
  6406=>"010001010",
  6407=>"101011111",
  6408=>"101011010",
  6409=>"001101010",
  6410=>"001010111",
  6411=>"100001110",
  6412=>"110110111",
  6413=>"000010000",
  6414=>"011011111",
  6415=>"010000110",
  6416=>"101100110",
  6417=>"010000001",
  6418=>"101101000",
  6419=>"110011100",
  6420=>"011011101",
  6421=>"100110001",
  6422=>"001001101",
  6423=>"101011011",
  6424=>"111101001",
  6425=>"011010000",
  6426=>"100000110",
  6427=>"110010100",
  6428=>"000000001",
  6429=>"010101110",
  6430=>"010010011",
  6431=>"010001111",
  6432=>"010001100",
  6433=>"011110000",
  6434=>"010111010",
  6435=>"101010100",
  6436=>"010000101",
  6437=>"101110110",
  6438=>"111101001",
  6439=>"111011100",
  6440=>"100111110",
  6441=>"010011101",
  6442=>"110010000",
  6443=>"010010110",
  6444=>"000111010",
  6445=>"111010100",
  6446=>"010000111",
  6447=>"100111011",
  6448=>"110010100",
  6449=>"001001000",
  6450=>"010010111",
  6451=>"110010011",
  6452=>"111111110",
  6453=>"000000110",
  6454=>"101100010",
  6455=>"111100101",
  6456=>"011011100",
  6457=>"001110010",
  6458=>"101110101",
  6459=>"011010110",
  6460=>"101111001",
  6461=>"010111000",
  6462=>"100111011",
  6463=>"110101100",
  6464=>"001000011",
  6465=>"101111000",
  6466=>"000101100",
  6467=>"111100100",
  6468=>"010000101",
  6469=>"010111101",
  6470=>"111110010",
  6471=>"110111100",
  6472=>"011000000",
  6473=>"110001001",
  6474=>"011100000",
  6475=>"000100011",
  6476=>"111110000",
  6477=>"101011000",
  6478=>"111111100",
  6479=>"110101001",
  6480=>"110101110",
  6481=>"001001100",
  6482=>"111010111",
  6483=>"001110011",
  6484=>"000000000",
  6485=>"111111010",
  6486=>"010110101",
  6487=>"011111011",
  6488=>"100001000",
  6489=>"111100110",
  6490=>"011100100",
  6491=>"100010001",
  6492=>"001001101",
  6493=>"001000001",
  6494=>"011101100",
  6495=>"000100110",
  6496=>"011111101",
  6497=>"101000001",
  6498=>"111100111",
  6499=>"000111011",
  6500=>"000111010",
  6501=>"100000010",
  6502=>"010101001",
  6503=>"110010111",
  6504=>"001101011",
  6505=>"011101100",
  6506=>"000011000",
  6507=>"010100010",
  6508=>"001001001",
  6509=>"111100011",
  6510=>"011111101",
  6511=>"011111010",
  6512=>"011010011",
  6513=>"010010001",
  6514=>"100101100",
  6515=>"111101000",
  6516=>"001111010",
  6517=>"011001001",
  6518=>"010101100",
  6519=>"000111010",
  6520=>"011000001",
  6521=>"110001110",
  6522=>"000001111",
  6523=>"000110000",
  6524=>"100111100",
  6525=>"111111111",
  6526=>"100011000",
  6527=>"111101001",
  6528=>"011011011",
  6529=>"100000001",
  6530=>"111001111",
  6531=>"000001000",
  6532=>"111101110",
  6533=>"101111100",
  6534=>"010000011",
  6535=>"110011000",
  6536=>"001000010",
  6537=>"100111110",
  6538=>"101000011",
  6539=>"000001100",
  6540=>"111100011",
  6541=>"100101100",
  6542=>"110110111",
  6543=>"111100101",
  6544=>"100100110",
  6545=>"001100100",
  6546=>"000111011",
  6547=>"100000010",
  6548=>"110101110",
  6549=>"000000000",
  6550=>"011100000",
  6551=>"011100000",
  6552=>"010011100",
  6553=>"011110111",
  6554=>"111101001",
  6555=>"101100100",
  6556=>"111000110",
  6557=>"001101010",
  6558=>"100011001",
  6559=>"101100101",
  6560=>"100101111",
  6561=>"000000110",
  6562=>"101011110",
  6563=>"000110011",
  6564=>"101110001",
  6565=>"101111001",
  6566=>"010000110",
  6567=>"011110101",
  6568=>"001100111",
  6569=>"010101100",
  6570=>"011011000",
  6571=>"000001001",
  6572=>"110110111",
  6573=>"111111010",
  6574=>"111111111",
  6575=>"100110000",
  6576=>"111000000",
  6577=>"001001001",
  6578=>"100101110",
  6579=>"011011101",
  6580=>"011011000",
  6581=>"000001111",
  6582=>"110100001",
  6583=>"001110000",
  6584=>"000111111",
  6585=>"001011101",
  6586=>"001000010",
  6587=>"101100111",
  6588=>"010001000",
  6589=>"101111101",
  6590=>"101111001",
  6591=>"001010001",
  6592=>"110110000",
  6593=>"010110000",
  6594=>"001010111",
  6595=>"010111011",
  6596=>"000001101",
  6597=>"010111000",
  6598=>"010011000",
  6599=>"110100111",
  6600=>"111111000",
  6601=>"010101100",
  6602=>"101000010",
  6603=>"110101101",
  6604=>"010011101",
  6605=>"001010010",
  6606=>"001100001",
  6607=>"111111000",
  6608=>"001101101",
  6609=>"001011100",
  6610=>"010110111",
  6611=>"010111011",
  6612=>"010111000",
  6613=>"000111111",
  6614=>"110111000",
  6615=>"000010001",
  6616=>"110010000",
  6617=>"010001110",
  6618=>"111000010",
  6619=>"010111100",
  6620=>"110010000",
  6621=>"010110111",
  6622=>"000010000",
  6623=>"010110011",
  6624=>"001111001",
  6625=>"110010111",
  6626=>"101100000",
  6627=>"001110101",
  6628=>"111000010",
  6629=>"110110111",
  6630=>"011000000",
  6631=>"011101101",
  6632=>"010000100",
  6633=>"111100101",
  6634=>"011011111",
  6635=>"010000111",
  6636=>"001000001",
  6637=>"110111011",
  6638=>"111110000",
  6639=>"010100101",
  6640=>"001100000",
  6641=>"110101101",
  6642=>"001111111",
  6643=>"001100001",
  6644=>"100001001",
  6645=>"010111100",
  6646=>"001001000",
  6647=>"111111110",
  6648=>"010011000",
  6649=>"110000101",
  6650=>"111000101",
  6651=>"010001001",
  6652=>"000001101",
  6653=>"000101100",
  6654=>"001100111",
  6655=>"101000111",
  6656=>"100101101",
  6657=>"110010111",
  6658=>"011101111",
  6659=>"100010001",
  6660=>"001001001",
  6661=>"100101000",
  6662=>"111111001",
  6663=>"010011001",
  6664=>"011110000",
  6665=>"001000011",
  6666=>"010001011",
  6667=>"101000001",
  6668=>"110001111",
  6669=>"000000001",
  6670=>"100101000",
  6671=>"110100100",
  6672=>"000000000",
  6673=>"011111000",
  6674=>"010111100",
  6675=>"100000001",
  6676=>"100001101",
  6677=>"000101010",
  6678=>"011011100",
  6679=>"100100101",
  6680=>"101111110",
  6681=>"010110101",
  6682=>"011010001",
  6683=>"101010101",
  6684=>"100000000",
  6685=>"000010001",
  6686=>"100001001",
  6687=>"000010111",
  6688=>"100000010",
  6689=>"010001111",
  6690=>"010000000",
  6691=>"001110100",
  6692=>"000011010",
  6693=>"001011011",
  6694=>"100100000",
  6695=>"111111001",
  6696=>"110110110",
  6697=>"100110101",
  6698=>"001001000",
  6699=>"001110110",
  6700=>"000000111",
  6701=>"001111111",
  6702=>"111011101",
  6703=>"000000001",
  6704=>"011000011",
  6705=>"011100001",
  6706=>"001000111",
  6707=>"011010110",
  6708=>"000000100",
  6709=>"010100111",
  6710=>"100011100",
  6711=>"010101000",
  6712=>"000001101",
  6713=>"110111110",
  6714=>"110010110",
  6715=>"011001000",
  6716=>"100110001",
  6717=>"111100110",
  6718=>"011101001",
  6719=>"110000000",
  6720=>"101011010",
  6721=>"110011001",
  6722=>"001000001",
  6723=>"111110010",
  6724=>"101110100",
  6725=>"000110111",
  6726=>"001110101",
  6727=>"011011000",
  6728=>"110111011",
  6729=>"101100101",
  6730=>"110100001",
  6731=>"000100101",
  6732=>"101111110",
  6733=>"000001101",
  6734=>"011110001",
  6735=>"001000111",
  6736=>"110000000",
  6737=>"100000000",
  6738=>"100111011",
  6739=>"000000100",
  6740=>"111010100",
  6741=>"010011100",
  6742=>"001010001",
  6743=>"010010001",
  6744=>"000101000",
  6745=>"111001001",
  6746=>"111001101",
  6747=>"111111100",
  6748=>"111000000",
  6749=>"111000010",
  6750=>"101100111",
  6751=>"000101001",
  6752=>"111001110",
  6753=>"011010011",
  6754=>"100111101",
  6755=>"111000001",
  6756=>"110110101",
  6757=>"010100111",
  6758=>"010101011",
  6759=>"111011111",
  6760=>"010011101",
  6761=>"011000011",
  6762=>"100110000",
  6763=>"001100101",
  6764=>"000010110",
  6765=>"001101011",
  6766=>"001000010",
  6767=>"111001100",
  6768=>"101111101",
  6769=>"001011101",
  6770=>"111010011",
  6771=>"001010001",
  6772=>"000001111",
  6773=>"101001100",
  6774=>"001101111",
  6775=>"001001000",
  6776=>"101100110",
  6777=>"100000000",
  6778=>"001001100",
  6779=>"100000101",
  6780=>"110011111",
  6781=>"000000001",
  6782=>"011010111",
  6783=>"010111010",
  6784=>"000010000",
  6785=>"101011110",
  6786=>"000001000",
  6787=>"000001101",
  6788=>"010000101",
  6789=>"000001010",
  6790=>"000101011",
  6791=>"010111011",
  6792=>"000100010",
  6793=>"111011001",
  6794=>"000111010",
  6795=>"111100011",
  6796=>"101110101",
  6797=>"110011111",
  6798=>"110110111",
  6799=>"010010100",
  6800=>"100110111",
  6801=>"000110110",
  6802=>"011011111",
  6803=>"010110001",
  6804=>"111000111",
  6805=>"011000010",
  6806=>"110011011",
  6807=>"111101010",
  6808=>"000011111",
  6809=>"010111111",
  6810=>"100000010",
  6811=>"010001000",
  6812=>"011011000",
  6813=>"010011001",
  6814=>"000010011",
  6815=>"100100100",
  6816=>"110100010",
  6817=>"100111010",
  6818=>"000000001",
  6819=>"101101010",
  6820=>"000001000",
  6821=>"000100111",
  6822=>"011011000",
  6823=>"101110001",
  6824=>"110000011",
  6825=>"111101000",
  6826=>"011100101",
  6827=>"100101100",
  6828=>"010110000",
  6829=>"011000111",
  6830=>"001110111",
  6831=>"110010010",
  6832=>"000100111",
  6833=>"010010100",
  6834=>"011010011",
  6835=>"110110011",
  6836=>"110010111",
  6837=>"111000101",
  6838=>"011001000",
  6839=>"010101011",
  6840=>"011001101",
  6841=>"110001001",
  6842=>"110010111",
  6843=>"101001111",
  6844=>"010111010",
  6845=>"000100000",
  6846=>"100110111",
  6847=>"101110110",
  6848=>"111110111",
  6849=>"000100111",
  6850=>"000011011",
  6851=>"101101100",
  6852=>"110010000",
  6853=>"100010101",
  6854=>"101011000",
  6855=>"110010100",
  6856=>"111010100",
  6857=>"010011010",
  6858=>"011011110",
  6859=>"100001111",
  6860=>"001011101",
  6861=>"000000101",
  6862=>"011110001",
  6863=>"000100111",
  6864=>"101001011",
  6865=>"110110110",
  6866=>"110010111",
  6867=>"001001000",
  6868=>"010010000",
  6869=>"110110001",
  6870=>"100101001",
  6871=>"010110111",
  6872=>"010111101",
  6873=>"101101010",
  6874=>"010000001",
  6875=>"100000010",
  6876=>"101101101",
  6877=>"100000011",
  6878=>"001100110",
  6879=>"001110101",
  6880=>"101000101",
  6881=>"001110100",
  6882=>"100101110",
  6883=>"000101010",
  6884=>"100111000",
  6885=>"111111001",
  6886=>"110111010",
  6887=>"000011110",
  6888=>"100100001",
  6889=>"101001101",
  6890=>"010100110",
  6891=>"011100000",
  6892=>"101000010",
  6893=>"101010101",
  6894=>"101010001",
  6895=>"001110000",
  6896=>"101110001",
  6897=>"010000111",
  6898=>"010111111",
  6899=>"111101111",
  6900=>"101111110",
  6901=>"011000010",
  6902=>"001101111",
  6903=>"011100101",
  6904=>"111100000",
  6905=>"100001001",
  6906=>"101110111",
  6907=>"111001011",
  6908=>"001000111",
  6909=>"011000101",
  6910=>"110000010",
  6911=>"010101111",
  6912=>"111010111",
  6913=>"000110011",
  6914=>"111001000",
  6915=>"110100010",
  6916=>"010110111",
  6917=>"000001000",
  6918=>"000000010",
  6919=>"100110100",
  6920=>"100001110",
  6921=>"000001111",
  6922=>"101100111",
  6923=>"000000001",
  6924=>"000011100",
  6925=>"100100111",
  6926=>"010010000",
  6927=>"111010000",
  6928=>"000001110",
  6929=>"001010100",
  6930=>"001111001",
  6931=>"100101011",
  6932=>"101001101",
  6933=>"111110101",
  6934=>"010001011",
  6935=>"111011111",
  6936=>"111001111",
  6937=>"100100101",
  6938=>"000010100",
  6939=>"110001000",
  6940=>"100011111",
  6941=>"001110110",
  6942=>"110001100",
  6943=>"000101100",
  6944=>"011000010",
  6945=>"001000010",
  6946=>"000011001",
  6947=>"011111011",
  6948=>"111110101",
  6949=>"110111011",
  6950=>"101001100",
  6951=>"011000100",
  6952=>"010101011",
  6953=>"110000001",
  6954=>"010000001",
  6955=>"001001101",
  6956=>"000000111",
  6957=>"000001011",
  6958=>"000001011",
  6959=>"111100011",
  6960=>"101000001",
  6961=>"000011010",
  6962=>"100111011",
  6963=>"110100100",
  6964=>"111111011",
  6965=>"110110100",
  6966=>"111110101",
  6967=>"001111110",
  6968=>"011111000",
  6969=>"101110001",
  6970=>"000110110",
  6971=>"101011100",
  6972=>"100001111",
  6973=>"001110001",
  6974=>"000100111",
  6975=>"001000000",
  6976=>"000001000",
  6977=>"100011000",
  6978=>"011000100",
  6979=>"111100010",
  6980=>"101011111",
  6981=>"001101101",
  6982=>"100010110",
  6983=>"001000101",
  6984=>"101001000",
  6985=>"011101001",
  6986=>"001100011",
  6987=>"000000001",
  6988=>"110111011",
  6989=>"100000001",
  6990=>"111100111",
  6991=>"110010011",
  6992=>"011111100",
  6993=>"110101111",
  6994=>"111111001",
  6995=>"001111110",
  6996=>"001011010",
  6997=>"101110100",
  6998=>"000110111",
  6999=>"111101000",
  7000=>"000001000",
  7001=>"101111000",
  7002=>"001100001",
  7003=>"101000101",
  7004=>"000100001",
  7005=>"010110011",
  7006=>"100111100",
  7007=>"000101000",
  7008=>"000010001",
  7009=>"111011011",
  7010=>"100000010",
  7011=>"011001101",
  7012=>"110111101",
  7013=>"001101000",
  7014=>"111001110",
  7015=>"100001111",
  7016=>"111110110",
  7017=>"001101101",
  7018=>"110100010",
  7019=>"101110000",
  7020=>"101110100",
  7021=>"000110100",
  7022=>"010100101",
  7023=>"100110011",
  7024=>"001001101",
  7025=>"100001110",
  7026=>"010111101",
  7027=>"001001110",
  7028=>"000100000",
  7029=>"100100101",
  7030=>"111100100",
  7031=>"111000010",
  7032=>"101011001",
  7033=>"011101110",
  7034=>"110001011",
  7035=>"011101011",
  7036=>"010000001",
  7037=>"011011100",
  7038=>"001011101",
  7039=>"110011110",
  7040=>"100100000",
  7041=>"100010011",
  7042=>"010011100",
  7043=>"110100011",
  7044=>"000001100",
  7045=>"100111100",
  7046=>"000110010",
  7047=>"100110100",
  7048=>"010101101",
  7049=>"111011111",
  7050=>"000011010",
  7051=>"110110010",
  7052=>"010100110",
  7053=>"001001111",
  7054=>"111110000",
  7055=>"011100110",
  7056=>"101111100",
  7057=>"100110010",
  7058=>"100111101",
  7059=>"011101100",
  7060=>"111001011",
  7061=>"111111000",
  7062=>"101100001",
  7063=>"001110010",
  7064=>"000111111",
  7065=>"111111111",
  7066=>"000010100",
  7067=>"001111111",
  7068=>"100101101",
  7069=>"000000001",
  7070=>"110111110",
  7071=>"001001110",
  7072=>"010110010",
  7073=>"101101111",
  7074=>"010101101",
  7075=>"011000100",
  7076=>"000011001",
  7077=>"011100110",
  7078=>"000000110",
  7079=>"011011101",
  7080=>"001001001",
  7081=>"101101010",
  7082=>"000111001",
  7083=>"111100001",
  7084=>"110100011",
  7085=>"000001000",
  7086=>"000100010",
  7087=>"111111011",
  7088=>"011010101",
  7089=>"001010001",
  7090=>"111111110",
  7091=>"000010010",
  7092=>"011100100",
  7093=>"000111011",
  7094=>"100011100",
  7095=>"000111011",
  7096=>"101101101",
  7097=>"100001000",
  7098=>"001000111",
  7099=>"100111111",
  7100=>"110101011",
  7101=>"100000000",
  7102=>"100011110",
  7103=>"001010011",
  7104=>"110000001",
  7105=>"010110010",
  7106=>"111011110",
  7107=>"111000000",
  7108=>"111101010",
  7109=>"000011011",
  7110=>"010110001",
  7111=>"100011010",
  7112=>"111100101",
  7113=>"111010100",
  7114=>"110011100",
  7115=>"100000010",
  7116=>"110111011",
  7117=>"111101011",
  7118=>"100011101",
  7119=>"000110101",
  7120=>"100100101",
  7121=>"001000011",
  7122=>"111000110",
  7123=>"100001110",
  7124=>"000111101",
  7125=>"101101011",
  7126=>"100101110",
  7127=>"010010111",
  7128=>"010000110",
  7129=>"100010110",
  7130=>"101011001",
  7131=>"010010011",
  7132=>"111001011",
  7133=>"110001101",
  7134=>"101111010",
  7135=>"101010111",
  7136=>"000000010",
  7137=>"111010011",
  7138=>"111001101",
  7139=>"111001000",
  7140=>"100010111",
  7141=>"110110011",
  7142=>"111001010",
  7143=>"111011110",
  7144=>"100000001",
  7145=>"110000110",
  7146=>"110110111",
  7147=>"000101100",
  7148=>"111001000",
  7149=>"001101000",
  7150=>"010111010",
  7151=>"011110011",
  7152=>"000000001",
  7153=>"101000000",
  7154=>"101000010",
  7155=>"100001110",
  7156=>"110011011",
  7157=>"011010010",
  7158=>"010100011",
  7159=>"000000011",
  7160=>"011111101",
  7161=>"000011000",
  7162=>"111111101",
  7163=>"011000110",
  7164=>"000100111",
  7165=>"000100010",
  7166=>"010011110",
  7167=>"011010111",
  7168=>"101110100",
  7169=>"110010111",
  7170=>"011010010",
  7171=>"111110001",
  7172=>"001001000",
  7173=>"000011101",
  7174=>"011000010",
  7175=>"000011011",
  7176=>"010100011",
  7177=>"001110010",
  7178=>"101100001",
  7179=>"110000101",
  7180=>"100011110",
  7181=>"100010011",
  7182=>"000011011",
  7183=>"111110101",
  7184=>"011111100",
  7185=>"100000000",
  7186=>"011110101",
  7187=>"001101001",
  7188=>"111010101",
  7189=>"110100101",
  7190=>"110110110",
  7191=>"100010001",
  7192=>"010011001",
  7193=>"101001111",
  7194=>"010100100",
  7195=>"110110111",
  7196=>"100001011",
  7197=>"011110100",
  7198=>"011010101",
  7199=>"101111101",
  7200=>"110011101",
  7201=>"100000111",
  7202=>"101001010",
  7203=>"011101000",
  7204=>"011001001",
  7205=>"001010100",
  7206=>"000100110",
  7207=>"111000101",
  7208=>"000010110",
  7209=>"101001110",
  7210=>"101011110",
  7211=>"000110110",
  7212=>"011011111",
  7213=>"111011000",
  7214=>"100001000",
  7215=>"100101000",
  7216=>"000111000",
  7217=>"101001100",
  7218=>"001001111",
  7219=>"010100000",
  7220=>"100100000",
  7221=>"011111010",
  7222=>"100111110",
  7223=>"010111010",
  7224=>"000001101",
  7225=>"101100001",
  7226=>"101101001",
  7227=>"100100001",
  7228=>"111100010",
  7229=>"110111001",
  7230=>"101001001",
  7231=>"001001001",
  7232=>"110100111",
  7233=>"010010100",
  7234=>"100011010",
  7235=>"110011101",
  7236=>"101101100",
  7237=>"000111101",
  7238=>"100100011",
  7239=>"101001000",
  7240=>"110011100",
  7241=>"001100100",
  7242=>"000111101",
  7243=>"111101001",
  7244=>"010101011",
  7245=>"111110110",
  7246=>"010000100",
  7247=>"111110101",
  7248=>"010101111",
  7249=>"111101101",
  7250=>"010110100",
  7251=>"110000100",
  7252=>"010010110",
  7253=>"110100001",
  7254=>"110110000",
  7255=>"010001001",
  7256=>"000100101",
  7257=>"101000110",
  7258=>"111100111",
  7259=>"100101111",
  7260=>"100111111",
  7261=>"000100011",
  7262=>"110010101",
  7263=>"001001111",
  7264=>"000011101",
  7265=>"101100100",
  7266=>"101111000",
  7267=>"111100000",
  7268=>"110110000",
  7269=>"100110101",
  7270=>"001101111",
  7271=>"001000010",
  7272=>"000111110",
  7273=>"100111101",
  7274=>"001101000",
  7275=>"111111001",
  7276=>"100001010",
  7277=>"001110100",
  7278=>"111100100",
  7279=>"111111110",
  7280=>"000001110",
  7281=>"111000110",
  7282=>"011001110",
  7283=>"101001011",
  7284=>"011100010",
  7285=>"100101011",
  7286=>"010011101",
  7287=>"100000000",
  7288=>"110110011",
  7289=>"101101000",
  7290=>"100001111",
  7291=>"010101101",
  7292=>"000000111",
  7293=>"010111011",
  7294=>"000110110",
  7295=>"111111011",
  7296=>"010110011",
  7297=>"101000100",
  7298=>"011100001",
  7299=>"100010110",
  7300=>"011000010",
  7301=>"100010100",
  7302=>"011010111",
  7303=>"111110101",
  7304=>"110000010",
  7305=>"110111110",
  7306=>"100101011",
  7307=>"111001100",
  7308=>"111000100",
  7309=>"110011001",
  7310=>"001011100",
  7311=>"111100111",
  7312=>"011001100",
  7313=>"010101000",
  7314=>"111001111",
  7315=>"111011011",
  7316=>"000110100",
  7317=>"000101111",
  7318=>"001000101",
  7319=>"000000101",
  7320=>"110011100",
  7321=>"010001101",
  7322=>"000101001",
  7323=>"101000101",
  7324=>"010010110",
  7325=>"111111100",
  7326=>"010011101",
  7327=>"110011100",
  7328=>"100010001",
  7329=>"000010111",
  7330=>"111001110",
  7331=>"000000010",
  7332=>"101000111",
  7333=>"001111110",
  7334=>"010101100",
  7335=>"010101010",
  7336=>"001011100",
  7337=>"000110100",
  7338=>"111101011",
  7339=>"011010101",
  7340=>"100011110",
  7341=>"100001110",
  7342=>"000000100",
  7343=>"001111001",
  7344=>"110111101",
  7345=>"111001010",
  7346=>"110011010",
  7347=>"001110110",
  7348=>"110110111",
  7349=>"001000111",
  7350=>"011001111",
  7351=>"011000100",
  7352=>"111000110",
  7353=>"101101001",
  7354=>"010010100",
  7355=>"011111011",
  7356=>"001010010",
  7357=>"110101101",
  7358=>"110110000",
  7359=>"110111001",
  7360=>"010000011",
  7361=>"010011101",
  7362=>"001000000",
  7363=>"001010111",
  7364=>"001101111",
  7365=>"111001001",
  7366=>"110011101",
  7367=>"111011000",
  7368=>"110001011",
  7369=>"011101110",
  7370=>"110111010",
  7371=>"011111011",
  7372=>"010101010",
  7373=>"101001111",
  7374=>"000000111",
  7375=>"001101000",
  7376=>"011000010",
  7377=>"100101000",
  7378=>"011000010",
  7379=>"001000011",
  7380=>"010111001",
  7381=>"110110100",
  7382=>"110010011",
  7383=>"000100000",
  7384=>"100111001",
  7385=>"100110001",
  7386=>"101001100",
  7387=>"110100000",
  7388=>"011001111",
  7389=>"101111110",
  7390=>"000101000",
  7391=>"011100000",
  7392=>"100000111",
  7393=>"111001110",
  7394=>"100101100",
  7395=>"100100001",
  7396=>"001000100",
  7397=>"101111110",
  7398=>"100111011",
  7399=>"000011110",
  7400=>"011101011",
  7401=>"111111011",
  7402=>"101111010",
  7403=>"101000101",
  7404=>"101101010",
  7405=>"100110111",
  7406=>"010010001",
  7407=>"111110000",
  7408=>"100010010",
  7409=>"001001010",
  7410=>"011100101",
  7411=>"101100111",
  7412=>"011011011",
  7413=>"100001000",
  7414=>"100111010",
  7415=>"111011000",
  7416=>"001000111",
  7417=>"110100010",
  7418=>"001111010",
  7419=>"001101010",
  7420=>"000001010",
  7421=>"000000011",
  7422=>"101001101",
  7423=>"100111011",
  7424=>"001001010",
  7425=>"011010111",
  7426=>"101101100",
  7427=>"100000011",
  7428=>"110000011",
  7429=>"010111110",
  7430=>"010010101",
  7431=>"100000101",
  7432=>"100101000",
  7433=>"100100011",
  7434=>"001101000",
  7435=>"010011100",
  7436=>"001001001",
  7437=>"000011001",
  7438=>"010010001",
  7439=>"000010111",
  7440=>"001110101",
  7441=>"000100011",
  7442=>"000001000",
  7443=>"100101101",
  7444=>"000110001",
  7445=>"011011011",
  7446=>"000100101",
  7447=>"011010111",
  7448=>"100101011",
  7449=>"101100010",
  7450=>"110100010",
  7451=>"000000111",
  7452=>"000010111",
  7453=>"100010100",
  7454=>"001110110",
  7455=>"000010110",
  7456=>"110000101",
  7457=>"110010000",
  7458=>"011110010",
  7459=>"101100111",
  7460=>"001011011",
  7461=>"100110101",
  7462=>"000011111",
  7463=>"010110101",
  7464=>"000001000",
  7465=>"011110010",
  7466=>"011111111",
  7467=>"101010111",
  7468=>"010100010",
  7469=>"001000001",
  7470=>"110000000",
  7471=>"101011101",
  7472=>"000001111",
  7473=>"000010000",
  7474=>"111111111",
  7475=>"100001100",
  7476=>"101001101",
  7477=>"100000011",
  7478=>"100001110",
  7479=>"000001001",
  7480=>"010001101",
  7481=>"101100111",
  7482=>"000111001",
  7483=>"000110000",
  7484=>"111001000",
  7485=>"011111110",
  7486=>"101000001",
  7487=>"101011100",
  7488=>"100101000",
  7489=>"001010000",
  7490=>"011111111",
  7491=>"001101100",
  7492=>"111011111",
  7493=>"101010011",
  7494=>"100011001",
  7495=>"101011110",
  7496=>"001000011",
  7497=>"011101011",
  7498=>"100110010",
  7499=>"111001010",
  7500=>"111101011",
  7501=>"100101011",
  7502=>"100000001",
  7503=>"001000010",
  7504=>"110110010",
  7505=>"110011001",
  7506=>"100101001",
  7507=>"000100011",
  7508=>"110010001",
  7509=>"101010000",
  7510=>"011010111",
  7511=>"100110011",
  7512=>"001001000",
  7513=>"001100100",
  7514=>"100010110",
  7515=>"111100000",
  7516=>"000110101",
  7517=>"010110100",
  7518=>"001001011",
  7519=>"000100110",
  7520=>"011110000",
  7521=>"011110101",
  7522=>"000010010",
  7523=>"110111110",
  7524=>"011000111",
  7525=>"010010110",
  7526=>"011101110",
  7527=>"111111001",
  7528=>"001000000",
  7529=>"111001110",
  7530=>"010001011",
  7531=>"101000010",
  7532=>"011100110",
  7533=>"100111101",
  7534=>"001001010",
  7535=>"011000011",
  7536=>"110101111",
  7537=>"111000000",
  7538=>"000011110",
  7539=>"000011001",
  7540=>"001110101",
  7541=>"111110101",
  7542=>"010101000",
  7543=>"010011111",
  7544=>"001101110",
  7545=>"100010010",
  7546=>"111010110",
  7547=>"111011011",
  7548=>"101111000",
  7549=>"001101011",
  7550=>"101010100",
  7551=>"101111011",
  7552=>"110111101",
  7553=>"101011101",
  7554=>"011000001",
  7555=>"100101101",
  7556=>"000011110",
  7557=>"000010011",
  7558=>"010010101",
  7559=>"001001000",
  7560=>"010001110",
  7561=>"000000011",
  7562=>"100010001",
  7563=>"111011000",
  7564=>"010100101",
  7565=>"101101100",
  7566=>"011000011",
  7567=>"001111110",
  7568=>"110001110",
  7569=>"011011100",
  7570=>"011100111",
  7571=>"101100001",
  7572=>"000001010",
  7573=>"000110010",
  7574=>"110101111",
  7575=>"100000111",
  7576=>"010011100",
  7577=>"011000100",
  7578=>"000001001",
  7579=>"001011110",
  7580=>"000000001",
  7581=>"111000110",
  7582=>"011001001",
  7583=>"110011000",
  7584=>"100010001",
  7585=>"110101000",
  7586=>"000100000",
  7587=>"111011000",
  7588=>"101111111",
  7589=>"110010010",
  7590=>"010011111",
  7591=>"001000111",
  7592=>"010001011",
  7593=>"111110101",
  7594=>"010001100",
  7595=>"111111111",
  7596=>"101110000",
  7597=>"111110011",
  7598=>"000001110",
  7599=>"010010100",
  7600=>"011011100",
  7601=>"001000100",
  7602=>"010000101",
  7603=>"010001000",
  7604=>"000011010",
  7605=>"010010100",
  7606=>"100100110",
  7607=>"001000110",
  7608=>"011011100",
  7609=>"100001111",
  7610=>"011001001",
  7611=>"101100111",
  7612=>"010010110",
  7613=>"111010110",
  7614=>"001010101",
  7615=>"110010110",
  7616=>"011110001",
  7617=>"011011100",
  7618=>"010101110",
  7619=>"110111101",
  7620=>"101110000",
  7621=>"011000101",
  7622=>"001010101",
  7623=>"000011011",
  7624=>"001001100",
  7625=>"010000111",
  7626=>"010000110",
  7627=>"001100100",
  7628=>"001000111",
  7629=>"100001101",
  7630=>"010011001",
  7631=>"000010000",
  7632=>"111011000",
  7633=>"001100010",
  7634=>"111101011",
  7635=>"111101000",
  7636=>"011011110",
  7637=>"011111001",
  7638=>"011100011",
  7639=>"111010100",
  7640=>"001001000",
  7641=>"101110110",
  7642=>"000110000",
  7643=>"111110101",
  7644=>"011100001",
  7645=>"101001000",
  7646=>"110100110",
  7647=>"101110101",
  7648=>"110111001",
  7649=>"100010100",
  7650=>"111110101",
  7651=>"110000100",
  7652=>"000110000",
  7653=>"011010001",
  7654=>"000011010",
  7655=>"010101101",
  7656=>"011011101",
  7657=>"100011011",
  7658=>"000111101",
  7659=>"101000111",
  7660=>"011000111",
  7661=>"011111001",
  7662=>"100110001",
  7663=>"011001110",
  7664=>"110111000",
  7665=>"011010101",
  7666=>"101011011",
  7667=>"110110100",
  7668=>"011000111",
  7669=>"000011010",
  7670=>"000011110",
  7671=>"100100111",
  7672=>"001011011",
  7673=>"111011000",
  7674=>"100001100",
  7675=>"111010011",
  7676=>"000010101",
  7677=>"000000000",
  7678=>"010000011",
  7679=>"011001111",
  7680=>"101101110",
  7681=>"010000101",
  7682=>"111110111",
  7683=>"001001100",
  7684=>"101101011",
  7685=>"010111000",
  7686=>"010101100",
  7687=>"100110011",
  7688=>"010001010",
  7689=>"001101101",
  7690=>"010000011",
  7691=>"101001111",
  7692=>"001101001",
  7693=>"110001000",
  7694=>"001011100",
  7695=>"011001110",
  7696=>"000010001",
  7697=>"010000100",
  7698=>"111001001",
  7699=>"111100101",
  7700=>"110010101",
  7701=>"000011011",
  7702=>"010111110",
  7703=>"100100010",
  7704=>"000100100",
  7705=>"110011101",
  7706=>"101100110",
  7707=>"011001010",
  7708=>"111101111",
  7709=>"000010011",
  7710=>"000000110",
  7711=>"110000000",
  7712=>"010011001",
  7713=>"100111010",
  7714=>"010101010",
  7715=>"001011110",
  7716=>"101101111",
  7717=>"111000000",
  7718=>"001110101",
  7719=>"000111001",
  7720=>"001001101",
  7721=>"010010010",
  7722=>"101111011",
  7723=>"001000100",
  7724=>"001000010",
  7725=>"101110101",
  7726=>"000101110",
  7727=>"011010011",
  7728=>"010010001",
  7729=>"001010111",
  7730=>"001010111",
  7731=>"011001100",
  7732=>"111101100",
  7733=>"011010111",
  7734=>"111011001",
  7735=>"111110010",
  7736=>"011110111",
  7737=>"101100010",
  7738=>"010110011",
  7739=>"110001011",
  7740=>"111000100",
  7741=>"001000100",
  7742=>"010110101",
  7743=>"100110000",
  7744=>"111111010",
  7745=>"111100010",
  7746=>"110010011",
  7747=>"010101100",
  7748=>"010100000",
  7749=>"000101101",
  7750=>"111111001",
  7751=>"100011100",
  7752=>"101101110",
  7753=>"111110000",
  7754=>"000100111",
  7755=>"100011111",
  7756=>"111110001",
  7757=>"000100101",
  7758=>"000101000",
  7759=>"100111011",
  7760=>"011000100",
  7761=>"111101101",
  7762=>"000010100",
  7763=>"111001111",
  7764=>"000010111",
  7765=>"000001111",
  7766=>"001110101",
  7767=>"000101010",
  7768=>"000011000",
  7769=>"111100111",
  7770=>"001100001",
  7771=>"101010000",
  7772=>"000000010",
  7773=>"000000000",
  7774=>"000101101",
  7775=>"110011001",
  7776=>"111010001",
  7777=>"111010111",
  7778=>"101100100",
  7779=>"010001011",
  7780=>"010101101",
  7781=>"000111101",
  7782=>"000011100",
  7783=>"000000010",
  7784=>"011110011",
  7785=>"100011000",
  7786=>"010001001",
  7787=>"111100110",
  7788=>"110011100",
  7789=>"110011110",
  7790=>"001100110",
  7791=>"000010001",
  7792=>"100010010",
  7793=>"111010011",
  7794=>"100101010",
  7795=>"101101101",
  7796=>"011000011",
  7797=>"111100101",
  7798=>"111101011",
  7799=>"110011001",
  7800=>"111110001",
  7801=>"101110001",
  7802=>"111100010",
  7803=>"100101110",
  7804=>"100011001",
  7805=>"110101000",
  7806=>"001000100",
  7807=>"010110000",
  7808=>"000101000",
  7809=>"101111101",
  7810=>"010101101",
  7811=>"001000100",
  7812=>"111101001",
  7813=>"101101111",
  7814=>"111110010",
  7815=>"011100011",
  7816=>"110010011",
  7817=>"111100010",
  7818=>"100101101",
  7819=>"001111100",
  7820=>"000111000",
  7821=>"110010011",
  7822=>"111111001",
  7823=>"101001001",
  7824=>"110010011",
  7825=>"111100101",
  7826=>"100110010",
  7827=>"011110111",
  7828=>"110100001",
  7829=>"000011100",
  7830=>"110010101",
  7831=>"001010001",
  7832=>"101010100",
  7833=>"110011110",
  7834=>"111101000",
  7835=>"010000011",
  7836=>"010000111",
  7837=>"101001101",
  7838=>"101010101",
  7839=>"110011100",
  7840=>"101110001",
  7841=>"111001011",
  7842=>"110010000",
  7843=>"111111101",
  7844=>"001101011",
  7845=>"111001011",
  7846=>"100010011",
  7847=>"001100101",
  7848=>"111011100",
  7849=>"111000110",
  7850=>"111010010",
  7851=>"101010001",
  7852=>"010001011",
  7853=>"000110010",
  7854=>"111010100",
  7855=>"100101100",
  7856=>"001010100",
  7857=>"001001100",
  7858=>"010011110",
  7859=>"011001011",
  7860=>"110111001",
  7861=>"011101001",
  7862=>"100111011",
  7863=>"001010001",
  7864=>"101001011",
  7865=>"011110111",
  7866=>"101111011",
  7867=>"010010000",
  7868=>"110100110",
  7869=>"011101000",
  7870=>"100011001",
  7871=>"100111011",
  7872=>"111110001",
  7873=>"110001011",
  7874=>"001101111",
  7875=>"111101010",
  7876=>"111111111",
  7877=>"101001100",
  7878=>"000100110",
  7879=>"001001110",
  7880=>"010000001",
  7881=>"011001001",
  7882=>"111101111",
  7883=>"011000110",
  7884=>"011110000",
  7885=>"000010010",
  7886=>"000000111",
  7887=>"011010010",
  7888=>"001110100",
  7889=>"001101100",
  7890=>"000101110",
  7891=>"011001011",
  7892=>"001100000",
  7893=>"000001111",
  7894=>"011100111",
  7895=>"001110101",
  7896=>"001000110",
  7897=>"001000111",
  7898=>"010110010",
  7899=>"111100110",
  7900=>"111101100",
  7901=>"010000000",
  7902=>"001001100",
  7903=>"001000000",
  7904=>"100110110",
  7905=>"000000000",
  7906=>"101100111",
  7907=>"000010011",
  7908=>"111111011",
  7909=>"011101000",
  7910=>"110110000",
  7911=>"011000111",
  7912=>"000101100",
  7913=>"111101100",
  7914=>"101110010",
  7915=>"110010011",
  7916=>"001100011",
  7917=>"011001111",
  7918=>"110000101",
  7919=>"111101110",
  7920=>"101111110",
  7921=>"001001010",
  7922=>"101110010",
  7923=>"010010000",
  7924=>"001010001",
  7925=>"100001010",
  7926=>"111001111",
  7927=>"011001001",
  7928=>"101100000",
  7929=>"110010010",
  7930=>"111111001",
  7931=>"011100111",
  7932=>"000011101",
  7933=>"100100110",
  7934=>"010111011",
  7935=>"001011000",
  7936=>"011101101",
  7937=>"111111001",
  7938=>"110110001",
  7939=>"101101001",
  7940=>"011001000",
  7941=>"101001110",
  7942=>"111110100",
  7943=>"110110100",
  7944=>"001110000",
  7945=>"000111000",
  7946=>"011110000",
  7947=>"001010001",
  7948=>"100010000",
  7949=>"001110100",
  7950=>"001000011",
  7951=>"000001001",
  7952=>"100000011",
  7953=>"001000011",
  7954=>"001001110",
  7955=>"010000011",
  7956=>"011100100",
  7957=>"000110011",
  7958=>"000001000",
  7959=>"110010111",
  7960=>"001001101",
  7961=>"010010001",
  7962=>"000000110",
  7963=>"001010000",
  7964=>"111100001",
  7965=>"010011001",
  7966=>"111011011",
  7967=>"000011110",
  7968=>"111100101",
  7969=>"110010001",
  7970=>"100011101",
  7971=>"000010010",
  7972=>"011001010",
  7973=>"100011100",
  7974=>"011001010",
  7975=>"010100100",
  7976=>"011101000",
  7977=>"001110110",
  7978=>"110000100",
  7979=>"110010100",
  7980=>"010111000",
  7981=>"001111010",
  7982=>"000001101",
  7983=>"101001000",
  7984=>"010000000",
  7985=>"101110001",
  7986=>"100000001",
  7987=>"000010111",
  7988=>"011011000",
  7989=>"110111100",
  7990=>"011111000",
  7991=>"111001011",
  7992=>"000101010",
  7993=>"110111000",
  7994=>"011011111",
  7995=>"111011101",
  7996=>"001000100",
  7997=>"101001110",
  7998=>"010010110",
  7999=>"101100000",
  8000=>"110011011",
  8001=>"100001011",
  8002=>"010000100",
  8003=>"110001000",
  8004=>"000101010",
  8005=>"011100111",
  8006=>"111000111",
  8007=>"000101001",
  8008=>"010110101",
  8009=>"000001110",
  8010=>"001011010",
  8011=>"111100000",
  8012=>"011011011",
  8013=>"011100100",
  8014=>"000110111",
  8015=>"011010100",
  8016=>"010001110",
  8017=>"000110110",
  8018=>"000101010",
  8019=>"111010010",
  8020=>"110101111",
  8021=>"000101100",
  8022=>"010111000",
  8023=>"110111111",
  8024=>"001000011",
  8025=>"010110111",
  8026=>"001100110",
  8027=>"110100001",
  8028=>"011010000",
  8029=>"100010011",
  8030=>"001000111",
  8031=>"000100100",
  8032=>"011000001",
  8033=>"110111101",
  8034=>"010000000",
  8035=>"011110101",
  8036=>"010001101",
  8037=>"101101111",
  8038=>"111100010",
  8039=>"100010111",
  8040=>"001100010",
  8041=>"001101001",
  8042=>"011000011",
  8043=>"011011100",
  8044=>"011000000",
  8045=>"110001011",
  8046=>"010000101",
  8047=>"100100110",
  8048=>"110110000",
  8049=>"111100011",
  8050=>"111101100",
  8051=>"010010011",
  8052=>"110010010",
  8053=>"101000101",
  8054=>"101001011",
  8055=>"010010000",
  8056=>"001001001",
  8057=>"010000010",
  8058=>"000101001",
  8059=>"011010000",
  8060=>"000000001",
  8061=>"111011110",
  8062=>"110111101",
  8063=>"110001101",
  8064=>"100011011",
  8065=>"100111011",
  8066=>"000001001",
  8067=>"111100011",
  8068=>"001000010",
  8069=>"001000000",
  8070=>"111011101",
  8071=>"011001101",
  8072=>"001011111",
  8073=>"011100000",
  8074=>"001000101",
  8075=>"000001101",
  8076=>"100000110",
  8077=>"010000101",
  8078=>"001011110",
  8079=>"110110111",
  8080=>"001011100",
  8081=>"010111101",
  8082=>"101100011",
  8083=>"111111011",
  8084=>"111110010",
  8085=>"111011100",
  8086=>"011010101",
  8087=>"001000110",
  8088=>"101001100",
  8089=>"100111111",
  8090=>"001100100",
  8091=>"110010011",
  8092=>"110010011",
  8093=>"011110110",
  8094=>"000100101",
  8095=>"101111000",
  8096=>"100101110",
  8097=>"011011100",
  8098=>"001101111",
  8099=>"111101000",
  8100=>"111111000",
  8101=>"001101100",
  8102=>"100001010",
  8103=>"010000010",
  8104=>"100011000",
  8105=>"000010101",
  8106=>"100111010",
  8107=>"001010101",
  8108=>"101110010",
  8109=>"111000101",
  8110=>"101100100",
  8111=>"101100111",
  8112=>"110000110",
  8113=>"111101000",
  8114=>"110011101",
  8115=>"000100000",
  8116=>"010110011",
  8117=>"001111100",
  8118=>"001100011",
  8119=>"111111110",
  8120=>"100000100",
  8121=>"000100100",
  8122=>"110101101",
  8123=>"000101000",
  8124=>"000010111",
  8125=>"000101110",
  8126=>"101100001",
  8127=>"000011000",
  8128=>"101111100",
  8129=>"000011110",
  8130=>"001001101",
  8131=>"010000011",
  8132=>"000000111",
  8133=>"111101001",
  8134=>"000111100",
  8135=>"000001010",
  8136=>"001010000",
  8137=>"111110100",
  8138=>"110000001",
  8139=>"110010000",
  8140=>"101100010",
  8141=>"010001111",
  8142=>"001110000",
  8143=>"111100100",
  8144=>"100000011",
  8145=>"011110111",
  8146=>"000101000",
  8147=>"110101010",
  8148=>"001100001",
  8149=>"010001000",
  8150=>"110001100",
  8151=>"000000001",
  8152=>"100110100",
  8153=>"110000000",
  8154=>"110001001",
  8155=>"101100110",
  8156=>"110000001",
  8157=>"001111010",
  8158=>"101111011",
  8159=>"101100011",
  8160=>"011111100",
  8161=>"101001111",
  8162=>"010000000",
  8163=>"001111100",
  8164=>"000011001",
  8165=>"110111001",
  8166=>"000100111",
  8167=>"000110000",
  8168=>"101100000",
  8169=>"100011110",
  8170=>"100011111",
  8171=>"011000101",
  8172=>"011100110",
  8173=>"110111101",
  8174=>"010100111",
  8175=>"011010001",
  8176=>"101010001",
  8177=>"110111010",
  8178=>"010000101",
  8179=>"000110011",
  8180=>"101101101",
  8181=>"110110000",
  8182=>"110110010",
  8183=>"111101110",
  8184=>"101010101",
  8185=>"110101001",
  8186=>"001110001",
  8187=>"000000110",
  8188=>"111101110",
  8189=>"010010110",
  8190=>"010111100",
  8191=>"111110101",
  8192=>"000010100",
  8193=>"011000100",
  8194=>"110010011",
  8195=>"000000000",
  8196=>"000000000",
  8197=>"100110110",
  8198=>"101110111",
  8199=>"000010100",
  8200=>"100010110",
  8201=>"001011100",
  8202=>"000001011",
  8203=>"110100010",
  8204=>"101100111",
  8205=>"000110001",
  8206=>"111010001",
  8207=>"000111110",
  8208=>"111100101",
  8209=>"000011000",
  8210=>"000001011",
  8211=>"010000100",
  8212=>"010001011",
  8213=>"011101101",
  8214=>"111111111",
  8215=>"000100010",
  8216=>"100101110",
  8217=>"100001100",
  8218=>"100110011",
  8219=>"011111100",
  8220=>"101110000",
  8221=>"101011101",
  8222=>"100110100",
  8223=>"101111111",
  8224=>"010000011",
  8225=>"110111011",
  8226=>"001100111",
  8227=>"101100011",
  8228=>"011011010",
  8229=>"011100000",
  8230=>"100010010",
  8231=>"010000001",
  8232=>"110000010",
  8233=>"001111101",
  8234=>"100010110",
  8235=>"101101001",
  8236=>"010110010",
  8237=>"100000111",
  8238=>"101000010",
  8239=>"111000110",
  8240=>"001010000",
  8241=>"110111101",
  8242=>"100110101",
  8243=>"110100100",
  8244=>"000010110",
  8245=>"000000010",
  8246=>"100000100",
  8247=>"010111011",
  8248=>"010111011",
  8249=>"101100100",
  8250=>"011000100",
  8251=>"010110100",
  8252=>"000001101",
  8253=>"001001001",
  8254=>"110000011",
  8255=>"000101001",
  8256=>"101101011",
  8257=>"001011101",
  8258=>"101110110",
  8259=>"101001110",
  8260=>"000100100",
  8261=>"100110100",
  8262=>"100100100",
  8263=>"001000101",
  8264=>"000010000",
  8265=>"101010010",
  8266=>"000111101",
  8267=>"010010100",
  8268=>"000001011",
  8269=>"010111100",
  8270=>"101000010",
  8271=>"110111000",
  8272=>"111011100",
  8273=>"000011000",
  8274=>"010111111",
  8275=>"001010001",
  8276=>"100110010",
  8277=>"010010100",
  8278=>"111001011",
  8279=>"010010001",
  8280=>"001010100",
  8281=>"000010011",
  8282=>"000000001",
  8283=>"001010000",
  8284=>"100100010",
  8285=>"100010011",
  8286=>"101010100",
  8287=>"000010011",
  8288=>"110101011",
  8289=>"001111111",
  8290=>"110011100",
  8291=>"001101000",
  8292=>"010110000",
  8293=>"110011011",
  8294=>"111011111",
  8295=>"000100011",
  8296=>"000111101",
  8297=>"111000000",
  8298=>"100010010",
  8299=>"010100110",
  8300=>"110001111",
  8301=>"010011000",
  8302=>"100100010",
  8303=>"011111111",
  8304=>"001000000",
  8305=>"010101001",
  8306=>"101011110",
  8307=>"111111000",
  8308=>"011010111",
  8309=>"011000101",
  8310=>"011000010",
  8311=>"101010111",
  8312=>"011111010",
  8313=>"111000101",
  8314=>"010001110",
  8315=>"100101001",
  8316=>"011000100",
  8317=>"011111001",
  8318=>"011010001",
  8319=>"011111101",
  8320=>"110001110",
  8321=>"010000101",
  8322=>"011101100",
  8323=>"000100010",
  8324=>"100100000",
  8325=>"001100101",
  8326=>"011101000",
  8327=>"100111111",
  8328=>"100100101",
  8329=>"111100011",
  8330=>"001011001",
  8331=>"010101101",
  8332=>"010111001",
  8333=>"101001111",
  8334=>"100101100",
  8335=>"001000001",
  8336=>"101101110",
  8337=>"011000000",
  8338=>"001011110",
  8339=>"110000101",
  8340=>"100111110",
  8341=>"101000011",
  8342=>"000000101",
  8343=>"011111011",
  8344=>"000001000",
  8345=>"101000000",
  8346=>"111011011",
  8347=>"011110001",
  8348=>"011001000",
  8349=>"010110110",
  8350=>"001001101",
  8351=>"000101111",
  8352=>"011101010",
  8353=>"110000011",
  8354=>"111111000",
  8355=>"001111111",
  8356=>"001110110",
  8357=>"000110000",
  8358=>"010011010",
  8359=>"100010100",
  8360=>"110000011",
  8361=>"100010111",
  8362=>"101011100",
  8363=>"110110100",
  8364=>"110100101",
  8365=>"001111001",
  8366=>"010001101",
  8367=>"001101111",
  8368=>"010011111",
  8369=>"101111100",
  8370=>"000001001",
  8371=>"011101001",
  8372=>"011000000",
  8373=>"101111000",
  8374=>"010110110",
  8375=>"100000011",
  8376=>"110100000",
  8377=>"010111111",
  8378=>"000010100",
  8379=>"101110101",
  8380=>"001010001",
  8381=>"100000110",
  8382=>"000000111",
  8383=>"011100001",
  8384=>"110110111",
  8385=>"001010010",
  8386=>"000010100",
  8387=>"001010000",
  8388=>"011000001",
  8389=>"000110110",
  8390=>"011111000",
  8391=>"101101111",
  8392=>"111000011",
  8393=>"111111011",
  8394=>"111000111",
  8395=>"111011001",
  8396=>"011010001",
  8397=>"110011111",
  8398=>"011100000",
  8399=>"110011100",
  8400=>"101011100",
  8401=>"000001100",
  8402=>"100110000",
  8403=>"110001010",
  8404=>"000111011",
  8405=>"010000000",
  8406=>"110100100",
  8407=>"110101100",
  8408=>"000101010",
  8409=>"011100000",
  8410=>"001110111",
  8411=>"011101110",
  8412=>"110101010",
  8413=>"010100011",
  8414=>"000110111",
  8415=>"000110101",
  8416=>"111001111",
  8417=>"100100000",
  8418=>"111001101",
  8419=>"011010011",
  8420=>"111110101",
  8421=>"111101011",
  8422=>"111011101",
  8423=>"000000101",
  8424=>"100011010",
  8425=>"111101100",
  8426=>"001111011",
  8427=>"000101100",
  8428=>"111110001",
  8429=>"001000101",
  8430=>"100000100",
  8431=>"011100001",
  8432=>"111110101",
  8433=>"100010001",
  8434=>"000100101",
  8435=>"111110101",
  8436=>"011010011",
  8437=>"011111100",
  8438=>"111010100",
  8439=>"101000001",
  8440=>"000000010",
  8441=>"001100101",
  8442=>"010000100",
  8443=>"101100110",
  8444=>"001000010",
  8445=>"011000010",
  8446=>"100000111",
  8447=>"010110010",
  8448=>"010101000",
  8449=>"011111110",
  8450=>"010100011",
  8451=>"111100110",
  8452=>"101111101",
  8453=>"101101100",
  8454=>"100111001",
  8455=>"101001001",
  8456=>"011111101",
  8457=>"011111111",
  8458=>"001010101",
  8459=>"101000001",
  8460=>"010011101",
  8461=>"101001011",
  8462=>"010010101",
  8463=>"000010111",
  8464=>"110000001",
  8465=>"001010010",
  8466=>"110101111",
  8467=>"010111000",
  8468=>"110111011",
  8469=>"100110100",
  8470=>"110100000",
  8471=>"011000100",
  8472=>"110000101",
  8473=>"100101100",
  8474=>"011100111",
  8475=>"111100100",
  8476=>"000010001",
  8477=>"010110010",
  8478=>"000011111",
  8479=>"110010111",
  8480=>"100101011",
  8481=>"111101101",
  8482=>"010011000",
  8483=>"100100101",
  8484=>"100010110",
  8485=>"111001111",
  8486=>"111000011",
  8487=>"011000010",
  8488=>"000110100",
  8489=>"010110011",
  8490=>"001000111",
  8491=>"001111111",
  8492=>"101001100",
  8493=>"110001100",
  8494=>"010000101",
  8495=>"000101101",
  8496=>"100001001",
  8497=>"001001000",
  8498=>"110100100",
  8499=>"010011000",
  8500=>"010100101",
  8501=>"100110001",
  8502=>"111111010",
  8503=>"001110100",
  8504=>"000010111",
  8505=>"110001101",
  8506=>"011100100",
  8507=>"101101000",
  8508=>"010010011",
  8509=>"000110100",
  8510=>"101011100",
  8511=>"111111010",
  8512=>"011000011",
  8513=>"110100101",
  8514=>"000001001",
  8515=>"110110101",
  8516=>"111100111",
  8517=>"001111000",
  8518=>"001110000",
  8519=>"100111010",
  8520=>"001101100",
  8521=>"100010100",
  8522=>"011101101",
  8523=>"100111100",
  8524=>"000111110",
  8525=>"011010000",
  8526=>"100001100",
  8527=>"101111001",
  8528=>"010101001",
  8529=>"000001111",
  8530=>"010010000",
  8531=>"010111100",
  8532=>"101101111",
  8533=>"001101110",
  8534=>"011110010",
  8535=>"010110101",
  8536=>"000000110",
  8537=>"000101010",
  8538=>"110101100",
  8539=>"001010110",
  8540=>"010001111",
  8541=>"100010011",
  8542=>"111011100",
  8543=>"010011000",
  8544=>"000111111",
  8545=>"111011100",
  8546=>"000010100",
  8547=>"000000000",
  8548=>"111101101",
  8549=>"001100000",
  8550=>"010011111",
  8551=>"110100100",
  8552=>"001101000",
  8553=>"100010001",
  8554=>"000100011",
  8555=>"000100001",
  8556=>"011010010",
  8557=>"110011100",
  8558=>"000010001",
  8559=>"100110111",
  8560=>"000011110",
  8561=>"111110001",
  8562=>"110111100",
  8563=>"111100101",
  8564=>"000010110",
  8565=>"000111110",
  8566=>"001001001",
  8567=>"001000110",
  8568=>"101110001",
  8569=>"100011100",
  8570=>"110110111",
  8571=>"110111110",
  8572=>"111111010",
  8573=>"010011111",
  8574=>"101000101",
  8575=>"100110011",
  8576=>"110010101",
  8577=>"111110101",
  8578=>"111100110",
  8579=>"111111011",
  8580=>"011001110",
  8581=>"010100110",
  8582=>"110110100",
  8583=>"011110110",
  8584=>"011111111",
  8585=>"101111111",
  8586=>"000001100",
  8587=>"010001011",
  8588=>"101100010",
  8589=>"101100111",
  8590=>"100100010",
  8591=>"111000010",
  8592=>"111110101",
  8593=>"110100101",
  8594=>"000100011",
  8595=>"100111101",
  8596=>"010110000",
  8597=>"111101000",
  8598=>"001101101",
  8599=>"111111111",
  8600=>"101010111",
  8601=>"100110101",
  8602=>"001100110",
  8603=>"000000100",
  8604=>"011110100",
  8605=>"111001100",
  8606=>"011010110",
  8607=>"110010111",
  8608=>"000011100",
  8609=>"100100111",
  8610=>"000100001",
  8611=>"000000000",
  8612=>"001001011",
  8613=>"010011000",
  8614=>"110000011",
  8615=>"010000100",
  8616=>"010000100",
  8617=>"111110001",
  8618=>"100011111",
  8619=>"111010101",
  8620=>"101111000",
  8621=>"100001101",
  8622=>"010101001",
  8623=>"111001001",
  8624=>"100111100",
  8625=>"001100001",
  8626=>"011101110",
  8627=>"100111110",
  8628=>"101110001",
  8629=>"011110110",
  8630=>"000100010",
  8631=>"110010011",
  8632=>"000111001",
  8633=>"100011000",
  8634=>"001011001",
  8635=>"100001100",
  8636=>"010101010",
  8637=>"100001111",
  8638=>"111100011",
  8639=>"110110011",
  8640=>"001001100",
  8641=>"000010011",
  8642=>"111101101",
  8643=>"010110001",
  8644=>"011001111",
  8645=>"000011001",
  8646=>"000101011",
  8647=>"011001110",
  8648=>"001011010",
  8649=>"011001001",
  8650=>"000110110",
  8651=>"001010010",
  8652=>"101011110",
  8653=>"000000001",
  8654=>"100111110",
  8655=>"000011000",
  8656=>"110000001",
  8657=>"000000000",
  8658=>"010100110",
  8659=>"110111011",
  8660=>"010101000",
  8661=>"010110100",
  8662=>"011001110",
  8663=>"110101110",
  8664=>"000100110",
  8665=>"111000100",
  8666=>"010110110",
  8667=>"110100000",
  8668=>"010100100",
  8669=>"101010000",
  8670=>"001110110",
  8671=>"110011000",
  8672=>"000001111",
  8673=>"000010100",
  8674=>"001001000",
  8675=>"111000111",
  8676=>"110010101",
  8677=>"111110101",
  8678=>"000000100",
  8679=>"000111000",
  8680=>"011001001",
  8681=>"111000111",
  8682=>"100010100",
  8683=>"101111000",
  8684=>"000110110",
  8685=>"101000110",
  8686=>"000101000",
  8687=>"101100010",
  8688=>"000101110",
  8689=>"001001111",
  8690=>"000110010",
  8691=>"101111000",
  8692=>"001000100",
  8693=>"110100100",
  8694=>"111100001",
  8695=>"000010011",
  8696=>"010101110",
  8697=>"110001011",
  8698=>"001100101",
  8699=>"000101110",
  8700=>"100101100",
  8701=>"100100100",
  8702=>"100111100",
  8703=>"101100110",
  8704=>"111111100",
  8705=>"110000001",
  8706=>"100111011",
  8707=>"101100010",
  8708=>"010111011",
  8709=>"110100110",
  8710=>"111100000",
  8711=>"000011000",
  8712=>"011101111",
  8713=>"110110111",
  8714=>"101010011",
  8715=>"010011101",
  8716=>"100011101",
  8717=>"011100011",
  8718=>"100001011",
  8719=>"011001110",
  8720=>"101111000",
  8721=>"101010010",
  8722=>"010111100",
  8723=>"111110101",
  8724=>"011000101",
  8725=>"101000000",
  8726=>"011010110",
  8727=>"000101000",
  8728=>"000001111",
  8729=>"000101111",
  8730=>"010010100",
  8731=>"101110110",
  8732=>"110010111",
  8733=>"000110111",
  8734=>"110000110",
  8735=>"110001001",
  8736=>"110010101",
  8737=>"111110111",
  8738=>"000000010",
  8739=>"000111101",
  8740=>"011011101",
  8741=>"010011100",
  8742=>"001001101",
  8743=>"010010000",
  8744=>"110100100",
  8745=>"000001110",
  8746=>"110110000",
  8747=>"100000111",
  8748=>"101101110",
  8749=>"100100011",
  8750=>"001101100",
  8751=>"001101110",
  8752=>"111111001",
  8753=>"101011111",
  8754=>"110111111",
  8755=>"000100000",
  8756=>"001010000",
  8757=>"001010010",
  8758=>"100000111",
  8759=>"110000110",
  8760=>"001001001",
  8761=>"000000001",
  8762=>"110010110",
  8763=>"110101111",
  8764=>"001100010",
  8765=>"001101000",
  8766=>"000110010",
  8767=>"101010000",
  8768=>"111011111",
  8769=>"110111110",
  8770=>"110000011",
  8771=>"010011011",
  8772=>"110101011",
  8773=>"110001010",
  8774=>"001001010",
  8775=>"010111010",
  8776=>"110111110",
  8777=>"111100111",
  8778=>"001011011",
  8779=>"010100011",
  8780=>"000010010",
  8781=>"101100000",
  8782=>"011100111",
  8783=>"001000011",
  8784=>"111000111",
  8785=>"001101101",
  8786=>"011101000",
  8787=>"100110010",
  8788=>"110000111",
  8789=>"001100001",
  8790=>"000100100",
  8791=>"000110111",
  8792=>"011100001",
  8793=>"111000111",
  8794=>"010110100",
  8795=>"000100110",
  8796=>"100100000",
  8797=>"001101111",
  8798=>"000011001",
  8799=>"101110110",
  8800=>"101010001",
  8801=>"100101111",
  8802=>"011001111",
  8803=>"111111001",
  8804=>"100001111",
  8805=>"100001010",
  8806=>"010000101",
  8807=>"101000110",
  8808=>"001100101",
  8809=>"111010011",
  8810=>"011000010",
  8811=>"001110000",
  8812=>"100111011",
  8813=>"010101011",
  8814=>"101000111",
  8815=>"000010001",
  8816=>"000000101",
  8817=>"010010011",
  8818=>"011111001",
  8819=>"101001000",
  8820=>"111000011",
  8821=>"110010010",
  8822=>"011100011",
  8823=>"011101001",
  8824=>"010010111",
  8825=>"101110100",
  8826=>"100000100",
  8827=>"001001011",
  8828=>"000000001",
  8829=>"011100001",
  8830=>"011101100",
  8831=>"111100110",
  8832=>"111110110",
  8833=>"011101101",
  8834=>"000111111",
  8835=>"101110100",
  8836=>"011011010",
  8837=>"000000110",
  8838=>"010011110",
  8839=>"010010000",
  8840=>"100101001",
  8841=>"101111100",
  8842=>"011111001",
  8843=>"001010010",
  8844=>"011100111",
  8845=>"111111111",
  8846=>"011011001",
  8847=>"010110011",
  8848=>"010011101",
  8849=>"111010101",
  8850=>"000011100",
  8851=>"100111111",
  8852=>"001011110",
  8853=>"110101100",
  8854=>"110111000",
  8855=>"100111101",
  8856=>"000000110",
  8857=>"010100101",
  8858=>"100001011",
  8859=>"101010110",
  8860=>"100100010",
  8861=>"010010000",
  8862=>"100001110",
  8863=>"010000101",
  8864=>"111101001",
  8865=>"111101110",
  8866=>"001101111",
  8867=>"011100110",
  8868=>"010101000",
  8869=>"011011110",
  8870=>"101100100",
  8871=>"010001100",
  8872=>"011010010",
  8873=>"111001100",
  8874=>"010000101",
  8875=>"011100010",
  8876=>"110111010",
  8877=>"011010100",
  8878=>"111011011",
  8879=>"111111110",
  8880=>"111001101",
  8881=>"010100110",
  8882=>"001010000",
  8883=>"101110100",
  8884=>"011101010",
  8885=>"110101010",
  8886=>"111111001",
  8887=>"011101011",
  8888=>"001111101",
  8889=>"001000111",
  8890=>"101000000",
  8891=>"110101110",
  8892=>"100001011",
  8893=>"000100011",
  8894=>"000100010",
  8895=>"101001010",
  8896=>"011110011",
  8897=>"001011111",
  8898=>"000111001",
  8899=>"011000110",
  8900=>"011100111",
  8901=>"010011100",
  8902=>"101111011",
  8903=>"011111011",
  8904=>"100010111",
  8905=>"010111100",
  8906=>"010001001",
  8907=>"110101010",
  8908=>"000010011",
  8909=>"000000000",
  8910=>"001100011",
  8911=>"110001010",
  8912=>"101110001",
  8913=>"001010100",
  8914=>"010110101",
  8915=>"011101101",
  8916=>"101001011",
  8917=>"010010111",
  8918=>"000011001",
  8919=>"011100000",
  8920=>"000110010",
  8921=>"001010011",
  8922=>"100110000",
  8923=>"101010001",
  8924=>"001110111",
  8925=>"111101110",
  8926=>"111000101",
  8927=>"011101110",
  8928=>"101110111",
  8929=>"001101101",
  8930=>"100001001",
  8931=>"110010101",
  8932=>"010100000",
  8933=>"011011010",
  8934=>"110110101",
  8935=>"010100010",
  8936=>"100000111",
  8937=>"111000110",
  8938=>"111110111",
  8939=>"110011111",
  8940=>"000001000",
  8941=>"010101011",
  8942=>"010110011",
  8943=>"101001101",
  8944=>"000011111",
  8945=>"010001101",
  8946=>"100011110",
  8947=>"100101110",
  8948=>"101011000",
  8949=>"010000010",
  8950=>"010100110",
  8951=>"111110101",
  8952=>"011110111",
  8953=>"000010101",
  8954=>"101011000",
  8955=>"010101111",
  8956=>"011010101",
  8957=>"011110010",
  8958=>"111011110",
  8959=>"011011111",
  8960=>"111111110",
  8961=>"100001001",
  8962=>"101110110",
  8963=>"011101101",
  8964=>"010101110",
  8965=>"010011110",
  8966=>"110111111",
  8967=>"000011100",
  8968=>"001001111",
  8969=>"110111001",
  8970=>"101110111",
  8971=>"100100111",
  8972=>"000000101",
  8973=>"111011010",
  8974=>"000011001",
  8975=>"101010110",
  8976=>"000111001",
  8977=>"001001100",
  8978=>"010001111",
  8979=>"111010101",
  8980=>"110010001",
  8981=>"000001100",
  8982=>"101100101",
  8983=>"000011110",
  8984=>"111101100",
  8985=>"100101111",
  8986=>"101110001",
  8987=>"101001010",
  8988=>"111111011",
  8989=>"001110111",
  8990=>"110011011",
  8991=>"101111010",
  8992=>"001000001",
  8993=>"011011000",
  8994=>"000110110",
  8995=>"000100010",
  8996=>"010000001",
  8997=>"110000110",
  8998=>"001011000",
  8999=>"010001010",
  9000=>"100101100",
  9001=>"000001101",
  9002=>"111111111",
  9003=>"100001111",
  9004=>"011111010",
  9005=>"110100001",
  9006=>"101100000",
  9007=>"111111110",
  9008=>"001010100",
  9009=>"101101101",
  9010=>"100101110",
  9011=>"001011010",
  9012=>"010000101",
  9013=>"100111111",
  9014=>"000010000",
  9015=>"000111110",
  9016=>"011011001",
  9017=>"100010011",
  9018=>"110100110",
  9019=>"110000001",
  9020=>"010111110",
  9021=>"011001001",
  9022=>"011100110",
  9023=>"011111110",
  9024=>"000001010",
  9025=>"100100111",
  9026=>"011110010",
  9027=>"011110101",
  9028=>"100100101",
  9029=>"111111000",
  9030=>"001010000",
  9031=>"111100111",
  9032=>"010110001",
  9033=>"101010001",
  9034=>"010101011",
  9035=>"011100010",
  9036=>"001101001",
  9037=>"111011101",
  9038=>"111000000",
  9039=>"110111011",
  9040=>"001111101",
  9041=>"000110101",
  9042=>"111000100",
  9043=>"000000101",
  9044=>"111001101",
  9045=>"100000110",
  9046=>"000001110",
  9047=>"000000000",
  9048=>"011010011",
  9049=>"010100010",
  9050=>"110111111",
  9051=>"100000101",
  9052=>"011101110",
  9053=>"111110000",
  9054=>"001011110",
  9055=>"100110100",
  9056=>"000010001",
  9057=>"011001100",
  9058=>"010111010",
  9059=>"001011000",
  9060=>"001011101",
  9061=>"011111100",
  9062=>"000101010",
  9063=>"100011111",
  9064=>"001011000",
  9065=>"111101110",
  9066=>"011011110",
  9067=>"111010011",
  9068=>"100001100",
  9069=>"111111111",
  9070=>"010101111",
  9071=>"011110001",
  9072=>"001010010",
  9073=>"111111110",
  9074=>"111101001",
  9075=>"101011111",
  9076=>"110111000",
  9077=>"111000010",
  9078=>"111110011",
  9079=>"011100010",
  9080=>"100001100",
  9081=>"101001010",
  9082=>"010001101",
  9083=>"100001000",
  9084=>"000001001",
  9085=>"000111111",
  9086=>"111000100",
  9087=>"110011111",
  9088=>"001000000",
  9089=>"100010011",
  9090=>"000101011",
  9091=>"111001010",
  9092=>"110100110",
  9093=>"010010001",
  9094=>"011000100",
  9095=>"111100011",
  9096=>"110101101",
  9097=>"000000010",
  9098=>"111100110",
  9099=>"110100101",
  9100=>"101100011",
  9101=>"001000010",
  9102=>"110110111",
  9103=>"111001100",
  9104=>"101010001",
  9105=>"110101000",
  9106=>"000001100",
  9107=>"111110100",
  9108=>"000111010",
  9109=>"110101101",
  9110=>"101011111",
  9111=>"011001110",
  9112=>"001000110",
  9113=>"011101100",
  9114=>"111011111",
  9115=>"000011001",
  9116=>"111011110",
  9117=>"110100000",
  9118=>"100010000",
  9119=>"010101101",
  9120=>"001000111",
  9121=>"111011010",
  9122=>"000001101",
  9123=>"110100000",
  9124=>"010010111",
  9125=>"110001010",
  9126=>"010100011",
  9127=>"011101100",
  9128=>"100100101",
  9129=>"010101010",
  9130=>"001111101",
  9131=>"000101111",
  9132=>"010011101",
  9133=>"001111011",
  9134=>"101110100",
  9135=>"000100011",
  9136=>"110101110",
  9137=>"100010000",
  9138=>"001101100",
  9139=>"010101100",
  9140=>"011111111",
  9141=>"111100011",
  9142=>"010111110",
  9143=>"100111110",
  9144=>"111001010",
  9145=>"001100010",
  9146=>"110110001",
  9147=>"101110110",
  9148=>"100000000",
  9149=>"100000000",
  9150=>"110101000",
  9151=>"010000101",
  9152=>"000101000",
  9153=>"010010001",
  9154=>"000100011",
  9155=>"101110110",
  9156=>"110000100",
  9157=>"010101110",
  9158=>"111000011",
  9159=>"010010111",
  9160=>"011011100",
  9161=>"001101111",
  9162=>"111001101",
  9163=>"100110111",
  9164=>"010001011",
  9165=>"111101011",
  9166=>"000100001",
  9167=>"011101011",
  9168=>"101110100",
  9169=>"011111101",
  9170=>"000010101",
  9171=>"011001000",
  9172=>"000110000",
  9173=>"111000101",
  9174=>"000011100",
  9175=>"000011111",
  9176=>"101010100",
  9177=>"001011010",
  9178=>"001011001",
  9179=>"111110010",
  9180=>"101011110",
  9181=>"110011101",
  9182=>"111111101",
  9183=>"111010110",
  9184=>"110100100",
  9185=>"000000110",
  9186=>"000100001",
  9187=>"111100111",
  9188=>"010001101",
  9189=>"111101000",
  9190=>"110011100",
  9191=>"100000110",
  9192=>"000001101",
  9193=>"010100010",
  9194=>"000010101",
  9195=>"100011010",
  9196=>"000001110",
  9197=>"011001111",
  9198=>"010010110",
  9199=>"111100101",
  9200=>"110010101",
  9201=>"111101100",
  9202=>"011001001",
  9203=>"100111001",
  9204=>"110111111",
  9205=>"000011010",
  9206=>"000100000",
  9207=>"010100011",
  9208=>"111110100",
  9209=>"110010011",
  9210=>"111111011",
  9211=>"010010111",
  9212=>"010001001",
  9213=>"010100000",
  9214=>"001111011",
  9215=>"010011010",
  9216=>"110001110",
  9217=>"100100000",
  9218=>"001110010",
  9219=>"101111011",
  9220=>"000011111",
  9221=>"000010001",
  9222=>"101101101",
  9223=>"001001010",
  9224=>"010010001",
  9225=>"000000001",
  9226=>"011100001",
  9227=>"111010010",
  9228=>"000011011",
  9229=>"111101111",
  9230=>"010101111",
  9231=>"001011000",
  9232=>"110110110",
  9233=>"101101000",
  9234=>"110101101",
  9235=>"001001110",
  9236=>"001101000",
  9237=>"000100111",
  9238=>"101010001",
  9239=>"110001110",
  9240=>"100000111",
  9241=>"010111010",
  9242=>"111010110",
  9243=>"010111110",
  9244=>"010111100",
  9245=>"101111010",
  9246=>"000010101",
  9247=>"101111100",
  9248=>"010011111",
  9249=>"010111001",
  9250=>"011000000",
  9251=>"001001111",
  9252=>"000001101",
  9253=>"111001010",
  9254=>"001101000",
  9255=>"111101010",
  9256=>"011100011",
  9257=>"011001111",
  9258=>"100000010",
  9259=>"000100111",
  9260=>"000100010",
  9261=>"010101011",
  9262=>"101111001",
  9263=>"001101000",
  9264=>"011010111",
  9265=>"011111000",
  9266=>"001111110",
  9267=>"010110001",
  9268=>"110111010",
  9269=>"100001101",
  9270=>"110111011",
  9271=>"011110000",
  9272=>"000000001",
  9273=>"011110000",
  9274=>"110110101",
  9275=>"011110110",
  9276=>"000100001",
  9277=>"110100010",
  9278=>"111011000",
  9279=>"001100011",
  9280=>"100110111",
  9281=>"111000111",
  9282=>"010000010",
  9283=>"000110100",
  9284=>"011001110",
  9285=>"000000110",
  9286=>"010100010",
  9287=>"100110111",
  9288=>"000011100",
  9289=>"011001011",
  9290=>"110001101",
  9291=>"110101111",
  9292=>"110110100",
  9293=>"011101011",
  9294=>"010011100",
  9295=>"101011000",
  9296=>"010100101",
  9297=>"000010011",
  9298=>"010000001",
  9299=>"100011001",
  9300=>"100000100",
  9301=>"000001011",
  9302=>"010011011",
  9303=>"000000010",
  9304=>"010100001",
  9305=>"000100101",
  9306=>"111011000",
  9307=>"100110110",
  9308=>"000000001",
  9309=>"100110000",
  9310=>"110000000",
  9311=>"010100100",
  9312=>"011011100",
  9313=>"110101011",
  9314=>"111100111",
  9315=>"011100010",
  9316=>"100110011",
  9317=>"000111100",
  9318=>"001101011",
  9319=>"000010110",
  9320=>"111010011",
  9321=>"001000001",
  9322=>"110110110",
  9323=>"111100110",
  9324=>"101000011",
  9325=>"001100010",
  9326=>"001001000",
  9327=>"011010001",
  9328=>"110110001",
  9329=>"001010000",
  9330=>"000010000",
  9331=>"110001110",
  9332=>"001010110",
  9333=>"010111101",
  9334=>"011110100",
  9335=>"111001011",
  9336=>"001011101",
  9337=>"101011100",
  9338=>"000010000",
  9339=>"001100100",
  9340=>"000010111",
  9341=>"010100010",
  9342=>"010110110",
  9343=>"010010010",
  9344=>"110101111",
  9345=>"000010000",
  9346=>"101100100",
  9347=>"011011101",
  9348=>"001000101",
  9349=>"001001000",
  9350=>"000000010",
  9351=>"011010100",
  9352=>"110111000",
  9353=>"000110101",
  9354=>"000001101",
  9355=>"101101001",
  9356=>"000001110",
  9357=>"010111001",
  9358=>"000011010",
  9359=>"100001101",
  9360=>"111001010",
  9361=>"111110011",
  9362=>"011111111",
  9363=>"011001101",
  9364=>"011100101",
  9365=>"111101110",
  9366=>"110001111",
  9367=>"010000001",
  9368=>"000010010",
  9369=>"100001000",
  9370=>"001111001",
  9371=>"001011011",
  9372=>"101011101",
  9373=>"000110001",
  9374=>"001000111",
  9375=>"101101011",
  9376=>"011000011",
  9377=>"011001010",
  9378=>"010000111",
  9379=>"000001000",
  9380=>"000010110",
  9381=>"000001011",
  9382=>"000110101",
  9383=>"101000001",
  9384=>"101011100",
  9385=>"011110101",
  9386=>"000100000",
  9387=>"010011111",
  9388=>"101000111",
  9389=>"110111101",
  9390=>"010110001",
  9391=>"111010110",
  9392=>"111111100",
  9393=>"000000100",
  9394=>"000000001",
  9395=>"011010001",
  9396=>"100111010",
  9397=>"111101111",
  9398=>"111011001",
  9399=>"001000101",
  9400=>"001010101",
  9401=>"110001100",
  9402=>"111000000",
  9403=>"001010000",
  9404=>"010101001",
  9405=>"101010101",
  9406=>"100010010",
  9407=>"110001000",
  9408=>"000000100",
  9409=>"010111100",
  9410=>"011001001",
  9411=>"000011110",
  9412=>"011101000",
  9413=>"111100110",
  9414=>"010000111",
  9415=>"001111011",
  9416=>"111011101",
  9417=>"100100111",
  9418=>"101000111",
  9419=>"001001100",
  9420=>"011001000",
  9421=>"111001111",
  9422=>"111111010",
  9423=>"010100011",
  9424=>"010000100",
  9425=>"000011111",
  9426=>"011100111",
  9427=>"010100000",
  9428=>"011101001",
  9429=>"010100100",
  9430=>"001101001",
  9431=>"000111110",
  9432=>"111011110",
  9433=>"110010000",
  9434=>"100111100",
  9435=>"111000110",
  9436=>"001001000",
  9437=>"110110110",
  9438=>"000100011",
  9439=>"111101010",
  9440=>"001000101",
  9441=>"110101011",
  9442=>"100010000",
  9443=>"011001100",
  9444=>"011101101",
  9445=>"101011101",
  9446=>"000001000",
  9447=>"110010101",
  9448=>"111100010",
  9449=>"001110101",
  9450=>"100011100",
  9451=>"011110100",
  9452=>"001100001",
  9453=>"011111011",
  9454=>"101011001",
  9455=>"100000011",
  9456=>"001001001",
  9457=>"000111101",
  9458=>"101101111",
  9459=>"010101001",
  9460=>"001101001",
  9461=>"000100101",
  9462=>"000100000",
  9463=>"111110111",
  9464=>"111100010",
  9465=>"011110000",
  9466=>"010111011",
  9467=>"000100100",
  9468=>"001101000",
  9469=>"000101001",
  9470=>"000010010",
  9471=>"001110100",
  9472=>"010011111",
  9473=>"101000001",
  9474=>"110001000",
  9475=>"011101111",
  9476=>"000010001",
  9477=>"010001010",
  9478=>"010000110",
  9479=>"111110001",
  9480=>"110111110",
  9481=>"001001111",
  9482=>"101110100",
  9483=>"110101011",
  9484=>"110000111",
  9485=>"100000010",
  9486=>"011010100",
  9487=>"000001001",
  9488=>"101111101",
  9489=>"001011010",
  9490=>"111100001",
  9491=>"011000110",
  9492=>"111111101",
  9493=>"000100100",
  9494=>"000100111",
  9495=>"101000111",
  9496=>"001010011",
  9497=>"111000100",
  9498=>"111110010",
  9499=>"010101100",
  9500=>"110001010",
  9501=>"101100110",
  9502=>"110111111",
  9503=>"010111001",
  9504=>"100010111",
  9505=>"101010010",
  9506=>"011101001",
  9507=>"100000100",
  9508=>"011111001",
  9509=>"011000001",
  9510=>"101000010",
  9511=>"011100000",
  9512=>"100001100",
  9513=>"010111110",
  9514=>"111100111",
  9515=>"010000111",
  9516=>"010111000",
  9517=>"101100001",
  9518=>"110110100",
  9519=>"000011000",
  9520=>"001000001",
  9521=>"111011111",
  9522=>"111100111",
  9523=>"010101110",
  9524=>"110100110",
  9525=>"011101111",
  9526=>"110010111",
  9527=>"000110111",
  9528=>"101100101",
  9529=>"011000111",
  9530=>"101001110",
  9531=>"100101000",
  9532=>"110000110",
  9533=>"101101110",
  9534=>"100100000",
  9535=>"111101000",
  9536=>"001000000",
  9537=>"011001011",
  9538=>"100010010",
  9539=>"101001001",
  9540=>"001000001",
  9541=>"111101011",
  9542=>"000000101",
  9543=>"101100111",
  9544=>"001100010",
  9545=>"001000110",
  9546=>"001001110",
  9547=>"000100100",
  9548=>"000010001",
  9549=>"010101001",
  9550=>"001101010",
  9551=>"110011100",
  9552=>"110010110",
  9553=>"101110001",
  9554=>"101000000",
  9555=>"110111001",
  9556=>"001011100",
  9557=>"001100000",
  9558=>"110111010",
  9559=>"001011100",
  9560=>"100001010",
  9561=>"000010011",
  9562=>"000101001",
  9563=>"000000010",
  9564=>"111011101",
  9565=>"010100111",
  9566=>"100011101",
  9567=>"100001101",
  9568=>"100001111",
  9569=>"111000111",
  9570=>"111100000",
  9571=>"000111001",
  9572=>"110100001",
  9573=>"011000000",
  9574=>"000100010",
  9575=>"110001110",
  9576=>"100010111",
  9577=>"000110100",
  9578=>"000110110",
  9579=>"000010001",
  9580=>"101001010",
  9581=>"111101010",
  9582=>"011110110",
  9583=>"001011001",
  9584=>"111001101",
  9585=>"011010000",
  9586=>"111111001",
  9587=>"001010001",
  9588=>"101110110",
  9589=>"001010110",
  9590=>"100100100",
  9591=>"000100101",
  9592=>"101110011",
  9593=>"110111011",
  9594=>"000100001",
  9595=>"111111000",
  9596=>"000010111",
  9597=>"111001010",
  9598=>"100001010",
  9599=>"111110001",
  9600=>"001111111",
  9601=>"001011100",
  9602=>"010101100",
  9603=>"101101101",
  9604=>"011101001",
  9605=>"010001000",
  9606=>"000101010",
  9607=>"011110101",
  9608=>"111011011",
  9609=>"000011101",
  9610=>"011010111",
  9611=>"110111011",
  9612=>"000101101",
  9613=>"011001010",
  9614=>"000001011",
  9615=>"111101000",
  9616=>"010100111",
  9617=>"000101011",
  9618=>"101001100",
  9619=>"111110011",
  9620=>"110100110",
  9621=>"000010100",
  9622=>"101110010",
  9623=>"000011111",
  9624=>"111111010",
  9625=>"011001001",
  9626=>"110110110",
  9627=>"000010110",
  9628=>"010100001",
  9629=>"000110001",
  9630=>"101001000",
  9631=>"100101011",
  9632=>"100000000",
  9633=>"101110011",
  9634=>"001110111",
  9635=>"010100011",
  9636=>"110011001",
  9637=>"010111100",
  9638=>"101010111",
  9639=>"010000011",
  9640=>"111110110",
  9641=>"010101111",
  9642=>"001100101",
  9643=>"000101101",
  9644=>"001010111",
  9645=>"000100010",
  9646=>"011100110",
  9647=>"101100010",
  9648=>"001110001",
  9649=>"000110110",
  9650=>"011110101",
  9651=>"101011000",
  9652=>"000011001",
  9653=>"111100111",
  9654=>"000000101",
  9655=>"000001111",
  9656=>"111111010",
  9657=>"110111111",
  9658=>"001011000",
  9659=>"101101111",
  9660=>"101101011",
  9661=>"110110000",
  9662=>"111101000",
  9663=>"001010000",
  9664=>"100001111",
  9665=>"001011111",
  9666=>"111110111",
  9667=>"100010000",
  9668=>"000100100",
  9669=>"010001001",
  9670=>"111011011",
  9671=>"011111010",
  9672=>"011100000",
  9673=>"010101101",
  9674=>"010111011",
  9675=>"011110001",
  9676=>"110111111",
  9677=>"100001101",
  9678=>"000010001",
  9679=>"110001011",
  9680=>"110111110",
  9681=>"100110000",
  9682=>"001010011",
  9683=>"011110111",
  9684=>"000011011",
  9685=>"001000111",
  9686=>"000100001",
  9687=>"110010110",
  9688=>"100110010",
  9689=>"010000101",
  9690=>"101110000",
  9691=>"110000010",
  9692=>"001100100",
  9693=>"101001111",
  9694=>"011111110",
  9695=>"010100011",
  9696=>"100010100",
  9697=>"011001010",
  9698=>"111001001",
  9699=>"110101101",
  9700=>"011001001",
  9701=>"001000011",
  9702=>"011100000",
  9703=>"101100010",
  9704=>"000001010",
  9705=>"111011110",
  9706=>"011111000",
  9707=>"000000110",
  9708=>"111000111",
  9709=>"110010110",
  9710=>"110001010",
  9711=>"011101011",
  9712=>"010111011",
  9713=>"111101011",
  9714=>"011011010",
  9715=>"011100011",
  9716=>"010001110",
  9717=>"010010000",
  9718=>"101111111",
  9719=>"110010100",
  9720=>"011101111",
  9721=>"001000100",
  9722=>"111010010",
  9723=>"100110100",
  9724=>"110001001",
  9725=>"111101010",
  9726=>"101010001",
  9727=>"101011011",
  9728=>"000010000",
  9729=>"100110111",
  9730=>"000110111",
  9731=>"101110110",
  9732=>"111011010",
  9733=>"110110111",
  9734=>"111111100",
  9735=>"100100111",
  9736=>"010110111",
  9737=>"000100001",
  9738=>"000100100",
  9739=>"011111000",
  9740=>"010011110",
  9741=>"100111101",
  9742=>"101000000",
  9743=>"001000110",
  9744=>"101001111",
  9745=>"001010000",
  9746=>"000101000",
  9747=>"100111011",
  9748=>"011101000",
  9749=>"001111000",
  9750=>"010111000",
  9751=>"110101010",
  9752=>"100011010",
  9753=>"001101000",
  9754=>"001000110",
  9755=>"000110110",
  9756=>"001110111",
  9757=>"011100011",
  9758=>"011101110",
  9759=>"010100101",
  9760=>"111001011",
  9761=>"111000010",
  9762=>"110001000",
  9763=>"110100011",
  9764=>"011001111",
  9765=>"010001011",
  9766=>"001111110",
  9767=>"011111111",
  9768=>"100000110",
  9769=>"100010000",
  9770=>"001000100",
  9771=>"011010011",
  9772=>"011110011",
  9773=>"110110111",
  9774=>"011011011",
  9775=>"101001000",
  9776=>"010000000",
  9777=>"111000010",
  9778=>"110100101",
  9779=>"000000110",
  9780=>"001011001",
  9781=>"111000001",
  9782=>"010000011",
  9783=>"111011101",
  9784=>"010001110",
  9785=>"110110110",
  9786=>"001010111",
  9787=>"111100101",
  9788=>"110111011",
  9789=>"000000110",
  9790=>"000100110",
  9791=>"011111000",
  9792=>"101010011",
  9793=>"110010100",
  9794=>"100000101",
  9795=>"000100100",
  9796=>"011111100",
  9797=>"011100011",
  9798=>"001010011",
  9799=>"100111101",
  9800=>"011011001",
  9801=>"010001110",
  9802=>"011110111",
  9803=>"101001111",
  9804=>"000010110",
  9805=>"011011010",
  9806=>"111011011",
  9807=>"111011101",
  9808=>"111101110",
  9809=>"011001010",
  9810=>"111100110",
  9811=>"111100000",
  9812=>"110110111",
  9813=>"010001100",
  9814=>"000000101",
  9815=>"011101101",
  9816=>"111011100",
  9817=>"001100100",
  9818=>"001100101",
  9819=>"010101101",
  9820=>"011100110",
  9821=>"100010110",
  9822=>"000011001",
  9823=>"011100110",
  9824=>"100001001",
  9825=>"000001110",
  9826=>"101001011",
  9827=>"111010011",
  9828=>"001110111",
  9829=>"111001000",
  9830=>"100111111",
  9831=>"110111111",
  9832=>"110010001",
  9833=>"001011001",
  9834=>"001100010",
  9835=>"100110010",
  9836=>"010100111",
  9837=>"000001001",
  9838=>"010110000",
  9839=>"001101101",
  9840=>"101101000",
  9841=>"110111110",
  9842=>"010001111",
  9843=>"101101001",
  9844=>"010001101",
  9845=>"110000100",
  9846=>"000011011",
  9847=>"101000001",
  9848=>"110110010",
  9849=>"111111101",
  9850=>"100011111",
  9851=>"001011110",
  9852=>"010101011",
  9853=>"011100000",
  9854=>"001101011",
  9855=>"100010000",
  9856=>"000011011",
  9857=>"011001110",
  9858=>"101100101",
  9859=>"000001000",
  9860=>"011101111",
  9861=>"010111101",
  9862=>"100101100",
  9863=>"010111110",
  9864=>"000010101",
  9865=>"011010000",
  9866=>"001010101",
  9867=>"011101010",
  9868=>"000110111",
  9869=>"000000101",
  9870=>"011001111",
  9871=>"000001101",
  9872=>"100101111",
  9873=>"111110010",
  9874=>"010110001",
  9875=>"001111010",
  9876=>"001011101",
  9877=>"111011110",
  9878=>"001101101",
  9879=>"100110000",
  9880=>"011011101",
  9881=>"000000000",
  9882=>"010110111",
  9883=>"110001101",
  9884=>"000100111",
  9885=>"011011110",
  9886=>"101101110",
  9887=>"100000001",
  9888=>"110000000",
  9889=>"001110111",
  9890=>"000001110",
  9891=>"000111010",
  9892=>"001001001",
  9893=>"111111111",
  9894=>"000000001",
  9895=>"001001100",
  9896=>"101001100",
  9897=>"000111110",
  9898=>"110101011",
  9899=>"011100010",
  9900=>"001010100",
  9901=>"010010100",
  9902=>"101100011",
  9903=>"100001000",
  9904=>"000110001",
  9905=>"110110101",
  9906=>"011100110",
  9907=>"011100001",
  9908=>"000011010",
  9909=>"101111100",
  9910=>"100110000",
  9911=>"100011110",
  9912=>"011110101",
  9913=>"000110111",
  9914=>"110001010",
  9915=>"100100101",
  9916=>"000000000",
  9917=>"011011110",
  9918=>"010100011",
  9919=>"000000111",
  9920=>"110000100",
  9921=>"101100100",
  9922=>"111110101",
  9923=>"110011110",
  9924=>"010000101",
  9925=>"111110000",
  9926=>"001000010",
  9927=>"100111100",
  9928=>"100011000",
  9929=>"100010011",
  9930=>"110111101",
  9931=>"100100110",
  9932=>"111011000",
  9933=>"001011111",
  9934=>"100100110",
  9935=>"101110010",
  9936=>"011001001",
  9937=>"100111101",
  9938=>"110011111",
  9939=>"101100011",
  9940=>"010010110",
  9941=>"000110000",
  9942=>"011110011",
  9943=>"000110000",
  9944=>"111111011",
  9945=>"100101100",
  9946=>"101110101",
  9947=>"011000000",
  9948=>"110100101",
  9949=>"101000011",
  9950=>"010011000",
  9951=>"001100101",
  9952=>"001011000",
  9953=>"011011001",
  9954=>"001011010",
  9955=>"010010100",
  9956=>"001110110",
  9957=>"010100110",
  9958=>"001110100",
  9959=>"110100001",
  9960=>"110000010",
  9961=>"100011111",
  9962=>"101111010",
  9963=>"010000110",
  9964=>"000001111",
  9965=>"000001001",
  9966=>"010010111",
  9967=>"110010001",
  9968=>"010111101",
  9969=>"011010000",
  9970=>"010011100",
  9971=>"111010000",
  9972=>"101011111",
  9973=>"111100101",
  9974=>"110111011",
  9975=>"111100011",
  9976=>"100010111",
  9977=>"001111100",
  9978=>"110000011",
  9979=>"010010110",
  9980=>"010111110",
  9981=>"011000110",
  9982=>"000110101",
  9983=>"011101011",
  9984=>"000001010",
  9985=>"110111010",
  9986=>"110110100",
  9987=>"000001010",
  9988=>"000111011",
  9989=>"000001000",
  9990=>"010001100",
  9991=>"011000010",
  9992=>"010011101",
  9993=>"001101011",
  9994=>"010011001",
  9995=>"111101000",
  9996=>"110100101",
  9997=>"011110100",
  9998=>"101110010",
  9999=>"011111110",
  10000=>"000001001",
  10001=>"101010101",
  10002=>"011111011",
  10003=>"100110110",
  10004=>"100110010",
  10005=>"010010001",
  10006=>"000001110",
  10007=>"110100001",
  10008=>"101110000",
  10009=>"010011001",
  10010=>"110010111",
  10011=>"110000000",
  10012=>"101100000",
  10013=>"110110001",
  10014=>"000010000",
  10015=>"101000110",
  10016=>"001011110",
  10017=>"110101011",
  10018=>"010011111",
  10019=>"011111101",
  10020=>"010111010",
  10021=>"111000100",
  10022=>"111001100",
  10023=>"001001011",
  10024=>"010110000",
  10025=>"100110110",
  10026=>"111001000",
  10027=>"111111110",
  10028=>"011000001",
  10029=>"101110001",
  10030=>"001010010",
  10031=>"000010011",
  10032=>"000010010",
  10033=>"001111010",
  10034=>"100110000",
  10035=>"110111100",
  10036=>"000101000",
  10037=>"101010010",
  10038=>"010000010",
  10039=>"111010011",
  10040=>"110101100",
  10041=>"111101000",
  10042=>"111001111",
  10043=>"000011010",
  10044=>"001100101",
  10045=>"111111000",
  10046=>"011101111",
  10047=>"100101011",
  10048=>"011111101",
  10049=>"010111001",
  10050=>"010101111",
  10051=>"010011110",
  10052=>"101010110",
  10053=>"110010100",
  10054=>"101000110",
  10055=>"101111000",
  10056=>"101101010",
  10057=>"111101110",
  10058=>"001010010",
  10059=>"110010111",
  10060=>"001110111",
  10061=>"100111110",
  10062=>"101101101",
  10063=>"100111000",
  10064=>"111000010",
  10065=>"011111000",
  10066=>"010010001",
  10067=>"101011101",
  10068=>"110110001",
  10069=>"011001001",
  10070=>"111010010",
  10071=>"110101111",
  10072=>"001000101",
  10073=>"100001111",
  10074=>"010010100",
  10075=>"101001101",
  10076=>"011001011",
  10077=>"101000110",
  10078=>"110101100",
  10079=>"000110110",
  10080=>"101011010",
  10081=>"100101010",
  10082=>"111100001",
  10083=>"111111011",
  10084=>"110001000",
  10085=>"101111111",
  10086=>"001001000",
  10087=>"010011101",
  10088=>"000000000",
  10089=>"011101010",
  10090=>"101000111",
  10091=>"100100101",
  10092=>"000001000",
  10093=>"101111010",
  10094=>"001100111",
  10095=>"010010001",
  10096=>"001001000",
  10097=>"101011011",
  10098=>"001110000",
  10099=>"010110010",
  10100=>"011010000",
  10101=>"001001001",
  10102=>"000110011",
  10103=>"001101111",
  10104=>"000111011",
  10105=>"100001111",
  10106=>"000000101",
  10107=>"101101110",
  10108=>"011110001",
  10109=>"111101100",
  10110=>"000010011",
  10111=>"100000001",
  10112=>"001001111",
  10113=>"110100110",
  10114=>"111001001",
  10115=>"110000001",
  10116=>"100110110",
  10117=>"110010100",
  10118=>"111100111",
  10119=>"001110010",
  10120=>"001101110",
  10121=>"101001010",
  10122=>"100010000",
  10123=>"101111000",
  10124=>"000011001",
  10125=>"101000011",
  10126=>"000001001",
  10127=>"110010001",
  10128=>"000001001",
  10129=>"011001110",
  10130=>"001100101",
  10131=>"000100011",
  10132=>"110111001",
  10133=>"110001110",
  10134=>"111111000",
  10135=>"010001001",
  10136=>"001001001",
  10137=>"010110001",
  10138=>"101100101",
  10139=>"011011011",
  10140=>"100010101",
  10141=>"000100001",
  10142=>"101011110",
  10143=>"001110101",
  10144=>"100100101",
  10145=>"101100001",
  10146=>"100111111",
  10147=>"101010001",
  10148=>"001100110",
  10149=>"101111010",
  10150=>"001110100",
  10151=>"111011010",
  10152=>"111111011",
  10153=>"011101110",
  10154=>"101110000",
  10155=>"000010000",
  10156=>"011001011",
  10157=>"100001101",
  10158=>"011010100",
  10159=>"111001101",
  10160=>"101100100",
  10161=>"000001111",
  10162=>"001011011",
  10163=>"011001110",
  10164=>"100010011",
  10165=>"011100111",
  10166=>"110001100",
  10167=>"101110000",
  10168=>"111011110",
  10169=>"111101101",
  10170=>"100110110",
  10171=>"110101111",
  10172=>"111110010",
  10173=>"010110000",
  10174=>"001110001",
  10175=>"000111001",
  10176=>"101001000",
  10177=>"111111111",
  10178=>"011110001",
  10179=>"110111011",
  10180=>"101110001",
  10181=>"001100100",
  10182=>"101101010",
  10183=>"100101000",
  10184=>"001010100",
  10185=>"001110010",
  10186=>"010101111",
  10187=>"000111111",
  10188=>"110000111",
  10189=>"101000111",
  10190=>"101101110",
  10191=>"001101001",
  10192=>"010010101",
  10193=>"111111001",
  10194=>"111000001",
  10195=>"101111111",
  10196=>"001001010",
  10197=>"100100100",
  10198=>"000111110",
  10199=>"001111111",
  10200=>"001011001",
  10201=>"001100000",
  10202=>"010011011",
  10203=>"111111001",
  10204=>"010110111",
  10205=>"110101001",
  10206=>"111010101",
  10207=>"011111011",
  10208=>"110000100",
  10209=>"110101010",
  10210=>"001010100",
  10211=>"101010111",
  10212=>"101011000",
  10213=>"101001110",
  10214=>"001011101",
  10215=>"000100101",
  10216=>"100100011",
  10217=>"011010100",
  10218=>"110101010",
  10219=>"010001011",
  10220=>"100100011",
  10221=>"001001100",
  10222=>"101111001",
  10223=>"101000110",
  10224=>"100111000",
  10225=>"000111001",
  10226=>"100100110",
  10227=>"101001010",
  10228=>"101010000",
  10229=>"011100001",
  10230=>"000101100",
  10231=>"110111110",
  10232=>"000100001",
  10233=>"110000110",
  10234=>"101010011",
  10235=>"101111100",
  10236=>"111000011",
  10237=>"100100001",
  10238=>"001101000",
  10239=>"100000101",
  10240=>"110001000",
  10241=>"110111011",
  10242=>"101100000",
  10243=>"101100000",
  10244=>"111101001",
  10245=>"101001100",
  10246=>"001011011",
  10247=>"110110111",
  10248=>"001001100",
  10249=>"110110000",
  10250=>"101000100",
  10251=>"111100000",
  10252=>"011010000",
  10253=>"000110101",
  10254=>"010010100",
  10255=>"101000010",
  10256=>"100110011",
  10257=>"100001111",
  10258=>"000100011",
  10259=>"011011001",
  10260=>"110101001",
  10261=>"011100001",
  10262=>"010010110",
  10263=>"101110100",
  10264=>"010100011",
  10265=>"110011011",
  10266=>"111101001",
  10267=>"101111001",
  10268=>"101010111",
  10269=>"001001100",
  10270=>"000011110",
  10271=>"001010111",
  10272=>"101110110",
  10273=>"010100001",
  10274=>"101001110",
  10275=>"110100100",
  10276=>"100111011",
  10277=>"010010111",
  10278=>"000001010",
  10279=>"001100011",
  10280=>"000000001",
  10281=>"111111010",
  10282=>"010111111",
  10283=>"101111010",
  10284=>"000000101",
  10285=>"100010001",
  10286=>"100100001",
  10287=>"111101100",
  10288=>"100101001",
  10289=>"111011111",
  10290=>"111000010",
  10291=>"101000000",
  10292=>"101011010",
  10293=>"101111100",
  10294=>"101000001",
  10295=>"011001100",
  10296=>"011010110",
  10297=>"100101100",
  10298=>"011111001",
  10299=>"001000000",
  10300=>"001001100",
  10301=>"001100010",
  10302=>"101101001",
  10303=>"110111000",
  10304=>"111101011",
  10305=>"101001110",
  10306=>"100110010",
  10307=>"000111000",
  10308=>"011010010",
  10309=>"100101101",
  10310=>"110110110",
  10311=>"111100100",
  10312=>"000001101",
  10313=>"011110100",
  10314=>"001011110",
  10315=>"011010101",
  10316=>"111111110",
  10317=>"101011011",
  10318=>"101010011",
  10319=>"011101111",
  10320=>"101101100",
  10321=>"001000111",
  10322=>"111110111",
  10323=>"100011011",
  10324=>"011000101",
  10325=>"100000000",
  10326=>"111010110",
  10327=>"000001010",
  10328=>"000111101",
  10329=>"101111010",
  10330=>"110110001",
  10331=>"000000101",
  10332=>"111000010",
  10333=>"101010011",
  10334=>"101001100",
  10335=>"011110101",
  10336=>"100101111",
  10337=>"011111011",
  10338=>"010011101",
  10339=>"011110000",
  10340=>"101011101",
  10341=>"001011110",
  10342=>"001101100",
  10343=>"101111100",
  10344=>"010001000",
  10345=>"111100111",
  10346=>"001001001",
  10347=>"110101010",
  10348=>"011010000",
  10349=>"111000011",
  10350=>"011110011",
  10351=>"010010100",
  10352=>"000101101",
  10353=>"011100001",
  10354=>"111100010",
  10355=>"000110010",
  10356=>"011110011",
  10357=>"111011101",
  10358=>"100011000",
  10359=>"100011001",
  10360=>"100111001",
  10361=>"010110110",
  10362=>"000011000",
  10363=>"010110100",
  10364=>"100110100",
  10365=>"100110010",
  10366=>"001000100",
  10367=>"101110011",
  10368=>"101110101",
  10369=>"011100000",
  10370=>"101001101",
  10371=>"111001011",
  10372=>"011010100",
  10373=>"111100001",
  10374=>"010011010",
  10375=>"000101011",
  10376=>"100001010",
  10377=>"101001100",
  10378=>"111100100",
  10379=>"111110111",
  10380=>"011100010",
  10381=>"101011010",
  10382=>"010001010",
  10383=>"110000000",
  10384=>"000100111",
  10385=>"000001110",
  10386=>"100111010",
  10387=>"010001100",
  10388=>"001110101",
  10389=>"111101101",
  10390=>"110000110",
  10391=>"000100100",
  10392=>"100100001",
  10393=>"000001000",
  10394=>"011100100",
  10395=>"000110010",
  10396=>"111001101",
  10397=>"000010111",
  10398=>"000000110",
  10399=>"011011010",
  10400=>"011000001",
  10401=>"101001011",
  10402=>"101100001",
  10403=>"110000000",
  10404=>"011001010",
  10405=>"001100010",
  10406=>"101000101",
  10407=>"110010110",
  10408=>"110011111",
  10409=>"100011101",
  10410=>"010111000",
  10411=>"000111011",
  10412=>"111111011",
  10413=>"111110110",
  10414=>"111001010",
  10415=>"010011100",
  10416=>"000101111",
  10417=>"110001010",
  10418=>"001010100",
  10419=>"110001001",
  10420=>"010110101",
  10421=>"000001001",
  10422=>"010010010",
  10423=>"100000010",
  10424=>"101100011",
  10425=>"001001000",
  10426=>"011110000",
  10427=>"110101111",
  10428=>"110110010",
  10429=>"101001011",
  10430=>"011000000",
  10431=>"110001111",
  10432=>"101001001",
  10433=>"110110010",
  10434=>"100110111",
  10435=>"101111100",
  10436=>"101100011",
  10437=>"110100010",
  10438=>"000000111",
  10439=>"101100010",
  10440=>"000110001",
  10441=>"010101100",
  10442=>"110011001",
  10443=>"111111110",
  10444=>"111101110",
  10445=>"010110101",
  10446=>"100000100",
  10447=>"011111111",
  10448=>"100111000",
  10449=>"110011000",
  10450=>"110011011",
  10451=>"001000001",
  10452=>"001111101",
  10453=>"011011010",
  10454=>"001111110",
  10455=>"000101110",
  10456=>"111010100",
  10457=>"011001101",
  10458=>"100101000",
  10459=>"111010110",
  10460=>"001011010",
  10461=>"010100001",
  10462=>"001001010",
  10463=>"011000000",
  10464=>"111011001",
  10465=>"011000101",
  10466=>"011101111",
  10467=>"110111110",
  10468=>"011100111",
  10469=>"100100100",
  10470=>"011000001",
  10471=>"110000101",
  10472=>"011111010",
  10473=>"010001110",
  10474=>"010000110",
  10475=>"001010110",
  10476=>"110101000",
  10477=>"001101010",
  10478=>"110011101",
  10479=>"101111111",
  10480=>"000001000",
  10481=>"001000000",
  10482=>"101001010",
  10483=>"100000110",
  10484=>"001000110",
  10485=>"001110000",
  10486=>"010100110",
  10487=>"100100010",
  10488=>"011000010",
  10489=>"000101110",
  10490=>"010111000",
  10491=>"101000011",
  10492=>"011001100",
  10493=>"100101100",
  10494=>"010001011",
  10495=>"000000111",
  10496=>"101110111",
  10497=>"001101001",
  10498=>"101000100",
  10499=>"101011011",
  10500=>"001110110",
  10501=>"111110101",
  10502=>"000000000",
  10503=>"011010111",
  10504=>"111001110",
  10505=>"010110100",
  10506=>"001010011",
  10507=>"010011111",
  10508=>"010011100",
  10509=>"100101000",
  10510=>"011110011",
  10511=>"111010101",
  10512=>"111101011",
  10513=>"111100101",
  10514=>"001010111",
  10515=>"001011011",
  10516=>"011101001",
  10517=>"001000110",
  10518=>"100001001",
  10519=>"100101100",
  10520=>"000111101",
  10521=>"001010101",
  10522=>"000000000",
  10523=>"010001100",
  10524=>"001000100",
  10525=>"111110011",
  10526=>"100010110",
  10527=>"110110101",
  10528=>"100100011",
  10529=>"111000001",
  10530=>"000001101",
  10531=>"101010010",
  10532=>"101111010",
  10533=>"011011000",
  10534=>"010111100",
  10535=>"100010001",
  10536=>"100101001",
  10537=>"111111010",
  10538=>"110000000",
  10539=>"111101100",
  10540=>"101100010",
  10541=>"000000110",
  10542=>"111100111",
  10543=>"000110000",
  10544=>"000110100",
  10545=>"100111011",
  10546=>"010101010",
  10547=>"111100101",
  10548=>"011000011",
  10549=>"101000101",
  10550=>"110000110",
  10551=>"111101111",
  10552=>"110100111",
  10553=>"100011011",
  10554=>"001111001",
  10555=>"101010110",
  10556=>"010000010",
  10557=>"101110100",
  10558=>"010011011",
  10559=>"100010011",
  10560=>"011011010",
  10561=>"111111011",
  10562=>"100001110",
  10563=>"010000100",
  10564=>"001010010",
  10565=>"110110001",
  10566=>"101000100",
  10567=>"110100010",
  10568=>"011011000",
  10569=>"100000011",
  10570=>"001111010",
  10571=>"011000110",
  10572=>"000010110",
  10573=>"010010000",
  10574=>"100111110",
  10575=>"010010100",
  10576=>"001100110",
  10577=>"011011111",
  10578=>"010001010",
  10579=>"111001010",
  10580=>"111000111",
  10581=>"010110101",
  10582=>"111110100",
  10583=>"100000000",
  10584=>"011000101",
  10585=>"011100111",
  10586=>"100010011",
  10587=>"011111101",
  10588=>"011101000",
  10589=>"101101101",
  10590=>"000110111",
  10591=>"001011001",
  10592=>"011000110",
  10593=>"100111001",
  10594=>"000101010",
  10595=>"000000110",
  10596=>"100011010",
  10597=>"011101000",
  10598=>"000100010",
  10599=>"000001000",
  10600=>"010010001",
  10601=>"111000011",
  10602=>"111001011",
  10603=>"101010101",
  10604=>"000100100",
  10605=>"001001000",
  10606=>"011000111",
  10607=>"001010000",
  10608=>"110001011",
  10609=>"000001100",
  10610=>"011010011",
  10611=>"001010101",
  10612=>"100100111",
  10613=>"101110111",
  10614=>"111010101",
  10615=>"000111010",
  10616=>"001000101",
  10617=>"110100101",
  10618=>"100110110",
  10619=>"001110101",
  10620=>"111110111",
  10621=>"101100110",
  10622=>"111110100",
  10623=>"110110011",
  10624=>"111101101",
  10625=>"101000111",
  10626=>"000000111",
  10627=>"101011000",
  10628=>"111000010",
  10629=>"010011100",
  10630=>"111000011",
  10631=>"001011000",
  10632=>"110111011",
  10633=>"001001010",
  10634=>"000100101",
  10635=>"110000011",
  10636=>"000100100",
  10637=>"100100000",
  10638=>"011001111",
  10639=>"011101101",
  10640=>"001111110",
  10641=>"110101100",
  10642=>"111111010",
  10643=>"100100000",
  10644=>"010001101",
  10645=>"100001001",
  10646=>"100000010",
  10647=>"100011010",
  10648=>"010100001",
  10649=>"110000100",
  10650=>"010110101",
  10651=>"001000101",
  10652=>"000000011",
  10653=>"000000010",
  10654=>"000010001",
  10655=>"001000000",
  10656=>"110101101",
  10657=>"011011001",
  10658=>"000010011",
  10659=>"100011001",
  10660=>"000000000",
  10661=>"000001001",
  10662=>"001001101",
  10663=>"010110010",
  10664=>"001110010",
  10665=>"001100010",
  10666=>"101000000",
  10667=>"001010101",
  10668=>"011001011",
  10669=>"010101111",
  10670=>"110100110",
  10671=>"101101011",
  10672=>"001100000",
  10673=>"011111010",
  10674=>"110011100",
  10675=>"000010111",
  10676=>"001101101",
  10677=>"101001000",
  10678=>"000011101",
  10679=>"101001101",
  10680=>"011001111",
  10681=>"001000111",
  10682=>"000000000",
  10683=>"111011111",
  10684=>"111011101",
  10685=>"000011001",
  10686=>"110001001",
  10687=>"110101001",
  10688=>"101100000",
  10689=>"100100010",
  10690=>"111000000",
  10691=>"011011100",
  10692=>"100001000",
  10693=>"100110001",
  10694=>"111100101",
  10695=>"101100001",
  10696=>"011101111",
  10697=>"100111010",
  10698=>"111111101",
  10699=>"000001000",
  10700=>"101000011",
  10701=>"001101001",
  10702=>"010001011",
  10703=>"010011001",
  10704=>"001111010",
  10705=>"000100110",
  10706=>"111111000",
  10707=>"100101001",
  10708=>"110110111",
  10709=>"011100110",
  10710=>"010101101",
  10711=>"110001101",
  10712=>"010010000",
  10713=>"011000101",
  10714=>"110101111",
  10715=>"100011111",
  10716=>"111111111",
  10717=>"010001010",
  10718=>"101110101",
  10719=>"111110000",
  10720=>"001010010",
  10721=>"011010000",
  10722=>"000000011",
  10723=>"001001000",
  10724=>"001111000",
  10725=>"100010001",
  10726=>"101110001",
  10727=>"100010001",
  10728=>"111001011",
  10729=>"101100001",
  10730=>"001100001",
  10731=>"000100111",
  10732=>"101111111",
  10733=>"110110001",
  10734=>"100101000",
  10735=>"010100000",
  10736=>"011011000",
  10737=>"010011110",
  10738=>"111000010",
  10739=>"000101011",
  10740=>"111001000",
  10741=>"010010100",
  10742=>"010000111",
  10743=>"111010111",
  10744=>"101011001",
  10745=>"011100110",
  10746=>"111101011",
  10747=>"011001100",
  10748=>"111000011",
  10749=>"000100101",
  10750=>"110011100",
  10751=>"111111111",
  10752=>"001100111",
  10753=>"010100110",
  10754=>"110110001",
  10755=>"110101101",
  10756=>"001101110",
  10757=>"111101010",
  10758=>"110010111",
  10759=>"001001000",
  10760=>"000001001",
  10761=>"010110110",
  10762=>"011101001",
  10763=>"001001010",
  10764=>"001111001",
  10765=>"000100010",
  10766=>"010001101",
  10767=>"101111000",
  10768=>"000101001",
  10769=>"011011111",
  10770=>"110111000",
  10771=>"100101001",
  10772=>"101110010",
  10773=>"011100010",
  10774=>"100011010",
  10775=>"100101110",
  10776=>"000001100",
  10777=>"001001111",
  10778=>"110110110",
  10779=>"000111110",
  10780=>"100110111",
  10781=>"000010101",
  10782=>"110001110",
  10783=>"110101111",
  10784=>"110001000",
  10785=>"111111101",
  10786=>"101010010",
  10787=>"001111011",
  10788=>"100111001",
  10789=>"100010000",
  10790=>"110100110",
  10791=>"101100111",
  10792=>"110000110",
  10793=>"111010000",
  10794=>"010111101",
  10795=>"010001000",
  10796=>"110010111",
  10797=>"111000000",
  10798=>"110000111",
  10799=>"000110011",
  10800=>"011100100",
  10801=>"111111101",
  10802=>"111001000",
  10803=>"000001000",
  10804=>"111101111",
  10805=>"111001111",
  10806=>"011101000",
  10807=>"010010010",
  10808=>"110000000",
  10809=>"101011001",
  10810=>"000001111",
  10811=>"011110010",
  10812=>"000011000",
  10813=>"101111000",
  10814=>"010101000",
  10815=>"000000010",
  10816=>"000111011",
  10817=>"000001101",
  10818=>"111100110",
  10819=>"011001111",
  10820=>"110111100",
  10821=>"010000011",
  10822=>"011001011",
  10823=>"010100001",
  10824=>"110100010",
  10825=>"010011100",
  10826=>"111010110",
  10827=>"111111111",
  10828=>"000101101",
  10829=>"100101000",
  10830=>"111010100",
  10831=>"001010101",
  10832=>"011010010",
  10833=>"101011100",
  10834=>"011101100",
  10835=>"110010010",
  10836=>"111010111",
  10837=>"110101110",
  10838=>"000110001",
  10839=>"101100100",
  10840=>"110110110",
  10841=>"100100000",
  10842=>"100011111",
  10843=>"001001010",
  10844=>"101101010",
  10845=>"011010000",
  10846=>"001110011",
  10847=>"000011110",
  10848=>"110000110",
  10849=>"100100100",
  10850=>"101001111",
  10851=>"111101111",
  10852=>"011011101",
  10853=>"011010101",
  10854=>"101100001",
  10855=>"011100011",
  10856=>"101101111",
  10857=>"010111001",
  10858=>"110110110",
  10859=>"101010011",
  10860=>"101000111",
  10861=>"010010010",
  10862=>"101100100",
  10863=>"001100110",
  10864=>"111101011",
  10865=>"000111011",
  10866=>"101111010",
  10867=>"000001100",
  10868=>"101010100",
  10869=>"111000110",
  10870=>"001010010",
  10871=>"010000110",
  10872=>"000011010",
  10873=>"111011011",
  10874=>"100111110",
  10875=>"010011111",
  10876=>"111110011",
  10877=>"001110100",
  10878=>"110101000",
  10879=>"010100010",
  10880=>"110111110",
  10881=>"111001001",
  10882=>"010110110",
  10883=>"010001001",
  10884=>"101011101",
  10885=>"010001111",
  10886=>"100110000",
  10887=>"111101111",
  10888=>"100101110",
  10889=>"111000100",
  10890=>"110011001",
  10891=>"100100111",
  10892=>"000110101",
  10893=>"110101010",
  10894=>"010110000",
  10895=>"000011011",
  10896=>"101001001",
  10897=>"000010101",
  10898=>"101011011",
  10899=>"000011011",
  10900=>"101010101",
  10901=>"001110000",
  10902=>"010000101",
  10903=>"011100011",
  10904=>"110010000",
  10905=>"010100101",
  10906=>"111110111",
  10907=>"110110111",
  10908=>"010100000",
  10909=>"001111111",
  10910=>"000100011",
  10911=>"111100111",
  10912=>"010000000",
  10913=>"001100000",
  10914=>"110011101",
  10915=>"011001010",
  10916=>"101001001",
  10917=>"000110100",
  10918=>"111101011",
  10919=>"110100010",
  10920=>"100001101",
  10921=>"101011100",
  10922=>"101000110",
  10923=>"110010101",
  10924=>"000010001",
  10925=>"010010101",
  10926=>"110110110",
  10927=>"101111101",
  10928=>"001011010",
  10929=>"101000111",
  10930=>"100100110",
  10931=>"111110101",
  10932=>"000101011",
  10933=>"110101111",
  10934=>"110101101",
  10935=>"111110100",
  10936=>"111011101",
  10937=>"000110110",
  10938=>"110001011",
  10939=>"010000011",
  10940=>"100000100",
  10941=>"111010111",
  10942=>"111011000",
  10943=>"101100011",
  10944=>"011111000",
  10945=>"010110110",
  10946=>"001101000",
  10947=>"100110110",
  10948=>"000111010",
  10949=>"000111010",
  10950=>"000000111",
  10951=>"101111000",
  10952=>"111111010",
  10953=>"110010101",
  10954=>"101111010",
  10955=>"001100000",
  10956=>"011010010",
  10957=>"011101001",
  10958=>"111011010",
  10959=>"110100111",
  10960=>"101010101",
  10961=>"110001011",
  10962=>"111001110",
  10963=>"101100001",
  10964=>"000011000",
  10965=>"101000011",
  10966=>"001001110",
  10967=>"100001101",
  10968=>"100001111",
  10969=>"001000100",
  10970=>"100100000",
  10971=>"000101100",
  10972=>"000000010",
  10973=>"001101011",
  10974=>"000100111",
  10975=>"010000011",
  10976=>"110101101",
  10977=>"001111001",
  10978=>"101111111",
  10979=>"101011010",
  10980=>"100101001",
  10981=>"110000001",
  10982=>"111110010",
  10983=>"111110001",
  10984=>"111010101",
  10985=>"100100111",
  10986=>"110111111",
  10987=>"100100111",
  10988=>"100101101",
  10989=>"110001100",
  10990=>"111010101",
  10991=>"110110101",
  10992=>"001101111",
  10993=>"000110101",
  10994=>"110010000",
  10995=>"111101011",
  10996=>"100110010",
  10997=>"001000000",
  10998=>"110110000",
  10999=>"110111010",
  11000=>"110010100",
  11001=>"001011110",
  11002=>"010110111",
  11003=>"011000100",
  11004=>"000111101",
  11005=>"010000110",
  11006=>"011001110",
  11007=>"010000100",
  11008=>"010000100",
  11009=>"110001110",
  11010=>"111111001",
  11011=>"000011000",
  11012=>"011110111",
  11013=>"110111000",
  11014=>"011010001",
  11015=>"001011001",
  11016=>"000111001",
  11017=>"001111111",
  11018=>"100011011",
  11019=>"011100111",
  11020=>"100000001",
  11021=>"001101010",
  11022=>"110000110",
  11023=>"011101001",
  11024=>"111100001",
  11025=>"000100000",
  11026=>"000101001",
  11027=>"100001010",
  11028=>"100111100",
  11029=>"110100110",
  11030=>"001010000",
  11031=>"110111000",
  11032=>"101110110",
  11033=>"110010110",
  11034=>"101010011",
  11035=>"110110101",
  11036=>"011101101",
  11037=>"001011100",
  11038=>"001010010",
  11039=>"001000110",
  11040=>"111011101",
  11041=>"101101101",
  11042=>"111000111",
  11043=>"111000000",
  11044=>"010000100",
  11045=>"000000100",
  11046=>"111010010",
  11047=>"001010110",
  11048=>"111101011",
  11049=>"110100101",
  11050=>"101110111",
  11051=>"001100111",
  11052=>"100101100",
  11053=>"000010001",
  11054=>"001000001",
  11055=>"011111010",
  11056=>"110110001",
  11057=>"111011101",
  11058=>"001100110",
  11059=>"011000000",
  11060=>"000001010",
  11061=>"011101010",
  11062=>"111100011",
  11063=>"111100000",
  11064=>"100000010",
  11065=>"000011010",
  11066=>"110010000",
  11067=>"000001110",
  11068=>"100000000",
  11069=>"111010001",
  11070=>"110111001",
  11071=>"011001111",
  11072=>"000000101",
  11073=>"000111101",
  11074=>"001011101",
  11075=>"001000110",
  11076=>"100101000",
  11077=>"101011010",
  11078=>"111101010",
  11079=>"101100001",
  11080=>"000100010",
  11081=>"110111100",
  11082=>"011000011",
  11083=>"001000010",
  11084=>"111111100",
  11085=>"100111111",
  11086=>"011101100",
  11087=>"111111110",
  11088=>"000001000",
  11089=>"100010101",
  11090=>"101111110",
  11091=>"110000001",
  11092=>"000110111",
  11093=>"101000011",
  11094=>"001100101",
  11095=>"001001000",
  11096=>"101010000",
  11097=>"000011101",
  11098=>"100110011",
  11099=>"001101111",
  11100=>"010111001",
  11101=>"111111111",
  11102=>"000101100",
  11103=>"110001101",
  11104=>"101111100",
  11105=>"101000101",
  11106=>"101010001",
  11107=>"001100111",
  11108=>"111000110",
  11109=>"011101011",
  11110=>"010010011",
  11111=>"011100101",
  11112=>"110000001",
  11113=>"110011010",
  11114=>"100001001",
  11115=>"111111000",
  11116=>"110001011",
  11117=>"001101110",
  11118=>"010010001",
  11119=>"000000111",
  11120=>"110001001",
  11121=>"111010111",
  11122=>"001001010",
  11123=>"101011110",
  11124=>"010010011",
  11125=>"101001000",
  11126=>"111011010",
  11127=>"101011111",
  11128=>"101001110",
  11129=>"111110001",
  11130=>"101110111",
  11131=>"100111100",
  11132=>"000011000",
  11133=>"111111111",
  11134=>"101000111",
  11135=>"011001011",
  11136=>"110000011",
  11137=>"000111100",
  11138=>"111111101",
  11139=>"111010111",
  11140=>"110100000",
  11141=>"011010000",
  11142=>"101110011",
  11143=>"000000101",
  11144=>"011101100",
  11145=>"001000111",
  11146=>"001100011",
  11147=>"111110111",
  11148=>"000000010",
  11149=>"110010011",
  11150=>"101101010",
  11151=>"011100010",
  11152=>"110101011",
  11153=>"100000110",
  11154=>"111111001",
  11155=>"111111011",
  11156=>"100001011",
  11157=>"011111011",
  11158=>"000011010",
  11159=>"010000110",
  11160=>"010000010",
  11161=>"000110110",
  11162=>"000100011",
  11163=>"001000001",
  11164=>"111110111",
  11165=>"101010110",
  11166=>"100100000",
  11167=>"101100011",
  11168=>"010101100",
  11169=>"001100010",
  11170=>"000011100",
  11171=>"011010010",
  11172=>"011010000",
  11173=>"010001001",
  11174=>"000011111",
  11175=>"001000110",
  11176=>"101010100",
  11177=>"000010010",
  11178=>"000100011",
  11179=>"011001010",
  11180=>"111011010",
  11181=>"001100111",
  11182=>"001010101",
  11183=>"101000100",
  11184=>"101111001",
  11185=>"000111110",
  11186=>"011000100",
  11187=>"000011000",
  11188=>"101100001",
  11189=>"011100101",
  11190=>"101100110",
  11191=>"101101100",
  11192=>"110010100",
  11193=>"000111010",
  11194=>"101011110",
  11195=>"100100101",
  11196=>"101001101",
  11197=>"000001101",
  11198=>"101110010",
  11199=>"001010101",
  11200=>"101111111",
  11201=>"110000101",
  11202=>"110011000",
  11203=>"000011100",
  11204=>"010101110",
  11205=>"010011011",
  11206=>"110000000",
  11207=>"101100100",
  11208=>"101000000",
  11209=>"111000111",
  11210=>"110000110",
  11211=>"011011010",
  11212=>"110010111",
  11213=>"010111100",
  11214=>"010111000",
  11215=>"000011001",
  11216=>"110001011",
  11217=>"011011001",
  11218=>"001111111",
  11219=>"101011011",
  11220=>"000001010",
  11221=>"001111000",
  11222=>"001110101",
  11223=>"111001010",
  11224=>"100001010",
  11225=>"101011111",
  11226=>"000011100",
  11227=>"101010000",
  11228=>"111010101",
  11229=>"001001001",
  11230=>"001000000",
  11231=>"010001000",
  11232=>"110011110",
  11233=>"111100000",
  11234=>"011001110",
  11235=>"100110011",
  11236=>"011011001",
  11237=>"011001001",
  11238=>"000011011",
  11239=>"111111000",
  11240=>"001001001",
  11241=>"100100000",
  11242=>"011111001",
  11243=>"101010011",
  11244=>"111110100",
  11245=>"011111110",
  11246=>"010010000",
  11247=>"000010011",
  11248=>"000111111",
  11249=>"000110001",
  11250=>"101011001",
  11251=>"100011111",
  11252=>"100111111",
  11253=>"101110100",
  11254=>"000001011",
  11255=>"100111111",
  11256=>"001110111",
  11257=>"111000100",
  11258=>"111101011",
  11259=>"100100000",
  11260=>"010110000",
  11261=>"111111000",
  11262=>"111000111",
  11263=>"011100000",
  11264=>"000010101",
  11265=>"110100111",
  11266=>"100011010",
  11267=>"110111100",
  11268=>"001111110",
  11269=>"101110001",
  11270=>"100110011",
  11271=>"000100100",
  11272=>"101110110",
  11273=>"110010110",
  11274=>"011100001",
  11275=>"000110010",
  11276=>"111101110",
  11277=>"001001011",
  11278=>"110010000",
  11279=>"111100010",
  11280=>"010101011",
  11281=>"001011010",
  11282=>"010000000",
  11283=>"110101111",
  11284=>"100100000",
  11285=>"111111101",
  11286=>"111001001",
  11287=>"001011100",
  11288=>"010001011",
  11289=>"011101010",
  11290=>"000100111",
  11291=>"000100010",
  11292=>"000101110",
  11293=>"001001001",
  11294=>"010001110",
  11295=>"011000110",
  11296=>"010000010",
  11297=>"110101010",
  11298=>"101111100",
  11299=>"111101111",
  11300=>"010000000",
  11301=>"000001011",
  11302=>"001011010",
  11303=>"111110100",
  11304=>"010111101",
  11305=>"101110010",
  11306=>"001001111",
  11307=>"011010100",
  11308=>"001000001",
  11309=>"011011011",
  11310=>"101110000",
  11311=>"111001011",
  11312=>"100001001",
  11313=>"000000111",
  11314=>"000100001",
  11315=>"101111111",
  11316=>"110010111",
  11317=>"111111100",
  11318=>"000100010",
  11319=>"111011010",
  11320=>"110110010",
  11321=>"011010111",
  11322=>"000100001",
  11323=>"111011001",
  11324=>"100001001",
  11325=>"010101010",
  11326=>"001100000",
  11327=>"110100111",
  11328=>"101111011",
  11329=>"000011000",
  11330=>"100101110",
  11331=>"010110101",
  11332=>"000011111",
  11333=>"000101001",
  11334=>"001010100",
  11335=>"101100011",
  11336=>"011101000",
  11337=>"111010111",
  11338=>"010010111",
  11339=>"000111111",
  11340=>"001100010",
  11341=>"110011001",
  11342=>"000101000",
  11343=>"011000010",
  11344=>"100111111",
  11345=>"000000001",
  11346=>"000110010",
  11347=>"000010010",
  11348=>"000100101",
  11349=>"010011000",
  11350=>"010100100",
  11351=>"000010000",
  11352=>"000110010",
  11353=>"101110100",
  11354=>"111010100",
  11355=>"111000101",
  11356=>"011001111",
  11357=>"000000100",
  11358=>"001010100",
  11359=>"010010100",
  11360=>"101000010",
  11361=>"000010110",
  11362=>"111010110",
  11363=>"000000001",
  11364=>"010101111",
  11365=>"000000111",
  11366=>"010010100",
  11367=>"001010000",
  11368=>"110111001",
  11369=>"001000111",
  11370=>"000001111",
  11371=>"010100100",
  11372=>"001000101",
  11373=>"011010010",
  11374=>"111001111",
  11375=>"111100101",
  11376=>"101001000",
  11377=>"111000110",
  11378=>"010001011",
  11379=>"010100100",
  11380=>"111010111",
  11381=>"011000011",
  11382=>"010101001",
  11383=>"000110111",
  11384=>"001000111",
  11385=>"000000100",
  11386=>"001001001",
  11387=>"100011110",
  11388=>"001001010",
  11389=>"110000100",
  11390=>"011000101",
  11391=>"000000001",
  11392=>"011000000",
  11393=>"001010010",
  11394=>"001111101",
  11395=>"010010110",
  11396=>"101010000",
  11397=>"010101111",
  11398=>"010100001",
  11399=>"111111101",
  11400=>"100110000",
  11401=>"111111111",
  11402=>"101001001",
  11403=>"011100101",
  11404=>"110000001",
  11405=>"111001001",
  11406=>"000001001",
  11407=>"100001001",
  11408=>"000011101",
  11409=>"010000001",
  11410=>"111111010",
  11411=>"100111111",
  11412=>"111111101",
  11413=>"000100110",
  11414=>"111100000",
  11415=>"010101011",
  11416=>"111010111",
  11417=>"011000000",
  11418=>"010110101",
  11419=>"001100010",
  11420=>"000101100",
  11421=>"111000100",
  11422=>"111000101",
  11423=>"000101000",
  11424=>"001110000",
  11425=>"000110111",
  11426=>"111011110",
  11427=>"101101101",
  11428=>"010011101",
  11429=>"100001011",
  11430=>"111000011",
  11431=>"111110111",
  11432=>"001000101",
  11433=>"000001011",
  11434=>"011111110",
  11435=>"100011111",
  11436=>"001100011",
  11437=>"011001100",
  11438=>"010101001",
  11439=>"101011010",
  11440=>"111111010",
  11441=>"110001011",
  11442=>"100111000",
  11443=>"101010100",
  11444=>"110110110",
  11445=>"101111011",
  11446=>"110110010",
  11447=>"001000100",
  11448=>"111011001",
  11449=>"000101111",
  11450=>"010101110",
  11451=>"000100110",
  11452=>"011001001",
  11453=>"001110010",
  11454=>"001010101",
  11455=>"000010111",
  11456=>"100101000",
  11457=>"111100111",
  11458=>"011111111",
  11459=>"000011110",
  11460=>"110000010",
  11461=>"011110101",
  11462=>"010110100",
  11463=>"001100110",
  11464=>"010001110",
  11465=>"011100110",
  11466=>"010001010",
  11467=>"111010011",
  11468=>"110010110",
  11469=>"000011110",
  11470=>"111111010",
  11471=>"111111001",
  11472=>"111101111",
  11473=>"000010111",
  11474=>"010010010",
  11475=>"000110010",
  11476=>"011000100",
  11477=>"101000000",
  11478=>"011111111",
  11479=>"100110110",
  11480=>"101111001",
  11481=>"110000111",
  11482=>"111100101",
  11483=>"010101101",
  11484=>"111111111",
  11485=>"110101111",
  11486=>"110001100",
  11487=>"000111100",
  11488=>"111111011",
  11489=>"011010011",
  11490=>"111111110",
  11491=>"001111111",
  11492=>"000000100",
  11493=>"000001101",
  11494=>"101010011",
  11495=>"100001111",
  11496=>"110011110",
  11497=>"110111000",
  11498=>"001110101",
  11499=>"110111100",
  11500=>"110111001",
  11501=>"101000001",
  11502=>"010111101",
  11503=>"000111110",
  11504=>"101000001",
  11505=>"011011011",
  11506=>"110110000",
  11507=>"100000000",
  11508=>"011101100",
  11509=>"001010010",
  11510=>"011110100",
  11511=>"011101111",
  11512=>"010011011",
  11513=>"110100101",
  11514=>"100101111",
  11515=>"011011000",
  11516=>"001101101",
  11517=>"011101010",
  11518=>"100101110",
  11519=>"000001010",
  11520=>"010111010",
  11521=>"011010100",
  11522=>"101101001",
  11523=>"011010100",
  11524=>"011011000",
  11525=>"011101101",
  11526=>"110011100",
  11527=>"110111000",
  11528=>"010000011",
  11529=>"011010011",
  11530=>"111010000",
  11531=>"111110000",
  11532=>"000100010",
  11533=>"111110010",
  11534=>"100011110",
  11535=>"000001010",
  11536=>"100110001",
  11537=>"111110111",
  11538=>"111011100",
  11539=>"110000010",
  11540=>"001011001",
  11541=>"000110000",
  11542=>"111110011",
  11543=>"110100100",
  11544=>"101000100",
  11545=>"110101001",
  11546=>"001111011",
  11547=>"111100111",
  11548=>"101100000",
  11549=>"010000000",
  11550=>"010101101",
  11551=>"101010110",
  11552=>"001011100",
  11553=>"111111100",
  11554=>"000010100",
  11555=>"111011001",
  11556=>"011000111",
  11557=>"010100100",
  11558=>"100000010",
  11559=>"010110111",
  11560=>"110110000",
  11561=>"010111101",
  11562=>"100100011",
  11563=>"001000100",
  11564=>"101111001",
  11565=>"000011010",
  11566=>"101111011",
  11567=>"001100011",
  11568=>"100100000",
  11569=>"100110011",
  11570=>"001111111",
  11571=>"001100011",
  11572=>"000000010",
  11573=>"001100000",
  11574=>"000001101",
  11575=>"101101111",
  11576=>"110000010",
  11577=>"010100000",
  11578=>"111011000",
  11579=>"111111011",
  11580=>"011101011",
  11581=>"001001110",
  11582=>"111111100",
  11583=>"111111111",
  11584=>"011101100",
  11585=>"011111000",
  11586=>"010111111",
  11587=>"000000000",
  11588=>"000100011",
  11589=>"100010111",
  11590=>"101111100",
  11591=>"101011110",
  11592=>"110110100",
  11593=>"111100000",
  11594=>"110011100",
  11595=>"110100110",
  11596=>"010010001",
  11597=>"001001101",
  11598=>"011100001",
  11599=>"011101100",
  11600=>"100000010",
  11601=>"100000001",
  11602=>"001011001",
  11603=>"001000011",
  11604=>"000111100",
  11605=>"000101111",
  11606=>"110010010",
  11607=>"110010110",
  11608=>"011010110",
  11609=>"110101100",
  11610=>"100011100",
  11611=>"110010101",
  11612=>"011110100",
  11613=>"111110101",
  11614=>"110111011",
  11615=>"011011100",
  11616=>"001111110",
  11617=>"111101100",
  11618=>"101000101",
  11619=>"000001111",
  11620=>"111101011",
  11621=>"000111010",
  11622=>"011000100",
  11623=>"100001100",
  11624=>"011010110",
  11625=>"000010100",
  11626=>"011100010",
  11627=>"011001100",
  11628=>"011110100",
  11629=>"100010011",
  11630=>"011110000",
  11631=>"101111101",
  11632=>"101001110",
  11633=>"011010101",
  11634=>"011001001",
  11635=>"011110000",
  11636=>"110101101",
  11637=>"001000111",
  11638=>"000000001",
  11639=>"110001000",
  11640=>"010011010",
  11641=>"111100001",
  11642=>"111000111",
  11643=>"001111010",
  11644=>"100111100",
  11645=>"110011000",
  11646=>"010000110",
  11647=>"011101000",
  11648=>"111011000",
  11649=>"001111101",
  11650=>"111101111",
  11651=>"000001101",
  11652=>"000101011",
  11653=>"101111111",
  11654=>"101111111",
  11655=>"110011001",
  11656=>"111001101",
  11657=>"010011001",
  11658=>"001011010",
  11659=>"111110011",
  11660=>"000001111",
  11661=>"110110000",
  11662=>"100011110",
  11663=>"010100100",
  11664=>"101010100",
  11665=>"110011000",
  11666=>"100001100",
  11667=>"100100110",
  11668=>"001010110",
  11669=>"001100110",
  11670=>"000101000",
  11671=>"110010100",
  11672=>"010001011",
  11673=>"010111101",
  11674=>"111111111",
  11675=>"001111011",
  11676=>"011010001",
  11677=>"101101110",
  11678=>"010001110",
  11679=>"010000010",
  11680=>"111110000",
  11681=>"111011101",
  11682=>"000110011",
  11683=>"100100100",
  11684=>"110110111",
  11685=>"001111000",
  11686=>"110101100",
  11687=>"011011111",
  11688=>"100111010",
  11689=>"110101010",
  11690=>"000110010",
  11691=>"111001111",
  11692=>"000011010",
  11693=>"010101010",
  11694=>"110111011",
  11695=>"100010010",
  11696=>"001101011",
  11697=>"101010000",
  11698=>"000001011",
  11699=>"000011010",
  11700=>"110110011",
  11701=>"100110001",
  11702=>"110110010",
  11703=>"001010111",
  11704=>"101111111",
  11705=>"011110011",
  11706=>"111011001",
  11707=>"110100000",
  11708=>"011101001",
  11709=>"100011001",
  11710=>"000111000",
  11711=>"110110100",
  11712=>"011101011",
  11713=>"111111011",
  11714=>"110001000",
  11715=>"110001110",
  11716=>"001100101",
  11717=>"000001000",
  11718=>"110000100",
  11719=>"100110111",
  11720=>"000001011",
  11721=>"101100000",
  11722=>"111111110",
  11723=>"111100000",
  11724=>"101110010",
  11725=>"011001011",
  11726=>"100101001",
  11727=>"110100111",
  11728=>"011000111",
  11729=>"011011001",
  11730=>"010011000",
  11731=>"100100110",
  11732=>"001000110",
  11733=>"110001000",
  11734=>"000101111",
  11735=>"000110110",
  11736=>"011001001",
  11737=>"010010000",
  11738=>"110101010",
  11739=>"111110111",
  11740=>"001100100",
  11741=>"010011011",
  11742=>"101010110",
  11743=>"100001000",
  11744=>"001000110",
  11745=>"110110000",
  11746=>"101001010",
  11747=>"100111110",
  11748=>"101011001",
  11749=>"010010110",
  11750=>"101001101",
  11751=>"011100111",
  11752=>"010111011",
  11753=>"011111101",
  11754=>"010101110",
  11755=>"111110010",
  11756=>"010100010",
  11757=>"100101101",
  11758=>"110110111",
  11759=>"011001101",
  11760=>"101100100",
  11761=>"100010111",
  11762=>"111111101",
  11763=>"011010000",
  11764=>"111101111",
  11765=>"000010111",
  11766=>"110000101",
  11767=>"100011111",
  11768=>"000110110",
  11769=>"101111111",
  11770=>"110111010",
  11771=>"101101100",
  11772=>"011000110",
  11773=>"110011101",
  11774=>"100000111",
  11775=>"110010100",
  11776=>"010000011",
  11777=>"000110100",
  11778=>"111111010",
  11779=>"010010001",
  11780=>"100110111",
  11781=>"001101010",
  11782=>"110000000",
  11783=>"010111000",
  11784=>"100000101",
  11785=>"111101001",
  11786=>"011010110",
  11787=>"001010001",
  11788=>"101010001",
  11789=>"100011011",
  11790=>"101111011",
  11791=>"100100111",
  11792=>"100100100",
  11793=>"101110011",
  11794=>"011001000",
  11795=>"111010010",
  11796=>"111001001",
  11797=>"000110111",
  11798=>"101111111",
  11799=>"000100011",
  11800=>"010100001",
  11801=>"111001011",
  11802=>"100111000",
  11803=>"101000101",
  11804=>"101110011",
  11805=>"011110010",
  11806=>"101110011",
  11807=>"001100101",
  11808=>"111111111",
  11809=>"110011101",
  11810=>"010011000",
  11811=>"010000001",
  11812=>"111010111",
  11813=>"010111110",
  11814=>"101110101",
  11815=>"100100101",
  11816=>"000110100",
  11817=>"101101000",
  11818=>"100101101",
  11819=>"010111010",
  11820=>"111101100",
  11821=>"100000100",
  11822=>"000010110",
  11823=>"001010011",
  11824=>"111100010",
  11825=>"001111110",
  11826=>"101111100",
  11827=>"100000001",
  11828=>"000110110",
  11829=>"010011100",
  11830=>"001010101",
  11831=>"101001000",
  11832=>"111111010",
  11833=>"111010110",
  11834=>"000100001",
  11835=>"011111010",
  11836=>"110001111",
  11837=>"011011010",
  11838=>"001101111",
  11839=>"010010011",
  11840=>"000110010",
  11841=>"011001111",
  11842=>"010010001",
  11843=>"000010011",
  11844=>"010010101",
  11845=>"111010101",
  11846=>"001000010",
  11847=>"111101010",
  11848=>"100110001",
  11849=>"100101000",
  11850=>"110010110",
  11851=>"111110000",
  11852=>"011110001",
  11853=>"001001100",
  11854=>"101111000",
  11855=>"101100010",
  11856=>"111010010",
  11857=>"111111100",
  11858=>"001001101",
  11859=>"001110000",
  11860=>"100011110",
  11861=>"111110010",
  11862=>"110101100",
  11863=>"001011011",
  11864=>"011110010",
  11865=>"000101000",
  11866=>"111001111",
  11867=>"101100010",
  11868=>"001001000",
  11869=>"000110100",
  11870=>"101001110",
  11871=>"100110101",
  11872=>"011000100",
  11873=>"110000001",
  11874=>"001010011",
  11875=>"100010011",
  11876=>"000100000",
  11877=>"001000011",
  11878=>"011011010",
  11879=>"000011001",
  11880=>"000010101",
  11881=>"110110011",
  11882=>"001111100",
  11883=>"000010010",
  11884=>"000001100",
  11885=>"010110001",
  11886=>"010010110",
  11887=>"011110011",
  11888=>"111111010",
  11889=>"101110111",
  11890=>"011011100",
  11891=>"000101010",
  11892=>"100010000",
  11893=>"011011000",
  11894=>"111000010",
  11895=>"100100100",
  11896=>"000011001",
  11897=>"001111101",
  11898=>"101001001",
  11899=>"100101111",
  11900=>"111101001",
  11901=>"011111011",
  11902=>"000001001",
  11903=>"100011100",
  11904=>"111010110",
  11905=>"111100000",
  11906=>"000001110",
  11907=>"101101001",
  11908=>"111111101",
  11909=>"100011100",
  11910=>"001011010",
  11911=>"101010011",
  11912=>"101100100",
  11913=>"010111100",
  11914=>"010010110",
  11915=>"001000011",
  11916=>"011000010",
  11917=>"101010011",
  11918=>"011000000",
  11919=>"000111000",
  11920=>"000000100",
  11921=>"001000101",
  11922=>"001011000",
  11923=>"001000110",
  11924=>"010010010",
  11925=>"011110011",
  11926=>"000111111",
  11927=>"110111100",
  11928=>"100010111",
  11929=>"001111000",
  11930=>"110001011",
  11931=>"010111000",
  11932=>"000000111",
  11933=>"111001111",
  11934=>"111001111",
  11935=>"011000001",
  11936=>"110010000",
  11937=>"111101111",
  11938=>"000100011",
  11939=>"100010100",
  11940=>"100010010",
  11941=>"101011110",
  11942=>"011000111",
  11943=>"101101111",
  11944=>"000001000",
  11945=>"111011000",
  11946=>"001000100",
  11947=>"111110000",
  11948=>"101000001",
  11949=>"010010011",
  11950=>"011011100",
  11951=>"001111100",
  11952=>"011000010",
  11953=>"010101000",
  11954=>"101001001",
  11955=>"011011101",
  11956=>"001000000",
  11957=>"010100011",
  11958=>"111111101",
  11959=>"111101000",
  11960=>"011110100",
  11961=>"100000010",
  11962=>"010110110",
  11963=>"111101110",
  11964=>"011100000",
  11965=>"010111011",
  11966=>"000111111",
  11967=>"001111111",
  11968=>"110001001",
  11969=>"000111010",
  11970=>"111111101",
  11971=>"011101001",
  11972=>"001100001",
  11973=>"101101100",
  11974=>"011110110",
  11975=>"110011011",
  11976=>"110101000",
  11977=>"110000001",
  11978=>"000111011",
  11979=>"101110101",
  11980=>"001111111",
  11981=>"111100111",
  11982=>"100010000",
  11983=>"011001010",
  11984=>"000000010",
  11985=>"110100110",
  11986=>"010001101",
  11987=>"100011000",
  11988=>"010101011",
  11989=>"001100011",
  11990=>"101000100",
  11991=>"111010010",
  11992=>"011000101",
  11993=>"000100110",
  11994=>"111111011",
  11995=>"000100001",
  11996=>"100011010",
  11997=>"101100111",
  11998=>"011001111",
  11999=>"100010100",
  12000=>"101110110",
  12001=>"100110110",
  12002=>"000000010",
  12003=>"000101110",
  12004=>"100000011",
  12005=>"100010000",
  12006=>"111011111",
  12007=>"000101001",
  12008=>"100101101",
  12009=>"001100101",
  12010=>"000011110",
  12011=>"100011101",
  12012=>"100011101",
  12013=>"010011101",
  12014=>"101101100",
  12015=>"100011110",
  12016=>"010010010",
  12017=>"001110010",
  12018=>"111011100",
  12019=>"110001100",
  12020=>"011010010",
  12021=>"011010110",
  12022=>"100010010",
  12023=>"101000010",
  12024=>"011111100",
  12025=>"100001100",
  12026=>"110000011",
  12027=>"110100000",
  12028=>"010111111",
  12029=>"101001010",
  12030=>"111011100",
  12031=>"100111001",
  12032=>"100101100",
  12033=>"011011110",
  12034=>"010100101",
  12035=>"110100100",
  12036=>"111111110",
  12037=>"010001000",
  12038=>"011010111",
  12039=>"100001011",
  12040=>"010010011",
  12041=>"011001111",
  12042=>"000101111",
  12043=>"010010100",
  12044=>"011101110",
  12045=>"011111001",
  12046=>"100010110",
  12047=>"111001101",
  12048=>"110101010",
  12049=>"001011111",
  12050=>"110010110",
  12051=>"011000100",
  12052=>"100010110",
  12053=>"110001111",
  12054=>"001110011",
  12055=>"101000101",
  12056=>"101111010",
  12057=>"011110001",
  12058=>"110100010",
  12059=>"100000000",
  12060=>"010011011",
  12061=>"000101111",
  12062=>"100100010",
  12063=>"111011000",
  12064=>"000111011",
  12065=>"011111100",
  12066=>"011100100",
  12067=>"010011011",
  12068=>"110000111",
  12069=>"000111000",
  12070=>"100100000",
  12071=>"000000100",
  12072=>"001110001",
  12073=>"111000101",
  12074=>"001100101",
  12075=>"101101001",
  12076=>"101100101",
  12077=>"100111111",
  12078=>"100110000",
  12079=>"010111101",
  12080=>"010100001",
  12081=>"111010001",
  12082=>"100010111",
  12083=>"001011100",
  12084=>"000001000",
  12085=>"011100000",
  12086=>"000011000",
  12087=>"100111011",
  12088=>"010100101",
  12089=>"100011000",
  12090=>"101101000",
  12091=>"000000100",
  12092=>"110001100",
  12093=>"001100100",
  12094=>"010010100",
  12095=>"111110101",
  12096=>"110101100",
  12097=>"000111111",
  12098=>"010101001",
  12099=>"101111110",
  12100=>"100101011",
  12101=>"010101001",
  12102=>"111110001",
  12103=>"000011011",
  12104=>"011111111",
  12105=>"110011000",
  12106=>"000100010",
  12107=>"001000011",
  12108=>"100101100",
  12109=>"001110010",
  12110=>"111101001",
  12111=>"000100010",
  12112=>"011100001",
  12113=>"100100000",
  12114=>"101011100",
  12115=>"110001010",
  12116=>"010001100",
  12117=>"110001100",
  12118=>"101100010",
  12119=>"110001100",
  12120=>"010011111",
  12121=>"010010001",
  12122=>"111011011",
  12123=>"000000111",
  12124=>"001100111",
  12125=>"110000001",
  12126=>"100111110",
  12127=>"011110110",
  12128=>"001010101",
  12129=>"101010111",
  12130=>"101111010",
  12131=>"000000000",
  12132=>"110000110",
  12133=>"110000110",
  12134=>"011101111",
  12135=>"111100011",
  12136=>"100011000",
  12137=>"100111000",
  12138=>"111010101",
  12139=>"010101000",
  12140=>"101010000",
  12141=>"011001100",
  12142=>"111011111",
  12143=>"010111111",
  12144=>"100000010",
  12145=>"110101111",
  12146=>"000010011",
  12147=>"000101000",
  12148=>"000101100",
  12149=>"111011101",
  12150=>"111110110",
  12151=>"011111111",
  12152=>"101100011",
  12153=>"101000100",
  12154=>"001011001",
  12155=>"111001001",
  12156=>"100000001",
  12157=>"001100001",
  12158=>"110000111",
  12159=>"011110000",
  12160=>"001011100",
  12161=>"011000001",
  12162=>"000101000",
  12163=>"100111010",
  12164=>"111111010",
  12165=>"101101000",
  12166=>"110010101",
  12167=>"011100000",
  12168=>"000000001",
  12169=>"101100000",
  12170=>"000000001",
  12171=>"111010100",
  12172=>"100101110",
  12173=>"011001111",
  12174=>"010110110",
  12175=>"100001101",
  12176=>"110101011",
  12177=>"000000000",
  12178=>"110100001",
  12179=>"101010011",
  12180=>"100100000",
  12181=>"110100101",
  12182=>"000000110",
  12183=>"111001011",
  12184=>"110111100",
  12185=>"000101000",
  12186=>"101111011",
  12187=>"011000110",
  12188=>"010101001",
  12189=>"110000110",
  12190=>"011111111",
  12191=>"001001111",
  12192=>"000001101",
  12193=>"111101101",
  12194=>"011110100",
  12195=>"110100101",
  12196=>"011110001",
  12197=>"011111011",
  12198=>"000101111",
  12199=>"010101011",
  12200=>"111101011",
  12201=>"101000000",
  12202=>"101001001",
  12203=>"111000000",
  12204=>"110110001",
  12205=>"100110101",
  12206=>"000000101",
  12207=>"000000110",
  12208=>"000001001",
  12209=>"111100111",
  12210=>"001100000",
  12211=>"010001101",
  12212=>"011100101",
  12213=>"000001100",
  12214=>"000010010",
  12215=>"111110011",
  12216=>"111001100",
  12217=>"000101110",
  12218=>"110011111",
  12219=>"111000010",
  12220=>"110101011",
  12221=>"100000000",
  12222=>"111111011",
  12223=>"011111010",
  12224=>"100001101",
  12225=>"110000101",
  12226=>"001110110",
  12227=>"000010100",
  12228=>"001101101",
  12229=>"010101000",
  12230=>"110010000",
  12231=>"111001011",
  12232=>"110010000",
  12233=>"110010011",
  12234=>"100110000",
  12235=>"100110000",
  12236=>"001101110",
  12237=>"000110010",
  12238=>"010111011",
  12239=>"011100111",
  12240=>"110011011",
  12241=>"111101100",
  12242=>"001111101",
  12243=>"100111010",
  12244=>"111100001",
  12245=>"111100111",
  12246=>"000001010",
  12247=>"100100111",
  12248=>"000001011",
  12249=>"011000111",
  12250=>"011001001",
  12251=>"111101101",
  12252=>"111111000",
  12253=>"111010111",
  12254=>"001011110",
  12255=>"101100010",
  12256=>"000011110",
  12257=>"000111110",
  12258=>"111100111",
  12259=>"101000011",
  12260=>"001111000",
  12261=>"100011010",
  12262=>"100001000",
  12263=>"010010111",
  12264=>"011110001",
  12265=>"101110100",
  12266=>"101010010",
  12267=>"011101110",
  12268=>"101101011",
  12269=>"010101110",
  12270=>"011011011",
  12271=>"010111001",
  12272=>"110100000",
  12273=>"011110100",
  12274=>"111110001",
  12275=>"110001100",
  12276=>"100010010",
  12277=>"011100011",
  12278=>"100011000",
  12279=>"111111011",
  12280=>"111100000",
  12281=>"000010000",
  12282=>"000010101",
  12283=>"111000010",
  12284=>"101000000",
  12285=>"110011000",
  12286=>"110001111",
  12287=>"011101100",
  12288=>"111110110",
  12289=>"110001010",
  12290=>"110110111",
  12291=>"100110111",
  12292=>"111100101",
  12293=>"100001001",
  12294=>"110010110",
  12295=>"100111110",
  12296=>"011110001",
  12297=>"111000110",
  12298=>"011101101",
  12299=>"011110000",
  12300=>"100101100",
  12301=>"010001010",
  12302=>"010101001",
  12303=>"101101001",
  12304=>"111111000",
  12305=>"100101000",
  12306=>"010111101",
  12307=>"011101101",
  12308=>"000011111",
  12309=>"110111010",
  12310=>"101101110",
  12311=>"000100010",
  12312=>"000000010",
  12313=>"111011011",
  12314=>"111101001",
  12315=>"110111111",
  12316=>"001000100",
  12317=>"010100000",
  12318=>"001110110",
  12319=>"110010110",
  12320=>"010110111",
  12321=>"001111001",
  12322=>"100011010",
  12323=>"000111100",
  12324=>"000111100",
  12325=>"000100111",
  12326=>"111010000",
  12327=>"001000001",
  12328=>"101100000",
  12329=>"000011111",
  12330=>"100000101",
  12331=>"110000101",
  12332=>"000100100",
  12333=>"100000001",
  12334=>"100011010",
  12335=>"111110111",
  12336=>"010001100",
  12337=>"011101110",
  12338=>"100001111",
  12339=>"111011100",
  12340=>"101001101",
  12341=>"101010010",
  12342=>"010010001",
  12343=>"100010101",
  12344=>"101011010",
  12345=>"000110001",
  12346=>"001001101",
  12347=>"100000110",
  12348=>"000111110",
  12349=>"010100111",
  12350=>"001001010",
  12351=>"000110111",
  12352=>"000000100",
  12353=>"010000000",
  12354=>"110011000",
  12355=>"101011101",
  12356=>"100001110",
  12357=>"011101110",
  12358=>"111000010",
  12359=>"100100111",
  12360=>"100100101",
  12361=>"001111000",
  12362=>"101010011",
  12363=>"101001100",
  12364=>"111101001",
  12365=>"111011111",
  12366=>"000101000",
  12367=>"111110001",
  12368=>"001101000",
  12369=>"000101001",
  12370=>"010010011",
  12371=>"110111000",
  12372=>"111110111",
  12373=>"111011000",
  12374=>"110000010",
  12375=>"100000111",
  12376=>"111100100",
  12377=>"010101110",
  12378=>"110010010",
  12379=>"111111001",
  12380=>"111011010",
  12381=>"001111111",
  12382=>"000011010",
  12383=>"101010000",
  12384=>"011000010",
  12385=>"111001011",
  12386=>"001111011",
  12387=>"011000000",
  12388=>"101100100",
  12389=>"110010110",
  12390=>"011110101",
  12391=>"111010110",
  12392=>"000110110",
  12393=>"001010111",
  12394=>"000010001",
  12395=>"100101100",
  12396=>"111100001",
  12397=>"010000010",
  12398=>"011011100",
  12399=>"010110010",
  12400=>"010000000",
  12401=>"111101000",
  12402=>"011001110",
  12403=>"100101100",
  12404=>"110000100",
  12405=>"110000111",
  12406=>"100110101",
  12407=>"110110011",
  12408=>"011001110",
  12409=>"001101000",
  12410=>"111100101",
  12411=>"101001010",
  12412=>"001001101",
  12413=>"101011000",
  12414=>"000011001",
  12415=>"101001111",
  12416=>"110001001",
  12417=>"111000111",
  12418=>"010010111",
  12419=>"110000001",
  12420=>"101000000",
  12421=>"010001000",
  12422=>"011100100",
  12423=>"011111111",
  12424=>"000001000",
  12425=>"000000000",
  12426=>"101010111",
  12427=>"001011010",
  12428=>"001001110",
  12429=>"010001000",
  12430=>"000011011",
  12431=>"001001011",
  12432=>"100110001",
  12433=>"000011101",
  12434=>"000011110",
  12435=>"111101101",
  12436=>"111000101",
  12437=>"110011100",
  12438=>"010000111",
  12439=>"101000100",
  12440=>"011100110",
  12441=>"000100110",
  12442=>"100101011",
  12443=>"001001000",
  12444=>"100010111",
  12445=>"000011011",
  12446=>"000100101",
  12447=>"010110101",
  12448=>"001110010",
  12449=>"100110010",
  12450=>"001011010",
  12451=>"110011011",
  12452=>"001011011",
  12453=>"000110010",
  12454=>"111110010",
  12455=>"111011011",
  12456=>"101010011",
  12457=>"111101000",
  12458=>"000101110",
  12459=>"110001011",
  12460=>"000000101",
  12461=>"010101101",
  12462=>"101110101",
  12463=>"100010111",
  12464=>"011101001",
  12465=>"000010000",
  12466=>"011100011",
  12467=>"101110001",
  12468=>"101101011",
  12469=>"010100000",
  12470=>"010011100",
  12471=>"001100000",
  12472=>"000000100",
  12473=>"000101001",
  12474=>"111010111",
  12475=>"001101110",
  12476=>"100011001",
  12477=>"000101011",
  12478=>"110010111",
  12479=>"101001100",
  12480=>"011000000",
  12481=>"010011101",
  12482=>"010111101",
  12483=>"010100000",
  12484=>"000101111",
  12485=>"101001111",
  12486=>"001000011",
  12487=>"100100001",
  12488=>"111111101",
  12489=>"011101010",
  12490=>"000110001",
  12491=>"011011100",
  12492=>"100110100",
  12493=>"011110111",
  12494=>"010111000",
  12495=>"111101010",
  12496=>"011100011",
  12497=>"110100111",
  12498=>"101111011",
  12499=>"001010100",
  12500=>"100110000",
  12501=>"001010010",
  12502=>"101100001",
  12503=>"000000000",
  12504=>"101111100",
  12505=>"010000100",
  12506=>"001101000",
  12507=>"010001000",
  12508=>"101000001",
  12509=>"101011101",
  12510=>"101101000",
  12511=>"101111100",
  12512=>"100101000",
  12513=>"101100001",
  12514=>"001111011",
  12515=>"000010100",
  12516=>"111010100",
  12517=>"101111001",
  12518=>"000001010",
  12519=>"111001110",
  12520=>"001001010",
  12521=>"101111010",
  12522=>"000011110",
  12523=>"111111101",
  12524=>"001101010",
  12525=>"011101110",
  12526=>"100011111",
  12527=>"100001000",
  12528=>"010111010",
  12529=>"110010010",
  12530=>"110000111",
  12531=>"100001001",
  12532=>"000101100",
  12533=>"000001010",
  12534=>"110010011",
  12535=>"010111001",
  12536=>"001100101",
  12537=>"111111110",
  12538=>"001001001",
  12539=>"101001010",
  12540=>"111100001",
  12541=>"100101001",
  12542=>"000111101",
  12543=>"111101010",
  12544=>"001011110",
  12545=>"010010001",
  12546=>"111000001",
  12547=>"100011110",
  12548=>"000111100",
  12549=>"001100100",
  12550=>"111111011",
  12551=>"100010101",
  12552=>"001100000",
  12553=>"001111100",
  12554=>"111011111",
  12555=>"110110111",
  12556=>"110110111",
  12557=>"010101010",
  12558=>"000001001",
  12559=>"111100100",
  12560=>"011101111",
  12561=>"101010001",
  12562=>"001100010",
  12563=>"010011010",
  12564=>"100101101",
  12565=>"001101101",
  12566=>"101100111",
  12567=>"110011001",
  12568=>"011100001",
  12569=>"010000101",
  12570=>"101110100",
  12571=>"011010000",
  12572=>"100111011",
  12573=>"110110000",
  12574=>"110101000",
  12575=>"001100101",
  12576=>"111100101",
  12577=>"110101000",
  12578=>"111000101",
  12579=>"000111011",
  12580=>"101100111",
  12581=>"111110100",
  12582=>"000100100",
  12583=>"111000010",
  12584=>"000100110",
  12585=>"010010111",
  12586=>"101000011",
  12587=>"011001101",
  12588=>"111100000",
  12589=>"111111101",
  12590=>"000001110",
  12591=>"000101000",
  12592=>"100100100",
  12593=>"010100101",
  12594=>"101110001",
  12595=>"001001101",
  12596=>"001100011",
  12597=>"110111000",
  12598=>"011110001",
  12599=>"001100000",
  12600=>"100101010",
  12601=>"101011001",
  12602=>"111001010",
  12603=>"000001011",
  12604=>"001101110",
  12605=>"011100000",
  12606=>"010010100",
  12607=>"010110000",
  12608=>"001001011",
  12609=>"101000011",
  12610=>"100101101",
  12611=>"010100010",
  12612=>"100100000",
  12613=>"010010011",
  12614=>"001010101",
  12615=>"000101101",
  12616=>"000111111",
  12617=>"001101011",
  12618=>"101011100",
  12619=>"111001110",
  12620=>"011000111",
  12621=>"110101010",
  12622=>"000010101",
  12623=>"010000000",
  12624=>"010001000",
  12625=>"001111000",
  12626=>"110011101",
  12627=>"010010101",
  12628=>"111100110",
  12629=>"000011101",
  12630=>"110111101",
  12631=>"111110000",
  12632=>"101101010",
  12633=>"001100110",
  12634=>"000100011",
  12635=>"100000011",
  12636=>"011111010",
  12637=>"000100010",
  12638=>"110101101",
  12639=>"010101111",
  12640=>"000010110",
  12641=>"110011101",
  12642=>"000010110",
  12643=>"010000101",
  12644=>"010010111",
  12645=>"000110110",
  12646=>"010011001",
  12647=>"000001000",
  12648=>"011010010",
  12649=>"111010101",
  12650=>"000010011",
  12651=>"001011011",
  12652=>"011000011",
  12653=>"101110110",
  12654=>"010010000",
  12655=>"001100011",
  12656=>"101001010",
  12657=>"010010010",
  12658=>"100001000",
  12659=>"010000111",
  12660=>"110101001",
  12661=>"110111100",
  12662=>"001010011",
  12663=>"011100000",
  12664=>"001101000",
  12665=>"100110001",
  12666=>"111100011",
  12667=>"010111011",
  12668=>"101011010",
  12669=>"101101001",
  12670=>"001011001",
  12671=>"101101100",
  12672=>"000101110",
  12673=>"010000001",
  12674=>"110111011",
  12675=>"111010111",
  12676=>"111110101",
  12677=>"000010000",
  12678=>"001000000",
  12679=>"000011101",
  12680=>"001000101",
  12681=>"100101101",
  12682=>"100000011",
  12683=>"100100011",
  12684=>"110111111",
  12685=>"110011001",
  12686=>"100100111",
  12687=>"101011100",
  12688=>"000100110",
  12689=>"000100101",
  12690=>"001110110",
  12691=>"001001100",
  12692=>"110000011",
  12693=>"010100011",
  12694=>"111010111",
  12695=>"001000100",
  12696=>"110110110",
  12697=>"000101001",
  12698=>"110001111",
  12699=>"100011111",
  12700=>"000001100",
  12701=>"111001111",
  12702=>"001111101",
  12703=>"000001111",
  12704=>"101011101",
  12705=>"011111011",
  12706=>"110000110",
  12707=>"010011010",
  12708=>"011000010",
  12709=>"000101110",
  12710=>"000111110",
  12711=>"000111010",
  12712=>"100000100",
  12713=>"001101100",
  12714=>"100000111",
  12715=>"000101110",
  12716=>"111001000",
  12717=>"100111100",
  12718=>"001100100",
  12719=>"111111001",
  12720=>"001001011",
  12721=>"010010011",
  12722=>"001111010",
  12723=>"101101100",
  12724=>"001111010",
  12725=>"100011001",
  12726=>"100000110",
  12727=>"100101100",
  12728=>"000110111",
  12729=>"011110100",
  12730=>"001011010",
  12731=>"110110101",
  12732=>"111010111",
  12733=>"100010111",
  12734=>"111110010",
  12735=>"001110001",
  12736=>"110111110",
  12737=>"110110010",
  12738=>"100111011",
  12739=>"001011000",
  12740=>"000011000",
  12741=>"111110001",
  12742=>"111111010",
  12743=>"001101000",
  12744=>"011001010",
  12745=>"000000011",
  12746=>"100000010",
  12747=>"101110111",
  12748=>"011100110",
  12749=>"001100011",
  12750=>"000000001",
  12751=>"111100100",
  12752=>"101100111",
  12753=>"100001110",
  12754=>"111110001",
  12755=>"000110111",
  12756=>"000001001",
  12757=>"001111110",
  12758=>"011101111",
  12759=>"000110101",
  12760=>"011111111",
  12761=>"011111111",
  12762=>"100011000",
  12763=>"110010110",
  12764=>"101110010",
  12765=>"000111000",
  12766=>"101101000",
  12767=>"100100110",
  12768=>"101111001",
  12769=>"001100101",
  12770=>"111101111",
  12771=>"001001100",
  12772=>"111101101",
  12773=>"110000111",
  12774=>"110011010",
  12775=>"111010101",
  12776=>"001001111",
  12777=>"101010101",
  12778=>"000000000",
  12779=>"011110100",
  12780=>"010100111",
  12781=>"100011000",
  12782=>"101011010",
  12783=>"000100000",
  12784=>"110101011",
  12785=>"000011011",
  12786=>"110111011",
  12787=>"001101000",
  12788=>"000110001",
  12789=>"011100000",
  12790=>"001110100",
  12791=>"110110011",
  12792=>"111010110",
  12793=>"000111010",
  12794=>"001110110",
  12795=>"000000110",
  12796=>"111100011",
  12797=>"110011111",
  12798=>"001011110",
  12799=>"100001111",
  12800=>"000101001",
  12801=>"111011100",
  12802=>"110110110",
  12803=>"110010111",
  12804=>"111101111",
  12805=>"011100100",
  12806=>"000001111",
  12807=>"010010101",
  12808=>"111001011",
  12809=>"101110101",
  12810=>"100111000",
  12811=>"010100010",
  12812=>"000100000",
  12813=>"101001011",
  12814=>"110111011",
  12815=>"110101100",
  12816=>"100001101",
  12817=>"111000111",
  12818=>"000010010",
  12819=>"001000100",
  12820=>"100010100",
  12821=>"010000100",
  12822=>"011110000",
  12823=>"001001111",
  12824=>"000000000",
  12825=>"001000110",
  12826=>"111100010",
  12827=>"001001010",
  12828=>"100100110",
  12829=>"000000000",
  12830=>"011001100",
  12831=>"110000001",
  12832=>"110001110",
  12833=>"100110001",
  12834=>"011110101",
  12835=>"001001101",
  12836=>"110101011",
  12837=>"101111101",
  12838=>"001100110",
  12839=>"100110011",
  12840=>"010110101",
  12841=>"100000001",
  12842=>"000001011",
  12843=>"010110011",
  12844=>"010011111",
  12845=>"001000000",
  12846=>"101111101",
  12847=>"101110011",
  12848=>"101111110",
  12849=>"110111110",
  12850=>"001001101",
  12851=>"000001110",
  12852=>"101001011",
  12853=>"010001000",
  12854=>"100000100",
  12855=>"101111111",
  12856=>"101000100",
  12857=>"001111100",
  12858=>"100011111",
  12859=>"111101010",
  12860=>"111010111",
  12861=>"100100110",
  12862=>"000011110",
  12863=>"111100000",
  12864=>"101010111",
  12865=>"100111110",
  12866=>"100111010",
  12867=>"001011001",
  12868=>"111011001",
  12869=>"111101011",
  12870=>"000001111",
  12871=>"101011100",
  12872=>"000001111",
  12873=>"101111010",
  12874=>"110011010",
  12875=>"101101000",
  12876=>"011100111",
  12877=>"100101000",
  12878=>"100001001",
  12879=>"001111011",
  12880=>"101010111",
  12881=>"011010110",
  12882=>"111011010",
  12883=>"111100001",
  12884=>"100010100",
  12885=>"001000110",
  12886=>"000000101",
  12887=>"100100000",
  12888=>"100001000",
  12889=>"110010100",
  12890=>"000001111",
  12891=>"010101101",
  12892=>"000111011",
  12893=>"111011100",
  12894=>"101000111",
  12895=>"111001110",
  12896=>"100000010",
  12897=>"001011010",
  12898=>"001110000",
  12899=>"010001010",
  12900=>"001001010",
  12901=>"110101111",
  12902=>"001101111",
  12903=>"000101011",
  12904=>"010111111",
  12905=>"111011111",
  12906=>"111001110",
  12907=>"010100111",
  12908=>"101011010",
  12909=>"010011100",
  12910=>"101011001",
  12911=>"111001111",
  12912=>"001001000",
  12913=>"001100000",
  12914=>"011000100",
  12915=>"000010000",
  12916=>"101111001",
  12917=>"110011010",
  12918=>"001111101",
  12919=>"101000100",
  12920=>"111110111",
  12921=>"110101001",
  12922=>"001100101",
  12923=>"101010101",
  12924=>"100011110",
  12925=>"110011001",
  12926=>"100010001",
  12927=>"010110101",
  12928=>"100110100",
  12929=>"001000010",
  12930=>"000000001",
  12931=>"111101111",
  12932=>"101110101",
  12933=>"110101111",
  12934=>"001110100",
  12935=>"010111110",
  12936=>"101000010",
  12937=>"010011000",
  12938=>"101111110",
  12939=>"101101110",
  12940=>"100011101",
  12941=>"011101001",
  12942=>"100110011",
  12943=>"000011010",
  12944=>"010001110",
  12945=>"110000111",
  12946=>"000100001",
  12947=>"111111111",
  12948=>"010110100",
  12949=>"110010110",
  12950=>"011010001",
  12951=>"111101100",
  12952=>"110010001",
  12953=>"111010101",
  12954=>"110110101",
  12955=>"101101010",
  12956=>"000010110",
  12957=>"010000010",
  12958=>"001111101",
  12959=>"000000110",
  12960=>"100100110",
  12961=>"110101000",
  12962=>"111110001",
  12963=>"110111110",
  12964=>"001001001",
  12965=>"101011000",
  12966=>"000110000",
  12967=>"101010101",
  12968=>"001000000",
  12969=>"111011000",
  12970=>"111011111",
  12971=>"011101001",
  12972=>"110011111",
  12973=>"001111111",
  12974=>"110000110",
  12975=>"001000001",
  12976=>"001011111",
  12977=>"100010111",
  12978=>"101111111",
  12979=>"100110011",
  12980=>"100000111",
  12981=>"101001110",
  12982=>"001001110",
  12983=>"000111111",
  12984=>"000001101",
  12985=>"101110100",
  12986=>"110010010",
  12987=>"000011111",
  12988=>"110000010",
  12989=>"001000000",
  12990=>"101000100",
  12991=>"101100111",
  12992=>"101000011",
  12993=>"111111010",
  12994=>"001100110",
  12995=>"001100011",
  12996=>"111000011",
  12997=>"100010000",
  12998=>"011110111",
  12999=>"100110001",
  13000=>"011100001",
  13001=>"110110110",
  13002=>"001101011",
  13003=>"101001001",
  13004=>"010011010",
  13005=>"100101100",
  13006=>"101100111",
  13007=>"010101101",
  13008=>"010111011",
  13009=>"100100101",
  13010=>"010110010",
  13011=>"011001101",
  13012=>"001001000",
  13013=>"110000101",
  13014=>"001110010",
  13015=>"010000101",
  13016=>"100000010",
  13017=>"011011100",
  13018=>"101010000",
  13019=>"101000100",
  13020=>"011111100",
  13021=>"010110010",
  13022=>"001110000",
  13023=>"110101101",
  13024=>"011001101",
  13025=>"110011000",
  13026=>"010011011",
  13027=>"000110011",
  13028=>"001100001",
  13029=>"100000110",
  13030=>"011010010",
  13031=>"101000100",
  13032=>"001000101",
  13033=>"101111111",
  13034=>"100110111",
  13035=>"111000000",
  13036=>"010011011",
  13037=>"100000000",
  13038=>"010011110",
  13039=>"000011001",
  13040=>"011101101",
  13041=>"000011100",
  13042=>"010101110",
  13043=>"010001111",
  13044=>"010010000",
  13045=>"011100010",
  13046=>"111001011",
  13047=>"111010000",
  13048=>"101110011",
  13049=>"111010011",
  13050=>"100100010",
  13051=>"100111010",
  13052=>"100010011",
  13053=>"011111101",
  13054=>"010000110",
  13055=>"001010001",
  13056=>"101111000",
  13057=>"011101111",
  13058=>"101101101",
  13059=>"110111100",
  13060=>"111011001",
  13061=>"110000101",
  13062=>"100100011",
  13063=>"111100010",
  13064=>"111000001",
  13065=>"110010000",
  13066=>"000001110",
  13067=>"001000110",
  13068=>"001110111",
  13069=>"000011100",
  13070=>"111111101",
  13071=>"000000100",
  13072=>"000000101",
  13073=>"001110010",
  13074=>"001011011",
  13075=>"110000001",
  13076=>"111001001",
  13077=>"010010111",
  13078=>"001010010",
  13079=>"001000001",
  13080=>"001001011",
  13081=>"111111010",
  13082=>"110000000",
  13083=>"110000001",
  13084=>"011001110",
  13085=>"000110001",
  13086=>"101111101",
  13087=>"111000001",
  13088=>"100001001",
  13089=>"100001000",
  13090=>"110000000",
  13091=>"101001010",
  13092=>"001010000",
  13093=>"000000000",
  13094=>"000100111",
  13095=>"010110010",
  13096=>"101100001",
  13097=>"100011111",
  13098=>"000001111",
  13099=>"001111010",
  13100=>"000011101",
  13101=>"000101101",
  13102=>"101110001",
  13103=>"111101001",
  13104=>"011101011",
  13105=>"111110100",
  13106=>"100100010",
  13107=>"011111111",
  13108=>"001100010",
  13109=>"000011101",
  13110=>"011111011",
  13111=>"110010000",
  13112=>"100001001",
  13113=>"110111111",
  13114=>"110001100",
  13115=>"011110110",
  13116=>"101001110",
  13117=>"001111101",
  13118=>"011101010",
  13119=>"110010010",
  13120=>"100100010",
  13121=>"100000011",
  13122=>"000111000",
  13123=>"001110110",
  13124=>"001001100",
  13125=>"000110000",
  13126=>"100010100",
  13127=>"001001010",
  13128=>"111010011",
  13129=>"011010010",
  13130=>"110011111",
  13131=>"110110110",
  13132=>"100001010",
  13133=>"101101000",
  13134=>"100000000",
  13135=>"110010010",
  13136=>"101000010",
  13137=>"100001001",
  13138=>"101100100",
  13139=>"111010010",
  13140=>"001000000",
  13141=>"110001001",
  13142=>"100111010",
  13143=>"110101111",
  13144=>"110111000",
  13145=>"001011010",
  13146=>"000110000",
  13147=>"111110000",
  13148=>"110010100",
  13149=>"001111010",
  13150=>"101111001",
  13151=>"100100110",
  13152=>"010001010",
  13153=>"110000100",
  13154=>"000000101",
  13155=>"111100000",
  13156=>"110100101",
  13157=>"001111101",
  13158=>"011011011",
  13159=>"010111000",
  13160=>"011010001",
  13161=>"000010001",
  13162=>"011011110",
  13163=>"101110110",
  13164=>"111100110",
  13165=>"101010010",
  13166=>"111001000",
  13167=>"011010001",
  13168=>"010111111",
  13169=>"101100100",
  13170=>"101011000",
  13171=>"101010111",
  13172=>"011100110",
  13173=>"001100000",
  13174=>"010111111",
  13175=>"010100101",
  13176=>"101001110",
  13177=>"101110001",
  13178=>"001101100",
  13179=>"111110010",
  13180=>"010101000",
  13181=>"110010000",
  13182=>"101100100",
  13183=>"110111010",
  13184=>"111011001",
  13185=>"100101001",
  13186=>"110001000",
  13187=>"101011100",
  13188=>"000010000",
  13189=>"111011011",
  13190=>"111010010",
  13191=>"110000000",
  13192=>"101111100",
  13193=>"010001010",
  13194=>"010010010",
  13195=>"100111110",
  13196=>"000101010",
  13197=>"011110000",
  13198=>"001100001",
  13199=>"110011100",
  13200=>"101000000",
  13201=>"011000001",
  13202=>"001000100",
  13203=>"100110001",
  13204=>"110000111",
  13205=>"001111101",
  13206=>"000011011",
  13207=>"110011110",
  13208=>"111110000",
  13209=>"000011011",
  13210=>"010101000",
  13211=>"100101110",
  13212=>"010011000",
  13213=>"111010111",
  13214=>"100000000",
  13215=>"101111111",
  13216=>"010011100",
  13217=>"000110111",
  13218=>"010111111",
  13219=>"011110000",
  13220=>"010111100",
  13221=>"001001001",
  13222=>"111111111",
  13223=>"101001000",
  13224=>"111111101",
  13225=>"100000000",
  13226=>"011110111",
  13227=>"000000000",
  13228=>"100111000",
  13229=>"010010010",
  13230=>"001110010",
  13231=>"100110010",
  13232=>"111100010",
  13233=>"111100101",
  13234=>"101001111",
  13235=>"010110010",
  13236=>"111100111",
  13237=>"011100110",
  13238=>"000000100",
  13239=>"011100001",
  13240=>"001101101",
  13241=>"111001110",
  13242=>"111110100",
  13243=>"011111111",
  13244=>"000000001",
  13245=>"110011100",
  13246=>"010010011",
  13247=>"111111100",
  13248=>"111111111",
  13249=>"010010110",
  13250=>"110111001",
  13251=>"001011100",
  13252=>"111110001",
  13253=>"011001101",
  13254=>"001110111",
  13255=>"100111101",
  13256=>"011011010",
  13257=>"110101010",
  13258=>"111101110",
  13259=>"011011101",
  13260=>"001001111",
  13261=>"001011101",
  13262=>"110000101",
  13263=>"101110100",
  13264=>"111100000",
  13265=>"100010010",
  13266=>"010001000",
  13267=>"000110111",
  13268=>"011010001",
  13269=>"001111111",
  13270=>"010010100",
  13271=>"011101000",
  13272=>"101001011",
  13273=>"000101111",
  13274=>"001010001",
  13275=>"111101000",
  13276=>"101011001",
  13277=>"100001111",
  13278=>"010101011",
  13279=>"000011011",
  13280=>"110100011",
  13281=>"000100101",
  13282=>"110110101",
  13283=>"100000000",
  13284=>"001110000",
  13285=>"111101111",
  13286=>"011111010",
  13287=>"010100000",
  13288=>"111010010",
  13289=>"110110011",
  13290=>"100000011",
  13291=>"111000100",
  13292=>"011110110",
  13293=>"010110011",
  13294=>"000101101",
  13295=>"010011000",
  13296=>"100010110",
  13297=>"100000000",
  13298=>"101000110",
  13299=>"001100101",
  13300=>"011011010",
  13301=>"111011111",
  13302=>"110001011",
  13303=>"000010111",
  13304=>"010010111",
  13305=>"101001101",
  13306=>"010011110",
  13307=>"110110111",
  13308=>"010001001",
  13309=>"000111101",
  13310=>"100011000",
  13311=>"000011110",
  13312=>"001000011",
  13313=>"010110100",
  13314=>"001110101",
  13315=>"110010010",
  13316=>"000000100",
  13317=>"010100000",
  13318=>"111011011",
  13319=>"110001111",
  13320=>"010011100",
  13321=>"010100000",
  13322=>"110101010",
  13323=>"100110100",
  13324=>"111010101",
  13325=>"101100010",
  13326=>"101010010",
  13327=>"000001101",
  13328=>"001101101",
  13329=>"001001000",
  13330=>"011000110",
  13331=>"110011010",
  13332=>"000001010",
  13333=>"011001011",
  13334=>"101110011",
  13335=>"000001100",
  13336=>"011111000",
  13337=>"011001110",
  13338=>"101100000",
  13339=>"101111111",
  13340=>"001000100",
  13341=>"110110101",
  13342=>"001011010",
  13343=>"100010110",
  13344=>"110010011",
  13345=>"000101111",
  13346=>"010111010",
  13347=>"010011111",
  13348=>"010000000",
  13349=>"110110111",
  13350=>"001110101",
  13351=>"100001101",
  13352=>"110010001",
  13353=>"100111000",
  13354=>"110111011",
  13355=>"001000100",
  13356=>"100010000",
  13357=>"011011111",
  13358=>"010101111",
  13359=>"000101111",
  13360=>"101001100",
  13361=>"101100011",
  13362=>"011001110",
  13363=>"111001111",
  13364=>"000110010",
  13365=>"000000000",
  13366=>"011000001",
  13367=>"110100010",
  13368=>"101100000",
  13369=>"010100000",
  13370=>"011101001",
  13371=>"111111110",
  13372=>"101111001",
  13373=>"110001000",
  13374=>"101110111",
  13375=>"101101100",
  13376=>"011101001",
  13377=>"101101101",
  13378=>"110001001",
  13379=>"001101001",
  13380=>"000111010",
  13381=>"111010001",
  13382=>"000010001",
  13383=>"001001000",
  13384=>"110101010",
  13385=>"011000101",
  13386=>"001010011",
  13387=>"111001101",
  13388=>"010101010",
  13389=>"001011100",
  13390=>"000100111",
  13391=>"000010100",
  13392=>"011100001",
  13393=>"000101100",
  13394=>"001011110",
  13395=>"111100110",
  13396=>"001100111",
  13397=>"001110010",
  13398=>"110000100",
  13399=>"011101110",
  13400=>"110101111",
  13401=>"101000100",
  13402=>"100000100",
  13403=>"100010011",
  13404=>"100011000",
  13405=>"000101000",
  13406=>"001000101",
  13407=>"110110000",
  13408=>"101100001",
  13409=>"001010010",
  13410=>"101101101",
  13411=>"000010001",
  13412=>"010010101",
  13413=>"101101000",
  13414=>"100111110",
  13415=>"001011010",
  13416=>"110010010",
  13417=>"101011010",
  13418=>"111000101",
  13419=>"011100011",
  13420=>"011111011",
  13421=>"110000001",
  13422=>"000011101",
  13423=>"110000111",
  13424=>"000000101",
  13425=>"101110101",
  13426=>"010001011",
  13427=>"101001101",
  13428=>"100011011",
  13429=>"001110111",
  13430=>"111100010",
  13431=>"101001111",
  13432=>"010111000",
  13433=>"111000101",
  13434=>"100001010",
  13435=>"000001111",
  13436=>"000101111",
  13437=>"000001101",
  13438=>"011110010",
  13439=>"100111110",
  13440=>"001010001",
  13441=>"110101000",
  13442=>"100001110",
  13443=>"101111111",
  13444=>"101010111",
  13445=>"101001101",
  13446=>"001010001",
  13447=>"001101011",
  13448=>"110000110",
  13449=>"001110001",
  13450=>"011011011",
  13451=>"011100011",
  13452=>"000101111",
  13453=>"110101010",
  13454=>"111101001",
  13455=>"000011111",
  13456=>"100011000",
  13457=>"101001010",
  13458=>"000010110",
  13459=>"001111101",
  13460=>"101101101",
  13461=>"111001000",
  13462=>"000101111",
  13463=>"011100101",
  13464=>"110110100",
  13465=>"001111010",
  13466=>"101110110",
  13467=>"101000110",
  13468=>"000011000",
  13469=>"011111000",
  13470=>"011110110",
  13471=>"110010011",
  13472=>"000101010",
  13473=>"110000000",
  13474=>"110111110",
  13475=>"100110010",
  13476=>"100011100",
  13477=>"101010001",
  13478=>"110010010",
  13479=>"111001001",
  13480=>"000000101",
  13481=>"100100010",
  13482=>"000110000",
  13483=>"011010001",
  13484=>"010011110",
  13485=>"111101010",
  13486=>"101101100",
  13487=>"001010100",
  13488=>"111101001",
  13489=>"111111110",
  13490=>"100001110",
  13491=>"011110001",
  13492=>"111101010",
  13493=>"001001100",
  13494=>"001001110",
  13495=>"110101010",
  13496=>"100100110",
  13497=>"001101101",
  13498=>"010010101",
  13499=>"011111111",
  13500=>"100111001",
  13501=>"111110000",
  13502=>"000010101",
  13503=>"101001010",
  13504=>"100001101",
  13505=>"000000101",
  13506=>"010111011",
  13507=>"011100010",
  13508=>"010111101",
  13509=>"101101001",
  13510=>"010001011",
  13511=>"110111111",
  13512=>"100000001",
  13513=>"010101110",
  13514=>"110000010",
  13515=>"011101001",
  13516=>"010011101",
  13517=>"000001000",
  13518=>"111000100",
  13519=>"000011000",
  13520=>"010010010",
  13521=>"001001000",
  13522=>"100000000",
  13523=>"110000101",
  13524=>"101000110",
  13525=>"011001001",
  13526=>"100001111",
  13527=>"000001111",
  13528=>"100010111",
  13529=>"001100010",
  13530=>"000010010",
  13531=>"100100011",
  13532=>"101000001",
  13533=>"011110111",
  13534=>"001000101",
  13535=>"111111110",
  13536=>"010011101",
  13537=>"110100101",
  13538=>"001000110",
  13539=>"100110010",
  13540=>"001100001",
  13541=>"010000100",
  13542=>"000011000",
  13543=>"100010001",
  13544=>"001011111",
  13545=>"100010001",
  13546=>"010011111",
  13547=>"000101111",
  13548=>"000001101",
  13549=>"010010111",
  13550=>"010100010",
  13551=>"110001111",
  13552=>"110100100",
  13553=>"111011111",
  13554=>"111111001",
  13555=>"100100010",
  13556=>"000110101",
  13557=>"111000100",
  13558=>"001111000",
  13559=>"001100010",
  13560=>"010001101",
  13561=>"001100101",
  13562=>"001111110",
  13563=>"011001001",
  13564=>"001100101",
  13565=>"111101000",
  13566=>"010010010",
  13567=>"101001000",
  13568=>"111010011",
  13569=>"111010001",
  13570=>"001001100",
  13571=>"010100000",
  13572=>"111100000",
  13573=>"101101111",
  13574=>"010000010",
  13575=>"001011101",
  13576=>"010111111",
  13577=>"000010000",
  13578=>"100110111",
  13579=>"010001010",
  13580=>"010001000",
  13581=>"111000001",
  13582=>"011000000",
  13583=>"110000110",
  13584=>"000101001",
  13585=>"001011101",
  13586=>"010000111",
  13587=>"100011011",
  13588=>"001010011",
  13589=>"000101010",
  13590=>"001000000",
  13591=>"011101100",
  13592=>"100100101",
  13593=>"110110101",
  13594=>"100000101",
  13595=>"101011010",
  13596=>"001001101",
  13597=>"011111001",
  13598=>"010110110",
  13599=>"001011010",
  13600=>"111010100",
  13601=>"100010011",
  13602=>"001011100",
  13603=>"000001111",
  13604=>"101010001",
  13605=>"011001110",
  13606=>"101101011",
  13607=>"100001000",
  13608=>"111010111",
  13609=>"010001000",
  13610=>"001000110",
  13611=>"111101101",
  13612=>"001110011",
  13613=>"100001010",
  13614=>"001000101",
  13615=>"011001111",
  13616=>"101100000",
  13617=>"100111111",
  13618=>"010100000",
  13619=>"000101011",
  13620=>"011010011",
  13621=>"001100010",
  13622=>"000010100",
  13623=>"101001111",
  13624=>"000000001",
  13625=>"101100111",
  13626=>"111110110",
  13627=>"100010000",
  13628=>"100100101",
  13629=>"111011000",
  13630=>"001100101",
  13631=>"110011100",
  13632=>"000110100",
  13633=>"001010000",
  13634=>"000010001",
  13635=>"010110000",
  13636=>"010000000",
  13637=>"010110010",
  13638=>"000000000",
  13639=>"100110100",
  13640=>"011000110",
  13641=>"010101000",
  13642=>"111101101",
  13643=>"011000011",
  13644=>"110100010",
  13645=>"110101110",
  13646=>"010010101",
  13647=>"011101101",
  13648=>"010000101",
  13649=>"111110010",
  13650=>"010010001",
  13651=>"110000001",
  13652=>"101010110",
  13653=>"000011101",
  13654=>"010101101",
  13655=>"000011101",
  13656=>"001001011",
  13657=>"010001001",
  13658=>"100100000",
  13659=>"000001110",
  13660=>"101011001",
  13661=>"110110001",
  13662=>"111110011",
  13663=>"011001001",
  13664=>"011111001",
  13665=>"011101100",
  13666=>"110111001",
  13667=>"100000101",
  13668=>"100101111",
  13669=>"000000110",
  13670=>"010110110",
  13671=>"011111111",
  13672=>"111110100",
  13673=>"010000011",
  13674=>"010110010",
  13675=>"000001101",
  13676=>"100000100",
  13677=>"000001100",
  13678=>"111010011",
  13679=>"010110011",
  13680=>"011010011",
  13681=>"110001001",
  13682=>"011000011",
  13683=>"100101101",
  13684=>"100100100",
  13685=>"101111011",
  13686=>"010101001",
  13687=>"011110010",
  13688=>"111100101",
  13689=>"000110010",
  13690=>"000001000",
  13691=>"011100001",
  13692=>"111011111",
  13693=>"001111100",
  13694=>"000000110",
  13695=>"110101100",
  13696=>"011001111",
  13697=>"000101011",
  13698=>"000000101",
  13699=>"001100001",
  13700=>"011101010",
  13701=>"100000100",
  13702=>"000110111",
  13703=>"000101010",
  13704=>"000110110",
  13705=>"011001001",
  13706=>"110010011",
  13707=>"111111101",
  13708=>"010011000",
  13709=>"011110001",
  13710=>"100001101",
  13711=>"101111111",
  13712=>"011111010",
  13713=>"010001000",
  13714=>"000011001",
  13715=>"111001001",
  13716=>"110100011",
  13717=>"000010110",
  13718=>"010000011",
  13719=>"110011100",
  13720=>"111100110",
  13721=>"000001101",
  13722=>"000001000",
  13723=>"111110101",
  13724=>"110010011",
  13725=>"011100000",
  13726=>"100110010",
  13727=>"100001101",
  13728=>"011100100",
  13729=>"111101001",
  13730=>"110111000",
  13731=>"000001000",
  13732=>"111011110",
  13733=>"111011110",
  13734=>"010010100",
  13735=>"111000000",
  13736=>"101011100",
  13737=>"011000010",
  13738=>"111000010",
  13739=>"010010111",
  13740=>"011111101",
  13741=>"011100011",
  13742=>"111010000",
  13743=>"011001010",
  13744=>"101110101",
  13745=>"100110010",
  13746=>"010000010",
  13747=>"111110111",
  13748=>"011110001",
  13749=>"001111110",
  13750=>"001101011",
  13751=>"111000001",
  13752=>"110111010",
  13753=>"100110111",
  13754=>"010000111",
  13755=>"001010001",
  13756=>"101111010",
  13757=>"001011000",
  13758=>"010100001",
  13759=>"101001001",
  13760=>"101010101",
  13761=>"100000010",
  13762=>"001001001",
  13763=>"001110111",
  13764=>"011111011",
  13765=>"101011001",
  13766=>"100101100",
  13767=>"010000111",
  13768=>"111111111",
  13769=>"111011001",
  13770=>"101001000",
  13771=>"001011011",
  13772=>"010100010",
  13773=>"010101111",
  13774=>"110100100",
  13775=>"101001000",
  13776=>"000110011",
  13777=>"110100101",
  13778=>"001101110",
  13779=>"010011100",
  13780=>"111101101",
  13781=>"100001111",
  13782=>"100110001",
  13783=>"110101011",
  13784=>"111101100",
  13785=>"110001100",
  13786=>"000000101",
  13787=>"011010000",
  13788=>"001110111",
  13789=>"001110001",
  13790=>"111000110",
  13791=>"111011100",
  13792=>"001111111",
  13793=>"011101001",
  13794=>"000010111",
  13795=>"110111111",
  13796=>"100000011",
  13797=>"101111101",
  13798=>"101100001",
  13799=>"110000101",
  13800=>"101001010",
  13801=>"011110011",
  13802=>"100001110",
  13803=>"101010111",
  13804=>"010010110",
  13805=>"000010001",
  13806=>"010110000",
  13807=>"010100010",
  13808=>"010110000",
  13809=>"000111001",
  13810=>"101101001",
  13811=>"001110101",
  13812=>"100110010",
  13813=>"111011100",
  13814=>"010010111",
  13815=>"100111111",
  13816=>"000010111",
  13817=>"000011101",
  13818=>"111001100",
  13819=>"000100011",
  13820=>"000001000",
  13821=>"001000101",
  13822=>"110101011",
  13823=>"101110000",
  13824=>"100100010",
  13825=>"110101001",
  13826=>"001001110",
  13827=>"010111100",
  13828=>"110100000",
  13829=>"101110010",
  13830=>"010000111",
  13831=>"000111110",
  13832=>"110011000",
  13833=>"000100010",
  13834=>"011110010",
  13835=>"101001000",
  13836=>"110001100",
  13837=>"101100000",
  13838=>"001000000",
  13839=>"110111001",
  13840=>"100010001",
  13841=>"000111101",
  13842=>"111000011",
  13843=>"011100010",
  13844=>"010000011",
  13845=>"000111001",
  13846=>"000000001",
  13847=>"101110001",
  13848=>"001011101",
  13849=>"011001110",
  13850=>"010101101",
  13851=>"011100011",
  13852=>"100011110",
  13853=>"111111010",
  13854=>"001001011",
  13855=>"011110011",
  13856=>"101010111",
  13857=>"000100011",
  13858=>"011101100",
  13859=>"101110100",
  13860=>"111100001",
  13861=>"111110010",
  13862=>"000000000",
  13863=>"010110111",
  13864=>"110011100",
  13865=>"000101111",
  13866=>"000111000",
  13867=>"011001011",
  13868=>"010110111",
  13869=>"110110101",
  13870=>"010101101",
  13871=>"111010111",
  13872=>"001000011",
  13873=>"000010001",
  13874=>"000101001",
  13875=>"110001101",
  13876=>"000111000",
  13877=>"100010111",
  13878=>"001111000",
  13879=>"111001101",
  13880=>"000101110",
  13881=>"000110110",
  13882=>"110100100",
  13883=>"010000011",
  13884=>"100001100",
  13885=>"010101000",
  13886=>"001010000",
  13887=>"010111010",
  13888=>"111000000",
  13889=>"101010111",
  13890=>"011110001",
  13891=>"101101001",
  13892=>"001101100",
  13893=>"100101111",
  13894=>"110110111",
  13895=>"110001000",
  13896=>"100011101",
  13897=>"111010001",
  13898=>"111110101",
  13899=>"001001111",
  13900=>"101011100",
  13901=>"011111000",
  13902=>"010001111",
  13903=>"000001001",
  13904=>"101100001",
  13905=>"101110111",
  13906=>"110101101",
  13907=>"011101000",
  13908=>"100000000",
  13909=>"010010100",
  13910=>"001001100",
  13911=>"111100011",
  13912=>"000100001",
  13913=>"010000001",
  13914=>"001000101",
  13915=>"100101110",
  13916=>"000110000",
  13917=>"000111001",
  13918=>"110010111",
  13919=>"000100111",
  13920=>"010000001",
  13921=>"110110110",
  13922=>"001010010",
  13923=>"111011101",
  13924=>"100101000",
  13925=>"000001001",
  13926=>"100010001",
  13927=>"100101101",
  13928=>"101000010",
  13929=>"110110010",
  13930=>"011011000",
  13931=>"010010011",
  13932=>"110010111",
  13933=>"110110011",
  13934=>"001011100",
  13935=>"100010100",
  13936=>"111011111",
  13937=>"010000010",
  13938=>"111000011",
  13939=>"101111100",
  13940=>"001100011",
  13941=>"111000001",
  13942=>"011000000",
  13943=>"100011111",
  13944=>"010010000",
  13945=>"111100001",
  13946=>"010110010",
  13947=>"011010100",
  13948=>"110000100",
  13949=>"011100010",
  13950=>"010001011",
  13951=>"101110001",
  13952=>"011010010",
  13953=>"110100101",
  13954=>"100010100",
  13955=>"011010110",
  13956=>"011001100",
  13957=>"100011010",
  13958=>"110101001",
  13959=>"010011001",
  13960=>"000110101",
  13961=>"011000100",
  13962=>"101010010",
  13963=>"101101100",
  13964=>"001000100",
  13965=>"001111110",
  13966=>"010000100",
  13967=>"001100000",
  13968=>"111110001",
  13969=>"000101110",
  13970=>"000110001",
  13971=>"101011111",
  13972=>"100000101",
  13973=>"100001100",
  13974=>"010100101",
  13975=>"100101111",
  13976=>"010000000",
  13977=>"001100101",
  13978=>"101100010",
  13979=>"110100000",
  13980=>"111010101",
  13981=>"101000010",
  13982=>"110001000",
  13983=>"011100110",
  13984=>"101001001",
  13985=>"011101100",
  13986=>"111100101",
  13987=>"100110000",
  13988=>"011001101",
  13989=>"110010100",
  13990=>"111111111",
  13991=>"110010100",
  13992=>"101011110",
  13993=>"000100000",
  13994=>"010110110",
  13995=>"111001100",
  13996=>"001010100",
  13997=>"010010000",
  13998=>"101101011",
  13999=>"000000010",
  14000=>"111100011",
  14001=>"110000101",
  14002=>"000011100",
  14003=>"010000110",
  14004=>"110100011",
  14005=>"001001011",
  14006=>"101010000",
  14007=>"010011110",
  14008=>"011101100",
  14009=>"111010110",
  14010=>"010100011",
  14011=>"011000100",
  14012=>"011101000",
  14013=>"100111101",
  14014=>"101100010",
  14015=>"001001011",
  14016=>"100010010",
  14017=>"011000100",
  14018=>"111000010",
  14019=>"000000110",
  14020=>"001000110",
  14021=>"000000011",
  14022=>"011111000",
  14023=>"000100000",
  14024=>"010010111",
  14025=>"010000100",
  14026=>"000111100",
  14027=>"101000011",
  14028=>"101001100",
  14029=>"001011101",
  14030=>"111111110",
  14031=>"101111100",
  14032=>"111111001",
  14033=>"111011000",
  14034=>"001001111",
  14035=>"011100000",
  14036=>"100101000",
  14037=>"010011101",
  14038=>"101011111",
  14039=>"000010000",
  14040=>"000111011",
  14041=>"000100110",
  14042=>"111010011",
  14043=>"101101110",
  14044=>"101100101",
  14045=>"111110111",
  14046=>"101101100",
  14047=>"010110101",
  14048=>"101111010",
  14049=>"001110111",
  14050=>"101111000",
  14051=>"000101110",
  14052=>"010011011",
  14053=>"000000111",
  14054=>"000110000",
  14055=>"101001001",
  14056=>"000100111",
  14057=>"001111000",
  14058=>"001011011",
  14059=>"100110011",
  14060=>"000101100",
  14061=>"000111011",
  14062=>"001001010",
  14063=>"111001101",
  14064=>"100001110",
  14065=>"000000100",
  14066=>"100010001",
  14067=>"111100111",
  14068=>"000001100",
  14069=>"110010100",
  14070=>"100110101",
  14071=>"110010100",
  14072=>"010110001",
  14073=>"001100101",
  14074=>"001110100",
  14075=>"001010000",
  14076=>"110111011",
  14077=>"100000000",
  14078=>"100100011",
  14079=>"100110000",
  14080=>"001010011",
  14081=>"101110100",
  14082=>"001111011",
  14083=>"101010001",
  14084=>"011111111",
  14085=>"100000100",
  14086=>"010100100",
  14087=>"100101001",
  14088=>"010010001",
  14089=>"111100100",
  14090=>"010001011",
  14091=>"000110010",
  14092=>"000010100",
  14093=>"000101100",
  14094=>"111010111",
  14095=>"111100001",
  14096=>"000100110",
  14097=>"010000010",
  14098=>"011000001",
  14099=>"001001010",
  14100=>"000101010",
  14101=>"000111010",
  14102=>"101001010",
  14103=>"110001001",
  14104=>"000011110",
  14105=>"001101010",
  14106=>"011011101",
  14107=>"001110100",
  14108=>"010000001",
  14109=>"000110010",
  14110=>"000000000",
  14111=>"010010100",
  14112=>"111111100",
  14113=>"110010011",
  14114=>"111100010",
  14115=>"111111001",
  14116=>"011000111",
  14117=>"011110011",
  14118=>"111010111",
  14119=>"101011100",
  14120=>"000001111",
  14121=>"111100000",
  14122=>"011010111",
  14123=>"010000101",
  14124=>"110001001",
  14125=>"000110011",
  14126=>"111011001",
  14127=>"001111100",
  14128=>"000001011",
  14129=>"101010110",
  14130=>"010000000",
  14131=>"010001100",
  14132=>"110011111",
  14133=>"111001100",
  14134=>"000000100",
  14135=>"011100100",
  14136=>"000001000",
  14137=>"010010100",
  14138=>"001001010",
  14139=>"111011000",
  14140=>"001000000",
  14141=>"000100000",
  14142=>"000101011",
  14143=>"111000100",
  14144=>"010011000",
  14145=>"100000011",
  14146=>"010110110",
  14147=>"011011001",
  14148=>"100010100",
  14149=>"011100111",
  14150=>"111010110",
  14151=>"100100100",
  14152=>"000000110",
  14153=>"110011011",
  14154=>"101101100",
  14155=>"111011100",
  14156=>"100000111",
  14157=>"000011000",
  14158=>"010011111",
  14159=>"100101111",
  14160=>"100110001",
  14161=>"100000001",
  14162=>"101110011",
  14163=>"000010000",
  14164=>"101001101",
  14165=>"110000000",
  14166=>"101010111",
  14167=>"000111000",
  14168=>"011101010",
  14169=>"001000011",
  14170=>"001010111",
  14171=>"000101100",
  14172=>"101000000",
  14173=>"000011001",
  14174=>"001011001",
  14175=>"001001000",
  14176=>"000111111",
  14177=>"110011100",
  14178=>"110010110",
  14179=>"111000111",
  14180=>"011000010",
  14181=>"111111010",
  14182=>"110010111",
  14183=>"000010111",
  14184=>"001000101",
  14185=>"101001101",
  14186=>"100111010",
  14187=>"011111001",
  14188=>"001010010",
  14189=>"101101010",
  14190=>"000001111",
  14191=>"010100110",
  14192=>"010111000",
  14193=>"001011110",
  14194=>"111111010",
  14195=>"111111100",
  14196=>"000110000",
  14197=>"110001110",
  14198=>"100100100",
  14199=>"001100000",
  14200=>"110110111",
  14201=>"001110111",
  14202=>"001101000",
  14203=>"100110111",
  14204=>"000101000",
  14205=>"000110101",
  14206=>"011000101",
  14207=>"110001110",
  14208=>"000100110",
  14209=>"100100111",
  14210=>"111101111",
  14211=>"111011100",
  14212=>"000100010",
  14213=>"001111000",
  14214=>"010101010",
  14215=>"111000010",
  14216=>"110000010",
  14217=>"100111100",
  14218=>"111111111",
  14219=>"100000111",
  14220=>"100001011",
  14221=>"111001000",
  14222=>"000010011",
  14223=>"111010000",
  14224=>"011100111",
  14225=>"111111111",
  14226=>"100010000",
  14227=>"100001000",
  14228=>"101010111",
  14229=>"000001110",
  14230=>"001100000",
  14231=>"011001100",
  14232=>"000100001",
  14233=>"111101111",
  14234=>"101001000",
  14235=>"001101101",
  14236=>"000010010",
  14237=>"000100110",
  14238=>"001110000",
  14239=>"111101101",
  14240=>"011110111",
  14241=>"000001111",
  14242=>"101110011",
  14243=>"010010101",
  14244=>"110010101",
  14245=>"111101001",
  14246=>"110010111",
  14247=>"011011010",
  14248=>"111101000",
  14249=>"110011011",
  14250=>"011010011",
  14251=>"101001000",
  14252=>"111011000",
  14253=>"000111001",
  14254=>"111101110",
  14255=>"010011011",
  14256=>"101100110",
  14257=>"100001111",
  14258=>"000000110",
  14259=>"101011110",
  14260=>"010010110",
  14261=>"001010100",
  14262=>"010000010",
  14263=>"110011011",
  14264=>"010000100",
  14265=>"001001010",
  14266=>"111110111",
  14267=>"111000011",
  14268=>"000001000",
  14269=>"001000000",
  14270=>"001011000",
  14271=>"010000000",
  14272=>"110100101",
  14273=>"000010010",
  14274=>"111001011",
  14275=>"100010010",
  14276=>"001111000",
  14277=>"110001010",
  14278=>"111110100",
  14279=>"001000100",
  14280=>"100010010",
  14281=>"111011101",
  14282=>"101001110",
  14283=>"011111111",
  14284=>"110010011",
  14285=>"100000100",
  14286=>"111000001",
  14287=>"000000111",
  14288=>"110111110",
  14289=>"000000000",
  14290=>"110111101",
  14291=>"110000000",
  14292=>"010111111",
  14293=>"010110001",
  14294=>"000010101",
  14295=>"100100001",
  14296=>"011001010",
  14297=>"001011101",
  14298=>"011010001",
  14299=>"110011001",
  14300=>"101011100",
  14301=>"010100111",
  14302=>"100011011",
  14303=>"001110100",
  14304=>"010100011",
  14305=>"110100111",
  14306=>"011111111",
  14307=>"001111001",
  14308=>"000001110",
  14309=>"111101101",
  14310=>"000010001",
  14311=>"010100010",
  14312=>"000110011",
  14313=>"100001000",
  14314=>"101100101",
  14315=>"011000000",
  14316=>"110000110",
  14317=>"011100100",
  14318=>"111100000",
  14319=>"111011000",
  14320=>"111101100",
  14321=>"110000100",
  14322=>"111011110",
  14323=>"000110011",
  14324=>"001000111",
  14325=>"111101000",
  14326=>"010000111",
  14327=>"000001010",
  14328=>"001110111",
  14329=>"100100010",
  14330=>"010110101",
  14331=>"000111110",
  14332=>"010100001",
  14333=>"000100111",
  14334=>"110111110",
  14335=>"001100110",
  14336=>"001111010",
  14337=>"000001000",
  14338=>"100110000",
  14339=>"010000111",
  14340=>"001100100",
  14341=>"101011011",
  14342=>"010100000",
  14343=>"100110001",
  14344=>"011000000",
  14345=>"011100101",
  14346=>"000101110",
  14347=>"010100110",
  14348=>"100100110",
  14349=>"110100110",
  14350=>"011001100",
  14351=>"110010011",
  14352=>"001100011",
  14353=>"101101111",
  14354=>"011111111",
  14355=>"100101001",
  14356=>"110011011",
  14357=>"100010001",
  14358=>"110010111",
  14359=>"011010100",
  14360=>"111100111",
  14361=>"111001111",
  14362=>"001110100",
  14363=>"110001011",
  14364=>"010101010",
  14365=>"111011111",
  14366=>"011001110",
  14367=>"010010101",
  14368=>"111111011",
  14369=>"000011100",
  14370=>"010101111",
  14371=>"010001000",
  14372=>"111111111",
  14373=>"111001001",
  14374=>"011100100",
  14375=>"111010010",
  14376=>"101101011",
  14377=>"010011110",
  14378=>"011111111",
  14379=>"110000110",
  14380=>"011111111",
  14381=>"111110111",
  14382=>"101100100",
  14383=>"101011000",
  14384=>"110111000",
  14385=>"000000100",
  14386=>"100000100",
  14387=>"000000110",
  14388=>"100000110",
  14389=>"010001100",
  14390=>"000110000",
  14391=>"011111000",
  14392=>"010011100",
  14393=>"101111000",
  14394=>"001111000",
  14395=>"100110101",
  14396=>"010111000",
  14397=>"011101011",
  14398=>"110101001",
  14399=>"010000011",
  14400=>"100000100",
  14401=>"101011110",
  14402=>"011010011",
  14403=>"001001000",
  14404=>"000011001",
  14405=>"000110010",
  14406=>"100111111",
  14407=>"110101011",
  14408=>"001100001",
  14409=>"111010011",
  14410=>"100110001",
  14411=>"110010011",
  14412=>"000011110",
  14413=>"001101101",
  14414=>"100001001",
  14415=>"111111101",
  14416=>"101000110",
  14417=>"111111110",
  14418=>"110101001",
  14419=>"101110010",
  14420=>"010111000",
  14421=>"000011000",
  14422=>"110010010",
  14423=>"011101111",
  14424=>"001100000",
  14425=>"101110010",
  14426=>"101110111",
  14427=>"001111001",
  14428=>"111111001",
  14429=>"101100110",
  14430=>"100110011",
  14431=>"100101110",
  14432=>"000001000",
  14433=>"011010001",
  14434=>"011101011",
  14435=>"000011100",
  14436=>"100101110",
  14437=>"101100100",
  14438=>"011011101",
  14439=>"100110000",
  14440=>"000010001",
  14441=>"000011010",
  14442=>"111001101",
  14443=>"100111100",
  14444=>"001101000",
  14445=>"111000011",
  14446=>"010001100",
  14447=>"001001000",
  14448=>"000100000",
  14449=>"010000001",
  14450=>"111111110",
  14451=>"000101110",
  14452=>"001110111",
  14453=>"001101111",
  14454=>"101101111",
  14455=>"011011001",
  14456=>"001111000",
  14457=>"001111011",
  14458=>"111111000",
  14459=>"001001101",
  14460=>"010100010",
  14461=>"000011110",
  14462=>"000111000",
  14463=>"001111100",
  14464=>"000000000",
  14465=>"110000111",
  14466=>"001000001",
  14467=>"110000100",
  14468=>"001100101",
  14469=>"011011100",
  14470=>"110110110",
  14471=>"011101110",
  14472=>"010001101",
  14473=>"101100101",
  14474=>"011000001",
  14475=>"011000110",
  14476=>"110101110",
  14477=>"110100000",
  14478=>"010000011",
  14479=>"000111101",
  14480=>"111111111",
  14481=>"100000011",
  14482=>"000110111",
  14483=>"000010001",
  14484=>"101111100",
  14485=>"001110101",
  14486=>"101111100",
  14487=>"100100010",
  14488=>"010011000",
  14489=>"011111111",
  14490=>"101101100",
  14491=>"001011011",
  14492=>"011001111",
  14493=>"000011000",
  14494=>"100001111",
  14495=>"100000010",
  14496=>"010010110",
  14497=>"111111010",
  14498=>"110000111",
  14499=>"101110111",
  14500=>"011001101",
  14501=>"101000010",
  14502=>"100010111",
  14503=>"001111010",
  14504=>"011111001",
  14505=>"100101110",
  14506=>"011011100",
  14507=>"011101010",
  14508=>"100111111",
  14509=>"001000001",
  14510=>"000000110",
  14511=>"000010011",
  14512=>"000011111",
  14513=>"101001000",
  14514=>"000010011",
  14515=>"001000101",
  14516=>"111011011",
  14517=>"001000001",
  14518=>"010001010",
  14519=>"010000100",
  14520=>"101001110",
  14521=>"011100011",
  14522=>"000010100",
  14523=>"010011110",
  14524=>"111011110",
  14525=>"011110100",
  14526=>"110110011",
  14527=>"111011011",
  14528=>"110110010",
  14529=>"100011010",
  14530=>"111010010",
  14531=>"110111111",
  14532=>"100111111",
  14533=>"101111100",
  14534=>"001001000",
  14535=>"000000010",
  14536=>"100011001",
  14537=>"101000010",
  14538=>"010100110",
  14539=>"010101001",
  14540=>"110001011",
  14541=>"001001101",
  14542=>"110111010",
  14543=>"001110000",
  14544=>"101000011",
  14545=>"101100100",
  14546=>"000100000",
  14547=>"011011001",
  14548=>"111001101",
  14549=>"011010111",
  14550=>"100010100",
  14551=>"100010110",
  14552=>"010000000",
  14553=>"111011110",
  14554=>"100011111",
  14555=>"100011101",
  14556=>"011011100",
  14557=>"010000110",
  14558=>"010100010",
  14559=>"011110110",
  14560=>"011101000",
  14561=>"011001001",
  14562=>"100011011",
  14563=>"001011001",
  14564=>"111111111",
  14565=>"011011111",
  14566=>"000001111",
  14567=>"001111111",
  14568=>"101101010",
  14569=>"000110111",
  14570=>"000111101",
  14571=>"000100011",
  14572=>"000001100",
  14573=>"000111101",
  14574=>"001000000",
  14575=>"110000110",
  14576=>"111010010",
  14577=>"101011100",
  14578=>"010000000",
  14579=>"111110110",
  14580=>"101011110",
  14581=>"110100011",
  14582=>"001101110",
  14583=>"000000010",
  14584=>"111011001",
  14585=>"010001011",
  14586=>"111010011",
  14587=>"100001000",
  14588=>"110000110",
  14589=>"010011010",
  14590=>"010110000",
  14591=>"111111110",
  14592=>"110111101",
  14593=>"100110010",
  14594=>"110011010",
  14595=>"100011011",
  14596=>"001100100",
  14597=>"010001001",
  14598=>"011001100",
  14599=>"011110100",
  14600=>"010010100",
  14601=>"001000010",
  14602=>"101110111",
  14603=>"101011101",
  14604=>"111001101",
  14605=>"000101110",
  14606=>"100100101",
  14607=>"110001101",
  14608=>"100010000",
  14609=>"010011010",
  14610=>"101110111",
  14611=>"110111110",
  14612=>"101001100",
  14613=>"100101110",
  14614=>"010101111",
  14615=>"000110000",
  14616=>"000110111",
  14617=>"010011001",
  14618=>"000100000",
  14619=>"011111101",
  14620=>"000000111",
  14621=>"000010100",
  14622=>"010011011",
  14623=>"011110000",
  14624=>"010010101",
  14625=>"010011001",
  14626=>"111010000",
  14627=>"000111101",
  14628=>"011010000",
  14629=>"000110001",
  14630=>"100101111",
  14631=>"101100110",
  14632=>"011101001",
  14633=>"101000110",
  14634=>"010111101",
  14635=>"110000010",
  14636=>"000011000",
  14637=>"111100011",
  14638=>"100000110",
  14639=>"000110001",
  14640=>"010001001",
  14641=>"111000110",
  14642=>"100110010",
  14643=>"010101101",
  14644=>"000011100",
  14645=>"111010111",
  14646=>"111110101",
  14647=>"111111101",
  14648=>"110110000",
  14649=>"110001101",
  14650=>"001010010",
  14651=>"010000010",
  14652=>"000110101",
  14653=>"100010100",
  14654=>"001000101",
  14655=>"110011011",
  14656=>"010000011",
  14657=>"000110001",
  14658=>"110111111",
  14659=>"101111100",
  14660=>"001010001",
  14661=>"011011000",
  14662=>"101110001",
  14663=>"101110010",
  14664=>"110100001",
  14665=>"001001000",
  14666=>"000001001",
  14667=>"010000110",
  14668=>"100001010",
  14669=>"100011111",
  14670=>"101100000",
  14671=>"000111000",
  14672=>"100000010",
  14673=>"000100100",
  14674=>"101101011",
  14675=>"111010011",
  14676=>"110101100",
  14677=>"100000010",
  14678=>"100110110",
  14679=>"110101001",
  14680=>"110110011",
  14681=>"010110010",
  14682=>"000100111",
  14683=>"111110010",
  14684=>"111011110",
  14685=>"011110100",
  14686=>"011111010",
  14687=>"100111100",
  14688=>"010101111",
  14689=>"110111111",
  14690=>"101111110",
  14691=>"000011010",
  14692=>"101101100",
  14693=>"000010011",
  14694=>"111100110",
  14695=>"111110101",
  14696=>"011110111",
  14697=>"000101000",
  14698=>"100010110",
  14699=>"010100100",
  14700=>"010111001",
  14701=>"101011001",
  14702=>"111001101",
  14703=>"111111111",
  14704=>"010010111",
  14705=>"100010000",
  14706=>"110010010",
  14707=>"010101101",
  14708=>"000011011",
  14709=>"101111000",
  14710=>"010101110",
  14711=>"110010000",
  14712=>"010100110",
  14713=>"001100001",
  14714=>"011000100",
  14715=>"010011000",
  14716=>"010100001",
  14717=>"101001111",
  14718=>"001001001",
  14719=>"010000010",
  14720=>"011001111",
  14721=>"010110010",
  14722=>"101110010",
  14723=>"000110011",
  14724=>"110011110",
  14725=>"100010111",
  14726=>"110001111",
  14727=>"010011001",
  14728=>"010110110",
  14729=>"101100111",
  14730=>"111000001",
  14731=>"011101010",
  14732=>"011010000",
  14733=>"100010010",
  14734=>"111001010",
  14735=>"010101010",
  14736=>"001011100",
  14737=>"011101110",
  14738=>"000110100",
  14739=>"110010101",
  14740=>"000001010",
  14741=>"101110111",
  14742=>"110111111",
  14743=>"001000010",
  14744=>"101110100",
  14745=>"000010000",
  14746=>"101010011",
  14747=>"111010111",
  14748=>"110111100",
  14749=>"101001011",
  14750=>"010011011",
  14751=>"010011111",
  14752=>"001010100",
  14753=>"101011010",
  14754=>"100000111",
  14755=>"000010000",
  14756=>"001100101",
  14757=>"101000110",
  14758=>"101010100",
  14759=>"000011011",
  14760=>"000000111",
  14761=>"001011001",
  14762=>"011110000",
  14763=>"101010111",
  14764=>"011001111",
  14765=>"111011100",
  14766=>"001000101",
  14767=>"001000001",
  14768=>"010001101",
  14769=>"001000001",
  14770=>"001011110",
  14771=>"000110110",
  14772=>"111000011",
  14773=>"111010001",
  14774=>"001001101",
  14775=>"100001011",
  14776=>"011100100",
  14777=>"010111001",
  14778=>"010010100",
  14779=>"101010010",
  14780=>"110111001",
  14781=>"110110111",
  14782=>"101000111",
  14783=>"010000011",
  14784=>"000101101",
  14785=>"001110100",
  14786=>"111100000",
  14787=>"010011000",
  14788=>"011011001",
  14789=>"110111001",
  14790=>"110001100",
  14791=>"001010000",
  14792=>"100111011",
  14793=>"110110001",
  14794=>"110010001",
  14795=>"010011000",
  14796=>"010000001",
  14797=>"001100111",
  14798=>"101001100",
  14799=>"111010010",
  14800=>"000011110",
  14801=>"001010000",
  14802=>"100101001",
  14803=>"000111010",
  14804=>"000011111",
  14805=>"100000111",
  14806=>"001110011",
  14807=>"000011000",
  14808=>"111010010",
  14809=>"100111001",
  14810=>"110001010",
  14811=>"110100110",
  14812=>"001000111",
  14813=>"000111011",
  14814=>"110000101",
  14815=>"001001010",
  14816=>"000011010",
  14817=>"111111001",
  14818=>"010011001",
  14819=>"100000100",
  14820=>"011101101",
  14821=>"101110000",
  14822=>"100000001",
  14823=>"110101000",
  14824=>"100000100",
  14825=>"010111011",
  14826=>"111010000",
  14827=>"110101111",
  14828=>"000110001",
  14829=>"000011101",
  14830=>"011000100",
  14831=>"001011001",
  14832=>"000011010",
  14833=>"111001011",
  14834=>"110110011",
  14835=>"100101100",
  14836=>"010100010",
  14837=>"110111101",
  14838=>"010001101",
  14839=>"011101011",
  14840=>"000100010",
  14841=>"011101101",
  14842=>"100001001",
  14843=>"101111010",
  14844=>"011001010",
  14845=>"111100101",
  14846=>"011010011",
  14847=>"010001000",
  14848=>"100001110",
  14849=>"001010000",
  14850=>"001011111",
  14851=>"000100011",
  14852=>"100111000",
  14853=>"011010101",
  14854=>"100101100",
  14855=>"001100001",
  14856=>"100110100",
  14857=>"100010001",
  14858=>"001000000",
  14859=>"000000010",
  14860=>"000010101",
  14861=>"010110100",
  14862=>"101011111",
  14863=>"101110000",
  14864=>"000111111",
  14865=>"000101000",
  14866=>"110110110",
  14867=>"111111011",
  14868=>"010110100",
  14869=>"011100100",
  14870=>"011000100",
  14871=>"100100110",
  14872=>"111000011",
  14873=>"001110011",
  14874=>"111011000",
  14875=>"110111001",
  14876=>"001100001",
  14877=>"100000010",
  14878=>"010001011",
  14879=>"001001101",
  14880=>"111101011",
  14881=>"100100010",
  14882=>"010100001",
  14883=>"001110101",
  14884=>"011110011",
  14885=>"010100100",
  14886=>"011001100",
  14887=>"110010011",
  14888=>"011000101",
  14889=>"011010110",
  14890=>"110100000",
  14891=>"001001101",
  14892=>"011101001",
  14893=>"000100000",
  14894=>"111010001",
  14895=>"100110100",
  14896=>"010101110",
  14897=>"111000010",
  14898=>"000001010",
  14899=>"000111110",
  14900=>"010110010",
  14901=>"000100010",
  14902=>"000111001",
  14903=>"100010001",
  14904=>"011101000",
  14905=>"110001101",
  14906=>"001100001",
  14907=>"000100111",
  14908=>"000011111",
  14909=>"000000000",
  14910=>"000001001",
  14911=>"110101100",
  14912=>"100100111",
  14913=>"110010001",
  14914=>"110010000",
  14915=>"000010010",
  14916=>"100000000",
  14917=>"100100111",
  14918=>"000100100",
  14919=>"111101011",
  14920=>"101110000",
  14921=>"000110000",
  14922=>"101101000",
  14923=>"010000101",
  14924=>"000001001",
  14925=>"110100110",
  14926=>"101111111",
  14927=>"100100010",
  14928=>"101011011",
  14929=>"100011000",
  14930=>"001000010",
  14931=>"010010001",
  14932=>"100001100",
  14933=>"000110000",
  14934=>"000110110",
  14935=>"001110010",
  14936=>"111000000",
  14937=>"110001001",
  14938=>"000101100",
  14939=>"100001110",
  14940=>"001011010",
  14941=>"010001100",
  14942=>"010011110",
  14943=>"011110001",
  14944=>"001011111",
  14945=>"001101010",
  14946=>"000011001",
  14947=>"011010101",
  14948=>"011001110",
  14949=>"111111100",
  14950=>"101010010",
  14951=>"010010010",
  14952=>"011001000",
  14953=>"001110001",
  14954=>"101011110",
  14955=>"000100011",
  14956=>"000100010",
  14957=>"100111010",
  14958=>"101011100",
  14959=>"000000000",
  14960=>"110100010",
  14961=>"100001100",
  14962=>"111000001",
  14963=>"000100011",
  14964=>"001101101",
  14965=>"110111011",
  14966=>"100010011",
  14967=>"110101000",
  14968=>"001010000",
  14969=>"011010011",
  14970=>"101100011",
  14971=>"101101000",
  14972=>"111100001",
  14973=>"000010111",
  14974=>"010110111",
  14975=>"000111011",
  14976=>"110000010",
  14977=>"011101001",
  14978=>"011001011",
  14979=>"001011001",
  14980=>"110100010",
  14981=>"100011010",
  14982=>"001010111",
  14983=>"100110110",
  14984=>"010010110",
  14985=>"100100101",
  14986=>"111110101",
  14987=>"110010010",
  14988=>"000000101",
  14989=>"101111110",
  14990=>"111111010",
  14991=>"001110000",
  14992=>"011111111",
  14993=>"011111101",
  14994=>"001011011",
  14995=>"011101111",
  14996=>"111010001",
  14997=>"000001110",
  14998=>"110000100",
  14999=>"100000111",
  15000=>"010001100",
  15001=>"001111011",
  15002=>"000100101",
  15003=>"110010100",
  15004=>"010001110",
  15005=>"001010001",
  15006=>"101010110",
  15007=>"110100010",
  15008=>"100100111",
  15009=>"010110101",
  15010=>"101110010",
  15011=>"101100100",
  15012=>"010101111",
  15013=>"001001101",
  15014=>"010001011",
  15015=>"011111101",
  15016=>"101010110",
  15017=>"001110010",
  15018=>"000001000",
  15019=>"111100000",
  15020=>"101110001",
  15021=>"001101101",
  15022=>"110001000",
  15023=>"110110101",
  15024=>"000111111",
  15025=>"000000000",
  15026=>"001011010",
  15027=>"101101001",
  15028=>"010010011",
  15029=>"110010001",
  15030=>"010111111",
  15031=>"000001010",
  15032=>"100110100",
  15033=>"000000110",
  15034=>"010111010",
  15035=>"101000110",
  15036=>"100101010",
  15037=>"111001001",
  15038=>"100001101",
  15039=>"000010110",
  15040=>"010011011",
  15041=>"110110110",
  15042=>"011001001",
  15043=>"100000111",
  15044=>"010000001",
  15045=>"001100111",
  15046=>"011110010",
  15047=>"111011010",
  15048=>"110000101",
  15049=>"011101001",
  15050=>"001110101",
  15051=>"100010100",
  15052=>"011010010",
  15053=>"100011010",
  15054=>"111011111",
  15055=>"001111011",
  15056=>"011100011",
  15057=>"001100011",
  15058=>"010111100",
  15059=>"011101000",
  15060=>"111111000",
  15061=>"000010010",
  15062=>"101010000",
  15063=>"111100100",
  15064=>"101011000",
  15065=>"100000101",
  15066=>"010111011",
  15067=>"101011101",
  15068=>"000101101",
  15069=>"010000010",
  15070=>"001100010",
  15071=>"000010000",
  15072=>"000100011",
  15073=>"010101110",
  15074=>"101100011",
  15075=>"110111011",
  15076=>"100010010",
  15077=>"101000100",
  15078=>"101111011",
  15079=>"001111000",
  15080=>"000101111",
  15081=>"110001001",
  15082=>"000110010",
  15083=>"010000011",
  15084=>"000000101",
  15085=>"011110110",
  15086=>"101011110",
  15087=>"110011101",
  15088=>"001000000",
  15089=>"111111111",
  15090=>"000000011",
  15091=>"010000111",
  15092=>"100111100",
  15093=>"100101110",
  15094=>"101001101",
  15095=>"011011010",
  15096=>"011101000",
  15097=>"111010111",
  15098=>"111011111",
  15099=>"010011001",
  15100=>"110110110",
  15101=>"110000001",
  15102=>"001101000",
  15103=>"010011001",
  15104=>"000101001",
  15105=>"010000111",
  15106=>"000100101",
  15107=>"000100000",
  15108=>"100111100",
  15109=>"011000010",
  15110=>"001010010",
  15111=>"110111101",
  15112=>"101011111",
  15113=>"000001100",
  15114=>"011111010",
  15115=>"000011100",
  15116=>"100001100",
  15117=>"010100101",
  15118=>"001010111",
  15119=>"111101011",
  15120=>"101111001",
  15121=>"001011011",
  15122=>"011000001",
  15123=>"110011101",
  15124=>"011000100",
  15125=>"100011100",
  15126=>"001010011",
  15127=>"100101000",
  15128=>"111111011",
  15129=>"011000001",
  15130=>"001000111",
  15131=>"001111010",
  15132=>"000001011",
  15133=>"000011000",
  15134=>"011001100",
  15135=>"110000001",
  15136=>"001111111",
  15137=>"111111011",
  15138=>"001100000",
  15139=>"101100011",
  15140=>"001001010",
  15141=>"001010010",
  15142=>"100111110",
  15143=>"101100110",
  15144=>"111000110",
  15145=>"010000101",
  15146=>"111011110",
  15147=>"100100101",
  15148=>"000001110",
  15149=>"100101000",
  15150=>"100111010",
  15151=>"110110101",
  15152=>"110011101",
  15153=>"000100110",
  15154=>"100100000",
  15155=>"111011010",
  15156=>"111110100",
  15157=>"100011000",
  15158=>"100011001",
  15159=>"000101011",
  15160=>"001000000",
  15161=>"000001011",
  15162=>"010110000",
  15163=>"101110010",
  15164=>"001000001",
  15165=>"000001001",
  15166=>"000000010",
  15167=>"101110011",
  15168=>"101000011",
  15169=>"001111110",
  15170=>"001001001",
  15171=>"100010100",
  15172=>"101101000",
  15173=>"000011101",
  15174=>"111101101",
  15175=>"011011001",
  15176=>"011000000",
  15177=>"001101010",
  15178=>"100010110",
  15179=>"101001001",
  15180=>"101100010",
  15181=>"001010101",
  15182=>"110010111",
  15183=>"100010000",
  15184=>"110110000",
  15185=>"110010100",
  15186=>"000000111",
  15187=>"000001111",
  15188=>"010001010",
  15189=>"100111011",
  15190=>"100000010",
  15191=>"010011010",
  15192=>"101010010",
  15193=>"010110011",
  15194=>"001111110",
  15195=>"111011000",
  15196=>"110110011",
  15197=>"101100100",
  15198=>"000110001",
  15199=>"101010001",
  15200=>"010000101",
  15201=>"111100100",
  15202=>"100100111",
  15203=>"010000001",
  15204=>"001001111",
  15205=>"101100001",
  15206=>"010000100",
  15207=>"101010000",
  15208=>"111000100",
  15209=>"000110000",
  15210=>"111010001",
  15211=>"100100101",
  15212=>"100100000",
  15213=>"110000001",
  15214=>"000001000",
  15215=>"110000101",
  15216=>"011000100",
  15217=>"010001001",
  15218=>"011011101",
  15219=>"010011101",
  15220=>"001100000",
  15221=>"010010000",
  15222=>"110100101",
  15223=>"101010101",
  15224=>"001001100",
  15225=>"100100101",
  15226=>"001011010",
  15227=>"011111010",
  15228=>"010001000",
  15229=>"110011010",
  15230=>"100001010",
  15231=>"000100011",
  15232=>"100011100",
  15233=>"100100110",
  15234=>"110011111",
  15235=>"001001011",
  15236=>"111010110",
  15237=>"111001110",
  15238=>"110111000",
  15239=>"001111100",
  15240=>"101100110",
  15241=>"000101011",
  15242=>"111100110",
  15243=>"000101011",
  15244=>"100110111",
  15245=>"110110100",
  15246=>"000110101",
  15247=>"010011110",
  15248=>"010011000",
  15249=>"111101001",
  15250=>"000001110",
  15251=>"101000011",
  15252=>"011100001",
  15253=>"001111111",
  15254=>"101011111",
  15255=>"011100010",
  15256=>"100011100",
  15257=>"101110001",
  15258=>"110110010",
  15259=>"001110010",
  15260=>"010001000",
  15261=>"001010000",
  15262=>"110000011",
  15263=>"101000111",
  15264=>"111000101",
  15265=>"010111111",
  15266=>"101110101",
  15267=>"010100101",
  15268=>"100100001",
  15269=>"111111011",
  15270=>"001011000",
  15271=>"000001000",
  15272=>"000010011",
  15273=>"111100101",
  15274=>"110010111",
  15275=>"101111011",
  15276=>"010010111",
  15277=>"100000111",
  15278=>"100010010",
  15279=>"101000010",
  15280=>"010101010",
  15281=>"011101011",
  15282=>"010011011",
  15283=>"000110100",
  15284=>"110111100",
  15285=>"000110001",
  15286=>"111011000",
  15287=>"001010110",
  15288=>"100111100",
  15289=>"011000000",
  15290=>"110010000",
  15291=>"111000101",
  15292=>"001100110",
  15293=>"010011110",
  15294=>"000110000",
  15295=>"011001001",
  15296=>"010110010",
  15297=>"000100001",
  15298=>"011101001",
  15299=>"000011011",
  15300=>"100010010",
  15301=>"010001000",
  15302=>"111110110",
  15303=>"110000111",
  15304=>"000000010",
  15305=>"000110000",
  15306=>"100101110",
  15307=>"100100011",
  15308=>"000011101",
  15309=>"010001110",
  15310=>"101010000",
  15311=>"000110011",
  15312=>"010111111",
  15313=>"111101111",
  15314=>"110111111",
  15315=>"111010000",
  15316=>"011100001",
  15317=>"100111001",
  15318=>"100011101",
  15319=>"010110000",
  15320=>"011010111",
  15321=>"010111100",
  15322=>"100001010",
  15323=>"001011000",
  15324=>"111101110",
  15325=>"100000110",
  15326=>"111011001",
  15327=>"110101011",
  15328=>"101100110",
  15329=>"001111101",
  15330=>"001001010",
  15331=>"010001111",
  15332=>"110011000",
  15333=>"111001000",
  15334=>"001001000",
  15335=>"100011010",
  15336=>"100010000",
  15337=>"100011010",
  15338=>"111001011",
  15339=>"001111111",
  15340=>"101000100",
  15341=>"100100001",
  15342=>"010110010",
  15343=>"100001111",
  15344=>"000110111",
  15345=>"101110101",
  15346=>"111111010",
  15347=>"111110101",
  15348=>"001001010",
  15349=>"000001100",
  15350=>"100101101",
  15351=>"110110111",
  15352=>"100111101",
  15353=>"110111101",
  15354=>"101011100",
  15355=>"101011111",
  15356=>"001001001",
  15357=>"101100100",
  15358=>"101110001",
  15359=>"011100011",
  15360=>"111111001",
  15361=>"010000000",
  15362=>"001011110",
  15363=>"001101110",
  15364=>"010011101",
  15365=>"101000111",
  15366=>"111111001",
  15367=>"101011111",
  15368=>"000101100",
  15369=>"000001110",
  15370=>"001110010",
  15371=>"011110000",
  15372=>"011011011",
  15373=>"101001001",
  15374=>"011100011",
  15375=>"000101000",
  15376=>"011111000",
  15377=>"001101011",
  15378=>"100111111",
  15379=>"010011011",
  15380=>"001001100",
  15381=>"010111111",
  15382=>"010101101",
  15383=>"000011000",
  15384=>"101000001",
  15385=>"111011011",
  15386=>"000000110",
  15387=>"111011010",
  15388=>"011111011",
  15389=>"000101010",
  15390=>"110101111",
  15391=>"010100010",
  15392=>"001100101",
  15393=>"100101000",
  15394=>"010101011",
  15395=>"101101110",
  15396=>"111100000",
  15397=>"111000000",
  15398=>"000001111",
  15399=>"111011100",
  15400=>"001100011",
  15401=>"011110010",
  15402=>"110101101",
  15403=>"000100011",
  15404=>"110000100",
  15405=>"100001010",
  15406=>"000011011",
  15407=>"100110011",
  15408=>"010101111",
  15409=>"111100000",
  15410=>"011101010",
  15411=>"100110101",
  15412=>"100011000",
  15413=>"011000010",
  15414=>"100000010",
  15415=>"110000010",
  15416=>"000011001",
  15417=>"001101100",
  15418=>"111101101",
  15419=>"011000011",
  15420=>"110101011",
  15421=>"010001010",
  15422=>"101111001",
  15423=>"101011111",
  15424=>"110101000",
  15425=>"101000100",
  15426=>"010010110",
  15427=>"111011101",
  15428=>"101100100",
  15429=>"100100101",
  15430=>"001100001",
  15431=>"000110111",
  15432=>"000100110",
  15433=>"110001010",
  15434=>"101000000",
  15435=>"001101111",
  15436=>"101001001",
  15437=>"111100111",
  15438=>"101101000",
  15439=>"000001111",
  15440=>"100110010",
  15441=>"000110001",
  15442=>"010101101",
  15443=>"000001011",
  15444=>"100001000",
  15445=>"101101010",
  15446=>"000011111",
  15447=>"001111101",
  15448=>"000101001",
  15449=>"001010111",
  15450=>"000011100",
  15451=>"001000110",
  15452=>"010011111",
  15453=>"000111101",
  15454=>"010000001",
  15455=>"001000101",
  15456=>"000001101",
  15457=>"111001011",
  15458=>"111001011",
  15459=>"010100010",
  15460=>"011100100",
  15461=>"010000100",
  15462=>"010001011",
  15463=>"100110010",
  15464=>"101010001",
  15465=>"010101101",
  15466=>"101100011",
  15467=>"001111101",
  15468=>"001111001",
  15469=>"000100110",
  15470=>"010001101",
  15471=>"111110011",
  15472=>"110010111",
  15473=>"010100001",
  15474=>"101111011",
  15475=>"011110000",
  15476=>"101111101",
  15477=>"001000100",
  15478=>"111110001",
  15479=>"010001010",
  15480=>"010101101",
  15481=>"100111010",
  15482=>"001001010",
  15483=>"100001110",
  15484=>"010000100",
  15485=>"011110100",
  15486=>"000000010",
  15487=>"100110101",
  15488=>"011000110",
  15489=>"011110101",
  15490=>"000111010",
  15491=>"000101110",
  15492=>"101000100",
  15493=>"001000011",
  15494=>"100000001",
  15495=>"010010010",
  15496=>"111111110",
  15497=>"001000000",
  15498=>"110011000",
  15499=>"110111001",
  15500=>"111101110",
  15501=>"110001011",
  15502=>"010110101",
  15503=>"110001100",
  15504=>"110011010",
  15505=>"001011000",
  15506=>"001010010",
  15507=>"111111111",
  15508=>"000011110",
  15509=>"101111111",
  15510=>"110010110",
  15511=>"000100010",
  15512=>"000000001",
  15513=>"111001110",
  15514=>"000010011",
  15515=>"101000110",
  15516=>"111100011",
  15517=>"100001001",
  15518=>"010011000",
  15519=>"011000110",
  15520=>"000100001",
  15521=>"000010100",
  15522=>"110111100",
  15523=>"100010000",
  15524=>"110011111",
  15525=>"110111100",
  15526=>"111101110",
  15527=>"010010010",
  15528=>"000111110",
  15529=>"011101000",
  15530=>"100001111",
  15531=>"101101101",
  15532=>"110000101",
  15533=>"101101100",
  15534=>"101111110",
  15535=>"110000101",
  15536=>"001010010",
  15537=>"111001100",
  15538=>"110101010",
  15539=>"000001011",
  15540=>"010011010",
  15541=>"111010001",
  15542=>"010000011",
  15543=>"011110000",
  15544=>"000001000",
  15545=>"111001111",
  15546=>"011010110",
  15547=>"000001000",
  15548=>"011100011",
  15549=>"110100000",
  15550=>"111101110",
  15551=>"010000100",
  15552=>"111011100",
  15553=>"110100100",
  15554=>"110110000",
  15555=>"011011101",
  15556=>"110010011",
  15557=>"001100001",
  15558=>"111101100",
  15559=>"101000100",
  15560=>"100011101",
  15561=>"000101101",
  15562=>"001111000",
  15563=>"100010111",
  15564=>"110100001",
  15565=>"111101011",
  15566=>"000000011",
  15567=>"111111111",
  15568=>"010010101",
  15569=>"000111001",
  15570=>"001101101",
  15571=>"000000100",
  15572=>"110001101",
  15573=>"001000101",
  15574=>"001101010",
  15575=>"001001101",
  15576=>"010110111",
  15577=>"111111110",
  15578=>"011100010",
  15579=>"000110011",
  15580=>"001101110",
  15581=>"000101110",
  15582=>"100101000",
  15583=>"010010011",
  15584=>"101000000",
  15585=>"010100101",
  15586=>"000011010",
  15587=>"101101000",
  15588=>"111100110",
  15589=>"011011011",
  15590=>"010111000",
  15591=>"001111010",
  15592=>"001100001",
  15593=>"011010001",
  15594=>"111010001",
  15595=>"001011000",
  15596=>"101000010",
  15597=>"111010011",
  15598=>"000000101",
  15599=>"110100010",
  15600=>"001011100",
  15601=>"010111111",
  15602=>"000011010",
  15603=>"101001111",
  15604=>"010010100",
  15605=>"101100110",
  15606=>"101110100",
  15607=>"010001010",
  15608=>"101000001",
  15609=>"011101101",
  15610=>"101011101",
  15611=>"001001010",
  15612=>"100010011",
  15613=>"000111000",
  15614=>"110110111",
  15615=>"111111001",
  15616=>"000000000",
  15617=>"100001001",
  15618=>"100111001",
  15619=>"001001110",
  15620=>"000001110",
  15621=>"110111100",
  15622=>"101101001",
  15623=>"000101100",
  15624=>"101100011",
  15625=>"001000001",
  15626=>"111011100",
  15627=>"101100100",
  15628=>"111111100",
  15629=>"101000111",
  15630=>"010101001",
  15631=>"010011001",
  15632=>"010010000",
  15633=>"100111100",
  15634=>"010000010",
  15635=>"110110100",
  15636=>"011011000",
  15637=>"011110011",
  15638=>"000101111",
  15639=>"010000111",
  15640=>"110101011",
  15641=>"111001011",
  15642=>"000010100",
  15643=>"111101100",
  15644=>"011011100",
  15645=>"111000000",
  15646=>"000111111",
  15647=>"001111100",
  15648=>"001110100",
  15649=>"110100110",
  15650=>"111000000",
  15651=>"110001110",
  15652=>"111000110",
  15653=>"010011010",
  15654=>"100110001",
  15655=>"111011011",
  15656=>"001001010",
  15657=>"100100111",
  15658=>"100000111",
  15659=>"111110001",
  15660=>"001000100",
  15661=>"110110100",
  15662=>"100111111",
  15663=>"000110101",
  15664=>"111100010",
  15665=>"010000000",
  15666=>"011011011",
  15667=>"011110110",
  15668=>"000010100",
  15669=>"001011011",
  15670=>"110000001",
  15671=>"010101101",
  15672=>"100101000",
  15673=>"001101010",
  15674=>"111101011",
  15675=>"110110100",
  15676=>"111111100",
  15677=>"110110110",
  15678=>"011110110",
  15679=>"110001110",
  15680=>"000111010",
  15681=>"000010100",
  15682=>"001001101",
  15683=>"001010000",
  15684=>"001110111",
  15685=>"110101001",
  15686=>"000000000",
  15687=>"001010001",
  15688=>"111110100",
  15689=>"111000100",
  15690=>"000010100",
  15691=>"100100011",
  15692=>"010101110",
  15693=>"111011111",
  15694=>"100100000",
  15695=>"000001110",
  15696=>"011110011",
  15697=>"100001000",
  15698=>"000010100",
  15699=>"011101010",
  15700=>"110010101",
  15701=>"100011101",
  15702=>"111101110",
  15703=>"110100111",
  15704=>"000100001",
  15705=>"000110110",
  15706=>"000101110",
  15707=>"111100000",
  15708=>"011011001",
  15709=>"001110010",
  15710=>"100000100",
  15711=>"101001110",
  15712=>"111100011",
  15713=>"111011110",
  15714=>"000000101",
  15715=>"101001011",
  15716=>"011001111",
  15717=>"010100110",
  15718=>"000010100",
  15719=>"110010111",
  15720=>"010110001",
  15721=>"000011011",
  15722=>"110100000",
  15723=>"011001000",
  15724=>"001011100",
  15725=>"100110100",
  15726=>"100110110",
  15727=>"101110100",
  15728=>"000110001",
  15729=>"010011111",
  15730=>"011100101",
  15731=>"110100111",
  15732=>"000101111",
  15733=>"100011011",
  15734=>"011001101",
  15735=>"111011010",
  15736=>"011101110",
  15737=>"000011010",
  15738=>"100000011",
  15739=>"001010000",
  15740=>"100010010",
  15741=>"100111101",
  15742=>"000100011",
  15743=>"010100100",
  15744=>"010000011",
  15745=>"100011110",
  15746=>"011111001",
  15747=>"110110101",
  15748=>"100110100",
  15749=>"111110110",
  15750=>"000011101",
  15751=>"000000101",
  15752=>"000010001",
  15753=>"001011010",
  15754=>"010010101",
  15755=>"101111101",
  15756=>"010110101",
  15757=>"111011000",
  15758=>"100001000",
  15759=>"101000101",
  15760=>"111101110",
  15761=>"111000000",
  15762=>"101101011",
  15763=>"101001100",
  15764=>"011111110",
  15765=>"100001111",
  15766=>"100001001",
  15767=>"111101110",
  15768=>"110101011",
  15769=>"101001101",
  15770=>"000000000",
  15771=>"110001100",
  15772=>"001100010",
  15773=>"011010101",
  15774=>"111001110",
  15775=>"010111000",
  15776=>"101000000",
  15777=>"110001000",
  15778=>"001000101",
  15779=>"110100111",
  15780=>"100010111",
  15781=>"000100010",
  15782=>"000000101",
  15783=>"111111101",
  15784=>"010111001",
  15785=>"001000111",
  15786=>"100101001",
  15787=>"011101010",
  15788=>"111111000",
  15789=>"110010011",
  15790=>"001001001",
  15791=>"111001000",
  15792=>"110000010",
  15793=>"101110011",
  15794=>"111110010",
  15795=>"001100001",
  15796=>"000101100",
  15797=>"100001101",
  15798=>"110101101",
  15799=>"000111001",
  15800=>"100011010",
  15801=>"010100011",
  15802=>"110110010",
  15803=>"101101101",
  15804=>"110010111",
  15805=>"010000001",
  15806=>"101101111",
  15807=>"110011110",
  15808=>"101000001",
  15809=>"010011011",
  15810=>"101100101",
  15811=>"110000111",
  15812=>"000010000",
  15813=>"101100000",
  15814=>"000010011",
  15815=>"111101000",
  15816=>"001001010",
  15817=>"110101000",
  15818=>"000010000",
  15819=>"010100110",
  15820=>"001111000",
  15821=>"111011001",
  15822=>"110000000",
  15823=>"110100110",
  15824=>"100111001",
  15825=>"111111101",
  15826=>"011111011",
  15827=>"000011110",
  15828=>"010011000",
  15829=>"100000011",
  15830=>"110000110",
  15831=>"011111000",
  15832=>"011001001",
  15833=>"011111001",
  15834=>"111101110",
  15835=>"111011101",
  15836=>"011010110",
  15837=>"010100100",
  15838=>"000110000",
  15839=>"011010100",
  15840=>"011000000",
  15841=>"100110010",
  15842=>"010110000",
  15843=>"110111111",
  15844=>"000110010",
  15845=>"001111011",
  15846=>"101110011",
  15847=>"101001011",
  15848=>"111001000",
  15849=>"111001111",
  15850=>"011010101",
  15851=>"110111010",
  15852=>"010101111",
  15853=>"111110000",
  15854=>"011001100",
  15855=>"100111011",
  15856=>"110100000",
  15857=>"110001111",
  15858=>"011011110",
  15859=>"010011100",
  15860=>"100101000",
  15861=>"000110001",
  15862=>"110000001",
  15863=>"111110010",
  15864=>"110011110",
  15865=>"110001100",
  15866=>"011111000",
  15867=>"100101111",
  15868=>"000101110",
  15869=>"111011100",
  15870=>"111000011",
  15871=>"010111001",
  15872=>"111010011",
  15873=>"111101001",
  15874=>"011011110",
  15875=>"010010101",
  15876=>"001111110",
  15877=>"001010000",
  15878=>"111101010",
  15879=>"000011001",
  15880=>"100101111",
  15881=>"111011111",
  15882=>"010101000",
  15883=>"110001100",
  15884=>"011011010",
  15885=>"110111110",
  15886=>"000000101",
  15887=>"011101011",
  15888=>"000101111",
  15889=>"000000010",
  15890=>"011101111",
  15891=>"000101000",
  15892=>"011001000",
  15893=>"101000101",
  15894=>"111001110",
  15895=>"111010111",
  15896=>"111110111",
  15897=>"000100111",
  15898=>"001100010",
  15899=>"100101100",
  15900=>"111000111",
  15901=>"101110111",
  15902=>"010011101",
  15903=>"101101111",
  15904=>"101000000",
  15905=>"111001110",
  15906=>"010001000",
  15907=>"111110001",
  15908=>"101111100",
  15909=>"011010111",
  15910=>"111010100",
  15911=>"010101101",
  15912=>"101100011",
  15913=>"111011010",
  15914=>"101001100",
  15915=>"101011000",
  15916=>"000010001",
  15917=>"100001110",
  15918=>"110100010",
  15919=>"011101101",
  15920=>"110001100",
  15921=>"001011101",
  15922=>"100010100",
  15923=>"101010001",
  15924=>"000000010",
  15925=>"100000100",
  15926=>"001111111",
  15927=>"001101010",
  15928=>"111100110",
  15929=>"110101010",
  15930=>"000101001",
  15931=>"100110111",
  15932=>"101011111",
  15933=>"100001000",
  15934=>"010100000",
  15935=>"111111001",
  15936=>"010110011",
  15937=>"100100001",
  15938=>"011101000",
  15939=>"000100000",
  15940=>"001000101",
  15941=>"101010011",
  15942=>"111000101",
  15943=>"001010111",
  15944=>"101000110",
  15945=>"011111010",
  15946=>"000101111",
  15947=>"011110111",
  15948=>"000010000",
  15949=>"101110111",
  15950=>"111011100",
  15951=>"001110001",
  15952=>"110111100",
  15953=>"000001110",
  15954=>"110111100",
  15955=>"011100000",
  15956=>"100100001",
  15957=>"101110110",
  15958=>"100100100",
  15959=>"100011011",
  15960=>"100111100",
  15961=>"100110011",
  15962=>"100001100",
  15963=>"010010111",
  15964=>"001100111",
  15965=>"001010011",
  15966=>"101111101",
  15967=>"000010000",
  15968=>"000010110",
  15969=>"101000001",
  15970=>"011110101",
  15971=>"100001011",
  15972=>"001101011",
  15973=>"000110010",
  15974=>"000001000",
  15975=>"001100001",
  15976=>"011111001",
  15977=>"010000100",
  15978=>"000101100",
  15979=>"101110000",
  15980=>"001111101",
  15981=>"101000101",
  15982=>"011110001",
  15983=>"100011001",
  15984=>"110110000",
  15985=>"010100110",
  15986=>"101110001",
  15987=>"101101011",
  15988=>"100110010",
  15989=>"111110000",
  15990=>"100001001",
  15991=>"100111011",
  15992=>"010101010",
  15993=>"001011101",
  15994=>"000000010",
  15995=>"111000111",
  15996=>"100111001",
  15997=>"000011010",
  15998=>"101101010",
  15999=>"100000101",
  16000=>"110111110",
  16001=>"011000010",
  16002=>"000001001",
  16003=>"001110100",
  16004=>"011011000",
  16005=>"100000010",
  16006=>"011101100",
  16007=>"111100110",
  16008=>"010100111",
  16009=>"010000000",
  16010=>"111000011",
  16011=>"110100111",
  16012=>"000100010",
  16013=>"010110001",
  16014=>"101010110",
  16015=>"100110001",
  16016=>"011111001",
  16017=>"111000110",
  16018=>"001000111",
  16019=>"011000110",
  16020=>"111000000",
  16021=>"100100111",
  16022=>"101101101",
  16023=>"101101000",
  16024=>"011101110",
  16025=>"100001101",
  16026=>"110101101",
  16027=>"000111011",
  16028=>"000010100",
  16029=>"000110000",
  16030=>"111100101",
  16031=>"100000000",
  16032=>"110110001",
  16033=>"010110001",
  16034=>"011011110",
  16035=>"100110011",
  16036=>"000011100",
  16037=>"111000110",
  16038=>"101100100",
  16039=>"001100111",
  16040=>"100010100",
  16041=>"111110100",
  16042=>"001001010",
  16043=>"010101010",
  16044=>"000010010",
  16045=>"011101000",
  16046=>"100100000",
  16047=>"011101011",
  16048=>"101101101",
  16049=>"000100100",
  16050=>"001000000",
  16051=>"000010010",
  16052=>"101110111",
  16053=>"010010101",
  16054=>"011101111",
  16055=>"010010100",
  16056=>"000111010",
  16057=>"010110000",
  16058=>"001111110",
  16059=>"011110111",
  16060=>"001100000",
  16061=>"011110001",
  16062=>"001111101",
  16063=>"100111001",
  16064=>"100000110",
  16065=>"011011111",
  16066=>"011111000",
  16067=>"110101000",
  16068=>"000000010",
  16069=>"100011011",
  16070=>"100011110",
  16071=>"101110111",
  16072=>"000010000",
  16073=>"001001001",
  16074=>"001111000",
  16075=>"000000010",
  16076=>"101111110",
  16077=>"001111111",
  16078=>"010100111",
  16079=>"100100001",
  16080=>"001111010",
  16081=>"001111101",
  16082=>"010111111",
  16083=>"110101010",
  16084=>"011101101",
  16085=>"100000111",
  16086=>"100000010",
  16087=>"100001110",
  16088=>"010100000",
  16089=>"110100000",
  16090=>"010111101",
  16091=>"111101010",
  16092=>"000111101",
  16093=>"010110011",
  16094=>"100001011",
  16095=>"111001001",
  16096=>"000011101",
  16097=>"100101101",
  16098=>"101001100",
  16099=>"100010110",
  16100=>"001000011",
  16101=>"000000101",
  16102=>"101110110",
  16103=>"001110110",
  16104=>"010001001",
  16105=>"101000010",
  16106=>"011000011",
  16107=>"000110000",
  16108=>"001010000",
  16109=>"000010100",
  16110=>"010101001",
  16111=>"001110100",
  16112=>"000111111",
  16113=>"101010001",
  16114=>"111100001",
  16115=>"001000101",
  16116=>"101100101",
  16117=>"100011000",
  16118=>"010000000",
  16119=>"001000100",
  16120=>"010110100",
  16121=>"101110011",
  16122=>"011101110",
  16123=>"110111000",
  16124=>"101101110",
  16125=>"000100101",
  16126=>"110010011",
  16127=>"010100000",
  16128=>"000110001",
  16129=>"010001111",
  16130=>"110001010",
  16131=>"001101000",
  16132=>"001010011",
  16133=>"000101011",
  16134=>"001010101",
  16135=>"110010000",
  16136=>"000000000",
  16137=>"001000011",
  16138=>"010001001",
  16139=>"101000000",
  16140=>"111111110",
  16141=>"101111111",
  16142=>"101010000",
  16143=>"001100000",
  16144=>"010010001",
  16145=>"110100010",
  16146=>"111110100",
  16147=>"110110101",
  16148=>"101101101",
  16149=>"011000100",
  16150=>"110000001",
  16151=>"100001011",
  16152=>"000011000",
  16153=>"000100101",
  16154=>"011101110",
  16155=>"111110100",
  16156=>"000101011",
  16157=>"010011000",
  16158=>"000010101",
  16159=>"010001101",
  16160=>"000101110",
  16161=>"111010000",
  16162=>"010000001",
  16163=>"111001001",
  16164=>"010110100",
  16165=>"110100100",
  16166=>"110010010",
  16167=>"101111010",
  16168=>"110111111",
  16169=>"010001110",
  16170=>"100011111",
  16171=>"010100101",
  16172=>"101000100",
  16173=>"100010001",
  16174=>"001100101",
  16175=>"000110011",
  16176=>"101011011",
  16177=>"000000100",
  16178=>"001001000",
  16179=>"011100111",
  16180=>"111110111",
  16181=>"000011011",
  16182=>"110001000",
  16183=>"001011000",
  16184=>"010001000",
  16185=>"101100101",
  16186=>"110010001",
  16187=>"100010010",
  16188=>"100111111",
  16189=>"001000000",
  16190=>"000101000",
  16191=>"000000000",
  16192=>"111110011",
  16193=>"101100100",
  16194=>"000101101",
  16195=>"001000110",
  16196=>"000110001",
  16197=>"101011010",
  16198=>"000011110",
  16199=>"010110011",
  16200=>"000001101",
  16201=>"111010011",
  16202=>"010001011",
  16203=>"011101001",
  16204=>"100001001",
  16205=>"010100110",
  16206=>"110110001",
  16207=>"000001011",
  16208=>"010110000",
  16209=>"101001000",
  16210=>"011000000",
  16211=>"101101010",
  16212=>"011110111",
  16213=>"111001001",
  16214=>"010010001",
  16215=>"110110111",
  16216=>"110000010",
  16217=>"111010101",
  16218=>"100111111",
  16219=>"100100111",
  16220=>"100011001",
  16221=>"111000100",
  16222=>"110011000",
  16223=>"000100010",
  16224=>"110001000",
  16225=>"010010100",
  16226=>"101111110",
  16227=>"011011000",
  16228=>"100010010",
  16229=>"100011000",
  16230=>"101010111",
  16231=>"001100000",
  16232=>"001010111",
  16233=>"000100000",
  16234=>"101110110",
  16235=>"110011111",
  16236=>"010101110",
  16237=>"001000011",
  16238=>"100100000",
  16239=>"100000111",
  16240=>"110101111",
  16241=>"101011110",
  16242=>"110010101",
  16243=>"111000001",
  16244=>"011100111",
  16245=>"111000110",
  16246=>"110000101",
  16247=>"011111010",
  16248=>"100101011",
  16249=>"110101000",
  16250=>"010010011",
  16251=>"101110100",
  16252=>"111001001",
  16253=>"001101100",
  16254=>"010111100",
  16255=>"101101101",
  16256=>"111000011",
  16257=>"111010001",
  16258=>"000111111",
  16259=>"010000010",
  16260=>"010111110",
  16261=>"011001001",
  16262=>"111010110",
  16263=>"100011110",
  16264=>"001110011",
  16265=>"011101000",
  16266=>"111010001",
  16267=>"110001010",
  16268=>"001110110",
  16269=>"011010010",
  16270=>"011010101",
  16271=>"001011111",
  16272=>"000000101",
  16273=>"000011111",
  16274=>"101111110",
  16275=>"111011000",
  16276=>"001101011",
  16277=>"010101000",
  16278=>"000010000",
  16279=>"011011110",
  16280=>"111011101",
  16281=>"010111000",
  16282=>"101100001",
  16283=>"001010010",
  16284=>"101110010",
  16285=>"111001111",
  16286=>"110000000",
  16287=>"111100001",
  16288=>"101110010",
  16289=>"101100010",
  16290=>"111111101",
  16291=>"101100010",
  16292=>"100101101",
  16293=>"001110111",
  16294=>"001111110",
  16295=>"011010110",
  16296=>"000101010",
  16297=>"000000100",
  16298=>"111111100",
  16299=>"111001011",
  16300=>"001110110",
  16301=>"010001001",
  16302=>"110010100",
  16303=>"000010000",
  16304=>"100111100",
  16305=>"111111110",
  16306=>"100110101",
  16307=>"000011010",
  16308=>"011000111",
  16309=>"000011100",
  16310=>"100111000",
  16311=>"110011110",
  16312=>"001100010",
  16313=>"011110000",
  16314=>"110000010",
  16315=>"101010010",
  16316=>"001001010",
  16317=>"111100110",
  16318=>"110110110",
  16319=>"110100110",
  16320=>"000110001",
  16321=>"000100011",
  16322=>"111011111",
  16323=>"101111001",
  16324=>"111001000",
  16325=>"100011100",
  16326=>"011011101",
  16327=>"101011111",
  16328=>"101011111",
  16329=>"111101100",
  16330=>"000010111",
  16331=>"011011001",
  16332=>"010100110",
  16333=>"000101100",
  16334=>"010000101",
  16335=>"000111000",
  16336=>"001110001",
  16337=>"010001000",
  16338=>"011000001",
  16339=>"010100111",
  16340=>"110010000",
  16341=>"010010101",
  16342=>"110111101",
  16343=>"100110110",
  16344=>"101011101",
  16345=>"011111011",
  16346=>"101100011",
  16347=>"110010010",
  16348=>"100000110",
  16349=>"111111111",
  16350=>"111001111",
  16351=>"010001100",
  16352=>"111001110",
  16353=>"011010101",
  16354=>"001100010",
  16355=>"010001011",
  16356=>"100010110",
  16357=>"001001101",
  16358=>"111010101",
  16359=>"000100101",
  16360=>"000001001",
  16361=>"000010001",
  16362=>"000001001",
  16363=>"010000111",
  16364=>"110000110",
  16365=>"111001100",
  16366=>"001001011",
  16367=>"100101110",
  16368=>"101011101",
  16369=>"011110000",
  16370=>"101001111",
  16371=>"000000001",
  16372=>"110001011",
  16373=>"001110101",
  16374=>"110010100",
  16375=>"100000111",
  16376=>"101101101",
  16377=>"101100110",
  16378=>"000110010",
  16379=>"110000110",
  16380=>"111010100",
  16381=>"011000010",
  16382=>"101110001",
  16383=>"010101010",
  16384=>"000100000",
  16385=>"111111101",
  16386=>"111011010",
  16387=>"011000110",
  16388=>"101101101",
  16389=>"110000011",
  16390=>"101000111",
  16391=>"111001000",
  16392=>"000111000",
  16393=>"010000101",
  16394=>"001101010",
  16395=>"011001111",
  16396=>"000101000",
  16397=>"110101110",
  16398=>"001000011",
  16399=>"001011011",
  16400=>"000110010",
  16401=>"000000111",
  16402=>"101000111",
  16403=>"001011101",
  16404=>"000100011",
  16405=>"011001010",
  16406=>"000011101",
  16407=>"011000010",
  16408=>"111001110",
  16409=>"000111111",
  16410=>"111001000",
  16411=>"100111111",
  16412=>"010001010",
  16413=>"100111101",
  16414=>"000101010",
  16415=>"100111000",
  16416=>"001101111",
  16417=>"010111011",
  16418=>"111011111",
  16419=>"110011000",
  16420=>"100101100",
  16421=>"000111011",
  16422=>"000110100",
  16423=>"111101100",
  16424=>"010000110",
  16425=>"000001010",
  16426=>"011110011",
  16427=>"001000001",
  16428=>"110000011",
  16429=>"100010010",
  16430=>"101001100",
  16431=>"010111010",
  16432=>"101000101",
  16433=>"011001100",
  16434=>"001000101",
  16435=>"010110010",
  16436=>"111111011",
  16437=>"110100000",
  16438=>"100010101",
  16439=>"001111110",
  16440=>"001011111",
  16441=>"010111011",
  16442=>"001001001",
  16443=>"100000110",
  16444=>"001110001",
  16445=>"101001110",
  16446=>"110001111",
  16447=>"000011010",
  16448=>"110111010",
  16449=>"000000110",
  16450=>"011100011",
  16451=>"110110000",
  16452=>"101100011",
  16453=>"001011001",
  16454=>"100100010",
  16455=>"000101010",
  16456=>"101111100",
  16457=>"011100010",
  16458=>"000111101",
  16459=>"110111111",
  16460=>"001111101",
  16461=>"111011111",
  16462=>"011101010",
  16463=>"001110001",
  16464=>"000111101",
  16465=>"010100010",
  16466=>"101001001",
  16467=>"011000000",
  16468=>"010000000",
  16469=>"110010011",
  16470=>"001001000",
  16471=>"000000000",
  16472=>"101011101",
  16473=>"010100101",
  16474=>"000011111",
  16475=>"001011001",
  16476=>"011111011",
  16477=>"100101111",
  16478=>"000001111",
  16479=>"101000001",
  16480=>"101100010",
  16481=>"111000101",
  16482=>"100001111",
  16483=>"001000100",
  16484=>"100000110",
  16485=>"001110001",
  16486=>"110101001",
  16487=>"111010100",
  16488=>"001000010",
  16489=>"111000111",
  16490=>"101101010",
  16491=>"111111101",
  16492=>"000000001",
  16493=>"111110100",
  16494=>"011101010",
  16495=>"100011001",
  16496=>"000011101",
  16497=>"101100111",
  16498=>"010001110",
  16499=>"010000001",
  16500=>"010100111",
  16501=>"010111000",
  16502=>"100100000",
  16503=>"111010111",
  16504=>"000001011",
  16505=>"000110111",
  16506=>"110001110",
  16507=>"011000000",
  16508=>"010010100",
  16509=>"101101100",
  16510=>"011100100",
  16511=>"101010001",
  16512=>"110100011",
  16513=>"011001011",
  16514=>"111000000",
  16515=>"010001000",
  16516=>"111011101",
  16517=>"101010001",
  16518=>"101111011",
  16519=>"000000000",
  16520=>"100010100",
  16521=>"101011011",
  16522=>"101001101",
  16523=>"010000001",
  16524=>"101100000",
  16525=>"010110101",
  16526=>"000001001",
  16527=>"110100000",
  16528=>"111001000",
  16529=>"110101111",
  16530=>"000010011",
  16531=>"100001101",
  16532=>"010101001",
  16533=>"110100110",
  16534=>"111110110",
  16535=>"111100100",
  16536=>"000010000",
  16537=>"110110101",
  16538=>"001110111",
  16539=>"001011011",
  16540=>"001111111",
  16541=>"010110111",
  16542=>"101100110",
  16543=>"101011011",
  16544=>"010111001",
  16545=>"011110111",
  16546=>"001011101",
  16547=>"110010111",
  16548=>"110100000",
  16549=>"011011101",
  16550=>"000101001",
  16551=>"000010001",
  16552=>"011000000",
  16553=>"001101001",
  16554=>"110010010",
  16555=>"101011101",
  16556=>"000100101",
  16557=>"000001011",
  16558=>"011100111",
  16559=>"000000001",
  16560=>"110101111",
  16561=>"000000010",
  16562=>"001000001",
  16563=>"111101000",
  16564=>"111010101",
  16565=>"000011000",
  16566=>"110010001",
  16567=>"011001000",
  16568=>"000000111",
  16569=>"011100101",
  16570=>"000111100",
  16571=>"101110101",
  16572=>"010001010",
  16573=>"111101111",
  16574=>"101110111",
  16575=>"100001010",
  16576=>"100110100",
  16577=>"100111010",
  16578=>"000010011",
  16579=>"001111101",
  16580=>"001000011",
  16581=>"100011010",
  16582=>"000001001",
  16583=>"110100101",
  16584=>"111011110",
  16585=>"000000011",
  16586=>"011100101",
  16587=>"010111111",
  16588=>"010110111",
  16589=>"001100110",
  16590=>"011111110",
  16591=>"101011100",
  16592=>"000000100",
  16593=>"010111011",
  16594=>"110101110",
  16595=>"111011010",
  16596=>"000010100",
  16597=>"011010011",
  16598=>"110001110",
  16599=>"111100010",
  16600=>"000010010",
  16601=>"101000101",
  16602=>"000110010",
  16603=>"100111001",
  16604=>"001010000",
  16605=>"011111101",
  16606=>"001001110",
  16607=>"011001111",
  16608=>"111010110",
  16609=>"100000010",
  16610=>"010110000",
  16611=>"011111110",
  16612=>"010001100",
  16613=>"000111101",
  16614=>"101000000",
  16615=>"111010001",
  16616=>"101010001",
  16617=>"001000100",
  16618=>"000010000",
  16619=>"101101000",
  16620=>"001011110",
  16621=>"010001001",
  16622=>"001110010",
  16623=>"000111011",
  16624=>"011010100",
  16625=>"101011000",
  16626=>"010010001",
  16627=>"011000101",
  16628=>"000110101",
  16629=>"000011101",
  16630=>"110100010",
  16631=>"000010000",
  16632=>"000001011",
  16633=>"011110001",
  16634=>"111010100",
  16635=>"001110010",
  16636=>"000101001",
  16637=>"010101000",
  16638=>"100111111",
  16639=>"100001101",
  16640=>"010111111",
  16641=>"000110001",
  16642=>"111001111",
  16643=>"010101111",
  16644=>"100110101",
  16645=>"000001100",
  16646=>"011011011",
  16647=>"001111001",
  16648=>"001000100",
  16649=>"101000100",
  16650=>"111110000",
  16651=>"001111101",
  16652=>"000010010",
  16653=>"111100110",
  16654=>"111111011",
  16655=>"000110010",
  16656=>"111000101",
  16657=>"101011111",
  16658=>"100100100",
  16659=>"110101101",
  16660=>"000000100",
  16661=>"101000010",
  16662=>"000000010",
  16663=>"001011011",
  16664=>"110001001",
  16665=>"001011001",
  16666=>"111011011",
  16667=>"101100000",
  16668=>"100101010",
  16669=>"101110000",
  16670=>"000100000",
  16671=>"001110111",
  16672=>"111001101",
  16673=>"000100111",
  16674=>"001101111",
  16675=>"110100011",
  16676=>"011110110",
  16677=>"000000111",
  16678=>"111101000",
  16679=>"110011011",
  16680=>"010010101",
  16681=>"111111110",
  16682=>"110101001",
  16683=>"100001011",
  16684=>"101101000",
  16685=>"010001101",
  16686=>"110100111",
  16687=>"100101011",
  16688=>"011110100",
  16689=>"101101110",
  16690=>"011010100",
  16691=>"011101111",
  16692=>"010011101",
  16693=>"011100100",
  16694=>"111110110",
  16695=>"101001100",
  16696=>"000000101",
  16697=>"011001100",
  16698=>"100110101",
  16699=>"011101101",
  16700=>"011100101",
  16701=>"010110101",
  16702=>"111001011",
  16703=>"010111010",
  16704=>"100100111",
  16705=>"100011001",
  16706=>"000100101",
  16707=>"110101101",
  16708=>"110101000",
  16709=>"100101000",
  16710=>"000001110",
  16711=>"000100001",
  16712=>"101000100",
  16713=>"001101011",
  16714=>"101000001",
  16715=>"000101101",
  16716=>"101010100",
  16717=>"101100101",
  16718=>"111111111",
  16719=>"000010010",
  16720=>"110101110",
  16721=>"111110000",
  16722=>"101100010",
  16723=>"010101000",
  16724=>"010011100",
  16725=>"100000100",
  16726=>"010000111",
  16727=>"001001011",
  16728=>"000000001",
  16729=>"001000011",
  16730=>"100010001",
  16731=>"010101100",
  16732=>"011011010",
  16733=>"010101010",
  16734=>"111001101",
  16735=>"010100001",
  16736=>"110011011",
  16737=>"100010000",
  16738=>"100000101",
  16739=>"100001001",
  16740=>"010100000",
  16741=>"001111100",
  16742=>"000101011",
  16743=>"110001100",
  16744=>"000111001",
  16745=>"100010000",
  16746=>"100100100",
  16747=>"000111011",
  16748=>"111010011",
  16749=>"100001111",
  16750=>"000101110",
  16751=>"001000100",
  16752=>"010010001",
  16753=>"110100000",
  16754=>"010000000",
  16755=>"111111111",
  16756=>"011111010",
  16757=>"101101010",
  16758=>"111100101",
  16759=>"100000000",
  16760=>"010000001",
  16761=>"000010111",
  16762=>"011100011",
  16763=>"101101111",
  16764=>"001100000",
  16765=>"111111100",
  16766=>"110110000",
  16767=>"100010010",
  16768=>"011000001",
  16769=>"000010001",
  16770=>"111101110",
  16771=>"000000011",
  16772=>"101111111",
  16773=>"000011010",
  16774=>"110011011",
  16775=>"101110000",
  16776=>"010001000",
  16777=>"000111010",
  16778=>"000000001",
  16779=>"011001100",
  16780=>"110000010",
  16781=>"000110101",
  16782=>"010000000",
  16783=>"110111011",
  16784=>"001101101",
  16785=>"011000000",
  16786=>"101001000",
  16787=>"101110011",
  16788=>"001111011",
  16789=>"011000110",
  16790=>"110110001",
  16791=>"110011110",
  16792=>"010010111",
  16793=>"100001011",
  16794=>"101110110",
  16795=>"101011011",
  16796=>"010111011",
  16797=>"100011001",
  16798=>"100011001",
  16799=>"101010110",
  16800=>"111111000",
  16801=>"001101001",
  16802=>"001100110",
  16803=>"101001110",
  16804=>"101000100",
  16805=>"110010010",
  16806=>"110111111",
  16807=>"001000001",
  16808=>"000110001",
  16809=>"101010001",
  16810=>"100000000",
  16811=>"001010011",
  16812=>"010000010",
  16813=>"111001110",
  16814=>"010100101",
  16815=>"100110100",
  16816=>"000011000",
  16817=>"111001110",
  16818=>"110111000",
  16819=>"001101111",
  16820=>"100100100",
  16821=>"110101010",
  16822=>"110001000",
  16823=>"101110110",
  16824=>"110000000",
  16825=>"110000110",
  16826=>"010111010",
  16827=>"100101000",
  16828=>"010011110",
  16829=>"110001111",
  16830=>"000001000",
  16831=>"011110101",
  16832=>"101100100",
  16833=>"101100011",
  16834=>"000011001",
  16835=>"000010110",
  16836=>"010001001",
  16837=>"101001110",
  16838=>"101001111",
  16839=>"111000111",
  16840=>"001010101",
  16841=>"101111110",
  16842=>"100001101",
  16843=>"001111111",
  16844=>"010000100",
  16845=>"011101100",
  16846=>"100110010",
  16847=>"010111010",
  16848=>"010001011",
  16849=>"110111000",
  16850=>"110001000",
  16851=>"000011011",
  16852=>"011010110",
  16853=>"100000101",
  16854=>"001101000",
  16855=>"100100111",
  16856=>"001011100",
  16857=>"011101110",
  16858=>"111011010",
  16859=>"001010110",
  16860=>"100110000",
  16861=>"001011111",
  16862=>"101111111",
  16863=>"110111011",
  16864=>"010010000",
  16865=>"010100011",
  16866=>"011100011",
  16867=>"111000100",
  16868=>"110010000",
  16869=>"010110010",
  16870=>"110110010",
  16871=>"001000101",
  16872=>"000111101",
  16873=>"010111000",
  16874=>"000101011",
  16875=>"110111101",
  16876=>"100000101",
  16877=>"101010001",
  16878=>"010000010",
  16879=>"110101011",
  16880=>"001111100",
  16881=>"101110010",
  16882=>"100111111",
  16883=>"110011010",
  16884=>"011100001",
  16885=>"111101011",
  16886=>"100110000",
  16887=>"101011100",
  16888=>"010111011",
  16889=>"111011100",
  16890=>"111100101",
  16891=>"000001101",
  16892=>"011000100",
  16893=>"101010111",
  16894=>"000000001",
  16895=>"010101000",
  16896=>"101111111",
  16897=>"000100101",
  16898=>"110011000",
  16899=>"010100001",
  16900=>"010101010",
  16901=>"011000000",
  16902=>"111000111",
  16903=>"101111011",
  16904=>"011000101",
  16905=>"000100000",
  16906=>"110101000",
  16907=>"000001111",
  16908=>"001001011",
  16909=>"001100011",
  16910=>"001000000",
  16911=>"000101101",
  16912=>"111101001",
  16913=>"100010001",
  16914=>"010100001",
  16915=>"110100010",
  16916=>"110111001",
  16917=>"001111011",
  16918=>"111011011",
  16919=>"011111010",
  16920=>"000101000",
  16921=>"001111111",
  16922=>"001001110",
  16923=>"100100011",
  16924=>"101010011",
  16925=>"101111001",
  16926=>"001011010",
  16927=>"111010000",
  16928=>"011100001",
  16929=>"010010101",
  16930=>"100000000",
  16931=>"110111010",
  16932=>"010011010",
  16933=>"111100111",
  16934=>"010011101",
  16935=>"001010011",
  16936=>"010001010",
  16937=>"011101110",
  16938=>"101100001",
  16939=>"110000111",
  16940=>"101011001",
  16941=>"000110101",
  16942=>"111110010",
  16943=>"011000111",
  16944=>"110000000",
  16945=>"111110100",
  16946=>"100010101",
  16947=>"000000011",
  16948=>"101101011",
  16949=>"001110000",
  16950=>"011111011",
  16951=>"101011101",
  16952=>"110010010",
  16953=>"111100010",
  16954=>"100110010",
  16955=>"111110000",
  16956=>"001101011",
  16957=>"000001100",
  16958=>"001000001",
  16959=>"001100101",
  16960=>"011100011",
  16961=>"000011111",
  16962=>"111101100",
  16963=>"001110000",
  16964=>"010001000",
  16965=>"110010001",
  16966=>"101000111",
  16967=>"000111110",
  16968=>"000110001",
  16969=>"100000100",
  16970=>"100100111",
  16971=>"111101010",
  16972=>"001010010",
  16973=>"011100101",
  16974=>"011001100",
  16975=>"000100011",
  16976=>"010100000",
  16977=>"101001001",
  16978=>"010000000",
  16979=>"101011110",
  16980=>"100010001",
  16981=>"001011101",
  16982=>"010001110",
  16983=>"100101110",
  16984=>"011100100",
  16985=>"010000000",
  16986=>"100011001",
  16987=>"001111000",
  16988=>"000000111",
  16989=>"001101000",
  16990=>"010011000",
  16991=>"111111000",
  16992=>"000101100",
  16993=>"000010000",
  16994=>"100001101",
  16995=>"101110010",
  16996=>"001011111",
  16997=>"111110010",
  16998=>"010101111",
  16999=>"101001101",
  17000=>"110010010",
  17001=>"011100101",
  17002=>"111011101",
  17003=>"000110001",
  17004=>"010000011",
  17005=>"111001100",
  17006=>"000000000",
  17007=>"111010000",
  17008=>"101000000",
  17009=>"001101010",
  17010=>"011101100",
  17011=>"010011111",
  17012=>"000110001",
  17013=>"000110000",
  17014=>"001101101",
  17015=>"100000111",
  17016=>"000111001",
  17017=>"101011001",
  17018=>"110010010",
  17019=>"110110001",
  17020=>"110000001",
  17021=>"101111100",
  17022=>"100100000",
  17023=>"001001111",
  17024=>"100000010",
  17025=>"111100101",
  17026=>"001101111",
  17027=>"010101011",
  17028=>"111110000",
  17029=>"000100011",
  17030=>"000010001",
  17031=>"100100001",
  17032=>"110100010",
  17033=>"100010111",
  17034=>"101001100",
  17035=>"011001000",
  17036=>"100100110",
  17037=>"100000010",
  17038=>"111111110",
  17039=>"100101111",
  17040=>"010000100",
  17041=>"110011100",
  17042=>"100110010",
  17043=>"100011001",
  17044=>"110011010",
  17045=>"101011011",
  17046=>"110001001",
  17047=>"010111010",
  17048=>"100000100",
  17049=>"010001000",
  17050=>"011011010",
  17051=>"010111111",
  17052=>"111100101",
  17053=>"110010001",
  17054=>"100010100",
  17055=>"110001011",
  17056=>"011010111",
  17057=>"110111011",
  17058=>"101100011",
  17059=>"100010010",
  17060=>"101001111",
  17061=>"010111000",
  17062=>"100001110",
  17063=>"100111111",
  17064=>"101011100",
  17065=>"010111110",
  17066=>"101101001",
  17067=>"110110011",
  17068=>"010000000",
  17069=>"001110011",
  17070=>"011111000",
  17071=>"010010101",
  17072=>"011000101",
  17073=>"100110001",
  17074=>"010100000",
  17075=>"000010100",
  17076=>"110111001",
  17077=>"111011111",
  17078=>"110101100",
  17079=>"101000111",
  17080=>"101011111",
  17081=>"100000111",
  17082=>"011110010",
  17083=>"010100101",
  17084=>"001010000",
  17085=>"110001010",
  17086=>"010101100",
  17087=>"000110110",
  17088=>"100000001",
  17089=>"110000010",
  17090=>"011111010",
  17091=>"000001101",
  17092=>"101000101",
  17093=>"010011000",
  17094=>"111110100",
  17095=>"010111100",
  17096=>"111000010",
  17097=>"111000000",
  17098=>"000010101",
  17099=>"000011010",
  17100=>"001100111",
  17101=>"011111100",
  17102=>"111100100",
  17103=>"101110110",
  17104=>"001100001",
  17105=>"101101100",
  17106=>"100110110",
  17107=>"111010010",
  17108=>"100000001",
  17109=>"010010010",
  17110=>"011111010",
  17111=>"000011000",
  17112=>"111111110",
  17113=>"100111100",
  17114=>"010110010",
  17115=>"000000011",
  17116=>"001101100",
  17117=>"111010001",
  17118=>"101111001",
  17119=>"011010101",
  17120=>"010001110",
  17121=>"001010111",
  17122=>"101110010",
  17123=>"100101111",
  17124=>"110001100",
  17125=>"000100111",
  17126=>"010011010",
  17127=>"011010101",
  17128=>"010010110",
  17129=>"001001100",
  17130=>"000010001",
  17131=>"111001011",
  17132=>"100001100",
  17133=>"100100011",
  17134=>"111001011",
  17135=>"000001100",
  17136=>"101111011",
  17137=>"111000111",
  17138=>"000011101",
  17139=>"100110011",
  17140=>"100111011",
  17141=>"011000110",
  17142=>"010100011",
  17143=>"011011111",
  17144=>"001011010",
  17145=>"100111111",
  17146=>"000010100",
  17147=>"111001100",
  17148=>"100110101",
  17149=>"101100001",
  17150=>"101111101",
  17151=>"100010000",
  17152=>"101000010",
  17153=>"000010010",
  17154=>"010111110",
  17155=>"001110101",
  17156=>"011111101",
  17157=>"011010001",
  17158=>"011011011",
  17159=>"111010100",
  17160=>"100110011",
  17161=>"000001111",
  17162=>"101110110",
  17163=>"111101011",
  17164=>"010001000",
  17165=>"001010111",
  17166=>"001000101",
  17167=>"110010100",
  17168=>"011000000",
  17169=>"001111101",
  17170=>"101011100",
  17171=>"011101001",
  17172=>"100111110",
  17173=>"000000100",
  17174=>"001101010",
  17175=>"001010011",
  17176=>"111010010",
  17177=>"111000100",
  17178=>"000100100",
  17179=>"110111110",
  17180=>"111101011",
  17181=>"110110011",
  17182=>"000101100",
  17183=>"111000101",
  17184=>"110101101",
  17185=>"000111101",
  17186=>"110101010",
  17187=>"000101010",
  17188=>"100001100",
  17189=>"101110100",
  17190=>"100101101",
  17191=>"100101011",
  17192=>"100000111",
  17193=>"000110100",
  17194=>"001111011",
  17195=>"111111111",
  17196=>"001111101",
  17197=>"000100000",
  17198=>"001000100",
  17199=>"101100000",
  17200=>"011100110",
  17201=>"000010110",
  17202=>"010111101",
  17203=>"101111101",
  17204=>"100101010",
  17205=>"110111000",
  17206=>"101101011",
  17207=>"101100001",
  17208=>"111100110",
  17209=>"111001110",
  17210=>"100001011",
  17211=>"011000100",
  17212=>"000110101",
  17213=>"111101101",
  17214=>"100000100",
  17215=>"001010000",
  17216=>"110111011",
  17217=>"100011110",
  17218=>"111011000",
  17219=>"110010001",
  17220=>"000001011",
  17221=>"101101111",
  17222=>"011100111",
  17223=>"000000010",
  17224=>"000010111",
  17225=>"000110111",
  17226=>"110111110",
  17227=>"101010011",
  17228=>"101110111",
  17229=>"010110001",
  17230=>"111111101",
  17231=>"110101111",
  17232=>"110100011",
  17233=>"101011010",
  17234=>"011100000",
  17235=>"111000000",
  17236=>"010000010",
  17237=>"000101000",
  17238=>"101000111",
  17239=>"000111010",
  17240=>"100000111",
  17241=>"000101101",
  17242=>"001011011",
  17243=>"111111100",
  17244=>"110010011",
  17245=>"100110110",
  17246=>"001111001",
  17247=>"000000010",
  17248=>"101000010",
  17249=>"110110110",
  17250=>"000001000",
  17251=>"111101101",
  17252=>"001000000",
  17253=>"101110000",
  17254=>"101110110",
  17255=>"001010010",
  17256=>"000010000",
  17257=>"011101000",
  17258=>"001110001",
  17259=>"001010000",
  17260=>"111010101",
  17261=>"011101111",
  17262=>"001011100",
  17263=>"011011111",
  17264=>"011001111",
  17265=>"011110111",
  17266=>"111011111",
  17267=>"111010000",
  17268=>"100101000",
  17269=>"001111110",
  17270=>"100100000",
  17271=>"000000011",
  17272=>"000100001",
  17273=>"001100010",
  17274=>"010111101",
  17275=>"111011010",
  17276=>"010000000",
  17277=>"010011101",
  17278=>"010011111",
  17279=>"000100110",
  17280=>"111110100",
  17281=>"100011110",
  17282=>"000010000",
  17283=>"101111100",
  17284=>"110101011",
  17285=>"110111010",
  17286=>"100110110",
  17287=>"000111010",
  17288=>"000110010",
  17289=>"100000100",
  17290=>"000010110",
  17291=>"001110010",
  17292=>"110110011",
  17293=>"110111000",
  17294=>"000101100",
  17295=>"100111111",
  17296=>"111000001",
  17297=>"101000011",
  17298=>"011010000",
  17299=>"010000111",
  17300=>"110100001",
  17301=>"011110001",
  17302=>"110000001",
  17303=>"001101011",
  17304=>"000000101",
  17305=>"100100110",
  17306=>"000000100",
  17307=>"000111010",
  17308=>"010001111",
  17309=>"111001100",
  17310=>"100011111",
  17311=>"000011011",
  17312=>"011001111",
  17313=>"100101111",
  17314=>"100001011",
  17315=>"001000000",
  17316=>"100110111",
  17317=>"110000101",
  17318=>"111001101",
  17319=>"010101110",
  17320=>"010101011",
  17321=>"100110010",
  17322=>"111110101",
  17323=>"001100111",
  17324=>"000001010",
  17325=>"010110000",
  17326=>"111001100",
  17327=>"111000111",
  17328=>"010100001",
  17329=>"010011110",
  17330=>"010100011",
  17331=>"101011001",
  17332=>"100010011",
  17333=>"111110110",
  17334=>"011110111",
  17335=>"000101010",
  17336=>"000001111",
  17337=>"010010001",
  17338=>"111110110",
  17339=>"110000111",
  17340=>"010011001",
  17341=>"111000001",
  17342=>"011110101",
  17343=>"000110011",
  17344=>"000101010",
  17345=>"110100010",
  17346=>"011001100",
  17347=>"110111011",
  17348=>"110000100",
  17349=>"000110001",
  17350=>"101101110",
  17351=>"111111000",
  17352=>"011100000",
  17353=>"000111111",
  17354=>"111110100",
  17355=>"100110000",
  17356=>"001110011",
  17357=>"100000001",
  17358=>"010110101",
  17359=>"000010011",
  17360=>"010111000",
  17361=>"000010001",
  17362=>"101110101",
  17363=>"000010100",
  17364=>"111110100",
  17365=>"111110011",
  17366=>"011010101",
  17367=>"011011010",
  17368=>"000000110",
  17369=>"101111001",
  17370=>"011111101",
  17371=>"101010100",
  17372=>"010011000",
  17373=>"111000000",
  17374=>"111010010",
  17375=>"000100010",
  17376=>"100000110",
  17377=>"010110101",
  17378=>"100111101",
  17379=>"110110010",
  17380=>"110100010",
  17381=>"000011100",
  17382=>"001000101",
  17383=>"101010111",
  17384=>"100011101",
  17385=>"000111011",
  17386=>"111000010",
  17387=>"110010110",
  17388=>"001001010",
  17389=>"000111000",
  17390=>"100111110",
  17391=>"001101000",
  17392=>"010110111",
  17393=>"101010011",
  17394=>"011000110",
  17395=>"110010001",
  17396=>"000000000",
  17397=>"011011010",
  17398=>"110110010",
  17399=>"001000010",
  17400=>"110100101",
  17401=>"111011111",
  17402=>"111101000",
  17403=>"111111001",
  17404=>"000010001",
  17405=>"011101101",
  17406=>"000111110",
  17407=>"111100100",
  17408=>"000111110",
  17409=>"110101101",
  17410=>"100010100",
  17411=>"000000101",
  17412=>"111110000",
  17413=>"011111010",
  17414=>"111110001",
  17415=>"010001100",
  17416=>"011111010",
  17417=>"111000110",
  17418=>"000101010",
  17419=>"111010111",
  17420=>"010100000",
  17421=>"101100111",
  17422=>"110000110",
  17423=>"000000010",
  17424=>"101100101",
  17425=>"101010111",
  17426=>"110111111",
  17427=>"101111010",
  17428=>"100100000",
  17429=>"110011000",
  17430=>"001001011",
  17431=>"010001001",
  17432=>"110111111",
  17433=>"000110111",
  17434=>"001001101",
  17435=>"001011011",
  17436=>"010101100",
  17437=>"010010000",
  17438=>"110011110",
  17439=>"000101110",
  17440=>"110111101",
  17441=>"111000000",
  17442=>"000000001",
  17443=>"000000001",
  17444=>"010111110",
  17445=>"100000011",
  17446=>"110010111",
  17447=>"101111000",
  17448=>"011010111",
  17449=>"000010100",
  17450=>"010110111",
  17451=>"011111010",
  17452=>"100000000",
  17453=>"110011011",
  17454=>"000111101",
  17455=>"010100100",
  17456=>"000001010",
  17457=>"010101000",
  17458=>"110000000",
  17459=>"011110001",
  17460=>"100110011",
  17461=>"011111100",
  17462=>"010011001",
  17463=>"010001101",
  17464=>"010100110",
  17465=>"010010000",
  17466=>"001010101",
  17467=>"111001111",
  17468=>"011010111",
  17469=>"111100101",
  17470=>"101001000",
  17471=>"101100011",
  17472=>"011000111",
  17473=>"011111101",
  17474=>"000100000",
  17475=>"101110011",
  17476=>"110010111",
  17477=>"000101110",
  17478=>"101000010",
  17479=>"101011011",
  17480=>"100110101",
  17481=>"100100101",
  17482=>"001001001",
  17483=>"111000111",
  17484=>"101001100",
  17485=>"010111100",
  17486=>"101000101",
  17487=>"110010010",
  17488=>"000010100",
  17489=>"111101011",
  17490=>"000001100",
  17491=>"111010001",
  17492=>"110100011",
  17493=>"011000000",
  17494=>"010111010",
  17495=>"001010011",
  17496=>"010101100",
  17497=>"010100111",
  17498=>"100010110",
  17499=>"011000101",
  17500=>"100101000",
  17501=>"011001000",
  17502=>"100000011",
  17503=>"001011010",
  17504=>"000010000",
  17505=>"011111011",
  17506=>"011100111",
  17507=>"110101011",
  17508=>"000110001",
  17509=>"100110100",
  17510=>"001111010",
  17511=>"010100011",
  17512=>"011000001",
  17513=>"110100000",
  17514=>"001001101",
  17515=>"100010011",
  17516=>"001001001",
  17517=>"111110001",
  17518=>"010111010",
  17519=>"100011001",
  17520=>"100100000",
  17521=>"110110111",
  17522=>"011100110",
  17523=>"010111100",
  17524=>"110011101",
  17525=>"101101101",
  17526=>"001010011",
  17527=>"111110010",
  17528=>"101101000",
  17529=>"110110011",
  17530=>"101010010",
  17531=>"010111011",
  17532=>"111011111",
  17533=>"100101011",
  17534=>"000001111",
  17535=>"010010110",
  17536=>"111100110",
  17537=>"101001011",
  17538=>"001010011",
  17539=>"011100110",
  17540=>"110001110",
  17541=>"001000011",
  17542=>"111111001",
  17543=>"110010011",
  17544=>"010000111",
  17545=>"000100000",
  17546=>"011001000",
  17547=>"111000101",
  17548=>"101111000",
  17549=>"011001000",
  17550=>"111101101",
  17551=>"101000010",
  17552=>"011110010",
  17553=>"111000111",
  17554=>"001001000",
  17555=>"111111101",
  17556=>"111100001",
  17557=>"010010011",
  17558=>"000010011",
  17559=>"100100111",
  17560=>"111001111",
  17561=>"110001110",
  17562=>"000000001",
  17563=>"100010010",
  17564=>"100110010",
  17565=>"101000001",
  17566=>"100000010",
  17567=>"001101011",
  17568=>"011011011",
  17569=>"111000110",
  17570=>"110100000",
  17571=>"100001110",
  17572=>"110001010",
  17573=>"111001101",
  17574=>"010001001",
  17575=>"000100010",
  17576=>"100011101",
  17577=>"111110111",
  17578=>"010001101",
  17579=>"101001101",
  17580=>"011110100",
  17581=>"101011011",
  17582=>"010110010",
  17583=>"101000111",
  17584=>"010101110",
  17585=>"000001001",
  17586=>"111111101",
  17587=>"001100001",
  17588=>"101010011",
  17589=>"111101011",
  17590=>"100100001",
  17591=>"110000011",
  17592=>"010000010",
  17593=>"001000011",
  17594=>"011000001",
  17595=>"101100011",
  17596=>"001001001",
  17597=>"101110000",
  17598=>"111111011",
  17599=>"011101000",
  17600=>"000100001",
  17601=>"010101011",
  17602=>"001011110",
  17603=>"100100110",
  17604=>"101110011",
  17605=>"000000100",
  17606=>"101011001",
  17607=>"101001001",
  17608=>"000100011",
  17609=>"100000100",
  17610=>"100011001",
  17611=>"001010010",
  17612=>"100100000",
  17613=>"100110010",
  17614=>"111100000",
  17615=>"011100100",
  17616=>"000111011",
  17617=>"011101010",
  17618=>"101010001",
  17619=>"001001111",
  17620=>"011101011",
  17621=>"001001000",
  17622=>"011111110",
  17623=>"001100010",
  17624=>"100100000",
  17625=>"100001100",
  17626=>"110000111",
  17627=>"001100001",
  17628=>"011101100",
  17629=>"001100101",
  17630=>"101100011",
  17631=>"001101100",
  17632=>"011000000",
  17633=>"100010001",
  17634=>"110011011",
  17635=>"001011000",
  17636=>"111011100",
  17637=>"001100011",
  17638=>"111110110",
  17639=>"111010111",
  17640=>"001110001",
  17641=>"010010101",
  17642=>"001001100",
  17643=>"010110100",
  17644=>"000000001",
  17645=>"100000011",
  17646=>"011010110",
  17647=>"000010000",
  17648=>"011101000",
  17649=>"111000111",
  17650=>"011000110",
  17651=>"100101001",
  17652=>"100000110",
  17653=>"100100110",
  17654=>"100100110",
  17655=>"011111110",
  17656=>"011011110",
  17657=>"111000110",
  17658=>"110011111",
  17659=>"011110101",
  17660=>"010010111",
  17661=>"111110000",
  17662=>"001100001",
  17663=>"101100110",
  17664=>"011001000",
  17665=>"101111100",
  17666=>"111111100",
  17667=>"010111111",
  17668=>"001100001",
  17669=>"110011101",
  17670=>"011111101",
  17671=>"110010100",
  17672=>"010110111",
  17673=>"100011001",
  17674=>"011111110",
  17675=>"110000101",
  17676=>"100010001",
  17677=>"000010001",
  17678=>"111010100",
  17679=>"101011111",
  17680=>"011000001",
  17681=>"001101001",
  17682=>"101111000",
  17683=>"111000100",
  17684=>"001100111",
  17685=>"000100111",
  17686=>"110000000",
  17687=>"011111010",
  17688=>"101001100",
  17689=>"001010000",
  17690=>"101110010",
  17691=>"001111000",
  17692=>"011101011",
  17693=>"111100000",
  17694=>"111000011",
  17695=>"000011001",
  17696=>"100100111",
  17697=>"100001001",
  17698=>"011111001",
  17699=>"101101011",
  17700=>"101000100",
  17701=>"100001101",
  17702=>"101001001",
  17703=>"101011001",
  17704=>"000110010",
  17705=>"011101110",
  17706=>"010011100",
  17707=>"000000000",
  17708=>"111011100",
  17709=>"111101000",
  17710=>"111111010",
  17711=>"101110011",
  17712=>"011001101",
  17713=>"100110011",
  17714=>"010110000",
  17715=>"010001000",
  17716=>"101011001",
  17717=>"111001010",
  17718=>"110010010",
  17719=>"001001100",
  17720=>"000000010",
  17721=>"101101001",
  17722=>"110111001",
  17723=>"001110100",
  17724=>"010001111",
  17725=>"001110010",
  17726=>"110100000",
  17727=>"000101111",
  17728=>"111101011",
  17729=>"110110000",
  17730=>"101111000",
  17731=>"000011111",
  17732=>"111011100",
  17733=>"101010111",
  17734=>"110010001",
  17735=>"011111111",
  17736=>"010010110",
  17737=>"001001001",
  17738=>"011011110",
  17739=>"000001010",
  17740=>"111010111",
  17741=>"100100011",
  17742=>"101001011",
  17743=>"111010011",
  17744=>"011001110",
  17745=>"001000100",
  17746=>"100100001",
  17747=>"000011100",
  17748=>"010100011",
  17749=>"010001101",
  17750=>"001001000",
  17751=>"001010000",
  17752=>"110100011",
  17753=>"000111110",
  17754=>"111110001",
  17755=>"010100001",
  17756=>"010110011",
  17757=>"011111011",
  17758=>"111000000",
  17759=>"000100001",
  17760=>"001010001",
  17761=>"111011110",
  17762=>"000111010",
  17763=>"000000011",
  17764=>"010010010",
  17765=>"110111000",
  17766=>"101111111",
  17767=>"111100111",
  17768=>"010111001",
  17769=>"000110111",
  17770=>"001001000",
  17771=>"001011110",
  17772=>"101010010",
  17773=>"011010000",
  17774=>"100011000",
  17775=>"110001111",
  17776=>"000000011",
  17777=>"111110010",
  17778=>"111111010",
  17779=>"010110101",
  17780=>"110001111",
  17781=>"000010011",
  17782=>"010011111",
  17783=>"101010000",
  17784=>"101000110",
  17785=>"111101011",
  17786=>"011100101",
  17787=>"100000100",
  17788=>"000100010",
  17789=>"110101010",
  17790=>"000001011",
  17791=>"000110101",
  17792=>"010111111",
  17793=>"101101000",
  17794=>"111101110",
  17795=>"111011101",
  17796=>"011111010",
  17797=>"111110111",
  17798=>"100001111",
  17799=>"001001011",
  17800=>"010010111",
  17801=>"010001100",
  17802=>"110000001",
  17803=>"000100000",
  17804=>"000001101",
  17805=>"101110100",
  17806=>"001100000",
  17807=>"110010101",
  17808=>"110101000",
  17809=>"001101101",
  17810=>"101000100",
  17811=>"110100011",
  17812=>"101011110",
  17813=>"000110001",
  17814=>"111110011",
  17815=>"000100001",
  17816=>"101111101",
  17817=>"010011001",
  17818=>"000111010",
  17819=>"111111010",
  17820=>"101011000",
  17821=>"000111010",
  17822=>"011000111",
  17823=>"110111101",
  17824=>"100111010",
  17825=>"111011000",
  17826=>"011001001",
  17827=>"011110011",
  17828=>"011010000",
  17829=>"110110111",
  17830=>"110111000",
  17831=>"110010100",
  17832=>"000001110",
  17833=>"110111100",
  17834=>"001011011",
  17835=>"000110110",
  17836=>"110100001",
  17837=>"100010111",
  17838=>"011000011",
  17839=>"011100000",
  17840=>"100100100",
  17841=>"110000001",
  17842=>"100010000",
  17843=>"011111101",
  17844=>"110110010",
  17845=>"100110001",
  17846=>"000110000",
  17847=>"100110010",
  17848=>"111111011",
  17849=>"001101111",
  17850=>"011010011",
  17851=>"100011001",
  17852=>"111101111",
  17853=>"000110110",
  17854=>"111110111",
  17855=>"100001001",
  17856=>"111010011",
  17857=>"101100101",
  17858=>"100010100",
  17859=>"111101011",
  17860=>"000001111",
  17861=>"010111101",
  17862=>"001010010",
  17863=>"011000000",
  17864=>"001101100",
  17865=>"010001101",
  17866=>"100001000",
  17867=>"010010001",
  17868=>"110011111",
  17869=>"000001000",
  17870=>"001010100",
  17871=>"000001000",
  17872=>"110111100",
  17873=>"011000010",
  17874=>"100111011",
  17875=>"000111000",
  17876=>"101011100",
  17877=>"001110010",
  17878=>"011111010",
  17879=>"111011011",
  17880=>"011001011",
  17881=>"101100001",
  17882=>"101110101",
  17883=>"011010100",
  17884=>"101110010",
  17885=>"110000100",
  17886=>"011100000",
  17887=>"101101100",
  17888=>"110101010",
  17889=>"111110110",
  17890=>"111001000",
  17891=>"110111000",
  17892=>"001000011",
  17893=>"000100101",
  17894=>"101111010",
  17895=>"110011001",
  17896=>"011100000",
  17897=>"111001000",
  17898=>"100101001",
  17899=>"011111101",
  17900=>"000110101",
  17901=>"000101010",
  17902=>"111001010",
  17903=>"110001101",
  17904=>"111110110",
  17905=>"000001101",
  17906=>"111100011",
  17907=>"000000001",
  17908=>"100101011",
  17909=>"111110111",
  17910=>"011010101",
  17911=>"111001100",
  17912=>"000001000",
  17913=>"100110000",
  17914=>"110011010",
  17915=>"011011010",
  17916=>"001101101",
  17917=>"110101110",
  17918=>"110111001",
  17919=>"000001110",
  17920=>"110101000",
  17921=>"001111110",
  17922=>"101010100",
  17923=>"000010111",
  17924=>"011100110",
  17925=>"101010101",
  17926=>"011001111",
  17927=>"110101011",
  17928=>"010011001",
  17929=>"100001000",
  17930=>"000101110",
  17931=>"111001110",
  17932=>"101001000",
  17933=>"001110000",
  17934=>"001011000",
  17935=>"100111000",
  17936=>"010001101",
  17937=>"000001011",
  17938=>"111011000",
  17939=>"010110010",
  17940=>"010010001",
  17941=>"100001110",
  17942=>"110011110",
  17943=>"100010010",
  17944=>"100101110",
  17945=>"101101001",
  17946=>"111010011",
  17947=>"011010111",
  17948=>"110111101",
  17949=>"001101101",
  17950=>"001010100",
  17951=>"111100110",
  17952=>"101011011",
  17953=>"111110000",
  17954=>"011011111",
  17955=>"000011000",
  17956=>"100111111",
  17957=>"110001001",
  17958=>"100000010",
  17959=>"010010100",
  17960=>"111001111",
  17961=>"100000111",
  17962=>"101100010",
  17963=>"110000101",
  17964=>"101010000",
  17965=>"101111111",
  17966=>"011100011",
  17967=>"000001101",
  17968=>"011001110",
  17969=>"111001010",
  17970=>"010001001",
  17971=>"010101011",
  17972=>"000110100",
  17973=>"001011111",
  17974=>"101100101",
  17975=>"010001010",
  17976=>"010101011",
  17977=>"111011000",
  17978=>"111010010",
  17979=>"110000100",
  17980=>"110111110",
  17981=>"111000101",
  17982=>"011101011",
  17983=>"000110100",
  17984=>"001111001",
  17985=>"000000010",
  17986=>"100100010",
  17987=>"000111001",
  17988=>"000010001",
  17989=>"001111110",
  17990=>"001000011",
  17991=>"001100100",
  17992=>"010101110",
  17993=>"111100010",
  17994=>"110001001",
  17995=>"111110010",
  17996=>"110001001",
  17997=>"001100001",
  17998=>"101111001",
  17999=>"011110111",
  18000=>"011000001",
  18001=>"001000000",
  18002=>"000110001",
  18003=>"110000010",
  18004=>"010001000",
  18005=>"011010101",
  18006=>"110110111",
  18007=>"110000110",
  18008=>"111100000",
  18009=>"001001110",
  18010=>"010100010",
  18011=>"001111110",
  18012=>"001111011",
  18013=>"101100100",
  18014=>"101010000",
  18015=>"111100000",
  18016=>"010101101",
  18017=>"111110111",
  18018=>"010010010",
  18019=>"001100110",
  18020=>"011000000",
  18021=>"001101000",
  18022=>"010000100",
  18023=>"010101010",
  18024=>"100011100",
  18025=>"111111011",
  18026=>"010110110",
  18027=>"011000101",
  18028=>"100100001",
  18029=>"011000011",
  18030=>"000001010",
  18031=>"111100001",
  18032=>"011101001",
  18033=>"100011100",
  18034=>"110000110",
  18035=>"001101111",
  18036=>"010001010",
  18037=>"100001000",
  18038=>"111011110",
  18039=>"100110001",
  18040=>"001000001",
  18041=>"011011011",
  18042=>"011000110",
  18043=>"000100111",
  18044=>"010000001",
  18045=>"000101110",
  18046=>"100001010",
  18047=>"001101111",
  18048=>"011100010",
  18049=>"110010010",
  18050=>"001000011",
  18051=>"110001110",
  18052=>"110011010",
  18053=>"100100000",
  18054=>"110000010",
  18055=>"010001111",
  18056=>"011101101",
  18057=>"010111110",
  18058=>"010111111",
  18059=>"100001100",
  18060=>"111111111",
  18061=>"010110101",
  18062=>"111001110",
  18063=>"000110000",
  18064=>"111100000",
  18065=>"011001110",
  18066=>"101111001",
  18067=>"011111000",
  18068=>"110100001",
  18069=>"010010100",
  18070=>"111001110",
  18071=>"101111111",
  18072=>"000110101",
  18073=>"111111111",
  18074=>"010000000",
  18075=>"111111110",
  18076=>"111000010",
  18077=>"101000011",
  18078=>"110110110",
  18079=>"001000110",
  18080=>"000010001",
  18081=>"111101110",
  18082=>"100110000",
  18083=>"110010001",
  18084=>"001011001",
  18085=>"101110010",
  18086=>"000111011",
  18087=>"001101100",
  18088=>"000000101",
  18089=>"000000100",
  18090=>"100000001",
  18091=>"010101010",
  18092=>"000101011",
  18093=>"010100110",
  18094=>"000000101",
  18095=>"000101100",
  18096=>"010001011",
  18097=>"011111010",
  18098=>"101001110",
  18099=>"001111000",
  18100=>"101110010",
  18101=>"001010111",
  18102=>"100001010",
  18103=>"111100100",
  18104=>"011010010",
  18105=>"011101000",
  18106=>"100000101",
  18107=>"100001000",
  18108=>"000001110",
  18109=>"111101101",
  18110=>"100101111",
  18111=>"001111010",
  18112=>"011111001",
  18113=>"100011101",
  18114=>"000111101",
  18115=>"000101010",
  18116=>"010001111",
  18117=>"110010101",
  18118=>"011100111",
  18119=>"111000111",
  18120=>"000100101",
  18121=>"000110100",
  18122=>"001101100",
  18123=>"010101111",
  18124=>"110110110",
  18125=>"100000000",
  18126=>"101001001",
  18127=>"111110110",
  18128=>"000001100",
  18129=>"010110011",
  18130=>"101011101",
  18131=>"000111110",
  18132=>"001000111",
  18133=>"111001011",
  18134=>"100010111",
  18135=>"011011100",
  18136=>"011111100",
  18137=>"101011110",
  18138=>"100001001",
  18139=>"000011011",
  18140=>"101110010",
  18141=>"001100011",
  18142=>"001101000",
  18143=>"000101010",
  18144=>"111111111",
  18145=>"000100001",
  18146=>"110010110",
  18147=>"000111010",
  18148=>"101100101",
  18149=>"000000000",
  18150=>"001110011",
  18151=>"110001010",
  18152=>"100101001",
  18153=>"110110111",
  18154=>"100100101",
  18155=>"110000011",
  18156=>"100111100",
  18157=>"000101011",
  18158=>"010101000",
  18159=>"110010100",
  18160=>"111110100",
  18161=>"000101000",
  18162=>"111001010",
  18163=>"011110111",
  18164=>"100001000",
  18165=>"011010111",
  18166=>"011111011",
  18167=>"001000010",
  18168=>"001000010",
  18169=>"011010000",
  18170=>"000011111",
  18171=>"100011001",
  18172=>"100111110",
  18173=>"001011110",
  18174=>"010111010",
  18175=>"100101001",
  18176=>"011111001",
  18177=>"011100100",
  18178=>"001000000",
  18179=>"010100000",
  18180=>"000010110",
  18181=>"100001010",
  18182=>"000110010",
  18183=>"010111111",
  18184=>"000011100",
  18185=>"100001000",
  18186=>"101101010",
  18187=>"000111001",
  18188=>"000010001",
  18189=>"001000011",
  18190=>"001000001",
  18191=>"111110100",
  18192=>"000011011",
  18193=>"001101000",
  18194=>"101110011",
  18195=>"111110111",
  18196=>"000001111",
  18197=>"111001111",
  18198=>"100011001",
  18199=>"000001110",
  18200=>"011111010",
  18201=>"001111001",
  18202=>"011101000",
  18203=>"000111000",
  18204=>"101100101",
  18205=>"111011011",
  18206=>"010000111",
  18207=>"100010111",
  18208=>"010101110",
  18209=>"011101011",
  18210=>"000000100",
  18211=>"100001010",
  18212=>"011011111",
  18213=>"010001001",
  18214=>"010110101",
  18215=>"000110111",
  18216=>"011001101",
  18217=>"010010000",
  18218=>"100111011",
  18219=>"000010011",
  18220=>"101000000",
  18221=>"111100101",
  18222=>"001111100",
  18223=>"100000011",
  18224=>"110001011",
  18225=>"101010111",
  18226=>"000110100",
  18227=>"010100010",
  18228=>"100100000",
  18229=>"111111110",
  18230=>"011100101",
  18231=>"100111101",
  18232=>"111110000",
  18233=>"000101100",
  18234=>"010110011",
  18235=>"001011010",
  18236=>"000001100",
  18237=>"011101101",
  18238=>"000010100",
  18239=>"000010101",
  18240=>"110001110",
  18241=>"010011100",
  18242=>"011100111",
  18243=>"000000001",
  18244=>"010010100",
  18245=>"010100110",
  18246=>"111100111",
  18247=>"001100111",
  18248=>"110101110",
  18249=>"101011000",
  18250=>"101000000",
  18251=>"001000111",
  18252=>"100100101",
  18253=>"110100100",
  18254=>"111000110",
  18255=>"011010100",
  18256=>"111110110",
  18257=>"000101000",
  18258=>"010101100",
  18259=>"010010011",
  18260=>"110011001",
  18261=>"000111110",
  18262=>"100010100",
  18263=>"111100111",
  18264=>"000111101",
  18265=>"000001100",
  18266=>"010010001",
  18267=>"101011000",
  18268=>"101111111",
  18269=>"011101011",
  18270=>"111100111",
  18271=>"100110001",
  18272=>"011100100",
  18273=>"110101111",
  18274=>"100100010",
  18275=>"100111010",
  18276=>"100011011",
  18277=>"010111111",
  18278=>"101000110",
  18279=>"101010111",
  18280=>"011011000",
  18281=>"001000101",
  18282=>"000010100",
  18283=>"111101101",
  18284=>"010010010",
  18285=>"110000100",
  18286=>"100100000",
  18287=>"111010011",
  18288=>"110000010",
  18289=>"111001010",
  18290=>"110111011",
  18291=>"110001111",
  18292=>"000000110",
  18293=>"110110110",
  18294=>"110001010",
  18295=>"001100011",
  18296=>"000001000",
  18297=>"101001011",
  18298=>"000011010",
  18299=>"010011000",
  18300=>"000001000",
  18301=>"000001110",
  18302=>"111100000",
  18303=>"100101010",
  18304=>"101101000",
  18305=>"101110110",
  18306=>"000111011",
  18307=>"111010110",
  18308=>"111101100",
  18309=>"111000100",
  18310=>"101101000",
  18311=>"100011010",
  18312=>"100000011",
  18313=>"001000011",
  18314=>"111000000",
  18315=>"001000011",
  18316=>"110001100",
  18317=>"110011011",
  18318=>"011010010",
  18319=>"001111111",
  18320=>"110111110",
  18321=>"111111101",
  18322=>"100001011",
  18323=>"111100110",
  18324=>"111010100",
  18325=>"101001110",
  18326=>"010011101",
  18327=>"001010010",
  18328=>"111000111",
  18329=>"000100111",
  18330=>"110110000",
  18331=>"101111101",
  18332=>"010100010",
  18333=>"101100110",
  18334=>"011011011",
  18335=>"101100011",
  18336=>"101110010",
  18337=>"100010101",
  18338=>"000001111",
  18339=>"100110011",
  18340=>"100001000",
  18341=>"101001110",
  18342=>"111011001",
  18343=>"000001110",
  18344=>"001001100",
  18345=>"101111110",
  18346=>"110001010",
  18347=>"010101111",
  18348=>"010110100",
  18349=>"001011000",
  18350=>"110010011",
  18351=>"010100010",
  18352=>"000001001",
  18353=>"000001111",
  18354=>"000100100",
  18355=>"001010110",
  18356=>"101001110",
  18357=>"101101100",
  18358=>"010010001",
  18359=>"111110011",
  18360=>"110000010",
  18361=>"110000000",
  18362=>"100100101",
  18363=>"101000001",
  18364=>"101101011",
  18365=>"010010111",
  18366=>"101000000",
  18367=>"100011110",
  18368=>"111000010",
  18369=>"111100110",
  18370=>"010110000",
  18371=>"100011110",
  18372=>"010001111",
  18373=>"111001110",
  18374=>"011110101",
  18375=>"011111111",
  18376=>"010011001",
  18377=>"011011001",
  18378=>"011000110",
  18379=>"111111100",
  18380=>"000000110",
  18381=>"110000101",
  18382=>"001010011",
  18383=>"000111011",
  18384=>"101111001",
  18385=>"101011111",
  18386=>"111111100",
  18387=>"101011111",
  18388=>"100010101",
  18389=>"011111111",
  18390=>"110101001",
  18391=>"000010000",
  18392=>"000010100",
  18393=>"111011110",
  18394=>"010111111",
  18395=>"010000110",
  18396=>"001001101",
  18397=>"010111001",
  18398=>"001101001",
  18399=>"101100000",
  18400=>"000010001",
  18401=>"010010111",
  18402=>"011001100",
  18403=>"101010111",
  18404=>"010001000",
  18405=>"110101000",
  18406=>"101111010",
  18407=>"001001010",
  18408=>"010111111",
  18409=>"111001111",
  18410=>"001110110",
  18411=>"000000100",
  18412=>"001010010",
  18413=>"001011101",
  18414=>"110101100",
  18415=>"000000110",
  18416=>"010111100",
  18417=>"110011111",
  18418=>"000101111",
  18419=>"101010010",
  18420=>"100110000",
  18421=>"011111100",
  18422=>"111011001",
  18423=>"000000010",
  18424=>"110111010",
  18425=>"001111001",
  18426=>"001110110",
  18427=>"000011011",
  18428=>"011101001",
  18429=>"000000000",
  18430=>"001101101",
  18431=>"110001101",
  18432=>"110000001",
  18433=>"000010111",
  18434=>"101010001",
  18435=>"000111000",
  18436=>"010000101",
  18437=>"110001001",
  18438=>"011110110",
  18439=>"101101001",
  18440=>"010010101",
  18441=>"100010011",
  18442=>"000011010",
  18443=>"110000101",
  18444=>"001101001",
  18445=>"010110111",
  18446=>"010000100",
  18447=>"100001101",
  18448=>"101111110",
  18449=>"111100000",
  18450=>"111011010",
  18451=>"110011000",
  18452=>"111001001",
  18453=>"000010111",
  18454=>"100010011",
  18455=>"000010011",
  18456=>"011000000",
  18457=>"001100001",
  18458=>"010011100",
  18459=>"010110111",
  18460=>"110100111",
  18461=>"101110010",
  18462=>"111010011",
  18463=>"110000000",
  18464=>"110011010",
  18465=>"111000100",
  18466=>"011000100",
  18467=>"100010101",
  18468=>"100001100",
  18469=>"011100001",
  18470=>"111110101",
  18471=>"010010011",
  18472=>"011100110",
  18473=>"001111101",
  18474=>"111111110",
  18475=>"000111101",
  18476=>"011111111",
  18477=>"100101010",
  18478=>"000010011",
  18479=>"001111010",
  18480=>"000000000",
  18481=>"000101110",
  18482=>"000101100",
  18483=>"011100100",
  18484=>"001000001",
  18485=>"000001000",
  18486=>"011010011",
  18487=>"011100100",
  18488=>"110111101",
  18489=>"011110010",
  18490=>"000011000",
  18491=>"000000101",
  18492=>"000101010",
  18493=>"110000100",
  18494=>"001011001",
  18495=>"010010011",
  18496=>"001100100",
  18497=>"010001101",
  18498=>"101010100",
  18499=>"110010100",
  18500=>"101001110",
  18501=>"110010001",
  18502=>"111011000",
  18503=>"011001000",
  18504=>"100110101",
  18505=>"011001100",
  18506=>"000111000",
  18507=>"001110011",
  18508=>"010011111",
  18509=>"010101100",
  18510=>"010111010",
  18511=>"010011111",
  18512=>"011001001",
  18513=>"011100010",
  18514=>"011000011",
  18515=>"001000000",
  18516=>"111011011",
  18517=>"010000000",
  18518=>"111010011",
  18519=>"100010010",
  18520=>"000111001",
  18521=>"011110101",
  18522=>"100011100",
  18523=>"100000101",
  18524=>"000001000",
  18525=>"010101010",
  18526=>"100111001",
  18527=>"010010001",
  18528=>"110001110",
  18529=>"010110010",
  18530=>"111111100",
  18531=>"101101101",
  18532=>"100000001",
  18533=>"101110101",
  18534=>"011010000",
  18535=>"101001100",
  18536=>"110110010",
  18537=>"000010011",
  18538=>"110001111",
  18539=>"100001000",
  18540=>"010001000",
  18541=>"110000111",
  18542=>"010111011",
  18543=>"000101011",
  18544=>"000010001",
  18545=>"010110011",
  18546=>"011100001",
  18547=>"000010110",
  18548=>"100011111",
  18549=>"010010011",
  18550=>"011101010",
  18551=>"000010001",
  18552=>"010101011",
  18553=>"000010000",
  18554=>"100011001",
  18555=>"110111110",
  18556=>"110101110",
  18557=>"011010110",
  18558=>"010110000",
  18559=>"001001110",
  18560=>"111010100",
  18561=>"001001000",
  18562=>"101110000",
  18563=>"010000011",
  18564=>"100110111",
  18565=>"001100110",
  18566=>"000000111",
  18567=>"110001110",
  18568=>"101010010",
  18569=>"010110111",
  18570=>"100101110",
  18571=>"001010000",
  18572=>"101100010",
  18573=>"010011100",
  18574=>"001100011",
  18575=>"100100001",
  18576=>"001001010",
  18577=>"101111111",
  18578=>"001000010",
  18579=>"100100101",
  18580=>"010000100",
  18581=>"000010101",
  18582=>"110011001",
  18583=>"110010101",
  18584=>"011001001",
  18585=>"101010001",
  18586=>"001010110",
  18587=>"111011101",
  18588=>"001001101",
  18589=>"001100011",
  18590=>"101010110",
  18591=>"011100111",
  18592=>"101101010",
  18593=>"000100100",
  18594=>"000001001",
  18595=>"000110100",
  18596=>"100001001",
  18597=>"100100111",
  18598=>"000000100",
  18599=>"110010111",
  18600=>"111010100",
  18601=>"100010101",
  18602=>"011001001",
  18603=>"100000001",
  18604=>"010010100",
  18605=>"000101100",
  18606=>"100011011",
  18607=>"000001010",
  18608=>"000101101",
  18609=>"000011100",
  18610=>"111011011",
  18611=>"000100010",
  18612=>"111101011",
  18613=>"011100101",
  18614=>"111101011",
  18615=>"110111010",
  18616=>"111000110",
  18617=>"111111011",
  18618=>"000110110",
  18619=>"111101111",
  18620=>"011010000",
  18621=>"110100010",
  18622=>"111110111",
  18623=>"100100011",
  18624=>"100111100",
  18625=>"010000101",
  18626=>"000101001",
  18627=>"001001011",
  18628=>"010111100",
  18629=>"011100010",
  18630=>"100101001",
  18631=>"111101111",
  18632=>"111011100",
  18633=>"001000010",
  18634=>"001000010",
  18635=>"111000101",
  18636=>"100001110",
  18637=>"100111011",
  18638=>"011010111",
  18639=>"010000001",
  18640=>"101111000",
  18641=>"110110011",
  18642=>"011010001",
  18643=>"110000110",
  18644=>"010110001",
  18645=>"011100100",
  18646=>"100101101",
  18647=>"001011111",
  18648=>"101010000",
  18649=>"001100010",
  18650=>"011011111",
  18651=>"111000010",
  18652=>"011101000",
  18653=>"111110110",
  18654=>"010101110",
  18655=>"011001010",
  18656=>"001000101",
  18657=>"000000011",
  18658=>"011001011",
  18659=>"000001100",
  18660=>"010111101",
  18661=>"000100110",
  18662=>"001100000",
  18663=>"001010100",
  18664=>"000000101",
  18665=>"011111111",
  18666=>"000001110",
  18667=>"001011011",
  18668=>"111110000",
  18669=>"000000001",
  18670=>"100001101",
  18671=>"011110010",
  18672=>"101011010",
  18673=>"010010111",
  18674=>"110110010",
  18675=>"001001000",
  18676=>"111101001",
  18677=>"101110001",
  18678=>"000010000",
  18679=>"101000001",
  18680=>"100101000",
  18681=>"011110000",
  18682=>"000001111",
  18683=>"111010101",
  18684=>"111010110",
  18685=>"000011010",
  18686=>"011101111",
  18687=>"010101101",
  18688=>"101001111",
  18689=>"011111110",
  18690=>"010001000",
  18691=>"011110110",
  18692=>"101011001",
  18693=>"000000111",
  18694=>"010100110",
  18695=>"110101111",
  18696=>"101000111",
  18697=>"100010010",
  18698=>"100111010",
  18699=>"100010001",
  18700=>"011101010",
  18701=>"000010001",
  18702=>"100101111",
  18703=>"011000000",
  18704=>"110110111",
  18705=>"011110010",
  18706=>"010010110",
  18707=>"011010011",
  18708=>"010110111",
  18709=>"110100101",
  18710=>"000100011",
  18711=>"101000100",
  18712=>"101111000",
  18713=>"110000011",
  18714=>"011001100",
  18715=>"001101111",
  18716=>"111111101",
  18717=>"001001110",
  18718=>"101111001",
  18719=>"101000000",
  18720=>"100000011",
  18721=>"010001100",
  18722=>"111011010",
  18723=>"000001110",
  18724=>"100001100",
  18725=>"001011000",
  18726=>"100011001",
  18727=>"011011000",
  18728=>"110011100",
  18729=>"100111010",
  18730=>"011111110",
  18731=>"111110010",
  18732=>"100000000",
  18733=>"100001100",
  18734=>"100101011",
  18735=>"011110110",
  18736=>"000101100",
  18737=>"101000010",
  18738=>"111101011",
  18739=>"010100010",
  18740=>"011011010",
  18741=>"010111010",
  18742=>"010100010",
  18743=>"100000011",
  18744=>"111100111",
  18745=>"001010111",
  18746=>"100001111",
  18747=>"110010111",
  18748=>"001001011",
  18749=>"001000110",
  18750=>"001000000",
  18751=>"000100010",
  18752=>"010011011",
  18753=>"011100010",
  18754=>"110001001",
  18755=>"001111101",
  18756=>"001001010",
  18757=>"001011011",
  18758=>"100101010",
  18759=>"100110101",
  18760=>"101101111",
  18761=>"011011000",
  18762=>"011011110",
  18763=>"001001110",
  18764=>"110011001",
  18765=>"100111101",
  18766=>"010111111",
  18767=>"001100101",
  18768=>"000001000",
  18769=>"000100101",
  18770=>"000001011",
  18771=>"100111100",
  18772=>"000100000",
  18773=>"101011110",
  18774=>"001000010",
  18775=>"000001010",
  18776=>"100000100",
  18777=>"010001001",
  18778=>"111010100",
  18779=>"110100001",
  18780=>"101101111",
  18781=>"000000110",
  18782=>"000101110",
  18783=>"011011000",
  18784=>"110101001",
  18785=>"001000110",
  18786=>"111111000",
  18787=>"001010111",
  18788=>"010000110",
  18789=>"110010000",
  18790=>"110000110",
  18791=>"001101101",
  18792=>"001000101",
  18793=>"100100000",
  18794=>"011100010",
  18795=>"111110001",
  18796=>"101111010",
  18797=>"000100110",
  18798=>"100000011",
  18799=>"100110110",
  18800=>"110100111",
  18801=>"011001110",
  18802=>"110100100",
  18803=>"011111101",
  18804=>"001101011",
  18805=>"000000011",
  18806=>"110100111",
  18807=>"101101100",
  18808=>"001010110",
  18809=>"000110100",
  18810=>"101110011",
  18811=>"001000001",
  18812=>"001101010",
  18813=>"011000010",
  18814=>"111101000",
  18815=>"001001101",
  18816=>"001110000",
  18817=>"110100010",
  18818=>"111101111",
  18819=>"001010001",
  18820=>"010001001",
  18821=>"111000111",
  18822=>"100011000",
  18823=>"101010111",
  18824=>"000010110",
  18825=>"000001101",
  18826=>"001110001",
  18827=>"101001110",
  18828=>"010011001",
  18829=>"011100110",
  18830=>"001011100",
  18831=>"011100000",
  18832=>"110000000",
  18833=>"010001100",
  18834=>"110100110",
  18835=>"111111011",
  18836=>"001111110",
  18837=>"010101001",
  18838=>"001101000",
  18839=>"011100111",
  18840=>"111101101",
  18841=>"101100110",
  18842=>"011010010",
  18843=>"010110110",
  18844=>"000101101",
  18845=>"000000110",
  18846=>"011011100",
  18847=>"101000111",
  18848=>"011000011",
  18849=>"000101111",
  18850=>"001110000",
  18851=>"110001111",
  18852=>"000111101",
  18853=>"111001011",
  18854=>"100111110",
  18855=>"011010111",
  18856=>"000001100",
  18857=>"101101110",
  18858=>"100010010",
  18859=>"001110110",
  18860=>"111110110",
  18861=>"001100001",
  18862=>"001010011",
  18863=>"111000101",
  18864=>"111001011",
  18865=>"010000100",
  18866=>"111100000",
  18867=>"000010110",
  18868=>"100111101",
  18869=>"000100010",
  18870=>"011000111",
  18871=>"001000001",
  18872=>"001000100",
  18873=>"101001001",
  18874=>"000010100",
  18875=>"110111100",
  18876=>"110110101",
  18877=>"000011111",
  18878=>"111100100",
  18879=>"010110111",
  18880=>"000010001",
  18881=>"000101010",
  18882=>"011010100",
  18883=>"101110110",
  18884=>"000000011",
  18885=>"010000101",
  18886=>"000001110",
  18887=>"011000101",
  18888=>"010110001",
  18889=>"000000000",
  18890=>"101110111",
  18891=>"111110100",
  18892=>"110100101",
  18893=>"001010100",
  18894=>"100001011",
  18895=>"010110110",
  18896=>"000000011",
  18897=>"010101011",
  18898=>"011100011",
  18899=>"010001000",
  18900=>"101110001",
  18901=>"101101000",
  18902=>"011010011",
  18903=>"000010001",
  18904=>"100101110",
  18905=>"001010110",
  18906=>"110010010",
  18907=>"101011100",
  18908=>"001110111",
  18909=>"111101101",
  18910=>"011101110",
  18911=>"110111110",
  18912=>"100110010",
  18913=>"010101011",
  18914=>"101001001",
  18915=>"101001111",
  18916=>"000100100",
  18917=>"101100001",
  18918=>"010001101",
  18919=>"010101011",
  18920=>"010101101",
  18921=>"000110110",
  18922=>"000000101",
  18923=>"000010000",
  18924=>"111100111",
  18925=>"100010111",
  18926=>"001101111",
  18927=>"110010000",
  18928=>"011101111",
  18929=>"000100010",
  18930=>"010111010",
  18931=>"001000010",
  18932=>"111010010",
  18933=>"100011010",
  18934=>"110000000",
  18935=>"010101111",
  18936=>"101011010",
  18937=>"111011001",
  18938=>"100011110",
  18939=>"011000111",
  18940=>"111011110",
  18941=>"000011000",
  18942=>"100110101",
  18943=>"110010111",
  18944=>"011100100",
  18945=>"110001000",
  18946=>"011001110",
  18947=>"010001010",
  18948=>"010101100",
  18949=>"110011110",
  18950=>"001111101",
  18951=>"111101010",
  18952=>"000011110",
  18953=>"110111110",
  18954=>"001010010",
  18955=>"011000110",
  18956=>"000111011",
  18957=>"100011111",
  18958=>"000110100",
  18959=>"000111111",
  18960=>"110100000",
  18961=>"000011010",
  18962=>"001111100",
  18963=>"011010101",
  18964=>"000011101",
  18965=>"100011100",
  18966=>"111110101",
  18967=>"010001111",
  18968=>"010001001",
  18969=>"100011100",
  18970=>"001010011",
  18971=>"110111010",
  18972=>"001101011",
  18973=>"100001100",
  18974=>"110011001",
  18975=>"111110010",
  18976=>"110110011",
  18977=>"111000110",
  18978=>"010000001",
  18979=>"101110000",
  18980=>"111111111",
  18981=>"000010111",
  18982=>"101110111",
  18983=>"010000010",
  18984=>"101100010",
  18985=>"111001000",
  18986=>"000000101",
  18987=>"100001010",
  18988=>"001110011",
  18989=>"110000100",
  18990=>"111011011",
  18991=>"111111100",
  18992=>"100110100",
  18993=>"011110001",
  18994=>"010101110",
  18995=>"000101111",
  18996=>"111001110",
  18997=>"001000001",
  18998=>"010101011",
  18999=>"101001011",
  19000=>"011011010",
  19001=>"000010000",
  19002=>"111000010",
  19003=>"110100000",
  19004=>"010001101",
  19005=>"000010000",
  19006=>"001101111",
  19007=>"000001101",
  19008=>"111001010",
  19009=>"010001110",
  19010=>"001000010",
  19011=>"111101011",
  19012=>"101001101",
  19013=>"000101000",
  19014=>"110001110",
  19015=>"001011100",
  19016=>"110100111",
  19017=>"100010011",
  19018=>"011001001",
  19019=>"000000000",
  19020=>"100100100",
  19021=>"000001110",
  19022=>"010001101",
  19023=>"010001100",
  19024=>"111000001",
  19025=>"011001111",
  19026=>"101100011",
  19027=>"011101001",
  19028=>"011101010",
  19029=>"011101000",
  19030=>"011000011",
  19031=>"110001000",
  19032=>"111110101",
  19033=>"010111100",
  19034=>"101011001",
  19035=>"001001100",
  19036=>"010101111",
  19037=>"100100100",
  19038=>"111010000",
  19039=>"100101010",
  19040=>"010010011",
  19041=>"100011011",
  19042=>"011001100",
  19043=>"101111110",
  19044=>"101100111",
  19045=>"111111001",
  19046=>"010001010",
  19047=>"011111010",
  19048=>"000010001",
  19049=>"000011101",
  19050=>"011010010",
  19051=>"000010100",
  19052=>"101110100",
  19053=>"010011010",
  19054=>"110000001",
  19055=>"110010101",
  19056=>"101110000",
  19057=>"100100100",
  19058=>"010000001",
  19059=>"010110110",
  19060=>"010111101",
  19061=>"100011111",
  19062=>"100011111",
  19063=>"100110001",
  19064=>"010111011",
  19065=>"010100101",
  19066=>"111011110",
  19067=>"110110111",
  19068=>"010010010",
  19069=>"011100011",
  19070=>"000000010",
  19071=>"101001111",
  19072=>"000000101",
  19073=>"111110000",
  19074=>"110110010",
  19075=>"001100010",
  19076=>"010001100",
  19077=>"110110101",
  19078=>"110010001",
  19079=>"001000101",
  19080=>"000101010",
  19081=>"001100001",
  19082=>"111100011",
  19083=>"100011101",
  19084=>"101011110",
  19085=>"101010001",
  19086=>"010101110",
  19087=>"101110110",
  19088=>"101100001",
  19089=>"100011101",
  19090=>"000011000",
  19091=>"000011011",
  19092=>"010010011",
  19093=>"110010100",
  19094=>"000110110",
  19095=>"101001000",
  19096=>"100111101",
  19097=>"100101010",
  19098=>"110111011",
  19099=>"011010100",
  19100=>"110000001",
  19101=>"111000011",
  19102=>"101001010",
  19103=>"100111000",
  19104=>"111100011",
  19105=>"111111100",
  19106=>"001010110",
  19107=>"110010000",
  19108=>"110011111",
  19109=>"000010100",
  19110=>"011011111",
  19111=>"101011000",
  19112=>"000000100",
  19113=>"000000011",
  19114=>"111011001",
  19115=>"110000000",
  19116=>"100100111",
  19117=>"011111000",
  19118=>"111010110",
  19119=>"101000111",
  19120=>"010010011",
  19121=>"100111000",
  19122=>"111010100",
  19123=>"100011111",
  19124=>"100111010",
  19125=>"101100101",
  19126=>"000000011",
  19127=>"011001000",
  19128=>"100001101",
  19129=>"001000010",
  19130=>"000111010",
  19131=>"000101010",
  19132=>"100000011",
  19133=>"111001001",
  19134=>"110110010",
  19135=>"011000111",
  19136=>"000110110",
  19137=>"110011011",
  19138=>"100101110",
  19139=>"101001101",
  19140=>"111100000",
  19141=>"100010111",
  19142=>"110100000",
  19143=>"010110010",
  19144=>"110001101",
  19145=>"010101110",
  19146=>"100010110",
  19147=>"011010100",
  19148=>"000010100",
  19149=>"010001000",
  19150=>"110110101",
  19151=>"110101010",
  19152=>"010110011",
  19153=>"011101101",
  19154=>"101011110",
  19155=>"010101111",
  19156=>"101101000",
  19157=>"110101011",
  19158=>"000010110",
  19159=>"000011000",
  19160=>"000011000",
  19161=>"100111011",
  19162=>"000111000",
  19163=>"001010001",
  19164=>"001111110",
  19165=>"011000000",
  19166=>"110001110",
  19167=>"000100110",
  19168=>"000011000",
  19169=>"100001010",
  19170=>"010110000",
  19171=>"000011001",
  19172=>"101100001",
  19173=>"111001010",
  19174=>"010101000",
  19175=>"001100101",
  19176=>"001101001",
  19177=>"001111100",
  19178=>"111010111",
  19179=>"011101110",
  19180=>"000100000",
  19181=>"110011111",
  19182=>"010110000",
  19183=>"011001010",
  19184=>"000000101",
  19185=>"000001010",
  19186=>"001011011",
  19187=>"101001001",
  19188=>"010000100",
  19189=>"000100001",
  19190=>"111101010",
  19191=>"010100110",
  19192=>"000010101",
  19193=>"010111111",
  19194=>"010000101",
  19195=>"110000011",
  19196=>"100110101",
  19197=>"110000010",
  19198=>"000000010",
  19199=>"000110101",
  19200=>"000110010",
  19201=>"101000111",
  19202=>"010100011",
  19203=>"010010111",
  19204=>"101101100",
  19205=>"101001110",
  19206=>"110101111",
  19207=>"001001101",
  19208=>"110110111",
  19209=>"010000010",
  19210=>"011110010",
  19211=>"010110001",
  19212=>"010000100",
  19213=>"101011000",
  19214=>"010110110",
  19215=>"011101011",
  19216=>"011010011",
  19217=>"100001001",
  19218=>"001001110",
  19219=>"111001010",
  19220=>"110010111",
  19221=>"001011110",
  19222=>"011000011",
  19223=>"111100010",
  19224=>"110111100",
  19225=>"110100011",
  19226=>"010010110",
  19227=>"110001011",
  19228=>"011101010",
  19229=>"001011110",
  19230=>"000001000",
  19231=>"110011000",
  19232=>"101111111",
  19233=>"001111111",
  19234=>"101101100",
  19235=>"110101110",
  19236=>"010010110",
  19237=>"001000000",
  19238=>"100011010",
  19239=>"000001110",
  19240=>"000010010",
  19241=>"010011111",
  19242=>"001011100",
  19243=>"011110101",
  19244=>"001001100",
  19245=>"010000000",
  19246=>"010101111",
  19247=>"101101001",
  19248=>"110001001",
  19249=>"100110100",
  19250=>"001111000",
  19251=>"010000011",
  19252=>"010110001",
  19253=>"100100110",
  19254=>"000100000",
  19255=>"010010001",
  19256=>"110001100",
  19257=>"111010110",
  19258=>"111101100",
  19259=>"111101110",
  19260=>"000000000",
  19261=>"000010000",
  19262=>"101101101",
  19263=>"111111100",
  19264=>"111001101",
  19265=>"100000001",
  19266=>"101010101",
  19267=>"000101010",
  19268=>"001100000",
  19269=>"100010111",
  19270=>"111101110",
  19271=>"100100000",
  19272=>"000101100",
  19273=>"000000010",
  19274=>"011011010",
  19275=>"010000110",
  19276=>"110100000",
  19277=>"000101011",
  19278=>"111001000",
  19279=>"001011000",
  19280=>"100011001",
  19281=>"011110101",
  19282=>"000010011",
  19283=>"100111111",
  19284=>"000001101",
  19285=>"010101110",
  19286=>"101110101",
  19287=>"101011010",
  19288=>"010111110",
  19289=>"101100111",
  19290=>"110100111",
  19291=>"111100010",
  19292=>"010111100",
  19293=>"000001100",
  19294=>"111111011",
  19295=>"010101000",
  19296=>"011001110",
  19297=>"100100111",
  19298=>"000010000",
  19299=>"110111000",
  19300=>"011000100",
  19301=>"110100000",
  19302=>"101000100",
  19303=>"100111100",
  19304=>"110110000",
  19305=>"111100110",
  19306=>"111101011",
  19307=>"101011010",
  19308=>"001111110",
  19309=>"000111011",
  19310=>"110011000",
  19311=>"000110001",
  19312=>"010000000",
  19313=>"110000101",
  19314=>"010010110",
  19315=>"101001100",
  19316=>"011000111",
  19317=>"100100000",
  19318=>"001011001",
  19319=>"100100011",
  19320=>"010100101",
  19321=>"110110100",
  19322=>"001100101",
  19323=>"001110011",
  19324=>"000100100",
  19325=>"010001001",
  19326=>"111000000",
  19327=>"100011100",
  19328=>"001011101",
  19329=>"110001110",
  19330=>"010001100",
  19331=>"101000111",
  19332=>"111101110",
  19333=>"101101011",
  19334=>"010100101",
  19335=>"100110100",
  19336=>"000111011",
  19337=>"101110001",
  19338=>"100011111",
  19339=>"110010000",
  19340=>"101100101",
  19341=>"010000100",
  19342=>"001110101",
  19343=>"101000111",
  19344=>"111110100",
  19345=>"111011101",
  19346=>"101100000",
  19347=>"100001011",
  19348=>"111111010",
  19349=>"101101011",
  19350=>"000100010",
  19351=>"011100111",
  19352=>"000000110",
  19353=>"101000100",
  19354=>"010011000",
  19355=>"110010000",
  19356=>"101111111",
  19357=>"011110111",
  19358=>"100110100",
  19359=>"011001001",
  19360=>"000101111",
  19361=>"010000000",
  19362=>"010101010",
  19363=>"011111111",
  19364=>"000000110",
  19365=>"011000101",
  19366=>"011111101",
  19367=>"010010101",
  19368=>"101000101",
  19369=>"011100110",
  19370=>"011100000",
  19371=>"101111101",
  19372=>"110000011",
  19373=>"100110111",
  19374=>"010000010",
  19375=>"100000110",
  19376=>"101010111",
  19377=>"001010000",
  19378=>"100111100",
  19379=>"100010001",
  19380=>"001011110",
  19381=>"101111101",
  19382=>"101001001",
  19383=>"000010111",
  19384=>"101000010",
  19385=>"110000000",
  19386=>"011101010",
  19387=>"010000111",
  19388=>"011010000",
  19389=>"001110011",
  19390=>"111101101",
  19391=>"000000010",
  19392=>"001100011",
  19393=>"000110100",
  19394=>"101111011",
  19395=>"111101001",
  19396=>"001010101",
  19397=>"000110011",
  19398=>"011001110",
  19399=>"000011000",
  19400=>"001100100",
  19401=>"011110101",
  19402=>"011000111",
  19403=>"010111110",
  19404=>"110111001",
  19405=>"111111001",
  19406=>"010011111",
  19407=>"110011000",
  19408=>"010010001",
  19409=>"111110110",
  19410=>"001100000",
  19411=>"010110001",
  19412=>"000010100",
  19413=>"000011011",
  19414=>"010101001",
  19415=>"000010010",
  19416=>"111000110",
  19417=>"011101010",
  19418=>"011001001",
  19419=>"010100110",
  19420=>"101101101",
  19421=>"000110011",
  19422=>"011100001",
  19423=>"011101001",
  19424=>"111100000",
  19425=>"000101000",
  19426=>"100001010",
  19427=>"100001010",
  19428=>"000000001",
  19429=>"100111111",
  19430=>"001110100",
  19431=>"100011001",
  19432=>"111101101",
  19433=>"011000010",
  19434=>"011000101",
  19435=>"011011110",
  19436=>"110010100",
  19437=>"000011100",
  19438=>"011101101",
  19439=>"000111011",
  19440=>"011110101",
  19441=>"100001110",
  19442=>"100010010",
  19443=>"011110110",
  19444=>"000000000",
  19445=>"001010100",
  19446=>"001010010",
  19447=>"111111111",
  19448=>"111000010",
  19449=>"000011100",
  19450=>"001100110",
  19451=>"010111010",
  19452=>"011110101",
  19453=>"000001000",
  19454=>"011111100",
  19455=>"111000111",
  19456=>"111111000",
  19457=>"010010110",
  19458=>"111101000",
  19459=>"100001101",
  19460=>"100001101",
  19461=>"011100111",
  19462=>"101110000",
  19463=>"010101100",
  19464=>"101000100",
  19465=>"111011011",
  19466=>"010011111",
  19467=>"011101010",
  19468=>"000000000",
  19469=>"001001011",
  19470=>"100011001",
  19471=>"010011101",
  19472=>"011010111",
  19473=>"000111001",
  19474=>"110101011",
  19475=>"110110111",
  19476=>"111110110",
  19477=>"100111110",
  19478=>"110111100",
  19479=>"111111100",
  19480=>"100111010",
  19481=>"011001110",
  19482=>"010000001",
  19483=>"111011011",
  19484=>"111000100",
  19485=>"110000101",
  19486=>"011101111",
  19487=>"110110011",
  19488=>"011111011",
  19489=>"000100101",
  19490=>"100011101",
  19491=>"011100101",
  19492=>"101011100",
  19493=>"101001010",
  19494=>"010111011",
  19495=>"100110001",
  19496=>"001011010",
  19497=>"101100100",
  19498=>"010011000",
  19499=>"110110001",
  19500=>"011000010",
  19501=>"111111001",
  19502=>"110110101",
  19503=>"111110011",
  19504=>"010101001",
  19505=>"100001011",
  19506=>"001010101",
  19507=>"111010011",
  19508=>"001010110",
  19509=>"001001101",
  19510=>"000110101",
  19511=>"110101110",
  19512=>"100000001",
  19513=>"000101100",
  19514=>"000110000",
  19515=>"100001000",
  19516=>"100000001",
  19517=>"111001100",
  19518=>"101100000",
  19519=>"011001010",
  19520=>"110110100",
  19521=>"000101001",
  19522=>"011111000",
  19523=>"001000001",
  19524=>"010010100",
  19525=>"001010100",
  19526=>"111110111",
  19527=>"001100110",
  19528=>"111001100",
  19529=>"001111000",
  19530=>"001101010",
  19531=>"010101000",
  19532=>"000111111",
  19533=>"010100011",
  19534=>"001010111",
  19535=>"100101000",
  19536=>"001100000",
  19537=>"110001011",
  19538=>"100000110",
  19539=>"001110000",
  19540=>"101001101",
  19541=>"011111101",
  19542=>"011100111",
  19543=>"000000010",
  19544=>"101110100",
  19545=>"101010000",
  19546=>"111011010",
  19547=>"110011010",
  19548=>"101111000",
  19549=>"000110011",
  19550=>"001111111",
  19551=>"010101001",
  19552=>"001100010",
  19553=>"100100001",
  19554=>"000110001",
  19555=>"000111111",
  19556=>"100001011",
  19557=>"001101001",
  19558=>"111010111",
  19559=>"001010110",
  19560=>"101011000",
  19561=>"100111000",
  19562=>"100110011",
  19563=>"011001011",
  19564=>"010011101",
  19565=>"110110101",
  19566=>"001110101",
  19567=>"000010111",
  19568=>"110010010",
  19569=>"111110010",
  19570=>"110001110",
  19571=>"100101111",
  19572=>"001111001",
  19573=>"110100000",
  19574=>"001000110",
  19575=>"101111001",
  19576=>"111111111",
  19577=>"010010000",
  19578=>"001110101",
  19579=>"010010000",
  19580=>"101001001",
  19581=>"010100110",
  19582=>"001000000",
  19583=>"100101001",
  19584=>"011100110",
  19585=>"010111011",
  19586=>"100010111",
  19587=>"000001100",
  19588=>"101011010",
  19589=>"000000010",
  19590=>"100010010",
  19591=>"000000001",
  19592=>"110000000",
  19593=>"100010101",
  19594=>"001010100",
  19595=>"011101101",
  19596=>"100000000",
  19597=>"011010010",
  19598=>"001000000",
  19599=>"111110110",
  19600=>"010100010",
  19601=>"111100001",
  19602=>"111111100",
  19603=>"100000100",
  19604=>"010000000",
  19605=>"111000001",
  19606=>"100010010",
  19607=>"011111001",
  19608=>"010001000",
  19609=>"110010010",
  19610=>"100001100",
  19611=>"001011001",
  19612=>"101010001",
  19613=>"111101011",
  19614=>"101011010",
  19615=>"001101000",
  19616=>"111101011",
  19617=>"011110000",
  19618=>"110010110",
  19619=>"000111000",
  19620=>"101001010",
  19621=>"111101100",
  19622=>"001001111",
  19623=>"101011111",
  19624=>"011101100",
  19625=>"111101000",
  19626=>"000010010",
  19627=>"001001110",
  19628=>"100000110",
  19629=>"011111101",
  19630=>"110100000",
  19631=>"000010010",
  19632=>"100011001",
  19633=>"111001111",
  19634=>"101111101",
  19635=>"001110000",
  19636=>"110111010",
  19637=>"100000010",
  19638=>"001011100",
  19639=>"011000101",
  19640=>"001001010",
  19641=>"101110111",
  19642=>"000101110",
  19643=>"000001010",
  19644=>"101101001",
  19645=>"111110101",
  19646=>"110110011",
  19647=>"110110110",
  19648=>"001011100",
  19649=>"110001111",
  19650=>"111011000",
  19651=>"101001110",
  19652=>"100110100",
  19653=>"001011001",
  19654=>"110100101",
  19655=>"111100010",
  19656=>"010010000",
  19657=>"010101100",
  19658=>"001101101",
  19659=>"101001010",
  19660=>"101000101",
  19661=>"110100011",
  19662=>"010010110",
  19663=>"101001101",
  19664=>"001011000",
  19665=>"001001011",
  19666=>"100100101",
  19667=>"000010011",
  19668=>"001011011",
  19669=>"110001100",
  19670=>"111101100",
  19671=>"111110000",
  19672=>"110101010",
  19673=>"001001111",
  19674=>"010111000",
  19675=>"011111100",
  19676=>"101000100",
  19677=>"000111110",
  19678=>"111100101",
  19679=>"001011000",
  19680=>"111101110",
  19681=>"110010100",
  19682=>"100000010",
  19683=>"001010001",
  19684=>"000100101",
  19685=>"110110000",
  19686=>"100010101",
  19687=>"010110100",
  19688=>"010110100",
  19689=>"110010111",
  19690=>"110101111",
  19691=>"000111110",
  19692=>"101000010",
  19693=>"100101110",
  19694=>"111101110",
  19695=>"001100101",
  19696=>"010000011",
  19697=>"011111101",
  19698=>"001000000",
  19699=>"011001000",
  19700=>"110010000",
  19701=>"011110100",
  19702=>"001010111",
  19703=>"101111100",
  19704=>"011110011",
  19705=>"110110100",
  19706=>"011101111",
  19707=>"110110000",
  19708=>"111100101",
  19709=>"000011101",
  19710=>"111100100",
  19711=>"111000110",
  19712=>"011000011",
  19713=>"010101110",
  19714=>"110011110",
  19715=>"111010101",
  19716=>"011101000",
  19717=>"110111010",
  19718=>"100001111",
  19719=>"011010011",
  19720=>"110110111",
  19721=>"001100000",
  19722=>"011111110",
  19723=>"001111110",
  19724=>"011110101",
  19725=>"000001001",
  19726=>"110101110",
  19727=>"011110111",
  19728=>"100100001",
  19729=>"010100100",
  19730=>"001111100",
  19731=>"111111101",
  19732=>"010101100",
  19733=>"101011110",
  19734=>"001101110",
  19735=>"101000001",
  19736=>"000011101",
  19737=>"000010000",
  19738=>"100011110",
  19739=>"110111010",
  19740=>"110001110",
  19741=>"011111111",
  19742=>"010111111",
  19743=>"010110000",
  19744=>"110000111",
  19745=>"111010001",
  19746=>"000111000",
  19747=>"001111011",
  19748=>"011100100",
  19749=>"100001010",
  19750=>"001111010",
  19751=>"111011111",
  19752=>"001001110",
  19753=>"010110000",
  19754=>"101011001",
  19755=>"101001111",
  19756=>"100110001",
  19757=>"000000000",
  19758=>"010001101",
  19759=>"000001100",
  19760=>"100111110",
  19761=>"011011100",
  19762=>"001010100",
  19763=>"100000110",
  19764=>"111110110",
  19765=>"000011010",
  19766=>"011111111",
  19767=>"000111010",
  19768=>"000111011",
  19769=>"110001111",
  19770=>"111001111",
  19771=>"001110000",
  19772=>"101011110",
  19773=>"111101100",
  19774=>"110100101",
  19775=>"010101110",
  19776=>"010100111",
  19777=>"001101101",
  19778=>"010101010",
  19779=>"101001111",
  19780=>"010000110",
  19781=>"011111111",
  19782=>"011011000",
  19783=>"110100001",
  19784=>"100010100",
  19785=>"011001001",
  19786=>"111000010",
  19787=>"001011100",
  19788=>"101110111",
  19789=>"110001000",
  19790=>"000100111",
  19791=>"111011111",
  19792=>"100000111",
  19793=>"011000011",
  19794=>"010000111",
  19795=>"110001001",
  19796=>"110111111",
  19797=>"101100011",
  19798=>"000001101",
  19799=>"100001101",
  19800=>"010010101",
  19801=>"111000010",
  19802=>"011000100",
  19803=>"100010111",
  19804=>"010001111",
  19805=>"100010110",
  19806=>"011101011",
  19807=>"000010010",
  19808=>"111110011",
  19809=>"010101010",
  19810=>"010101000",
  19811=>"111110111",
  19812=>"001010000",
  19813=>"110100011",
  19814=>"000111001",
  19815=>"010100111",
  19816=>"000111001",
  19817=>"011101000",
  19818=>"100110001",
  19819=>"000100110",
  19820=>"010000100",
  19821=>"100111100",
  19822=>"001101101",
  19823=>"011011100",
  19824=>"110111110",
  19825=>"010000011",
  19826=>"101110111",
  19827=>"000000101",
  19828=>"101101111",
  19829=>"110111000",
  19830=>"111100011",
  19831=>"011000110",
  19832=>"101011000",
  19833=>"010110101",
  19834=>"101010110",
  19835=>"010101011",
  19836=>"000000111",
  19837=>"000100010",
  19838=>"010110010",
  19839=>"101100110",
  19840=>"100101000",
  19841=>"111111000",
  19842=>"001000011",
  19843=>"010111010",
  19844=>"010001000",
  19845=>"001001010",
  19846=>"001111000",
  19847=>"111111001",
  19848=>"110010110",
  19849=>"100100101",
  19850=>"010101000",
  19851=>"001000100",
  19852=>"110010101",
  19853=>"011101100",
  19854=>"110001011",
  19855=>"100010001",
  19856=>"011011010",
  19857=>"110100010",
  19858=>"101111011",
  19859=>"000101111",
  19860=>"101111010",
  19861=>"011010011",
  19862=>"011011011",
  19863=>"010000100",
  19864=>"000101101",
  19865=>"100110110",
  19866=>"110011100",
  19867=>"010111100",
  19868=>"010011100",
  19869=>"111101101",
  19870=>"011011100",
  19871=>"010000001",
  19872=>"100100110",
  19873=>"101000100",
  19874=>"100111010",
  19875=>"010011011",
  19876=>"100011100",
  19877=>"000010011",
  19878=>"011000100",
  19879=>"001010110",
  19880=>"000100100",
  19881=>"010101010",
  19882=>"111101101",
  19883=>"100100101",
  19884=>"010100111",
  19885=>"100111011",
  19886=>"100010001",
  19887=>"100010100",
  19888=>"101000000",
  19889=>"001000101",
  19890=>"111101110",
  19891=>"011111110",
  19892=>"001001010",
  19893=>"000100110",
  19894=>"111011110",
  19895=>"101001110",
  19896=>"010110010",
  19897=>"011001111",
  19898=>"000000001",
  19899=>"110000101",
  19900=>"101110111",
  19901=>"010011010",
  19902=>"110110101",
  19903=>"111100011",
  19904=>"000011010",
  19905=>"010110101",
  19906=>"000101101",
  19907=>"111000111",
  19908=>"000111100",
  19909=>"101111111",
  19910=>"001100011",
  19911=>"111110000",
  19912=>"111110001",
  19913=>"001010101",
  19914=>"010101110",
  19915=>"010111000",
  19916=>"011010110",
  19917=>"010100010",
  19918=>"100100110",
  19919=>"111000100",
  19920=>"000001100",
  19921=>"110000111",
  19922=>"010000100",
  19923=>"011010011",
  19924=>"110101110",
  19925=>"010101010",
  19926=>"011110101",
  19927=>"101110100",
  19928=>"100001110",
  19929=>"001000000",
  19930=>"001000111",
  19931=>"110000011",
  19932=>"000010001",
  19933=>"100011011",
  19934=>"011010011",
  19935=>"110001101",
  19936=>"011000001",
  19937=>"101111010",
  19938=>"001011001",
  19939=>"010111111",
  19940=>"100100110",
  19941=>"101110111",
  19942=>"111101101",
  19943=>"011000000",
  19944=>"100100001",
  19945=>"110100010",
  19946=>"010000111",
  19947=>"111010001",
  19948=>"111010001",
  19949=>"111100000",
  19950=>"001100101",
  19951=>"111001010",
  19952=>"101000101",
  19953=>"000000100",
  19954=>"111010010",
  19955=>"101111010",
  19956=>"110101100",
  19957=>"100000011",
  19958=>"111101100",
  19959=>"110110000",
  19960=>"010011001",
  19961=>"001000101",
  19962=>"010111011",
  19963=>"010111001",
  19964=>"001010100",
  19965=>"011110111",
  19966=>"110010000",
  19967=>"000000010",
  19968=>"010110010",
  19969=>"111101010",
  19970=>"001011010",
  19971=>"111001101",
  19972=>"000000011",
  19973=>"110101100",
  19974=>"010011000",
  19975=>"101101011",
  19976=>"000110010",
  19977=>"101110110",
  19978=>"110010101",
  19979=>"001111011",
  19980=>"011010100",
  19981=>"000001001",
  19982=>"110001111",
  19983=>"010100111",
  19984=>"101011010",
  19985=>"001010010",
  19986=>"000110000",
  19987=>"110001010",
  19988=>"110010111",
  19989=>"001101111",
  19990=>"101010000",
  19991=>"101001000",
  19992=>"010011101",
  19993=>"101001110",
  19994=>"001010000",
  19995=>"000000010",
  19996=>"111111100",
  19997=>"001001011",
  19998=>"001010101",
  19999=>"101110010",
  20000=>"000010111",
  20001=>"111111101",
  20002=>"001001101",
  20003=>"010010000",
  20004=>"101011101",
  20005=>"110001100",
  20006=>"010111110",
  20007=>"000010000",
  20008=>"001100000",
  20009=>"100110100",
  20010=>"100010110",
  20011=>"001100000",
  20012=>"101111010",
  20013=>"111100101",
  20014=>"001101111",
  20015=>"111100001",
  20016=>"010000000",
  20017=>"011000101",
  20018=>"010010001",
  20019=>"011011111",
  20020=>"111001000",
  20021=>"000010111",
  20022=>"100101101",
  20023=>"101110010",
  20024=>"011001000",
  20025=>"100010111",
  20026=>"010110111",
  20027=>"111011001",
  20028=>"110000010",
  20029=>"101011001",
  20030=>"000000111",
  20031=>"110011110",
  20032=>"111010001",
  20033=>"101010111",
  20034=>"110101110",
  20035=>"101001000",
  20036=>"000001110",
  20037=>"100010011",
  20038=>"000010101",
  20039=>"011100100",
  20040=>"101100010",
  20041=>"001100100",
  20042=>"010100111",
  20043=>"110011011",
  20044=>"111111000",
  20045=>"000001000",
  20046=>"001000011",
  20047=>"111100110",
  20048=>"011000011",
  20049=>"110100001",
  20050=>"011001101",
  20051=>"010000011",
  20052=>"100100111",
  20053=>"000000111",
  20054=>"001001011",
  20055=>"111010100",
  20056=>"100000101",
  20057=>"110001000",
  20058=>"110111111",
  20059=>"111010011",
  20060=>"001101011",
  20061=>"111110111",
  20062=>"010111000",
  20063=>"110011010",
  20064=>"111011100",
  20065=>"011110010",
  20066=>"001010000",
  20067=>"001011100",
  20068=>"111110110",
  20069=>"001100111",
  20070=>"000001101",
  20071=>"000110010",
  20072=>"100100110",
  20073=>"011110100",
  20074=>"101110001",
  20075=>"101101110",
  20076=>"000011011",
  20077=>"110110111",
  20078=>"111010010",
  20079=>"111010010",
  20080=>"001111101",
  20081=>"010110101",
  20082=>"001000001",
  20083=>"111110001",
  20084=>"010010001",
  20085=>"111111001",
  20086=>"110001010",
  20087=>"111110011",
  20088=>"001110000",
  20089=>"010000000",
  20090=>"010011110",
  20091=>"111111011",
  20092=>"010101000",
  20093=>"010110000",
  20094=>"011010000",
  20095=>"000110100",
  20096=>"101101011",
  20097=>"111101111",
  20098=>"001101101",
  20099=>"001000011",
  20100=>"100010001",
  20101=>"011101010",
  20102=>"011111101",
  20103=>"011100011",
  20104=>"100000000",
  20105=>"010011111",
  20106=>"101110001",
  20107=>"101100010",
  20108=>"001101010",
  20109=>"000000010",
  20110=>"110000000",
  20111=>"000100110",
  20112=>"001000011",
  20113=>"011000011",
  20114=>"010011001",
  20115=>"001101000",
  20116=>"000100011",
  20117=>"001110010",
  20118=>"001011101",
  20119=>"110010111",
  20120=>"011101001",
  20121=>"001111010",
  20122=>"100000110",
  20123=>"001110101",
  20124=>"111000001",
  20125=>"000011100",
  20126=>"011010110",
  20127=>"001110111",
  20128=>"111011111",
  20129=>"110111101",
  20130=>"000011001",
  20131=>"100111000",
  20132=>"011010010",
  20133=>"001000010",
  20134=>"001101011",
  20135=>"101010000",
  20136=>"001111011",
  20137=>"111110010",
  20138=>"100010100",
  20139=>"000001000",
  20140=>"000111101",
  20141=>"110111010",
  20142=>"111111100",
  20143=>"111011001",
  20144=>"100001010",
  20145=>"000101000",
  20146=>"001110011",
  20147=>"110111101",
  20148=>"011111000",
  20149=>"101111101",
  20150=>"100111101",
  20151=>"001000100",
  20152=>"011110100",
  20153=>"010110110",
  20154=>"011001000",
  20155=>"110000010",
  20156=>"100110110",
  20157=>"101011101",
  20158=>"111101010",
  20159=>"110100001",
  20160=>"101101000",
  20161=>"111000010",
  20162=>"000011011",
  20163=>"010001111",
  20164=>"010111000",
  20165=>"011010011",
  20166=>"101011100",
  20167=>"000001011",
  20168=>"001011010",
  20169=>"000010011",
  20170=>"001001000",
  20171=>"110111011",
  20172=>"101000001",
  20173=>"011010111",
  20174=>"100010111",
  20175=>"101101001",
  20176=>"110011111",
  20177=>"110110111",
  20178=>"101000010",
  20179=>"101100101",
  20180=>"100110001",
  20181=>"011001010",
  20182=>"001100010",
  20183=>"111111011",
  20184=>"111001101",
  20185=>"110100100",
  20186=>"110000100",
  20187=>"101010010",
  20188=>"001000011",
  20189=>"110001111",
  20190=>"011010100",
  20191=>"001100011",
  20192=>"100100101",
  20193=>"100001001",
  20194=>"101111111",
  20195=>"110011010",
  20196=>"001001000",
  20197=>"011110101",
  20198=>"010010101",
  20199=>"000011010",
  20200=>"000110011",
  20201=>"001011110",
  20202=>"101110100",
  20203=>"011010001",
  20204=>"011001001",
  20205=>"000111101",
  20206=>"000001101",
  20207=>"011100010",
  20208=>"111001101",
  20209=>"100011011",
  20210=>"000110111",
  20211=>"010110100",
  20212=>"101010011",
  20213=>"000011000",
  20214=>"010111101",
  20215=>"111101101",
  20216=>"110001100",
  20217=>"100111101",
  20218=>"100001010",
  20219=>"010100000",
  20220=>"111101000",
  20221=>"001111101",
  20222=>"101001110",
  20223=>"100011010",
  20224=>"011111111",
  20225=>"011000001",
  20226=>"111010000",
  20227=>"000000110",
  20228=>"101010001",
  20229=>"110010110",
  20230=>"010101001",
  20231=>"001001001",
  20232=>"010000111",
  20233=>"101111111",
  20234=>"110101001",
  20235=>"000111000",
  20236=>"011000000",
  20237=>"101111001",
  20238=>"111110110",
  20239=>"010101000",
  20240=>"011011111",
  20241=>"010111100",
  20242=>"010000101",
  20243=>"100000100",
  20244=>"000011010",
  20245=>"001110101",
  20246=>"010011011",
  20247=>"001111101",
  20248=>"101011100",
  20249=>"001101000",
  20250=>"101110000",
  20251=>"110011111",
  20252=>"000000101",
  20253=>"011010001",
  20254=>"101101011",
  20255=>"101110101",
  20256=>"000001010",
  20257=>"001101101",
  20258=>"000101011",
  20259=>"111000111",
  20260=>"010100001",
  20261=>"001110010",
  20262=>"101101011",
  20263=>"101110001",
  20264=>"110100111",
  20265=>"010111101",
  20266=>"010001010",
  20267=>"000110000",
  20268=>"101011111",
  20269=>"100111001",
  20270=>"011110111",
  20271=>"010101111",
  20272=>"100100110",
  20273=>"100001011",
  20274=>"001001101",
  20275=>"101110000",
  20276=>"001011101",
  20277=>"101110010",
  20278=>"111101000",
  20279=>"001010001",
  20280=>"000000010",
  20281=>"000111010",
  20282=>"110111110",
  20283=>"101111101",
  20284=>"000000010",
  20285=>"001101000",
  20286=>"100101011",
  20287=>"011110000",
  20288=>"111011000",
  20289=>"101010110",
  20290=>"000111101",
  20291=>"111111010",
  20292=>"111111110",
  20293=>"000110101",
  20294=>"100000011",
  20295=>"011111111",
  20296=>"001111001",
  20297=>"110111101",
  20298=>"001101110",
  20299=>"101000101",
  20300=>"100011110",
  20301=>"011111100",
  20302=>"001110101",
  20303=>"100001101",
  20304=>"010101010",
  20305=>"011001011",
  20306=>"110100011",
  20307=>"100010110",
  20308=>"000101001",
  20309=>"011100111",
  20310=>"000101101",
  20311=>"110101001",
  20312=>"101110000",
  20313=>"110000110",
  20314=>"111111000",
  20315=>"000001010",
  20316=>"000100000",
  20317=>"110010000",
  20318=>"010000000",
  20319=>"111011101",
  20320=>"001000001",
  20321=>"000011010",
  20322=>"001011100",
  20323=>"111110010",
  20324=>"101110111",
  20325=>"100001110",
  20326=>"111101100",
  20327=>"100110101",
  20328=>"001011000",
  20329=>"000010101",
  20330=>"101001111",
  20331=>"000000010",
  20332=>"011111010",
  20333=>"111010110",
  20334=>"111010001",
  20335=>"111001111",
  20336=>"010000101",
  20337=>"001011001",
  20338=>"000000100",
  20339=>"110001100",
  20340=>"001101011",
  20341=>"010100111",
  20342=>"111100111",
  20343=>"110010100",
  20344=>"110010110",
  20345=>"100011110",
  20346=>"011001010",
  20347=>"100111001",
  20348=>"011000101",
  20349=>"011000000",
  20350=>"011000000",
  20351=>"001010110",
  20352=>"110110100",
  20353=>"011111100",
  20354=>"110101000",
  20355=>"100111011",
  20356=>"000111010",
  20357=>"001010010",
  20358=>"000000010",
  20359=>"001100111",
  20360=>"101000101",
  20361=>"101001011",
  20362=>"101001000",
  20363=>"001011011",
  20364=>"001000101",
  20365=>"111111100",
  20366=>"110110000",
  20367=>"011000111",
  20368=>"100101001",
  20369=>"110101001",
  20370=>"110000000",
  20371=>"100001011",
  20372=>"001011010",
  20373=>"000111001",
  20374=>"000000101",
  20375=>"011011001",
  20376=>"001111100",
  20377=>"110111110",
  20378=>"001000110",
  20379=>"110101000",
  20380=>"101010101",
  20381=>"001101010",
  20382=>"011000111",
  20383=>"111101111",
  20384=>"100110101",
  20385=>"111010101",
  20386=>"011010100",
  20387=>"111100111",
  20388=>"110001000",
  20389=>"000010011",
  20390=>"100100110",
  20391=>"101111001",
  20392=>"111001110",
  20393=>"101111111",
  20394=>"111000001",
  20395=>"100100000",
  20396=>"100001011",
  20397=>"111111110",
  20398=>"100111101",
  20399=>"110000110",
  20400=>"010101010",
  20401=>"010000000",
  20402=>"101100100",
  20403=>"001001001",
  20404=>"011010001",
  20405=>"100100011",
  20406=>"110110101",
  20407=>"010111001",
  20408=>"111100101",
  20409=>"011110110",
  20410=>"000001101",
  20411=>"111010001",
  20412=>"101000111",
  20413=>"010000001",
  20414=>"110001111",
  20415=>"011101110",
  20416=>"110011011",
  20417=>"000110101",
  20418=>"100010011",
  20419=>"001000110",
  20420=>"000010100",
  20421=>"101010100",
  20422=>"101100010",
  20423=>"101010000",
  20424=>"000110000",
  20425=>"111110111",
  20426=>"010110110",
  20427=>"111001100",
  20428=>"010100100",
  20429=>"010010101",
  20430=>"101100011",
  20431=>"111010111",
  20432=>"001011110",
  20433=>"001001100",
  20434=>"101010010",
  20435=>"010000110",
  20436=>"110101100",
  20437=>"010010000",
  20438=>"110011000",
  20439=>"111011001",
  20440=>"000001001",
  20441=>"110101001",
  20442=>"111101110",
  20443=>"001101110",
  20444=>"100011010",
  20445=>"110111000",
  20446=>"111011110",
  20447=>"000010000",
  20448=>"101101010",
  20449=>"100100101",
  20450=>"111010001",
  20451=>"101000000",
  20452=>"000010010",
  20453=>"010010111",
  20454=>"111101101",
  20455=>"110010000",
  20456=>"100101010",
  20457=>"001001011",
  20458=>"100111111",
  20459=>"000011110",
  20460=>"011101110",
  20461=>"011011011",
  20462=>"011110001",
  20463=>"111111011",
  20464=>"000010110",
  20465=>"111110000",
  20466=>"010001111",
  20467=>"010001101",
  20468=>"000011111",
  20469=>"000001001",
  20470=>"011100000",
  20471=>"011101101",
  20472=>"101001010",
  20473=>"111100010",
  20474=>"101001101",
  20475=>"111000100",
  20476=>"101101001",
  20477=>"101100101",
  20478=>"101111011",
  20479=>"000111010",
  20480=>"100011111",
  20481=>"100000000",
  20482=>"111110101",
  20483=>"111111100",
  20484=>"001000111",
  20485=>"110011000",
  20486=>"000010100",
  20487=>"100000110",
  20488=>"001110000",
  20489=>"000001100",
  20490=>"101111000",
  20491=>"000100110",
  20492=>"000001111",
  20493=>"000110110",
  20494=>"011101001",
  20495=>"010100101",
  20496=>"000010110",
  20497=>"010111110",
  20498=>"010010000",
  20499=>"101011000",
  20500=>"101001000",
  20501=>"001000110",
  20502=>"011010011",
  20503=>"000101100",
  20504=>"101101000",
  20505=>"001001010",
  20506=>"011010000",
  20507=>"110000101",
  20508=>"110111001",
  20509=>"000011011",
  20510=>"010110001",
  20511=>"111011101",
  20512=>"111010101",
  20513=>"100111100",
  20514=>"100000000",
  20515=>"110010100",
  20516=>"001111101",
  20517=>"101000010",
  20518=>"011001111",
  20519=>"011011101",
  20520=>"100011000",
  20521=>"111011100",
  20522=>"111011101",
  20523=>"100101011",
  20524=>"111100100",
  20525=>"000010010",
  20526=>"111111101",
  20527=>"000101000",
  20528=>"010110010",
  20529=>"000000111",
  20530=>"101010111",
  20531=>"111100001",
  20532=>"101010000",
  20533=>"100001011",
  20534=>"000001100",
  20535=>"100111111",
  20536=>"001000010",
  20537=>"011100100",
  20538=>"010111011",
  20539=>"110010000",
  20540=>"110111011",
  20541=>"000010011",
  20542=>"011111000",
  20543=>"111001010",
  20544=>"101110110",
  20545=>"101101110",
  20546=>"011110110",
  20547=>"111010011",
  20548=>"010100001",
  20549=>"001011000",
  20550=>"011111101",
  20551=>"100010100",
  20552=>"011111000",
  20553=>"101101101",
  20554=>"111000111",
  20555=>"011011100",
  20556=>"000000001",
  20557=>"111011000",
  20558=>"010110111",
  20559=>"000000011",
  20560=>"101101000",
  20561=>"010010011",
  20562=>"100100111",
  20563=>"001100010",
  20564=>"110001001",
  20565=>"110010101",
  20566=>"110111011",
  20567=>"110100010",
  20568=>"011100101",
  20569=>"011101001",
  20570=>"110000100",
  20571=>"000001001",
  20572=>"110011010",
  20573=>"101101100",
  20574=>"010110100",
  20575=>"000000000",
  20576=>"001100000",
  20577=>"000000110",
  20578=>"111100110",
  20579=>"010011010",
  20580=>"111100101",
  20581=>"011000110",
  20582=>"111110000",
  20583=>"001111111",
  20584=>"110110010",
  20585=>"110011101",
  20586=>"011110111",
  20587=>"010010001",
  20588=>"101100010",
  20589=>"100110000",
  20590=>"101011000",
  20591=>"011100111",
  20592=>"010001100",
  20593=>"110001110",
  20594=>"110110011",
  20595=>"111010101",
  20596=>"110011010",
  20597=>"110101001",
  20598=>"111000101",
  20599=>"011101101",
  20600=>"110000001",
  20601=>"001000000",
  20602=>"101001000",
  20603=>"100110000",
  20604=>"010111111",
  20605=>"110001111",
  20606=>"110110001",
  20607=>"000011111",
  20608=>"100110010",
  20609=>"111101110",
  20610=>"101000011",
  20611=>"010101000",
  20612=>"101010100",
  20613=>"101101101",
  20614=>"111100001",
  20615=>"011111011",
  20616=>"000010110",
  20617=>"001111111",
  20618=>"101100001",
  20619=>"010101001",
  20620=>"111101111",
  20621=>"000100111",
  20622=>"000011001",
  20623=>"000010100",
  20624=>"100101110",
  20625=>"011010011",
  20626=>"101110000",
  20627=>"011011111",
  20628=>"010011011",
  20629=>"011100100",
  20630=>"000010101",
  20631=>"111111010",
  20632=>"111000001",
  20633=>"110001101",
  20634=>"001010001",
  20635=>"111100111",
  20636=>"100110000",
  20637=>"011110101",
  20638=>"101001101",
  20639=>"011001100",
  20640=>"011110010",
  20641=>"000010000",
  20642=>"001100011",
  20643=>"111110100",
  20644=>"111001011",
  20645=>"101001110",
  20646=>"001100110",
  20647=>"100000101",
  20648=>"111100110",
  20649=>"110111111",
  20650=>"100101001",
  20651=>"100000110",
  20652=>"010100000",
  20653=>"111111011",
  20654=>"100110001",
  20655=>"010100011",
  20656=>"010011101",
  20657=>"100100100",
  20658=>"000111001",
  20659=>"101000010",
  20660=>"110001110",
  20661=>"110111110",
  20662=>"100101110",
  20663=>"001011101",
  20664=>"011100100",
  20665=>"100100100",
  20666=>"110110110",
  20667=>"000011010",
  20668=>"101011101",
  20669=>"101010000",
  20670=>"100111001",
  20671=>"100001101",
  20672=>"011011001",
  20673=>"000111110",
  20674=>"110011111",
  20675=>"100010011",
  20676=>"101110000",
  20677=>"100001001",
  20678=>"010011101",
  20679=>"101100110",
  20680=>"111011011",
  20681=>"000111011",
  20682=>"101011011",
  20683=>"101101110",
  20684=>"011011010",
  20685=>"010110100",
  20686=>"101101011",
  20687=>"001000000",
  20688=>"011110110",
  20689=>"110001100",
  20690=>"001110111",
  20691=>"011101011",
  20692=>"101100001",
  20693=>"011000011",
  20694=>"000110111",
  20695=>"100010101",
  20696=>"111111001",
  20697=>"000110011",
  20698=>"111001000",
  20699=>"010010001",
  20700=>"111000001",
  20701=>"000000100",
  20702=>"111101011",
  20703=>"010111101",
  20704=>"101100011",
  20705=>"110011110",
  20706=>"000110101",
  20707=>"000001010",
  20708=>"100010010",
  20709=>"001110111",
  20710=>"111111000",
  20711=>"001100101",
  20712=>"011010110",
  20713=>"000101101",
  20714=>"001111010",
  20715=>"000000100",
  20716=>"010010010",
  20717=>"000101010",
  20718=>"000001110",
  20719=>"101010111",
  20720=>"101011001",
  20721=>"001111100",
  20722=>"011010011",
  20723=>"111000100",
  20724=>"011000010",
  20725=>"100100010",
  20726=>"110001100",
  20727=>"100010100",
  20728=>"001000101",
  20729=>"010010000",
  20730=>"001000111",
  20731=>"100001011",
  20732=>"001110010",
  20733=>"001001001",
  20734=>"011011110",
  20735=>"011001001",
  20736=>"110111001",
  20737=>"010010111",
  20738=>"111010011",
  20739=>"011110100",
  20740=>"111100100",
  20741=>"110101010",
  20742=>"110110101",
  20743=>"000111100",
  20744=>"110010011",
  20745=>"100100011",
  20746=>"010100111",
  20747=>"100100000",
  20748=>"001100000",
  20749=>"000001010",
  20750=>"001110110",
  20751=>"010101101",
  20752=>"110110110",
  20753=>"101010110",
  20754=>"100000111",
  20755=>"101111110",
  20756=>"110110111",
  20757=>"101100000",
  20758=>"100110000",
  20759=>"101011010",
  20760=>"101010100",
  20761=>"011110001",
  20762=>"110011011",
  20763=>"111111001",
  20764=>"110000011",
  20765=>"010010100",
  20766=>"001000011",
  20767=>"001001001",
  20768=>"100110010",
  20769=>"000001011",
  20770=>"101001011",
  20771=>"000010101",
  20772=>"010010101",
  20773=>"000001111",
  20774=>"000000110",
  20775=>"011110000",
  20776=>"100011110",
  20777=>"101011010",
  20778=>"100100100",
  20779=>"110101110",
  20780=>"110111111",
  20781=>"010100011",
  20782=>"110101111",
  20783=>"111111111",
  20784=>"000111110",
  20785=>"010111111",
  20786=>"110100000",
  20787=>"101010101",
  20788=>"000000001",
  20789=>"111101011",
  20790=>"100110100",
  20791=>"111110101",
  20792=>"000011110",
  20793=>"000010011",
  20794=>"100101000",
  20795=>"011010010",
  20796=>"011011010",
  20797=>"101110110",
  20798=>"011100000",
  20799=>"001010100",
  20800=>"010110000",
  20801=>"101100101",
  20802=>"101100100",
  20803=>"001101100",
  20804=>"111101100",
  20805=>"101100000",
  20806=>"111101110",
  20807=>"000111000",
  20808=>"110010101",
  20809=>"100000100",
  20810=>"100101111",
  20811=>"110111100",
  20812=>"011110011",
  20813=>"110000001",
  20814=>"110100110",
  20815=>"110010110",
  20816=>"010011010",
  20817=>"100000010",
  20818=>"111100000",
  20819=>"101101000",
  20820=>"110000101",
  20821=>"110001110",
  20822=>"000010011",
  20823=>"010011111",
  20824=>"110001001",
  20825=>"000111101",
  20826=>"010111100",
  20827=>"110011010",
  20828=>"000111000",
  20829=>"111100110",
  20830=>"010100110",
  20831=>"111110011",
  20832=>"111011101",
  20833=>"011010111",
  20834=>"001001011",
  20835=>"000000000",
  20836=>"101100000",
  20837=>"101000011",
  20838=>"110111011",
  20839=>"000000010",
  20840=>"110100111",
  20841=>"010111011",
  20842=>"100010100",
  20843=>"110001100",
  20844=>"100001001",
  20845=>"000100011",
  20846=>"100100001",
  20847=>"001010001",
  20848=>"111011110",
  20849=>"111100000",
  20850=>"100010001",
  20851=>"010111101",
  20852=>"100111001",
  20853=>"110001010",
  20854=>"010000010",
  20855=>"001011001",
  20856=>"010001010",
  20857=>"111101111",
  20858=>"000101000",
  20859=>"011101100",
  20860=>"111010100",
  20861=>"000110011",
  20862=>"000101100",
  20863=>"000000101",
  20864=>"110000110",
  20865=>"000000011",
  20866=>"100111010",
  20867=>"000000010",
  20868=>"110110000",
  20869=>"001111000",
  20870=>"001100010",
  20871=>"100101101",
  20872=>"101100101",
  20873=>"110000101",
  20874=>"011101000",
  20875=>"001111111",
  20876=>"111100100",
  20877=>"000110100",
  20878=>"111101111",
  20879=>"101110001",
  20880=>"101000101",
  20881=>"111000101",
  20882=>"000100000",
  20883=>"101010010",
  20884=>"110110011",
  20885=>"101010111",
  20886=>"100010000",
  20887=>"001000111",
  20888=>"011011111",
  20889=>"000100000",
  20890=>"000001011",
  20891=>"110100001",
  20892=>"110000011",
  20893=>"111101010",
  20894=>"100000000",
  20895=>"110010010",
  20896=>"001101011",
  20897=>"110100011",
  20898=>"011000101",
  20899=>"011001101",
  20900=>"110101100",
  20901=>"000101110",
  20902=>"110100011",
  20903=>"101011000",
  20904=>"000110011",
  20905=>"000010000",
  20906=>"100001101",
  20907=>"010011110",
  20908=>"011010011",
  20909=>"110101011",
  20910=>"101101110",
  20911=>"010001100",
  20912=>"010101000",
  20913=>"101001000",
  20914=>"000100110",
  20915=>"100010111",
  20916=>"111011001",
  20917=>"111001010",
  20918=>"000101000",
  20919=>"110011001",
  20920=>"100100110",
  20921=>"001111101",
  20922=>"010010010",
  20923=>"101100111",
  20924=>"101101101",
  20925=>"000101100",
  20926=>"100001111",
  20927=>"000101110",
  20928=>"010001011",
  20929=>"001100110",
  20930=>"101010100",
  20931=>"100111011",
  20932=>"011110101",
  20933=>"101010010",
  20934=>"010110001",
  20935=>"010101101",
  20936=>"001001001",
  20937=>"101010001",
  20938=>"111010011",
  20939=>"001101111",
  20940=>"001010101",
  20941=>"110101000",
  20942=>"101101000",
  20943=>"111000010",
  20944=>"001100010",
  20945=>"001100011",
  20946=>"011011011",
  20947=>"101111101",
  20948=>"101000010",
  20949=>"000100101",
  20950=>"011001100",
  20951=>"111111000",
  20952=>"111010010",
  20953=>"001011100",
  20954=>"100010000",
  20955=>"011111111",
  20956=>"011100101",
  20957=>"001000001",
  20958=>"110100001",
  20959=>"010100000",
  20960=>"010000001",
  20961=>"000011001",
  20962=>"001000101",
  20963=>"111001000",
  20964=>"010110100",
  20965=>"100111010",
  20966=>"110000010",
  20967=>"000000110",
  20968=>"010000110",
  20969=>"101110001",
  20970=>"101110001",
  20971=>"010110101",
  20972=>"011001001",
  20973=>"110001011",
  20974=>"110100011",
  20975=>"011101000",
  20976=>"011110001",
  20977=>"010110001",
  20978=>"100010000",
  20979=>"000000001",
  20980=>"110001100",
  20981=>"010101110",
  20982=>"110010001",
  20983=>"110011001",
  20984=>"000100010",
  20985=>"001001000",
  20986=>"110100111",
  20987=>"010000110",
  20988=>"110011101",
  20989=>"110011000",
  20990=>"111010101",
  20991=>"100000100",
  20992=>"001001010",
  20993=>"001010100",
  20994=>"010111110",
  20995=>"000011111",
  20996=>"000100000",
  20997=>"001001111",
  20998=>"010011111",
  20999=>"111101011",
  21000=>"000110110",
  21001=>"100011100",
  21002=>"000010110",
  21003=>"111010101",
  21004=>"101110000",
  21005=>"010100110",
  21006=>"100010101",
  21007=>"101101101",
  21008=>"011001110",
  21009=>"011111011",
  21010=>"000100100",
  21011=>"011100101",
  21012=>"000010001",
  21013=>"010111011",
  21014=>"111111111",
  21015=>"000111001",
  21016=>"000000110",
  21017=>"011100111",
  21018=>"111011110",
  21019=>"101111110",
  21020=>"001000000",
  21021=>"100100011",
  21022=>"011001000",
  21023=>"000101010",
  21024=>"110111001",
  21025=>"101000111",
  21026=>"111001110",
  21027=>"001000101",
  21028=>"000011011",
  21029=>"011001011",
  21030=>"100101111",
  21031=>"011100000",
  21032=>"100011000",
  21033=>"101100101",
  21034=>"111110110",
  21035=>"111100110",
  21036=>"100110110",
  21037=>"100000111",
  21038=>"000101010",
  21039=>"110110000",
  21040=>"001100010",
  21041=>"011110000",
  21042=>"010011010",
  21043=>"011100000",
  21044=>"001100000",
  21045=>"111111110",
  21046=>"100011100",
  21047=>"010011011",
  21048=>"110111001",
  21049=>"101001001",
  21050=>"000001110",
  21051=>"111001100",
  21052=>"111110011",
  21053=>"001100111",
  21054=>"011111100",
  21055=>"101100100",
  21056=>"110010001",
  21057=>"101011011",
  21058=>"101110010",
  21059=>"101100111",
  21060=>"010000110",
  21061=>"111100101",
  21062=>"111101001",
  21063=>"100010111",
  21064=>"010100001",
  21065=>"110111110",
  21066=>"100000110",
  21067=>"011100011",
  21068=>"101011110",
  21069=>"001110110",
  21070=>"101101101",
  21071=>"001110000",
  21072=>"111000010",
  21073=>"010001000",
  21074=>"010110110",
  21075=>"000001000",
  21076=>"001001110",
  21077=>"100100000",
  21078=>"011000100",
  21079=>"001110111",
  21080=>"111001101",
  21081=>"101111111",
  21082=>"100001110",
  21083=>"000110000",
  21084=>"100111010",
  21085=>"000100011",
  21086=>"101110101",
  21087=>"100000110",
  21088=>"000001000",
  21089=>"000101110",
  21090=>"111010110",
  21091=>"100010000",
  21092=>"011010111",
  21093=>"001010001",
  21094=>"011101111",
  21095=>"100001111",
  21096=>"000111000",
  21097=>"111010111",
  21098=>"000000001",
  21099=>"000101000",
  21100=>"000011111",
  21101=>"110001111",
  21102=>"000100101",
  21103=>"111110011",
  21104=>"111111001",
  21105=>"110110110",
  21106=>"111100011",
  21107=>"011010000",
  21108=>"000001011",
  21109=>"011110100",
  21110=>"000011100",
  21111=>"000011111",
  21112=>"110000010",
  21113=>"000011101",
  21114=>"001101000",
  21115=>"111101011",
  21116=>"111100000",
  21117=>"110000001",
  21118=>"000001000",
  21119=>"111101000",
  21120=>"000000000",
  21121=>"010100011",
  21122=>"111100111",
  21123=>"100100010",
  21124=>"101101001",
  21125=>"110001000",
  21126=>"110010011",
  21127=>"110011000",
  21128=>"001110010",
  21129=>"000010100",
  21130=>"111101110",
  21131=>"110011110",
  21132=>"001101110",
  21133=>"010011001",
  21134=>"111010010",
  21135=>"110010101",
  21136=>"001001011",
  21137=>"111111010",
  21138=>"100001001",
  21139=>"101001000",
  21140=>"111111000",
  21141=>"110101101",
  21142=>"110000101",
  21143=>"100101011",
  21144=>"010101010",
  21145=>"111100100",
  21146=>"001111010",
  21147=>"001101101",
  21148=>"101000010",
  21149=>"111000101",
  21150=>"101101111",
  21151=>"110010011",
  21152=>"101000101",
  21153=>"011101000",
  21154=>"100110101",
  21155=>"000111111",
  21156=>"111111010",
  21157=>"000000100",
  21158=>"010000100",
  21159=>"001001011",
  21160=>"100111011",
  21161=>"001111001",
  21162=>"111100111",
  21163=>"101001100",
  21164=>"000010010",
  21165=>"110100001",
  21166=>"111101001",
  21167=>"011000100",
  21168=>"101101110",
  21169=>"000111010",
  21170=>"110100111",
  21171=>"001010010",
  21172=>"111010000",
  21173=>"011010111",
  21174=>"010110110",
  21175=>"101001000",
  21176=>"001010111",
  21177=>"000101010",
  21178=>"000100001",
  21179=>"001111010",
  21180=>"001000100",
  21181=>"010110100",
  21182=>"011100001",
  21183=>"010101101",
  21184=>"110101111",
  21185=>"000110100",
  21186=>"111111011",
  21187=>"101011111",
  21188=>"010110111",
  21189=>"010011101",
  21190=>"001001110",
  21191=>"101000100",
  21192=>"010101100",
  21193=>"101110010",
  21194=>"111001010",
  21195=>"110100000",
  21196=>"000101110",
  21197=>"111011111",
  21198=>"110001000",
  21199=>"101100000",
  21200=>"111011010",
  21201=>"111011111",
  21202=>"110010101",
  21203=>"000001011",
  21204=>"010001011",
  21205=>"000110000",
  21206=>"011000001",
  21207=>"010111100",
  21208=>"101010010",
  21209=>"110010100",
  21210=>"011110111",
  21211=>"111100111",
  21212=>"100101111",
  21213=>"100101001",
  21214=>"010011100",
  21215=>"001110011",
  21216=>"100101000",
  21217=>"111000101",
  21218=>"010001110",
  21219=>"111010111",
  21220=>"111010101",
  21221=>"011001011",
  21222=>"000010000",
  21223=>"001001000",
  21224=>"100010110",
  21225=>"011010000",
  21226=>"100101101",
  21227=>"100000001",
  21228=>"111100100",
  21229=>"010001100",
  21230=>"111100100",
  21231=>"110000110",
  21232=>"010011110",
  21233=>"110101011",
  21234=>"110101011",
  21235=>"011000000",
  21236=>"101001001",
  21237=>"101111110",
  21238=>"110011001",
  21239=>"100111101",
  21240=>"110111011",
  21241=>"100011011",
  21242=>"011001001",
  21243=>"010101110",
  21244=>"011010000",
  21245=>"101100001",
  21246=>"010010010",
  21247=>"110000110",
  21248=>"110010101",
  21249=>"110010011",
  21250=>"011111100",
  21251=>"101100001",
  21252=>"100001100",
  21253=>"110100011",
  21254=>"010111001",
  21255=>"001011000",
  21256=>"011011101",
  21257=>"111100111",
  21258=>"000011011",
  21259=>"101001010",
  21260=>"101001000",
  21261=>"111011000",
  21262=>"100010001",
  21263=>"100001110",
  21264=>"001010010",
  21265=>"000100100",
  21266=>"010101001",
  21267=>"100010001",
  21268=>"011010010",
  21269=>"001000001",
  21270=>"010110010",
  21271=>"111000000",
  21272=>"111000101",
  21273=>"100111110",
  21274=>"110100010",
  21275=>"101111011",
  21276=>"100011100",
  21277=>"101010111",
  21278=>"110001010",
  21279=>"001111000",
  21280=>"111110110",
  21281=>"100100011",
  21282=>"101011101",
  21283=>"000101100",
  21284=>"011010101",
  21285=>"010101010",
  21286=>"001110011",
  21287=>"010010010",
  21288=>"000011100",
  21289=>"110111001",
  21290=>"111100110",
  21291=>"011011110",
  21292=>"111100001",
  21293=>"010110001",
  21294=>"100100111",
  21295=>"000110101",
  21296=>"000011101",
  21297=>"110011110",
  21298=>"101011100",
  21299=>"000101100",
  21300=>"111011100",
  21301=>"110100010",
  21302=>"100000000",
  21303=>"001010110",
  21304=>"100010001",
  21305=>"010010110",
  21306=>"100001111",
  21307=>"001101001",
  21308=>"011110101",
  21309=>"101111101",
  21310=>"000000010",
  21311=>"011000001",
  21312=>"000011101",
  21313=>"001001010",
  21314=>"100000000",
  21315=>"010000100",
  21316=>"000110010",
  21317=>"000101101",
  21318=>"011111001",
  21319=>"110100011",
  21320=>"111110000",
  21321=>"100010000",
  21322=>"110100110",
  21323=>"100101000",
  21324=>"111100011",
  21325=>"110011101",
  21326=>"111111110",
  21327=>"001110000",
  21328=>"100101111",
  21329=>"000000011",
  21330=>"010000110",
  21331=>"001000111",
  21332=>"111000010",
  21333=>"010011100",
  21334=>"011100111",
  21335=>"100110100",
  21336=>"100011000",
  21337=>"011001101",
  21338=>"010111000",
  21339=>"010101111",
  21340=>"111111111",
  21341=>"010111000",
  21342=>"010010100",
  21343=>"101110010",
  21344=>"101100100",
  21345=>"111111101",
  21346=>"101011000",
  21347=>"001111110",
  21348=>"101010111",
  21349=>"111100001",
  21350=>"010000000",
  21351=>"111011110",
  21352=>"110100110",
  21353=>"100001100",
  21354=>"100001110",
  21355=>"101001011",
  21356=>"001101011",
  21357=>"101101100",
  21358=>"100111100",
  21359=>"000011111",
  21360=>"111110111",
  21361=>"101010010",
  21362=>"000011000",
  21363=>"000011100",
  21364=>"001010000",
  21365=>"111100100",
  21366=>"110010110",
  21367=>"011011011",
  21368=>"011011000",
  21369=>"110101101",
  21370=>"011001000",
  21371=>"001101010",
  21372=>"111110110",
  21373=>"111011001",
  21374=>"111010101",
  21375=>"110010101",
  21376=>"011110010",
  21377=>"100010001",
  21378=>"000010011",
  21379=>"110101011",
  21380=>"100110100",
  21381=>"011011001",
  21382=>"111111111",
  21383=>"000010010",
  21384=>"110011111",
  21385=>"100001111",
  21386=>"000011111",
  21387=>"111011101",
  21388=>"110111011",
  21389=>"110101000",
  21390=>"010110100",
  21391=>"000000001",
  21392=>"101100110",
  21393=>"001000110",
  21394=>"101001110",
  21395=>"110111000",
  21396=>"000000000",
  21397=>"010101010",
  21398=>"001010111",
  21399=>"000100100",
  21400=>"100011010",
  21401=>"011001000",
  21402=>"101001111",
  21403=>"001011011",
  21404=>"000000010",
  21405=>"001011011",
  21406=>"010110010",
  21407=>"000100011",
  21408=>"011011000",
  21409=>"010101001",
  21410=>"100011010",
  21411=>"110011101",
  21412=>"110010000",
  21413=>"111010111",
  21414=>"101010000",
  21415=>"001110001",
  21416=>"010100000",
  21417=>"000000100",
  21418=>"110110010",
  21419=>"000011011",
  21420=>"100011011",
  21421=>"110101001",
  21422=>"001111110",
  21423=>"111110111",
  21424=>"100010110",
  21425=>"111101000",
  21426=>"001011011",
  21427=>"010000010",
  21428=>"011100000",
  21429=>"111110110",
  21430=>"011110011",
  21431=>"100111011",
  21432=>"111110101",
  21433=>"101010111",
  21434=>"011100001",
  21435=>"011101000",
  21436=>"000100100",
  21437=>"101100001",
  21438=>"000001110",
  21439=>"000111111",
  21440=>"111010110",
  21441=>"001001000",
  21442=>"100100011",
  21443=>"100100001",
  21444=>"010100001",
  21445=>"100110111",
  21446=>"001001011",
  21447=>"000111000",
  21448=>"100110000",
  21449=>"000000100",
  21450=>"110010011",
  21451=>"010011110",
  21452=>"110100111",
  21453=>"100111101",
  21454=>"000010100",
  21455=>"001010011",
  21456=>"110100110",
  21457=>"110011100",
  21458=>"110110101",
  21459=>"011100110",
  21460=>"011001111",
  21461=>"001110110",
  21462=>"100001001",
  21463=>"101000011",
  21464=>"011111101",
  21465=>"001110101",
  21466=>"001011000",
  21467=>"110011100",
  21468=>"101101011",
  21469=>"011100111",
  21470=>"011100010",
  21471=>"011100011",
  21472=>"000111111",
  21473=>"011011010",
  21474=>"101101111",
  21475=>"111010001",
  21476=>"000001111",
  21477=>"000110001",
  21478=>"001110110",
  21479=>"101011100",
  21480=>"011000100",
  21481=>"011010110",
  21482=>"101110000",
  21483=>"000110011",
  21484=>"101011111",
  21485=>"100111101",
  21486=>"010110111",
  21487=>"001110110",
  21488=>"111011111",
  21489=>"010011011",
  21490=>"000000000",
  21491=>"011000010",
  21492=>"000010010",
  21493=>"101010111",
  21494=>"110100110",
  21495=>"000001000",
  21496=>"011101001",
  21497=>"011110001",
  21498=>"110000011",
  21499=>"110011101",
  21500=>"010011111",
  21501=>"011111110",
  21502=>"010101011",
  21503=>"000011011",
  21504=>"010110101",
  21505=>"100110111",
  21506=>"110101100",
  21507=>"111111110",
  21508=>"100111001",
  21509=>"000101011",
  21510=>"110111101",
  21511=>"100110001",
  21512=>"011111111",
  21513=>"101101110",
  21514=>"110011001",
  21515=>"010001001",
  21516=>"000011000",
  21517=>"100111000",
  21518=>"100010001",
  21519=>"011111110",
  21520=>"111010000",
  21521=>"110101010",
  21522=>"111000111",
  21523=>"011101000",
  21524=>"100110111",
  21525=>"011100111",
  21526=>"000001000",
  21527=>"110000101",
  21528=>"000010110",
  21529=>"001111110",
  21530=>"100111010",
  21531=>"001010101",
  21532=>"111001010",
  21533=>"010010100",
  21534=>"011101011",
  21535=>"001000000",
  21536=>"110000011",
  21537=>"100001101",
  21538=>"100011101",
  21539=>"101000001",
  21540=>"110010011",
  21541=>"011010110",
  21542=>"001100100",
  21543=>"001101111",
  21544=>"100000001",
  21545=>"010010010",
  21546=>"001010010",
  21547=>"111001010",
  21548=>"110000110",
  21549=>"111010101",
  21550=>"000010101",
  21551=>"100100010",
  21552=>"011011011",
  21553=>"010010010",
  21554=>"110001100",
  21555=>"101001110",
  21556=>"010011101",
  21557=>"011110001",
  21558=>"010110001",
  21559=>"000111101",
  21560=>"011001101",
  21561=>"110010101",
  21562=>"010011100",
  21563=>"110000011",
  21564=>"111111100",
  21565=>"111101010",
  21566=>"101011101",
  21567=>"010101110",
  21568=>"010111000",
  21569=>"011010000",
  21570=>"100000001",
  21571=>"011100000",
  21572=>"010010010",
  21573=>"010110101",
  21574=>"011111001",
  21575=>"011111001",
  21576=>"000111100",
  21577=>"101100111",
  21578=>"100010000",
  21579=>"110011000",
  21580=>"010000011",
  21581=>"011100011",
  21582=>"000001010",
  21583=>"000010101",
  21584=>"101001000",
  21585=>"001001011",
  21586=>"111011101",
  21587=>"101110011",
  21588=>"011001100",
  21589=>"101101101",
  21590=>"100010111",
  21591=>"010010111",
  21592=>"111010111",
  21593=>"101010011",
  21594=>"010010000",
  21595=>"000100101",
  21596=>"111011111",
  21597=>"100100000",
  21598=>"100101101",
  21599=>"111100001",
  21600=>"001101010",
  21601=>"001110001",
  21602=>"001000110",
  21603=>"001001100",
  21604=>"111100101",
  21605=>"100011010",
  21606=>"110010001",
  21607=>"111000011",
  21608=>"001001111",
  21609=>"000110111",
  21610=>"010111110",
  21611=>"001100101",
  21612=>"111111010",
  21613=>"010010010",
  21614=>"010010110",
  21615=>"111001101",
  21616=>"010111101",
  21617=>"001000000",
  21618=>"101010011",
  21619=>"110010111",
  21620=>"100000111",
  21621=>"000001001",
  21622=>"100100101",
  21623=>"000011000",
  21624=>"101100110",
  21625=>"001010000",
  21626=>"111110111",
  21627=>"111100110",
  21628=>"010100000",
  21629=>"110101110",
  21630=>"111100101",
  21631=>"101011001",
  21632=>"010001100",
  21633=>"110000001",
  21634=>"110010011",
  21635=>"110101111",
  21636=>"111111010",
  21637=>"000110000",
  21638=>"011011100",
  21639=>"001110010",
  21640=>"010010111",
  21641=>"010001010",
  21642=>"111111100",
  21643=>"110111101",
  21644=>"011011000",
  21645=>"000001010",
  21646=>"111101111",
  21647=>"110110010",
  21648=>"010000110",
  21649=>"010111100",
  21650=>"011000000",
  21651=>"000010000",
  21652=>"011100101",
  21653=>"110110100",
  21654=>"001100011",
  21655=>"110101000",
  21656=>"100111111",
  21657=>"111010101",
  21658=>"000010011",
  21659=>"101111001",
  21660=>"101000000",
  21661=>"111010010",
  21662=>"111011011",
  21663=>"010010100",
  21664=>"001110011",
  21665=>"101110100",
  21666=>"011010011",
  21667=>"110010010",
  21668=>"000011111",
  21669=>"011001100",
  21670=>"001001001",
  21671=>"100010000",
  21672=>"001101110",
  21673=>"000010010",
  21674=>"001101101",
  21675=>"011111110",
  21676=>"011110001",
  21677=>"011110010",
  21678=>"001010100",
  21679=>"111101001",
  21680=>"001011001",
  21681=>"110101000",
  21682=>"111101100",
  21683=>"110101111",
  21684=>"111111101",
  21685=>"011011001",
  21686=>"110111111",
  21687=>"010100010",
  21688=>"101011000",
  21689=>"001110110",
  21690=>"011110011",
  21691=>"011110101",
  21692=>"001110101",
  21693=>"111100100",
  21694=>"001001111",
  21695=>"101111101",
  21696=>"101001011",
  21697=>"011101001",
  21698=>"001100111",
  21699=>"100110100",
  21700=>"000010100",
  21701=>"111100110",
  21702=>"000010000",
  21703=>"100011110",
  21704=>"111001111",
  21705=>"001111001",
  21706=>"110111010",
  21707=>"100101110",
  21708=>"010100010",
  21709=>"010100011",
  21710=>"001110111",
  21711=>"000000100",
  21712=>"001001101",
  21713=>"011111100",
  21714=>"010000001",
  21715=>"011010001",
  21716=>"010011010",
  21717=>"111001000",
  21718=>"100111011",
  21719=>"011001011",
  21720=>"111010000",
  21721=>"011110101",
  21722=>"111000000",
  21723=>"101001011",
  21724=>"110011100",
  21725=>"001110100",
  21726=>"110101010",
  21727=>"010100100",
  21728=>"101101001",
  21729=>"001000110",
  21730=>"111010011",
  21731=>"010100001",
  21732=>"010111101",
  21733=>"101010011",
  21734=>"000000000",
  21735=>"110101101",
  21736=>"110110000",
  21737=>"100111101",
  21738=>"100011000",
  21739=>"010010000",
  21740=>"110111001",
  21741=>"001011001",
  21742=>"000010100",
  21743=>"001010010",
  21744=>"010110110",
  21745=>"000010001",
  21746=>"110010110",
  21747=>"110110111",
  21748=>"000111011",
  21749=>"000011010",
  21750=>"111101010",
  21751=>"000110010",
  21752=>"110010111",
  21753=>"001010011",
  21754=>"110011001",
  21755=>"110101010",
  21756=>"010011110",
  21757=>"010110111",
  21758=>"010111110",
  21759=>"100111010",
  21760=>"111101010",
  21761=>"001011100",
  21762=>"101000001",
  21763=>"111100111",
  21764=>"110001010",
  21765=>"111001100",
  21766=>"101100010",
  21767=>"010100111",
  21768=>"100101001",
  21769=>"001001110",
  21770=>"001111100",
  21771=>"000111100",
  21772=>"101001101",
  21773=>"111110101",
  21774=>"100100000",
  21775=>"001011110",
  21776=>"110000001",
  21777=>"001010010",
  21778=>"110100111",
  21779=>"111100111",
  21780=>"110001000",
  21781=>"010010100",
  21782=>"001001101",
  21783=>"011100001",
  21784=>"100011001",
  21785=>"001100010",
  21786=>"010010111",
  21787=>"010011011",
  21788=>"011101110",
  21789=>"111000100",
  21790=>"011101100",
  21791=>"100001111",
  21792=>"101101101",
  21793=>"001011001",
  21794=>"001110101",
  21795=>"111111000",
  21796=>"100011110",
  21797=>"000100110",
  21798=>"100100010",
  21799=>"111000001",
  21800=>"010000001",
  21801=>"100001111",
  21802=>"111010110",
  21803=>"111000101",
  21804=>"010000110",
  21805=>"001000001",
  21806=>"110100010",
  21807=>"111110101",
  21808=>"110101101",
  21809=>"111011111",
  21810=>"010101010",
  21811=>"100110111",
  21812=>"111010000",
  21813=>"101111101",
  21814=>"011101111",
  21815=>"010100001",
  21816=>"110100011",
  21817=>"100101011",
  21818=>"000100011",
  21819=>"000011110",
  21820=>"101101111",
  21821=>"000011101",
  21822=>"011101100",
  21823=>"011010000",
  21824=>"001110111",
  21825=>"110111111",
  21826=>"000111100",
  21827=>"110110111",
  21828=>"101101101",
  21829=>"010011111",
  21830=>"101010010",
  21831=>"100101110",
  21832=>"010101011",
  21833=>"000110100",
  21834=>"011100001",
  21835=>"111010011",
  21836=>"000111000",
  21837=>"001100101",
  21838=>"001101001",
  21839=>"100111110",
  21840=>"110101111",
  21841=>"110111101",
  21842=>"000101010",
  21843=>"110111010",
  21844=>"100101110",
  21845=>"001111101",
  21846=>"000101001",
  21847=>"101011001",
  21848=>"101000111",
  21849=>"110101101",
  21850=>"100001101",
  21851=>"110001101",
  21852=>"000100110",
  21853=>"010100110",
  21854=>"011001100",
  21855=>"001101100",
  21856=>"001010111",
  21857=>"100011111",
  21858=>"010011100",
  21859=>"110011110",
  21860=>"001101001",
  21861=>"011100010",
  21862=>"110101000",
  21863=>"101010110",
  21864=>"110110011",
  21865=>"010001100",
  21866=>"111101000",
  21867=>"111100010",
  21868=>"011100111",
  21869=>"110101010",
  21870=>"001000000",
  21871=>"010011100",
  21872=>"001000010",
  21873=>"100010100",
  21874=>"100001011",
  21875=>"110011111",
  21876=>"000100100",
  21877=>"011011010",
  21878=>"011110110",
  21879=>"010110010",
  21880=>"100100000",
  21881=>"011101100",
  21882=>"100000110",
  21883=>"111011100",
  21884=>"110100010",
  21885=>"000100000",
  21886=>"011010111",
  21887=>"001101011",
  21888=>"010101011",
  21889=>"000000111",
  21890=>"001111111",
  21891=>"011001001",
  21892=>"100100011",
  21893=>"000000100",
  21894=>"111101110",
  21895=>"000101010",
  21896=>"011100101",
  21897=>"000100110",
  21898=>"101011111",
  21899=>"001000010",
  21900=>"110101101",
  21901=>"110001100",
  21902=>"010100000",
  21903=>"100110101",
  21904=>"011101111",
  21905=>"010100100",
  21906=>"000100010",
  21907=>"000000010",
  21908=>"101011111",
  21909=>"001110100",
  21910=>"000010111",
  21911=>"000111001",
  21912=>"001110100",
  21913=>"010111001",
  21914=>"110101111",
  21915=>"000001101",
  21916=>"000011100",
  21917=>"011111011",
  21918=>"111010101",
  21919=>"000011110",
  21920=>"000110111",
  21921=>"001010010",
  21922=>"000010001",
  21923=>"110100010",
  21924=>"010100000",
  21925=>"111100101",
  21926=>"011111001",
  21927=>"011110011",
  21928=>"000011001",
  21929=>"000001000",
  21930=>"011110111",
  21931=>"111001011",
  21932=>"001001000",
  21933=>"011010110",
  21934=>"100101111",
  21935=>"001101110",
  21936=>"000001111",
  21937=>"000101101",
  21938=>"110100101",
  21939=>"110011011",
  21940=>"000011010",
  21941=>"000101011",
  21942=>"101011100",
  21943=>"011000000",
  21944=>"101100100",
  21945=>"110110010",
  21946=>"010000011",
  21947=>"101101110",
  21948=>"100011000",
  21949=>"010111100",
  21950=>"101011100",
  21951=>"111110010",
  21952=>"111100110",
  21953=>"111111010",
  21954=>"111000001",
  21955=>"000100101",
  21956=>"000000101",
  21957=>"111000101",
  21958=>"010010111",
  21959=>"101001000",
  21960=>"000001100",
  21961=>"001101100",
  21962=>"010100000",
  21963=>"000101011",
  21964=>"010010001",
  21965=>"101101100",
  21966=>"010101010",
  21967=>"111110001",
  21968=>"000100110",
  21969=>"011111001",
  21970=>"100001101",
  21971=>"001011010",
  21972=>"000111000",
  21973=>"001000010",
  21974=>"011111110",
  21975=>"111111101",
  21976=>"011101000",
  21977=>"111111000",
  21978=>"001101011",
  21979=>"000111111",
  21980=>"011000101",
  21981=>"010001100",
  21982=>"111100010",
  21983=>"011011100",
  21984=>"011110000",
  21985=>"001011001",
  21986=>"111110110",
  21987=>"110000110",
  21988=>"000100110",
  21989=>"010011101",
  21990=>"001011011",
  21991=>"001001000",
  21992=>"110100001",
  21993=>"000101110",
  21994=>"000011100",
  21995=>"110011010",
  21996=>"010110011",
  21997=>"011111100",
  21998=>"010011110",
  21999=>"000011101",
  22000=>"010011101",
  22001=>"010101100",
  22002=>"111001010",
  22003=>"011101010",
  22004=>"000010000",
  22005=>"011101000",
  22006=>"111111001",
  22007=>"010001001",
  22008=>"110001101",
  22009=>"110111110",
  22010=>"000001110",
  22011=>"000110111",
  22012=>"001101010",
  22013=>"100001000",
  22014=>"110000001",
  22015=>"110111000",
  22016=>"101100000",
  22017=>"011001100",
  22018=>"010100010",
  22019=>"010011010",
  22020=>"010101110",
  22021=>"001000100",
  22022=>"010001111",
  22023=>"010100100",
  22024=>"110001110",
  22025=>"111011000",
  22026=>"011101100",
  22027=>"010011010",
  22028=>"100001100",
  22029=>"111111000",
  22030=>"000001111",
  22031=>"010111101",
  22032=>"011110101",
  22033=>"010001001",
  22034=>"010100010",
  22035=>"110000001",
  22036=>"010011001",
  22037=>"110110010",
  22038=>"001111111",
  22039=>"111101100",
  22040=>"111110100",
  22041=>"011010101",
  22042=>"001001011",
  22043=>"110000101",
  22044=>"111000100",
  22045=>"100111001",
  22046=>"001000011",
  22047=>"101001001",
  22048=>"100100001",
  22049=>"111010110",
  22050=>"001110011",
  22051=>"001010000",
  22052=>"000011101",
  22053=>"010011010",
  22054=>"100010110",
  22055=>"000111011",
  22056=>"011111000",
  22057=>"101111010",
  22058=>"110100011",
  22059=>"111100010",
  22060=>"110111110",
  22061=>"111000001",
  22062=>"110110100",
  22063=>"100110011",
  22064=>"100010001",
  22065=>"110011010",
  22066=>"000001101",
  22067=>"100011111",
  22068=>"101100101",
  22069=>"101111001",
  22070=>"111000101",
  22071=>"011110000",
  22072=>"100111010",
  22073=>"110110111",
  22074=>"101011000",
  22075=>"011100110",
  22076=>"011010100",
  22077=>"010000010",
  22078=>"100101111",
  22079=>"101100011",
  22080=>"010010000",
  22081=>"010011100",
  22082=>"111000001",
  22083=>"111110110",
  22084=>"000000001",
  22085=>"001010001",
  22086=>"000111001",
  22087=>"111111010",
  22088=>"001101000",
  22089=>"111101000",
  22090=>"001100000",
  22091=>"001011010",
  22092=>"101011111",
  22093=>"001100001",
  22094=>"111100111",
  22095=>"100101100",
  22096=>"000010001",
  22097=>"010100000",
  22098=>"000001110",
  22099=>"100001001",
  22100=>"101110000",
  22101=>"111000000",
  22102=>"101101101",
  22103=>"000111111",
  22104=>"111111110",
  22105=>"011000000",
  22106=>"111100101",
  22107=>"101100101",
  22108=>"100101001",
  22109=>"010010000",
  22110=>"100010010",
  22111=>"001110001",
  22112=>"110001101",
  22113=>"111010000",
  22114=>"100010110",
  22115=>"000000111",
  22116=>"101001011",
  22117=>"001100001",
  22118=>"100100010",
  22119=>"111000010",
  22120=>"010101101",
  22121=>"101011010",
  22122=>"001111101",
  22123=>"000000000",
  22124=>"111111111",
  22125=>"111101111",
  22126=>"010011110",
  22127=>"110000110",
  22128=>"001110010",
  22129=>"011011001",
  22130=>"110110001",
  22131=>"110100110",
  22132=>"101010010",
  22133=>"000100000",
  22134=>"010001000",
  22135=>"010110000",
  22136=>"110111001",
  22137=>"111100101",
  22138=>"100011011",
  22139=>"011101101",
  22140=>"110001000",
  22141=>"110011111",
  22142=>"010100000",
  22143=>"100011011",
  22144=>"011001100",
  22145=>"110100000",
  22146=>"011101100",
  22147=>"111101100",
  22148=>"010101111",
  22149=>"111000110",
  22150=>"111111101",
  22151=>"000101111",
  22152=>"011001011",
  22153=>"011010111",
  22154=>"110000010",
  22155=>"110001000",
  22156=>"111101001",
  22157=>"000110110",
  22158=>"110010000",
  22159=>"101000111",
  22160=>"111111111",
  22161=>"100000101",
  22162=>"100100000",
  22163=>"001111000",
  22164=>"011100010",
  22165=>"000001010",
  22166=>"101011001",
  22167=>"111001000",
  22168=>"000110001",
  22169=>"100000100",
  22170=>"101000101",
  22171=>"101111001",
  22172=>"000000000",
  22173=>"111101011",
  22174=>"110001000",
  22175=>"001111010",
  22176=>"000110011",
  22177=>"100111000",
  22178=>"100100000",
  22179=>"011010111",
  22180=>"001001001",
  22181=>"001000101",
  22182=>"111110100",
  22183=>"111101001",
  22184=>"011110000",
  22185=>"000101001",
  22186=>"000001000",
  22187=>"110111101",
  22188=>"001110101",
  22189=>"110100010",
  22190=>"111110001",
  22191=>"101101010",
  22192=>"100000010",
  22193=>"100001111",
  22194=>"111111010",
  22195=>"001110000",
  22196=>"010001001",
  22197=>"101001000",
  22198=>"110111101",
  22199=>"000100011",
  22200=>"110010001",
  22201=>"100101111",
  22202=>"000111010",
  22203=>"011011000",
  22204=>"111101101",
  22205=>"101011001",
  22206=>"111111100",
  22207=>"011111000",
  22208=>"110000111",
  22209=>"110111111",
  22210=>"000000101",
  22211=>"001111000",
  22212=>"000000010",
  22213=>"101001110",
  22214=>"010100100",
  22215=>"101111011",
  22216=>"100111110",
  22217=>"110110010",
  22218=>"100010001",
  22219=>"001111010",
  22220=>"010100101",
  22221=>"000001101",
  22222=>"011010110",
  22223=>"011110001",
  22224=>"101000010",
  22225=>"010111001",
  22226=>"010100101",
  22227=>"011101000",
  22228=>"011111101",
  22229=>"111000001",
  22230=>"011011101",
  22231=>"010001010",
  22232=>"111000001",
  22233=>"101000000",
  22234=>"101110111",
  22235=>"001000111",
  22236=>"010000101",
  22237=>"000000110",
  22238=>"100000100",
  22239=>"001000001",
  22240=>"100001010",
  22241=>"111001111",
  22242=>"110010001",
  22243=>"110011100",
  22244=>"000011000",
  22245=>"010111011",
  22246=>"100110100",
  22247=>"111100000",
  22248=>"111111011",
  22249=>"011001010",
  22250=>"110100000",
  22251=>"101000010",
  22252=>"101101100",
  22253=>"011101011",
  22254=>"000111101",
  22255=>"001001011",
  22256=>"000011011",
  22257=>"101100101",
  22258=>"010010110",
  22259=>"001000010",
  22260=>"111101110",
  22261=>"111110101",
  22262=>"011000100",
  22263=>"001000011",
  22264=>"010011101",
  22265=>"001101000",
  22266=>"100101111",
  22267=>"010110001",
  22268=>"000100110",
  22269=>"101101010",
  22270=>"111001110",
  22271=>"001101101",
  22272=>"000001011",
  22273=>"011011001",
  22274=>"101001100",
  22275=>"001101001",
  22276=>"011111100",
  22277=>"110000010",
  22278=>"101011100",
  22279=>"001010000",
  22280=>"001100100",
  22281=>"000101110",
  22282=>"001000011",
  22283=>"101000110",
  22284=>"010111101",
  22285=>"100110000",
  22286=>"110100011",
  22287=>"000000101",
  22288=>"000010010",
  22289=>"100101000",
  22290=>"110011110",
  22291=>"110011100",
  22292=>"010011100",
  22293=>"110101100",
  22294=>"111110000",
  22295=>"110000000",
  22296=>"011000001",
  22297=>"101111111",
  22298=>"001101011",
  22299=>"000100111",
  22300=>"000110110",
  22301=>"110000011",
  22302=>"110111110",
  22303=>"001101111",
  22304=>"011110110",
  22305=>"010010001",
  22306=>"000011111",
  22307=>"101000001",
  22308=>"111100001",
  22309=>"010111011",
  22310=>"110111000",
  22311=>"100010110",
  22312=>"000011000",
  22313=>"111110001",
  22314=>"111001111",
  22315=>"110111000",
  22316=>"100000100",
  22317=>"100000010",
  22318=>"000111011",
  22319=>"111110101",
  22320=>"111010101",
  22321=>"101011001",
  22322=>"100110011",
  22323=>"001001100",
  22324=>"000011010",
  22325=>"010111001",
  22326=>"000111110",
  22327=>"011111110",
  22328=>"000000100",
  22329=>"110010011",
  22330=>"011010101",
  22331=>"001111000",
  22332=>"111100110",
  22333=>"001000111",
  22334=>"100110001",
  22335=>"011001000",
  22336=>"101100110",
  22337=>"011010001",
  22338=>"011010011",
  22339=>"000011010",
  22340=>"001000001",
  22341=>"111100101",
  22342=>"001001011",
  22343=>"000011000",
  22344=>"111100010",
  22345=>"111110001",
  22346=>"011100011",
  22347=>"111010101",
  22348=>"101010010",
  22349=>"000000000",
  22350=>"011011111",
  22351=>"000000110",
  22352=>"011101010",
  22353=>"001010000",
  22354=>"111010000",
  22355=>"110100110",
  22356=>"111011010",
  22357=>"101110110",
  22358=>"100010110",
  22359=>"110001011",
  22360=>"110100101",
  22361=>"010011101",
  22362=>"010100101",
  22363=>"000100101",
  22364=>"001001111",
  22365=>"110010111",
  22366=>"000111000",
  22367=>"001101000",
  22368=>"001000110",
  22369=>"010110110",
  22370=>"110001100",
  22371=>"011111000",
  22372=>"010110110",
  22373=>"011001100",
  22374=>"100101001",
  22375=>"011101011",
  22376=>"010101010",
  22377=>"101010111",
  22378=>"000100010",
  22379=>"011101101",
  22380=>"110101000",
  22381=>"110100100",
  22382=>"110010110",
  22383=>"010011110",
  22384=>"111011001",
  22385=>"001110110",
  22386=>"100011010",
  22387=>"001101010",
  22388=>"101010001",
  22389=>"100001111",
  22390=>"010001010",
  22391=>"001111000",
  22392=>"010110011",
  22393=>"100001110",
  22394=>"001011001",
  22395=>"010110111",
  22396=>"011010011",
  22397=>"010001000",
  22398=>"110010111",
  22399=>"010010101",
  22400=>"101010010",
  22401=>"011110100",
  22402=>"000001101",
  22403=>"101000101",
  22404=>"110100101",
  22405=>"100000010",
  22406=>"000101011",
  22407=>"001101000",
  22408=>"110110101",
  22409=>"111101000",
  22410=>"111010111",
  22411=>"001111100",
  22412=>"110001000",
  22413=>"010001001",
  22414=>"010101110",
  22415=>"001000111",
  22416=>"110101010",
  22417=>"100010100",
  22418=>"011110000",
  22419=>"110010100",
  22420=>"011000111",
  22421=>"111001110",
  22422=>"001011110",
  22423=>"110001110",
  22424=>"100000100",
  22425=>"000101010",
  22426=>"101101011",
  22427=>"011101100",
  22428=>"010000111",
  22429=>"010010011",
  22430=>"100101000",
  22431=>"011000110",
  22432=>"001101001",
  22433=>"111011101",
  22434=>"001101010",
  22435=>"000000100",
  22436=>"101000111",
  22437=>"001110100",
  22438=>"001110111",
  22439=>"000110100",
  22440=>"001001000",
  22441=>"000011011",
  22442=>"110101101",
  22443=>"010001001",
  22444=>"010010101",
  22445=>"111100101",
  22446=>"011001001",
  22447=>"100001110",
  22448=>"111111000",
  22449=>"100010010",
  22450=>"010001110",
  22451=>"110000011",
  22452=>"100110101",
  22453=>"100110000",
  22454=>"000111000",
  22455=>"000010011",
  22456=>"110100100",
  22457=>"100001100",
  22458=>"100101111",
  22459=>"101111100",
  22460=>"000000011",
  22461=>"001110010",
  22462=>"111101001",
  22463=>"000000000",
  22464=>"000000011",
  22465=>"010111110",
  22466=>"111001010",
  22467=>"000100011",
  22468=>"110110001",
  22469=>"111010110",
  22470=>"100010001",
  22471=>"000111011",
  22472=>"001000100",
  22473=>"000110111",
  22474=>"000100100",
  22475=>"101010001",
  22476=>"100111000",
  22477=>"100000111",
  22478=>"111100010",
  22479=>"110101100",
  22480=>"011101111",
  22481=>"001101100",
  22482=>"001001101",
  22483=>"100011100",
  22484=>"011010011",
  22485=>"101101111",
  22486=>"000100101",
  22487=>"111100100",
  22488=>"011111100",
  22489=>"001001000",
  22490=>"000110111",
  22491=>"100111000",
  22492=>"001001100",
  22493=>"100100001",
  22494=>"010111100",
  22495=>"101111111",
  22496=>"111110101",
  22497=>"101110000",
  22498=>"101001100",
  22499=>"010001000",
  22500=>"011110000",
  22501=>"111011000",
  22502=>"010101100",
  22503=>"111010000",
  22504=>"011001100",
  22505=>"101100101",
  22506=>"100011100",
  22507=>"101000110",
  22508=>"111111001",
  22509=>"010010010",
  22510=>"000111100",
  22511=>"111000101",
  22512=>"101110000",
  22513=>"111001001",
  22514=>"111001001",
  22515=>"000101000",
  22516=>"101101001",
  22517=>"011111100",
  22518=>"001010000",
  22519=>"110000100",
  22520=>"011110110",
  22521=>"110111000",
  22522=>"101101100",
  22523=>"010110110",
  22524=>"110001101",
  22525=>"011001000",
  22526=>"110101001",
  22527=>"110010111",
  22528=>"001101010",
  22529=>"010010000",
  22530=>"001110001",
  22531=>"010010110",
  22532=>"110001110",
  22533=>"101011101",
  22534=>"110001101",
  22535=>"100010011",
  22536=>"000101100",
  22537=>"110110110",
  22538=>"100000100",
  22539=>"110001111",
  22540=>"101101110",
  22541=>"100001000",
  22542=>"111010001",
  22543=>"101110110",
  22544=>"111110010",
  22545=>"001011101",
  22546=>"111010101",
  22547=>"110000001",
  22548=>"000111101",
  22549=>"101010011",
  22550=>"011010011",
  22551=>"111100000",
  22552=>"110010001",
  22553=>"011100001",
  22554=>"011001111",
  22555=>"011011000",
  22556=>"101000011",
  22557=>"100111000",
  22558=>"100000001",
  22559=>"111110010",
  22560=>"111000011",
  22561=>"010011011",
  22562=>"000001000",
  22563=>"111101001",
  22564=>"111011010",
  22565=>"100010110",
  22566=>"000100100",
  22567=>"000011110",
  22568=>"000001010",
  22569=>"100110001",
  22570=>"111100001",
  22571=>"111111101",
  22572=>"011001000",
  22573=>"111001101",
  22574=>"001100000",
  22575=>"001011110",
  22576=>"110100111",
  22577=>"001001101",
  22578=>"111011110",
  22579=>"010111111",
  22580=>"010101001",
  22581=>"000111010",
  22582=>"110001011",
  22583=>"111010000",
  22584=>"101101000",
  22585=>"110111110",
  22586=>"111110011",
  22587=>"100010110",
  22588=>"011110010",
  22589=>"000000111",
  22590=>"000110110",
  22591=>"001011010",
  22592=>"000101001",
  22593=>"101001111",
  22594=>"110101101",
  22595=>"100100001",
  22596=>"101010010",
  22597=>"001111011",
  22598=>"010111111",
  22599=>"101100111",
  22600=>"110111110",
  22601=>"010110001",
  22602=>"100101011",
  22603=>"000000111",
  22604=>"000110100",
  22605=>"011101011",
  22606=>"101001001",
  22607=>"111100011",
  22608=>"111111111",
  22609=>"010001100",
  22610=>"111101011",
  22611=>"000011100",
  22612=>"111000100",
  22613=>"000000111",
  22614=>"000111010",
  22615=>"100100100",
  22616=>"111000100",
  22617=>"100010110",
  22618=>"011001101",
  22619=>"000010000",
  22620=>"011010001",
  22621=>"110100111",
  22622=>"110010001",
  22623=>"001000001",
  22624=>"011101100",
  22625=>"101100000",
  22626=>"111011010",
  22627=>"010011010",
  22628=>"100100101",
  22629=>"010011100",
  22630=>"001001111",
  22631=>"001100001",
  22632=>"110101100",
  22633=>"001001010",
  22634=>"001101010",
  22635=>"100010100",
  22636=>"011100111",
  22637=>"001100100",
  22638=>"011011110",
  22639=>"100110111",
  22640=>"001001001",
  22641=>"111001111",
  22642=>"001110001",
  22643=>"000010101",
  22644=>"010110100",
  22645=>"001000101",
  22646=>"101110110",
  22647=>"000000001",
  22648=>"011101100",
  22649=>"000000011",
  22650=>"110111100",
  22651=>"100110000",
  22652=>"110001011",
  22653=>"100010100",
  22654=>"000100110",
  22655=>"110010111",
  22656=>"000110001",
  22657=>"000010010",
  22658=>"111101000",
  22659=>"001101111",
  22660=>"010110001",
  22661=>"001110111",
  22662=>"010100010",
  22663=>"100111111",
  22664=>"011100010",
  22665=>"101011001",
  22666=>"100101100",
  22667=>"011010110",
  22668=>"000011110",
  22669=>"111000111",
  22670=>"111101100",
  22671=>"110000001",
  22672=>"000010010",
  22673=>"010101011",
  22674=>"000100101",
  22675=>"000000110",
  22676=>"110001111",
  22677=>"001111100",
  22678=>"001001101",
  22679=>"100010001",
  22680=>"110001000",
  22681=>"000000110",
  22682=>"101111011",
  22683=>"110001010",
  22684=>"010000100",
  22685=>"100101110",
  22686=>"101010111",
  22687=>"101101011",
  22688=>"110000011",
  22689=>"110110110",
  22690=>"111100010",
  22691=>"110101111",
  22692=>"110010000",
  22693=>"101101111",
  22694=>"110111000",
  22695=>"111010100",
  22696=>"011001001",
  22697=>"110010010",
  22698=>"010000010",
  22699=>"110111000",
  22700=>"011000101",
  22701=>"111110000",
  22702=>"100101100",
  22703=>"111110010",
  22704=>"111101001",
  22705=>"001110111",
  22706=>"001100111",
  22707=>"111110000",
  22708=>"000101011",
  22709=>"110001101",
  22710=>"111101100",
  22711=>"110010011",
  22712=>"011000000",
  22713=>"110011100",
  22714=>"111111011",
  22715=>"010011110",
  22716=>"101101010",
  22717=>"111110110",
  22718=>"011100000",
  22719=>"011000101",
  22720=>"110100111",
  22721=>"100101100",
  22722=>"000000011",
  22723=>"110001001",
  22724=>"011111110",
  22725=>"100110001",
  22726=>"011110101",
  22727=>"011010101",
  22728=>"111000000",
  22729=>"001001110",
  22730=>"100111001",
  22731=>"001111111",
  22732=>"001010110",
  22733=>"100101010",
  22734=>"010100010",
  22735=>"111111100",
  22736=>"100100101",
  22737=>"101110100",
  22738=>"000101011",
  22739=>"011100101",
  22740=>"001010111",
  22741=>"101000110",
  22742=>"100001000",
  22743=>"000001110",
  22744=>"001101011",
  22745=>"001010101",
  22746=>"001011111",
  22747=>"011010000",
  22748=>"100101000",
  22749=>"110001110",
  22750=>"100110001",
  22751=>"010001000",
  22752=>"110101000",
  22753=>"011100010",
  22754=>"010001110",
  22755=>"000101101",
  22756=>"110111100",
  22757=>"101101011",
  22758=>"000000010",
  22759=>"111110011",
  22760=>"100000001",
  22761=>"101101000",
  22762=>"000111101",
  22763=>"000000001",
  22764=>"111100011",
  22765=>"100001000",
  22766=>"010111001",
  22767=>"100011101",
  22768=>"111111110",
  22769=>"010000010",
  22770=>"010100100",
  22771=>"101000111",
  22772=>"001000111",
  22773=>"000000101",
  22774=>"001110000",
  22775=>"111101000",
  22776=>"101000110",
  22777=>"100011000",
  22778=>"010010101",
  22779=>"111111110",
  22780=>"101011110",
  22781=>"000100101",
  22782=>"000100100",
  22783=>"010110100",
  22784=>"110100010",
  22785=>"001011101",
  22786=>"111001111",
  22787=>"101011010",
  22788=>"001101010",
  22789=>"001000011",
  22790=>"101101111",
  22791=>"110110101",
  22792=>"001010110",
  22793=>"011011111",
  22794=>"011111001",
  22795=>"010011011",
  22796=>"000011010",
  22797=>"001101100",
  22798=>"100111101",
  22799=>"100001011",
  22800=>"110010001",
  22801=>"101101111",
  22802=>"111101101",
  22803=>"000000010",
  22804=>"110101011",
  22805=>"000101101",
  22806=>"010110001",
  22807=>"111110011",
  22808=>"010101001",
  22809=>"110100110",
  22810=>"000010010",
  22811=>"111111011",
  22812=>"111011111",
  22813=>"111100101",
  22814=>"011000010",
  22815=>"100001101",
  22816=>"000000110",
  22817=>"110100100",
  22818=>"010010101",
  22819=>"110101000",
  22820=>"001101001",
  22821=>"010111111",
  22822=>"000000000",
  22823=>"001010001",
  22824=>"111101111",
  22825=>"110000001",
  22826=>"011111110",
  22827=>"011110001",
  22828=>"011000111",
  22829=>"111000000",
  22830=>"001101010",
  22831=>"001111000",
  22832=>"111001010",
  22833=>"100100110",
  22834=>"010001101",
  22835=>"011111010",
  22836=>"001010110",
  22837=>"110100100",
  22838=>"001011000",
  22839=>"110110001",
  22840=>"100101011",
  22841=>"010110111",
  22842=>"101111101",
  22843=>"011010000",
  22844=>"111010000",
  22845=>"000000000",
  22846=>"100000001",
  22847=>"110101001",
  22848=>"110000101",
  22849=>"101111000",
  22850=>"000010000",
  22851=>"011010001",
  22852=>"011100100",
  22853=>"110101001",
  22854=>"010000000",
  22855=>"100001000",
  22856=>"001010100",
  22857=>"101111101",
  22858=>"010001010",
  22859=>"111101011",
  22860=>"111110101",
  22861=>"010011001",
  22862=>"100010001",
  22863=>"111111010",
  22864=>"100100110",
  22865=>"110011100",
  22866=>"001101011",
  22867=>"111110101",
  22868=>"110001001",
  22869=>"101001101",
  22870=>"100000011",
  22871=>"011111110",
  22872=>"001011110",
  22873=>"000011101",
  22874=>"001101111",
  22875=>"100110010",
  22876=>"001000100",
  22877=>"001000100",
  22878=>"010101001",
  22879=>"000110100",
  22880=>"111011110",
  22881=>"110001100",
  22882=>"000011101",
  22883=>"101010110",
  22884=>"110110001",
  22885=>"011010111",
  22886=>"111111000",
  22887=>"100110011",
  22888=>"010010101",
  22889=>"010011000",
  22890=>"001011110",
  22891=>"100011111",
  22892=>"101001100",
  22893=>"111111001",
  22894=>"110000001",
  22895=>"110001011",
  22896=>"100000110",
  22897=>"111010100",
  22898=>"111111000",
  22899=>"100101010",
  22900=>"001101000",
  22901=>"011000001",
  22902=>"000000011",
  22903=>"000001010",
  22904=>"110000111",
  22905=>"000000010",
  22906=>"000000001",
  22907=>"101100000",
  22908=>"110100101",
  22909=>"011101100",
  22910=>"011100000",
  22911=>"110100100",
  22912=>"110000000",
  22913=>"000000101",
  22914=>"011000011",
  22915=>"010110000",
  22916=>"001111111",
  22917=>"011110111",
  22918=>"101110101",
  22919=>"100100010",
  22920=>"111111101",
  22921=>"110111110",
  22922=>"100101000",
  22923=>"111011011",
  22924=>"000100011",
  22925=>"111001100",
  22926=>"000010111",
  22927=>"000000101",
  22928=>"101001110",
  22929=>"100100001",
  22930=>"101100011",
  22931=>"101111000",
  22932=>"011001101",
  22933=>"110101110",
  22934=>"010110010",
  22935=>"010011000",
  22936=>"100111010",
  22937=>"110110001",
  22938=>"001001101",
  22939=>"001000000",
  22940=>"101000000",
  22941=>"000101110",
  22942=>"001111101",
  22943=>"011010010",
  22944=>"000110101",
  22945=>"010101010",
  22946=>"110110100",
  22947=>"111010011",
  22948=>"011001101",
  22949=>"101000100",
  22950=>"111010011",
  22951=>"010100101",
  22952=>"111010100",
  22953=>"000110101",
  22954=>"100100100",
  22955=>"010100100",
  22956=>"100110010",
  22957=>"010111000",
  22958=>"000010000",
  22959=>"001110010",
  22960=>"101111100",
  22961=>"011011110",
  22962=>"001111111",
  22963=>"010101000",
  22964=>"110011111",
  22965=>"101110111",
  22966=>"100010000",
  22967=>"110101010",
  22968=>"011101110",
  22969=>"111010111",
  22970=>"110011110",
  22971=>"111110011",
  22972=>"100110000",
  22973=>"110110010",
  22974=>"101000000",
  22975=>"001100001",
  22976=>"111011000",
  22977=>"100100000",
  22978=>"101010110",
  22979=>"100110010",
  22980=>"101100100",
  22981=>"011011011",
  22982=>"011011101",
  22983=>"100011011",
  22984=>"001001110",
  22985=>"111111000",
  22986=>"011100011",
  22987=>"000101100",
  22988=>"100101111",
  22989=>"000101101",
  22990=>"101101101",
  22991=>"000111111",
  22992=>"101010001",
  22993=>"010111010",
  22994=>"011110000",
  22995=>"111101100",
  22996=>"110010111",
  22997=>"101010011",
  22998=>"010110000",
  22999=>"001100010",
  23000=>"010011100",
  23001=>"101100111",
  23002=>"100011100",
  23003=>"011000100",
  23004=>"010001111",
  23005=>"110111000",
  23006=>"111101001",
  23007=>"101001011",
  23008=>"101001100",
  23009=>"101011111",
  23010=>"000000100",
  23011=>"010000011",
  23012=>"111001011",
  23013=>"100010010",
  23014=>"110111100",
  23015=>"001101000",
  23016=>"111000110",
  23017=>"010101011",
  23018=>"110110111",
  23019=>"100000101",
  23020=>"000100110",
  23021=>"110101111",
  23022=>"011101001",
  23023=>"101100100",
  23024=>"001011100",
  23025=>"000001001",
  23026=>"110011000",
  23027=>"000000010",
  23028=>"001111100",
  23029=>"000100001",
  23030=>"100100011",
  23031=>"100100011",
  23032=>"101100000",
  23033=>"000001010",
  23034=>"101011010",
  23035=>"011101100",
  23036=>"110011101",
  23037=>"001001101",
  23038=>"100111110",
  23039=>"001001001",
  23040=>"001101111",
  23041=>"000001000",
  23042=>"111000111",
  23043=>"100000000",
  23044=>"101000110",
  23045=>"010110110",
  23046=>"010101101",
  23047=>"110000101",
  23048=>"100001101",
  23049=>"000101011",
  23050=>"010111111",
  23051=>"111110111",
  23052=>"111011111",
  23053=>"001000011",
  23054=>"011110101",
  23055=>"101000100",
  23056=>"100110011",
  23057=>"111100000",
  23058=>"111101010",
  23059=>"011101110",
  23060=>"001111100",
  23061=>"010011100",
  23062=>"110111000",
  23063=>"100010010",
  23064=>"101101000",
  23065=>"100000001",
  23066=>"000000001",
  23067=>"110101101",
  23068=>"001100000",
  23069=>"010011000",
  23070=>"011000000",
  23071=>"111001010",
  23072=>"110000000",
  23073=>"000001000",
  23074=>"010110010",
  23075=>"000011101",
  23076=>"101001010",
  23077=>"011111110",
  23078=>"110000001",
  23079=>"000100101",
  23080=>"110010000",
  23081=>"001011101",
  23082=>"100100100",
  23083=>"000101001",
  23084=>"110010111",
  23085=>"111100011",
  23086=>"101110100",
  23087=>"101111110",
  23088=>"110001110",
  23089=>"101011000",
  23090=>"000010101",
  23091=>"101011100",
  23092=>"011100011",
  23093=>"011110101",
  23094=>"110100110",
  23095=>"011100111",
  23096=>"100000010",
  23097=>"010010101",
  23098=>"011000111",
  23099=>"100011101",
  23100=>"001010101",
  23101=>"110110101",
  23102=>"110110100",
  23103=>"100001001",
  23104=>"111111110",
  23105=>"001110110",
  23106=>"000010101",
  23107=>"001001101",
  23108=>"110010100",
  23109=>"111110000",
  23110=>"110001001",
  23111=>"000110111",
  23112=>"011011000",
  23113=>"011000000",
  23114=>"011010100",
  23115=>"100000011",
  23116=>"110011000",
  23117=>"111000100",
  23118=>"001011000",
  23119=>"100001111",
  23120=>"100101011",
  23121=>"110110000",
  23122=>"001100010",
  23123=>"111111101",
  23124=>"111110101",
  23125=>"010100000",
  23126=>"100101010",
  23127=>"110111100",
  23128=>"101111101",
  23129=>"001111110",
  23130=>"101101001",
  23131=>"001001011",
  23132=>"001010000",
  23133=>"001010010",
  23134=>"100101010",
  23135=>"110101011",
  23136=>"110010010",
  23137=>"010110001",
  23138=>"010010110",
  23139=>"001010000",
  23140=>"111001001",
  23141=>"111001110",
  23142=>"101011111",
  23143=>"001010010",
  23144=>"000001000",
  23145=>"100001100",
  23146=>"110000110",
  23147=>"110011111",
  23148=>"110111011",
  23149=>"111101001",
  23150=>"101101101",
  23151=>"100010111",
  23152=>"000000100",
  23153=>"000001001",
  23154=>"110100101",
  23155=>"010001101",
  23156=>"101001111",
  23157=>"010011001",
  23158=>"011001000",
  23159=>"101010110",
  23160=>"110000011",
  23161=>"011100100",
  23162=>"111001100",
  23163=>"101000010",
  23164=>"011001110",
  23165=>"011100111",
  23166=>"100101011",
  23167=>"110000010",
  23168=>"100011110",
  23169=>"001010001",
  23170=>"010000000",
  23171=>"010100110",
  23172=>"111000101",
  23173=>"010010111",
  23174=>"100111100",
  23175=>"100011011",
  23176=>"011100101",
  23177=>"100000110",
  23178=>"000101110",
  23179=>"110101011",
  23180=>"001011001",
  23181=>"111100000",
  23182=>"110001010",
  23183=>"111101111",
  23184=>"010010010",
  23185=>"010110011",
  23186=>"101101111",
  23187=>"111011000",
  23188=>"001111010",
  23189=>"001011111",
  23190=>"011000100",
  23191=>"111101110",
  23192=>"101000110",
  23193=>"001001000",
  23194=>"100010111",
  23195=>"111101100",
  23196=>"010001010",
  23197=>"010010010",
  23198=>"110011101",
  23199=>"000100110",
  23200=>"110110001",
  23201=>"101011000",
  23202=>"011101011",
  23203=>"000111011",
  23204=>"011001101",
  23205=>"110010110",
  23206=>"010000000",
  23207=>"001100000",
  23208=>"000001001",
  23209=>"011101101",
  23210=>"010100001",
  23211=>"010001001",
  23212=>"010000100",
  23213=>"011110111",
  23214=>"111000010",
  23215=>"001001011",
  23216=>"001111000",
  23217=>"011101010",
  23218=>"100000101",
  23219=>"110010000",
  23220=>"000010100",
  23221=>"110000011",
  23222=>"011101100",
  23223=>"000111111",
  23224=>"111010011",
  23225=>"010011011",
  23226=>"010111000",
  23227=>"100001100",
  23228=>"011101001",
  23229=>"000100001",
  23230=>"100000000",
  23231=>"000010110",
  23232=>"010110011",
  23233=>"010010011",
  23234=>"101100000",
  23235=>"001101100",
  23236=>"010000011",
  23237=>"111001001",
  23238=>"011101010",
  23239=>"100111110",
  23240=>"100110010",
  23241=>"111100010",
  23242=>"001000010",
  23243=>"101000111",
  23244=>"011110011",
  23245=>"101011010",
  23246=>"001001001",
  23247=>"000000110",
  23248=>"000111010",
  23249=>"110100011",
  23250=>"101111010",
  23251=>"111110111",
  23252=>"101101100",
  23253=>"010111111",
  23254=>"110111101",
  23255=>"101110100",
  23256=>"000110011",
  23257=>"100000011",
  23258=>"010000111",
  23259=>"111001101",
  23260=>"000000000",
  23261=>"100101101",
  23262=>"001001101",
  23263=>"111000000",
  23264=>"110111001",
  23265=>"100100110",
  23266=>"100010001",
  23267=>"010010111",
  23268=>"000001001",
  23269=>"011101001",
  23270=>"110011000",
  23271=>"111001011",
  23272=>"111101000",
  23273=>"011000000",
  23274=>"101000101",
  23275=>"010011111",
  23276=>"011101010",
  23277=>"100000110",
  23278=>"011111110",
  23279=>"110100001",
  23280=>"001001010",
  23281=>"101000000",
  23282=>"010100001",
  23283=>"111011110",
  23284=>"101010000",
  23285=>"000110001",
  23286=>"011111000",
  23287=>"000100000",
  23288=>"000000100",
  23289=>"101110000",
  23290=>"110001010",
  23291=>"101100110",
  23292=>"000001010",
  23293=>"000000100",
  23294=>"011101100",
  23295=>"110000000",
  23296=>"110001001",
  23297=>"101101101",
  23298=>"111001001",
  23299=>"111010010",
  23300=>"011111110",
  23301=>"010111111",
  23302=>"111101001",
  23303=>"111111111",
  23304=>"010100000",
  23305=>"011110000",
  23306=>"001110110",
  23307=>"000011111",
  23308=>"011111100",
  23309=>"100011001",
  23310=>"000011110",
  23311=>"010101110",
  23312=>"000000011",
  23313=>"010100110",
  23314=>"011111111",
  23315=>"100011110",
  23316=>"101101111",
  23317=>"010011011",
  23318=>"111010111",
  23319=>"011111101",
  23320=>"000000001",
  23321=>"001110011",
  23322=>"101111111",
  23323=>"010000101",
  23324=>"100111001",
  23325=>"111100111",
  23326=>"100010110",
  23327=>"111000011",
  23328=>"000010110",
  23329=>"001110001",
  23330=>"110001100",
  23331=>"101110110",
  23332=>"111011011",
  23333=>"010101000",
  23334=>"100100011",
  23335=>"111110111",
  23336=>"010000001",
  23337=>"110000000",
  23338=>"100011110",
  23339=>"011101011",
  23340=>"000001111",
  23341=>"100011100",
  23342=>"001001010",
  23343=>"100110110",
  23344=>"000100010",
  23345=>"101000110",
  23346=>"100110001",
  23347=>"011111011",
  23348=>"001111000",
  23349=>"110011010",
  23350=>"110001011",
  23351=>"111101101",
  23352=>"001101100",
  23353=>"111101111",
  23354=>"101100101",
  23355=>"000010001",
  23356=>"001110000",
  23357=>"001100001",
  23358=>"111110100",
  23359=>"011010001",
  23360=>"000101110",
  23361=>"100000011",
  23362=>"010101011",
  23363=>"110100110",
  23364=>"000010101",
  23365=>"011111000",
  23366=>"111101111",
  23367=>"100011000",
  23368=>"101100000",
  23369=>"000100001",
  23370=>"001111001",
  23371=>"110000010",
  23372=>"111111101",
  23373=>"110010110",
  23374=>"110111100",
  23375=>"101011110",
  23376=>"101110101",
  23377=>"010110000",
  23378=>"010010110",
  23379=>"100010101",
  23380=>"000100001",
  23381=>"001001110",
  23382=>"011110110",
  23383=>"101101000",
  23384=>"000011000",
  23385=>"111111101",
  23386=>"111010110",
  23387=>"100111110",
  23388=>"110111101",
  23389=>"000011101",
  23390=>"110101001",
  23391=>"100111010",
  23392=>"001101111",
  23393=>"111000100",
  23394=>"100000010",
  23395=>"101000101",
  23396=>"111010101",
  23397=>"011110101",
  23398=>"100000101",
  23399=>"011101100",
  23400=>"101010001",
  23401=>"111010010",
  23402=>"000110101",
  23403=>"100100001",
  23404=>"111111110",
  23405=>"000101000",
  23406=>"101111111",
  23407=>"110110111",
  23408=>"000100000",
  23409=>"101001110",
  23410=>"100110000",
  23411=>"010101101",
  23412=>"101010111",
  23413=>"010011111",
  23414=>"101011101",
  23415=>"111101100",
  23416=>"001100010",
  23417=>"101111101",
  23418=>"000011100",
  23419=>"101101000",
  23420=>"100110000",
  23421=>"001101000",
  23422=>"000100011",
  23423=>"101011011",
  23424=>"000100000",
  23425=>"000111101",
  23426=>"000100000",
  23427=>"110010110",
  23428=>"111110111",
  23429=>"110010100",
  23430=>"000110101",
  23431=>"110000111",
  23432=>"111110101",
  23433=>"100000100",
  23434=>"100100000",
  23435=>"011011100",
  23436=>"101001100",
  23437=>"000101010",
  23438=>"000001010",
  23439=>"000101110",
  23440=>"000110100",
  23441=>"110110001",
  23442=>"010001110",
  23443=>"001011100",
  23444=>"011111000",
  23445=>"111111001",
  23446=>"011000001",
  23447=>"100100101",
  23448=>"010101101",
  23449=>"100001011",
  23450=>"010100100",
  23451=>"101100101",
  23452=>"001010001",
  23453=>"110111001",
  23454=>"001010101",
  23455=>"010000111",
  23456=>"100000000",
  23457=>"001111111",
  23458=>"110110100",
  23459=>"111110111",
  23460=>"001000000",
  23461=>"111111101",
  23462=>"111110101",
  23463=>"101100011",
  23464=>"111010101",
  23465=>"011101010",
  23466=>"101101010",
  23467=>"110010111",
  23468=>"010010011",
  23469=>"000111101",
  23470=>"111110110",
  23471=>"111110110",
  23472=>"011111011",
  23473=>"101110000",
  23474=>"100101101",
  23475=>"001001010",
  23476=>"001111000",
  23477=>"111110110",
  23478=>"101101011",
  23479=>"011011000",
  23480=>"110001011",
  23481=>"011100000",
  23482=>"001001010",
  23483=>"001010100",
  23484=>"101011000",
  23485=>"010101110",
  23486=>"000010110",
  23487=>"101010000",
  23488=>"101001000",
  23489=>"011110101",
  23490=>"011111011",
  23491=>"001010010",
  23492=>"001110101",
  23493=>"001111000",
  23494=>"001001011",
  23495=>"011100001",
  23496=>"010110111",
  23497=>"101000111",
  23498=>"111111111",
  23499=>"111001010",
  23500=>"110000000",
  23501=>"111100111",
  23502=>"000110100",
  23503=>"001111101",
  23504=>"110001001",
  23505=>"111000110",
  23506=>"010011111",
  23507=>"001101111",
  23508=>"101100001",
  23509=>"100110001",
  23510=>"100111011",
  23511=>"100011001",
  23512=>"000100001",
  23513=>"000000101",
  23514=>"000000000",
  23515=>"010111010",
  23516=>"100011000",
  23517=>"001011100",
  23518=>"111000100",
  23519=>"001010100",
  23520=>"111011001",
  23521=>"011011111",
  23522=>"100111100",
  23523=>"000000111",
  23524=>"010100001",
  23525=>"011010010",
  23526=>"111111100",
  23527=>"111101111",
  23528=>"100010011",
  23529=>"001010011",
  23530=>"101011001",
  23531=>"111101110",
  23532=>"110100011",
  23533=>"011001011",
  23534=>"111111001",
  23535=>"010110100",
  23536=>"011110111",
  23537=>"000111010",
  23538=>"000110011",
  23539=>"000110010",
  23540=>"100000100",
  23541=>"011111010",
  23542=>"010011000",
  23543=>"011100100",
  23544=>"111110001",
  23545=>"100101001",
  23546=>"010101111",
  23547=>"110100110",
  23548=>"111110101",
  23549=>"000101100",
  23550=>"011000100",
  23551=>"010001011",
  23552=>"100000101",
  23553=>"001011001",
  23554=>"010111000",
  23555=>"100010001",
  23556=>"110010101",
  23557=>"110101000",
  23558=>"000010000",
  23559=>"101000000",
  23560=>"101100101",
  23561=>"110111000",
  23562=>"011110100",
  23563=>"010110011",
  23564=>"110000101",
  23565=>"110010001",
  23566=>"010100010",
  23567=>"101110100",
  23568=>"100111100",
  23569=>"100100001",
  23570=>"001011101",
  23571=>"101111011",
  23572=>"011111100",
  23573=>"101001111",
  23574=>"110010100",
  23575=>"110111000",
  23576=>"000111000",
  23577=>"010100000",
  23578=>"100111101",
  23579=>"010010100",
  23580=>"110001000",
  23581=>"110010000",
  23582=>"010010001",
  23583=>"100111000",
  23584=>"000001101",
  23585=>"100100000",
  23586=>"100011111",
  23587=>"111001010",
  23588=>"011111010",
  23589=>"101111011",
  23590=>"110100000",
  23591=>"001001010",
  23592=>"100010011",
  23593=>"001110000",
  23594=>"110111100",
  23595=>"110111100",
  23596=>"010110000",
  23597=>"111001110",
  23598=>"111000000",
  23599=>"101000101",
  23600=>"000011011",
  23601=>"001100101",
  23602=>"111101111",
  23603=>"011101011",
  23604=>"111110000",
  23605=>"111001100",
  23606=>"011010011",
  23607=>"111110101",
  23608=>"101110000",
  23609=>"010000010",
  23610=>"000010110",
  23611=>"111001111",
  23612=>"001100010",
  23613=>"001011011",
  23614=>"100010101",
  23615=>"111101001",
  23616=>"101011011",
  23617=>"110100011",
  23618=>"111010000",
  23619=>"000011111",
  23620=>"110011001",
  23621=>"110110011",
  23622=>"010111110",
  23623=>"111110111",
  23624=>"100101011",
  23625=>"011000011",
  23626=>"101101010",
  23627=>"001001100",
  23628=>"111110111",
  23629=>"110111001",
  23630=>"111001111",
  23631=>"101100101",
  23632=>"011100111",
  23633=>"111001101",
  23634=>"100100001",
  23635=>"011010111",
  23636=>"000110001",
  23637=>"010100100",
  23638=>"010100000",
  23639=>"001001011",
  23640=>"111111010",
  23641=>"101011101",
  23642=>"110110000",
  23643=>"001011111",
  23644=>"000011000",
  23645=>"111111001",
  23646=>"110010110",
  23647=>"111101101",
  23648=>"001100001",
  23649=>"111110100",
  23650=>"011010100",
  23651=>"101100000",
  23652=>"111110110",
  23653=>"010000110",
  23654=>"100010001",
  23655=>"100000110",
  23656=>"000001110",
  23657=>"011010111",
  23658=>"100110000",
  23659=>"100110000",
  23660=>"000101011",
  23661=>"100100100",
  23662=>"110000011",
  23663=>"010011000",
  23664=>"011001110",
  23665=>"010001101",
  23666=>"111000000",
  23667=>"011000111",
  23668=>"111010001",
  23669=>"010111000",
  23670=>"111011111",
  23671=>"111000000",
  23672=>"110010111",
  23673=>"100011010",
  23674=>"111101011",
  23675=>"010010110",
  23676=>"101101111",
  23677=>"011011111",
  23678=>"010101010",
  23679=>"001001110",
  23680=>"101100011",
  23681=>"111111010",
  23682=>"111101001",
  23683=>"000011000",
  23684=>"110111111",
  23685=>"111101001",
  23686=>"111101011",
  23687=>"000100111",
  23688=>"111000101",
  23689=>"000101110",
  23690=>"001101011",
  23691=>"001011011",
  23692=>"111100110",
  23693=>"110111111",
  23694=>"110110110",
  23695=>"000001010",
  23696=>"111111010",
  23697=>"001010100",
  23698=>"010000101",
  23699=>"111110011",
  23700=>"010110011",
  23701=>"000110000",
  23702=>"101010101",
  23703=>"001100001",
  23704=>"001110010",
  23705=>"011001011",
  23706=>"010101101",
  23707=>"100101101",
  23708=>"000011000",
  23709=>"000100000",
  23710=>"010100011",
  23711=>"011100110",
  23712=>"110010011",
  23713=>"100011100",
  23714=>"010010000",
  23715=>"100111101",
  23716=>"011100011",
  23717=>"100010110",
  23718=>"111001011",
  23719=>"001111110",
  23720=>"011000111",
  23721=>"011010101",
  23722=>"110101110",
  23723=>"111100011",
  23724=>"011010111",
  23725=>"011111101",
  23726=>"010000011",
  23727=>"111110101",
  23728=>"110111101",
  23729=>"010001011",
  23730=>"100110000",
  23731=>"010111000",
  23732=>"001011011",
  23733=>"111101110",
  23734=>"111100110",
  23735=>"101101001",
  23736=>"011110110",
  23737=>"111111011",
  23738=>"111101101",
  23739=>"111011111",
  23740=>"101011010",
  23741=>"101110111",
  23742=>"101111001",
  23743=>"001001001",
  23744=>"100100000",
  23745=>"000101101",
  23746=>"001111110",
  23747=>"010011000",
  23748=>"001001100",
  23749=>"011101110",
  23750=>"110110111",
  23751=>"110010110",
  23752=>"111010100",
  23753=>"010001010",
  23754=>"010011011",
  23755=>"110001100",
  23756=>"111000011",
  23757=>"010100100",
  23758=>"100011110",
  23759=>"010100010",
  23760=>"100001110",
  23761=>"111001110",
  23762=>"000001000",
  23763=>"100100110",
  23764=>"110101010",
  23765=>"101110110",
  23766=>"111000000",
  23767=>"101010011",
  23768=>"011111000",
  23769=>"100110101",
  23770=>"110010000",
  23771=>"111000100",
  23772=>"001000010",
  23773=>"010001010",
  23774=>"101111101",
  23775=>"001110110",
  23776=>"110101100",
  23777=>"110100100",
  23778=>"111110000",
  23779=>"011100100",
  23780=>"110010011",
  23781=>"111010101",
  23782=>"111110111",
  23783=>"111111110",
  23784=>"011011011",
  23785=>"110001111",
  23786=>"001010111",
  23787=>"000100000",
  23788=>"000111001",
  23789=>"011001101",
  23790=>"000001000",
  23791=>"110101101",
  23792=>"011010100",
  23793=>"101111110",
  23794=>"010110100",
  23795=>"010101001",
  23796=>"111001110",
  23797=>"000101111",
  23798=>"100110010",
  23799=>"101000001",
  23800=>"000110001",
  23801=>"011010100",
  23802=>"101001011",
  23803=>"101001111",
  23804=>"001001000",
  23805=>"011010101",
  23806=>"100101010",
  23807=>"101110011",
  23808=>"011010010",
  23809=>"010111000",
  23810=>"010011001",
  23811=>"110011110",
  23812=>"010000001",
  23813=>"000011011",
  23814=>"110111110",
  23815=>"110010100",
  23816=>"010010000",
  23817=>"000110111",
  23818=>"111000111",
  23819=>"110101100",
  23820=>"100001010",
  23821=>"110111110",
  23822=>"001010000",
  23823=>"110010100",
  23824=>"100000001",
  23825=>"100010110",
  23826=>"010111110",
  23827=>"011110010",
  23828=>"011010111",
  23829=>"010000101",
  23830=>"101100100",
  23831=>"000111011",
  23832=>"011110010",
  23833=>"011101000",
  23834=>"110101010",
  23835=>"001100001",
  23836=>"001101001",
  23837=>"010010111",
  23838=>"100100110",
  23839=>"011100101",
  23840=>"001111100",
  23841=>"000000101",
  23842=>"001101101",
  23843=>"101110110",
  23844=>"000111010",
  23845=>"110010011",
  23846=>"001000001",
  23847=>"110110001",
  23848=>"110100010",
  23849=>"011100111",
  23850=>"000010110",
  23851=>"010010100",
  23852=>"000000101",
  23853=>"111101111",
  23854=>"010001111",
  23855=>"010110010",
  23856=>"110110000",
  23857=>"100000011",
  23858=>"101101100",
  23859=>"000010111",
  23860=>"100000111",
  23861=>"000000001",
  23862=>"001000110",
  23863=>"011110011",
  23864=>"111111111",
  23865=>"110010001",
  23866=>"101100001",
  23867=>"000011000",
  23868=>"111110101",
  23869=>"001010100",
  23870=>"110110001",
  23871=>"110011001",
  23872=>"001000001",
  23873=>"000000000",
  23874=>"111100101",
  23875=>"111001100",
  23876=>"111101111",
  23877=>"001100110",
  23878=>"110011011",
  23879=>"000000011",
  23880=>"101110110",
  23881=>"110010111",
  23882=>"010101001",
  23883=>"000101000",
  23884=>"111011010",
  23885=>"100010000",
  23886=>"010011000",
  23887=>"010110111",
  23888=>"101111111",
  23889=>"111111011",
  23890=>"110110011",
  23891=>"000010100",
  23892=>"001001110",
  23893=>"000011001",
  23894=>"001101011",
  23895=>"110110100",
  23896=>"110001100",
  23897=>"100011010",
  23898=>"111110111",
  23899=>"100001010",
  23900=>"011110100",
  23901=>"101101110",
  23902=>"010000001",
  23903=>"011010001",
  23904=>"111111110",
  23905=>"011110010",
  23906=>"001100110",
  23907=>"101010000",
  23908=>"010010001",
  23909=>"011011000",
  23910=>"111010000",
  23911=>"111110011",
  23912=>"011011100",
  23913=>"111001110",
  23914=>"010111011",
  23915=>"110110110",
  23916=>"110011111",
  23917=>"001000110",
  23918=>"101110100",
  23919=>"110111101",
  23920=>"110110010",
  23921=>"110101111",
  23922=>"110011001",
  23923=>"001100000",
  23924=>"111011000",
  23925=>"111011011",
  23926=>"000011001",
  23927=>"111000001",
  23928=>"010011000",
  23929=>"011001110",
  23930=>"111110111",
  23931=>"000100100",
  23932=>"110001100",
  23933=>"101110111",
  23934=>"111111110",
  23935=>"111100111",
  23936=>"100101100",
  23937=>"110101011",
  23938=>"010010000",
  23939=>"000100111",
  23940=>"101110110",
  23941=>"100100011",
  23942=>"010101111",
  23943=>"111001001",
  23944=>"000011111",
  23945=>"111010110",
  23946=>"000011000",
  23947=>"000010101",
  23948=>"010001101",
  23949=>"111101111",
  23950=>"001101101",
  23951=>"111111000",
  23952=>"011000111",
  23953=>"111111111",
  23954=>"100001011",
  23955=>"101111011",
  23956=>"000110011",
  23957=>"010000010",
  23958=>"010100101",
  23959=>"011101001",
  23960=>"010100100",
  23961=>"000001111",
  23962=>"000100000",
  23963=>"111100000",
  23964=>"101100111",
  23965=>"110111110",
  23966=>"100010101",
  23967=>"111111001",
  23968=>"101101111",
  23969=>"000000101",
  23970=>"010110100",
  23971=>"001100111",
  23972=>"111001111",
  23973=>"001100000",
  23974=>"011100111",
  23975=>"000000010",
  23976=>"000100101",
  23977=>"101011111",
  23978=>"000010110",
  23979=>"000100101",
  23980=>"011100111",
  23981=>"001001111",
  23982=>"011111111",
  23983=>"011011110",
  23984=>"101100000",
  23985=>"111110100",
  23986=>"011111110",
  23987=>"000101000",
  23988=>"101100111",
  23989=>"101101101",
  23990=>"000110100",
  23991=>"000001011",
  23992=>"000100001",
  23993=>"101111000",
  23994=>"101001111",
  23995=>"010011000",
  23996=>"011101000",
  23997=>"111100101",
  23998=>"110000111",
  23999=>"101000101",
  24000=>"100101110",
  24001=>"110101010",
  24002=>"001101000",
  24003=>"011010110",
  24004=>"010011101",
  24005=>"100101001",
  24006=>"011101000",
  24007=>"110001111",
  24008=>"101110111",
  24009=>"110001001",
  24010=>"000111111",
  24011=>"100001011",
  24012=>"010110111",
  24013=>"000001110",
  24014=>"111101100",
  24015=>"110011110",
  24016=>"010101000",
  24017=>"011101111",
  24018=>"100101101",
  24019=>"101011110",
  24020=>"000101011",
  24021=>"110001000",
  24022=>"010000111",
  24023=>"101111100",
  24024=>"111000110",
  24025=>"111101110",
  24026=>"100111110",
  24027=>"000100011",
  24028=>"000100100",
  24029=>"110011101",
  24030=>"010001011",
  24031=>"100010110",
  24032=>"110111100",
  24033=>"110101110",
  24034=>"111111111",
  24035=>"011111100",
  24036=>"000001010",
  24037=>"000000010",
  24038=>"000100010",
  24039=>"111010101",
  24040=>"010001011",
  24041=>"110000100",
  24042=>"010100011",
  24043=>"000101000",
  24044=>"101000111",
  24045=>"010111111",
  24046=>"010001111",
  24047=>"001111011",
  24048=>"001101100",
  24049=>"101010000",
  24050=>"110100110",
  24051=>"001010111",
  24052=>"110101001",
  24053=>"111010110",
  24054=>"000001001",
  24055=>"000111010",
  24056=>"111111101",
  24057=>"011110100",
  24058=>"010111110",
  24059=>"101001101",
  24060=>"111011001",
  24061=>"000001111",
  24062=>"010101110",
  24063=>"000000011",
  24064=>"110110111",
  24065=>"111000101",
  24066=>"110101000",
  24067=>"001000001",
  24068=>"101011101",
  24069=>"101100000",
  24070=>"011011111",
  24071=>"110011011",
  24072=>"001001011",
  24073=>"001100100",
  24074=>"101111100",
  24075=>"111000000",
  24076=>"001111111",
  24077=>"101111001",
  24078=>"000100110",
  24079=>"111000100",
  24080=>"011010001",
  24081=>"000100101",
  24082=>"011111101",
  24083=>"100010111",
  24084=>"010000011",
  24085=>"010001101",
  24086=>"010110011",
  24087=>"011001001",
  24088=>"111111111",
  24089=>"111011001",
  24090=>"111011011",
  24091=>"101100010",
  24092=>"001100110",
  24093=>"101011001",
  24094=>"100000010",
  24095=>"000000000",
  24096=>"100100000",
  24097=>"100001001",
  24098=>"101010001",
  24099=>"110000010",
  24100=>"101100100",
  24101=>"101100001",
  24102=>"100001101",
  24103=>"101010100",
  24104=>"011101011",
  24105=>"000001011",
  24106=>"110110111",
  24107=>"111110001",
  24108=>"110111011",
  24109=>"100000110",
  24110=>"101010000",
  24111=>"000001010",
  24112=>"011011001",
  24113=>"110110010",
  24114=>"010101100",
  24115=>"100000101",
  24116=>"011111001",
  24117=>"000110001",
  24118=>"010100100",
  24119=>"011011010",
  24120=>"110111000",
  24121=>"011010000",
  24122=>"011010110",
  24123=>"100010001",
  24124=>"000111011",
  24125=>"100011111",
  24126=>"010100010",
  24127=>"000000011",
  24128=>"011100101",
  24129=>"101010110",
  24130=>"110101111",
  24131=>"011000110",
  24132=>"111111001",
  24133=>"100011010",
  24134=>"000000000",
  24135=>"010010111",
  24136=>"001010010",
  24137=>"000001111",
  24138=>"111101011",
  24139=>"101011010",
  24140=>"010100001",
  24141=>"001111111",
  24142=>"101101011",
  24143=>"110000000",
  24144=>"011110111",
  24145=>"101001001",
  24146=>"100000001",
  24147=>"101010100",
  24148=>"101110000",
  24149=>"001000001",
  24150=>"100010011",
  24151=>"110000001",
  24152=>"001111111",
  24153=>"100110101",
  24154=>"000000011",
  24155=>"100111100",
  24156=>"111110000",
  24157=>"100000100",
  24158=>"000111101",
  24159=>"010101100",
  24160=>"001000011",
  24161=>"001010011",
  24162=>"110100101",
  24163=>"111010000",
  24164=>"101010100",
  24165=>"101110001",
  24166=>"001110110",
  24167=>"100001100",
  24168=>"001000111",
  24169=>"000100000",
  24170=>"010111111",
  24171=>"111100111",
  24172=>"100110000",
  24173=>"111101000",
  24174=>"110000000",
  24175=>"011110100",
  24176=>"001111110",
  24177=>"011000111",
  24178=>"011101010",
  24179=>"100000100",
  24180=>"101010101",
  24181=>"000100100",
  24182=>"011010011",
  24183=>"110101010",
  24184=>"101110000",
  24185=>"111101100",
  24186=>"110011010",
  24187=>"011010001",
  24188=>"010100100",
  24189=>"000001011",
  24190=>"000000001",
  24191=>"000011010",
  24192=>"000000111",
  24193=>"101000111",
  24194=>"110111010",
  24195=>"000011111",
  24196=>"110100111",
  24197=>"110011001",
  24198=>"001001010",
  24199=>"100011110",
  24200=>"001001000",
  24201=>"000101100",
  24202=>"001001101",
  24203=>"100111011",
  24204=>"101101010",
  24205=>"100001111",
  24206=>"101111001",
  24207=>"010010100",
  24208=>"010110111",
  24209=>"010010110",
  24210=>"101001100",
  24211=>"100110101",
  24212=>"011101000",
  24213=>"101011110",
  24214=>"100001000",
  24215=>"000010011",
  24216=>"010111010",
  24217=>"010000110",
  24218=>"010001110",
  24219=>"101011101",
  24220=>"011110101",
  24221=>"000101110",
  24222=>"011000000",
  24223=>"000111011",
  24224=>"001000100",
  24225=>"100000100",
  24226=>"110010011",
  24227=>"010101110",
  24228=>"111001100",
  24229=>"000001000",
  24230=>"110110010",
  24231=>"001000100",
  24232=>"000000000",
  24233=>"101000111",
  24234=>"110100111",
  24235=>"001010011",
  24236=>"110011001",
  24237=>"110110001",
  24238=>"110000000",
  24239=>"010110001",
  24240=>"100111100",
  24241=>"100000110",
  24242=>"111000111",
  24243=>"111111110",
  24244=>"111100100",
  24245=>"101001011",
  24246=>"001001100",
  24247=>"100011111",
  24248=>"100101110",
  24249=>"001010011",
  24250=>"110010110",
  24251=>"001000000",
  24252=>"101100100",
  24253=>"010111110",
  24254=>"000101111",
  24255=>"011111001",
  24256=>"001010111",
  24257=>"000100100",
  24258=>"011000011",
  24259=>"100101111",
  24260=>"000110101",
  24261=>"000111011",
  24262=>"011010101",
  24263=>"100001110",
  24264=>"010101110",
  24265=>"110001001",
  24266=>"001101001",
  24267=>"100101010",
  24268=>"011100110",
  24269=>"011000110",
  24270=>"001111000",
  24271=>"010001011",
  24272=>"111000011",
  24273=>"001111010",
  24274=>"011000001",
  24275=>"100110101",
  24276=>"101101010",
  24277=>"100000010",
  24278=>"111011111",
  24279=>"101101110",
  24280=>"000010000",
  24281=>"001011000",
  24282=>"111111100",
  24283=>"110000010",
  24284=>"000100110",
  24285=>"011110000",
  24286=>"100101100",
  24287=>"101111010",
  24288=>"101111011",
  24289=>"100011111",
  24290=>"000000000",
  24291=>"101001000",
  24292=>"110110110",
  24293=>"100110100",
  24294=>"000001000",
  24295=>"101011010",
  24296=>"100101000",
  24297=>"100100000",
  24298=>"011111111",
  24299=>"111111111",
  24300=>"001010101",
  24301=>"111011010",
  24302=>"001011000",
  24303=>"001011110",
  24304=>"111111110",
  24305=>"000000101",
  24306=>"110100100",
  24307=>"000001010",
  24308=>"000101100",
  24309=>"000010010",
  24310=>"110101101",
  24311=>"100010100",
  24312=>"101110011",
  24313=>"011011101",
  24314=>"011010110",
  24315=>"111101110",
  24316=>"101100111",
  24317=>"001101110",
  24318=>"010011000",
  24319=>"000100110",
  24320=>"011010011",
  24321=>"101001110",
  24322=>"000100111",
  24323=>"100011010",
  24324=>"001100000",
  24325=>"010110100",
  24326=>"110110110",
  24327=>"110000101",
  24328=>"001111101",
  24329=>"111011010",
  24330=>"111101001",
  24331=>"001000000",
  24332=>"011111111",
  24333=>"011101001",
  24334=>"101010000",
  24335=>"000000001",
  24336=>"111110001",
  24337=>"100001010",
  24338=>"010110000",
  24339=>"111000010",
  24340=>"100010101",
  24341=>"010100110",
  24342=>"101010111",
  24343=>"100111011",
  24344=>"001101100",
  24345=>"000000001",
  24346=>"101010111",
  24347=>"000101000",
  24348=>"101010000",
  24349=>"111101111",
  24350=>"101110111",
  24351=>"011110000",
  24352=>"110100010",
  24353=>"101011110",
  24354=>"001000100",
  24355=>"011001100",
  24356=>"111011100",
  24357=>"101110111",
  24358=>"011111101",
  24359=>"111010110",
  24360=>"000000011",
  24361=>"010101001",
  24362=>"001011111",
  24363=>"101100000",
  24364=>"010010100",
  24365=>"000000000",
  24366=>"111111011",
  24367=>"110101000",
  24368=>"010001001",
  24369=>"000100001",
  24370=>"101110011",
  24371=>"011110000",
  24372=>"011110011",
  24373=>"011010110",
  24374=>"001001001",
  24375=>"110011011",
  24376=>"101001000",
  24377=>"000010010",
  24378=>"111001000",
  24379=>"100010001",
  24380=>"100110001",
  24381=>"000011000",
  24382=>"001000010",
  24383=>"000111110",
  24384=>"000011000",
  24385=>"111011100",
  24386=>"010110110",
  24387=>"111100101",
  24388=>"101000100",
  24389=>"111110101",
  24390=>"000010011",
  24391=>"000001001",
  24392=>"110111010",
  24393=>"000001001",
  24394=>"100111101",
  24395=>"100010000",
  24396=>"010111010",
  24397=>"100010001",
  24398=>"001110111",
  24399=>"110100101",
  24400=>"101100111",
  24401=>"101001100",
  24402=>"001001111",
  24403=>"110101100",
  24404=>"101110101",
  24405=>"010101100",
  24406=>"101001111",
  24407=>"100000000",
  24408=>"000010010",
  24409=>"001011101",
  24410=>"100001100",
  24411=>"101101001",
  24412=>"011010111",
  24413=>"000001111",
  24414=>"111110011",
  24415=>"000000100",
  24416=>"101110110",
  24417=>"111100100",
  24418=>"101111100",
  24419=>"001010111",
  24420=>"111010111",
  24421=>"100000100",
  24422=>"010101111",
  24423=>"000001000",
  24424=>"100101100",
  24425=>"010000111",
  24426=>"000100001",
  24427=>"110000000",
  24428=>"011110010",
  24429=>"001001001",
  24430=>"100100001",
  24431=>"100011100",
  24432=>"000111101",
  24433=>"001000000",
  24434=>"011001010",
  24435=>"100001001",
  24436=>"001010011",
  24437=>"000001000",
  24438=>"111001000",
  24439=>"011011110",
  24440=>"001000010",
  24441=>"110011011",
  24442=>"100111010",
  24443=>"000110111",
  24444=>"111111101",
  24445=>"011001011",
  24446=>"100011000",
  24447=>"100110110",
  24448=>"000010100",
  24449=>"100000101",
  24450=>"000101000",
  24451=>"100100011",
  24452=>"010111111",
  24453=>"101000100",
  24454=>"101010111",
  24455=>"101000001",
  24456=>"111001110",
  24457=>"101011100",
  24458=>"100110000",
  24459=>"111100011",
  24460=>"110010110",
  24461=>"110011100",
  24462=>"000010100",
  24463=>"000111110",
  24464=>"000011101",
  24465=>"110001110",
  24466=>"000011110",
  24467=>"111010101",
  24468=>"110000000",
  24469=>"110101101",
  24470=>"011011000",
  24471=>"000000011",
  24472=>"011111110",
  24473=>"101001010",
  24474=>"110111100",
  24475=>"101000010",
  24476=>"101011100",
  24477=>"000010000",
  24478=>"100010111",
  24479=>"001000001",
  24480=>"010001100",
  24481=>"101110111",
  24482=>"001001001",
  24483=>"101101111",
  24484=>"100101111",
  24485=>"110100000",
  24486=>"111010000",
  24487=>"110001001",
  24488=>"011011101",
  24489=>"001111100",
  24490=>"100010011",
  24491=>"100110011",
  24492=>"110110110",
  24493=>"010000101",
  24494=>"010000000",
  24495=>"010101010",
  24496=>"011101010",
  24497=>"111010111",
  24498=>"011010011",
  24499=>"010101110",
  24500=>"001010001",
  24501=>"111001000",
  24502=>"011111101",
  24503=>"110000110",
  24504=>"011101111",
  24505=>"001010010",
  24506=>"110010000",
  24507=>"001111010",
  24508=>"001110100",
  24509=>"001001111",
  24510=>"000001000",
  24511=>"101100111",
  24512=>"010010100",
  24513=>"101111100",
  24514=>"111100111",
  24515=>"011100000",
  24516=>"010101010",
  24517=>"010000001",
  24518=>"001000001",
  24519=>"100011100",
  24520=>"010101000",
  24521=>"110000101",
  24522=>"111100111",
  24523=>"100100100",
  24524=>"101000001",
  24525=>"101101011",
  24526=>"010011110",
  24527=>"111001111",
  24528=>"000111001",
  24529=>"101010100",
  24530=>"011110011",
  24531=>"001101001",
  24532=>"111101110",
  24533=>"110011100",
  24534=>"010110011",
  24535=>"111010010",
  24536=>"101100000",
  24537=>"011111110",
  24538=>"111111001",
  24539=>"001101101",
  24540=>"101001111",
  24541=>"000000000",
  24542=>"111000110",
  24543=>"110001111",
  24544=>"101100011",
  24545=>"011110110",
  24546=>"100011110",
  24547=>"011111010",
  24548=>"111001111",
  24549=>"101000101",
  24550=>"011010111",
  24551=>"001001001",
  24552=>"011010110",
  24553=>"110010011",
  24554=>"011011101",
  24555=>"100010111",
  24556=>"100000011",
  24557=>"111110011",
  24558=>"110100001",
  24559=>"000011100",
  24560=>"111101011",
  24561=>"101000010",
  24562=>"011001101",
  24563=>"110110100",
  24564=>"100000110",
  24565=>"110001100",
  24566=>"000110010",
  24567=>"110111010",
  24568=>"011101100",
  24569=>"100100000",
  24570=>"101110111",
  24571=>"111100011",
  24572=>"001001100",
  24573=>"010001110",
  24574=>"101110000",
  24575=>"110001110",
  24576=>"110011101",
  24577=>"110011011",
  24578=>"101110010",
  24579=>"111100000",
  24580=>"110110010",
  24581=>"010100000",
  24582=>"110011100",
  24583=>"011101000",
  24584=>"100000001",
  24585=>"100001000",
  24586=>"001010001",
  24587=>"101000000",
  24588=>"110011110",
  24589=>"010100011",
  24590=>"110011011",
  24591=>"110111000",
  24592=>"000010000",
  24593=>"111101100",
  24594=>"010001000",
  24595=>"100001001",
  24596=>"001100100",
  24597=>"010101100",
  24598=>"001101010",
  24599=>"000110111",
  24600=>"001010001",
  24601=>"001100001",
  24602=>"100000100",
  24603=>"001010001",
  24604=>"010100111",
  24605=>"100101101",
  24606=>"011001000",
  24607=>"010000000",
  24608=>"010110001",
  24609=>"111000000",
  24610=>"001000001",
  24611=>"001110010",
  24612=>"010110100",
  24613=>"011001011",
  24614=>"101000100",
  24615=>"001010100",
  24616=>"001100111",
  24617=>"111011111",
  24618=>"010100111",
  24619=>"110001000",
  24620=>"111101100",
  24621=>"000010001",
  24622=>"110110011",
  24623=>"101101110",
  24624=>"111001011",
  24625=>"100011101",
  24626=>"000101110",
  24627=>"000011110",
  24628=>"101111101",
  24629=>"110001110",
  24630=>"000101110",
  24631=>"100100110",
  24632=>"010000111",
  24633=>"000010011",
  24634=>"000011110",
  24635=>"000011010",
  24636=>"111010101",
  24637=>"011110001",
  24638=>"011010100",
  24639=>"100010100",
  24640=>"110111111",
  24641=>"101000010",
  24642=>"101001111",
  24643=>"011010110",
  24644=>"001011100",
  24645=>"001110101",
  24646=>"001010011",
  24647=>"000110000",
  24648=>"010001001",
  24649=>"110010100",
  24650=>"101110100",
  24651=>"110110101",
  24652=>"100011001",
  24653=>"111110101",
  24654=>"111011000",
  24655=>"011100110",
  24656=>"110110101",
  24657=>"110011011",
  24658=>"110000111",
  24659=>"110101100",
  24660=>"011101010",
  24661=>"011101011",
  24662=>"001110101",
  24663=>"100111110",
  24664=>"111000111",
  24665=>"000000001",
  24666=>"000011100",
  24667=>"011000010",
  24668=>"111001011",
  24669=>"100110001",
  24670=>"110001000",
  24671=>"110001010",
  24672=>"000110101",
  24673=>"000101011",
  24674=>"110000100",
  24675=>"110010010",
  24676=>"000111110",
  24677=>"010011001",
  24678=>"100110010",
  24679=>"101010100",
  24680=>"101001010",
  24681=>"101111111",
  24682=>"010000100",
  24683=>"000000001",
  24684=>"100011110",
  24685=>"011111011",
  24686=>"010101111",
  24687=>"001011001",
  24688=>"110000101",
  24689=>"101011001",
  24690=>"001111000",
  24691=>"001111010",
  24692=>"010010010",
  24693=>"110110000",
  24694=>"000110010",
  24695=>"000010001",
  24696=>"101010011",
  24697=>"000001011",
  24698=>"101000001",
  24699=>"000000100",
  24700=>"011111000",
  24701=>"111101001",
  24702=>"011000011",
  24703=>"101111101",
  24704=>"100101011",
  24705=>"110101101",
  24706=>"100001001",
  24707=>"010000011",
  24708=>"101110110",
  24709=>"101101010",
  24710=>"110100110",
  24711=>"010000100",
  24712=>"011010100",
  24713=>"011101111",
  24714=>"100011000",
  24715=>"110100011",
  24716=>"000011101",
  24717=>"101000111",
  24718=>"010100110",
  24719=>"101100011",
  24720=>"110100111",
  24721=>"100100110",
  24722=>"110000100",
  24723=>"100001100",
  24724=>"011001010",
  24725=>"000101100",
  24726=>"010111101",
  24727=>"110101101",
  24728=>"000111111",
  24729=>"001001110",
  24730=>"110001001",
  24731=>"011100111",
  24732=>"101101010",
  24733=>"011001000",
  24734=>"011011111",
  24735=>"000010011",
  24736=>"001000000",
  24737=>"011011010",
  24738=>"110010100",
  24739=>"011101110",
  24740=>"000000001",
  24741=>"000100010",
  24742=>"011010001",
  24743=>"100101001",
  24744=>"011000101",
  24745=>"001100011",
  24746=>"110010110",
  24747=>"011100010",
  24748=>"111111110",
  24749=>"111010011",
  24750=>"110110101",
  24751=>"010010010",
  24752=>"101001110",
  24753=>"010110001",
  24754=>"100010110",
  24755=>"110010110",
  24756=>"000111010",
  24757=>"010101010",
  24758=>"110110010",
  24759=>"001001010",
  24760=>"101001100",
  24761=>"010101001",
  24762=>"000011011",
  24763=>"111111111",
  24764=>"000010101",
  24765=>"110010001",
  24766=>"001000100",
  24767=>"111100110",
  24768=>"101010010",
  24769=>"110101000",
  24770=>"101100110",
  24771=>"000010101",
  24772=>"000000111",
  24773=>"100100000",
  24774=>"011000010",
  24775=>"111110111",
  24776=>"010101111",
  24777=>"011101111",
  24778=>"100110001",
  24779=>"010110010",
  24780=>"000101010",
  24781=>"011010101",
  24782=>"101111100",
  24783=>"110010011",
  24784=>"000110011",
  24785=>"011011000",
  24786=>"111011011",
  24787=>"101111100",
  24788=>"010010101",
  24789=>"001111101",
  24790=>"100101001",
  24791=>"010101011",
  24792=>"011111111",
  24793=>"111001111",
  24794=>"101001110",
  24795=>"011010010",
  24796=>"011000011",
  24797=>"100110111",
  24798=>"111100110",
  24799=>"100101100",
  24800=>"101000110",
  24801=>"100010111",
  24802=>"101101010",
  24803=>"111010100",
  24804=>"101010010",
  24805=>"101010010",
  24806=>"111110011",
  24807=>"011110111",
  24808=>"000011000",
  24809=>"110100101",
  24810=>"110000000",
  24811=>"000110010",
  24812=>"100011000",
  24813=>"000010110",
  24814=>"100000101",
  24815=>"101100001",
  24816=>"000010110",
  24817=>"000000100",
  24818=>"010011011",
  24819=>"011100010",
  24820=>"110111001",
  24821=>"001101110",
  24822=>"011111111",
  24823=>"011010010",
  24824=>"000110101",
  24825=>"010101000",
  24826=>"011111010",
  24827=>"100101000",
  24828=>"111000010",
  24829=>"001100101",
  24830=>"111110001",
  24831=>"100000110",
  24832=>"000100000",
  24833=>"010001101",
  24834=>"001100011",
  24835=>"110010001",
  24836=>"011011010",
  24837=>"010111010",
  24838=>"111110110",
  24839=>"111010111",
  24840=>"001110000",
  24841=>"011011000",
  24842=>"111000100",
  24843=>"000111110",
  24844=>"110100100",
  24845=>"010011010",
  24846=>"010001101",
  24847=>"010000101",
  24848=>"000010111",
  24849=>"000110001",
  24850=>"110111001",
  24851=>"000000100",
  24852=>"110100111",
  24853=>"001101111",
  24854=>"100010100",
  24855=>"011001010",
  24856=>"010000010",
  24857=>"110100110",
  24858=>"000000001",
  24859=>"011010111",
  24860=>"010011100",
  24861=>"101100111",
  24862=>"001011100",
  24863=>"000101000",
  24864=>"000000011",
  24865=>"001110110",
  24866=>"000010111",
  24867=>"100001011",
  24868=>"011001000",
  24869=>"011000100",
  24870=>"001111111",
  24871=>"011100001",
  24872=>"101011001",
  24873=>"010100011",
  24874=>"010000100",
  24875=>"000101111",
  24876=>"011101011",
  24877=>"100000100",
  24878=>"111111110",
  24879=>"001110111",
  24880=>"010100000",
  24881=>"101010110",
  24882=>"110110010",
  24883=>"001010000",
  24884=>"011011110",
  24885=>"001001001",
  24886=>"100111000",
  24887=>"001111010",
  24888=>"000001010",
  24889=>"000101011",
  24890=>"000111011",
  24891=>"010110100",
  24892=>"100101001",
  24893=>"111011101",
  24894=>"010001111",
  24895=>"110011111",
  24896=>"110010011",
  24897=>"100000000",
  24898=>"000011000",
  24899=>"000111101",
  24900=>"100101011",
  24901=>"000110110",
  24902=>"101001001",
  24903=>"001100110",
  24904=>"001001001",
  24905=>"111101010",
  24906=>"000111101",
  24907=>"100000000",
  24908=>"100110011",
  24909=>"001101010",
  24910=>"000011101",
  24911=>"001000011",
  24912=>"001011101",
  24913=>"101110110",
  24914=>"010110001",
  24915=>"101010001",
  24916=>"011000001",
  24917=>"111010010",
  24918=>"110001000",
  24919=>"111001001",
  24920=>"010011111",
  24921=>"001010000",
  24922=>"111101010",
  24923=>"000000101",
  24924=>"111111011",
  24925=>"000101110",
  24926=>"010000111",
  24927=>"111101010",
  24928=>"000011011",
  24929=>"000010101",
  24930=>"011010111",
  24931=>"100000000",
  24932=>"011010101",
  24933=>"100101011",
  24934=>"110000011",
  24935=>"100111011",
  24936=>"111100000",
  24937=>"110001000",
  24938=>"110001000",
  24939=>"011101111",
  24940=>"101010000",
  24941=>"001110111",
  24942=>"101001111",
  24943=>"100001101",
  24944=>"011110001",
  24945=>"011000010",
  24946=>"101110100",
  24947=>"101100001",
  24948=>"100100110",
  24949=>"001101011",
  24950=>"111010000",
  24951=>"111111101",
  24952=>"010000101",
  24953=>"110010001",
  24954=>"000011010",
  24955=>"001101010",
  24956=>"011101101",
  24957=>"001100110",
  24958=>"111000001",
  24959=>"010110011",
  24960=>"111010010",
  24961=>"000110100",
  24962=>"001110000",
  24963=>"001001110",
  24964=>"101011011",
  24965=>"111110010",
  24966=>"000111010",
  24967=>"001000001",
  24968=>"000101101",
  24969=>"011011010",
  24970=>"000101000",
  24971=>"001011101",
  24972=>"101010110",
  24973=>"101000010",
  24974=>"001011000",
  24975=>"010001010",
  24976=>"111100101",
  24977=>"100100010",
  24978=>"011001001",
  24979=>"011000011",
  24980=>"101000111",
  24981=>"000100111",
  24982=>"000001111",
  24983=>"001110000",
  24984=>"100101000",
  24985=>"111001010",
  24986=>"100111111",
  24987=>"101010001",
  24988=>"101111011",
  24989=>"111111111",
  24990=>"010100100",
  24991=>"110001100",
  24992=>"010010000",
  24993=>"110111111",
  24994=>"110101001",
  24995=>"100001001",
  24996=>"111010000",
  24997=>"010111000",
  24998=>"110101110",
  24999=>"011001110",
  25000=>"001000100",
  25001=>"000100001",
  25002=>"000000100",
  25003=>"000101010",
  25004=>"111000110",
  25005=>"001101011",
  25006=>"011101000",
  25007=>"100000000",
  25008=>"100101110",
  25009=>"010101010",
  25010=>"111111111",
  25011=>"100100010",
  25012=>"010110101",
  25013=>"010000001",
  25014=>"001110010",
  25015=>"100001010",
  25016=>"101001011",
  25017=>"100100000",
  25018=>"001100000",
  25019=>"010000011",
  25020=>"010001101",
  25021=>"010111111",
  25022=>"010111100",
  25023=>"001010000",
  25024=>"010011001",
  25025=>"010111110",
  25026=>"111101000",
  25027=>"111010100",
  25028=>"011010010",
  25029=>"110001101",
  25030=>"001101101",
  25031=>"111101011",
  25032=>"110111010",
  25033=>"110111101",
  25034=>"010010100",
  25035=>"001011010",
  25036=>"010010000",
  25037=>"101011110",
  25038=>"111111011",
  25039=>"110010011",
  25040=>"000110100",
  25041=>"011110010",
  25042=>"001110011",
  25043=>"101011111",
  25044=>"001011100",
  25045=>"010010010",
  25046=>"000010000",
  25047=>"111010001",
  25048=>"110011011",
  25049=>"110100110",
  25050=>"010111001",
  25051=>"100111101",
  25052=>"100000010",
  25053=>"111101110",
  25054=>"101101101",
  25055=>"101100000",
  25056=>"000000111",
  25057=>"010100001",
  25058=>"010100000",
  25059=>"101100110",
  25060=>"100001010",
  25061=>"100101110",
  25062=>"100010111",
  25063=>"100000011",
  25064=>"000010000",
  25065=>"000001111",
  25066=>"110101010",
  25067=>"110010001",
  25068=>"101000111",
  25069=>"011111100",
  25070=>"111001001",
  25071=>"011000111",
  25072=>"000111001",
  25073=>"100111100",
  25074=>"100011011",
  25075=>"010111010",
  25076=>"110010110",
  25077=>"111101100",
  25078=>"100011001",
  25079=>"001001000",
  25080=>"110001111",
  25081=>"100001000",
  25082=>"111110001",
  25083=>"111001011",
  25084=>"100101101",
  25085=>"000010000",
  25086=>"110111000",
  25087=>"111000101",
  25088=>"110111011",
  25089=>"011100011",
  25090=>"110010001",
  25091=>"101011010",
  25092=>"011101011",
  25093=>"110111000",
  25094=>"001111111",
  25095=>"001111000",
  25096=>"011111101",
  25097=>"101111000",
  25098=>"100001001",
  25099=>"000011001",
  25100=>"000111110",
  25101=>"100001100",
  25102=>"110001000",
  25103=>"001001001",
  25104=>"101011100",
  25105=>"001010100",
  25106=>"011001100",
  25107=>"101100100",
  25108=>"100110000",
  25109=>"101010110",
  25110=>"100001111",
  25111=>"110100000",
  25112=>"110111010",
  25113=>"001000001",
  25114=>"101100101",
  25115=>"011000111",
  25116=>"000001001",
  25117=>"110111101",
  25118=>"001000010",
  25119=>"110010100",
  25120=>"011011001",
  25121=>"101100011",
  25122=>"110101010",
  25123=>"011110011",
  25124=>"001111111",
  25125=>"000110011",
  25126=>"111000111",
  25127=>"000011011",
  25128=>"110010110",
  25129=>"011011011",
  25130=>"011010101",
  25131=>"101000110",
  25132=>"101110111",
  25133=>"101101110",
  25134=>"011000000",
  25135=>"110111110",
  25136=>"010000101",
  25137=>"110001110",
  25138=>"010110101",
  25139=>"000000111",
  25140=>"111100001",
  25141=>"000001110",
  25142=>"101100010",
  25143=>"110000101",
  25144=>"001111110",
  25145=>"000010011",
  25146=>"011110111",
  25147=>"011110111",
  25148=>"000110101",
  25149=>"000000111",
  25150=>"101000000",
  25151=>"010001010",
  25152=>"110010101",
  25153=>"010111101",
  25154=>"001111111",
  25155=>"011101101",
  25156=>"010100000",
  25157=>"110110101",
  25158=>"001000111",
  25159=>"011101101",
  25160=>"001001111",
  25161=>"110110111",
  25162=>"011011001",
  25163=>"101100000",
  25164=>"001100110",
  25165=>"100111000",
  25166=>"100010111",
  25167=>"000101001",
  25168=>"111110100",
  25169=>"001111010",
  25170=>"110100101",
  25171=>"011001100",
  25172=>"001000000",
  25173=>"110000000",
  25174=>"100111100",
  25175=>"010100111",
  25176=>"000010101",
  25177=>"111110011",
  25178=>"000001100",
  25179=>"000000010",
  25180=>"100010011",
  25181=>"010000001",
  25182=>"001101101",
  25183=>"011001011",
  25184=>"010000010",
  25185=>"101111001",
  25186=>"100101010",
  25187=>"101001010",
  25188=>"000000000",
  25189=>"101101100",
  25190=>"111111100",
  25191=>"110001011",
  25192=>"111110001",
  25193=>"010111111",
  25194=>"100010011",
  25195=>"100001000",
  25196=>"111101110",
  25197=>"111001001",
  25198=>"000100110",
  25199=>"110011010",
  25200=>"110011010",
  25201=>"100001100",
  25202=>"111001111",
  25203=>"110011010",
  25204=>"100110000",
  25205=>"000000001",
  25206=>"001111110",
  25207=>"100110110",
  25208=>"100000110",
  25209=>"101101011",
  25210=>"111101101",
  25211=>"100100011",
  25212=>"111011101",
  25213=>"100010001",
  25214=>"110111010",
  25215=>"011010111",
  25216=>"000000110",
  25217=>"000000010",
  25218=>"010000111",
  25219=>"010001000",
  25220=>"010010110",
  25221=>"100100101",
  25222=>"100001101",
  25223=>"110011000",
  25224=>"110011001",
  25225=>"110010111",
  25226=>"111110000",
  25227=>"011100000",
  25228=>"111100111",
  25229=>"100010001",
  25230=>"010101000",
  25231=>"100000011",
  25232=>"010001110",
  25233=>"111000011",
  25234=>"001100001",
  25235=>"000000101",
  25236=>"110101011",
  25237=>"101101011",
  25238=>"110011011",
  25239=>"010100011",
  25240=>"000101010",
  25241=>"001011000",
  25242=>"101011110",
  25243=>"100010111",
  25244=>"000011010",
  25245=>"011101011",
  25246=>"001011000",
  25247=>"011001100",
  25248=>"110001111",
  25249=>"101001000",
  25250=>"101110000",
  25251=>"111001110",
  25252=>"110000110",
  25253=>"010001100",
  25254=>"100000111",
  25255=>"000010000",
  25256=>"101110111",
  25257=>"001100110",
  25258=>"100000001",
  25259=>"110100011",
  25260=>"011000011",
  25261=>"010111101",
  25262=>"000000001",
  25263=>"101011101",
  25264=>"001110010",
  25265=>"100111010",
  25266=>"100101011",
  25267=>"100101100",
  25268=>"000001001",
  25269=>"011011001",
  25270=>"000101101",
  25271=>"010010011",
  25272=>"100101010",
  25273=>"010001110",
  25274=>"011100100",
  25275=>"011010000",
  25276=>"001011101",
  25277=>"111111010",
  25278=>"111101100",
  25279=>"011001000",
  25280=>"001111110",
  25281=>"011100111",
  25282=>"000000010",
  25283=>"111011110",
  25284=>"010101100",
  25285=>"110001110",
  25286=>"111001111",
  25287=>"010101000",
  25288=>"010000100",
  25289=>"010111000",
  25290=>"011101001",
  25291=>"000001100",
  25292=>"100010010",
  25293=>"110000000",
  25294=>"100110100",
  25295=>"111110010",
  25296=>"101100111",
  25297=>"000011101",
  25298=>"101110111",
  25299=>"111011101",
  25300=>"001000000",
  25301=>"000101000",
  25302=>"111111011",
  25303=>"111110110",
  25304=>"101001101",
  25305=>"000010001",
  25306=>"100000001",
  25307=>"100101001",
  25308=>"011111100",
  25309=>"001100011",
  25310=>"010000100",
  25311=>"011010011",
  25312=>"000000001",
  25313=>"011110011",
  25314=>"011110110",
  25315=>"011010001",
  25316=>"100011011",
  25317=>"011000111",
  25318=>"000011001",
  25319=>"010001000",
  25320=>"000111010",
  25321=>"111010001",
  25322=>"010111011",
  25323=>"100001010",
  25324=>"000011011",
  25325=>"000010110",
  25326=>"111110010",
  25327=>"100010100",
  25328=>"111011000",
  25329=>"001110110",
  25330=>"110011000",
  25331=>"110011101",
  25332=>"001010011",
  25333=>"110100111",
  25334=>"010101100",
  25335=>"011111101",
  25336=>"001110001",
  25337=>"000101111",
  25338=>"000110001",
  25339=>"111011100",
  25340=>"011110111",
  25341=>"010001110",
  25342=>"101110010",
  25343=>"011110110",
  25344=>"101010100",
  25345=>"010000011",
  25346=>"101001110",
  25347=>"101100011",
  25348=>"101100011",
  25349=>"001000001",
  25350=>"010101100",
  25351=>"101110011",
  25352=>"111101000",
  25353=>"110000110",
  25354=>"011011000",
  25355=>"100001111",
  25356=>"110101011",
  25357=>"001101010",
  25358=>"100011011",
  25359=>"011000000",
  25360=>"011001010",
  25361=>"001100101",
  25362=>"111100001",
  25363=>"110110011",
  25364=>"011001001",
  25365=>"000010100",
  25366=>"010001000",
  25367=>"110011000",
  25368=>"111101100",
  25369=>"010000100",
  25370=>"001100100",
  25371=>"111101001",
  25372=>"011001001",
  25373=>"001110000",
  25374=>"101111000",
  25375=>"101000010",
  25376=>"111010011",
  25377=>"010100100",
  25378=>"011110100",
  25379=>"101010010",
  25380=>"011000001",
  25381=>"110101111",
  25382=>"101111100",
  25383=>"100010101",
  25384=>"011101101",
  25385=>"001001101",
  25386=>"011110010",
  25387=>"000111100",
  25388=>"000010100",
  25389=>"000000001",
  25390=>"111100101",
  25391=>"011000101",
  25392=>"110000110",
  25393=>"110101110",
  25394=>"100010000",
  25395=>"001001100",
  25396=>"011010001",
  25397=>"010011110",
  25398=>"101011101",
  25399=>"010001101",
  25400=>"000010111",
  25401=>"101110111",
  25402=>"001001011",
  25403=>"001100101",
  25404=>"101101101",
  25405=>"000000000",
  25406=>"110101011",
  25407=>"100010001",
  25408=>"110100011",
  25409=>"001110101",
  25410=>"100111100",
  25411=>"001001011",
  25412=>"010011111",
  25413=>"000000010",
  25414=>"011100000",
  25415=>"000110000",
  25416=>"011110000",
  25417=>"110101111",
  25418=>"100001000",
  25419=>"111100100",
  25420=>"101110111",
  25421=>"101011010",
  25422=>"001101001",
  25423=>"001110011",
  25424=>"111001111",
  25425=>"101110111",
  25426=>"110110110",
  25427=>"111100000",
  25428=>"111000001",
  25429=>"000111010",
  25430=>"000001010",
  25431=>"001011001",
  25432=>"000111111",
  25433=>"000101111",
  25434=>"101100010",
  25435=>"110111110",
  25436=>"110000011",
  25437=>"011101100",
  25438=>"101000000",
  25439=>"000101111",
  25440=>"101100001",
  25441=>"111110101",
  25442=>"110010000",
  25443=>"101100110",
  25444=>"001101100",
  25445=>"110000111",
  25446=>"001101010",
  25447=>"010110000",
  25448=>"111010110",
  25449=>"101111110",
  25450=>"101101100",
  25451=>"110100010",
  25452=>"001000011",
  25453=>"001001000",
  25454=>"010111000",
  25455=>"101110110",
  25456=>"101001010",
  25457=>"010001101",
  25458=>"111100111",
  25459=>"111011000",
  25460=>"101111110",
  25461=>"000000000",
  25462=>"000111101",
  25463=>"001101011",
  25464=>"111010010",
  25465=>"101001001",
  25466=>"011110100",
  25467=>"100101011",
  25468=>"000111011",
  25469=>"100101001",
  25470=>"011000101",
  25471=>"111000111",
  25472=>"001110000",
  25473=>"100110111",
  25474=>"110001011",
  25475=>"001011111",
  25476=>"100000111",
  25477=>"100010110",
  25478=>"010000001",
  25479=>"101101000",
  25480=>"000010110",
  25481=>"101011001",
  25482=>"100110110",
  25483=>"101101111",
  25484=>"000000000",
  25485=>"110101011",
  25486=>"000011011",
  25487=>"001011010",
  25488=>"101100010",
  25489=>"001101110",
  25490=>"011110000",
  25491=>"000000100",
  25492=>"100000011",
  25493=>"110110110",
  25494=>"000011011",
  25495=>"011010101",
  25496=>"000100000",
  25497=>"111001110",
  25498=>"000101111",
  25499=>"001000101",
  25500=>"001100111",
  25501=>"010111110",
  25502=>"110101010",
  25503=>"101001110",
  25504=>"011001001",
  25505=>"010110001",
  25506=>"111001110",
  25507=>"000010110",
  25508=>"101110111",
  25509=>"110111011",
  25510=>"111101000",
  25511=>"000110110",
  25512=>"011110100",
  25513=>"000100101",
  25514=>"100000110",
  25515=>"001011100",
  25516=>"000101111",
  25517=>"011001010",
  25518=>"101010011",
  25519=>"110101011",
  25520=>"100010010",
  25521=>"000101010",
  25522=>"110111101",
  25523=>"100101011",
  25524=>"011110011",
  25525=>"011011100",
  25526=>"000011010",
  25527=>"110111011",
  25528=>"011111100",
  25529=>"000000110",
  25530=>"111011111",
  25531=>"010100110",
  25532=>"110010101",
  25533=>"011011010",
  25534=>"010111111",
  25535=>"111100001",
  25536=>"111101111",
  25537=>"101000011",
  25538=>"001000101",
  25539=>"111111111",
  25540=>"000101101",
  25541=>"010011110",
  25542=>"010110101",
  25543=>"111110010",
  25544=>"111001100",
  25545=>"100110001",
  25546=>"001010100",
  25547=>"100001111",
  25548=>"000101111",
  25549=>"111101101",
  25550=>"011110110",
  25551=>"011100000",
  25552=>"100011001",
  25553=>"110010001",
  25554=>"001011011",
  25555=>"011110111",
  25556=>"000011000",
  25557=>"101000111",
  25558=>"010001000",
  25559=>"010101110",
  25560=>"100010001",
  25561=>"001001011",
  25562=>"110100110",
  25563=>"010010110",
  25564=>"000010111",
  25565=>"000100000",
  25566=>"010000011",
  25567=>"111011111",
  25568=>"110000101",
  25569=>"101000011",
  25570=>"101000000",
  25571=>"110010000",
  25572=>"000001111",
  25573=>"001011100",
  25574=>"000101111",
  25575=>"111000100",
  25576=>"001001101",
  25577=>"001111100",
  25578=>"111010001",
  25579=>"110100001",
  25580=>"011000111",
  25581=>"101101001",
  25582=>"001001011",
  25583=>"101011100",
  25584=>"001100100",
  25585=>"111001110",
  25586=>"001011010",
  25587=>"101110110",
  25588=>"111010111",
  25589=>"111101100",
  25590=>"101101111",
  25591=>"100001111",
  25592=>"010010110",
  25593=>"000111010",
  25594=>"110001010",
  25595=>"110010101",
  25596=>"111001010",
  25597=>"100010100",
  25598=>"111101111",
  25599=>"111000100",
  25600=>"110010000",
  25601=>"001110101",
  25602=>"010000111",
  25603=>"010100000",
  25604=>"010100010",
  25605=>"001110011",
  25606=>"111001101",
  25607=>"100111001",
  25608=>"111010110",
  25609=>"001011001",
  25610=>"101111111",
  25611=>"101010010",
  25612=>"010011000",
  25613=>"101101010",
  25614=>"011101110",
  25615=>"010001001",
  25616=>"110010101",
  25617=>"010100011",
  25618=>"101001111",
  25619=>"100011011",
  25620=>"111101001",
  25621=>"100001010",
  25622=>"100110100",
  25623=>"100101011",
  25624=>"111100111",
  25625=>"111101000",
  25626=>"111110100",
  25627=>"110101110",
  25628=>"011101000",
  25629=>"000110110",
  25630=>"100100011",
  25631=>"011010011",
  25632=>"100000000",
  25633=>"001010110",
  25634=>"110111001",
  25635=>"111011010",
  25636=>"110001011",
  25637=>"001101111",
  25638=>"111000011",
  25639=>"011010010",
  25640=>"010100011",
  25641=>"110100111",
  25642=>"010110001",
  25643=>"011111011",
  25644=>"000001100",
  25645=>"011111110",
  25646=>"000111111",
  25647=>"011101111",
  25648=>"110111001",
  25649=>"011101010",
  25650=>"101110111",
  25651=>"000110101",
  25652=>"101111011",
  25653=>"001000001",
  25654=>"101010001",
  25655=>"001010111",
  25656=>"001101110",
  25657=>"110101000",
  25658=>"111111111",
  25659=>"111011111",
  25660=>"000101001",
  25661=>"010100000",
  25662=>"010001101",
  25663=>"001110011",
  25664=>"111100111",
  25665=>"001010111",
  25666=>"110110011",
  25667=>"110110101",
  25668=>"110011000",
  25669=>"111010000",
  25670=>"011100010",
  25671=>"010101000",
  25672=>"101111110",
  25673=>"101100101",
  25674=>"000000010",
  25675=>"000111011",
  25676=>"100110011",
  25677=>"100001111",
  25678=>"101101001",
  25679=>"110000110",
  25680=>"000011000",
  25681=>"010010100",
  25682=>"101110100",
  25683=>"110000010",
  25684=>"100001010",
  25685=>"011101011",
  25686=>"111001010",
  25687=>"011111010",
  25688=>"011110001",
  25689=>"111100001",
  25690=>"000001001",
  25691=>"100011100",
  25692=>"001100000",
  25693=>"101010001",
  25694=>"001100100",
  25695=>"000000101",
  25696=>"011101000",
  25697=>"111010111",
  25698=>"001110010",
  25699=>"010001110",
  25700=>"101011110",
  25701=>"011000111",
  25702=>"011001001",
  25703=>"101101101",
  25704=>"000000000",
  25705=>"001001010",
  25706=>"000101011",
  25707=>"110010100",
  25708=>"111100111",
  25709=>"000001111",
  25710=>"011000100",
  25711=>"111000100",
  25712=>"000110010",
  25713=>"000111101",
  25714=>"010001000",
  25715=>"000101110",
  25716=>"001101101",
  25717=>"101100110",
  25718=>"110000111",
  25719=>"011101010",
  25720=>"011101111",
  25721=>"111011111",
  25722=>"111011001",
  25723=>"110001100",
  25724=>"010111101",
  25725=>"001110100",
  25726=>"001000101",
  25727=>"110100101",
  25728=>"110010010",
  25729=>"000010110",
  25730=>"101011001",
  25731=>"001101111",
  25732=>"000010000",
  25733=>"101010100",
  25734=>"011001110",
  25735=>"001100010",
  25736=>"100111110",
  25737=>"110101100",
  25738=>"001110001",
  25739=>"010100101",
  25740=>"111110110",
  25741=>"111101110",
  25742=>"111001011",
  25743=>"010001111",
  25744=>"111101010",
  25745=>"100010010",
  25746=>"100101111",
  25747=>"111010011",
  25748=>"100001011",
  25749=>"000101011",
  25750=>"111100101",
  25751=>"100001100",
  25752=>"011101101",
  25753=>"001011111",
  25754=>"100001101",
  25755=>"000000101",
  25756=>"111111111",
  25757=>"000000010",
  25758=>"101101000",
  25759=>"101000100",
  25760=>"110001100",
  25761=>"111010100",
  25762=>"111111010",
  25763=>"110000101",
  25764=>"001100100",
  25765=>"111111100",
  25766=>"101100101",
  25767=>"010110000",
  25768=>"100110111",
  25769=>"001010000",
  25770=>"110111101",
  25771=>"111100100",
  25772=>"111000011",
  25773=>"110101010",
  25774=>"000101010",
  25775=>"000000011",
  25776=>"011011110",
  25777=>"010001011",
  25778=>"011000110",
  25779=>"111011010",
  25780=>"100001101",
  25781=>"001001001",
  25782=>"010010011",
  25783=>"110011000",
  25784=>"011001011",
  25785=>"110010101",
  25786=>"111100010",
  25787=>"101111010",
  25788=>"111100010",
  25789=>"011011100",
  25790=>"000110111",
  25791=>"001001010",
  25792=>"111100101",
  25793=>"011000010",
  25794=>"001011001",
  25795=>"011011101",
  25796=>"010011010",
  25797=>"001011001",
  25798=>"011110111",
  25799=>"010001001",
  25800=>"000001010",
  25801=>"011110011",
  25802=>"101111101",
  25803=>"101001110",
  25804=>"011001110",
  25805=>"000101100",
  25806=>"000111001",
  25807=>"010011001",
  25808=>"111100110",
  25809=>"111111001",
  25810=>"001110000",
  25811=>"100110000",
  25812=>"111010011",
  25813=>"100101001",
  25814=>"001001110",
  25815=>"001110000",
  25816=>"000000011",
  25817=>"000100111",
  25818=>"001010010",
  25819=>"010001001",
  25820=>"111101100",
  25821=>"010001111",
  25822=>"000000010",
  25823=>"011111101",
  25824=>"101101010",
  25825=>"111011111",
  25826=>"001100001",
  25827=>"011000100",
  25828=>"110001110",
  25829=>"011010001",
  25830=>"101011010",
  25831=>"111101110",
  25832=>"001111010",
  25833=>"100011010",
  25834=>"100101000",
  25835=>"011000011",
  25836=>"001101100",
  25837=>"010100101",
  25838=>"100100110",
  25839=>"110111101",
  25840=>"110101011",
  25841=>"111110100",
  25842=>"101011011",
  25843=>"111110111",
  25844=>"001010001",
  25845=>"110110110",
  25846=>"101100010",
  25847=>"000010110",
  25848=>"111100111",
  25849=>"001011000",
  25850=>"000110110",
  25851=>"000000110",
  25852=>"000001110",
  25853=>"111101111",
  25854=>"111111000",
  25855=>"101100001",
  25856=>"011010100",
  25857=>"000101001",
  25858=>"001011010",
  25859=>"100101011",
  25860=>"000101011",
  25861=>"100011001",
  25862=>"100011001",
  25863=>"001110010",
  25864=>"010011100",
  25865=>"110001100",
  25866=>"010001100",
  25867=>"001011100",
  25868=>"011111111",
  25869=>"011111001",
  25870=>"110110100",
  25871=>"110000011",
  25872=>"111011010",
  25873=>"110100000",
  25874=>"011110110",
  25875=>"011110110",
  25876=>"101000100",
  25877=>"101001100",
  25878=>"110010001",
  25879=>"101101100",
  25880=>"100100001",
  25881=>"011011011",
  25882=>"110101011",
  25883=>"000000010",
  25884=>"100000110",
  25885=>"110000110",
  25886=>"010100001",
  25887=>"011000011",
  25888=>"100101000",
  25889=>"001001101",
  25890=>"000010001",
  25891=>"010101000",
  25892=>"001001010",
  25893=>"100110011",
  25894=>"010111011",
  25895=>"110000101",
  25896=>"100100111",
  25897=>"001000000",
  25898=>"001001001",
  25899=>"100010000",
  25900=>"100010111",
  25901=>"001000010",
  25902=>"011101000",
  25903=>"001110101",
  25904=>"001100111",
  25905=>"110011100",
  25906=>"000111111",
  25907=>"101111010",
  25908=>"100101001",
  25909=>"100011011",
  25910=>"000101011",
  25911=>"110000100",
  25912=>"101001001",
  25913=>"110010000",
  25914=>"010101100",
  25915=>"000101000",
  25916=>"011110110",
  25917=>"010110111",
  25918=>"110110011",
  25919=>"011000011",
  25920=>"101100010",
  25921=>"111000110",
  25922=>"001101000",
  25923=>"101110101",
  25924=>"010001110",
  25925=>"000110001",
  25926=>"011010011",
  25927=>"000100011",
  25928=>"001010001",
  25929=>"111101010",
  25930=>"111010110",
  25931=>"101010111",
  25932=>"100011000",
  25933=>"111100110",
  25934=>"101000100",
  25935=>"000000110",
  25936=>"011110001",
  25937=>"101111110",
  25938=>"011011101",
  25939=>"100000111",
  25940=>"000010110",
  25941=>"101100011",
  25942=>"101100001",
  25943=>"101011110",
  25944=>"010000001",
  25945=>"101001000",
  25946=>"100011100",
  25947=>"000111100",
  25948=>"101100111",
  25949=>"111100100",
  25950=>"111101111",
  25951=>"000101011",
  25952=>"111000110",
  25953=>"011000111",
  25954=>"100010110",
  25955=>"010011111",
  25956=>"101010111",
  25957=>"010001111",
  25958=>"100010011",
  25959=>"111011100",
  25960=>"000100011",
  25961=>"000001101",
  25962=>"011100011",
  25963=>"000101011",
  25964=>"100101000",
  25965=>"011110011",
  25966=>"111110011",
  25967=>"110110101",
  25968=>"101001001",
  25969=>"101001111",
  25970=>"010111101",
  25971=>"101000010",
  25972=>"110101011",
  25973=>"011111100",
  25974=>"111011000",
  25975=>"001100101",
  25976=>"000011001",
  25977=>"101011101",
  25978=>"100111010",
  25979=>"010101000",
  25980=>"100001011",
  25981=>"101000111",
  25982=>"111100000",
  25983=>"110101111",
  25984=>"011111101",
  25985=>"001110011",
  25986=>"110001100",
  25987=>"011011111",
  25988=>"111111011",
  25989=>"100101000",
  25990=>"101110110",
  25991=>"110001111",
  25992=>"110010010",
  25993=>"111101000",
  25994=>"111010111",
  25995=>"010100110",
  25996=>"001010000",
  25997=>"111001000",
  25998=>"111011011",
  25999=>"000110010",
  26000=>"010111000",
  26001=>"001011101",
  26002=>"000011110",
  26003=>"010010010",
  26004=>"000101011",
  26005=>"101000000",
  26006=>"111010011",
  26007=>"001011001",
  26008=>"000101011",
  26009=>"100111011",
  26010=>"011000001",
  26011=>"100111000",
  26012=>"110110101",
  26013=>"101101001",
  26014=>"110101110",
  26015=>"111101100",
  26016=>"100110100",
  26017=>"011010001",
  26018=>"101010110",
  26019=>"110110000",
  26020=>"111101100",
  26021=>"000101000",
  26022=>"110101011",
  26023=>"101111011",
  26024=>"000100101",
  26025=>"010011101",
  26026=>"011100010",
  26027=>"011010010",
  26028=>"111011000",
  26029=>"011010111",
  26030=>"001000000",
  26031=>"011110010",
  26032=>"000001101",
  26033=>"100100011",
  26034=>"010000111",
  26035=>"000000001",
  26036=>"011110011",
  26037=>"101011101",
  26038=>"101011100",
  26039=>"011100110",
  26040=>"001111000",
  26041=>"010101001",
  26042=>"010010010",
  26043=>"110110000",
  26044=>"010100011",
  26045=>"001011001",
  26046=>"000011000",
  26047=>"111101011",
  26048=>"001000111",
  26049=>"111000010",
  26050=>"001110010",
  26051=>"110001000",
  26052=>"001111100",
  26053=>"111110000",
  26054=>"111011001",
  26055=>"000001000",
  26056=>"010011011",
  26057=>"100111111",
  26058=>"000001010",
  26059=>"111000110",
  26060=>"001011001",
  26061=>"010111000",
  26062=>"011001110",
  26063=>"001011000",
  26064=>"100110001",
  26065=>"110111100",
  26066=>"100100000",
  26067=>"010111100",
  26068=>"100110111",
  26069=>"110000000",
  26070=>"111110000",
  26071=>"100011111",
  26072=>"110110110",
  26073=>"100011111",
  26074=>"111111111",
  26075=>"001101010",
  26076=>"011101011",
  26077=>"110110111",
  26078=>"001000001",
  26079=>"000100101",
  26080=>"000111011",
  26081=>"000000011",
  26082=>"111011100",
  26083=>"111011011",
  26084=>"010110101",
  26085=>"100110011",
  26086=>"001100000",
  26087=>"110011001",
  26088=>"100001110",
  26089=>"110101111",
  26090=>"000111100",
  26091=>"110100001",
  26092=>"111010111",
  26093=>"000100110",
  26094=>"101010000",
  26095=>"111011100",
  26096=>"010110111",
  26097=>"110101001",
  26098=>"101111111",
  26099=>"001100111",
  26100=>"110000111",
  26101=>"000010000",
  26102=>"111101011",
  26103=>"010100010",
  26104=>"000010011",
  26105=>"010110000",
  26106=>"100110111",
  26107=>"110001001",
  26108=>"000000110",
  26109=>"011111101",
  26110=>"110010110",
  26111=>"101100000",
  26112=>"101111010",
  26113=>"000100011",
  26114=>"101111010",
  26115=>"001010000",
  26116=>"111111111",
  26117=>"000111101",
  26118=>"101101101",
  26119=>"101001111",
  26120=>"011011010",
  26121=>"011100111",
  26122=>"011100110",
  26123=>"000110101",
  26124=>"101100100",
  26125=>"110111111",
  26126=>"000001011",
  26127=>"101010111",
  26128=>"001001101",
  26129=>"000000100",
  26130=>"111000001",
  26131=>"010111001",
  26132=>"110000000",
  26133=>"100000101",
  26134=>"100111100",
  26135=>"111110111",
  26136=>"111101001",
  26137=>"001100011",
  26138=>"100011101",
  26139=>"010101010",
  26140=>"110001001",
  26141=>"000001001",
  26142=>"001101101",
  26143=>"100100001",
  26144=>"101110010",
  26145=>"101111100",
  26146=>"001110000",
  26147=>"011010101",
  26148=>"001000101",
  26149=>"111111111",
  26150=>"110001101",
  26151=>"100101100",
  26152=>"100101000",
  26153=>"011111011",
  26154=>"000100101",
  26155=>"010011100",
  26156=>"011111110",
  26157=>"111110111",
  26158=>"001111000",
  26159=>"110001011",
  26160=>"110010011",
  26161=>"101101011",
  26162=>"110110010",
  26163=>"000100000",
  26164=>"010000110",
  26165=>"110111011",
  26166=>"011101100",
  26167=>"001010001",
  26168=>"001000000",
  26169=>"001101111",
  26170=>"011100100",
  26171=>"010011101",
  26172=>"001011100",
  26173=>"000011001",
  26174=>"100101000",
  26175=>"100101101",
  26176=>"101111001",
  26177=>"100110011",
  26178=>"100010111",
  26179=>"111000101",
  26180=>"101000000",
  26181=>"101000111",
  26182=>"111100000",
  26183=>"101001010",
  26184=>"000111000",
  26185=>"111010001",
  26186=>"110011111",
  26187=>"100110001",
  26188=>"000011000",
  26189=>"111101101",
  26190=>"010111110",
  26191=>"111101101",
  26192=>"111100011",
  26193=>"000100010",
  26194=>"101001011",
  26195=>"000110010",
  26196=>"110010111",
  26197=>"010001011",
  26198=>"011110101",
  26199=>"010110110",
  26200=>"011010101",
  26201=>"111110010",
  26202=>"001011110",
  26203=>"100111111",
  26204=>"010111000",
  26205=>"101110011",
  26206=>"000000110",
  26207=>"110011011",
  26208=>"100011110",
  26209=>"000000010",
  26210=>"100111111",
  26211=>"110010011",
  26212=>"111111010",
  26213=>"011100011",
  26214=>"011101011",
  26215=>"011010110",
  26216=>"110100101",
  26217=>"001010010",
  26218=>"001101100",
  26219=>"000011011",
  26220=>"001100110",
  26221=>"000000010",
  26222=>"111011001",
  26223=>"010111111",
  26224=>"111001100",
  26225=>"101001011",
  26226=>"001101111",
  26227=>"111011011",
  26228=>"100000101",
  26229=>"010010001",
  26230=>"101010100",
  26231=>"100100100",
  26232=>"000111000",
  26233=>"001111001",
  26234=>"010110101",
  26235=>"010101100",
  26236=>"111111001",
  26237=>"001011001",
  26238=>"111101111",
  26239=>"011100101",
  26240=>"001010011",
  26241=>"011111100",
  26242=>"011001001",
  26243=>"011000000",
  26244=>"011011010",
  26245=>"000000001",
  26246=>"100110100",
  26247=>"001010110",
  26248=>"100101000",
  26249=>"101000110",
  26250=>"010010010",
  26251=>"110000000",
  26252=>"010101011",
  26253=>"011010101",
  26254=>"010001000",
  26255=>"010101010",
  26256=>"110111001",
  26257=>"110001101",
  26258=>"110101010",
  26259=>"011010000",
  26260=>"000111011",
  26261=>"111101001",
  26262=>"011000111",
  26263=>"001001101",
  26264=>"001100100",
  26265=>"001000110",
  26266=>"100000010",
  26267=>"001110000",
  26268=>"100011010",
  26269=>"000000010",
  26270=>"011010111",
  26271=>"100010100",
  26272=>"101100010",
  26273=>"111101000",
  26274=>"110110110",
  26275=>"000100011",
  26276=>"101110100",
  26277=>"011101110",
  26278=>"110110000",
  26279=>"010010010",
  26280=>"100010110",
  26281=>"000001101",
  26282=>"000100011",
  26283=>"100111011",
  26284=>"010111001",
  26285=>"011110100",
  26286=>"111101011",
  26287=>"101101111",
  26288=>"001100110",
  26289=>"111000100",
  26290=>"100110001",
  26291=>"000100001",
  26292=>"110010110",
  26293=>"010011100",
  26294=>"001001100",
  26295=>"000100010",
  26296=>"000111001",
  26297=>"110011000",
  26298=>"100011100",
  26299=>"000010100",
  26300=>"111010010",
  26301=>"111100011",
  26302=>"111010000",
  26303=>"010000111",
  26304=>"010010111",
  26305=>"111010000",
  26306=>"111110011",
  26307=>"010010101",
  26308=>"100100101",
  26309=>"011000111",
  26310=>"011100010",
  26311=>"000000000",
  26312=>"011010101",
  26313=>"110100001",
  26314=>"101100101",
  26315=>"110001101",
  26316=>"000100010",
  26317=>"110100001",
  26318=>"110011010",
  26319=>"000000000",
  26320=>"000100010",
  26321=>"000000011",
  26322=>"001000111",
  26323=>"011100100",
  26324=>"100010111",
  26325=>"101111000",
  26326=>"101001110",
  26327=>"000001101",
  26328=>"111011001",
  26329=>"111001100",
  26330=>"101110010",
  26331=>"100010101",
  26332=>"000000001",
  26333=>"000010011",
  26334=>"010011111",
  26335=>"011000001",
  26336=>"100000000",
  26337=>"111110000",
  26338=>"101111111",
  26339=>"000111000",
  26340=>"001000000",
  26341=>"101100110",
  26342=>"001010001",
  26343=>"100111100",
  26344=>"000000001",
  26345=>"101110111",
  26346=>"111111111",
  26347=>"100111000",
  26348=>"000000001",
  26349=>"011110111",
  26350=>"000111110",
  26351=>"111100011",
  26352=>"110010111",
  26353=>"010111011",
  26354=>"110000100",
  26355=>"100010100",
  26356=>"011100000",
  26357=>"100100110",
  26358=>"011001111",
  26359=>"000000001",
  26360=>"010111000",
  26361=>"001100011",
  26362=>"010111000",
  26363=>"111100100",
  26364=>"100010101",
  26365=>"010101011",
  26366=>"100011100",
  26367=>"000001101",
  26368=>"000100100",
  26369=>"110100100",
  26370=>"101100011",
  26371=>"101100111",
  26372=>"101000010",
  26373=>"011001000",
  26374=>"001011110",
  26375=>"011100011",
  26376=>"010100010",
  26377=>"001010111",
  26378=>"110111000",
  26379=>"111011101",
  26380=>"111001100",
  26381=>"100110000",
  26382=>"010011001",
  26383=>"110110100",
  26384=>"010110110",
  26385=>"111010100",
  26386=>"000001011",
  26387=>"101011111",
  26388=>"110110101",
  26389=>"111100110",
  26390=>"100111110",
  26391=>"010101000",
  26392=>"001001000",
  26393=>"001101000",
  26394=>"110010110",
  26395=>"100001110",
  26396=>"011101010",
  26397=>"110011111",
  26398=>"101000001",
  26399=>"010101011",
  26400=>"011111110",
  26401=>"100100100",
  26402=>"111111101",
  26403=>"011000110",
  26404=>"011110110",
  26405=>"110011101",
  26406=>"010001100",
  26407=>"101001011",
  26408=>"100111110",
  26409=>"111010010",
  26410=>"011011010",
  26411=>"111101111",
  26412=>"010101000",
  26413=>"000101111",
  26414=>"110110100",
  26415=>"110000100",
  26416=>"101010011",
  26417=>"000100011",
  26418=>"010000010",
  26419=>"110101100",
  26420=>"110010000",
  26421=>"100110111",
  26422=>"100001110",
  26423=>"001110101",
  26424=>"010101011",
  26425=>"000101011",
  26426=>"001011101",
  26427=>"001000101",
  26428=>"010010110",
  26429=>"000001110",
  26430=>"111010010",
  26431=>"101011110",
  26432=>"100011111",
  26433=>"011100011",
  26434=>"001111101",
  26435=>"000101000",
  26436=>"100101010",
  26437=>"110110010",
  26438=>"000001001",
  26439=>"100000010",
  26440=>"000011001",
  26441=>"110101000",
  26442=>"101000000",
  26443=>"110110101",
  26444=>"110011100",
  26445=>"111101101",
  26446=>"001110110",
  26447=>"111100010",
  26448=>"111000110",
  26449=>"100001011",
  26450=>"011010111",
  26451=>"010001111",
  26452=>"101100010",
  26453=>"000101101",
  26454=>"111000101",
  26455=>"011011111",
  26456=>"011011111",
  26457=>"000110100",
  26458=>"010000001",
  26459=>"100100101",
  26460=>"001111100",
  26461=>"101110001",
  26462=>"001001101",
  26463=>"100100101",
  26464=>"000101000",
  26465=>"101111000",
  26466=>"110111010",
  26467=>"001000000",
  26468=>"110011000",
  26469=>"100000001",
  26470=>"100001000",
  26471=>"010011001",
  26472=>"001010101",
  26473=>"111111010",
  26474=>"110110000",
  26475=>"011111110",
  26476=>"000101100",
  26477=>"001001101",
  26478=>"000100001",
  26479=>"011000101",
  26480=>"110111111",
  26481=>"000000101",
  26482=>"101110011",
  26483=>"111100101",
  26484=>"000011010",
  26485=>"010111100",
  26486=>"010101000",
  26487=>"101011100",
  26488=>"110111010",
  26489=>"000000101",
  26490=>"110101110",
  26491=>"000101001",
  26492=>"000010110",
  26493=>"011010010",
  26494=>"101110111",
  26495=>"101110111",
  26496=>"010111101",
  26497=>"101010110",
  26498=>"010110001",
  26499=>"111010110",
  26500=>"110011011",
  26501=>"110101111",
  26502=>"000010110",
  26503=>"111001010",
  26504=>"011101101",
  26505=>"101011101",
  26506=>"100111101",
  26507=>"011010001",
  26508=>"111110010",
  26509=>"001101101",
  26510=>"101100001",
  26511=>"101101101",
  26512=>"000101110",
  26513=>"111001001",
  26514=>"010000101",
  26515=>"110000101",
  26516=>"010010001",
  26517=>"010000001",
  26518=>"111100100",
  26519=>"000110000",
  26520=>"111000101",
  26521=>"111101001",
  26522=>"101000101",
  26523=>"000011111",
  26524=>"010101111",
  26525=>"110010110",
  26526=>"001111110",
  26527=>"110111111",
  26528=>"100100100",
  26529=>"001101001",
  26530=>"101011010",
  26531=>"010100010",
  26532=>"111110110",
  26533=>"110110111",
  26534=>"000100001",
  26535=>"000110000",
  26536=>"001100001",
  26537=>"111010111",
  26538=>"011001000",
  26539=>"001110011",
  26540=>"001010000",
  26541=>"100010111",
  26542=>"101001101",
  26543=>"001111111",
  26544=>"110011011",
  26545=>"111100010",
  26546=>"011011111",
  26547=>"111000011",
  26548=>"101110111",
  26549=>"100101011",
  26550=>"001011010",
  26551=>"101100111",
  26552=>"110110001",
  26553=>"100101000",
  26554=>"010011001",
  26555=>"000000011",
  26556=>"111010100",
  26557=>"001100011",
  26558=>"100011000",
  26559=>"110110001",
  26560=>"011100001",
  26561=>"111001110",
  26562=>"011101000",
  26563=>"011101100",
  26564=>"011100010",
  26565=>"110101111",
  26566=>"101101011",
  26567=>"110111011",
  26568=>"011100010",
  26569=>"010100010",
  26570=>"001110110",
  26571=>"100001001",
  26572=>"111100010",
  26573=>"110010100",
  26574=>"100010001",
  26575=>"100101011",
  26576=>"001110001",
  26577=>"011110110",
  26578=>"001100110",
  26579=>"010000000",
  26580=>"000011101",
  26581=>"001101011",
  26582=>"000001010",
  26583=>"010101011",
  26584=>"111111001",
  26585=>"101100011",
  26586=>"110110011",
  26587=>"001100000",
  26588=>"000000111",
  26589=>"000101100",
  26590=>"111111100",
  26591=>"100111111",
  26592=>"011010100",
  26593=>"101000111",
  26594=>"000111000",
  26595=>"101111010",
  26596=>"101000000",
  26597=>"111101101",
  26598=>"100100110",
  26599=>"001010010",
  26600=>"101001101",
  26601=>"101010000",
  26602=>"010110000",
  26603=>"110011110",
  26604=>"010001000",
  26605=>"010100000",
  26606=>"000100001",
  26607=>"000010110",
  26608=>"001011111",
  26609=>"011001101",
  26610=>"100101110",
  26611=>"100011000",
  26612=>"111110101",
  26613=>"011010000",
  26614=>"001110101",
  26615=>"010001001",
  26616=>"011001100",
  26617=>"010000010",
  26618=>"101000110",
  26619=>"110100000",
  26620=>"000100010",
  26621=>"101010001",
  26622=>"111100011",
  26623=>"100011100",
  26624=>"001110001",
  26625=>"100110011",
  26626=>"100111100",
  26627=>"110101100",
  26628=>"110111100",
  26629=>"010100000",
  26630=>"001010110",
  26631=>"001000111",
  26632=>"010111011",
  26633=>"101100011",
  26634=>"101001110",
  26635=>"111111111",
  26636=>"110000001",
  26637=>"010010111",
  26638=>"001001011",
  26639=>"010100111",
  26640=>"010110111",
  26641=>"001000110",
  26642=>"100001000",
  26643=>"011101100",
  26644=>"010101001",
  26645=>"000110111",
  26646=>"111101100",
  26647=>"000100110",
  26648=>"111011100",
  26649=>"000010010",
  26650=>"111001010",
  26651=>"010101010",
  26652=>"000001111",
  26653=>"111111111",
  26654=>"100110101",
  26655=>"010010101",
  26656=>"111000101",
  26657=>"001111010",
  26658=>"001010000",
  26659=>"101110001",
  26660=>"010100011",
  26661=>"000011011",
  26662=>"100100010",
  26663=>"111111111",
  26664=>"001101010",
  26665=>"010110101",
  26666=>"010110000",
  26667=>"001100000",
  26668=>"110011000",
  26669=>"111011110",
  26670=>"101100000",
  26671=>"111011010",
  26672=>"000110000",
  26673=>"111000010",
  26674=>"001110111",
  26675=>"000100110",
  26676=>"000110100",
  26677=>"100010110",
  26678=>"100111101",
  26679=>"001101011",
  26680=>"000001110",
  26681=>"101000111",
  26682=>"000011111",
  26683=>"000010000",
  26684=>"111010000",
  26685=>"010011110",
  26686=>"011101000",
  26687=>"010110100",
  26688=>"111110100",
  26689=>"000101100",
  26690=>"101111000",
  26691=>"100000110",
  26692=>"001011000",
  26693=>"001011101",
  26694=>"010111101",
  26695=>"010111000",
  26696=>"001100011",
  26697=>"011111001",
  26698=>"101111010",
  26699=>"101011000",
  26700=>"010111111",
  26701=>"110011100",
  26702=>"000100000",
  26703=>"100001011",
  26704=>"010100001",
  26705=>"100000000",
  26706=>"101100000",
  26707=>"000110110",
  26708=>"110000111",
  26709=>"001100000",
  26710=>"000111000",
  26711=>"001101010",
  26712=>"010011001",
  26713=>"110101101",
  26714=>"100011010",
  26715=>"110001000",
  26716=>"110100110",
  26717=>"000001111",
  26718=>"010001111",
  26719=>"000100011",
  26720=>"010000111",
  26721=>"000100111",
  26722=>"111101011",
  26723=>"000110000",
  26724=>"101001000",
  26725=>"100011111",
  26726=>"011110011",
  26727=>"000110111",
  26728=>"001100101",
  26729=>"010101011",
  26730=>"011001011",
  26731=>"001110100",
  26732=>"111101011",
  26733=>"100110010",
  26734=>"011111110",
  26735=>"101001001",
  26736=>"001000111",
  26737=>"101000100",
  26738=>"110011110",
  26739=>"010011100",
  26740=>"110110011",
  26741=>"110111011",
  26742=>"111100001",
  26743=>"111011000",
  26744=>"111011000",
  26745=>"011001111",
  26746=>"111001000",
  26747=>"010111001",
  26748=>"110101101",
  26749=>"010010101",
  26750=>"110000011",
  26751=>"001111111",
  26752=>"111001001",
  26753=>"000010000",
  26754=>"000010010",
  26755=>"110001000",
  26756=>"101001001",
  26757=>"111000010",
  26758=>"111000010",
  26759=>"110110001",
  26760=>"010100111",
  26761=>"001000010",
  26762=>"110001001",
  26763=>"100010011",
  26764=>"111111000",
  26765=>"111100111",
  26766=>"100111000",
  26767=>"100011000",
  26768=>"001010110",
  26769=>"011001000",
  26770=>"101011000",
  26771=>"100001011",
  26772=>"000001010",
  26773=>"010110010",
  26774=>"100001010",
  26775=>"111000011",
  26776=>"000010111",
  26777=>"011011110",
  26778=>"101101111",
  26779=>"101000111",
  26780=>"100100010",
  26781=>"100010001",
  26782=>"110011011",
  26783=>"010101000",
  26784=>"101100100",
  26785=>"011101010",
  26786=>"100000111",
  26787=>"110100110",
  26788=>"111010111",
  26789=>"101111110",
  26790=>"000000000",
  26791=>"010111010",
  26792=>"110000010",
  26793=>"111110011",
  26794=>"011000010",
  26795=>"000111001",
  26796=>"101111111",
  26797=>"110001010",
  26798=>"101100000",
  26799=>"100111000",
  26800=>"011111101",
  26801=>"110100101",
  26802=>"011000110",
  26803=>"001101111",
  26804=>"010001000",
  26805=>"000111100",
  26806=>"110000010",
  26807=>"100011100",
  26808=>"011010111",
  26809=>"101001001",
  26810=>"001100010",
  26811=>"000001011",
  26812=>"010010010",
  26813=>"001110010",
  26814=>"110110001",
  26815=>"111100100",
  26816=>"010111111",
  26817=>"100010010",
  26818=>"111010000",
  26819=>"101110000",
  26820=>"101011101",
  26821=>"000100001",
  26822=>"101101110",
  26823=>"001001111",
  26824=>"111100110",
  26825=>"101110010",
  26826=>"010101001",
  26827=>"001100110",
  26828=>"010110100",
  26829=>"111000011",
  26830=>"100101001",
  26831=>"001010000",
  26832=>"110000010",
  26833=>"101100101",
  26834=>"001000101",
  26835=>"010001111",
  26836=>"101011100",
  26837=>"010111001",
  26838=>"110111101",
  26839=>"011011011",
  26840=>"011010100",
  26841=>"111010000",
  26842=>"010000100",
  26843=>"011011101",
  26844=>"000110001",
  26845=>"101010110",
  26846=>"101100110",
  26847=>"111011011",
  26848=>"001010111",
  26849=>"000001100",
  26850=>"100011101",
  26851=>"110000000",
  26852=>"000011111",
  26853=>"110000010",
  26854=>"100000110",
  26855=>"010001100",
  26856=>"000010011",
  26857=>"011111100",
  26858=>"111111001",
  26859=>"000100111",
  26860=>"010000111",
  26861=>"101101111",
  26862=>"001001010",
  26863=>"001000110",
  26864=>"101110100",
  26865=>"010100101",
  26866=>"011100011",
  26867=>"101011011",
  26868=>"001111101",
  26869=>"110101010",
  26870=>"101101001",
  26871=>"000000011",
  26872=>"011001011",
  26873=>"101110000",
  26874=>"011111101",
  26875=>"000110111",
  26876=>"000011010",
  26877=>"111011000",
  26878=>"000101000",
  26879=>"101011101",
  26880=>"011101010",
  26881=>"101111110",
  26882=>"101011001",
  26883=>"001100111",
  26884=>"000111011",
  26885=>"011101001",
  26886=>"011110101",
  26887=>"011100011",
  26888=>"100001001",
  26889=>"001110101",
  26890=>"000000110",
  26891=>"110101000",
  26892=>"100100100",
  26893=>"101101001",
  26894=>"001100000",
  26895=>"100101011",
  26896=>"000100001",
  26897=>"100011110",
  26898=>"011110110",
  26899=>"010001110",
  26900=>"110101010",
  26901=>"111010101",
  26902=>"100001110",
  26903=>"100101110",
  26904=>"010011101",
  26905=>"001101001",
  26906=>"000111101",
  26907=>"010100011",
  26908=>"110010010",
  26909=>"001000110",
  26910=>"000110110",
  26911=>"010110111",
  26912=>"001001110",
  26913=>"110111111",
  26914=>"011110100",
  26915=>"100100110",
  26916=>"000111011",
  26917=>"100001110",
  26918=>"011100100",
  26919=>"010000100",
  26920=>"101110101",
  26921=>"100010101",
  26922=>"001001010",
  26923=>"110000010",
  26924=>"011111011",
  26925=>"110000001",
  26926=>"011010110",
  26927=>"100000101",
  26928=>"111000110",
  26929=>"010000101",
  26930=>"010110011",
  26931=>"110011000",
  26932=>"100100000",
  26933=>"010100001",
  26934=>"111101110",
  26935=>"110000001",
  26936=>"011011100",
  26937=>"111100110",
  26938=>"011010010",
  26939=>"111001000",
  26940=>"001000101",
  26941=>"111110111",
  26942=>"101001011",
  26943=>"111001001",
  26944=>"111111010",
  26945=>"100100011",
  26946=>"110110010",
  26947=>"101101011",
  26948=>"110100001",
  26949=>"100001100",
  26950=>"011101111",
  26951=>"000010011",
  26952=>"011100010",
  26953=>"111001110",
  26954=>"101011100",
  26955=>"110011010",
  26956=>"011111001",
  26957=>"111110111",
  26958=>"011111001",
  26959=>"100010001",
  26960=>"101001100",
  26961=>"110100001",
  26962=>"000111011",
  26963=>"001000010",
  26964=>"100000111",
  26965=>"101100001",
  26966=>"110000101",
  26967=>"100011111",
  26968=>"011111111",
  26969=>"001100100",
  26970=>"001100000",
  26971=>"010010101",
  26972=>"100000111",
  26973=>"010100000",
  26974=>"001110010",
  26975=>"011110110",
  26976=>"010100110",
  26977=>"010000010",
  26978=>"101001101",
  26979=>"101000111",
  26980=>"111000111",
  26981=>"101011011",
  26982=>"111011101",
  26983=>"011011101",
  26984=>"011111011",
  26985=>"010100111",
  26986=>"111111111",
  26987=>"001100101",
  26988=>"110010110",
  26989=>"110100111",
  26990=>"000000111",
  26991=>"011100000",
  26992=>"001110011",
  26993=>"000010010",
  26994=>"010111110",
  26995=>"000000100",
  26996=>"101010110",
  26997=>"110001001",
  26998=>"010010111",
  26999=>"010000010",
  27000=>"000100101",
  27001=>"000010011",
  27002=>"100110101",
  27003=>"011101110",
  27004=>"000101001",
  27005=>"010011101",
  27006=>"011110010",
  27007=>"100111001",
  27008=>"101000111",
  27009=>"111010000",
  27010=>"001101100",
  27011=>"000001110",
  27012=>"010111100",
  27013=>"001010000",
  27014=>"001111011",
  27015=>"111011010",
  27016=>"000111101",
  27017=>"100000010",
  27018=>"111111101",
  27019=>"000110011",
  27020=>"100000111",
  27021=>"001001011",
  27022=>"111010101",
  27023=>"111100100",
  27024=>"010111101",
  27025=>"001000010",
  27026=>"001000111",
  27027=>"111010010",
  27028=>"100001010",
  27029=>"001100001",
  27030=>"000100000",
  27031=>"100000011",
  27032=>"111101110",
  27033=>"000111011",
  27034=>"101110011",
  27035=>"101100111",
  27036=>"010110001",
  27037=>"011101101",
  27038=>"010000000",
  27039=>"111000110",
  27040=>"101100001",
  27041=>"101001111",
  27042=>"000110000",
  27043=>"110100111",
  27044=>"010011100",
  27045=>"110000010",
  27046=>"000111111",
  27047=>"011001101",
  27048=>"001111111",
  27049=>"101101001",
  27050=>"111100101",
  27051=>"000100101",
  27052=>"011011110",
  27053=>"011011011",
  27054=>"100010001",
  27055=>"011000000",
  27056=>"000010011",
  27057=>"110101110",
  27058=>"011101101",
  27059=>"000100111",
  27060=>"101111010",
  27061=>"000111011",
  27062=>"100100111",
  27063=>"011110101",
  27064=>"100111001",
  27065=>"100110000",
  27066=>"001000001",
  27067=>"101110111",
  27068=>"111010001",
  27069=>"100001111",
  27070=>"101001010",
  27071=>"110011000",
  27072=>"011000100",
  27073=>"001111100",
  27074=>"100010100",
  27075=>"011100000",
  27076=>"101110101",
  27077=>"110101011",
  27078=>"111100101",
  27079=>"000000011",
  27080=>"010011111",
  27081=>"100110010",
  27082=>"000100010",
  27083=>"010011101",
  27084=>"010001010",
  27085=>"111000100",
  27086=>"100111001",
  27087=>"111000111",
  27088=>"001101100",
  27089=>"101010010",
  27090=>"110010011",
  27091=>"110101010",
  27092=>"001001001",
  27093=>"001001110",
  27094=>"000100110",
  27095=>"000011101",
  27096=>"100111100",
  27097=>"101100011",
  27098=>"110101001",
  27099=>"101110111",
  27100=>"010010010",
  27101=>"101010100",
  27102=>"111001111",
  27103=>"110111111",
  27104=>"110111110",
  27105=>"100010110",
  27106=>"000100010",
  27107=>"000110011",
  27108=>"100101010",
  27109=>"011100000",
  27110=>"000000101",
  27111=>"100011101",
  27112=>"110001111",
  27113=>"001010001",
  27114=>"011001111",
  27115=>"000001111",
  27116=>"011011001",
  27117=>"011010100",
  27118=>"001001000",
  27119=>"111000001",
  27120=>"011101000",
  27121=>"111101111",
  27122=>"110110010",
  27123=>"011010010",
  27124=>"110010110",
  27125=>"001000001",
  27126=>"001101010",
  27127=>"110110011",
  27128=>"000000011",
  27129=>"111001000",
  27130=>"100010011",
  27131=>"110011001",
  27132=>"100000101",
  27133=>"111000010",
  27134=>"011110010",
  27135=>"110001011",
  27136=>"111101010",
  27137=>"111111111",
  27138=>"011010101",
  27139=>"101010100",
  27140=>"101111111",
  27141=>"010000101",
  27142=>"000011100",
  27143=>"100001000",
  27144=>"111101001",
  27145=>"010101101",
  27146=>"110111111",
  27147=>"010110100",
  27148=>"000110110",
  27149=>"101010111",
  27150=>"001011100",
  27151=>"100101010",
  27152=>"011100010",
  27153=>"100110100",
  27154=>"010001111",
  27155=>"111101101",
  27156=>"100101101",
  27157=>"011000100",
  27158=>"000010000",
  27159=>"111110011",
  27160=>"001110001",
  27161=>"001101010",
  27162=>"011111000",
  27163=>"011111100",
  27164=>"000010010",
  27165=>"011001110",
  27166=>"111000001",
  27167=>"111110000",
  27168=>"110100100",
  27169=>"001111110",
  27170=>"100011000",
  27171=>"101010011",
  27172=>"011101101",
  27173=>"011101111",
  27174=>"110010010",
  27175=>"100011000",
  27176=>"010001110",
  27177=>"111001110",
  27178=>"100010001",
  27179=>"011001101",
  27180=>"010010001",
  27181=>"110000010",
  27182=>"101111001",
  27183=>"011101011",
  27184=>"011110001",
  27185=>"111111001",
  27186=>"001110100",
  27187=>"101010100",
  27188=>"011010111",
  27189=>"101000100",
  27190=>"000001011",
  27191=>"110011100",
  27192=>"110011010",
  27193=>"111111000",
  27194=>"011101100",
  27195=>"000110101",
  27196=>"111100111",
  27197=>"100001010",
  27198=>"101001110",
  27199=>"011000010",
  27200=>"110111011",
  27201=>"100010100",
  27202=>"100000001",
  27203=>"010110001",
  27204=>"101001101",
  27205=>"101011000",
  27206=>"000100001",
  27207=>"001000010",
  27208=>"101101011",
  27209=>"011001100",
  27210=>"110111100",
  27211=>"101001110",
  27212=>"011011100",
  27213=>"010000110",
  27214=>"110100000",
  27215=>"011101001",
  27216=>"001001110",
  27217=>"110111001",
  27218=>"111101110",
  27219=>"101011000",
  27220=>"110111110",
  27221=>"011001000",
  27222=>"000010000",
  27223=>"000000111",
  27224=>"111001010",
  27225=>"101011001",
  27226=>"001110110",
  27227=>"100001000",
  27228=>"101000100",
  27229=>"100001000",
  27230=>"000101111",
  27231=>"101100100",
  27232=>"000011000",
  27233=>"000010101",
  27234=>"000011011",
  27235=>"100100001",
  27236=>"110011100",
  27237=>"001011101",
  27238=>"010111111",
  27239=>"010000010",
  27240=>"111101100",
  27241=>"111000110",
  27242=>"011100100",
  27243=>"000001011",
  27244=>"001101001",
  27245=>"011011111",
  27246=>"011111111",
  27247=>"100111001",
  27248=>"000100000",
  27249=>"001111100",
  27250=>"000101000",
  27251=>"110110101",
  27252=>"010000111",
  27253=>"100011011",
  27254=>"100001011",
  27255=>"001011011",
  27256=>"011000100",
  27257=>"110010010",
  27258=>"010001000",
  27259=>"000011100",
  27260=>"001001010",
  27261=>"111100111",
  27262=>"110101001",
  27263=>"000100011",
  27264=>"101111011",
  27265=>"010000000",
  27266=>"000000111",
  27267=>"101111001",
  27268=>"100001100",
  27269=>"010011101",
  27270=>"011011111",
  27271=>"010000011",
  27272=>"001010100",
  27273=>"001101000",
  27274=>"010000101",
  27275=>"111111101",
  27276=>"101001100",
  27277=>"010100000",
  27278=>"011110000",
  27279=>"011011111",
  27280=>"111100001",
  27281=>"100001101",
  27282=>"010010111",
  27283=>"111111001",
  27284=>"111100110",
  27285=>"100001101",
  27286=>"100010001",
  27287=>"101001000",
  27288=>"010001101",
  27289=>"101011101",
  27290=>"001110101",
  27291=>"101111111",
  27292=>"110000011",
  27293=>"101010011",
  27294=>"000010001",
  27295=>"101011100",
  27296=>"011101110",
  27297=>"010001010",
  27298=>"111101111",
  27299=>"000000001",
  27300=>"100000001",
  27301=>"100001110",
  27302=>"101100011",
  27303=>"000000001",
  27304=>"011010000",
  27305=>"100100111",
  27306=>"001111101",
  27307=>"010110110",
  27308=>"000010110",
  27309=>"010011001",
  27310=>"101100000",
  27311=>"100100010",
  27312=>"010001110",
  27313=>"011011010",
  27314=>"111111001",
  27315=>"011001000",
  27316=>"011100010",
  27317=>"011101000",
  27318=>"101001011",
  27319=>"101101011",
  27320=>"100000110",
  27321=>"111001010",
  27322=>"100000001",
  27323=>"110000101",
  27324=>"000110000",
  27325=>"000011111",
  27326=>"110001111",
  27327=>"000010110",
  27328=>"100010011",
  27329=>"001001010",
  27330=>"100111111",
  27331=>"010001010",
  27332=>"100101111",
  27333=>"010101110",
  27334=>"010111010",
  27335=>"101000001",
  27336=>"110101100",
  27337=>"011000001",
  27338=>"001000001",
  27339=>"011011011",
  27340=>"101111100",
  27341=>"010100111",
  27342=>"110101001",
  27343=>"000001100",
  27344=>"111111011",
  27345=>"010010000",
  27346=>"010011111",
  27347=>"000100101",
  27348=>"101110111",
  27349=>"001000111",
  27350=>"000011100",
  27351=>"100010000",
  27352=>"001001110",
  27353=>"000010001",
  27354=>"010000000",
  27355=>"110100111",
  27356=>"101001011",
  27357=>"100101100",
  27358=>"011000101",
  27359=>"001010111",
  27360=>"101011101",
  27361=>"000110001",
  27362=>"110101010",
  27363=>"000000110",
  27364=>"101110101",
  27365=>"010100000",
  27366=>"101010010",
  27367=>"100000000",
  27368=>"000001000",
  27369=>"111101101",
  27370=>"010110110",
  27371=>"101101110",
  27372=>"001111100",
  27373=>"101000110",
  27374=>"110100001",
  27375=>"010100011",
  27376=>"110000111",
  27377=>"111100100",
  27378=>"101010111",
  27379=>"100101110",
  27380=>"110101011",
  27381=>"001110100",
  27382=>"011000111",
  27383=>"111000010",
  27384=>"110000000",
  27385=>"111010001",
  27386=>"001011110",
  27387=>"011011000",
  27388=>"110011101",
  27389=>"101111011",
  27390=>"010010000",
  27391=>"010100100",
  27392=>"100011010",
  27393=>"010111001",
  27394=>"111110000",
  27395=>"101111001",
  27396=>"010110100",
  27397=>"100010011",
  27398=>"000111011",
  27399=>"001100011",
  27400=>"001100010",
  27401=>"011001011",
  27402=>"110011011",
  27403=>"010001010",
  27404=>"010111011",
  27405=>"000000000",
  27406=>"111111001",
  27407=>"000011001",
  27408=>"010001101",
  27409=>"110101101",
  27410=>"001010011",
  27411=>"001101001",
  27412=>"110111111",
  27413=>"001010011",
  27414=>"001101111",
  27415=>"000000011",
  27416=>"110001010",
  27417=>"110110010",
  27418=>"101111011",
  27419=>"011010101",
  27420=>"010101111",
  27421=>"010110001",
  27422=>"100011010",
  27423=>"101001010",
  27424=>"111111100",
  27425=>"011000010",
  27426=>"001100000",
  27427=>"110011001",
  27428=>"100000000",
  27429=>"110100001",
  27430=>"100100011",
  27431=>"010010101",
  27432=>"101011101",
  27433=>"000011111",
  27434=>"110100101",
  27435=>"111110000",
  27436=>"001101011",
  27437=>"001101011",
  27438=>"010111000",
  27439=>"111111010",
  27440=>"111000100",
  27441=>"000000011",
  27442=>"001100010",
  27443=>"001111100",
  27444=>"010100000",
  27445=>"010111101",
  27446=>"011000000",
  27447=>"000000101",
  27448=>"100011010",
  27449=>"000110001",
  27450=>"101110100",
  27451=>"010101110",
  27452=>"001000000",
  27453=>"110101001",
  27454=>"101001010",
  27455=>"010101110",
  27456=>"010001000",
  27457=>"111001001",
  27458=>"111000110",
  27459=>"010010111",
  27460=>"111110000",
  27461=>"101101110",
  27462=>"101111100",
  27463=>"010101101",
  27464=>"111010011",
  27465=>"110111111",
  27466=>"110110001",
  27467=>"100111101",
  27468=>"100000100",
  27469=>"101010010",
  27470=>"111011001",
  27471=>"001000011",
  27472=>"111100110",
  27473=>"001000110",
  27474=>"101001011",
  27475=>"011000000",
  27476=>"000000011",
  27477=>"010100011",
  27478=>"011001100",
  27479=>"100011000",
  27480=>"110011110",
  27481=>"110110110",
  27482=>"001000110",
  27483=>"101001011",
  27484=>"000101101",
  27485=>"110001000",
  27486=>"000100100",
  27487=>"001010011",
  27488=>"011001011",
  27489=>"010000011",
  27490=>"101111101",
  27491=>"010111110",
  27492=>"101010000",
  27493=>"110101101",
  27494=>"011100100",
  27495=>"110111010",
  27496=>"000110001",
  27497=>"111001111",
  27498=>"001001010",
  27499=>"100110111",
  27500=>"010010100",
  27501=>"101100001",
  27502=>"000101111",
  27503=>"100111011",
  27504=>"011101011",
  27505=>"100111101",
  27506=>"010100101",
  27507=>"100100000",
  27508=>"110111100",
  27509=>"010010101",
  27510=>"111010101",
  27511=>"101000101",
  27512=>"001111010",
  27513=>"000000111",
  27514=>"111010111",
  27515=>"011101110",
  27516=>"010000001",
  27517=>"100000001",
  27518=>"101000000",
  27519=>"110000000",
  27520=>"110111001",
  27521=>"001000111",
  27522=>"010111001",
  27523=>"000000101",
  27524=>"001110111",
  27525=>"110110011",
  27526=>"110011101",
  27527=>"110110100",
  27528=>"011111011",
  27529=>"000010001",
  27530=>"110101100",
  27531=>"011011011",
  27532=>"110001100",
  27533=>"110100101",
  27534=>"011000100",
  27535=>"101101111",
  27536=>"001100010",
  27537=>"010100100",
  27538=>"000001010",
  27539=>"101000010",
  27540=>"110101010",
  27541=>"000011101",
  27542=>"100101111",
  27543=>"111110110",
  27544=>"110111000",
  27545=>"100101101",
  27546=>"111000001",
  27547=>"000110010",
  27548=>"100101011",
  27549=>"110101110",
  27550=>"110101111",
  27551=>"000010100",
  27552=>"010011110",
  27553=>"001000111",
  27554=>"001111100",
  27555=>"011100010",
  27556=>"000001011",
  27557=>"101011101",
  27558=>"001101101",
  27559=>"011110001",
  27560=>"100110001",
  27561=>"011100110",
  27562=>"011111110",
  27563=>"101011111",
  27564=>"111101111",
  27565=>"101010010",
  27566=>"100100010",
  27567=>"001000100",
  27568=>"010011010",
  27569=>"111101100",
  27570=>"011000001",
  27571=>"000110011",
  27572=>"111001100",
  27573=>"101000111",
  27574=>"010000001",
  27575=>"001001110",
  27576=>"000000101",
  27577=>"001100010",
  27578=>"011001110",
  27579=>"101110100",
  27580=>"011000100",
  27581=>"100000110",
  27582=>"110101000",
  27583=>"000100000",
  27584=>"000000001",
  27585=>"000110001",
  27586=>"111101010",
  27587=>"101100000",
  27588=>"110101010",
  27589=>"001011111",
  27590=>"111110100",
  27591=>"111110000",
  27592=>"100010110",
  27593=>"001101010",
  27594=>"101001100",
  27595=>"001101011",
  27596=>"101100100",
  27597=>"010100111",
  27598=>"111110010",
  27599=>"011111010",
  27600=>"101111110",
  27601=>"011100010",
  27602=>"100000111",
  27603=>"100011001",
  27604=>"101110100",
  27605=>"001111110",
  27606=>"110000111",
  27607=>"110010101",
  27608=>"100000100",
  27609=>"100011010",
  27610=>"001001000",
  27611=>"100100001",
  27612=>"101000001",
  27613=>"100011111",
  27614=>"100101111",
  27615=>"001111101",
  27616=>"000000101",
  27617=>"001011101",
  27618=>"001101101",
  27619=>"101101100",
  27620=>"010100011",
  27621=>"000100011",
  27622=>"100111000",
  27623=>"000000111",
  27624=>"100101000",
  27625=>"111111011",
  27626=>"101110100",
  27627=>"110111111",
  27628=>"010110001",
  27629=>"101000011",
  27630=>"000001111",
  27631=>"010101011",
  27632=>"001001010",
  27633=>"010000011",
  27634=>"001100100",
  27635=>"101000101",
  27636=>"100100111",
  27637=>"010011100",
  27638=>"101010110",
  27639=>"011111011",
  27640=>"100110011",
  27641=>"000010000",
  27642=>"011101000",
  27643=>"011101110",
  27644=>"100100000",
  27645=>"010110110",
  27646=>"010111011",
  27647=>"001001101",
  27648=>"100001101",
  27649=>"110011001",
  27650=>"010100111",
  27651=>"111011110",
  27652=>"101000100",
  27653=>"010000000",
  27654=>"101010001",
  27655=>"001100000",
  27656=>"111000110",
  27657=>"101011001",
  27658=>"000010111",
  27659=>"101101001",
  27660=>"110110000",
  27661=>"011011010",
  27662=>"010111101",
  27663=>"001111000",
  27664=>"110001100",
  27665=>"000111010",
  27666=>"000000010",
  27667=>"100010111",
  27668=>"011010001",
  27669=>"010000111",
  27670=>"110011000",
  27671=>"010110100",
  27672=>"111110000",
  27673=>"101011110",
  27674=>"000001001",
  27675=>"101010011",
  27676=>"110111110",
  27677=>"000000111",
  27678=>"110010110",
  27679=>"111001100",
  27680=>"001100101",
  27681=>"101110010",
  27682=>"000101100",
  27683=>"000110100",
  27684=>"111011000",
  27685=>"010000111",
  27686=>"101011000",
  27687=>"110110001",
  27688=>"000100100",
  27689=>"101100111",
  27690=>"010100011",
  27691=>"000001001",
  27692=>"101110101",
  27693=>"001100001",
  27694=>"000101111",
  27695=>"010010000",
  27696=>"101101000",
  27697=>"000010111",
  27698=>"110010101",
  27699=>"000010011",
  27700=>"111000001",
  27701=>"111110001",
  27702=>"000100000",
  27703=>"010000010",
  27704=>"000100001",
  27705=>"001101001",
  27706=>"010010100",
  27707=>"011010100",
  27708=>"101101000",
  27709=>"101110111",
  27710=>"100000001",
  27711=>"110100101",
  27712=>"111100011",
  27713=>"110011110",
  27714=>"001000001",
  27715=>"110001010",
  27716=>"000110001",
  27717=>"000000000",
  27718=>"110000011",
  27719=>"010000000",
  27720=>"101111111",
  27721=>"100110101",
  27722=>"010110010",
  27723=>"111101010",
  27724=>"010100001",
  27725=>"000110001",
  27726=>"010100111",
  27727=>"000101101",
  27728=>"000011010",
  27729=>"111000010",
  27730=>"000100101",
  27731=>"110101011",
  27732=>"110001011",
  27733=>"110100011",
  27734=>"111100100",
  27735=>"101101000",
  27736=>"111100000",
  27737=>"100001110",
  27738=>"110011000",
  27739=>"111110100",
  27740=>"111001000",
  27741=>"001111001",
  27742=>"001011110",
  27743=>"001100010",
  27744=>"001001011",
  27745=>"001100000",
  27746=>"001100110",
  27747=>"101001010",
  27748=>"100100101",
  27749=>"110100001",
  27750=>"111001010",
  27751=>"110110100",
  27752=>"000010010",
  27753=>"100000010",
  27754=>"010101111",
  27755=>"011101001",
  27756=>"010111100",
  27757=>"001001010",
  27758=>"001110101",
  27759=>"001010101",
  27760=>"101100111",
  27761=>"100101100",
  27762=>"011000000",
  27763=>"101111110",
  27764=>"110101100",
  27765=>"110110000",
  27766=>"111010001",
  27767=>"001000111",
  27768=>"001101110",
  27769=>"101001000",
  27770=>"111111011",
  27771=>"010000010",
  27772=>"100001011",
  27773=>"010001010",
  27774=>"010001111",
  27775=>"111011000",
  27776=>"010010001",
  27777=>"010110011",
  27778=>"100110110",
  27779=>"001111110",
  27780=>"101000101",
  27781=>"101000000",
  27782=>"111010111",
  27783=>"000100010",
  27784=>"000001010",
  27785=>"110111011",
  27786=>"000001100",
  27787=>"001010100",
  27788=>"100110001",
  27789=>"000011111",
  27790=>"111110100",
  27791=>"000111110",
  27792=>"111111111",
  27793=>"110000011",
  27794=>"110111000",
  27795=>"110011110",
  27796=>"001000001",
  27797=>"000111010",
  27798=>"101001100",
  27799=>"010011000",
  27800=>"000111011",
  27801=>"010111111",
  27802=>"001000100",
  27803=>"110101000",
  27804=>"100010001",
  27805=>"110010000",
  27806=>"001010101",
  27807=>"001000001",
  27808=>"110111111",
  27809=>"100000101",
  27810=>"011101101",
  27811=>"000001000",
  27812=>"010010011",
  27813=>"111011100",
  27814=>"000010001",
  27815=>"111010000",
  27816=>"000010010",
  27817=>"001110111",
  27818=>"001110100",
  27819=>"000100110",
  27820=>"010101010",
  27821=>"010010110",
  27822=>"010011011",
  27823=>"110010000",
  27824=>"100010111",
  27825=>"101110010",
  27826=>"111010011",
  27827=>"110110011",
  27828=>"010000100",
  27829=>"000101101",
  27830=>"110101110",
  27831=>"101101110",
  27832=>"001110100",
  27833=>"001000110",
  27834=>"100010001",
  27835=>"110000101",
  27836=>"011100011",
  27837=>"010110001",
  27838=>"101011100",
  27839=>"110101110",
  27840=>"000010111",
  27841=>"111011001",
  27842=>"111011010",
  27843=>"001011111",
  27844=>"100100110",
  27845=>"100110011",
  27846=>"010011101",
  27847=>"111110100",
  27848=>"000001111",
  27849=>"100101100",
  27850=>"111110001",
  27851=>"000100011",
  27852=>"101001111",
  27853=>"011011101",
  27854=>"101110111",
  27855=>"010101011",
  27856=>"000010010",
  27857=>"111000001",
  27858=>"111100000",
  27859=>"110101100",
  27860=>"100001010",
  27861=>"000010110",
  27862=>"101010110",
  27863=>"001000111",
  27864=>"000001101",
  27865=>"011011111",
  27866=>"010111011",
  27867=>"111111010",
  27868=>"000100111",
  27869=>"011110101",
  27870=>"110011011",
  27871=>"100101000",
  27872=>"011001001",
  27873=>"000101011",
  27874=>"010111000",
  27875=>"111000100",
  27876=>"111111110",
  27877=>"101001100",
  27878=>"111101111",
  27879=>"111011100",
  27880=>"001010011",
  27881=>"010100000",
  27882=>"110001000",
  27883=>"101101110",
  27884=>"101101010",
  27885=>"000100100",
  27886=>"001111010",
  27887=>"100100111",
  27888=>"111100010",
  27889=>"010001010",
  27890=>"011000000",
  27891=>"101111010",
  27892=>"111110100",
  27893=>"111111111",
  27894=>"100110111",
  27895=>"110101111",
  27896=>"011110001",
  27897=>"010001001",
  27898=>"010001100",
  27899=>"110000010",
  27900=>"000000111",
  27901=>"011101110",
  27902=>"101000000",
  27903=>"011101000",
  27904=>"110000010",
  27905=>"011110011",
  27906=>"110000111",
  27907=>"111001010",
  27908=>"010111101",
  27909=>"100110100",
  27910=>"011111110",
  27911=>"100011000",
  27912=>"010110100",
  27913=>"000000100",
  27914=>"110110101",
  27915=>"110110001",
  27916=>"100100001",
  27917=>"100111111",
  27918=>"010001011",
  27919=>"011000100",
  27920=>"110010100",
  27921=>"000001110",
  27922=>"100010001",
  27923=>"110001010",
  27924=>"111110100",
  27925=>"101110101",
  27926=>"110101110",
  27927=>"010111101",
  27928=>"000010001",
  27929=>"000011001",
  27930=>"110010111",
  27931=>"000010000",
  27932=>"000001111",
  27933=>"011001110",
  27934=>"001010011",
  27935=>"101100001",
  27936=>"110110000",
  27937=>"000101000",
  27938=>"110010000",
  27939=>"010111110",
  27940=>"101110101",
  27941=>"011011100",
  27942=>"100000001",
  27943=>"011001010",
  27944=>"011001111",
  27945=>"001110111",
  27946=>"001011001",
  27947=>"011101001",
  27948=>"000111011",
  27949=>"110001100",
  27950=>"000010000",
  27951=>"101000111",
  27952=>"101110100",
  27953=>"111101111",
  27954=>"001000010",
  27955=>"111100010",
  27956=>"000100000",
  27957=>"101100111",
  27958=>"110111100",
  27959=>"011011000",
  27960=>"000111111",
  27961=>"101011000",
  27962=>"010001110",
  27963=>"100111000",
  27964=>"111101000",
  27965=>"110011001",
  27966=>"001011010",
  27967=>"011110000",
  27968=>"010111111",
  27969=>"001000101",
  27970=>"011010110",
  27971=>"110100011",
  27972=>"000111111",
  27973=>"110110000",
  27974=>"111111001",
  27975=>"111010111",
  27976=>"111110000",
  27977=>"010011100",
  27978=>"011000110",
  27979=>"000101101",
  27980=>"001001100",
  27981=>"101011011",
  27982=>"000100010",
  27983=>"011111100",
  27984=>"001111110",
  27985=>"010110000",
  27986=>"000111001",
  27987=>"001001111",
  27988=>"111000010",
  27989=>"000000111",
  27990=>"000101011",
  27991=>"001000111",
  27992=>"001110110",
  27993=>"000001011",
  27994=>"011101100",
  27995=>"110000011",
  27996=>"111011011",
  27997=>"111110010",
  27998=>"011000001",
  27999=>"010001000",
  28000=>"110100100",
  28001=>"011011101",
  28002=>"001110011",
  28003=>"000000101",
  28004=>"010011001",
  28005=>"101010000",
  28006=>"110111000",
  28007=>"001000000",
  28008=>"000101000",
  28009=>"011111100",
  28010=>"101111011",
  28011=>"000000010",
  28012=>"101011110",
  28013=>"010100000",
  28014=>"100110101",
  28015=>"001100101",
  28016=>"101110111",
  28017=>"011111100",
  28018=>"001010100",
  28019=>"100101011",
  28020=>"110001110",
  28021=>"010101101",
  28022=>"100101010",
  28023=>"011000011",
  28024=>"100010110",
  28025=>"101111111",
  28026=>"000111110",
  28027=>"011110001",
  28028=>"011010100",
  28029=>"011010111",
  28030=>"001101010",
  28031=>"011001100",
  28032=>"010001011",
  28033=>"000010100",
  28034=>"111010111",
  28035=>"011010000",
  28036=>"001100111",
  28037=>"110101101",
  28038=>"010000001",
  28039=>"011111110",
  28040=>"100101011",
  28041=>"111011111",
  28042=>"100111010",
  28043=>"111111000",
  28044=>"111100010",
  28045=>"001001011",
  28046=>"101011100",
  28047=>"111101010",
  28048=>"000010111",
  28049=>"001001100",
  28050=>"011110000",
  28051=>"000010110",
  28052=>"010000101",
  28053=>"000101010",
  28054=>"100001101",
  28055=>"010000000",
  28056=>"100110100",
  28057=>"111110101",
  28058=>"111001110",
  28059=>"100001110",
  28060=>"001110100",
  28061=>"100111010",
  28062=>"101101001",
  28063=>"010000111",
  28064=>"111101110",
  28065=>"101100001",
  28066=>"000000110",
  28067=>"010101101",
  28068=>"100011110",
  28069=>"100100111",
  28070=>"101001100",
  28071=>"100111100",
  28072=>"011011000",
  28073=>"010100001",
  28074=>"000000010",
  28075=>"000010101",
  28076=>"111011111",
  28077=>"001011110",
  28078=>"100001101",
  28079=>"101100000",
  28080=>"010011010",
  28081=>"001100100",
  28082=>"111010001",
  28083=>"101001110",
  28084=>"000011011",
  28085=>"000010101",
  28086=>"001110001",
  28087=>"100111010",
  28088=>"110111100",
  28089=>"000111111",
  28090=>"101110011",
  28091=>"010100100",
  28092=>"001000101",
  28093=>"101101100",
  28094=>"100101000",
  28095=>"111101011",
  28096=>"101010011",
  28097=>"111111100",
  28098=>"000000110",
  28099=>"010000110",
  28100=>"011110000",
  28101=>"000010110",
  28102=>"000011010",
  28103=>"011001111",
  28104=>"010110000",
  28105=>"010000110",
  28106=>"000110110",
  28107=>"110111001",
  28108=>"100010010",
  28109=>"111010001",
  28110=>"111000001",
  28111=>"000101100",
  28112=>"001011010",
  28113=>"100111110",
  28114=>"000101001",
  28115=>"111110101",
  28116=>"101010111",
  28117=>"101100000",
  28118=>"110110100",
  28119=>"110101010",
  28120=>"011010011",
  28121=>"010011111",
  28122=>"100111000",
  28123=>"010001111",
  28124=>"010100111",
  28125=>"100100110",
  28126=>"011100011",
  28127=>"000110110",
  28128=>"011110000",
  28129=>"010101001",
  28130=>"110001100",
  28131=>"101000000",
  28132=>"000110111",
  28133=>"110010001",
  28134=>"111010110",
  28135=>"010000110",
  28136=>"011001000",
  28137=>"001001001",
  28138=>"100110011",
  28139=>"100111100",
  28140=>"100010110",
  28141=>"101010010",
  28142=>"111101000",
  28143=>"001011110",
  28144=>"111011011",
  28145=>"001111111",
  28146=>"010110000",
  28147=>"110010101",
  28148=>"000110100",
  28149=>"010011010",
  28150=>"111111110",
  28151=>"011110010",
  28152=>"100010011",
  28153=>"100000011",
  28154=>"111010000",
  28155=>"111101110",
  28156=>"100101011",
  28157=>"111000111",
  28158=>"000011000",
  28159=>"101001000",
  28160=>"111100001",
  28161=>"001000111",
  28162=>"010011010",
  28163=>"010010000",
  28164=>"001011010",
  28165=>"000110011",
  28166=>"111110000",
  28167=>"001110011",
  28168=>"000001101",
  28169=>"010001001",
  28170=>"000010100",
  28171=>"000100011",
  28172=>"011000011",
  28173=>"001000010",
  28174=>"000000111",
  28175=>"001100010",
  28176=>"001000001",
  28177=>"100100010",
  28178=>"111011000",
  28179=>"010000010",
  28180=>"001010010",
  28181=>"111010111",
  28182=>"110001000",
  28183=>"010100001",
  28184=>"101111110",
  28185=>"111101110",
  28186=>"101001001",
  28187=>"010000110",
  28188=>"110101111",
  28189=>"010111010",
  28190=>"111101111",
  28191=>"100011100",
  28192=>"011101010",
  28193=>"100010111",
  28194=>"000110000",
  28195=>"001000001",
  28196=>"100110110",
  28197=>"010110110",
  28198=>"010010100",
  28199=>"100011000",
  28200=>"101000001",
  28201=>"000110110",
  28202=>"000100010",
  28203=>"111011010",
  28204=>"011001100",
  28205=>"110101010",
  28206=>"011011100",
  28207=>"000000010",
  28208=>"111000000",
  28209=>"110010010",
  28210=>"000010101",
  28211=>"011000001",
  28212=>"111010111",
  28213=>"001000011",
  28214=>"000101111",
  28215=>"110111000",
  28216=>"010010100",
  28217=>"101100000",
  28218=>"110010001",
  28219=>"000010100",
  28220=>"110010011",
  28221=>"001100111",
  28222=>"110101100",
  28223=>"001000001",
  28224=>"000101001",
  28225=>"110010110",
  28226=>"011110010",
  28227=>"101111100",
  28228=>"110110001",
  28229=>"011000001",
  28230=>"001001100",
  28231=>"000010111",
  28232=>"110110100",
  28233=>"100111000",
  28234=>"111100110",
  28235=>"111111111",
  28236=>"111000001",
  28237=>"101101001",
  28238=>"100100110",
  28239=>"011100000",
  28240=>"010000011",
  28241=>"000000000",
  28242=>"111111001",
  28243=>"100010000",
  28244=>"101010100",
  28245=>"111111111",
  28246=>"010010010",
  28247=>"101110000",
  28248=>"110011111",
  28249=>"000010001",
  28250=>"011101011",
  28251=>"111101100",
  28252=>"101110000",
  28253=>"011010101",
  28254=>"111101011",
  28255=>"111000101",
  28256=>"100011111",
  28257=>"010100110",
  28258=>"100011011",
  28259=>"111010011",
  28260=>"011010101",
  28261=>"101011001",
  28262=>"111101100",
  28263=>"110000001",
  28264=>"100100000",
  28265=>"011000110",
  28266=>"111101001",
  28267=>"000001011",
  28268=>"100101000",
  28269=>"100011110",
  28270=>"100001000",
  28271=>"111101100",
  28272=>"101110100",
  28273=>"001110011",
  28274=>"100101110",
  28275=>"101000111",
  28276=>"110100110",
  28277=>"111010110",
  28278=>"011110110",
  28279=>"100111100",
  28280=>"100100011",
  28281=>"101110001",
  28282=>"100010011",
  28283=>"010000011",
  28284=>"000010000",
  28285=>"110111000",
  28286=>"011111100",
  28287=>"010001010",
  28288=>"111011000",
  28289=>"111010100",
  28290=>"100110011",
  28291=>"101001001",
  28292=>"101111000",
  28293=>"111000001",
  28294=>"001111100",
  28295=>"101111111",
  28296=>"001000000",
  28297=>"010001011",
  28298=>"101011001",
  28299=>"010111000",
  28300=>"110111101",
  28301=>"000101001",
  28302=>"010011111",
  28303=>"010001101",
  28304=>"110110111",
  28305=>"010100100",
  28306=>"110101011",
  28307=>"111110110",
  28308=>"101001000",
  28309=>"110100100",
  28310=>"111100110",
  28311=>"011001111",
  28312=>"010011101",
  28313=>"110000100",
  28314=>"110010111",
  28315=>"110000010",
  28316=>"100100110",
  28317=>"001000100",
  28318=>"010110101",
  28319=>"001000000",
  28320=>"111110000",
  28321=>"100100011",
  28322=>"111010001",
  28323=>"011100100",
  28324=>"110000000",
  28325=>"110010111",
  28326=>"110011000",
  28327=>"101111010",
  28328=>"111100111",
  28329=>"101101010",
  28330=>"100000100",
  28331=>"000000111",
  28332=>"011011111",
  28333=>"111100001",
  28334=>"111011110",
  28335=>"010111011",
  28336=>"110110001",
  28337=>"110011011",
  28338=>"010011010",
  28339=>"010110011",
  28340=>"001111001",
  28341=>"100000011",
  28342=>"110000101",
  28343=>"100000000",
  28344=>"100101000",
  28345=>"011011001",
  28346=>"011010011",
  28347=>"101110011",
  28348=>"011001101",
  28349=>"100010010",
  28350=>"101100101",
  28351=>"110010000",
  28352=>"010000001",
  28353=>"001011010",
  28354=>"101000010",
  28355=>"111011100",
  28356=>"100111000",
  28357=>"100110000",
  28358=>"010100000",
  28359=>"100110110",
  28360=>"010100000",
  28361=>"111000110",
  28362=>"011011001",
  28363=>"100110001",
  28364=>"001001110",
  28365=>"011011110",
  28366=>"101011110",
  28367=>"100011000",
  28368=>"000001100",
  28369=>"011101011",
  28370=>"000111101",
  28371=>"101111010",
  28372=>"111100011",
  28373=>"000111111",
  28374=>"111000001",
  28375=>"000010000",
  28376=>"110111110",
  28377=>"011001010",
  28378=>"010010011",
  28379=>"110111101",
  28380=>"000001101",
  28381=>"100111111",
  28382=>"010100011",
  28383=>"101011111",
  28384=>"010001111",
  28385=>"011110110",
  28386=>"110111011",
  28387=>"110100000",
  28388=>"110100111",
  28389=>"101101100",
  28390=>"000001111",
  28391=>"111011101",
  28392=>"111100001",
  28393=>"101110100",
  28394=>"010001011",
  28395=>"100110100",
  28396=>"011100101",
  28397=>"000111110",
  28398=>"110010100",
  28399=>"101100101",
  28400=>"010010001",
  28401=>"010000011",
  28402=>"111111000",
  28403=>"100100110",
  28404=>"100101110",
  28405=>"100110011",
  28406=>"011010101",
  28407=>"011011000",
  28408=>"011011111",
  28409=>"101001000",
  28410=>"100000011",
  28411=>"001001111",
  28412=>"101001110",
  28413=>"011101010",
  28414=>"011000000",
  28415=>"001100100",
  28416=>"011000001",
  28417=>"110010000",
  28418=>"011010010",
  28419=>"000110001",
  28420=>"101000110",
  28421=>"101000111",
  28422=>"101110001",
  28423=>"010110101",
  28424=>"110111010",
  28425=>"110000001",
  28426=>"000111001",
  28427=>"111011010",
  28428=>"110001010",
  28429=>"011011111",
  28430=>"010101101",
  28431=>"010010000",
  28432=>"000011011",
  28433=>"101011000",
  28434=>"001100110",
  28435=>"101001000",
  28436=>"010000011",
  28437=>"110110001",
  28438=>"001111000",
  28439=>"111001000",
  28440=>"101100101",
  28441=>"110110000",
  28442=>"010111011",
  28443=>"011011000",
  28444=>"010010010",
  28445=>"001100100",
  28446=>"110100010",
  28447=>"010011111",
  28448=>"100110101",
  28449=>"001011111",
  28450=>"010101001",
  28451=>"101011110",
  28452=>"011111101",
  28453=>"010000000",
  28454=>"001011111",
  28455=>"101000000",
  28456=>"110101011",
  28457=>"101000011",
  28458=>"011000110",
  28459=>"011000001",
  28460=>"011001000",
  28461=>"011010111",
  28462=>"110011101",
  28463=>"111010111",
  28464=>"101000001",
  28465=>"101010000",
  28466=>"000001010",
  28467=>"110100101",
  28468=>"111110001",
  28469=>"100100100",
  28470=>"011100101",
  28471=>"001100010",
  28472=>"100110101",
  28473=>"100011100",
  28474=>"000101100",
  28475=>"010000000",
  28476=>"111111100",
  28477=>"000111111",
  28478=>"101101010",
  28479=>"100110010",
  28480=>"011001111",
  28481=>"000001010",
  28482=>"101011101",
  28483=>"101100010",
  28484=>"111011000",
  28485=>"101100111",
  28486=>"101010011",
  28487=>"010010101",
  28488=>"101100101",
  28489=>"100110000",
  28490=>"000101110",
  28491=>"100100000",
  28492=>"111011000",
  28493=>"111111110",
  28494=>"011100110",
  28495=>"111110100",
  28496=>"101111010",
  28497=>"011010111",
  28498=>"110000111",
  28499=>"110010110",
  28500=>"011010100",
  28501=>"011110011",
  28502=>"000001101",
  28503=>"001001111",
  28504=>"100010110",
  28505=>"001100010",
  28506=>"001000101",
  28507=>"101000100",
  28508=>"000010000",
  28509=>"011111101",
  28510=>"100000010",
  28511=>"100101010",
  28512=>"001010010",
  28513=>"100100100",
  28514=>"001000010",
  28515=>"101100110",
  28516=>"111010100",
  28517=>"011010000",
  28518=>"000100101",
  28519=>"111110111",
  28520=>"101101111",
  28521=>"111000010",
  28522=>"100010101",
  28523=>"000001000",
  28524=>"111011011",
  28525=>"101111000",
  28526=>"011101010",
  28527=>"110101100",
  28528=>"010010110",
  28529=>"010110000",
  28530=>"011010001",
  28531=>"000111110",
  28532=>"110101010",
  28533=>"000111010",
  28534=>"100111101",
  28535=>"001010001",
  28536=>"111111110",
  28537=>"001101101",
  28538=>"010000011",
  28539=>"001010101",
  28540=>"010111000",
  28541=>"110110101",
  28542=>"000001011",
  28543=>"101011101",
  28544=>"111011011",
  28545=>"011111010",
  28546=>"001111011",
  28547=>"001101101",
  28548=>"100011110",
  28549=>"011011001",
  28550=>"000110010",
  28551=>"011100001",
  28552=>"010000000",
  28553=>"101111100",
  28554=>"000101000",
  28555=>"000000010",
  28556=>"101100110",
  28557=>"011101001",
  28558=>"010011000",
  28559=>"100100001",
  28560=>"110101001",
  28561=>"000001000",
  28562=>"101000111",
  28563=>"000110110",
  28564=>"000010110",
  28565=>"000110000",
  28566=>"010100110",
  28567=>"101010001",
  28568=>"001110101",
  28569=>"100100110",
  28570=>"111100110",
  28571=>"101101001",
  28572=>"011011101",
  28573=>"110111110",
  28574=>"100100111",
  28575=>"011101110",
  28576=>"101001101",
  28577=>"111111100",
  28578=>"111101101",
  28579=>"000110010",
  28580=>"000101000",
  28581=>"001011000",
  28582=>"111111111",
  28583=>"110110011",
  28584=>"101001110",
  28585=>"101101000",
  28586=>"011111100",
  28587=>"000100111",
  28588=>"111101101",
  28589=>"000111000",
  28590=>"111010111",
  28591=>"111000101",
  28592=>"111010001",
  28593=>"011101111",
  28594=>"000111110",
  28595=>"010101111",
  28596=>"100011000",
  28597=>"011101010",
  28598=>"110110011",
  28599=>"101011111",
  28600=>"001000011",
  28601=>"111010110",
  28602=>"111010101",
  28603=>"110011001",
  28604=>"101101001",
  28605=>"111010110",
  28606=>"110101111",
  28607=>"110111101",
  28608=>"001001100",
  28609=>"010010111",
  28610=>"000010011",
  28611=>"000000010",
  28612=>"100000010",
  28613=>"001111011",
  28614=>"011110110",
  28615=>"010111011",
  28616=>"010111110",
  28617=>"011011110",
  28618=>"101000000",
  28619=>"110011111",
  28620=>"010100110",
  28621=>"001001000",
  28622=>"001000010",
  28623=>"111011101",
  28624=>"100110100",
  28625=>"011110111",
  28626=>"010001101",
  28627=>"001000000",
  28628=>"111100101",
  28629=>"111000101",
  28630=>"101111011",
  28631=>"101011011",
  28632=>"010000000",
  28633=>"110000111",
  28634=>"111111100",
  28635=>"100111111",
  28636=>"100111010",
  28637=>"111011111",
  28638=>"001100111",
  28639=>"001011111",
  28640=>"100110000",
  28641=>"001111111",
  28642=>"000010100",
  28643=>"100010110",
  28644=>"000101100",
  28645=>"111110100",
  28646=>"110110110",
  28647=>"111101010",
  28648=>"110110101",
  28649=>"111111010",
  28650=>"100010110",
  28651=>"100100000",
  28652=>"011010011",
  28653=>"100011100",
  28654=>"001111010",
  28655=>"101100000",
  28656=>"001001111",
  28657=>"111001011",
  28658=>"111011110",
  28659=>"110001100",
  28660=>"010011001",
  28661=>"101100101",
  28662=>"011010111",
  28663=>"000110001",
  28664=>"101000111",
  28665=>"001010111",
  28666=>"010101001",
  28667=>"001000010",
  28668=>"110100000",
  28669=>"000101000",
  28670=>"001001001",
  28671=>"001010000",
  28672=>"001011000",
  28673=>"010000001",
  28674=>"101000010",
  28675=>"100001010",
  28676=>"111011000",
  28677=>"100001010",
  28678=>"101110001",
  28679=>"101011000",
  28680=>"101000100",
  28681=>"010001010",
  28682=>"010010010",
  28683=>"011111011",
  28684=>"000101111",
  28685=>"011111011",
  28686=>"110010101",
  28687=>"111000011",
  28688=>"110100001",
  28689=>"001001100",
  28690=>"110110110",
  28691=>"001001110",
  28692=>"100111001",
  28693=>"101000000",
  28694=>"000000001",
  28695=>"010000101",
  28696=>"010011011",
  28697=>"010000111",
  28698=>"010110001",
  28699=>"110010111",
  28700=>"010100010",
  28701=>"000111000",
  28702=>"011000110",
  28703=>"101001001",
  28704=>"000101100",
  28705=>"110101111",
  28706=>"000010111",
  28707=>"001010111",
  28708=>"000100000",
  28709=>"011011010",
  28710=>"100011010",
  28711=>"001110010",
  28712=>"010111001",
  28713=>"110001101",
  28714=>"011110011",
  28715=>"100000100",
  28716=>"100001001",
  28717=>"010011110",
  28718=>"100110101",
  28719=>"101111001",
  28720=>"100111111",
  28721=>"110010010",
  28722=>"010111001",
  28723=>"011000000",
  28724=>"001110011",
  28725=>"110000010",
  28726=>"111010011",
  28727=>"001110001",
  28728=>"011100101",
  28729=>"001000110",
  28730=>"110000001",
  28731=>"111100011",
  28732=>"100100101",
  28733=>"100110110",
  28734=>"001010101",
  28735=>"100001100",
  28736=>"111101001",
  28737=>"000010110",
  28738=>"000001000",
  28739=>"000111110",
  28740=>"001010110",
  28741=>"111000000",
  28742=>"011001111",
  28743=>"011110010",
  28744=>"000001010",
  28745=>"000110100",
  28746=>"110001000",
  28747=>"010111100",
  28748=>"001111111",
  28749=>"101010011",
  28750=>"111000110",
  28751=>"000010000",
  28752=>"001100000",
  28753=>"100000110",
  28754=>"010001111",
  28755=>"010100010",
  28756=>"000011110",
  28757=>"011110110",
  28758=>"110010000",
  28759=>"010110001",
  28760=>"001000001",
  28761=>"111010010",
  28762=>"011100100",
  28763=>"001101010",
  28764=>"010000110",
  28765=>"110001100",
  28766=>"000100011",
  28767=>"000110111",
  28768=>"010110011",
  28769=>"001011001",
  28770=>"111100111",
  28771=>"011111111",
  28772=>"011110001",
  28773=>"111100110",
  28774=>"111111010",
  28775=>"100110111",
  28776=>"000011001",
  28777=>"011101111",
  28778=>"000101011",
  28779=>"011000001",
  28780=>"100011001",
  28781=>"111011011",
  28782=>"011010011",
  28783=>"000111100",
  28784=>"111000010",
  28785=>"001101111",
  28786=>"001101110",
  28787=>"011100011",
  28788=>"000000000",
  28789=>"000101011",
  28790=>"100001110",
  28791=>"010100111",
  28792=>"000000101",
  28793=>"011101010",
  28794=>"010010010",
  28795=>"000000011",
  28796=>"110001100",
  28797=>"001101000",
  28798=>"010000100",
  28799=>"111011011",
  28800=>"110100101",
  28801=>"010100000",
  28802=>"111101111",
  28803=>"100110101",
  28804=>"000010110",
  28805=>"110000011",
  28806=>"111010110",
  28807=>"000111011",
  28808=>"010100000",
  28809=>"101001011",
  28810=>"000000101",
  28811=>"111101101",
  28812=>"111000010",
  28813=>"100100011",
  28814=>"010010100",
  28815=>"001010011",
  28816=>"000110101",
  28817=>"011010011",
  28818=>"110100001",
  28819=>"111011111",
  28820=>"000010100",
  28821=>"011011010",
  28822=>"001010001",
  28823=>"001010110",
  28824=>"110100100",
  28825=>"001111001",
  28826=>"101101000",
  28827=>"010111000",
  28828=>"010001001",
  28829=>"111000100",
  28830=>"001001010",
  28831=>"101111111",
  28832=>"100011101",
  28833=>"110101111",
  28834=>"001100001",
  28835=>"101101111",
  28836=>"101010011",
  28837=>"000010111",
  28838=>"010110000",
  28839=>"000110010",
  28840=>"101001000",
  28841=>"101101000",
  28842=>"111111010",
  28843=>"100110101",
  28844=>"010111011",
  28845=>"010101001",
  28846=>"111001010",
  28847=>"111100110",
  28848=>"001001010",
  28849=>"001010100",
  28850=>"011101001",
  28851=>"000000010",
  28852=>"010000101",
  28853=>"111110100",
  28854=>"001001000",
  28855=>"011011011",
  28856=>"010011011",
  28857=>"001101100",
  28858=>"010101100",
  28859=>"000010011",
  28860=>"000110100",
  28861=>"101111001",
  28862=>"101010001",
  28863=>"001011110",
  28864=>"111001101",
  28865=>"000110110",
  28866=>"000110011",
  28867=>"011110111",
  28868=>"111110110",
  28869=>"010110000",
  28870=>"001111111",
  28871=>"000111111",
  28872=>"111001010",
  28873=>"101100101",
  28874=>"011111111",
  28875=>"101100000",
  28876=>"011001010",
  28877=>"000001100",
  28878=>"110010101",
  28879=>"010011001",
  28880=>"000000001",
  28881=>"010101111",
  28882=>"000000100",
  28883=>"000100011",
  28884=>"110011100",
  28885=>"000011111",
  28886=>"100101010",
  28887=>"100110100",
  28888=>"111101000",
  28889=>"100000110",
  28890=>"100010010",
  28891=>"100010010",
  28892=>"110011010",
  28893=>"111001011",
  28894=>"000000100",
  28895=>"001000100",
  28896=>"010101001",
  28897=>"010101001",
  28898=>"100100011",
  28899=>"101111110",
  28900=>"111000111",
  28901=>"101110100",
  28902=>"110001000",
  28903=>"000010100",
  28904=>"000000011",
  28905=>"000101110",
  28906=>"000001000",
  28907=>"001111110",
  28908=>"111110000",
  28909=>"001011110",
  28910=>"011001010",
  28911=>"001011000",
  28912=>"001100111",
  28913=>"101111011",
  28914=>"011001001",
  28915=>"000010001",
  28916=>"100011101",
  28917=>"111111001",
  28918=>"110111000",
  28919=>"010000000",
  28920=>"001010100",
  28921=>"001101010",
  28922=>"111000100",
  28923=>"100101001",
  28924=>"111000100",
  28925=>"000111000",
  28926=>"011011101",
  28927=>"011111101",
  28928=>"111000011",
  28929=>"110010101",
  28930=>"010000000",
  28931=>"000110100",
  28932=>"100101001",
  28933=>"001011000",
  28934=>"111110100",
  28935=>"101001001",
  28936=>"000110111",
  28937=>"101000000",
  28938=>"001100000",
  28939=>"011111111",
  28940=>"010100111",
  28941=>"000000001",
  28942=>"000101001",
  28943=>"001101010",
  28944=>"011000010",
  28945=>"110001110",
  28946=>"000010001",
  28947=>"000010001",
  28948=>"000110010",
  28949=>"100001110",
  28950=>"111010100",
  28951=>"000111000",
  28952=>"000101101",
  28953=>"000100110",
  28954=>"000001100",
  28955=>"100101101",
  28956=>"000011010",
  28957=>"000000101",
  28958=>"000110101",
  28959=>"010100000",
  28960=>"110000010",
  28961=>"101111100",
  28962=>"100110111",
  28963=>"110111111",
  28964=>"101011101",
  28965=>"111110010",
  28966=>"111011000",
  28967=>"010011111",
  28968=>"111001000",
  28969=>"111111111",
  28970=>"000111000",
  28971=>"110011100",
  28972=>"000000110",
  28973=>"111111101",
  28974=>"001011101",
  28975=>"001110111",
  28976=>"110001110",
  28977=>"101000000",
  28978=>"010100110",
  28979=>"001100011",
  28980=>"110001001",
  28981=>"000011010",
  28982=>"111110111",
  28983=>"010010101",
  28984=>"001110000",
  28985=>"111101101",
  28986=>"010100000",
  28987=>"111010011",
  28988=>"111101111",
  28989=>"000100000",
  28990=>"111101110",
  28991=>"101111110",
  28992=>"001011010",
  28993=>"010101001",
  28994=>"111111111",
  28995=>"001000100",
  28996=>"000011100",
  28997=>"010010100",
  28998=>"010111101",
  28999=>"110001001",
  29000=>"000010111",
  29001=>"000001111",
  29002=>"001001101",
  29003=>"000011100",
  29004=>"111010100",
  29005=>"110001001",
  29006=>"110001100",
  29007=>"011000010",
  29008=>"100011010",
  29009=>"001100011",
  29010=>"101011101",
  29011=>"100000000",
  29012=>"000010110",
  29013=>"111010011",
  29014=>"111110010",
  29015=>"111111110",
  29016=>"100000011",
  29017=>"101000011",
  29018=>"110111111",
  29019=>"111110111",
  29020=>"101101001",
  29021=>"011111110",
  29022=>"110001010",
  29023=>"010110001",
  29024=>"000011101",
  29025=>"111100110",
  29026=>"111100001",
  29027=>"001010011",
  29028=>"010110101",
  29029=>"010100000",
  29030=>"000011001",
  29031=>"111010011",
  29032=>"100011110",
  29033=>"110000011",
  29034=>"010001101",
  29035=>"010101110",
  29036=>"100001100",
  29037=>"001011010",
  29038=>"100000100",
  29039=>"000001011",
  29040=>"100010011",
  29041=>"111110000",
  29042=>"010000001",
  29043=>"100100111",
  29044=>"010110101",
  29045=>"011001000",
  29046=>"101100011",
  29047=>"010111010",
  29048=>"001010011",
  29049=>"001110010",
  29050=>"110011111",
  29051=>"100001101",
  29052=>"001111001",
  29053=>"110101111",
  29054=>"100111000",
  29055=>"111100000",
  29056=>"100101100",
  29057=>"101011101",
  29058=>"001101000",
  29059=>"101000110",
  29060=>"000100010",
  29061=>"001110101",
  29062=>"111011010",
  29063=>"000101001",
  29064=>"000001000",
  29065=>"001101100",
  29066=>"000100111",
  29067=>"010001110",
  29068=>"010101111",
  29069=>"010001011",
  29070=>"111000110",
  29071=>"000000100",
  29072=>"010001001",
  29073=>"111111001",
  29074=>"101101010",
  29075=>"000011000",
  29076=>"000101101",
  29077=>"000011111",
  29078=>"111111111",
  29079=>"110111010",
  29080=>"100110001",
  29081=>"001000110",
  29082=>"010100011",
  29083=>"011010011",
  29084=>"111101001",
  29085=>"101111011",
  29086=>"010010100",
  29087=>"011111111",
  29088=>"110100011",
  29089=>"101001010",
  29090=>"100010111",
  29091=>"000101000",
  29092=>"100110101",
  29093=>"011000011",
  29094=>"001011110",
  29095=>"010101111",
  29096=>"011010101",
  29097=>"111111001",
  29098=>"110011001",
  29099=>"101110110",
  29100=>"101100010",
  29101=>"111010001",
  29102=>"000000100",
  29103=>"011100000",
  29104=>"101011101",
  29105=>"000011001",
  29106=>"000001000",
  29107=>"110010000",
  29108=>"101100100",
  29109=>"111011010",
  29110=>"010101100",
  29111=>"011001001",
  29112=>"010001100",
  29113=>"001101011",
  29114=>"000001011",
  29115=>"111101110",
  29116=>"111100110",
  29117=>"100001000",
  29118=>"001001001",
  29119=>"001110000",
  29120=>"110000000",
  29121=>"001000011",
  29122=>"100100001",
  29123=>"110100000",
  29124=>"000010010",
  29125=>"101010011",
  29126=>"101010110",
  29127=>"111001010",
  29128=>"000000000",
  29129=>"100010100",
  29130=>"000101101",
  29131=>"111111010",
  29132=>"100010000",
  29133=>"000001001",
  29134=>"000011111",
  29135=>"100001000",
  29136=>"111111000",
  29137=>"111111111",
  29138=>"111001111",
  29139=>"010111001",
  29140=>"011110000",
  29141=>"100111010",
  29142=>"010111101",
  29143=>"001011001",
  29144=>"101101001",
  29145=>"100001001",
  29146=>"001111100",
  29147=>"101110111",
  29148=>"111010101",
  29149=>"111001100",
  29150=>"111001101",
  29151=>"001111111",
  29152=>"101001001",
  29153=>"011101000",
  29154=>"111111000",
  29155=>"000111101",
  29156=>"011011000",
  29157=>"001000011",
  29158=>"100011000",
  29159=>"111100000",
  29160=>"011110010",
  29161=>"000101000",
  29162=>"110010100",
  29163=>"111001000",
  29164=>"010011100",
  29165=>"010001000",
  29166=>"010101010",
  29167=>"011101010",
  29168=>"011000000",
  29169=>"011001100",
  29170=>"011011011",
  29171=>"110100100",
  29172=>"111010110",
  29173=>"001010000",
  29174=>"011001001",
  29175=>"111000100",
  29176=>"000000000",
  29177=>"001001001",
  29178=>"111011110",
  29179=>"001001011",
  29180=>"010101101",
  29181=>"010100111",
  29182=>"100111100",
  29183=>"011011101",
  29184=>"010010010",
  29185=>"110001101",
  29186=>"011000011",
  29187=>"001101000",
  29188=>"000001000",
  29189=>"010000101",
  29190=>"110111011",
  29191=>"110000100",
  29192=>"010101001",
  29193=>"100011101",
  29194=>"010010110",
  29195=>"101000011",
  29196=>"000010000",
  29197=>"001100001",
  29198=>"001100000",
  29199=>"100110010",
  29200=>"111101100",
  29201=>"101111101",
  29202=>"110111100",
  29203=>"011111011",
  29204=>"100000110",
  29205=>"100100110",
  29206=>"100111011",
  29207=>"011011011",
  29208=>"110111000",
  29209=>"101110001",
  29210=>"010110110",
  29211=>"000010111",
  29212=>"110010011",
  29213=>"001100001",
  29214=>"101011111",
  29215=>"000110001",
  29216=>"000001001",
  29217=>"111010000",
  29218=>"010110010",
  29219=>"000101010",
  29220=>"101111111",
  29221=>"110000000",
  29222=>"110010101",
  29223=>"010101111",
  29224=>"001101001",
  29225=>"110001001",
  29226=>"001000001",
  29227=>"001010100",
  29228=>"111111111",
  29229=>"110000000",
  29230=>"111101000",
  29231=>"101011011",
  29232=>"100110001",
  29233=>"101111001",
  29234=>"111001011",
  29235=>"010010110",
  29236=>"010100000",
  29237=>"001001010",
  29238=>"010110101",
  29239=>"100111000",
  29240=>"010100011",
  29241=>"110010011",
  29242=>"001001000",
  29243=>"001011000",
  29244=>"001101111",
  29245=>"110101001",
  29246=>"010011000",
  29247=>"010111100",
  29248=>"001101011",
  29249=>"101101010",
  29250=>"100100011",
  29251=>"000100101",
  29252=>"011111111",
  29253=>"011101000",
  29254=>"010000101",
  29255=>"010011010",
  29256=>"011001111",
  29257=>"110110110",
  29258=>"001110010",
  29259=>"111010010",
  29260=>"100000101",
  29261=>"111000111",
  29262=>"100010000",
  29263=>"100001110",
  29264=>"110110010",
  29265=>"111001000",
  29266=>"010000001",
  29267=>"010111111",
  29268=>"011001110",
  29269=>"001010110",
  29270=>"010100011",
  29271=>"110110000",
  29272=>"001000110",
  29273=>"011011010",
  29274=>"111001100",
  29275=>"111011110",
  29276=>"110111110",
  29277=>"001011000",
  29278=>"000011111",
  29279=>"110010001",
  29280=>"110001000",
  29281=>"111001001",
  29282=>"100011001",
  29283=>"000100000",
  29284=>"000100000",
  29285=>"110111011",
  29286=>"010111011",
  29287=>"000101000",
  29288=>"111100110",
  29289=>"110010111",
  29290=>"011001010",
  29291=>"110101110",
  29292=>"011101101",
  29293=>"111111001",
  29294=>"000000000",
  29295=>"010011101",
  29296=>"101101001",
  29297=>"111110010",
  29298=>"010111111",
  29299=>"110011010",
  29300=>"100001011",
  29301=>"010000100",
  29302=>"110100110",
  29303=>"111111100",
  29304=>"001001110",
  29305=>"010110000",
  29306=>"000111001",
  29307=>"101101100",
  29308=>"100110101",
  29309=>"100010011",
  29310=>"000010101",
  29311=>"100000101",
  29312=>"101111101",
  29313=>"110100001",
  29314=>"010110111",
  29315=>"000100110",
  29316=>"111110100",
  29317=>"101111010",
  29318=>"100111111",
  29319=>"111101111",
  29320=>"000111010",
  29321=>"001110101",
  29322=>"110111011",
  29323=>"111100011",
  29324=>"111011101",
  29325=>"101011100",
  29326=>"010110100",
  29327=>"100100001",
  29328=>"101111000",
  29329=>"011100100",
  29330=>"111010111",
  29331=>"100110000",
  29332=>"010110001",
  29333=>"001101111",
  29334=>"000000011",
  29335=>"100101111",
  29336=>"010111011",
  29337=>"100010000",
  29338=>"110100110",
  29339=>"110111111",
  29340=>"010111001",
  29341=>"011100001",
  29342=>"000110110",
  29343=>"000010000",
  29344=>"111101011",
  29345=>"100000100",
  29346=>"111100101",
  29347=>"110001101",
  29348=>"001011000",
  29349=>"101010111",
  29350=>"000101110",
  29351=>"100011011",
  29352=>"101011111",
  29353=>"011110110",
  29354=>"010001110",
  29355=>"010110100",
  29356=>"010110101",
  29357=>"101010000",
  29358=>"000001100",
  29359=>"011010010",
  29360=>"111000001",
  29361=>"011101110",
  29362=>"110011001",
  29363=>"110101110",
  29364=>"101010000",
  29365=>"010101110",
  29366=>"110001000",
  29367=>"000010101",
  29368=>"010011110",
  29369=>"001101110",
  29370=>"111101101",
  29371=>"110111101",
  29372=>"110101111",
  29373=>"001011011",
  29374=>"011101101",
  29375=>"110000000",
  29376=>"101100010",
  29377=>"011110111",
  29378=>"111101100",
  29379=>"010011000",
  29380=>"010001001",
  29381=>"101010101",
  29382=>"100101011",
  29383=>"110101110",
  29384=>"110100100",
  29385=>"011111000",
  29386=>"001100111",
  29387=>"010110010",
  29388=>"111111010",
  29389=>"000011101",
  29390=>"001111111",
  29391=>"010001100",
  29392=>"001101001",
  29393=>"101101101",
  29394=>"000010011",
  29395=>"011000110",
  29396=>"100000011",
  29397=>"000011010",
  29398=>"100111011",
  29399=>"011011011",
  29400=>"001010110",
  29401=>"101000011",
  29402=>"011000101",
  29403=>"101110001",
  29404=>"101101111",
  29405=>"000100101",
  29406=>"101100111",
  29407=>"100110010",
  29408=>"111100100",
  29409=>"111010110",
  29410=>"101100010",
  29411=>"111110101",
  29412=>"100010101",
  29413=>"111111110",
  29414=>"000010001",
  29415=>"000010010",
  29416=>"010000100",
  29417=>"000100101",
  29418=>"010110010",
  29419=>"001001000",
  29420=>"101110111",
  29421=>"101110100",
  29422=>"000010001",
  29423=>"100000001",
  29424=>"010111110",
  29425=>"011010110",
  29426=>"100101100",
  29427=>"100000100",
  29428=>"111000010",
  29429=>"010000100",
  29430=>"110111100",
  29431=>"000101101",
  29432=>"110101110",
  29433=>"110100001",
  29434=>"110100000",
  29435=>"101010000",
  29436=>"011001101",
  29437=>"101101101",
  29438=>"100011110",
  29439=>"000001010",
  29440=>"100110000",
  29441=>"110110110",
  29442=>"010010101",
  29443=>"000100111",
  29444=>"011110000",
  29445=>"100110000",
  29446=>"000011110",
  29447=>"010100010",
  29448=>"111111011",
  29449=>"011000111",
  29450=>"111110000",
  29451=>"100100001",
  29452=>"000110000",
  29453=>"111111111",
  29454=>"110010111",
  29455=>"111001000",
  29456=>"111101111",
  29457=>"000010001",
  29458=>"110101011",
  29459=>"001111010",
  29460=>"011100100",
  29461=>"110111100",
  29462=>"101011100",
  29463=>"111101111",
  29464=>"101001011",
  29465=>"000000100",
  29466=>"000110000",
  29467=>"000111100",
  29468=>"101010000",
  29469=>"101111011",
  29470=>"101010101",
  29471=>"011010110",
  29472=>"001000011",
  29473=>"101101100",
  29474=>"010010001",
  29475=>"111001111",
  29476=>"110110000",
  29477=>"001010000",
  29478=>"100010111",
  29479=>"010010100",
  29480=>"011100011",
  29481=>"100011100",
  29482=>"000010101",
  29483=>"000000010",
  29484=>"011011001",
  29485=>"101010111",
  29486=>"111110000",
  29487=>"001111110",
  29488=>"101101100",
  29489=>"100000111",
  29490=>"111100101",
  29491=>"111001110",
  29492=>"110011111",
  29493=>"110100011",
  29494=>"111001001",
  29495=>"001010101",
  29496=>"101010110",
  29497=>"000001000",
  29498=>"100000110",
  29499=>"011101011",
  29500=>"010010101",
  29501=>"101110001",
  29502=>"101000001",
  29503=>"011110111",
  29504=>"110100000",
  29505=>"010011110",
  29506=>"000001101",
  29507=>"110110110",
  29508=>"011000001",
  29509=>"001010011",
  29510=>"011011101",
  29511=>"111011111",
  29512=>"010011100",
  29513=>"110011000",
  29514=>"111100111",
  29515=>"001001001",
  29516=>"101000010",
  29517=>"010011000",
  29518=>"011111100",
  29519=>"101010000",
  29520=>"000100101",
  29521=>"100011111",
  29522=>"110000010",
  29523=>"010101110",
  29524=>"110101001",
  29525=>"101001100",
  29526=>"000111000",
  29527=>"010111010",
  29528=>"011010000",
  29529=>"010001000",
  29530=>"011111110",
  29531=>"011100001",
  29532=>"011111110",
  29533=>"100010101",
  29534=>"011110111",
  29535=>"011100110",
  29536=>"110010101",
  29537=>"001000100",
  29538=>"011111111",
  29539=>"111001001",
  29540=>"010001010",
  29541=>"110111000",
  29542=>"000001001",
  29543=>"100111010",
  29544=>"100111100",
  29545=>"101011000",
  29546=>"000111010",
  29547=>"011100101",
  29548=>"010010001",
  29549=>"011010010",
  29550=>"111010001",
  29551=>"011111100",
  29552=>"110111111",
  29553=>"110011111",
  29554=>"010100011",
  29555=>"100001111",
  29556=>"010111011",
  29557=>"101101001",
  29558=>"010111010",
  29559=>"110111110",
  29560=>"111011010",
  29561=>"011110010",
  29562=>"011010001",
  29563=>"111000001",
  29564=>"110110111",
  29565=>"101000100",
  29566=>"010111100",
  29567=>"001100000",
  29568=>"011010110",
  29569=>"010110110",
  29570=>"100101111",
  29571=>"010011010",
  29572=>"011110100",
  29573=>"001001010",
  29574=>"011011011",
  29575=>"001010010",
  29576=>"111111110",
  29577=>"011111100",
  29578=>"000100010",
  29579=>"001100000",
  29580=>"110101110",
  29581=>"001001111",
  29582=>"001111000",
  29583=>"100000010",
  29584=>"110010110",
  29585=>"110010110",
  29586=>"101101000",
  29587=>"110011000",
  29588=>"010110101",
  29589=>"011010110",
  29590=>"101100100",
  29591=>"111101101",
  29592=>"101010011",
  29593=>"010001001",
  29594=>"100010110",
  29595=>"011110101",
  29596=>"001100001",
  29597=>"100101111",
  29598=>"010101111",
  29599=>"011011010",
  29600=>"101101110",
  29601=>"011111101",
  29602=>"111001100",
  29603=>"110111101",
  29604=>"101100001",
  29605=>"001110101",
  29606=>"000010101",
  29607=>"010100001",
  29608=>"000010010",
  29609=>"000001011",
  29610=>"011011110",
  29611=>"111110001",
  29612=>"100001110",
  29613=>"010001111",
  29614=>"110110011",
  29615=>"011010111",
  29616=>"000110101",
  29617=>"010110011",
  29618=>"011100101",
  29619=>"110001011",
  29620=>"111001000",
  29621=>"001000010",
  29622=>"101010000",
  29623=>"010101000",
  29624=>"110000100",
  29625=>"110000110",
  29626=>"001100011",
  29627=>"000000000",
  29628=>"010110100",
  29629=>"101010100",
  29630=>"000101100",
  29631=>"001011101",
  29632=>"000101101",
  29633=>"100000101",
  29634=>"101100000",
  29635=>"101010110",
  29636=>"000000111",
  29637=>"101001011",
  29638=>"100011100",
  29639=>"011000110",
  29640=>"001001010",
  29641=>"100100100",
  29642=>"000000010",
  29643=>"000111100",
  29644=>"100101111",
  29645=>"000010001",
  29646=>"001110110",
  29647=>"111101011",
  29648=>"100111110",
  29649=>"110011001",
  29650=>"101110110",
  29651=>"011010101",
  29652=>"010110010",
  29653=>"001111101",
  29654=>"111100101",
  29655=>"011001110",
  29656=>"000000101",
  29657=>"000000100",
  29658=>"001000011",
  29659=>"111001111",
  29660=>"000101001",
  29661=>"110010101",
  29662=>"000001110",
  29663=>"100000001",
  29664=>"010101101",
  29665=>"001100101",
  29666=>"100010001",
  29667=>"110010110",
  29668=>"000111101",
  29669=>"100001000",
  29670=>"100110001",
  29671=>"010001001",
  29672=>"111100010",
  29673=>"100111011",
  29674=>"010111000",
  29675=>"001100111",
  29676=>"001011111",
  29677=>"010001001",
  29678=>"000010101",
  29679=>"001001110",
  29680=>"000011000",
  29681=>"100100100",
  29682=>"011101101",
  29683=>"000111111",
  29684=>"111110101",
  29685=>"001001101",
  29686=>"110000010",
  29687=>"011101110",
  29688=>"111011000",
  29689=>"000100011",
  29690=>"101100001",
  29691=>"010110111",
  29692=>"010101010",
  29693=>"101111000",
  29694=>"111011010",
  29695=>"000111111",
  29696=>"001101110",
  29697=>"010100010",
  29698=>"011100101",
  29699=>"011001000",
  29700=>"011001000",
  29701=>"010011000",
  29702=>"000001100",
  29703=>"110011100",
  29704=>"110111100",
  29705=>"101000110",
  29706=>"001001101",
  29707=>"100111000",
  29708=>"000111100",
  29709=>"011000011",
  29710=>"010100000",
  29711=>"101011001",
  29712=>"001001111",
  29713=>"001100100",
  29714=>"000011110",
  29715=>"001111111",
  29716=>"010010111",
  29717=>"011011111",
  29718=>"001111010",
  29719=>"000100011",
  29720=>"101000111",
  29721=>"000001110",
  29722=>"100000001",
  29723=>"010000101",
  29724=>"011010110",
  29725=>"110001000",
  29726=>"011110000",
  29727=>"100100001",
  29728=>"101010011",
  29729=>"010101001",
  29730=>"001110010",
  29731=>"111001001",
  29732=>"110010010",
  29733=>"110001010",
  29734=>"001101100",
  29735=>"101000110",
  29736=>"111011001",
  29737=>"101001010",
  29738=>"010011110",
  29739=>"000100000",
  29740=>"110111001",
  29741=>"011111100",
  29742=>"011000011",
  29743=>"000001111",
  29744=>"101100010",
  29745=>"110010010",
  29746=>"011010000",
  29747=>"100010001",
  29748=>"010001111",
  29749=>"110101101",
  29750=>"000000010",
  29751=>"111000011",
  29752=>"010100100",
  29753=>"011111111",
  29754=>"011100001",
  29755=>"011010101",
  29756=>"100011100",
  29757=>"100110001",
  29758=>"100110001",
  29759=>"110111100",
  29760=>"101110101",
  29761=>"010011100",
  29762=>"010000101",
  29763=>"001111000",
  29764=>"011001000",
  29765=>"110001010",
  29766=>"010010101",
  29767=>"110001010",
  29768=>"011010111",
  29769=>"000001101",
  29770=>"000000011",
  29771=>"000000110",
  29772=>"101101100",
  29773=>"111101100",
  29774=>"011010110",
  29775=>"100000011",
  29776=>"111001101",
  29777=>"100011110",
  29778=>"001110100",
  29779=>"100001100",
  29780=>"100010001",
  29781=>"110100000",
  29782=>"100110100",
  29783=>"111101011",
  29784=>"101011111",
  29785=>"010000100",
  29786=>"000000011",
  29787=>"100011000",
  29788=>"100000110",
  29789=>"011010010",
  29790=>"110000010",
  29791=>"010011100",
  29792=>"110011011",
  29793=>"000011100",
  29794=>"010010101",
  29795=>"111111101",
  29796=>"100011101",
  29797=>"111010011",
  29798=>"011001011",
  29799=>"111000111",
  29800=>"101000100",
  29801=>"010100100",
  29802=>"110011000",
  29803=>"001110110",
  29804=>"011110110",
  29805=>"111000010",
  29806=>"010010111",
  29807=>"011001110",
  29808=>"100001101",
  29809=>"111010010",
  29810=>"110011001",
  29811=>"110011010",
  29812=>"011010111",
  29813=>"111100010",
  29814=>"100100001",
  29815=>"111011010",
  29816=>"001001100",
  29817=>"000010010",
  29818=>"011010010",
  29819=>"100011101",
  29820=>"101100010",
  29821=>"001111100",
  29822=>"000001010",
  29823=>"101111010",
  29824=>"011000001",
  29825=>"011010111",
  29826=>"000101010",
  29827=>"100110110",
  29828=>"111101110",
  29829=>"100110111",
  29830=>"000101101",
  29831=>"010010000",
  29832=>"011110100",
  29833=>"001110000",
  29834=>"100000110",
  29835=>"111101110",
  29836=>"111110111",
  29837=>"111010100",
  29838=>"000011111",
  29839=>"101100100",
  29840=>"011111101",
  29841=>"110000010",
  29842=>"111100100",
  29843=>"110010010",
  29844=>"000100000",
  29845=>"110101001",
  29846=>"111001011",
  29847=>"110111011",
  29848=>"010001011",
  29849=>"100111100",
  29850=>"110001101",
  29851=>"011000001",
  29852=>"100101110",
  29853=>"111010000",
  29854=>"011110010",
  29855=>"101001110",
  29856=>"011100010",
  29857=>"010110010",
  29858=>"100000100",
  29859=>"110111100",
  29860=>"011011001",
  29861=>"000001000",
  29862=>"100010010",
  29863=>"001100110",
  29864=>"010111000",
  29865=>"110001100",
  29866=>"001110000",
  29867=>"111101101",
  29868=>"111100010",
  29869=>"000011001",
  29870=>"001101011",
  29871=>"011110000",
  29872=>"010111000",
  29873=>"010100110",
  29874=>"000001010",
  29875=>"101111111",
  29876=>"111000110",
  29877=>"100010000",
  29878=>"000101100",
  29879=>"011101011",
  29880=>"100001011",
  29881=>"001100000",
  29882=>"111110110",
  29883=>"010011110",
  29884=>"111010011",
  29885=>"111001101",
  29886=>"100011010",
  29887=>"001010000",
  29888=>"011001101",
  29889=>"000111110",
  29890=>"101000010",
  29891=>"011100101",
  29892=>"000111110",
  29893=>"000101010",
  29894=>"111001100",
  29895=>"001011100",
  29896=>"001110101",
  29897=>"100100101",
  29898=>"101100100",
  29899=>"001101110",
  29900=>"010001101",
  29901=>"100110101",
  29902=>"110100010",
  29903=>"010111100",
  29904=>"011011100",
  29905=>"011110111",
  29906=>"010100110",
  29907=>"010100111",
  29908=>"010101011",
  29909=>"110110100",
  29910=>"010001100",
  29911=>"101111111",
  29912=>"101001011",
  29913=>"011111110",
  29914=>"011001010",
  29915=>"000110100",
  29916=>"000101110",
  29917=>"000111010",
  29918=>"101001011",
  29919=>"111100011",
  29920=>"111000011",
  29921=>"000011001",
  29922=>"010000000",
  29923=>"000101000",
  29924=>"111001111",
  29925=>"010011100",
  29926=>"101000000",
  29927=>"010000011",
  29928=>"011100000",
  29929=>"010110011",
  29930=>"001000101",
  29931=>"000100100",
  29932=>"010010100",
  29933=>"111011000",
  29934=>"100001111",
  29935=>"011101011",
  29936=>"000111000",
  29937=>"001011101",
  29938=>"001001001",
  29939=>"000010000",
  29940=>"101111001",
  29941=>"010001100",
  29942=>"110000111",
  29943=>"111010100",
  29944=>"110110111",
  29945=>"101101100",
  29946=>"001001101",
  29947=>"000011110",
  29948=>"011111101",
  29949=>"000100000",
  29950=>"001100111",
  29951=>"001110101",
  29952=>"001011000",
  29953=>"110000111",
  29954=>"110101100",
  29955=>"101111010",
  29956=>"011000101",
  29957=>"001100001",
  29958=>"011010001",
  29959=>"100011110",
  29960=>"100011110",
  29961=>"010111101",
  29962=>"101010110",
  29963=>"010101010",
  29964=>"011010000",
  29965=>"010010101",
  29966=>"111100110",
  29967=>"000101000",
  29968=>"111101000",
  29969=>"101010101",
  29970=>"100010100",
  29971=>"011101000",
  29972=>"100001111",
  29973=>"001100001",
  29974=>"110000010",
  29975=>"111110001",
  29976=>"000000000",
  29977=>"100110000",
  29978=>"001011011",
  29979=>"101001010",
  29980=>"000111011",
  29981=>"111011001",
  29982=>"111101001",
  29983=>"011011111",
  29984=>"100010011",
  29985=>"000101011",
  29986=>"000001111",
  29987=>"110100110",
  29988=>"110000110",
  29989=>"001110010",
  29990=>"010110010",
  29991=>"000110100",
  29992=>"110010011",
  29993=>"011101100",
  29994=>"101011001",
  29995=>"111110110",
  29996=>"010100110",
  29997=>"001000111",
  29998=>"110011101",
  29999=>"001100101",
  30000=>"110000011",
  30001=>"011101101",
  30002=>"100100000",
  30003=>"100000100",
  30004=>"100111011",
  30005=>"011101101",
  30006=>"001001001",
  30007=>"100101011",
  30008=>"110011110",
  30009=>"110110010",
  30010=>"001000110",
  30011=>"100010011",
  30012=>"111110001",
  30013=>"011100000",
  30014=>"110100011",
  30015=>"011010110",
  30016=>"011100110",
  30017=>"101011010",
  30018=>"011001101",
  30019=>"010100000",
  30020=>"110010110",
  30021=>"110100100",
  30022=>"100110000",
  30023=>"110000011",
  30024=>"110000000",
  30025=>"011001100",
  30026=>"001000101",
  30027=>"010100010",
  30028=>"110101111",
  30029=>"101111111",
  30030=>"111011110",
  30031=>"111111011",
  30032=>"000011011",
  30033=>"110010011",
  30034=>"111101001",
  30035=>"110110001",
  30036=>"000110001",
  30037=>"011000111",
  30038=>"101001110",
  30039=>"100101111",
  30040=>"011100100",
  30041=>"100110111",
  30042=>"100000101",
  30043=>"000100100",
  30044=>"111011100",
  30045=>"010111110",
  30046=>"000110011",
  30047=>"101100001",
  30048=>"001101110",
  30049=>"011001110",
  30050=>"001111011",
  30051=>"100110101",
  30052=>"010001101",
  30053=>"101001011",
  30054=>"100110001",
  30055=>"111011010",
  30056=>"101101001",
  30057=>"000011000",
  30058=>"110001000",
  30059=>"011010100",
  30060=>"111011100",
  30061=>"000001000",
  30062=>"110010001",
  30063=>"001111011",
  30064=>"000111011",
  30065=>"110011111",
  30066=>"111101101",
  30067=>"111110011",
  30068=>"110101110",
  30069=>"100100111",
  30070=>"001000110",
  30071=>"111010001",
  30072=>"000101010",
  30073=>"001110010",
  30074=>"101110100",
  30075=>"000111111",
  30076=>"000111011",
  30077=>"100101101",
  30078=>"111110011",
  30079=>"101110000",
  30080=>"011100000",
  30081=>"000100110",
  30082=>"101110011",
  30083=>"000101100",
  30084=>"111010110",
  30085=>"111110110",
  30086=>"111101100",
  30087=>"110000110",
  30088=>"101000000",
  30089=>"011010111",
  30090=>"001100001",
  30091=>"010011010",
  30092=>"000000000",
  30093=>"101011010",
  30094=>"110000111",
  30095=>"001100100",
  30096=>"111111100",
  30097=>"001011111",
  30098=>"110110111",
  30099=>"101101000",
  30100=>"110100011",
  30101=>"101100111",
  30102=>"000111111",
  30103=>"010011001",
  30104=>"110111001",
  30105=>"010001110",
  30106=>"000011001",
  30107=>"010101010",
  30108=>"101101111",
  30109=>"101000001",
  30110=>"111110111",
  30111=>"101011110",
  30112=>"000001101",
  30113=>"001101101",
  30114=>"001011101",
  30115=>"100111110",
  30116=>"100001101",
  30117=>"100100000",
  30118=>"100110111",
  30119=>"111100001",
  30120=>"101100111",
  30121=>"110010000",
  30122=>"100111010",
  30123=>"010001001",
  30124=>"000000000",
  30125=>"110100000",
  30126=>"011010101",
  30127=>"100100000",
  30128=>"101110010",
  30129=>"011010001",
  30130=>"100011101",
  30131=>"111001001",
  30132=>"000010100",
  30133=>"110101101",
  30134=>"111011101",
  30135=>"100100001",
  30136=>"000101001",
  30137=>"110010010",
  30138=>"100101100",
  30139=>"001010000",
  30140=>"000110001",
  30141=>"001100011",
  30142=>"111011010",
  30143=>"000100001",
  30144=>"101000010",
  30145=>"010011100",
  30146=>"010111011",
  30147=>"111001100",
  30148=>"100010010",
  30149=>"010110111",
  30150=>"011000101",
  30151=>"101100001",
  30152=>"001100010",
  30153=>"011000101",
  30154=>"111110100",
  30155=>"110111011",
  30156=>"111111011",
  30157=>"110010001",
  30158=>"101100010",
  30159=>"100111111",
  30160=>"011010001",
  30161=>"000110110",
  30162=>"010011101",
  30163=>"010100001",
  30164=>"111010000",
  30165=>"111111100",
  30166=>"011100001",
  30167=>"011100101",
  30168=>"111101011",
  30169=>"010000101",
  30170=>"001110110",
  30171=>"101000010",
  30172=>"000011010",
  30173=>"111011110",
  30174=>"101000100",
  30175=>"010011110",
  30176=>"101111000",
  30177=>"010010010",
  30178=>"001000011",
  30179=>"101011111",
  30180=>"011111100",
  30181=>"101010000",
  30182=>"110010110",
  30183=>"101011001",
  30184=>"100000100",
  30185=>"101000000",
  30186=>"101110101",
  30187=>"000000001",
  30188=>"101011001",
  30189=>"000010010",
  30190=>"000010101",
  30191=>"101000001",
  30192=>"110100100",
  30193=>"000010010",
  30194=>"100001011",
  30195=>"000000010",
  30196=>"111010001",
  30197=>"001100000",
  30198=>"110100000",
  30199=>"110111011",
  30200=>"010000001",
  30201=>"000001001",
  30202=>"010100101",
  30203=>"111100101",
  30204=>"000110101",
  30205=>"110110001",
  30206=>"101010101",
  30207=>"100001010",
  30208=>"110110100",
  30209=>"010101100",
  30210=>"001111100",
  30211=>"100101011",
  30212=>"110111001",
  30213=>"110001001",
  30214=>"111010000",
  30215=>"111101110",
  30216=>"000010101",
  30217=>"001011010",
  30218=>"000111110",
  30219=>"001001111",
  30220=>"011111001",
  30221=>"101101011",
  30222=>"000000110",
  30223=>"101100100",
  30224=>"100000001",
  30225=>"001001010",
  30226=>"110110101",
  30227=>"111010011",
  30228=>"101011010",
  30229=>"001010011",
  30230=>"100001010",
  30231=>"100011100",
  30232=>"101001111",
  30233=>"001010000",
  30234=>"001011111",
  30235=>"111100100",
  30236=>"010010110",
  30237=>"011111000",
  30238=>"000010011",
  30239=>"000110111",
  30240=>"010000111",
  30241=>"100010100",
  30242=>"100010010",
  30243=>"100110011",
  30244=>"010001000",
  30245=>"111110011",
  30246=>"000111110",
  30247=>"011010100",
  30248=>"001101001",
  30249=>"000011101",
  30250=>"000000010",
  30251=>"000111101",
  30252=>"111101000",
  30253=>"011100010",
  30254=>"010001010",
  30255=>"011110010",
  30256=>"001101001",
  30257=>"000111101",
  30258=>"011110010",
  30259=>"100110101",
  30260=>"100111110",
  30261=>"000010111",
  30262=>"001011000",
  30263=>"110111101",
  30264=>"000011110",
  30265=>"110110001",
  30266=>"110101011",
  30267=>"000100111",
  30268=>"001001011",
  30269=>"101011010",
  30270=>"000000011",
  30271=>"101100110",
  30272=>"000011100",
  30273=>"100110110",
  30274=>"000010011",
  30275=>"000111010",
  30276=>"010101100",
  30277=>"000110110",
  30278=>"010001110",
  30279=>"011001110",
  30280=>"010101100",
  30281=>"000000010",
  30282=>"101101111",
  30283=>"101111010",
  30284=>"100000011",
  30285=>"000010011",
  30286=>"100001001",
  30287=>"010110111",
  30288=>"011101011",
  30289=>"100000010",
  30290=>"001110101",
  30291=>"010010011",
  30292=>"110000111",
  30293=>"010111010",
  30294=>"111011100",
  30295=>"000100000",
  30296=>"110010100",
  30297=>"101010101",
  30298=>"100000010",
  30299=>"110111101",
  30300=>"001110010",
  30301=>"000010010",
  30302=>"100001001",
  30303=>"101111100",
  30304=>"010000100",
  30305=>"010000011",
  30306=>"101000001",
  30307=>"110001001",
  30308=>"110011011",
  30309=>"111111010",
  30310=>"110110101",
  30311=>"111001100",
  30312=>"110011010",
  30313=>"100011101",
  30314=>"000101111",
  30315=>"000100011",
  30316=>"011010010",
  30317=>"111011011",
  30318=>"101110010",
  30319=>"111011000",
  30320=>"010100010",
  30321=>"011010101",
  30322=>"100110101",
  30323=>"110101000",
  30324=>"010010010",
  30325=>"111001101",
  30326=>"101111011",
  30327=>"000011101",
  30328=>"000000010",
  30329=>"001101101",
  30330=>"001111110",
  30331=>"110011100",
  30332=>"111110000",
  30333=>"101100001",
  30334=>"000110000",
  30335=>"000001101",
  30336=>"101000100",
  30337=>"111111001",
  30338=>"011010110",
  30339=>"010010010",
  30340=>"011111000",
  30341=>"001100110",
  30342=>"101111010",
  30343=>"111010111",
  30344=>"011101110",
  30345=>"010010010",
  30346=>"100110010",
  30347=>"011011111",
  30348=>"111011010",
  30349=>"110010000",
  30350=>"111101100",
  30351=>"100000000",
  30352=>"101101100",
  30353=>"111100111",
  30354=>"010100110",
  30355=>"011011000",
  30356=>"110011100",
  30357=>"000001001",
  30358=>"010101011",
  30359=>"011010101",
  30360=>"110001001",
  30361=>"100000110",
  30362=>"100011001",
  30363=>"101001101",
  30364=>"000001011",
  30365=>"001110101",
  30366=>"100000101",
  30367=>"100101111",
  30368=>"110100001",
  30369=>"111010100",
  30370=>"011111100",
  30371=>"001111011",
  30372=>"100010101",
  30373=>"011001010",
  30374=>"010000000",
  30375=>"101100101",
  30376=>"000100010",
  30377=>"000101010",
  30378=>"010100100",
  30379=>"000001100",
  30380=>"110100111",
  30381=>"110001110",
  30382=>"001100011",
  30383=>"001011001",
  30384=>"110011001",
  30385=>"011100110",
  30386=>"000100100",
  30387=>"011101011",
  30388=>"001010101",
  30389=>"001101111",
  30390=>"000010001",
  30391=>"110111110",
  30392=>"011101111",
  30393=>"010011100",
  30394=>"100101001",
  30395=>"101001101",
  30396=>"010100000",
  30397=>"000001011",
  30398=>"010010110",
  30399=>"011111011",
  30400=>"000010100",
  30401=>"010000101",
  30402=>"101000100",
  30403=>"000011000",
  30404=>"110000000",
  30405=>"011001001",
  30406=>"001110111",
  30407=>"001111101",
  30408=>"110000100",
  30409=>"010011000",
  30410=>"010011001",
  30411=>"111100100",
  30412=>"101000110",
  30413=>"011100000",
  30414=>"111001010",
  30415=>"010100011",
  30416=>"111101111",
  30417=>"100000110",
  30418=>"110101010",
  30419=>"000001100",
  30420=>"011010110",
  30421=>"101010011",
  30422=>"010001001",
  30423=>"000011000",
  30424=>"011101001",
  30425=>"111010101",
  30426=>"110001100",
  30427=>"011000001",
  30428=>"010110011",
  30429=>"110001111",
  30430=>"110010111",
  30431=>"111110011",
  30432=>"011010000",
  30433=>"110101101",
  30434=>"100111010",
  30435=>"110110001",
  30436=>"101101010",
  30437=>"011111001",
  30438=>"110100110",
  30439=>"100110111",
  30440=>"011110010",
  30441=>"110011100",
  30442=>"100110101",
  30443=>"110001101",
  30444=>"010000010",
  30445=>"001001010",
  30446=>"111000110",
  30447=>"001011011",
  30448=>"101111001",
  30449=>"111001110",
  30450=>"001010011",
  30451=>"111110001",
  30452=>"010011000",
  30453=>"101001011",
  30454=>"000000101",
  30455=>"100110110",
  30456=>"110110001",
  30457=>"000101011",
  30458=>"001010001",
  30459=>"101111101",
  30460=>"011101010",
  30461=>"101000001",
  30462=>"010000111",
  30463=>"010011101",
  30464=>"111101110",
  30465=>"110100100",
  30466=>"111101100",
  30467=>"000011010",
  30468=>"001011011",
  30469=>"000101010",
  30470=>"101001010",
  30471=>"010000010",
  30472=>"111111101",
  30473=>"111000010",
  30474=>"101001011",
  30475=>"111010010",
  30476=>"011001010",
  30477=>"110110101",
  30478=>"010000110",
  30479=>"001000101",
  30480=>"110010011",
  30481=>"101110100",
  30482=>"000000110",
  30483=>"001100011",
  30484=>"001111111",
  30485=>"101001111",
  30486=>"111010010",
  30487=>"101111011",
  30488=>"010011000",
  30489=>"111111000",
  30490=>"100110111",
  30491=>"101101011",
  30492=>"111011110",
  30493=>"000101100",
  30494=>"101000010",
  30495=>"011100010",
  30496=>"001010100",
  30497=>"101011101",
  30498=>"100100111",
  30499=>"000000111",
  30500=>"010101000",
  30501=>"000110011",
  30502=>"101110111",
  30503=>"101110000",
  30504=>"111011011",
  30505=>"100101000",
  30506=>"101010110",
  30507=>"101010100",
  30508=>"111101001",
  30509=>"001011001",
  30510=>"010111101",
  30511=>"010001000",
  30512=>"010111011",
  30513=>"001111001",
  30514=>"001000110",
  30515=>"110111010",
  30516=>"100000011",
  30517=>"010100011",
  30518=>"100111011",
  30519=>"011111001",
  30520=>"001000101",
  30521=>"011101100",
  30522=>"111010100",
  30523=>"000111000",
  30524=>"111101010",
  30525=>"101001111",
  30526=>"011010010",
  30527=>"100110010",
  30528=>"011011111",
  30529=>"110111111",
  30530=>"100100100",
  30531=>"011010000",
  30532=>"001001011",
  30533=>"000110101",
  30534=>"011111110",
  30535=>"010001101",
  30536=>"110000111",
  30537=>"111001011",
  30538=>"000101010",
  30539=>"101011001",
  30540=>"111100001",
  30541=>"000111100",
  30542=>"101000111",
  30543=>"100011101",
  30544=>"011110001",
  30545=>"000001000",
  30546=>"001101011",
  30547=>"110001011",
  30548=>"100001011",
  30549=>"010010111",
  30550=>"111010000",
  30551=>"010101011",
  30552=>"011010010",
  30553=>"111011100",
  30554=>"001110101",
  30555=>"001001101",
  30556=>"010001011",
  30557=>"101001110",
  30558=>"011101111",
  30559=>"010111000",
  30560=>"100001000",
  30561=>"000000000",
  30562=>"011101001",
  30563=>"100101111",
  30564=>"010110101",
  30565=>"101001000",
  30566=>"110000101",
  30567=>"010101010",
  30568=>"001100101",
  30569=>"100111010",
  30570=>"111111111",
  30571=>"010011111",
  30572=>"010100000",
  30573=>"011100100",
  30574=>"011000000",
  30575=>"100100001",
  30576=>"011011010",
  30577=>"000111010",
  30578=>"101100001",
  30579=>"000111111",
  30580=>"000101100",
  30581=>"101010111",
  30582=>"010100100",
  30583=>"110000011",
  30584=>"011100000",
  30585=>"001101000",
  30586=>"100110110",
  30587=>"000111100",
  30588=>"011011010",
  30589=>"010000100",
  30590=>"001100001",
  30591=>"001001110",
  30592=>"110011101",
  30593=>"110000100",
  30594=>"000100101",
  30595=>"000101101",
  30596=>"011010010",
  30597=>"010010111",
  30598=>"011010011",
  30599=>"001111000",
  30600=>"100010100",
  30601=>"001010110",
  30602=>"101000101",
  30603=>"000000000",
  30604=>"111101010",
  30605=>"100000001",
  30606=>"111110010",
  30607=>"101111001",
  30608=>"110011110",
  30609=>"111101011",
  30610=>"010100001",
  30611=>"100100011",
  30612=>"000000101",
  30613=>"100011100",
  30614=>"100101000",
  30615=>"010111000",
  30616=>"110100111",
  30617=>"101100001",
  30618=>"001100100",
  30619=>"110101110",
  30620=>"011100110",
  30621=>"100001011",
  30622=>"111100011",
  30623=>"011011000",
  30624=>"001110001",
  30625=>"100100101",
  30626=>"000111001",
  30627=>"000010001",
  30628=>"000101000",
  30629=>"111000010",
  30630=>"010001000",
  30631=>"000011010",
  30632=>"011101011",
  30633=>"111100000",
  30634=>"000011111",
  30635=>"100010110",
  30636=>"101111010",
  30637=>"101100001",
  30638=>"000101111",
  30639=>"100010010",
  30640=>"000010110",
  30641=>"000101000",
  30642=>"001100001",
  30643=>"011111100",
  30644=>"100100000",
  30645=>"000111111",
  30646=>"101111000",
  30647=>"001111111",
  30648=>"101010001",
  30649=>"110001001",
  30650=>"100001010",
  30651=>"100100101",
  30652=>"010101010",
  30653=>"000101010",
  30654=>"011100100",
  30655=>"010010011",
  30656=>"001001100",
  30657=>"101110011",
  30658=>"111111011",
  30659=>"110011101",
  30660=>"100010110",
  30661=>"011000001",
  30662=>"110101001",
  30663=>"100010101",
  30664=>"110101000",
  30665=>"010000000",
  30666=>"000111001",
  30667=>"011001001",
  30668=>"010111010",
  30669=>"010100000",
  30670=>"100011110",
  30671=>"111001110",
  30672=>"011101011",
  30673=>"110100111",
  30674=>"010100000",
  30675=>"000110001",
  30676=>"100111100",
  30677=>"011101001",
  30678=>"010100111",
  30679=>"011100001",
  30680=>"100000001",
  30681=>"101001111",
  30682=>"100011010",
  30683=>"110111111",
  30684=>"101011010",
  30685=>"101011000",
  30686=>"110000111",
  30687=>"011100111",
  30688=>"110100010",
  30689=>"011111011",
  30690=>"001000001",
  30691=>"010001011",
  30692=>"100000110",
  30693=>"011010001",
  30694=>"000001010",
  30695=>"000010100",
  30696=>"110101111",
  30697=>"011000011",
  30698=>"010000000",
  30699=>"100000001",
  30700=>"110101101",
  30701=>"100010111",
  30702=>"010100000",
  30703=>"110110001",
  30704=>"001000111",
  30705=>"011110011",
  30706=>"101111001",
  30707=>"110001101",
  30708=>"011000000",
  30709=>"001000100",
  30710=>"000010010",
  30711=>"111111001",
  30712=>"101010110",
  30713=>"011001010",
  30714=>"111011011",
  30715=>"101101001",
  30716=>"100000110",
  30717=>"111111101",
  30718=>"000111110",
  30719=>"101000101",
  30720=>"000110001",
  30721=>"000110010",
  30722=>"001010000",
  30723=>"000101010",
  30724=>"000001000",
  30725=>"010110011",
  30726=>"000000100",
  30727=>"000010001",
  30728=>"111000001",
  30729=>"001110101",
  30730=>"111000011",
  30731=>"010001111",
  30732=>"010000011",
  30733=>"111101001",
  30734=>"011000000",
  30735=>"010000101",
  30736=>"110011001",
  30737=>"010001101",
  30738=>"111011110",
  30739=>"100111000",
  30740=>"111111111",
  30741=>"011000011",
  30742=>"001010110",
  30743=>"010111111",
  30744=>"101000111",
  30745=>"011011100",
  30746=>"011011001",
  30747=>"010001010",
  30748=>"111011111",
  30749=>"111010111",
  30750=>"100110110",
  30751=>"010101010",
  30752=>"011110010",
  30753=>"110100110",
  30754=>"110111000",
  30755=>"010110001",
  30756=>"010000000",
  30757=>"000001010",
  30758=>"000000011",
  30759=>"000000110",
  30760=>"110001011",
  30761=>"000111010",
  30762=>"010010000",
  30763=>"111111011",
  30764=>"111111000",
  30765=>"010011011",
  30766=>"000000111",
  30767=>"100110111",
  30768=>"101000111",
  30769=>"001110000",
  30770=>"010010000",
  30771=>"000000111",
  30772=>"110101111",
  30773=>"101001010",
  30774=>"101010010",
  30775=>"111001101",
  30776=>"000011010",
  30777=>"101011101",
  30778=>"000001000",
  30779=>"001110011",
  30780=>"111001001",
  30781=>"001110000",
  30782=>"011111110",
  30783=>"111010000",
  30784=>"101010001",
  30785=>"000000100",
  30786=>"111111000",
  30787=>"101111100",
  30788=>"111110000",
  30789=>"101110010",
  30790=>"110010010",
  30791=>"110001000",
  30792=>"001111000",
  30793=>"001100100",
  30794=>"000001011",
  30795=>"010100000",
  30796=>"110000111",
  30797=>"111110111",
  30798=>"111011000",
  30799=>"110100100",
  30800=>"000110111",
  30801=>"011100101",
  30802=>"000111111",
  30803=>"111011111",
  30804=>"101010001",
  30805=>"010000010",
  30806=>"011111110",
  30807=>"001111101",
  30808=>"111001001",
  30809=>"101101100",
  30810=>"101100100",
  30811=>"111010000",
  30812=>"011101101",
  30813=>"101100101",
  30814=>"000111000",
  30815=>"000100000",
  30816=>"011010010",
  30817=>"011101111",
  30818=>"100110011",
  30819=>"001001011",
  30820=>"000111010",
  30821=>"011010001",
  30822=>"100011001",
  30823=>"110010011",
  30824=>"111101010",
  30825=>"111101011",
  30826=>"101110000",
  30827=>"001011000",
  30828=>"101011100",
  30829=>"100000010",
  30830=>"011111100",
  30831=>"001011010",
  30832=>"011110100",
  30833=>"111101011",
  30834=>"111111001",
  30835=>"110000011",
  30836=>"000011011",
  30837=>"111010100",
  30838=>"101101001",
  30839=>"110000011",
  30840=>"011001000",
  30841=>"000000000",
  30842=>"010111111",
  30843=>"000010010",
  30844=>"011000011",
  30845=>"110000101",
  30846=>"011000101",
  30847=>"111011011",
  30848=>"001000010",
  30849=>"001011100",
  30850=>"111010001",
  30851=>"111101000",
  30852=>"110001000",
  30853=>"000100011",
  30854=>"001001111",
  30855=>"101001011",
  30856=>"000110101",
  30857=>"001111111",
  30858=>"011110010",
  30859=>"001110001",
  30860=>"101101100",
  30861=>"110110011",
  30862=>"001100100",
  30863=>"000011101",
  30864=>"000001011",
  30865=>"010001100",
  30866=>"100101001",
  30867=>"110110100",
  30868=>"100101111",
  30869=>"001111101",
  30870=>"110011001",
  30871=>"100001011",
  30872=>"000101011",
  30873=>"010011010",
  30874=>"001010000",
  30875=>"100100011",
  30876=>"001101010",
  30877=>"011100100",
  30878=>"000100111",
  30879=>"101101000",
  30880=>"101100111",
  30881=>"001000000",
  30882=>"110011101",
  30883=>"010000011",
  30884=>"111111010",
  30885=>"100111001",
  30886=>"111101010",
  30887=>"101000011",
  30888=>"111111111",
  30889=>"111011110",
  30890=>"010100010",
  30891=>"111001100",
  30892=>"101111110",
  30893=>"111111101",
  30894=>"010010000",
  30895=>"001111110",
  30896=>"001010000",
  30897=>"111000110",
  30898=>"100101001",
  30899=>"111010000",
  30900=>"011111001",
  30901=>"100000111",
  30902=>"111111111",
  30903=>"111001111",
  30904=>"111000010",
  30905=>"001011100",
  30906=>"111111111",
  30907=>"111000101",
  30908=>"000100000",
  30909=>"000110111",
  30910=>"011100111",
  30911=>"101010001",
  30912=>"111100111",
  30913=>"100100011",
  30914=>"000101000",
  30915=>"000110011",
  30916=>"000000110",
  30917=>"000101001",
  30918=>"110110000",
  30919=>"110101111",
  30920=>"001010001",
  30921=>"111101010",
  30922=>"111001100",
  30923=>"001100111",
  30924=>"100001011",
  30925=>"101010011",
  30926=>"001001000",
  30927=>"011011001",
  30928=>"001001000",
  30929=>"110010000",
  30930=>"001001110",
  30931=>"000010100",
  30932=>"101111001",
  30933=>"001101000",
  30934=>"100111100",
  30935=>"010110110",
  30936=>"010111001",
  30937=>"110010010",
  30938=>"110110001",
  30939=>"100101001",
  30940=>"111010110",
  30941=>"010010011",
  30942=>"010011010",
  30943=>"010001010",
  30944=>"111101111",
  30945=>"110110101",
  30946=>"010010100",
  30947=>"100101100",
  30948=>"111001011",
  30949=>"110111101",
  30950=>"010100101",
  30951=>"010110111",
  30952=>"100111001",
  30953=>"101001010",
  30954=>"110000111",
  30955=>"001000101",
  30956=>"100011000",
  30957=>"011001101",
  30958=>"001011001",
  30959=>"011001001",
  30960=>"010010111",
  30961=>"101111111",
  30962=>"110100000",
  30963=>"000001001",
  30964=>"001111000",
  30965=>"000111111",
  30966=>"100011011",
  30967=>"000001001",
  30968=>"100011011",
  30969=>"010010011",
  30970=>"100101010",
  30971=>"111111010",
  30972=>"110100101",
  30973=>"000001110",
  30974=>"011011000",
  30975=>"110100000",
  30976=>"101101101",
  30977=>"110000011",
  30978=>"110011111",
  30979=>"010110000",
  30980=>"001011100",
  30981=>"001101111",
  30982=>"111001100",
  30983=>"000011011",
  30984=>"100000010",
  30985=>"100000011",
  30986=>"110001101",
  30987=>"000101001",
  30988=>"011110011",
  30989=>"101101111",
  30990=>"100000101",
  30991=>"101011000",
  30992=>"010101111",
  30993=>"010100011",
  30994=>"111010001",
  30995=>"010111111",
  30996=>"101000101",
  30997=>"100111110",
  30998=>"101100111",
  30999=>"111001010",
  31000=>"000001010",
  31001=>"100000010",
  31002=>"010000110",
  31003=>"111100000",
  31004=>"111000011",
  31005=>"100010110",
  31006=>"110111111",
  31007=>"110101100",
  31008=>"110100011",
  31009=>"001011010",
  31010=>"011011011",
  31011=>"101000001",
  31012=>"000001011",
  31013=>"100010011",
  31014=>"100001001",
  31015=>"001010111",
  31016=>"010101011",
  31017=>"110010111",
  31018=>"111101100",
  31019=>"110101010",
  31020=>"000111010",
  31021=>"101001101",
  31022=>"010010000",
  31023=>"111010111",
  31024=>"001010000",
  31025=>"000010010",
  31026=>"011110000",
  31027=>"011010100",
  31028=>"110011010",
  31029=>"010000010",
  31030=>"000000010",
  31031=>"000111110",
  31032=>"001011101",
  31033=>"100110001",
  31034=>"010001110",
  31035=>"011111111",
  31036=>"001110001",
  31037=>"110101111",
  31038=>"000100001",
  31039=>"000111000",
  31040=>"111111111",
  31041=>"000010101",
  31042=>"000000110",
  31043=>"001101111",
  31044=>"000111101",
  31045=>"001110001",
  31046=>"110001101",
  31047=>"110111110",
  31048=>"111011100",
  31049=>"110000101",
  31050=>"001000110",
  31051=>"111101110",
  31052=>"101101011",
  31053=>"100001001",
  31054=>"111000101",
  31055=>"010111001",
  31056=>"110101011",
  31057=>"100101000",
  31058=>"000110001",
  31059=>"101100001",
  31060=>"000001010",
  31061=>"010001110",
  31062=>"100011000",
  31063=>"100011011",
  31064=>"100010000",
  31065=>"010010101",
  31066=>"111100111",
  31067=>"011011010",
  31068=>"101101100",
  31069=>"010001111",
  31070=>"111000000",
  31071=>"110010010",
  31072=>"011111010",
  31073=>"001011001",
  31074=>"001000010",
  31075=>"001001110",
  31076=>"101100101",
  31077=>"001100100",
  31078=>"111100100",
  31079=>"000000010",
  31080=>"010011011",
  31081=>"000001011",
  31082=>"110111101",
  31083=>"111110010",
  31084=>"010000010",
  31085=>"110011101",
  31086=>"110010110",
  31087=>"000000001",
  31088=>"000100011",
  31089=>"111101101",
  31090=>"001101001",
  31091=>"110000000",
  31092=>"101100100",
  31093=>"110000101",
  31094=>"001010001",
  31095=>"110000111",
  31096=>"101111101",
  31097=>"101111001",
  31098=>"000100111",
  31099=>"000101100",
  31100=>"111111101",
  31101=>"011110010",
  31102=>"100010010",
  31103=>"101000111",
  31104=>"011100010",
  31105=>"001100001",
  31106=>"010110111",
  31107=>"110000001",
  31108=>"111101000",
  31109=>"000000001",
  31110=>"011110010",
  31111=>"000110000",
  31112=>"000010111",
  31113=>"000110111",
  31114=>"111101000",
  31115=>"001111100",
  31116=>"010101100",
  31117=>"010011001",
  31118=>"101010101",
  31119=>"011111010",
  31120=>"110011001",
  31121=>"001000100",
  31122=>"010011111",
  31123=>"110101010",
  31124=>"101111111",
  31125=>"000010000",
  31126=>"011110011",
  31127=>"111010101",
  31128=>"110010000",
  31129=>"000100101",
  31130=>"000100101",
  31131=>"100100010",
  31132=>"000010001",
  31133=>"001000110",
  31134=>"001000010",
  31135=>"111101110",
  31136=>"010110011",
  31137=>"010111011",
  31138=>"101111001",
  31139=>"010010111",
  31140=>"101110000",
  31141=>"111100001",
  31142=>"010010100",
  31143=>"001000111",
  31144=>"100100111",
  31145=>"010010000",
  31146=>"111101101",
  31147=>"001110010",
  31148=>"011111010",
  31149=>"000010100",
  31150=>"000111101",
  31151=>"101110101",
  31152=>"000110100",
  31153=>"001110011",
  31154=>"000101000",
  31155=>"001000011",
  31156=>"011011101",
  31157=>"011111101",
  31158=>"011101001",
  31159=>"010011101",
  31160=>"101101000",
  31161=>"100110100",
  31162=>"011111101",
  31163=>"011111101",
  31164=>"011000101",
  31165=>"000011011",
  31166=>"111011110",
  31167=>"001010000",
  31168=>"100001010",
  31169=>"010100110",
  31170=>"001110100",
  31171=>"011001001",
  31172=>"110110111",
  31173=>"100001111",
  31174=>"111111011",
  31175=>"101110000",
  31176=>"100000001",
  31177=>"001100101",
  31178=>"000000000",
  31179=>"110101011",
  31180=>"101101000",
  31181=>"110101110",
  31182=>"100000101",
  31183=>"011110100",
  31184=>"111111111",
  31185=>"010110000",
  31186=>"001101110",
  31187=>"101101010",
  31188=>"011101111",
  31189=>"010110001",
  31190=>"010100001",
  31191=>"001000010",
  31192=>"001011011",
  31193=>"001111101",
  31194=>"011111001",
  31195=>"111010010",
  31196=>"101010010",
  31197=>"011111010",
  31198=>"001001100",
  31199=>"011000001",
  31200=>"011110110",
  31201=>"011010000",
  31202=>"011100100",
  31203=>"010011000",
  31204=>"101101111",
  31205=>"101000011",
  31206=>"010011011",
  31207=>"100000001",
  31208=>"110111001",
  31209=>"001111110",
  31210=>"011000010",
  31211=>"101000100",
  31212=>"010010110",
  31213=>"111101000",
  31214=>"111001101",
  31215=>"000010010",
  31216=>"110101110",
  31217=>"000011001",
  31218=>"000010100",
  31219=>"011011100",
  31220=>"101100010",
  31221=>"100111010",
  31222=>"101000011",
  31223=>"000000000",
  31224=>"100101111",
  31225=>"011101010",
  31226=>"101010101",
  31227=>"111111111",
  31228=>"001001100",
  31229=>"110111101",
  31230=>"011111001",
  31231=>"000010101",
  31232=>"100011111",
  31233=>"001100110",
  31234=>"101001001",
  31235=>"100100110",
  31236=>"011101011",
  31237=>"011001001",
  31238=>"000100010",
  31239=>"010000111",
  31240=>"111000110",
  31241=>"111110111",
  31242=>"110100110",
  31243=>"100011000",
  31244=>"011011101",
  31245=>"110010111",
  31246=>"000100100",
  31247=>"011111111",
  31248=>"011101010",
  31249=>"010111101",
  31250=>"000111101",
  31251=>"010010011",
  31252=>"010001000",
  31253=>"111101001",
  31254=>"011000000",
  31255=>"001111101",
  31256=>"101001100",
  31257=>"100000011",
  31258=>"111010011",
  31259=>"101000000",
  31260=>"000001111",
  31261=>"000000000",
  31262=>"001111110",
  31263=>"111011110",
  31264=>"100110000",
  31265=>"001001101",
  31266=>"100001101",
  31267=>"111110101",
  31268=>"010110001",
  31269=>"000101001",
  31270=>"011101001",
  31271=>"100001110",
  31272=>"000000001",
  31273=>"100101100",
  31274=>"011011000",
  31275=>"100100110",
  31276=>"010110101",
  31277=>"111001100",
  31278=>"000100110",
  31279=>"000000101",
  31280=>"010110110",
  31281=>"000001111",
  31282=>"001111000",
  31283=>"110110111",
  31284=>"100111011",
  31285=>"011000110",
  31286=>"111100111",
  31287=>"101111111",
  31288=>"101000000",
  31289=>"100111010",
  31290=>"011001110",
  31291=>"000000110",
  31292=>"110110000",
  31293=>"111100000",
  31294=>"000011001",
  31295=>"111011000",
  31296=>"101100100",
  31297=>"011111101",
  31298=>"111001100",
  31299=>"010111001",
  31300=>"101100101",
  31301=>"101010101",
  31302=>"110111000",
  31303=>"000001110",
  31304=>"110101100",
  31305=>"010100110",
  31306=>"110110011",
  31307=>"100100010",
  31308=>"111110000",
  31309=>"000000111",
  31310=>"100111111",
  31311=>"100011110",
  31312=>"111000010",
  31313=>"111010001",
  31314=>"101001111",
  31315=>"100000110",
  31316=>"001011011",
  31317=>"000010101",
  31318=>"010011010",
  31319=>"010110101",
  31320=>"101000000",
  31321=>"100110011",
  31322=>"001011010",
  31323=>"001011000",
  31324=>"000000000",
  31325=>"100100110",
  31326=>"011010101",
  31327=>"111100000",
  31328=>"101001100",
  31329=>"001001111",
  31330=>"111101101",
  31331=>"100100001",
  31332=>"101000101",
  31333=>"001000011",
  31334=>"101000011",
  31335=>"100011101",
  31336=>"011100010",
  31337=>"110001000",
  31338=>"110010010",
  31339=>"010011100",
  31340=>"010001100",
  31341=>"011101100",
  31342=>"101111110",
  31343=>"111011111",
  31344=>"010101011",
  31345=>"100110110",
  31346=>"011101101",
  31347=>"011101011",
  31348=>"101111111",
  31349=>"000011010",
  31350=>"111111110",
  31351=>"011000101",
  31352=>"111000100",
  31353=>"111110100",
  31354=>"011000011",
  31355=>"011001011",
  31356=>"001000001",
  31357=>"110101001",
  31358=>"111000100",
  31359=>"010111100",
  31360=>"010111111",
  31361=>"100110000",
  31362=>"011100001",
  31363=>"100100001",
  31364=>"100110110",
  31365=>"110000111",
  31366=>"110110010",
  31367=>"011100000",
  31368=>"111110111",
  31369=>"000000010",
  31370=>"100101000",
  31371=>"000110011",
  31372=>"011000000",
  31373=>"000000010",
  31374=>"010001110",
  31375=>"010000101",
  31376=>"101001111",
  31377=>"101010101",
  31378=>"100001010",
  31379=>"101111111",
  31380=>"101010100",
  31381=>"001111000",
  31382=>"001000110",
  31383=>"110110000",
  31384=>"101011111",
  31385=>"111010000",
  31386=>"001011000",
  31387=>"110001100",
  31388=>"001000010",
  31389=>"101001111",
  31390=>"000110000",
  31391=>"111001000",
  31392=>"010110010",
  31393=>"010100111",
  31394=>"111011001",
  31395=>"101011010",
  31396=>"100001001",
  31397=>"011011011",
  31398=>"111110000",
  31399=>"100110011",
  31400=>"000101110",
  31401=>"010110101",
  31402=>"110100100",
  31403=>"000000000",
  31404=>"011111010",
  31405=>"000110110",
  31406=>"010000011",
  31407=>"111100011",
  31408=>"100111011",
  31409=>"010010000",
  31410=>"101011001",
  31411=>"011010110",
  31412=>"010111000",
  31413=>"011111100",
  31414=>"101000001",
  31415=>"101100100",
  31416=>"100001000",
  31417=>"000101011",
  31418=>"101111000",
  31419=>"000000101",
  31420=>"010110011",
  31421=>"110111000",
  31422=>"000010000",
  31423=>"110001111",
  31424=>"101010010",
  31425=>"100101100",
  31426=>"111100110",
  31427=>"100000000",
  31428=>"110100100",
  31429=>"000001110",
  31430=>"111010000",
  31431=>"000100110",
  31432=>"010010100",
  31433=>"100011100",
  31434=>"101000110",
  31435=>"110111000",
  31436=>"001101101",
  31437=>"110111011",
  31438=>"100100110",
  31439=>"101101111",
  31440=>"111111111",
  31441=>"001010100",
  31442=>"000010011",
  31443=>"100101001",
  31444=>"110001100",
  31445=>"101000001",
  31446=>"101000101",
  31447=>"110000111",
  31448=>"100100111",
  31449=>"111001011",
  31450=>"001011101",
  31451=>"000011000",
  31452=>"111000011",
  31453=>"100010001",
  31454=>"110100011",
  31455=>"111000111",
  31456=>"011101111",
  31457=>"011011001",
  31458=>"000001100",
  31459=>"000000100",
  31460=>"100001101",
  31461=>"000011011",
  31462=>"010100001",
  31463=>"010101001",
  31464=>"100011101",
  31465=>"100010110",
  31466=>"010101010",
  31467=>"111010000",
  31468=>"101011001",
  31469=>"110111110",
  31470=>"100011101",
  31471=>"100000011",
  31472=>"000101111",
  31473=>"111111110",
  31474=>"111110111",
  31475=>"000001011",
  31476=>"011011110",
  31477=>"110101100",
  31478=>"111010000",
  31479=>"000101000",
  31480=>"001010011",
  31481=>"001111010",
  31482=>"100101100",
  31483=>"100011010",
  31484=>"000010101",
  31485=>"011101000",
  31486=>"000011100",
  31487=>"101011011",
  31488=>"011111111",
  31489=>"111111101",
  31490=>"101010111",
  31491=>"101000101",
  31492=>"010000100",
  31493=>"000010000",
  31494=>"010110010",
  31495=>"111001100",
  31496=>"110010000",
  31497=>"100110111",
  31498=>"010100010",
  31499=>"000000001",
  31500=>"011110110",
  31501=>"011111010",
  31502=>"011010111",
  31503=>"100110111",
  31504=>"101010000",
  31505=>"111111100",
  31506=>"110000010",
  31507=>"101000000",
  31508=>"001011110",
  31509=>"111110011",
  31510=>"111100000",
  31511=>"110001001",
  31512=>"000010001",
  31513=>"011100100",
  31514=>"111000100",
  31515=>"001101000",
  31516=>"011001111",
  31517=>"111111011",
  31518=>"110010110",
  31519=>"101111101",
  31520=>"001010110",
  31521=>"100001001",
  31522=>"010000000",
  31523=>"001101101",
  31524=>"001110100",
  31525=>"110010001",
  31526=>"010010011",
  31527=>"111100110",
  31528=>"100110011",
  31529=>"100111011",
  31530=>"110110011",
  31531=>"100010110",
  31532=>"110100101",
  31533=>"111101011",
  31534=>"011000000",
  31535=>"100000011",
  31536=>"110001010",
  31537=>"111111110",
  31538=>"100010000",
  31539=>"100111110",
  31540=>"110111111",
  31541=>"100100100",
  31542=>"010101010",
  31543=>"100001010",
  31544=>"011110100",
  31545=>"000011001",
  31546=>"111110010",
  31547=>"011001011",
  31548=>"110001010",
  31549=>"101101001",
  31550=>"011010000",
  31551=>"000011000",
  31552=>"110000000",
  31553=>"101111001",
  31554=>"001001001",
  31555=>"101001011",
  31556=>"100001110",
  31557=>"010101111",
  31558=>"100000011",
  31559=>"100111111",
  31560=>"000110110",
  31561=>"100101100",
  31562=>"110010001",
  31563=>"101110000",
  31564=>"101010010",
  31565=>"111011010",
  31566=>"000000110",
  31567=>"001011001",
  31568=>"010111001",
  31569=>"011001110",
  31570=>"001110110",
  31571=>"000010001",
  31572=>"010010100",
  31573=>"111110101",
  31574=>"101011001",
  31575=>"010001001",
  31576=>"101101101",
  31577=>"111010010",
  31578=>"110000000",
  31579=>"010001000",
  31580=>"110001011",
  31581=>"111111011",
  31582=>"010000111",
  31583=>"111111000",
  31584=>"111101000",
  31585=>"101000111",
  31586=>"101000111",
  31587=>"011111001",
  31588=>"101100011",
  31589=>"000001010",
  31590=>"111110111",
  31591=>"101010000",
  31592=>"011110011",
  31593=>"111111011",
  31594=>"100010000",
  31595=>"001110101",
  31596=>"000100011",
  31597=>"010111011",
  31598=>"101111011",
  31599=>"111011101",
  31600=>"011011111",
  31601=>"101001111",
  31602=>"100001000",
  31603=>"101000011",
  31604=>"000001011",
  31605=>"010001011",
  31606=>"010011000",
  31607=>"001110000",
  31608=>"010011110",
  31609=>"100111001",
  31610=>"101100101",
  31611=>"110111111",
  31612=>"110011011",
  31613=>"011101000",
  31614=>"110110001",
  31615=>"001101100",
  31616=>"001101001",
  31617=>"000001010",
  31618=>"011010010",
  31619=>"000011010",
  31620=>"111101101",
  31621=>"111001111",
  31622=>"000001000",
  31623=>"010110100",
  31624=>"000011010",
  31625=>"111111001",
  31626=>"000010101",
  31627=>"111101000",
  31628=>"010010000",
  31629=>"100111001",
  31630=>"000100101",
  31631=>"001111011",
  31632=>"000110111",
  31633=>"010101100",
  31634=>"100001000",
  31635=>"111100010",
  31636=>"111100101",
  31637=>"110110001",
  31638=>"110011010",
  31639=>"010101000",
  31640=>"110000001",
  31641=>"111010110",
  31642=>"011000011",
  31643=>"001110100",
  31644=>"100111000",
  31645=>"101111101",
  31646=>"011111111",
  31647=>"000111101",
  31648=>"000101000",
  31649=>"000001101",
  31650=>"110011100",
  31651=>"000000001",
  31652=>"110100001",
  31653=>"100110101",
  31654=>"100100101",
  31655=>"000000110",
  31656=>"101001111",
  31657=>"010000000",
  31658=>"111100010",
  31659=>"000000100",
  31660=>"111001010",
  31661=>"110010000",
  31662=>"001110110",
  31663=>"111110111",
  31664=>"101111010",
  31665=>"011001000",
  31666=>"100100010",
  31667=>"111101100",
  31668=>"000001111",
  31669=>"111000111",
  31670=>"111110001",
  31671=>"011000011",
  31672=>"000101101",
  31673=>"101000111",
  31674=>"001101111",
  31675=>"111001110",
  31676=>"101101011",
  31677=>"110111011",
  31678=>"100111001",
  31679=>"000000110",
  31680=>"100001000",
  31681=>"110010010",
  31682=>"001001011",
  31683=>"001110110",
  31684=>"001101111",
  31685=>"000111111",
  31686=>"110100010",
  31687=>"101110111",
  31688=>"000110011",
  31689=>"110000100",
  31690=>"011000001",
  31691=>"010101101",
  31692=>"100000111",
  31693=>"000110000",
  31694=>"111010110",
  31695=>"100111101",
  31696=>"110100011",
  31697=>"010101101",
  31698=>"010001110",
  31699=>"010000000",
  31700=>"001101100",
  31701=>"110000101",
  31702=>"000100001",
  31703=>"000111100",
  31704=>"100010000",
  31705=>"001011000",
  31706=>"110001001",
  31707=>"010000110",
  31708=>"001110011",
  31709=>"000110001",
  31710=>"100110100",
  31711=>"100000111",
  31712=>"101000111",
  31713=>"101011110",
  31714=>"101101111",
  31715=>"001111010",
  31716=>"000000000",
  31717=>"010010110",
  31718=>"111011001",
  31719=>"100010000",
  31720=>"000000001",
  31721=>"010101011",
  31722=>"001010100",
  31723=>"001011000",
  31724=>"000010101",
  31725=>"011111000",
  31726=>"001000011",
  31727=>"011010111",
  31728=>"101000010",
  31729=>"101001110",
  31730=>"001101100",
  31731=>"110110001",
  31732=>"111101100",
  31733=>"001110100",
  31734=>"011111100",
  31735=>"001110010",
  31736=>"011010011",
  31737=>"011100000",
  31738=>"100000100",
  31739=>"110001111",
  31740=>"111001111",
  31741=>"010001010",
  31742=>"101000001",
  31743=>"000101101",
  31744=>"111111011",
  31745=>"100111100",
  31746=>"011101101",
  31747=>"100101110",
  31748=>"111111011",
  31749=>"100000101",
  31750=>"101000110",
  31751=>"001010110",
  31752=>"111101110",
  31753=>"101111011",
  31754=>"011110001",
  31755=>"000110011",
  31756=>"000000011",
  31757=>"101011001",
  31758=>"010001110",
  31759=>"110101111",
  31760=>"111100000",
  31761=>"010110100",
  31762=>"100111100",
  31763=>"101000011",
  31764=>"101100100",
  31765=>"000110100",
  31766=>"101111001",
  31767=>"111100111",
  31768=>"111111010",
  31769=>"000100000",
  31770=>"011000100",
  31771=>"010110111",
  31772=>"101010000",
  31773=>"100010111",
  31774=>"010110010",
  31775=>"001000100",
  31776=>"011000001",
  31777=>"000000100",
  31778=>"111110110",
  31779=>"111110001",
  31780=>"001110011",
  31781=>"001000010",
  31782=>"111011100",
  31783=>"000101010",
  31784=>"010101110",
  31785=>"000111111",
  31786=>"111011100",
  31787=>"111001101",
  31788=>"000000000",
  31789=>"010000101",
  31790=>"110110110",
  31791=>"001111001",
  31792=>"010000100",
  31793=>"101101110",
  31794=>"011001100",
  31795=>"001011100",
  31796=>"111001100",
  31797=>"000001010",
  31798=>"010001000",
  31799=>"100110011",
  31800=>"111100011",
  31801=>"110111111",
  31802=>"000110111",
  31803=>"111000011",
  31804=>"000110100",
  31805=>"101010111",
  31806=>"110101001",
  31807=>"101000100",
  31808=>"111101000",
  31809=>"110001001",
  31810=>"010001000",
  31811=>"010011111",
  31812=>"100111000",
  31813=>"101101111",
  31814=>"111101010",
  31815=>"011101001",
  31816=>"100010010",
  31817=>"000000100",
  31818=>"001000100",
  31819=>"000000010",
  31820=>"000101001",
  31821=>"000000001",
  31822=>"000111010",
  31823=>"101011000",
  31824=>"001000010",
  31825=>"111110011",
  31826=>"101010100",
  31827=>"111111010",
  31828=>"101110110",
  31829=>"010010111",
  31830=>"110001010",
  31831=>"101011110",
  31832=>"011111111",
  31833=>"111100010",
  31834=>"111011111",
  31835=>"011000111",
  31836=>"100001110",
  31837=>"000111001",
  31838=>"010110100",
  31839=>"101100110",
  31840=>"110110110",
  31841=>"110010110",
  31842=>"100101111",
  31843=>"101111110",
  31844=>"001001111",
  31845=>"111111000",
  31846=>"111101001",
  31847=>"111001100",
  31848=>"111011110",
  31849=>"110100101",
  31850=>"000000101",
  31851=>"101111010",
  31852=>"101100001",
  31853=>"011110010",
  31854=>"111101110",
  31855=>"111111111",
  31856=>"111101100",
  31857=>"110011101",
  31858=>"010000010",
  31859=>"100100111",
  31860=>"110011001",
  31861=>"011011101",
  31862=>"000101111",
  31863=>"100100100",
  31864=>"101010101",
  31865=>"011000100",
  31866=>"110010001",
  31867=>"101111011",
  31868=>"000011100",
  31869=>"101010110",
  31870=>"111101001",
  31871=>"101100010",
  31872=>"100000010",
  31873=>"100110001",
  31874=>"101000001",
  31875=>"000101100",
  31876=>"000010000",
  31877=>"101001010",
  31878=>"000111001",
  31879=>"000101111",
  31880=>"110000111",
  31881=>"011110011",
  31882=>"000110000",
  31883=>"110011110",
  31884=>"011001101",
  31885=>"001001000",
  31886=>"101100000",
  31887=>"010011011",
  31888=>"111100101",
  31889=>"111000100",
  31890=>"001000010",
  31891=>"111101111",
  31892=>"010100001",
  31893=>"101101000",
  31894=>"111111100",
  31895=>"001000101",
  31896=>"100110101",
  31897=>"011101100",
  31898=>"010001000",
  31899=>"000000001",
  31900=>"100010111",
  31901=>"001110000",
  31902=>"000110010",
  31903=>"000011111",
  31904=>"010001111",
  31905=>"100000010",
  31906=>"100000110",
  31907=>"000011100",
  31908=>"010010010",
  31909=>"101010001",
  31910=>"010100100",
  31911=>"101110001",
  31912=>"011111011",
  31913=>"111100110",
  31914=>"001111000",
  31915=>"011100011",
  31916=>"000001110",
  31917=>"011101011",
  31918=>"110101001",
  31919=>"111100000",
  31920=>"001000110",
  31921=>"010110100",
  31922=>"101001011",
  31923=>"010000101",
  31924=>"010111101",
  31925=>"000111000",
  31926=>"111111111",
  31927=>"010101110",
  31928=>"111001111",
  31929=>"101100111",
  31930=>"111100111",
  31931=>"111110000",
  31932=>"011110110",
  31933=>"000001010",
  31934=>"011001101",
  31935=>"111001010",
  31936=>"011011000",
  31937=>"001011011",
  31938=>"010100000",
  31939=>"110001101",
  31940=>"111011001",
  31941=>"100111000",
  31942=>"001000011",
  31943=>"000111001",
  31944=>"011110011",
  31945=>"111010000",
  31946=>"101101101",
  31947=>"010111101",
  31948=>"000101100",
  31949=>"100101000",
  31950=>"011101110",
  31951=>"110001100",
  31952=>"010101001",
  31953=>"000100000",
  31954=>"000011101",
  31955=>"111111001",
  31956=>"110101011",
  31957=>"000000001",
  31958=>"000010001",
  31959=>"011000001",
  31960=>"101001111",
  31961=>"100110110",
  31962=>"001101101",
  31963=>"001110000",
  31964=>"100110100",
  31965=>"100110101",
  31966=>"011111111",
  31967=>"110010111",
  31968=>"100011010",
  31969=>"000110000",
  31970=>"001000000",
  31971=>"011100000",
  31972=>"010001110",
  31973=>"001011110",
  31974=>"010110011",
  31975=>"001101111",
  31976=>"101110011",
  31977=>"001000010",
  31978=>"010100010",
  31979=>"001011100",
  31980=>"000101001",
  31981=>"101000010",
  31982=>"001100011",
  31983=>"011110000",
  31984=>"111101001",
  31985=>"010000010",
  31986=>"101111001",
  31987=>"100001110",
  31988=>"000001100",
  31989=>"110000000",
  31990=>"111001000",
  31991=>"001111100",
  31992=>"111110111",
  31993=>"001111000",
  31994=>"110011100",
  31995=>"101011110",
  31996=>"100010000",
  31997=>"100100000",
  31998=>"010101011",
  31999=>"100001011",
  32000=>"110100100",
  32001=>"111010011",
  32002=>"111000111",
  32003=>"010111110",
  32004=>"001000000",
  32005=>"111011001",
  32006=>"011111100",
  32007=>"101000110",
  32008=>"111111110",
  32009=>"111101011",
  32010=>"101010110",
  32011=>"000111110",
  32012=>"000100000",
  32013=>"101001001",
  32014=>"100110000",
  32015=>"011111110",
  32016=>"110111000",
  32017=>"000011010",
  32018=>"111111101",
  32019=>"111111001",
  32020=>"111100001",
  32021=>"001010010",
  32022=>"110111001",
  32023=>"101110111",
  32024=>"100100010",
  32025=>"010011010",
  32026=>"010000100",
  32027=>"000001011",
  32028=>"000110111",
  32029=>"111100100",
  32030=>"000101101",
  32031=>"111101111",
  32032=>"010111110",
  32033=>"000011101",
  32034=>"000001100",
  32035=>"110010011",
  32036=>"010001001",
  32037=>"100000110",
  32038=>"111111111",
  32039=>"001100001",
  32040=>"000010000",
  32041=>"011111100",
  32042=>"000010111",
  32043=>"011101100",
  32044=>"000110001",
  32045=>"000111100",
  32046=>"000100111",
  32047=>"011100011",
  32048=>"011000011",
  32049=>"111110111",
  32050=>"000100110",
  32051=>"101101011",
  32052=>"111011011",
  32053=>"001100000",
  32054=>"010110001",
  32055=>"010010000",
  32056=>"101010101",
  32057=>"011011000",
  32058=>"111010100",
  32059=>"000010011",
  32060=>"000101111",
  32061=>"010000010",
  32062=>"110111110",
  32063=>"111000100",
  32064=>"100000111",
  32065=>"111100001",
  32066=>"010000111",
  32067=>"100000011",
  32068=>"100001100",
  32069=>"100110011",
  32070=>"110011101",
  32071=>"100001011",
  32072=>"110100110",
  32073=>"010101000",
  32074=>"111111000",
  32075=>"001010000",
  32076=>"000100101",
  32077=>"001000010",
  32078=>"100101111",
  32079=>"110011011",
  32080=>"011000110",
  32081=>"000100111",
  32082=>"000000000",
  32083=>"111110110",
  32084=>"101100011",
  32085=>"010011101",
  32086=>"100000110",
  32087=>"011100001",
  32088=>"101010110",
  32089=>"010000011",
  32090=>"010100010",
  32091=>"100010001",
  32092=>"001010101",
  32093=>"001101010",
  32094=>"001100011",
  32095=>"110011010",
  32096=>"010011101",
  32097=>"011010000",
  32098=>"010100101",
  32099=>"011010111",
  32100=>"100111001",
  32101=>"001000010",
  32102=>"001000110",
  32103=>"010000000",
  32104=>"011100111",
  32105=>"111111011",
  32106=>"001011010",
  32107=>"101110011",
  32108=>"000100111",
  32109=>"100111000",
  32110=>"100001110",
  32111=>"011111010",
  32112=>"110001011",
  32113=>"101000101",
  32114=>"100001101",
  32115=>"110001000",
  32116=>"101101111",
  32117=>"110010101",
  32118=>"011110111",
  32119=>"101100111",
  32120=>"010001011",
  32121=>"001101101",
  32122=>"001111111",
  32123=>"100000011",
  32124=>"001000000",
  32125=>"010000010",
  32126=>"110100111",
  32127=>"001111010",
  32128=>"100000110",
  32129=>"010010011",
  32130=>"100101000",
  32131=>"010000111",
  32132=>"100010000",
  32133=>"110111000",
  32134=>"111111000",
  32135=>"111010101",
  32136=>"001001000",
  32137=>"000000101",
  32138=>"010100011",
  32139=>"010001100",
  32140=>"111100111",
  32141=>"101110011",
  32142=>"011001001",
  32143=>"000111000",
  32144=>"101100101",
  32145=>"001100101",
  32146=>"110110110",
  32147=>"010010101",
  32148=>"011101011",
  32149=>"110101011",
  32150=>"100111011",
  32151=>"100000000",
  32152=>"101111011",
  32153=>"011110110",
  32154=>"110111111",
  32155=>"011010010",
  32156=>"111011110",
  32157=>"101101010",
  32158=>"110110111",
  32159=>"110001000",
  32160=>"011101101",
  32161=>"001000111",
  32162=>"010000100",
  32163=>"001101011",
  32164=>"010011101",
  32165=>"111100011",
  32166=>"000000001",
  32167=>"101110010",
  32168=>"111010100",
  32169=>"000100001",
  32170=>"111110100",
  32171=>"000101000",
  32172=>"101001000",
  32173=>"000110111",
  32174=>"000001011",
  32175=>"010101101",
  32176=>"010010010",
  32177=>"011011111",
  32178=>"001111000",
  32179=>"000011111",
  32180=>"110001001",
  32181=>"101111010",
  32182=>"001001100",
  32183=>"000001101",
  32184=>"100011110",
  32185=>"101010010",
  32186=>"111011001",
  32187=>"100110100",
  32188=>"000101010",
  32189=>"110111111",
  32190=>"010011110",
  32191=>"000110111",
  32192=>"110100100",
  32193=>"010000110",
  32194=>"011010010",
  32195=>"111001101",
  32196=>"100110111",
  32197=>"110000110",
  32198=>"011110000",
  32199=>"110110000",
  32200=>"011101011",
  32201=>"000010001",
  32202=>"111011011",
  32203=>"111110111",
  32204=>"111001011",
  32205=>"100011010",
  32206=>"000111001",
  32207=>"001010011",
  32208=>"000100100",
  32209=>"111010111",
  32210=>"111010101",
  32211=>"001100000",
  32212=>"001001000",
  32213=>"011000010",
  32214=>"000111100",
  32215=>"111010101",
  32216=>"001111100",
  32217=>"001110010",
  32218=>"100001001",
  32219=>"100011011",
  32220=>"101000001",
  32221=>"000100110",
  32222=>"111111011",
  32223=>"010011011",
  32224=>"001000110",
  32225=>"011111010",
  32226=>"000111010",
  32227=>"110101110",
  32228=>"101101100",
  32229=>"011111111",
  32230=>"010100000",
  32231=>"011011000",
  32232=>"101011000",
  32233=>"010100001",
  32234=>"010011010",
  32235=>"000000101",
  32236=>"110000010",
  32237=>"101101111",
  32238=>"010111111",
  32239=>"011001001",
  32240=>"110101101",
  32241=>"000111100",
  32242=>"001100111",
  32243=>"011100000",
  32244=>"111100111",
  32245=>"110110011",
  32246=>"101111000",
  32247=>"111011011",
  32248=>"111110101",
  32249=>"100011010",
  32250=>"001101001",
  32251=>"000001110",
  32252=>"101101011",
  32253=>"111001011",
  32254=>"101110100",
  32255=>"011000111",
  32256=>"010011010",
  32257=>"101100011",
  32258=>"111011010",
  32259=>"100101111",
  32260=>"101001111",
  32261=>"001111110",
  32262=>"011001010",
  32263=>"010110010",
  32264=>"010010100",
  32265=>"011011011",
  32266=>"111000010",
  32267=>"101110010",
  32268=>"010001000",
  32269=>"110110110",
  32270=>"011000011",
  32271=>"111110001",
  32272=>"100101100",
  32273=>"110110110",
  32274=>"011010101",
  32275=>"000100111",
  32276=>"101001000",
  32277=>"000100101",
  32278=>"100101100",
  32279=>"001010010",
  32280=>"010101011",
  32281=>"000100011",
  32282=>"011000001",
  32283=>"001100001",
  32284=>"001000010",
  32285=>"100000010",
  32286=>"001011110",
  32287=>"000100000",
  32288=>"101101100",
  32289=>"100010010",
  32290=>"111111110",
  32291=>"010101001",
  32292=>"111011010",
  32293=>"100111100",
  32294=>"001001100",
  32295=>"000100100",
  32296=>"100101111",
  32297=>"110001111",
  32298=>"100110000",
  32299=>"100111101",
  32300=>"001110111",
  32301=>"010010111",
  32302=>"110100001",
  32303=>"011100100",
  32304=>"011101110",
  32305=>"111011010",
  32306=>"100000100",
  32307=>"111110101",
  32308=>"100100101",
  32309=>"001011111",
  32310=>"111001101",
  32311=>"110100110",
  32312=>"111111101",
  32313=>"010101110",
  32314=>"000100000",
  32315=>"010110000",
  32316=>"101010100",
  32317=>"001100000",
  32318=>"000110110",
  32319=>"000000011",
  32320=>"111100110",
  32321=>"101100000",
  32322=>"111101110",
  32323=>"110111000",
  32324=>"010101100",
  32325=>"011001111",
  32326=>"000100001",
  32327=>"100010011",
  32328=>"111010110",
  32329=>"010000011",
  32330=>"110100001",
  32331=>"000000101",
  32332=>"101010110",
  32333=>"100001101",
  32334=>"111101000",
  32335=>"001011111",
  32336=>"000010011",
  32337=>"001101011",
  32338=>"101110011",
  32339=>"010110001",
  32340=>"100011010",
  32341=>"100010010",
  32342=>"100011011",
  32343=>"111010011",
  32344=>"000100100",
  32345=>"011101100",
  32346=>"111010111",
  32347=>"111110011",
  32348=>"000010000",
  32349=>"001000110",
  32350=>"000101000",
  32351=>"000111000",
  32352=>"011010101",
  32353=>"000001101",
  32354=>"001100110",
  32355=>"101111111",
  32356=>"111010100",
  32357=>"000000001",
  32358=>"000111010",
  32359=>"100101111",
  32360=>"110110001",
  32361=>"100001100",
  32362=>"000001010",
  32363=>"000111111",
  32364=>"111101100",
  32365=>"100001000",
  32366=>"000101010",
  32367=>"110110100",
  32368=>"100010110",
  32369=>"010101110",
  32370=>"011111010",
  32371=>"000001100",
  32372=>"011101001",
  32373=>"111101101",
  32374=>"001000010",
  32375=>"111111000",
  32376=>"000000000",
  32377=>"001011100",
  32378=>"101011100",
  32379=>"010001111",
  32380=>"110010111",
  32381=>"001001000",
  32382=>"101101010",
  32383=>"100100110",
  32384=>"001110011",
  32385=>"000101101",
  32386=>"100101010",
  32387=>"101110111",
  32388=>"011000000",
  32389=>"000111011",
  32390=>"001010010",
  32391=>"111011010",
  32392=>"000100000",
  32393=>"100100010",
  32394=>"100011100",
  32395=>"101111000",
  32396=>"100001110",
  32397=>"011010111",
  32398=>"011110111",
  32399=>"100111101",
  32400=>"010000000",
  32401=>"100010001",
  32402=>"001011010",
  32403=>"111001101",
  32404=>"010000011",
  32405=>"010000101",
  32406=>"010010000",
  32407=>"111011000",
  32408=>"101011101",
  32409=>"100111000",
  32410=>"101111110",
  32411=>"001111000",
  32412=>"010111010",
  32413=>"011101100",
  32414=>"000111110",
  32415=>"011011110",
  32416=>"011011100",
  32417=>"010101010",
  32418=>"101011110",
  32419=>"010000011",
  32420=>"100110010",
  32421=>"010001010",
  32422=>"100000100",
  32423=>"001000101",
  32424=>"011110110",
  32425=>"111011101",
  32426=>"100001010",
  32427=>"011010100",
  32428=>"111010110",
  32429=>"000101001",
  32430=>"100111010",
  32431=>"000110001",
  32432=>"111110100",
  32433=>"000001101",
  32434=>"000111000",
  32435=>"001111000",
  32436=>"011101101",
  32437=>"011000110",
  32438=>"110001001",
  32439=>"001001100",
  32440=>"000010110",
  32441=>"001011111",
  32442=>"010110100",
  32443=>"011001100",
  32444=>"100001111",
  32445=>"101001101",
  32446=>"101101111",
  32447=>"010100101",
  32448=>"000111011",
  32449=>"011101101",
  32450=>"000011001",
  32451=>"100110110",
  32452=>"010001000",
  32453=>"110001100",
  32454=>"111101111",
  32455=>"000000100",
  32456=>"101111111",
  32457=>"100111110",
  32458=>"101011111",
  32459=>"000110110",
  32460=>"101110000",
  32461=>"101110111",
  32462=>"000011100",
  32463=>"011110011",
  32464=>"010101000",
  32465=>"100100011",
  32466=>"100001011",
  32467=>"011000001",
  32468=>"111110101",
  32469=>"010100100",
  32470=>"101001111",
  32471=>"110001000",
  32472=>"100001011",
  32473=>"110001011",
  32474=>"101100110",
  32475=>"100111001",
  32476=>"100010111",
  32477=>"011111000",
  32478=>"000110100",
  32479=>"000010100",
  32480=>"000011111",
  32481=>"111101110",
  32482=>"111111110",
  32483=>"001110111",
  32484=>"110010110",
  32485=>"111100000",
  32486=>"000010101",
  32487=>"111110011",
  32488=>"001111011",
  32489=>"110101010",
  32490=>"111000100",
  32491=>"101110110",
  32492=>"011010111",
  32493=>"100111000",
  32494=>"101111110",
  32495=>"111111101",
  32496=>"000110010",
  32497=>"010111111",
  32498=>"000101011",
  32499=>"101000001",
  32500=>"110000101",
  32501=>"011101110",
  32502=>"111010011",
  32503=>"000000000",
  32504=>"111100011",
  32505=>"000000000",
  32506=>"110101001",
  32507=>"010000110",
  32508=>"001101010",
  32509=>"011010000",
  32510=>"111110111",
  32511=>"111101010",
  32512=>"011000110",
  32513=>"101010100",
  32514=>"001111001",
  32515=>"101111111",
  32516=>"000101001",
  32517=>"000100111",
  32518=>"000101100",
  32519=>"011001110",
  32520=>"110000010",
  32521=>"100101000",
  32522=>"110100000",
  32523=>"111101100",
  32524=>"001111010",
  32525=>"111110000",
  32526=>"011000111",
  32527=>"010111000",
  32528=>"000100000",
  32529=>"101001101",
  32530=>"001101110",
  32531=>"000111000",
  32532=>"000101101",
  32533=>"000011101",
  32534=>"001010001",
  32535=>"010011111",
  32536=>"001001111",
  32537=>"011000011",
  32538=>"110011000",
  32539=>"110101010",
  32540=>"000101110",
  32541=>"011100100",
  32542=>"100101000",
  32543=>"111011010",
  32544=>"011011111",
  32545=>"001010010",
  32546=>"011011111",
  32547=>"001000110",
  32548=>"110011100",
  32549=>"100010011",
  32550=>"111100111",
  32551=>"010100101",
  32552=>"010101110",
  32553=>"001011101",
  32554=>"001101011",
  32555=>"000010011",
  32556=>"101111110",
  32557=>"111111111",
  32558=>"001010110",
  32559=>"111110110",
  32560=>"111001110",
  32561=>"101000001",
  32562=>"111011010",
  32563=>"001010010",
  32564=>"011000000",
  32565=>"011111000",
  32566=>"100111010",
  32567=>"001110111",
  32568=>"110011000",
  32569=>"001111100",
  32570=>"000100100",
  32571=>"011111000",
  32572=>"001110110",
  32573=>"001110101",
  32574=>"011001001",
  32575=>"101100111",
  32576=>"100100010",
  32577=>"101010000",
  32578=>"011100001",
  32579=>"110110100",
  32580=>"010001111",
  32581=>"010011110",
  32582=>"100110101",
  32583=>"110001100",
  32584=>"111111011",
  32585=>"110000110",
  32586=>"111100010",
  32587=>"111000000",
  32588=>"101101001",
  32589=>"011100000",
  32590=>"100001100",
  32591=>"001000010",
  32592=>"101100111",
  32593=>"010001001",
  32594=>"000101010",
  32595=>"010010101",
  32596=>"000101001",
  32597=>"001111000",
  32598=>"001001110",
  32599=>"011011011",
  32600=>"010111000",
  32601=>"111111011",
  32602=>"011010010",
  32603=>"100101101",
  32604=>"111000001",
  32605=>"001000110",
  32606=>"110110101",
  32607=>"101010101",
  32608=>"110000000",
  32609=>"001110111",
  32610=>"101111011",
  32611=>"111011001",
  32612=>"010101010",
  32613=>"000110110",
  32614=>"010101111",
  32615=>"010001011",
  32616=>"000100100",
  32617=>"011010011",
  32618=>"000100010",
  32619=>"100100001",
  32620=>"110110110",
  32621=>"101100000",
  32622=>"000100101",
  32623=>"001011100",
  32624=>"110111011",
  32625=>"010001010",
  32626=>"110001000",
  32627=>"110000100",
  32628=>"010001010",
  32629=>"011010011",
  32630=>"010001111",
  32631=>"000000011",
  32632=>"010001000",
  32633=>"111100101",
  32634=>"111111100",
  32635=>"111000001",
  32636=>"111101001",
  32637=>"100101011",
  32638=>"000001111",
  32639=>"010111111",
  32640=>"111010000",
  32641=>"010010011",
  32642=>"000000101",
  32643=>"000010111",
  32644=>"101010010",
  32645=>"100101011",
  32646=>"000010110",
  32647=>"010011110",
  32648=>"100110111",
  32649=>"111000001",
  32650=>"111100000",
  32651=>"001011000",
  32652=>"000011010",
  32653=>"011000101",
  32654=>"011000011",
  32655=>"100110101",
  32656=>"101100000",
  32657=>"010101100",
  32658=>"100000011",
  32659=>"011001110",
  32660=>"111000111",
  32661=>"101010010",
  32662=>"001000000",
  32663=>"110011111",
  32664=>"101011010",
  32665=>"000110011",
  32666=>"010111110",
  32667=>"101100010",
  32668=>"110010111",
  32669=>"101001001",
  32670=>"000101110",
  32671=>"010010111",
  32672=>"101101010",
  32673=>"001110000",
  32674=>"010111001",
  32675=>"000101000",
  32676=>"011110101",
  32677=>"111000011",
  32678=>"011100011",
  32679=>"101100110",
  32680=>"100101001",
  32681=>"111011011",
  32682=>"101111011",
  32683=>"100110011",
  32684=>"101111101",
  32685=>"111011101",
  32686=>"010100000",
  32687=>"100101101",
  32688=>"001111011",
  32689=>"010111000",
  32690=>"010010001",
  32691=>"110010010",
  32692=>"000100000",
  32693=>"101110101",
  32694=>"000001011",
  32695=>"000110000",
  32696=>"101100101",
  32697=>"000100110",
  32698=>"110000111",
  32699=>"010100101",
  32700=>"001001000",
  32701=>"000111000",
  32702=>"000000001",
  32703=>"001101001",
  32704=>"011111111",
  32705=>"000110101",
  32706=>"001001110",
  32707=>"000101111",
  32708=>"101110101",
  32709=>"011100101",
  32710=>"010111010",
  32711=>"011010001",
  32712=>"010111100",
  32713=>"010101001",
  32714=>"001001000",
  32715=>"011110111",
  32716=>"000110101",
  32717=>"100100111",
  32718=>"111101111",
  32719=>"000111000",
  32720=>"000111000",
  32721=>"100111000",
  32722=>"000011110",
  32723=>"011010000",
  32724=>"111110101",
  32725=>"010111011",
  32726=>"110000011",
  32727=>"001000101",
  32728=>"010111010",
  32729=>"011101101",
  32730=>"000001110",
  32731=>"110111010",
  32732=>"111000110",
  32733=>"011110011",
  32734=>"111001101",
  32735=>"000000100",
  32736=>"011001011",
  32737=>"000001000",
  32738=>"100001011",
  32739=>"110110010",
  32740=>"000110101",
  32741=>"111101110",
  32742=>"011000111",
  32743=>"111100111",
  32744=>"010111011",
  32745=>"100110111",
  32746=>"101111010",
  32747=>"000010011",
  32748=>"010101001",
  32749=>"111010000",
  32750=>"111000000",
  32751=>"011111010",
  32752=>"100111000",
  32753=>"101101101",
  32754=>"101011111",
  32755=>"010110110",
  32756=>"111011001",
  32757=>"111110011",
  32758=>"010101110",
  32759=>"001001010",
  32760=>"100010000",
  32761=>"111111111",
  32762=>"111010010",
  32763=>"010000011",
  32764=>"111101011",
  32765=>"000101011",
  32766=>"010101110",
  32767=>"011100111",
  32768=>"000101001",
  32769=>"101101011",
  32770=>"110101110",
  32771=>"001110110",
  32772=>"110010110",
  32773=>"100000100",
  32774=>"101100101",
  32775=>"111100111",
  32776=>"011101100",
  32777=>"010001010",
  32778=>"000011110",
  32779=>"000110000",
  32780=>"001001111",
  32781=>"001110100",
  32782=>"111100111",
  32783=>"101000100",
  32784=>"011100111",
  32785=>"110100000",
  32786=>"101001010",
  32787=>"000100001",
  32788=>"000000000",
  32789=>"011010111",
  32790=>"100110000",
  32791=>"000000101",
  32792=>"010110011",
  32793=>"011010011",
  32794=>"111110011",
  32795=>"000011101",
  32796=>"011000101",
  32797=>"110100011",
  32798=>"010001000",
  32799=>"000101011",
  32800=>"110111111",
  32801=>"001111011",
  32802=>"101001000",
  32803=>"010101110",
  32804=>"110000111",
  32805=>"001011100",
  32806=>"001010001",
  32807=>"101011001",
  32808=>"001011111",
  32809=>"111100110",
  32810=>"011110111",
  32811=>"110000000",
  32812=>"001110111",
  32813=>"000001101",
  32814=>"100100010",
  32815=>"111101111",
  32816=>"011110111",
  32817=>"100100001",
  32818=>"000110010",
  32819=>"001100110",
  32820=>"110111101",
  32821=>"001011011",
  32822=>"010000011",
  32823=>"011111100",
  32824=>"001000100",
  32825=>"111111011",
  32826=>"111000000",
  32827=>"100100011",
  32828=>"110010001",
  32829=>"100110101",
  32830=>"101011000",
  32831=>"100011100",
  32832=>"101011101",
  32833=>"000010000",
  32834=>"101001011",
  32835=>"001100011",
  32836=>"011011011",
  32837=>"001110110",
  32838=>"101100111",
  32839=>"000001000",
  32840=>"100000110",
  32841=>"011001010",
  32842=>"001001010",
  32843=>"010111101",
  32844=>"001000001",
  32845=>"111111111",
  32846=>"100100000",
  32847=>"000000110",
  32848=>"111001000",
  32849=>"101010011",
  32850=>"001000001",
  32851=>"000111000",
  32852=>"011110100",
  32853=>"001011000",
  32854=>"010101110",
  32855=>"001111111",
  32856=>"111110010",
  32857=>"000111111",
  32858=>"001111001",
  32859=>"001011010",
  32860=>"010101111",
  32861=>"110100000",
  32862=>"111011001",
  32863=>"000010001",
  32864=>"011100111",
  32865=>"001000000",
  32866=>"010011000",
  32867=>"000100001",
  32868=>"111010000",
  32869=>"111101010",
  32870=>"110100011",
  32871=>"101110010",
  32872=>"000110111",
  32873=>"010111001",
  32874=>"011101111",
  32875=>"001111000",
  32876=>"111000111",
  32877=>"010011111",
  32878=>"101011100",
  32879=>"101110100",
  32880=>"010000001",
  32881=>"111101000",
  32882=>"100000110",
  32883=>"110011101",
  32884=>"100111011",
  32885=>"010001101",
  32886=>"001011011",
  32887=>"001001001",
  32888=>"010111011",
  32889=>"111110010",
  32890=>"110001100",
  32891=>"100000000",
  32892=>"000001111",
  32893=>"100010000",
  32894=>"100110001",
  32895=>"100110101",
  32896=>"100000010",
  32897=>"011011011",
  32898=>"111100101",
  32899=>"000011111",
  32900=>"101000000",
  32901=>"001000111",
  32902=>"011110000",
  32903=>"111110111",
  32904=>"101010101",
  32905=>"001000001",
  32906=>"000001001",
  32907=>"010111111",
  32908=>"111111110",
  32909=>"111010101",
  32910=>"100011101",
  32911=>"110101011",
  32912=>"000110000",
  32913=>"110011110",
  32914=>"000000111",
  32915=>"111001100",
  32916=>"111101111",
  32917=>"000000000",
  32918=>"000010100",
  32919=>"001101111",
  32920=>"010101010",
  32921=>"100010110",
  32922=>"100011011",
  32923=>"101111111",
  32924=>"110111010",
  32925=>"101100101",
  32926=>"000000000",
  32927=>"100110101",
  32928=>"010001011",
  32929=>"010010001",
  32930=>"010110100",
  32931=>"010110010",
  32932=>"111100000",
  32933=>"001000001",
  32934=>"110101011",
  32935=>"000100000",
  32936=>"000101000",
  32937=>"110110000",
  32938=>"100110010",
  32939=>"001011100",
  32940=>"011111111",
  32941=>"110010000",
  32942=>"110110001",
  32943=>"110000111",
  32944=>"000000001",
  32945=>"100111111",
  32946=>"101101101",
  32947=>"010000001",
  32948=>"011100100",
  32949=>"001001011",
  32950=>"101101111",
  32951=>"110011110",
  32952=>"001001111",
  32953=>"101110111",
  32954=>"000000100",
  32955=>"101000101",
  32956=>"101001010",
  32957=>"110001111",
  32958=>"000001101",
  32959=>"110110000",
  32960=>"110011101",
  32961=>"100001011",
  32962=>"101101100",
  32963=>"010111111",
  32964=>"111000010",
  32965=>"100010111",
  32966=>"001111000",
  32967=>"100111010",
  32968=>"101001111",
  32969=>"100110001",
  32970=>"100000111",
  32971=>"001011100",
  32972=>"101111000",
  32973=>"011011011",
  32974=>"001000000",
  32975=>"100010110",
  32976=>"101001100",
  32977=>"110100010",
  32978=>"001111101",
  32979=>"110010011",
  32980=>"010100101",
  32981=>"111001011",
  32982=>"111001100",
  32983=>"110101010",
  32984=>"101000000",
  32985=>"100100011",
  32986=>"000010000",
  32987=>"011110000",
  32988=>"010101110",
  32989=>"001000100",
  32990=>"110001111",
  32991=>"010001101",
  32992=>"111101110",
  32993=>"101011111",
  32994=>"011010001",
  32995=>"111101010",
  32996=>"010111010",
  32997=>"000110100",
  32998=>"010100110",
  32999=>"001000111",
  33000=>"011101011",
  33001=>"000011000",
  33002=>"010100011",
  33003=>"000010100",
  33004=>"100101110",
  33005=>"101111101",
  33006=>"000111100",
  33007=>"000010000",
  33008=>"011001111",
  33009=>"010000010",
  33010=>"010010000",
  33011=>"011111001",
  33012=>"100000110",
  33013=>"010001111",
  33014=>"100001000",
  33015=>"000000010",
  33016=>"101000011",
  33017=>"000000010",
  33018=>"110001110",
  33019=>"001000100",
  33020=>"010101000",
  33021=>"101101000",
  33022=>"011000100",
  33023=>"100001010",
  33024=>"000011000",
  33025=>"011011011",
  33026=>"110000001",
  33027=>"010001110",
  33028=>"001101110",
  33029=>"100011011",
  33030=>"100000110",
  33031=>"000100101",
  33032=>"001101010",
  33033=>"110101001",
  33034=>"000111010",
  33035=>"000011010",
  33036=>"010011101",
  33037=>"000110010",
  33038=>"011000000",
  33039=>"111001100",
  33040=>"011111111",
  33041=>"000010010",
  33042=>"110110110",
  33043=>"100110000",
  33044=>"001000011",
  33045=>"010100111",
  33046=>"100011111",
  33047=>"101111110",
  33048=>"100000001",
  33049=>"011010110",
  33050=>"111010001",
  33051=>"100111110",
  33052=>"111111000",
  33053=>"010011010",
  33054=>"010110010",
  33055=>"000001111",
  33056=>"001101101",
  33057=>"000110010",
  33058=>"000111111",
  33059=>"011001000",
  33060=>"101011111",
  33061=>"110110101",
  33062=>"000010110",
  33063=>"101111000",
  33064=>"001100000",
  33065=>"001101010",
  33066=>"110110100",
  33067=>"011100101",
  33068=>"101000100",
  33069=>"011101011",
  33070=>"000110111",
  33071=>"111000001",
  33072=>"011100101",
  33073=>"000001001",
  33074=>"100100001",
  33075=>"011101110",
  33076=>"010000100",
  33077=>"101010100",
  33078=>"010100000",
  33079=>"010110000",
  33080=>"100001101",
  33081=>"110111000",
  33082=>"110011011",
  33083=>"110100000",
  33084=>"100000110",
  33085=>"000101101",
  33086=>"111100010",
  33087=>"001100010",
  33088=>"000110001",
  33089=>"111100000",
  33090=>"001110110",
  33091=>"101100111",
  33092=>"010111111",
  33093=>"110100111",
  33094=>"100001101",
  33095=>"101101101",
  33096=>"000010110",
  33097=>"100001100",
  33098=>"100100111",
  33099=>"000000000",
  33100=>"101101011",
  33101=>"100101101",
  33102=>"011000000",
  33103=>"110000100",
  33104=>"111000001",
  33105=>"011010110",
  33106=>"000100101",
  33107=>"101010110",
  33108=>"010111011",
  33109=>"111100110",
  33110=>"100101100",
  33111=>"000101100",
  33112=>"110000000",
  33113=>"011000100",
  33114=>"000110111",
  33115=>"001100100",
  33116=>"011011000",
  33117=>"001011101",
  33118=>"110001010",
  33119=>"001000111",
  33120=>"101000001",
  33121=>"001001111",
  33122=>"010101000",
  33123=>"000000001",
  33124=>"010110100",
  33125=>"011001011",
  33126=>"010101001",
  33127=>"000000001",
  33128=>"010111010",
  33129=>"001100001",
  33130=>"100011001",
  33131=>"100101001",
  33132=>"001010011",
  33133=>"110101001",
  33134=>"101011110",
  33135=>"100001010",
  33136=>"011111010",
  33137=>"111111111",
  33138=>"000010101",
  33139=>"001101101",
  33140=>"100000010",
  33141=>"001101011",
  33142=>"111100011",
  33143=>"011100001",
  33144=>"101111111",
  33145=>"110000010",
  33146=>"010101000",
  33147=>"110000101",
  33148=>"111000111",
  33149=>"111111100",
  33150=>"011000101",
  33151=>"101101000",
  33152=>"001000110",
  33153=>"001110001",
  33154=>"010111101",
  33155=>"111100100",
  33156=>"110000110",
  33157=>"100110101",
  33158=>"111010100",
  33159=>"010110111",
  33160=>"101001110",
  33161=>"000100101",
  33162=>"110111100",
  33163=>"110010000",
  33164=>"100111011",
  33165=>"111001001",
  33166=>"010110111",
  33167=>"101010010",
  33168=>"110101010",
  33169=>"000100011",
  33170=>"001101110",
  33171=>"010111010",
  33172=>"010000101",
  33173=>"101100001",
  33174=>"100010110",
  33175=>"111111011",
  33176=>"001000100",
  33177=>"001100011",
  33178=>"100011111",
  33179=>"011000011",
  33180=>"011110110",
  33181=>"110001110",
  33182=>"111111010",
  33183=>"101011010",
  33184=>"000100000",
  33185=>"100110000",
  33186=>"111000101",
  33187=>"111111111",
  33188=>"111001011",
  33189=>"000111001",
  33190=>"001001111",
  33191=>"101000000",
  33192=>"110101101",
  33193=>"100110011",
  33194=>"110100011",
  33195=>"111111101",
  33196=>"001010110",
  33197=>"101001001",
  33198=>"101010110",
  33199=>"010000010",
  33200=>"001000001",
  33201=>"011000100",
  33202=>"000011000",
  33203=>"100011111",
  33204=>"101100101",
  33205=>"010100101",
  33206=>"100100000",
  33207=>"001001011",
  33208=>"100110100",
  33209=>"100101100",
  33210=>"001001001",
  33211=>"100101100",
  33212=>"001101001",
  33213=>"011000111",
  33214=>"011100010",
  33215=>"011111011",
  33216=>"111011100",
  33217=>"011100101",
  33218=>"000100001",
  33219=>"001001101",
  33220=>"100100000",
  33221=>"101010001",
  33222=>"011110010",
  33223=>"110010111",
  33224=>"011001100",
  33225=>"001001001",
  33226=>"010000101",
  33227=>"000100101",
  33228=>"001111110",
  33229=>"010101111",
  33230=>"000100000",
  33231=>"011000101",
  33232=>"111011001",
  33233=>"000110101",
  33234=>"111001100",
  33235=>"000101001",
  33236=>"110111110",
  33237=>"011000110",
  33238=>"111111100",
  33239=>"100001001",
  33240=>"100001100",
  33241=>"101000101",
  33242=>"100111000",
  33243=>"011101001",
  33244=>"001001000",
  33245=>"001001101",
  33246=>"001110011",
  33247=>"010000100",
  33248=>"101010110",
  33249=>"000100000",
  33250=>"110100110",
  33251=>"011101101",
  33252=>"111001101",
  33253=>"110011101",
  33254=>"010000111",
  33255=>"101011010",
  33256=>"100000111",
  33257=>"010100110",
  33258=>"001111100",
  33259=>"000111001",
  33260=>"011010010",
  33261=>"010010011",
  33262=>"000111110",
  33263=>"110111001",
  33264=>"001110000",
  33265=>"001010000",
  33266=>"001011100",
  33267=>"000001100",
  33268=>"001000001",
  33269=>"010110001",
  33270=>"111000101",
  33271=>"101001110",
  33272=>"000110001",
  33273=>"011011000",
  33274=>"001110011",
  33275=>"011011110",
  33276=>"111101010",
  33277=>"000110111",
  33278=>"111000111",
  33279=>"011110010",
  33280=>"000101000",
  33281=>"011001010",
  33282=>"000000010",
  33283=>"001011100",
  33284=>"111001011",
  33285=>"110000101",
  33286=>"001001011",
  33287=>"000101101",
  33288=>"101001000",
  33289=>"110101111",
  33290=>"110001011",
  33291=>"011100000",
  33292=>"000010000",
  33293=>"101111101",
  33294=>"101010001",
  33295=>"011010111",
  33296=>"011111111",
  33297=>"000101100",
  33298=>"111000001",
  33299=>"000000010",
  33300=>"101100100",
  33301=>"011110000",
  33302=>"001000000",
  33303=>"100000101",
  33304=>"101111100",
  33305=>"101001000",
  33306=>"011010111",
  33307=>"001101010",
  33308=>"001000000",
  33309=>"101001010",
  33310=>"110010000",
  33311=>"111101011",
  33312=>"111000111",
  33313=>"000111100",
  33314=>"000100011",
  33315=>"100011010",
  33316=>"110110100",
  33317=>"001101100",
  33318=>"001101111",
  33319=>"001000000",
  33320=>"101010000",
  33321=>"100101101",
  33322=>"111001101",
  33323=>"011010000",
  33324=>"000111010",
  33325=>"110101000",
  33326=>"001110100",
  33327=>"000010000",
  33328=>"110011000",
  33329=>"011101010",
  33330=>"111110111",
  33331=>"000001000",
  33332=>"101110100",
  33333=>"001100110",
  33334=>"110100011",
  33335=>"010101000",
  33336=>"111000000",
  33337=>"111100101",
  33338=>"000001011",
  33339=>"101011100",
  33340=>"111011100",
  33341=>"000001110",
  33342=>"010000011",
  33343=>"110010111",
  33344=>"010100111",
  33345=>"100110001",
  33346=>"100110001",
  33347=>"010000011",
  33348=>"011011111",
  33349=>"111011101",
  33350=>"101111010",
  33351=>"010101011",
  33352=>"001000001",
  33353=>"111011111",
  33354=>"100100101",
  33355=>"100001101",
  33356=>"100110011",
  33357=>"110001101",
  33358=>"010111010",
  33359=>"110110001",
  33360=>"111001110",
  33361=>"000001000",
  33362=>"100000001",
  33363=>"001011000",
  33364=>"011000011",
  33365=>"001011110",
  33366=>"100111101",
  33367=>"011111010",
  33368=>"101001111",
  33369=>"101101001",
  33370=>"010101011",
  33371=>"100000100",
  33372=>"100001011",
  33373=>"101001011",
  33374=>"100101100",
  33375=>"001100010",
  33376=>"100100001",
  33377=>"011111101",
  33378=>"100100100",
  33379=>"100000010",
  33380=>"100001010",
  33381=>"100101100",
  33382=>"001110101",
  33383=>"011100100",
  33384=>"010100000",
  33385=>"110000100",
  33386=>"011001110",
  33387=>"101011100",
  33388=>"110000010",
  33389=>"011101001",
  33390=>"000010100",
  33391=>"100000101",
  33392=>"111000110",
  33393=>"011111101",
  33394=>"000000100",
  33395=>"011001111",
  33396=>"001000011",
  33397=>"000010011",
  33398=>"100010100",
  33399=>"010111101",
  33400=>"111110101",
  33401=>"011100000",
  33402=>"100000000",
  33403=>"000110001",
  33404=>"001010101",
  33405=>"100000101",
  33406=>"100100000",
  33407=>"000011000",
  33408=>"110011011",
  33409=>"000000000",
  33410=>"001101001",
  33411=>"111111100",
  33412=>"101001010",
  33413=>"110100000",
  33414=>"000011110",
  33415=>"100101000",
  33416=>"011001000",
  33417=>"111010110",
  33418=>"111111001",
  33419=>"010011000",
  33420=>"111110101",
  33421=>"011001101",
  33422=>"010111110",
  33423=>"110110001",
  33424=>"011011010",
  33425=>"110101100",
  33426=>"110011111",
  33427=>"111101010",
  33428=>"010011100",
  33429=>"000010101",
  33430=>"000000000",
  33431=>"110111100",
  33432=>"111111101",
  33433=>"001011110",
  33434=>"100001101",
  33435=>"011001101",
  33436=>"111000001",
  33437=>"001001010",
  33438=>"000100111",
  33439=>"001101111",
  33440=>"101101111",
  33441=>"000001100",
  33442=>"001110001",
  33443=>"110110000",
  33444=>"111011000",
  33445=>"011011011",
  33446=>"101011000",
  33447=>"000100101",
  33448=>"111101011",
  33449=>"000000100",
  33450=>"101110111",
  33451=>"011001010",
  33452=>"100010100",
  33453=>"001100000",
  33454=>"101110000",
  33455=>"001011000",
  33456=>"101010000",
  33457=>"000011011",
  33458=>"100000100",
  33459=>"111011101",
  33460=>"100001011",
  33461=>"001001011",
  33462=>"110100000",
  33463=>"000111100",
  33464=>"010000101",
  33465=>"010000011",
  33466=>"001100000",
  33467=>"100011011",
  33468=>"100011111",
  33469=>"100010011",
  33470=>"011010011",
  33471=>"011011011",
  33472=>"100000111",
  33473=>"000001011",
  33474=>"100111010",
  33475=>"011010000",
  33476=>"000000011",
  33477=>"000111010",
  33478=>"011111110",
  33479=>"110001100",
  33480=>"110111111",
  33481=>"001001110",
  33482=>"001111101",
  33483=>"001100100",
  33484=>"000000001",
  33485=>"001110100",
  33486=>"000110111",
  33487=>"100100000",
  33488=>"111110111",
  33489=>"110111110",
  33490=>"001110111",
  33491=>"111001110",
  33492=>"001010010",
  33493=>"100000100",
  33494=>"001101001",
  33495=>"101101101",
  33496=>"010011110",
  33497=>"011100011",
  33498=>"100110000",
  33499=>"101001101",
  33500=>"101000001",
  33501=>"000000000",
  33502=>"111100000",
  33503=>"001101000",
  33504=>"111011110",
  33505=>"010010010",
  33506=>"001100100",
  33507=>"101001100",
  33508=>"100100011",
  33509=>"010100101",
  33510=>"111000000",
  33511=>"011101110",
  33512=>"010001100",
  33513=>"110111100",
  33514=>"001111110",
  33515=>"001011001",
  33516=>"000000011",
  33517=>"100111110",
  33518=>"001110001",
  33519=>"110110100",
  33520=>"001110111",
  33521=>"101011000",
  33522=>"111000100",
  33523=>"010111010",
  33524=>"110000001",
  33525=>"000100000",
  33526=>"000110110",
  33527=>"101010110",
  33528=>"000000010",
  33529=>"001000101",
  33530=>"000100000",
  33531=>"011100101",
  33532=>"000110111",
  33533=>"100011101",
  33534=>"101111101",
  33535=>"100000110",
  33536=>"100110100",
  33537=>"101011100",
  33538=>"101101110",
  33539=>"000001010",
  33540=>"011001100",
  33541=>"100000101",
  33542=>"100010000",
  33543=>"010100001",
  33544=>"000010011",
  33545=>"111111111",
  33546=>"001101100",
  33547=>"011101101",
  33548=>"000100110",
  33549=>"111110001",
  33550=>"001011101",
  33551=>"011101111",
  33552=>"111110110",
  33553=>"101101100",
  33554=>"010001001",
  33555=>"110100011",
  33556=>"101001100",
  33557=>"110100100",
  33558=>"000101011",
  33559=>"001010110",
  33560=>"111101011",
  33561=>"001110100",
  33562=>"000001001",
  33563=>"001100101",
  33564=>"100011000",
  33565=>"010010011",
  33566=>"100111110",
  33567=>"100001010",
  33568=>"111101010",
  33569=>"111000111",
  33570=>"111100001",
  33571=>"010100011",
  33572=>"111000111",
  33573=>"110111111",
  33574=>"110111000",
  33575=>"010110111",
  33576=>"111001110",
  33577=>"001001000",
  33578=>"000110001",
  33579=>"101100111",
  33580=>"000010001",
  33581=>"111110111",
  33582=>"100101111",
  33583=>"000111001",
  33584=>"111010001",
  33585=>"000001001",
  33586=>"101110001",
  33587=>"111000110",
  33588=>"001011010",
  33589=>"000000010",
  33590=>"010000101",
  33591=>"001010101",
  33592=>"110100000",
  33593=>"111010110",
  33594=>"010010011",
  33595=>"010100000",
  33596=>"110101011",
  33597=>"001010011",
  33598=>"100100101",
  33599=>"010111101",
  33600=>"000101010",
  33601=>"101010100",
  33602=>"010111111",
  33603=>"101101100",
  33604=>"011001011",
  33605=>"000111010",
  33606=>"101001010",
  33607=>"011001011",
  33608=>"100101110",
  33609=>"011110100",
  33610=>"011110101",
  33611=>"000110001",
  33612=>"111001011",
  33613=>"000111010",
  33614=>"000100000",
  33615=>"001101100",
  33616=>"000100100",
  33617=>"101010111",
  33618=>"010001000",
  33619=>"011010011",
  33620=>"000101101",
  33621=>"010000000",
  33622=>"110010011",
  33623=>"110001101",
  33624=>"010101001",
  33625=>"000100010",
  33626=>"010000111",
  33627=>"101111101",
  33628=>"110111011",
  33629=>"100000011",
  33630=>"101101110",
  33631=>"111001111",
  33632=>"110110011",
  33633=>"101000100",
  33634=>"100100011",
  33635=>"100000110",
  33636=>"111100010",
  33637=>"011110101",
  33638=>"011001000",
  33639=>"111111110",
  33640=>"100110111",
  33641=>"111101011",
  33642=>"011011011",
  33643=>"001011111",
  33644=>"111001011",
  33645=>"010110101",
  33646=>"100000111",
  33647=>"100111010",
  33648=>"110011110",
  33649=>"111100111",
  33650=>"110011100",
  33651=>"101000110",
  33652=>"000011010",
  33653=>"000101111",
  33654=>"111001111",
  33655=>"111011001",
  33656=>"000111111",
  33657=>"010110010",
  33658=>"011010110",
  33659=>"100001010",
  33660=>"000001101",
  33661=>"111010001",
  33662=>"101111110",
  33663=>"010110100",
  33664=>"101000010",
  33665=>"100010100",
  33666=>"010100110",
  33667=>"111000110",
  33668=>"001010110",
  33669=>"100011101",
  33670=>"011000011",
  33671=>"011101110",
  33672=>"101000001",
  33673=>"010011101",
  33674=>"011101010",
  33675=>"101100100",
  33676=>"000010010",
  33677=>"110010010",
  33678=>"000101101",
  33679=>"100101000",
  33680=>"100110111",
  33681=>"100010011",
  33682=>"100010101",
  33683=>"111100010",
  33684=>"001010101",
  33685=>"101100111",
  33686=>"111000001",
  33687=>"100001101",
  33688=>"011011000",
  33689=>"011010001",
  33690=>"011001000",
  33691=>"000101110",
  33692=>"001001011",
  33693=>"111101001",
  33694=>"010010111",
  33695=>"000111000",
  33696=>"011111101",
  33697=>"011011100",
  33698=>"010110100",
  33699=>"010010011",
  33700=>"100011001",
  33701=>"111011010",
  33702=>"100111001",
  33703=>"000000000",
  33704=>"110001011",
  33705=>"101010001",
  33706=>"011110110",
  33707=>"001010101",
  33708=>"011110011",
  33709=>"101000010",
  33710=>"110110000",
  33711=>"011000000",
  33712=>"010000101",
  33713=>"011000011",
  33714=>"110101110",
  33715=>"001000110",
  33716=>"011110000",
  33717=>"010010000",
  33718=>"000100011",
  33719=>"000111000",
  33720=>"100010011",
  33721=>"010100111",
  33722=>"001110100",
  33723=>"010101100",
  33724=>"110100010",
  33725=>"010010001",
  33726=>"111000101",
  33727=>"011001001",
  33728=>"101110111",
  33729=>"101111010",
  33730=>"010101100",
  33731=>"010011110",
  33732=>"100100001",
  33733=>"001011101",
  33734=>"010101011",
  33735=>"100100011",
  33736=>"001001010",
  33737=>"101011001",
  33738=>"010101001",
  33739=>"101011001",
  33740=>"001101000",
  33741=>"010001110",
  33742=>"000111101",
  33743=>"101000000",
  33744=>"001001111",
  33745=>"101001001",
  33746=>"111001010",
  33747=>"000100000",
  33748=>"001100101",
  33749=>"111011110",
  33750=>"110000111",
  33751=>"001000000",
  33752=>"001000001",
  33753=>"100000001",
  33754=>"111000001",
  33755=>"010100100",
  33756=>"101001110",
  33757=>"000000101",
  33758=>"101111101",
  33759=>"010110001",
  33760=>"011001101",
  33761=>"000101010",
  33762=>"101101110",
  33763=>"011100011",
  33764=>"000000010",
  33765=>"000000010",
  33766=>"101000101",
  33767=>"000010001",
  33768=>"000100110",
  33769=>"010111011",
  33770=>"000111010",
  33771=>"000001100",
  33772=>"000111100",
  33773=>"000011010",
  33774=>"111010101",
  33775=>"111011010",
  33776=>"010110100",
  33777=>"011001010",
  33778=>"010111111",
  33779=>"001000100",
  33780=>"001010000",
  33781=>"100010011",
  33782=>"100000111",
  33783=>"010111000",
  33784=>"000110011",
  33785=>"000110011",
  33786=>"111110110",
  33787=>"110010100",
  33788=>"110110111",
  33789=>"011110100",
  33790=>"001000100",
  33791=>"011111100",
  33792=>"100101001",
  33793=>"101000101",
  33794=>"001101110",
  33795=>"111110001",
  33796=>"011111110",
  33797=>"110101100",
  33798=>"000111010",
  33799=>"111011001",
  33800=>"011010100",
  33801=>"110101110",
  33802=>"001100100",
  33803=>"010010001",
  33804=>"000111010",
  33805=>"101000010",
  33806=>"010100101",
  33807=>"010010110",
  33808=>"001000000",
  33809=>"000011100",
  33810=>"100111111",
  33811=>"000011101",
  33812=>"101000011",
  33813=>"010010100",
  33814=>"001001101",
  33815=>"001000111",
  33816=>"011001100",
  33817=>"111100100",
  33818=>"101100000",
  33819=>"001010010",
  33820=>"101001100",
  33821=>"111010001",
  33822=>"000010000",
  33823=>"001101110",
  33824=>"100100101",
  33825=>"110011010",
  33826=>"111100000",
  33827=>"001111100",
  33828=>"001011010",
  33829=>"100010110",
  33830=>"101011111",
  33831=>"111010111",
  33832=>"100001001",
  33833=>"000111001",
  33834=>"000111101",
  33835=>"111001011",
  33836=>"110000110",
  33837=>"100000100",
  33838=>"110001110",
  33839=>"111110100",
  33840=>"100110001",
  33841=>"001011100",
  33842=>"110110001",
  33843=>"000100100",
  33844=>"000101111",
  33845=>"001101010",
  33846=>"001011111",
  33847=>"101100001",
  33848=>"010001001",
  33849=>"111001101",
  33850=>"100110111",
  33851=>"101001100",
  33852=>"100100000",
  33853=>"000001010",
  33854=>"111111100",
  33855=>"010111101",
  33856=>"110101101",
  33857=>"001011010",
  33858=>"010000111",
  33859=>"001101001",
  33860=>"011000110",
  33861=>"001000110",
  33862=>"111111111",
  33863=>"010100110",
  33864=>"110100011",
  33865=>"101100100",
  33866=>"011001001",
  33867=>"011110110",
  33868=>"001010010",
  33869=>"101111111",
  33870=>"011001110",
  33871=>"110010001",
  33872=>"001010011",
  33873=>"101101110",
  33874=>"000101011",
  33875=>"001010000",
  33876=>"001001100",
  33877=>"001100111",
  33878=>"000011000",
  33879=>"000101010",
  33880=>"011001010",
  33881=>"000001001",
  33882=>"111000010",
  33883=>"000001111",
  33884=>"000010001",
  33885=>"100101110",
  33886=>"010010001",
  33887=>"110011001",
  33888=>"101001010",
  33889=>"001000000",
  33890=>"100010001",
  33891=>"101001011",
  33892=>"001000000",
  33893=>"110011100",
  33894=>"110011001",
  33895=>"010100110",
  33896=>"100010011",
  33897=>"101001010",
  33898=>"010011010",
  33899=>"010000010",
  33900=>"010111111",
  33901=>"000110100",
  33902=>"111101000",
  33903=>"111111011",
  33904=>"100100111",
  33905=>"011011010",
  33906=>"110101101",
  33907=>"100001111",
  33908=>"111111001",
  33909=>"100010010",
  33910=>"100111000",
  33911=>"100101111",
  33912=>"010110010",
  33913=>"001111011",
  33914=>"110010000",
  33915=>"000000000",
  33916=>"110111100",
  33917=>"110100010",
  33918=>"111011100",
  33919=>"000011011",
  33920=>"111111111",
  33921=>"010000010",
  33922=>"100101011",
  33923=>"100000001",
  33924=>"000000011",
  33925=>"010111011",
  33926=>"110010110",
  33927=>"001110001",
  33928=>"000010000",
  33929=>"001101010",
  33930=>"000100100",
  33931=>"111001100",
  33932=>"001010011",
  33933=>"110001101",
  33934=>"010011100",
  33935=>"101001000",
  33936=>"011010110",
  33937=>"111110000",
  33938=>"000010011",
  33939=>"100010101",
  33940=>"011110010",
  33941=>"110111101",
  33942=>"000001001",
  33943=>"000000101",
  33944=>"100000111",
  33945=>"010101101",
  33946=>"011111111",
  33947=>"111010110",
  33948=>"101101110",
  33949=>"010111011",
  33950=>"001110001",
  33951=>"011011000",
  33952=>"000011111",
  33953=>"011101101",
  33954=>"110100010",
  33955=>"001000111",
  33956=>"110010010",
  33957=>"111100010",
  33958=>"100100001",
  33959=>"001010000",
  33960=>"100101011",
  33961=>"011001011",
  33962=>"000000010",
  33963=>"110100110",
  33964=>"100011110",
  33965=>"011101000",
  33966=>"111101111",
  33967=>"111001111",
  33968=>"011011011",
  33969=>"010001011",
  33970=>"001001101",
  33971=>"110101000",
  33972=>"111010101",
  33973=>"011010110",
  33974=>"111111111",
  33975=>"100011100",
  33976=>"000111100",
  33977=>"010011010",
  33978=>"110000111",
  33979=>"011100110",
  33980=>"110010011",
  33981=>"111111100",
  33982=>"011110111",
  33983=>"100011011",
  33984=>"101011010",
  33985=>"110110110",
  33986=>"000001111",
  33987=>"110000010",
  33988=>"100110010",
  33989=>"000101111",
  33990=>"100011100",
  33991=>"000100001",
  33992=>"100010001",
  33993=>"100010000",
  33994=>"001000101",
  33995=>"110101011",
  33996=>"110110110",
  33997=>"001001011",
  33998=>"000100011",
  33999=>"000110011",
  34000=>"100100011",
  34001=>"100111001",
  34002=>"000111111",
  34003=>"010110101",
  34004=>"000000001",
  34005=>"000101001",
  34006=>"101001110",
  34007=>"100011110",
  34008=>"100100000",
  34009=>"000100111",
  34010=>"000001000",
  34011=>"010011010",
  34012=>"011100000",
  34013=>"100010100",
  34014=>"011111001",
  34015=>"010000110",
  34016=>"100001011",
  34017=>"111011110",
  34018=>"011100000",
  34019=>"000000100",
  34020=>"110000000",
  34021=>"101101101",
  34022=>"100110001",
  34023=>"010001010",
  34024=>"101011010",
  34025=>"000011010",
  34026=>"110000111",
  34027=>"011101000",
  34028=>"010010110",
  34029=>"101001110",
  34030=>"100011000",
  34031=>"110010001",
  34032=>"101110010",
  34033=>"001011000",
  34034=>"101001011",
  34035=>"011011001",
  34036=>"010010100",
  34037=>"001010011",
  34038=>"110001001",
  34039=>"101001110",
  34040=>"001110011",
  34041=>"001110101",
  34042=>"000001010",
  34043=>"101000001",
  34044=>"011111001",
  34045=>"011110010",
  34046=>"101010111",
  34047=>"011101111",
  34048=>"100001000",
  34049=>"001001000",
  34050=>"000100100",
  34051=>"110011010",
  34052=>"100001111",
  34053=>"011010110",
  34054=>"000010111",
  34055=>"101101001",
  34056=>"101110100",
  34057=>"100101000",
  34058=>"110011011",
  34059=>"100110110",
  34060=>"000110011",
  34061=>"000110000",
  34062=>"101001101",
  34063=>"000000100",
  34064=>"000010110",
  34065=>"010011000",
  34066=>"110111001",
  34067=>"111000011",
  34068=>"111010111",
  34069=>"001101101",
  34070=>"011001000",
  34071=>"011010111",
  34072=>"101100111",
  34073=>"100011010",
  34074=>"110100100",
  34075=>"111111111",
  34076=>"000001100",
  34077=>"000100100",
  34078=>"110000001",
  34079=>"000101111",
  34080=>"110011000",
  34081=>"000101100",
  34082=>"100110000",
  34083=>"000011001",
  34084=>"001010010",
  34085=>"001010001",
  34086=>"000011011",
  34087=>"111010000",
  34088=>"001100011",
  34089=>"001000111",
  34090=>"111010010",
  34091=>"000111010",
  34092=>"111000010",
  34093=>"111110010",
  34094=>"111100111",
  34095=>"000011010",
  34096=>"000110110",
  34097=>"010000100",
  34098=>"010110101",
  34099=>"100011011",
  34100=>"111010001",
  34101=>"101100010",
  34102=>"010010111",
  34103=>"010100100",
  34104=>"010000000",
  34105=>"000010111",
  34106=>"101110000",
  34107=>"000010010",
  34108=>"100001100",
  34109=>"100101010",
  34110=>"010000100",
  34111=>"101000100",
  34112=>"101001011",
  34113=>"001011101",
  34114=>"011110010",
  34115=>"101101100",
  34116=>"011010000",
  34117=>"000000000",
  34118=>"111000100",
  34119=>"110100110",
  34120=>"110001010",
  34121=>"000010011",
  34122=>"110010110",
  34123=>"001001111",
  34124=>"011001110",
  34125=>"001010001",
  34126=>"110011000",
  34127=>"101010100",
  34128=>"000100010",
  34129=>"000011111",
  34130=>"111100010",
  34131=>"110001010",
  34132=>"101110111",
  34133=>"111011010",
  34134=>"100100010",
  34135=>"001010001",
  34136=>"010000010",
  34137=>"111010111",
  34138=>"010010101",
  34139=>"100011110",
  34140=>"111011110",
  34141=>"001110000",
  34142=>"111101111",
  34143=>"000100101",
  34144=>"001011101",
  34145=>"011001000",
  34146=>"011000100",
  34147=>"011111000",
  34148=>"001000111",
  34149=>"111011011",
  34150=>"111111000",
  34151=>"111101001",
  34152=>"101000000",
  34153=>"011110101",
  34154=>"000100100",
  34155=>"011001111",
  34156=>"010100110",
  34157=>"011010000",
  34158=>"000111001",
  34159=>"111100100",
  34160=>"010101001",
  34161=>"011111110",
  34162=>"110110000",
  34163=>"000110000",
  34164=>"011100001",
  34165=>"111000100",
  34166=>"101110010",
  34167=>"100100010",
  34168=>"010000000",
  34169=>"000111011",
  34170=>"000000001",
  34171=>"010100011",
  34172=>"110101000",
  34173=>"100010101",
  34174=>"010010011",
  34175=>"110000001",
  34176=>"100001011",
  34177=>"011000000",
  34178=>"011101000",
  34179=>"011110011",
  34180=>"001110111",
  34181=>"011010011",
  34182=>"010111000",
  34183=>"011011100",
  34184=>"100100111",
  34185=>"000010001",
  34186=>"110111110",
  34187=>"111101010",
  34188=>"000010111",
  34189=>"110111100",
  34190=>"100011011",
  34191=>"011011100",
  34192=>"110001000",
  34193=>"011101111",
  34194=>"011010010",
  34195=>"010101110",
  34196=>"010100011",
  34197=>"111001111",
  34198=>"000001010",
  34199=>"000111111",
  34200=>"001111011",
  34201=>"111001101",
  34202=>"111001000",
  34203=>"100001001",
  34204=>"110110000",
  34205=>"011001111",
  34206=>"010110101",
  34207=>"001001010",
  34208=>"101010110",
  34209=>"000001111",
  34210=>"010001110",
  34211=>"011110111",
  34212=>"110001010",
  34213=>"110000100",
  34214=>"111100100",
  34215=>"010001000",
  34216=>"001101010",
  34217=>"111101001",
  34218=>"101110110",
  34219=>"100001101",
  34220=>"000010111",
  34221=>"000110110",
  34222=>"101100011",
  34223=>"001001101",
  34224=>"110010010",
  34225=>"101010111",
  34226=>"000101101",
  34227=>"011011001",
  34228=>"100000000",
  34229=>"101101101",
  34230=>"110101111",
  34231=>"010111010",
  34232=>"111100011",
  34233=>"111110111",
  34234=>"100010101",
  34235=>"101011100",
  34236=>"000001001",
  34237=>"110110010",
  34238=>"111000011",
  34239=>"100111101",
  34240=>"100111111",
  34241=>"011010101",
  34242=>"100101010",
  34243=>"100100111",
  34244=>"101111011",
  34245=>"001000001",
  34246=>"100011010",
  34247=>"101000001",
  34248=>"110011110",
  34249=>"000100101",
  34250=>"110011111",
  34251=>"010111010",
  34252=>"100101001",
  34253=>"101011000",
  34254=>"101001000",
  34255=>"101010011",
  34256=>"101010010",
  34257=>"000010000",
  34258=>"100000100",
  34259=>"010000110",
  34260=>"000000010",
  34261=>"010111111",
  34262=>"010010110",
  34263=>"011010010",
  34264=>"101101010",
  34265=>"111111100",
  34266=>"010010000",
  34267=>"010000010",
  34268=>"100110100",
  34269=>"010101101",
  34270=>"101101011",
  34271=>"001111110",
  34272=>"101110110",
  34273=>"111001010",
  34274=>"110010010",
  34275=>"110101010",
  34276=>"100011100",
  34277=>"101000010",
  34278=>"110001001",
  34279=>"011011011",
  34280=>"010001010",
  34281=>"101100001",
  34282=>"110111011",
  34283=>"000000011",
  34284=>"100101101",
  34285=>"000001011",
  34286=>"111001100",
  34287=>"110000000",
  34288=>"101000100",
  34289=>"111011101",
  34290=>"010011100",
  34291=>"000100111",
  34292=>"110101001",
  34293=>"011100000",
  34294=>"000111101",
  34295=>"101110100",
  34296=>"110010100",
  34297=>"011001110",
  34298=>"111111101",
  34299=>"111010010",
  34300=>"111101001",
  34301=>"000101110",
  34302=>"000110111",
  34303=>"001001111",
  34304=>"000110000",
  34305=>"110100100",
  34306=>"110111111",
  34307=>"010111110",
  34308=>"111111101",
  34309=>"011011010",
  34310=>"100011111",
  34311=>"100010000",
  34312=>"100101011",
  34313=>"000111100",
  34314=>"101000100",
  34315=>"111000100",
  34316=>"000110010",
  34317=>"101000000",
  34318=>"000110000",
  34319=>"110111001",
  34320=>"101100110",
  34321=>"001101111",
  34322=>"111101100",
  34323=>"100111001",
  34324=>"110001001",
  34325=>"111101101",
  34326=>"100111100",
  34327=>"101001111",
  34328=>"000000010",
  34329=>"110100110",
  34330=>"011101011",
  34331=>"100111001",
  34332=>"001100111",
  34333=>"011001011",
  34334=>"011000001",
  34335=>"100000000",
  34336=>"100111111",
  34337=>"101100001",
  34338=>"000000011",
  34339=>"100110001",
  34340=>"101111001",
  34341=>"110001101",
  34342=>"011100101",
  34343=>"000001100",
  34344=>"001001111",
  34345=>"011011011",
  34346=>"010010001",
  34347=>"011101111",
  34348=>"001110110",
  34349=>"011001001",
  34350=>"111110101",
  34351=>"010111100",
  34352=>"000000000",
  34353=>"111100011",
  34354=>"100001101",
  34355=>"110010101",
  34356=>"000101011",
  34357=>"001011011",
  34358=>"011101100",
  34359=>"000101111",
  34360=>"101011110",
  34361=>"000001000",
  34362=>"101001001",
  34363=>"111101110",
  34364=>"010001110",
  34365=>"010111001",
  34366=>"101101100",
  34367=>"010111001",
  34368=>"110000100",
  34369=>"100101101",
  34370=>"110111100",
  34371=>"110001100",
  34372=>"110111111",
  34373=>"001011110",
  34374=>"111010011",
  34375=>"000001111",
  34376=>"010001011",
  34377=>"111100110",
  34378=>"111110110",
  34379=>"000010010",
  34380=>"111100111",
  34381=>"000000110",
  34382=>"001011000",
  34383=>"001101100",
  34384=>"111111011",
  34385=>"010011000",
  34386=>"110001000",
  34387=>"100011111",
  34388=>"011010110",
  34389=>"000010001",
  34390=>"000000000",
  34391=>"011101010",
  34392=>"100110110",
  34393=>"110110100",
  34394=>"111100111",
  34395=>"000101101",
  34396=>"001001011",
  34397=>"101000001",
  34398=>"101111011",
  34399=>"110110010",
  34400=>"000101100",
  34401=>"001111001",
  34402=>"010001011",
  34403=>"001101001",
  34404=>"101001001",
  34405=>"010101001",
  34406=>"011111010",
  34407=>"011111010",
  34408=>"010010011",
  34409=>"100101000",
  34410=>"000111000",
  34411=>"011001011",
  34412=>"110110011",
  34413=>"101000001",
  34414=>"111101110",
  34415=>"001011011",
  34416=>"111101010",
  34417=>"000101100",
  34418=>"111101100",
  34419=>"011000101",
  34420=>"000111111",
  34421=>"101010111",
  34422=>"000011010",
  34423=>"110001011",
  34424=>"110001011",
  34425=>"100111110",
  34426=>"101110100",
  34427=>"001100011",
  34428=>"111101010",
  34429=>"100010001",
  34430=>"100110011",
  34431=>"000011010",
  34432=>"010111111",
  34433=>"100010110",
  34434=>"000100110",
  34435=>"001100111",
  34436=>"100001111",
  34437=>"010010111",
  34438=>"111111011",
  34439=>"101100000",
  34440=>"000111101",
  34441=>"011000000",
  34442=>"110111110",
  34443=>"100001000",
  34444=>"010000000",
  34445=>"110010011",
  34446=>"100110101",
  34447=>"000100010",
  34448=>"101100001",
  34449=>"000000000",
  34450=>"110001100",
  34451=>"111100010",
  34452=>"111111101",
  34453=>"011111010",
  34454=>"011010011",
  34455=>"010101001",
  34456=>"000001000",
  34457=>"010011000",
  34458=>"100010111",
  34459=>"111001100",
  34460=>"000100111",
  34461=>"001000010",
  34462=>"001111011",
  34463=>"100000001",
  34464=>"101010010",
  34465=>"101111001",
  34466=>"111111000",
  34467=>"110001010",
  34468=>"001111000",
  34469=>"010001111",
  34470=>"001001110",
  34471=>"000000000",
  34472=>"110011011",
  34473=>"001111111",
  34474=>"111011110",
  34475=>"110001010",
  34476=>"000000101",
  34477=>"101110000",
  34478=>"101101000",
  34479=>"000101011",
  34480=>"000010100",
  34481=>"000101110",
  34482=>"001001110",
  34483=>"010011010",
  34484=>"110011101",
  34485=>"011111101",
  34486=>"011110110",
  34487=>"000101100",
  34488=>"110011101",
  34489=>"011011011",
  34490=>"001110100",
  34491=>"100110010",
  34492=>"010100110",
  34493=>"011000011",
  34494=>"000011001",
  34495=>"110010100",
  34496=>"000011001",
  34497=>"001001111",
  34498=>"010011100",
  34499=>"000000011",
  34500=>"010000111",
  34501=>"000000001",
  34502=>"010100100",
  34503=>"010110110",
  34504=>"010100111",
  34505=>"011001011",
  34506=>"110011111",
  34507=>"111010011",
  34508=>"001001011",
  34509=>"111000100",
  34510=>"101111010",
  34511=>"111111010",
  34512=>"111100001",
  34513=>"111011010",
  34514=>"100010001",
  34515=>"000100011",
  34516=>"101100001",
  34517=>"111011001",
  34518=>"001001000",
  34519=>"001100110",
  34520=>"000011100",
  34521=>"101111010",
  34522=>"000001000",
  34523=>"111100001",
  34524=>"101010000",
  34525=>"111110000",
  34526=>"011001001",
  34527=>"011011011",
  34528=>"011001111",
  34529=>"001001110",
  34530=>"111000011",
  34531=>"110000010",
  34532=>"001001110",
  34533=>"001011101",
  34534=>"000101110",
  34535=>"001000010",
  34536=>"100101101",
  34537=>"000100011",
  34538=>"010010100",
  34539=>"000110111",
  34540=>"000000101",
  34541=>"100011010",
  34542=>"110111110",
  34543=>"010010001",
  34544=>"100111000",
  34545=>"111001110",
  34546=>"010001101",
  34547=>"011000000",
  34548=>"100111101",
  34549=>"001101101",
  34550=>"110111111",
  34551=>"011010010",
  34552=>"101101101",
  34553=>"001011111",
  34554=>"010010011",
  34555=>"000000011",
  34556=>"110100010",
  34557=>"010101001",
  34558=>"001011111",
  34559=>"101110111",
  34560=>"010000010",
  34561=>"001111100",
  34562=>"001111000",
  34563=>"111101101",
  34564=>"101011111",
  34565=>"101010100",
  34566=>"000100100",
  34567=>"101001001",
  34568=>"100000010",
  34569=>"110101000",
  34570=>"111101011",
  34571=>"010110101",
  34572=>"010011111",
  34573=>"010101000",
  34574=>"100110100",
  34575=>"111010011",
  34576=>"000010000",
  34577=>"010000100",
  34578=>"011110101",
  34579=>"011010111",
  34580=>"110111000",
  34581=>"100010000",
  34582=>"000001001",
  34583=>"010001011",
  34584=>"000111101",
  34585=>"101010000",
  34586=>"101111110",
  34587=>"001110110",
  34588=>"100001000",
  34589=>"010101000",
  34590=>"010010010",
  34591=>"101110000",
  34592=>"101101111",
  34593=>"001000000",
  34594=>"111000110",
  34595=>"010110101",
  34596=>"011100111",
  34597=>"101010110",
  34598=>"111010001",
  34599=>"011001011",
  34600=>"010111111",
  34601=>"010110000",
  34602=>"111000000",
  34603=>"100111010",
  34604=>"011000111",
  34605=>"000111000",
  34606=>"110110101",
  34607=>"101110110",
  34608=>"000111110",
  34609=>"101101110",
  34610=>"100100010",
  34611=>"100000000",
  34612=>"111000000",
  34613=>"111100000",
  34614=>"110111010",
  34615=>"011110110",
  34616=>"110010011",
  34617=>"001100101",
  34618=>"001101000",
  34619=>"011111011",
  34620=>"010101011",
  34621=>"100000001",
  34622=>"010000001",
  34623=>"001101111",
  34624=>"101100110",
  34625=>"001000000",
  34626=>"111101000",
  34627=>"001110001",
  34628=>"100000100",
  34629=>"011100011",
  34630=>"001001101",
  34631=>"010110000",
  34632=>"001101001",
  34633=>"001101100",
  34634=>"110110111",
  34635=>"110000000",
  34636=>"111000001",
  34637=>"100010000",
  34638=>"100011001",
  34639=>"101001111",
  34640=>"110111111",
  34641=>"011101111",
  34642=>"000100000",
  34643=>"011110001",
  34644=>"010110111",
  34645=>"100111101",
  34646=>"000011111",
  34647=>"101011101",
  34648=>"000110000",
  34649=>"011110000",
  34650=>"011110100",
  34651=>"000001101",
  34652=>"101101101",
  34653=>"001001111",
  34654=>"110100001",
  34655=>"010111111",
  34656=>"111001010",
  34657=>"000101111",
  34658=>"000101111",
  34659=>"101011111",
  34660=>"111110110",
  34661=>"000010001",
  34662=>"011111011",
  34663=>"110101000",
  34664=>"000000110",
  34665=>"001111110",
  34666=>"011011000",
  34667=>"010101110",
  34668=>"000000000",
  34669=>"111101101",
  34670=>"110111001",
  34671=>"110011001",
  34672=>"101100110",
  34673=>"111100110",
  34674=>"000010110",
  34675=>"001011111",
  34676=>"001100100",
  34677=>"110100010",
  34678=>"010000101",
  34679=>"101100100",
  34680=>"110000000",
  34681=>"110000010",
  34682=>"111111000",
  34683=>"010000001",
  34684=>"000110010",
  34685=>"001111100",
  34686=>"001000111",
  34687=>"010000100",
  34688=>"111001001",
  34689=>"000101011",
  34690=>"011111011",
  34691=>"111101000",
  34692=>"000111010",
  34693=>"010001100",
  34694=>"000111000",
  34695=>"010001101",
  34696=>"010110110",
  34697=>"110001101",
  34698=>"101111000",
  34699=>"000101001",
  34700=>"110000011",
  34701=>"001100110",
  34702=>"000100011",
  34703=>"110010111",
  34704=>"000011001",
  34705=>"101110011",
  34706=>"000001000",
  34707=>"111000100",
  34708=>"101111001",
  34709=>"100111110",
  34710=>"101011001",
  34711=>"011110001",
  34712=>"011111001",
  34713=>"100010001",
  34714=>"110101010",
  34715=>"000100101",
  34716=>"000010110",
  34717=>"110101111",
  34718=>"110011110",
  34719=>"100110011",
  34720=>"101100111",
  34721=>"010100011",
  34722=>"100101000",
  34723=>"001010100",
  34724=>"100100000",
  34725=>"000111111",
  34726=>"100101100",
  34727=>"101001110",
  34728=>"110010110",
  34729=>"001011010",
  34730=>"111100010",
  34731=>"011000010",
  34732=>"100000110",
  34733=>"111000001",
  34734=>"011000001",
  34735=>"101011010",
  34736=>"011000110",
  34737=>"001000101",
  34738=>"010000000",
  34739=>"011101100",
  34740=>"010010111",
  34741=>"010111100",
  34742=>"011001111",
  34743=>"110001011",
  34744=>"111110111",
  34745=>"100000110",
  34746=>"000001000",
  34747=>"111111101",
  34748=>"111101101",
  34749=>"100101101",
  34750=>"110011001",
  34751=>"000000011",
  34752=>"111001000",
  34753=>"101001100",
  34754=>"101000001",
  34755=>"101010000",
  34756=>"011001111",
  34757=>"100011110",
  34758=>"001111111",
  34759=>"101101001",
  34760=>"100111011",
  34761=>"011111010",
  34762=>"101001011",
  34763=>"111110111",
  34764=>"011000100",
  34765=>"110001111",
  34766=>"010110111",
  34767=>"100110110",
  34768=>"011110101",
  34769=>"000000000",
  34770=>"011000011",
  34771=>"101101101",
  34772=>"111101101",
  34773=>"010101000",
  34774=>"010000100",
  34775=>"110011101",
  34776=>"100111111",
  34777=>"100110111",
  34778=>"001011000",
  34779=>"001110001",
  34780=>"101111010",
  34781=>"001111011",
  34782=>"001100101",
  34783=>"100100101",
  34784=>"111111001",
  34785=>"011100100",
  34786=>"001101110",
  34787=>"000100110",
  34788=>"100100101",
  34789=>"000000100",
  34790=>"010111001",
  34791=>"101101011",
  34792=>"000100001",
  34793=>"001011110",
  34794=>"010110011",
  34795=>"100100000",
  34796=>"001001011",
  34797=>"101011000",
  34798=>"100000111",
  34799=>"011100010",
  34800=>"110001000",
  34801=>"110110000",
  34802=>"000110101",
  34803=>"111001111",
  34804=>"010000000",
  34805=>"000110011",
  34806=>"001011011",
  34807=>"101110011",
  34808=>"000010111",
  34809=>"010110100",
  34810=>"000000100",
  34811=>"101010001",
  34812=>"010011011",
  34813=>"101110101",
  34814=>"001010011",
  34815=>"001001001",
  34816=>"010111001",
  34817=>"111000111",
  34818=>"110100111",
  34819=>"010100011",
  34820=>"001011100",
  34821=>"011110011",
  34822=>"100000000",
  34823=>"110101011",
  34824=>"001001010",
  34825=>"001011000",
  34826=>"111100010",
  34827=>"100000111",
  34828=>"011001011",
  34829=>"001110011",
  34830=>"001110001",
  34831=>"101000111",
  34832=>"010101000",
  34833=>"110100110",
  34834=>"110000111",
  34835=>"011001111",
  34836=>"000101111",
  34837=>"001000100",
  34838=>"000011110",
  34839=>"100001001",
  34840=>"010001111",
  34841=>"001010111",
  34842=>"110100101",
  34843=>"011101100",
  34844=>"011100110",
  34845=>"100011110",
  34846=>"011111101",
  34847=>"011011001",
  34848=>"111110110",
  34849=>"101100101",
  34850=>"000010000",
  34851=>"100110001",
  34852=>"110001001",
  34853=>"000111000",
  34854=>"101101010",
  34855=>"001111000",
  34856=>"101111111",
  34857=>"100010111",
  34858=>"110001100",
  34859=>"001101011",
  34860=>"110101100",
  34861=>"000110010",
  34862=>"110001001",
  34863=>"111000000",
  34864=>"101001011",
  34865=>"010100000",
  34866=>"001110101",
  34867=>"111001010",
  34868=>"001011110",
  34869=>"100001101",
  34870=>"011110001",
  34871=>"110111100",
  34872=>"001001000",
  34873=>"100000010",
  34874=>"111000011",
  34875=>"011011001",
  34876=>"000000100",
  34877=>"010101001",
  34878=>"011011001",
  34879=>"100101111",
  34880=>"011110110",
  34881=>"011111101",
  34882=>"100010111",
  34883=>"010011101",
  34884=>"010011000",
  34885=>"101101001",
  34886=>"110110010",
  34887=>"010111100",
  34888=>"101011101",
  34889=>"010110101",
  34890=>"000000000",
  34891=>"000001000",
  34892=>"001001001",
  34893=>"110001100",
  34894=>"011011001",
  34895=>"010010101",
  34896=>"011011101",
  34897=>"100000110",
  34898=>"100001101",
  34899=>"000110101",
  34900=>"100100100",
  34901=>"101110100",
  34902=>"110010110",
  34903=>"111011101",
  34904=>"111001011",
  34905=>"110000111",
  34906=>"001001110",
  34907=>"100001001",
  34908=>"000111001",
  34909=>"001001001",
  34910=>"111010000",
  34911=>"101100100",
  34912=>"110110000",
  34913=>"001011101",
  34914=>"011001100",
  34915=>"010010000",
  34916=>"110000011",
  34917=>"001000011",
  34918=>"101001110",
  34919=>"011011011",
  34920=>"100000101",
  34921=>"110011010",
  34922=>"111011000",
  34923=>"100010011",
  34924=>"110011100",
  34925=>"100101000",
  34926=>"011000111",
  34927=>"011101000",
  34928=>"110011111",
  34929=>"000101110",
  34930=>"110111001",
  34931=>"100001011",
  34932=>"010010001",
  34933=>"110100111",
  34934=>"000111101",
  34935=>"111010111",
  34936=>"000110111",
  34937=>"001101001",
  34938=>"101110001",
  34939=>"011001010",
  34940=>"001011010",
  34941=>"011111001",
  34942=>"001011011",
  34943=>"100111111",
  34944=>"000100011",
  34945=>"011000001",
  34946=>"101011110",
  34947=>"100001111",
  34948=>"000111111",
  34949=>"100101001",
  34950=>"101100010",
  34951=>"110111011",
  34952=>"111001100",
  34953=>"101011100",
  34954=>"111111110",
  34955=>"010001110",
  34956=>"110101111",
  34957=>"001110110",
  34958=>"000010011",
  34959=>"010000100",
  34960=>"001101011",
  34961=>"100001110",
  34962=>"111010001",
  34963=>"011100110",
  34964=>"001000100",
  34965=>"011101000",
  34966=>"111111001",
  34967=>"010100011",
  34968=>"101100000",
  34969=>"011101010",
  34970=>"110000111",
  34971=>"000111000",
  34972=>"000101100",
  34973=>"110100010",
  34974=>"010010110",
  34975=>"011011110",
  34976=>"100011000",
  34977=>"011100000",
  34978=>"100101010",
  34979=>"000110011",
  34980=>"100110111",
  34981=>"010000011",
  34982=>"100000000",
  34983=>"000001000",
  34984=>"000011011",
  34985=>"111111110",
  34986=>"100011100",
  34987=>"111111011",
  34988=>"100100010",
  34989=>"111100001",
  34990=>"111101001",
  34991=>"000000110",
  34992=>"010001010",
  34993=>"001011111",
  34994=>"000001011",
  34995=>"010110100",
  34996=>"110010010",
  34997=>"011100000",
  34998=>"100011011",
  34999=>"110001110",
  35000=>"100001000",
  35001=>"000101101",
  35002=>"010000101",
  35003=>"010010110",
  35004=>"100001111",
  35005=>"100100010",
  35006=>"001101101",
  35007=>"001111000",
  35008=>"101011111",
  35009=>"011111111",
  35010=>"100010101",
  35011=>"101110100",
  35012=>"001100010",
  35013=>"111001111",
  35014=>"111101101",
  35015=>"111111111",
  35016=>"110011000",
  35017=>"111110011",
  35018=>"101010010",
  35019=>"001011000",
  35020=>"000110011",
  35021=>"000100111",
  35022=>"010111001",
  35023=>"011001111",
  35024=>"111100100",
  35025=>"111100000",
  35026=>"110111001",
  35027=>"001010011",
  35028=>"001001110",
  35029=>"000000111",
  35030=>"110010000",
  35031=>"101000110",
  35032=>"011010100",
  35033=>"111100100",
  35034=>"001011000",
  35035=>"011000010",
  35036=>"110111101",
  35037=>"010101101",
  35038=>"001001010",
  35039=>"101100111",
  35040=>"011001101",
  35041=>"010000110",
  35042=>"011010000",
  35043=>"010000100",
  35044=>"000010000",
  35045=>"111100110",
  35046=>"010000110",
  35047=>"111011000",
  35048=>"001101001",
  35049=>"000000011",
  35050=>"110011011",
  35051=>"100011000",
  35052=>"100100011",
  35053=>"011001110",
  35054=>"011001010",
  35055=>"101101010",
  35056=>"100011010",
  35057=>"101111111",
  35058=>"001101111",
  35059=>"001111011",
  35060=>"110111001",
  35061=>"111101011",
  35062=>"001001001",
  35063=>"000000100",
  35064=>"110000110",
  35065=>"110000010",
  35066=>"011110011",
  35067=>"001001001",
  35068=>"001110101",
  35069=>"111111010",
  35070=>"011000100",
  35071=>"111001111",
  35072=>"110001111",
  35073=>"100001110",
  35074=>"111010101",
  35075=>"110100100",
  35076=>"100000001",
  35077=>"000001101",
  35078=>"001101011",
  35079=>"000111111",
  35080=>"000001111",
  35081=>"000011101",
  35082=>"000101011",
  35083=>"011011000",
  35084=>"011100001",
  35085=>"110010101",
  35086=>"001101001",
  35087=>"011011010",
  35088=>"010001111",
  35089=>"000011111",
  35090=>"000001011",
  35091=>"111111100",
  35092=>"111000101",
  35093=>"000011011",
  35094=>"110011001",
  35095=>"100100110",
  35096=>"100111110",
  35097=>"010100011",
  35098=>"000001101",
  35099=>"010110101",
  35100=>"000000001",
  35101=>"111000000",
  35102=>"111000110",
  35103=>"010111100",
  35104=>"111101101",
  35105=>"011111001",
  35106=>"111010110",
  35107=>"100000011",
  35108=>"100110011",
  35109=>"001101000",
  35110=>"001000000",
  35111=>"001100000",
  35112=>"001100100",
  35113=>"000111110",
  35114=>"100110111",
  35115=>"010010010",
  35116=>"111101011",
  35117=>"001011011",
  35118=>"101011111",
  35119=>"111000010",
  35120=>"011100011",
  35121=>"110111101",
  35122=>"110010101",
  35123=>"000111000",
  35124=>"001001001",
  35125=>"001011001",
  35126=>"011100111",
  35127=>"011100101",
  35128=>"001001011",
  35129=>"101001001",
  35130=>"111000101",
  35131=>"011010111",
  35132=>"110111001",
  35133=>"010111010",
  35134=>"010100100",
  35135=>"101001111",
  35136=>"001000000",
  35137=>"000010011",
  35138=>"100101110",
  35139=>"000110101",
  35140=>"000110000",
  35141=>"001010010",
  35142=>"010000000",
  35143=>"101001001",
  35144=>"100000100",
  35145=>"011111100",
  35146=>"000010111",
  35147=>"101101100",
  35148=>"000000010",
  35149=>"011011010",
  35150=>"000000010",
  35151=>"011011100",
  35152=>"000101001",
  35153=>"110001000",
  35154=>"100001100",
  35155=>"101110101",
  35156=>"110010110",
  35157=>"000000110",
  35158=>"001111010",
  35159=>"001111000",
  35160=>"000100100",
  35161=>"101000111",
  35162=>"100001101",
  35163=>"011000111",
  35164=>"010110011",
  35165=>"111001100",
  35166=>"001010100",
  35167=>"011000011",
  35168=>"111100011",
  35169=>"100010111",
  35170=>"000010110",
  35171=>"101101111",
  35172=>"001111101",
  35173=>"011111001",
  35174=>"000001110",
  35175=>"110110110",
  35176=>"000010100",
  35177=>"000001111",
  35178=>"001100100",
  35179=>"001000111",
  35180=>"110011101",
  35181=>"000101110",
  35182=>"011011000",
  35183=>"000100101",
  35184=>"001010110",
  35185=>"000100011",
  35186=>"110010011",
  35187=>"101010011",
  35188=>"101111000",
  35189=>"001001100",
  35190=>"010001000",
  35191=>"101010011",
  35192=>"100010010",
  35193=>"100100110",
  35194=>"001111101",
  35195=>"000100101",
  35196=>"010011110",
  35197=>"101111011",
  35198=>"001100001",
  35199=>"110001100",
  35200=>"101101010",
  35201=>"101001010",
  35202=>"010100010",
  35203=>"001100010",
  35204=>"000110011",
  35205=>"001011000",
  35206=>"011010000",
  35207=>"010011000",
  35208=>"000111010",
  35209=>"011010100",
  35210=>"001000110",
  35211=>"111101101",
  35212=>"010010000",
  35213=>"100000011",
  35214=>"101101001",
  35215=>"001100010",
  35216=>"001001110",
  35217=>"011100101",
  35218=>"010111010",
  35219=>"110100000",
  35220=>"010011110",
  35221=>"111010010",
  35222=>"101100100",
  35223=>"001101001",
  35224=>"001100000",
  35225=>"001011011",
  35226=>"001001000",
  35227=>"111110001",
  35228=>"001011011",
  35229=>"101001111",
  35230=>"001100101",
  35231=>"001110011",
  35232=>"111001010",
  35233=>"100111111",
  35234=>"010110101",
  35235=>"110100001",
  35236=>"011011011",
  35237=>"000010100",
  35238=>"100011000",
  35239=>"111110000",
  35240=>"011110101",
  35241=>"010011101",
  35242=>"001101100",
  35243=>"000011001",
  35244=>"011011110",
  35245=>"101110111",
  35246=>"101000010",
  35247=>"010101011",
  35248=>"010100100",
  35249=>"111110100",
  35250=>"100010000",
  35251=>"000001011",
  35252=>"111101101",
  35253=>"111011011",
  35254=>"001111010",
  35255=>"101111110",
  35256=>"100011100",
  35257=>"100000000",
  35258=>"000010010",
  35259=>"101001001",
  35260=>"010101101",
  35261=>"011101101",
  35262=>"011010110",
  35263=>"001000101",
  35264=>"100010010",
  35265=>"100100000",
  35266=>"110010001",
  35267=>"011100001",
  35268=>"010000100",
  35269=>"010110111",
  35270=>"110100101",
  35271=>"101001110",
  35272=>"110101010",
  35273=>"101101110",
  35274=>"111001100",
  35275=>"000011101",
  35276=>"010100010",
  35277=>"000111001",
  35278=>"100111110",
  35279=>"010101010",
  35280=>"000010000",
  35281=>"100100111",
  35282=>"011111101",
  35283=>"111000001",
  35284=>"110100011",
  35285=>"010000011",
  35286=>"110101111",
  35287=>"111000101",
  35288=>"001111001",
  35289=>"001001011",
  35290=>"010000010",
  35291=>"110011000",
  35292=>"111111011",
  35293=>"001100011",
  35294=>"010101010",
  35295=>"111000100",
  35296=>"001011110",
  35297=>"001111000",
  35298=>"101011010",
  35299=>"110111001",
  35300=>"000001001",
  35301=>"100100111",
  35302=>"000011101",
  35303=>"111111101",
  35304=>"010000000",
  35305=>"101010000",
  35306=>"001100011",
  35307=>"111100110",
  35308=>"110011011",
  35309=>"001100011",
  35310=>"110010000",
  35311=>"101101000",
  35312=>"001110100",
  35313=>"101001100",
  35314=>"111011100",
  35315=>"000101100",
  35316=>"110111101",
  35317=>"110110110",
  35318=>"111101010",
  35319=>"101001111",
  35320=>"111001101",
  35321=>"111110101",
  35322=>"100001100",
  35323=>"000011101",
  35324=>"101001100",
  35325=>"000100000",
  35326=>"001010011",
  35327=>"010000000",
  35328=>"101001100",
  35329=>"101001010",
  35330=>"000000000",
  35331=>"011101010",
  35332=>"010001111",
  35333=>"111001010",
  35334=>"101110001",
  35335=>"010011110",
  35336=>"011001101",
  35337=>"111011100",
  35338=>"111100111",
  35339=>"000001001",
  35340=>"100100001",
  35341=>"011111011",
  35342=>"111110000",
  35343=>"111100000",
  35344=>"000110101",
  35345=>"011111111",
  35346=>"110011110",
  35347=>"100101000",
  35348=>"010000111",
  35349=>"111011010",
  35350=>"000010001",
  35351=>"111101001",
  35352=>"001011101",
  35353=>"111001010",
  35354=>"111001001",
  35355=>"000010110",
  35356=>"110101110",
  35357=>"011001110",
  35358=>"000001011",
  35359=>"000100111",
  35360=>"110010011",
  35361=>"111100000",
  35362=>"101000111",
  35363=>"011101011",
  35364=>"110100101",
  35365=>"111011001",
  35366=>"010011010",
  35367=>"100010001",
  35368=>"110001001",
  35369=>"011111010",
  35370=>"010110011",
  35371=>"110111100",
  35372=>"000101001",
  35373=>"100000010",
  35374=>"101111101",
  35375=>"110101000",
  35376=>"010101110",
  35377=>"001010011",
  35378=>"000011100",
  35379=>"110111011",
  35380=>"100111111",
  35381=>"100100110",
  35382=>"101110011",
  35383=>"100100101",
  35384=>"011010011",
  35385=>"000101010",
  35386=>"010011001",
  35387=>"101101011",
  35388=>"100111111",
  35389=>"101001111",
  35390=>"011000101",
  35391=>"110110100",
  35392=>"101111011",
  35393=>"000111111",
  35394=>"101001110",
  35395=>"010001011",
  35396=>"000100101",
  35397=>"110001010",
  35398=>"110001000",
  35399=>"010110101",
  35400=>"010100001",
  35401=>"011101101",
  35402=>"100001000",
  35403=>"101001100",
  35404=>"011100111",
  35405=>"000100101",
  35406=>"111010101",
  35407=>"011111011",
  35408=>"100011111",
  35409=>"110001001",
  35410=>"111001110",
  35411=>"001110101",
  35412=>"000000111",
  35413=>"001010010",
  35414=>"110000111",
  35415=>"011000111",
  35416=>"000111101",
  35417=>"011011111",
  35418=>"011010000",
  35419=>"011100010",
  35420=>"001010001",
  35421=>"101010001",
  35422=>"000110110",
  35423=>"111100010",
  35424=>"110111011",
  35425=>"001011000",
  35426=>"011001010",
  35427=>"110111001",
  35428=>"100111010",
  35429=>"001100110",
  35430=>"101111110",
  35431=>"100101100",
  35432=>"010010111",
  35433=>"000010110",
  35434=>"000100010",
  35435=>"001100000",
  35436=>"001100001",
  35437=>"010101101",
  35438=>"111101110",
  35439=>"110001001",
  35440=>"011101010",
  35441=>"101000101",
  35442=>"110110010",
  35443=>"101100000",
  35444=>"001010001",
  35445=>"110000101",
  35446=>"111011000",
  35447=>"010011101",
  35448=>"101110101",
  35449=>"110111001",
  35450=>"001011010",
  35451=>"100011100",
  35452=>"101100110",
  35453=>"110011010",
  35454=>"101000001",
  35455=>"110011101",
  35456=>"000001111",
  35457=>"101000100",
  35458=>"010111010",
  35459=>"000110110",
  35460=>"100100000",
  35461=>"001000101",
  35462=>"110111110",
  35463=>"100100101",
  35464=>"010100001",
  35465=>"110000011",
  35466=>"000000010",
  35467=>"101100100",
  35468=>"011000110",
  35469=>"111111001",
  35470=>"011111000",
  35471=>"000011010",
  35472=>"011101011",
  35473=>"001010000",
  35474=>"000011000",
  35475=>"000000001",
  35476=>"101001110",
  35477=>"001001110",
  35478=>"101100011",
  35479=>"101111011",
  35480=>"111010000",
  35481=>"011100111",
  35482=>"100001110",
  35483=>"110011001",
  35484=>"110100100",
  35485=>"100000110",
  35486=>"010000000",
  35487=>"010111000",
  35488=>"000011100",
  35489=>"111010000",
  35490=>"111110110",
  35491=>"110111001",
  35492=>"101011001",
  35493=>"011100011",
  35494=>"111111111",
  35495=>"001111111",
  35496=>"111110111",
  35497=>"100101000",
  35498=>"011110111",
  35499=>"000010010",
  35500=>"000111110",
  35501=>"100001011",
  35502=>"110011101",
  35503=>"101101000",
  35504=>"101001000",
  35505=>"001110100",
  35506=>"010010011",
  35507=>"100110111",
  35508=>"101100100",
  35509=>"010100110",
  35510=>"000011000",
  35511=>"101000001",
  35512=>"000100110",
  35513=>"001011110",
  35514=>"010110111",
  35515=>"111111100",
  35516=>"101000010",
  35517=>"110111100",
  35518=>"010111001",
  35519=>"000001110",
  35520=>"111100101",
  35521=>"111001010",
  35522=>"101000101",
  35523=>"000000001",
  35524=>"111000111",
  35525=>"010110001",
  35526=>"100110101",
  35527=>"010100011",
  35528=>"110111111",
  35529=>"001001000",
  35530=>"100100101",
  35531=>"000001001",
  35532=>"010100100",
  35533=>"010101010",
  35534=>"110110111",
  35535=>"101011101",
  35536=>"000110101",
  35537=>"011010100",
  35538=>"111011001",
  35539=>"100100111",
  35540=>"011111000",
  35541=>"010100010",
  35542=>"010101111",
  35543=>"111010000",
  35544=>"100010010",
  35545=>"111110011",
  35546=>"101100110",
  35547=>"011010101",
  35548=>"001001001",
  35549=>"110001101",
  35550=>"000110101",
  35551=>"011111111",
  35552=>"001100011",
  35553=>"111100000",
  35554=>"011000011",
  35555=>"111011010",
  35556=>"000100111",
  35557=>"110100111",
  35558=>"101000000",
  35559=>"110010010",
  35560=>"000010110",
  35561=>"001110010",
  35562=>"011110110",
  35563=>"100011000",
  35564=>"001100001",
  35565=>"100010101",
  35566=>"001101100",
  35567=>"111011111",
  35568=>"111111111",
  35569=>"110110000",
  35570=>"000001101",
  35571=>"101000001",
  35572=>"011110101",
  35573=>"001000111",
  35574=>"101001100",
  35575=>"010010111",
  35576=>"111100111",
  35577=>"011000000",
  35578=>"000011000",
  35579=>"101001010",
  35580=>"110111001",
  35581=>"110111010",
  35582=>"101001011",
  35583=>"011110110",
  35584=>"010001111",
  35585=>"100101101",
  35586=>"011001010",
  35587=>"001110100",
  35588=>"110110010",
  35589=>"101101011",
  35590=>"111000110",
  35591=>"011100101",
  35592=>"101001101",
  35593=>"111111101",
  35594=>"111101001",
  35595=>"100101000",
  35596=>"001011101",
  35597=>"010000100",
  35598=>"011000110",
  35599=>"001110111",
  35600=>"100111111",
  35601=>"101010001",
  35602=>"010000000",
  35603=>"110001100",
  35604=>"011001111",
  35605=>"000111000",
  35606=>"111001011",
  35607=>"100001001",
  35608=>"011011000",
  35609=>"000000001",
  35610=>"000010111",
  35611=>"100000101",
  35612=>"110101000",
  35613=>"100011000",
  35614=>"110000111",
  35615=>"111110010",
  35616=>"100111010",
  35617=>"111011010",
  35618=>"100000111",
  35619=>"010010111",
  35620=>"011001000",
  35621=>"111100100",
  35622=>"100011111",
  35623=>"100111000",
  35624=>"001010101",
  35625=>"001001001",
  35626=>"000111110",
  35627=>"100101001",
  35628=>"100100010",
  35629=>"000110100",
  35630=>"001001111",
  35631=>"100011001",
  35632=>"000001000",
  35633=>"101101111",
  35634=>"011010011",
  35635=>"101010101",
  35636=>"111111111",
  35637=>"000000111",
  35638=>"011111101",
  35639=>"100111000",
  35640=>"101101010",
  35641=>"111101000",
  35642=>"011011000",
  35643=>"101010001",
  35644=>"110001000",
  35645=>"111000000",
  35646=>"011111010",
  35647=>"011011110",
  35648=>"001110000",
  35649=>"111011100",
  35650=>"111101100",
  35651=>"111000110",
  35652=>"101001001",
  35653=>"001011011",
  35654=>"011100101",
  35655=>"111111100",
  35656=>"010011001",
  35657=>"101000111",
  35658=>"011101001",
  35659=>"000001110",
  35660=>"110111110",
  35661=>"110101011",
  35662=>"000110111",
  35663=>"111011110",
  35664=>"101101111",
  35665=>"000001000",
  35666=>"101010110",
  35667=>"001010000",
  35668=>"010100001",
  35669=>"001100011",
  35670=>"001111000",
  35671=>"001100100",
  35672=>"110110111",
  35673=>"110011000",
  35674=>"110001100",
  35675=>"011111100",
  35676=>"111010000",
  35677=>"001011100",
  35678=>"110100111",
  35679=>"100000100",
  35680=>"100000011",
  35681=>"100110010",
  35682=>"001000100",
  35683=>"111111101",
  35684=>"001001011",
  35685=>"010000001",
  35686=>"011111001",
  35687=>"101101001",
  35688=>"101010001",
  35689=>"101000001",
  35690=>"100000101",
  35691=>"101000000",
  35692=>"110110011",
  35693=>"011001000",
  35694=>"000011001",
  35695=>"110111110",
  35696=>"010101011",
  35697=>"010101010",
  35698=>"101110100",
  35699=>"100000011",
  35700=>"000010101",
  35701=>"000101010",
  35702=>"011011001",
  35703=>"101001100",
  35704=>"001001111",
  35705=>"000110110",
  35706=>"000011000",
  35707=>"000100111",
  35708=>"101110010",
  35709=>"001111101",
  35710=>"111001001",
  35711=>"010110000",
  35712=>"000110000",
  35713=>"010011110",
  35714=>"110100011",
  35715=>"101101100",
  35716=>"011110000",
  35717=>"011111101",
  35718=>"000111010",
  35719=>"010101011",
  35720=>"100111100",
  35721=>"000101011",
  35722=>"100110000",
  35723=>"010010011",
  35724=>"100100000",
  35725=>"100010111",
  35726=>"000100110",
  35727=>"001000001",
  35728=>"101101111",
  35729=>"001111011",
  35730=>"101111101",
  35731=>"011000010",
  35732=>"111111110",
  35733=>"001100110",
  35734=>"000011110",
  35735=>"011011011",
  35736=>"001111111",
  35737=>"001001000",
  35738=>"100110100",
  35739=>"111000100",
  35740=>"010000011",
  35741=>"011110010",
  35742=>"110000110",
  35743=>"111011111",
  35744=>"011111001",
  35745=>"011100000",
  35746=>"011110001",
  35747=>"110110010",
  35748=>"000111111",
  35749=>"010011001",
  35750=>"010100000",
  35751=>"110010010",
  35752=>"001110000",
  35753=>"100000000",
  35754=>"010111111",
  35755=>"000011111",
  35756=>"011011110",
  35757=>"011010101",
  35758=>"101000100",
  35759=>"001001110",
  35760=>"110001111",
  35761=>"000110110",
  35762=>"111001101",
  35763=>"100101101",
  35764=>"100011001",
  35765=>"101100000",
  35766=>"011100100",
  35767=>"111100111",
  35768=>"001111000",
  35769=>"010110010",
  35770=>"110100101",
  35771=>"100011000",
  35772=>"011010010",
  35773=>"001001101",
  35774=>"010110001",
  35775=>"100101000",
  35776=>"001111000",
  35777=>"001101100",
  35778=>"000101101",
  35779=>"010101011",
  35780=>"101100111",
  35781=>"001110001",
  35782=>"011110010",
  35783=>"111100001",
  35784=>"010001001",
  35785=>"011111011",
  35786=>"010010001",
  35787=>"101001100",
  35788=>"100010011",
  35789=>"010100011",
  35790=>"001111101",
  35791=>"000011100",
  35792=>"011111011",
  35793=>"000110000",
  35794=>"101011011",
  35795=>"010101110",
  35796=>"111101101",
  35797=>"011101011",
  35798=>"000000000",
  35799=>"110010110",
  35800=>"000010001",
  35801=>"110001101",
  35802=>"101000000",
  35803=>"111010001",
  35804=>"100001101",
  35805=>"000100101",
  35806=>"101010010",
  35807=>"000000000",
  35808=>"000000010",
  35809=>"101101011",
  35810=>"000011111",
  35811=>"000100010",
  35812=>"001011111",
  35813=>"111101111",
  35814=>"011011010",
  35815=>"111001111",
  35816=>"000001000",
  35817=>"010011110",
  35818=>"000010000",
  35819=>"111000010",
  35820=>"011010000",
  35821=>"101000110",
  35822=>"110110111",
  35823=>"100000100",
  35824=>"011011000",
  35825=>"111111100",
  35826=>"001110110",
  35827=>"111101010",
  35828=>"001001000",
  35829=>"101101100",
  35830=>"101000101",
  35831=>"000010111",
  35832=>"011001000",
  35833=>"011111010",
  35834=>"110001000",
  35835=>"100010011",
  35836=>"110100101",
  35837=>"111100110",
  35838=>"101011110",
  35839=>"110110111",
  35840=>"101000011",
  35841=>"011111110",
  35842=>"100100100",
  35843=>"011100100",
  35844=>"000110111",
  35845=>"111010010",
  35846=>"101100101",
  35847=>"011011111",
  35848=>"100111011",
  35849=>"001111010",
  35850=>"100001011",
  35851=>"010111011",
  35852=>"111001101",
  35853=>"000000101",
  35854=>"111011101",
  35855=>"101001010",
  35856=>"000111110",
  35857=>"001000001",
  35858=>"100011110",
  35859=>"101101111",
  35860=>"010000000",
  35861=>"111010100",
  35862=>"111100011",
  35863=>"000010000",
  35864=>"110001111",
  35865=>"000000000",
  35866=>"011111011",
  35867=>"000111111",
  35868=>"110101101",
  35869=>"000010110",
  35870=>"110001110",
  35871=>"010110000",
  35872=>"110111111",
  35873=>"010101111",
  35874=>"001111110",
  35875=>"110000100",
  35876=>"001011111",
  35877=>"001010111",
  35878=>"111000010",
  35879=>"110111100",
  35880=>"011111010",
  35881=>"000001010",
  35882=>"110111111",
  35883=>"001100011",
  35884=>"100110100",
  35885=>"100010001",
  35886=>"000111111",
  35887=>"010001101",
  35888=>"101111111",
  35889=>"101101111",
  35890=>"001010001",
  35891=>"111110111",
  35892=>"101000010",
  35893=>"100001101",
  35894=>"100100000",
  35895=>"101110001",
  35896=>"000001111",
  35897=>"001100010",
  35898=>"001011001",
  35899=>"100000111",
  35900=>"011111110",
  35901=>"001100010",
  35902=>"001011000",
  35903=>"010001101",
  35904=>"110111110",
  35905=>"101000110",
  35906=>"110101011",
  35907=>"101101011",
  35908=>"100100101",
  35909=>"101010010",
  35910=>"110110110",
  35911=>"100011010",
  35912=>"110110010",
  35913=>"011110111",
  35914=>"001111101",
  35915=>"000100001",
  35916=>"001111000",
  35917=>"000001100",
  35918=>"011110001",
  35919=>"101110001",
  35920=>"101110011",
  35921=>"000010110",
  35922=>"100010000",
  35923=>"000110110",
  35924=>"101111010",
  35925=>"111100111",
  35926=>"010010100",
  35927=>"001011000",
  35928=>"000010010",
  35929=>"110101100",
  35930=>"001101010",
  35931=>"011000000",
  35932=>"001000011",
  35933=>"001011000",
  35934=>"101001100",
  35935=>"010011101",
  35936=>"000010011",
  35937=>"110111011",
  35938=>"010011011",
  35939=>"111100011",
  35940=>"101011100",
  35941=>"110010101",
  35942=>"111011101",
  35943=>"001111101",
  35944=>"000110000",
  35945=>"011000011",
  35946=>"101000000",
  35947=>"011101001",
  35948=>"001101111",
  35949=>"110110001",
  35950=>"110111010",
  35951=>"000101110",
  35952=>"111111100",
  35953=>"011001000",
  35954=>"011111010",
  35955=>"110001110",
  35956=>"110101000",
  35957=>"110011100",
  35958=>"101000011",
  35959=>"100011001",
  35960=>"010011111",
  35961=>"010001001",
  35962=>"110010011",
  35963=>"000001010",
  35964=>"001000010",
  35965=>"001001000",
  35966=>"110110110",
  35967=>"101110111",
  35968=>"011100110",
  35969=>"000111111",
  35970=>"001000001",
  35971=>"111101101",
  35972=>"100110000",
  35973=>"001100011",
  35974=>"111110101",
  35975=>"001001111",
  35976=>"011101110",
  35977=>"101001000",
  35978=>"111010010",
  35979=>"010110000",
  35980=>"010011000",
  35981=>"000111001",
  35982=>"100101010",
  35983=>"100100101",
  35984=>"111110110",
  35985=>"110101001",
  35986=>"101011000",
  35987=>"001011011",
  35988=>"110111011",
  35989=>"100101001",
  35990=>"010001100",
  35991=>"001110110",
  35992=>"100110010",
  35993=>"111000010",
  35994=>"100011111",
  35995=>"011000000",
  35996=>"111111110",
  35997=>"100001100",
  35998=>"001100011",
  35999=>"010101101",
  36000=>"011111010",
  36001=>"100000001",
  36002=>"110101100",
  36003=>"010000111",
  36004=>"100111000",
  36005=>"101111111",
  36006=>"100101010",
  36007=>"010000101",
  36008=>"110010000",
  36009=>"101111110",
  36010=>"100111100",
  36011=>"111110111",
  36012=>"010010010",
  36013=>"001110111",
  36014=>"000101101",
  36015=>"000010011",
  36016=>"000011011",
  36017=>"001010001",
  36018=>"001100111",
  36019=>"110011110",
  36020=>"001000010",
  36021=>"100000000",
  36022=>"101000111",
  36023=>"001011000",
  36024=>"110010001",
  36025=>"110000101",
  36026=>"000011101",
  36027=>"100010011",
  36028=>"110000100",
  36029=>"111100011",
  36030=>"111100001",
  36031=>"000000000",
  36032=>"001110111",
  36033=>"100101000",
  36034=>"000001001",
  36035=>"111111101",
  36036=>"111110001",
  36037=>"111000111",
  36038=>"000011100",
  36039=>"100100111",
  36040=>"010010010",
  36041=>"000110001",
  36042=>"000010100",
  36043=>"100110111",
  36044=>"111001000",
  36045=>"101001011",
  36046=>"001110001",
  36047=>"001111001",
  36048=>"011110000",
  36049=>"100010010",
  36050=>"110100010",
  36051=>"010111101",
  36052=>"101000010",
  36053=>"101101111",
  36054=>"001001100",
  36055=>"110010011",
  36056=>"000111001",
  36057=>"001101010",
  36058=>"010000111",
  36059=>"100010100",
  36060=>"111011110",
  36061=>"110000000",
  36062=>"111001111",
  36063=>"011101011",
  36064=>"011100000",
  36065=>"010110001",
  36066=>"101111100",
  36067=>"001010100",
  36068=>"110010101",
  36069=>"011111100",
  36070=>"111101001",
  36071=>"111011100",
  36072=>"011110011",
  36073=>"111000111",
  36074=>"011000110",
  36075=>"010111001",
  36076=>"010001110",
  36077=>"001111010",
  36078=>"110101000",
  36079=>"001110000",
  36080=>"000010000",
  36081=>"110000000",
  36082=>"111100110",
  36083=>"100100111",
  36084=>"010010101",
  36085=>"110000000",
  36086=>"010000111",
  36087=>"000000011",
  36088=>"011001111",
  36089=>"001001111",
  36090=>"101100101",
  36091=>"101000111",
  36092=>"011111100",
  36093=>"011110100",
  36094=>"111110011",
  36095=>"100101101",
  36096=>"011110010",
  36097=>"000100011",
  36098=>"100110111",
  36099=>"101000000",
  36100=>"101111110",
  36101=>"001011101",
  36102=>"011101010",
  36103=>"100110010",
  36104=>"011111111",
  36105=>"000001000",
  36106=>"110001000",
  36107=>"011100010",
  36108=>"000110001",
  36109=>"010001111",
  36110=>"010101011",
  36111=>"111010010",
  36112=>"111111100",
  36113=>"111111111",
  36114=>"010010011",
  36115=>"001010111",
  36116=>"111001110",
  36117=>"101001100",
  36118=>"100110000",
  36119=>"001000101",
  36120=>"110110110",
  36121=>"011100100",
  36122=>"100100000",
  36123=>"101011010",
  36124=>"110101110",
  36125=>"010001011",
  36126=>"100001111",
  36127=>"000000010",
  36128=>"101000000",
  36129=>"110111010",
  36130=>"011110001",
  36131=>"000001001",
  36132=>"010110001",
  36133=>"111010101",
  36134=>"101100011",
  36135=>"000111100",
  36136=>"111110010",
  36137=>"110111100",
  36138=>"100010111",
  36139=>"000101001",
  36140=>"010001011",
  36141=>"001010110",
  36142=>"111100101",
  36143=>"111010110",
  36144=>"101011001",
  36145=>"110100100",
  36146=>"111010100",
  36147=>"111000111",
  36148=>"100011110",
  36149=>"101000100",
  36150=>"000001000",
  36151=>"100010000",
  36152=>"011110100",
  36153=>"011011001",
  36154=>"001101011",
  36155=>"000100001",
  36156=>"101001111",
  36157=>"001011111",
  36158=>"110110100",
  36159=>"110110111",
  36160=>"011011000",
  36161=>"010000101",
  36162=>"000100101",
  36163=>"111000010",
  36164=>"110110110",
  36165=>"111111111",
  36166=>"110101000",
  36167=>"100000010",
  36168=>"111110001",
  36169=>"010000010",
  36170=>"001111100",
  36171=>"100101000",
  36172=>"100011110",
  36173=>"110011001",
  36174=>"001100100",
  36175=>"110111110",
  36176=>"111001101",
  36177=>"011100100",
  36178=>"100011101",
  36179=>"110101101",
  36180=>"000100001",
  36181=>"111111000",
  36182=>"110100101",
  36183=>"010000010",
  36184=>"001111110",
  36185=>"011011100",
  36186=>"101011011",
  36187=>"110100110",
  36188=>"011101101",
  36189=>"010000010",
  36190=>"001011011",
  36191=>"000000000",
  36192=>"011101110",
  36193=>"010010010",
  36194=>"101001100",
  36195=>"010010010",
  36196=>"101011110",
  36197=>"110011101",
  36198=>"100001111",
  36199=>"110011110",
  36200=>"101101000",
  36201=>"100111011",
  36202=>"100100101",
  36203=>"000011000",
  36204=>"011111001",
  36205=>"101101011",
  36206=>"011100001",
  36207=>"010111000",
  36208=>"011010100",
  36209=>"000101100",
  36210=>"100110101",
  36211=>"110010111",
  36212=>"110000000",
  36213=>"000111011",
  36214=>"001001101",
  36215=>"101101101",
  36216=>"010000110",
  36217=>"011100110",
  36218=>"001011101",
  36219=>"000000000",
  36220=>"000001100",
  36221=>"011001100",
  36222=>"101111110",
  36223=>"110000011",
  36224=>"010011110",
  36225=>"011010011",
  36226=>"011011111",
  36227=>"000000001",
  36228=>"001101100",
  36229=>"110101000",
  36230=>"001011100",
  36231=>"110110010",
  36232=>"001100110",
  36233=>"000001100",
  36234=>"100110011",
  36235=>"110110000",
  36236=>"010011011",
  36237=>"110100100",
  36238=>"101010010",
  36239=>"101000000",
  36240=>"000010111",
  36241=>"111001101",
  36242=>"000000110",
  36243=>"000111110",
  36244=>"101000011",
  36245=>"100101010",
  36246=>"011010111",
  36247=>"011100010",
  36248=>"110110001",
  36249=>"010011001",
  36250=>"010100011",
  36251=>"100000011",
  36252=>"100000011",
  36253=>"011011010",
  36254=>"100110001",
  36255=>"000010110",
  36256=>"101101101",
  36257=>"011011011",
  36258=>"011000010",
  36259=>"000000011",
  36260=>"000001110",
  36261=>"110110111",
  36262=>"100010010",
  36263=>"000000101",
  36264=>"001001010",
  36265=>"000100011",
  36266=>"011000001",
  36267=>"110001101",
  36268=>"000100111",
  36269=>"010001100",
  36270=>"001010000",
  36271=>"000111010",
  36272=>"101100000",
  36273=>"000001110",
  36274=>"001000100",
  36275=>"001000001",
  36276=>"110111011",
  36277=>"110010011",
  36278=>"001110101",
  36279=>"111000111",
  36280=>"001010100",
  36281=>"000011011",
  36282=>"001001111",
  36283=>"011001101",
  36284=>"101110010",
  36285=>"101110110",
  36286=>"010101101",
  36287=>"000110011",
  36288=>"111011001",
  36289=>"010100000",
  36290=>"010111000",
  36291=>"001010010",
  36292=>"100000000",
  36293=>"101100001",
  36294=>"101010101",
  36295=>"101101100",
  36296=>"001110110",
  36297=>"011001101",
  36298=>"011101110",
  36299=>"001111111",
  36300=>"101010111",
  36301=>"000001001",
  36302=>"111000001",
  36303=>"010001001",
  36304=>"100111010",
  36305=>"101101101",
  36306=>"110111110",
  36307=>"001001010",
  36308=>"111111011",
  36309=>"000000010",
  36310=>"001110010",
  36311=>"000110001",
  36312=>"000011101",
  36313=>"111100111",
  36314=>"000111011",
  36315=>"001001100",
  36316=>"111100001",
  36317=>"001101101",
  36318=>"001010000",
  36319=>"001110001",
  36320=>"111000101",
  36321=>"101010011",
  36322=>"011000111",
  36323=>"001000000",
  36324=>"111001011",
  36325=>"011110101",
  36326=>"101101001",
  36327=>"100001111",
  36328=>"010010011",
  36329=>"110010100",
  36330=>"110001101",
  36331=>"000001101",
  36332=>"100110101",
  36333=>"000011100",
  36334=>"001000111",
  36335=>"000000111",
  36336=>"110010100",
  36337=>"011101111",
  36338=>"100011001",
  36339=>"011010000",
  36340=>"101111000",
  36341=>"010001111",
  36342=>"111011000",
  36343=>"000100101",
  36344=>"110111000",
  36345=>"111000110",
  36346=>"100001011",
  36347=>"000011011",
  36348=>"011110011",
  36349=>"110111011",
  36350=>"000111001",
  36351=>"111000000",
  36352=>"010100001",
  36353=>"100101000",
  36354=>"001100010",
  36355=>"111010011",
  36356=>"011101000",
  36357=>"000111000",
  36358=>"111110110",
  36359=>"001111000",
  36360=>"001010110",
  36361=>"110100101",
  36362=>"111111100",
  36363=>"000110000",
  36364=>"001010010",
  36365=>"100110011",
  36366=>"101000100",
  36367=>"010111001",
  36368=>"011110011",
  36369=>"000100100",
  36370=>"011100010",
  36371=>"110111111",
  36372=>"100110001",
  36373=>"000001100",
  36374=>"000110111",
  36375=>"110110001",
  36376=>"110001110",
  36377=>"110110000",
  36378=>"011000000",
  36379=>"010010100",
  36380=>"011000001",
  36381=>"100101000",
  36382=>"001011110",
  36383=>"100010110",
  36384=>"001000011",
  36385=>"010110001",
  36386=>"111110111",
  36387=>"111011010",
  36388=>"001001000",
  36389=>"110000011",
  36390=>"111011001",
  36391=>"011011010",
  36392=>"100010100",
  36393=>"110110001",
  36394=>"000100000",
  36395=>"010000011",
  36396=>"000101011",
  36397=>"010010011",
  36398=>"100100000",
  36399=>"011010010",
  36400=>"011101101",
  36401=>"000001111",
  36402=>"110001111",
  36403=>"111001111",
  36404=>"111000100",
  36405=>"000010110",
  36406=>"011001111",
  36407=>"001010011",
  36408=>"000110011",
  36409=>"001110111",
  36410=>"010001001",
  36411=>"101110101",
  36412=>"011000100",
  36413=>"111111001",
  36414=>"001100001",
  36415=>"110101101",
  36416=>"110111111",
  36417=>"001000011",
  36418=>"001011001",
  36419=>"001101101",
  36420=>"101111111",
  36421=>"101001101",
  36422=>"001100100",
  36423=>"101101101",
  36424=>"000000101",
  36425=>"101100001",
  36426=>"100001111",
  36427=>"100011010",
  36428=>"110101001",
  36429=>"100100001",
  36430=>"000000001",
  36431=>"001001111",
  36432=>"110111110",
  36433=>"010010110",
  36434=>"011111101",
  36435=>"110000001",
  36436=>"000010100",
  36437=>"101000100",
  36438=>"001001111",
  36439=>"001011111",
  36440=>"110110100",
  36441=>"101010001",
  36442=>"101100001",
  36443=>"011000000",
  36444=>"011011110",
  36445=>"000010101",
  36446=>"100000001",
  36447=>"101111100",
  36448=>"110000101",
  36449=>"010010101",
  36450=>"100001000",
  36451=>"011100011",
  36452=>"000010000",
  36453=>"011000010",
  36454=>"010101100",
  36455=>"111110110",
  36456=>"110001110",
  36457=>"111011000",
  36458=>"001011111",
  36459=>"101100111",
  36460=>"001001001",
  36461=>"010111000",
  36462=>"011111111",
  36463=>"110000010",
  36464=>"001110001",
  36465=>"000001010",
  36466=>"011010001",
  36467=>"111010111",
  36468=>"110000010",
  36469=>"000100011",
  36470=>"101100001",
  36471=>"111110100",
  36472=>"010100001",
  36473=>"011101101",
  36474=>"100000111",
  36475=>"111001011",
  36476=>"101110011",
  36477=>"001010101",
  36478=>"101100000",
  36479=>"110101110",
  36480=>"111111001",
  36481=>"110000110",
  36482=>"111010111",
  36483=>"010011110",
  36484=>"111110110",
  36485=>"101100000",
  36486=>"011111011",
  36487=>"110000010",
  36488=>"100101101",
  36489=>"010111111",
  36490=>"111110101",
  36491=>"110101001",
  36492=>"100110100",
  36493=>"110000110",
  36494=>"100001110",
  36495=>"111111100",
  36496=>"001111011",
  36497=>"001001010",
  36498=>"010010001",
  36499=>"100010001",
  36500=>"101110000",
  36501=>"010111100",
  36502=>"101000101",
  36503=>"101100101",
  36504=>"110011001",
  36505=>"110000000",
  36506=>"111010111",
  36507=>"101111110",
  36508=>"101011111",
  36509=>"110000010",
  36510=>"111010001",
  36511=>"101101011",
  36512=>"000111001",
  36513=>"011100000",
  36514=>"010010111",
  36515=>"100000110",
  36516=>"011000111",
  36517=>"001100111",
  36518=>"000100001",
  36519=>"011001000",
  36520=>"000000100",
  36521=>"010000000",
  36522=>"101111110",
  36523=>"111101110",
  36524=>"010011110",
  36525=>"100000000",
  36526=>"110101000",
  36527=>"011000000",
  36528=>"010000011",
  36529=>"111000100",
  36530=>"101001001",
  36531=>"110011101",
  36532=>"101101110",
  36533=>"001111100",
  36534=>"010010010",
  36535=>"000000111",
  36536=>"110011010",
  36537=>"001011110",
  36538=>"010010010",
  36539=>"110001100",
  36540=>"011111101",
  36541=>"011000101",
  36542=>"000000010",
  36543=>"000001001",
  36544=>"010110001",
  36545=>"111010011",
  36546=>"000101111",
  36547=>"100001101",
  36548=>"000100101",
  36549=>"000111101",
  36550=>"010000001",
  36551=>"101101101",
  36552=>"111110101",
  36553=>"001001110",
  36554=>"011111101",
  36555=>"010111101",
  36556=>"100110011",
  36557=>"001000011",
  36558=>"011011011",
  36559=>"001100111",
  36560=>"010000101",
  36561=>"111110000",
  36562=>"001000000",
  36563=>"000100010",
  36564=>"100101001",
  36565=>"010000001",
  36566=>"101001010",
  36567=>"010011000",
  36568=>"000011000",
  36569=>"110001000",
  36570=>"001101110",
  36571=>"001001011",
  36572=>"111101000",
  36573=>"111001100",
  36574=>"010100010",
  36575=>"001110110",
  36576=>"111001110",
  36577=>"100011100",
  36578=>"011010001",
  36579=>"100110101",
  36580=>"010111111",
  36581=>"111110101",
  36582=>"100011110",
  36583=>"110110101",
  36584=>"100010010",
  36585=>"110111111",
  36586=>"010111101",
  36587=>"100100110",
  36588=>"000100011",
  36589=>"111101111",
  36590=>"111111111",
  36591=>"000011010",
  36592=>"000100111",
  36593=>"010110100",
  36594=>"011101101",
  36595=>"111001000",
  36596=>"101010010",
  36597=>"110000110",
  36598=>"111111000",
  36599=>"011000000",
  36600=>"110010010",
  36601=>"110000110",
  36602=>"000111111",
  36603=>"111011110",
  36604=>"110000001",
  36605=>"101111000",
  36606=>"110010001",
  36607=>"111000000",
  36608=>"110111000",
  36609=>"001100110",
  36610=>"100101110",
  36611=>"100000110",
  36612=>"101000100",
  36613=>"111110001",
  36614=>"010111110",
  36615=>"100100001",
  36616=>"001111110",
  36617=>"000001111",
  36618=>"011000110",
  36619=>"101010011",
  36620=>"011101100",
  36621=>"101000011",
  36622=>"001000011",
  36623=>"101001011",
  36624=>"111100110",
  36625=>"001000010",
  36626=>"101110001",
  36627=>"110000001",
  36628=>"001111110",
  36629=>"000110101",
  36630=>"100011001",
  36631=>"000010000",
  36632=>"110001000",
  36633=>"100101100",
  36634=>"011000001",
  36635=>"000001000",
  36636=>"111010000",
  36637=>"110100010",
  36638=>"001111010",
  36639=>"110110110",
  36640=>"101100111",
  36641=>"011000000",
  36642=>"100110010",
  36643=>"111100000",
  36644=>"001110101",
  36645=>"000001010",
  36646=>"100101110",
  36647=>"100001101",
  36648=>"010011101",
  36649=>"111001100",
  36650=>"110110011",
  36651=>"101011100",
  36652=>"110101000",
  36653=>"000011000",
  36654=>"100001011",
  36655=>"101001011",
  36656=>"000100110",
  36657=>"110001110",
  36658=>"111110000",
  36659=>"000000010",
  36660=>"111101010",
  36661=>"011101110",
  36662=>"000011010",
  36663=>"000101100",
  36664=>"000111000",
  36665=>"100110011",
  36666=>"001000010",
  36667=>"101000000",
  36668=>"011101001",
  36669=>"011011010",
  36670=>"001100001",
  36671=>"010010110",
  36672=>"111100101",
  36673=>"001111101",
  36674=>"110111101",
  36675=>"101010001",
  36676=>"101010001",
  36677=>"110111101",
  36678=>"101101011",
  36679=>"111101010",
  36680=>"101101110",
  36681=>"000011001",
  36682=>"011001011",
  36683=>"001101011",
  36684=>"111111000",
  36685=>"001010110",
  36686=>"000001011",
  36687=>"101101100",
  36688=>"110110001",
  36689=>"001110111",
  36690=>"111111110",
  36691=>"000010000",
  36692=>"100101010",
  36693=>"110011001",
  36694=>"011010101",
  36695=>"010101101",
  36696=>"111001000",
  36697=>"010010100",
  36698=>"110111101",
  36699=>"011100000",
  36700=>"111101010",
  36701=>"001000000",
  36702=>"110110110",
  36703=>"000010000",
  36704=>"100010111",
  36705=>"001001001",
  36706=>"010110000",
  36707=>"011100101",
  36708=>"001000000",
  36709=>"110100110",
  36710=>"010000100",
  36711=>"111100100",
  36712=>"111111000",
  36713=>"010010000",
  36714=>"010010001",
  36715=>"101010110",
  36716=>"111100011",
  36717=>"001111000",
  36718=>"000001100",
  36719=>"100010110",
  36720=>"010001111",
  36721=>"011001111",
  36722=>"111001001",
  36723=>"101000110",
  36724=>"110110100",
  36725=>"000110001",
  36726=>"010000101",
  36727=>"011110111",
  36728=>"111011011",
  36729=>"000010010",
  36730=>"101101010",
  36731=>"010000110",
  36732=>"111010111",
  36733=>"101001110",
  36734=>"100111110",
  36735=>"011101110",
  36736=>"100100010",
  36737=>"011000011",
  36738=>"111001010",
  36739=>"101000001",
  36740=>"000001001",
  36741=>"111010110",
  36742=>"010011110",
  36743=>"010100001",
  36744=>"110101001",
  36745=>"100000101",
  36746=>"001000100",
  36747=>"111110111",
  36748=>"011101000",
  36749=>"000000010",
  36750=>"101101011",
  36751=>"100001100",
  36752=>"110100001",
  36753=>"101110110",
  36754=>"001111110",
  36755=>"110011111",
  36756=>"110100010",
  36757=>"101110111",
  36758=>"111011111",
  36759=>"000001111",
  36760=>"011000000",
  36761=>"001010011",
  36762=>"111010010",
  36763=>"100101110",
  36764=>"110000100",
  36765=>"001000001",
  36766=>"001100011",
  36767=>"110001010",
  36768=>"100101001",
  36769=>"011000111",
  36770=>"110111111",
  36771=>"100111011",
  36772=>"100111111",
  36773=>"111010100",
  36774=>"111010001",
  36775=>"011101011",
  36776=>"000100010",
  36777=>"011001001",
  36778=>"011010100",
  36779=>"110011000",
  36780=>"000101101",
  36781=>"010010000",
  36782=>"101110001",
  36783=>"000010111",
  36784=>"010010011",
  36785=>"000010101",
  36786=>"000110000",
  36787=>"110101000",
  36788=>"010010011",
  36789=>"110111110",
  36790=>"001100010",
  36791=>"101001000",
  36792=>"110000111",
  36793=>"001111011",
  36794=>"001001011",
  36795=>"100010000",
  36796=>"010001010",
  36797=>"100101000",
  36798=>"101100101",
  36799=>"000000110",
  36800=>"110110001",
  36801=>"101100110",
  36802=>"111110101",
  36803=>"100000101",
  36804=>"110100101",
  36805=>"101110111",
  36806=>"100100101",
  36807=>"110101110",
  36808=>"000110010",
  36809=>"011011000",
  36810=>"010111110",
  36811=>"100111111",
  36812=>"110101000",
  36813=>"100100100",
  36814=>"010101011",
  36815=>"010100000",
  36816=>"111001110",
  36817=>"000000110",
  36818=>"010100101",
  36819=>"000100000",
  36820=>"001010010",
  36821=>"110110010",
  36822=>"011110000",
  36823=>"111110011",
  36824=>"101110110",
  36825=>"011100011",
  36826=>"000011000",
  36827=>"110111001",
  36828=>"100100110",
  36829=>"111111100",
  36830=>"111100011",
  36831=>"100100111",
  36832=>"010000011",
  36833=>"100011110",
  36834=>"011010010",
  36835=>"110001011",
  36836=>"000000010",
  36837=>"010001001",
  36838=>"000111110",
  36839=>"001001010",
  36840=>"111001101",
  36841=>"001010011",
  36842=>"010110001",
  36843=>"100100111",
  36844=>"101000000",
  36845=>"011110001",
  36846=>"001000101",
  36847=>"000100111",
  36848=>"110111011",
  36849=>"011000001",
  36850=>"111001101",
  36851=>"010010000",
  36852=>"010101110",
  36853=>"000110101",
  36854=>"110000101",
  36855=>"000010011",
  36856=>"001111000",
  36857=>"100010101",
  36858=>"101101001",
  36859=>"110111010",
  36860=>"111101001",
  36861=>"010110100",
  36862=>"011100110",
  36863=>"111111010",
  36864=>"011100001",
  36865=>"000001000",
  36866=>"000110111",
  36867=>"000100001",
  36868=>"001000101",
  36869=>"101010010",
  36870=>"001111010",
  36871=>"010101110",
  36872=>"110100000",
  36873=>"001101001",
  36874=>"000010000",
  36875=>"101100010",
  36876=>"000111001",
  36877=>"010110011",
  36878=>"000010011",
  36879=>"010100010",
  36880=>"110101101",
  36881=>"000110100",
  36882=>"011101001",
  36883=>"001001101",
  36884=>"110011010",
  36885=>"100110100",
  36886=>"011010101",
  36887=>"000000000",
  36888=>"111100001",
  36889=>"010101001",
  36890=>"100110111",
  36891=>"010001100",
  36892=>"000110011",
  36893=>"101110101",
  36894=>"110011100",
  36895=>"100101110",
  36896=>"100011011",
  36897=>"001101001",
  36898=>"101010010",
  36899=>"100010100",
  36900=>"001101100",
  36901=>"001101101",
  36902=>"110100111",
  36903=>"011010111",
  36904=>"101101000",
  36905=>"010101100",
  36906=>"111101101",
  36907=>"110011101",
  36908=>"111111111",
  36909=>"111111101",
  36910=>"010010011",
  36911=>"010100100",
  36912=>"101010110",
  36913=>"000000010",
  36914=>"010011011",
  36915=>"110100010",
  36916=>"011110111",
  36917=>"110100100",
  36918=>"110001110",
  36919=>"111011010",
  36920=>"010000001",
  36921=>"111101111",
  36922=>"001101100",
  36923=>"010010101",
  36924=>"101000010",
  36925=>"111100111",
  36926=>"111011111",
  36927=>"011010110",
  36928=>"001010111",
  36929=>"101001001",
  36930=>"110001111",
  36931=>"100001110",
  36932=>"001110001",
  36933=>"011100010",
  36934=>"010111011",
  36935=>"110111100",
  36936=>"011110011",
  36937=>"110010101",
  36938=>"001010110",
  36939=>"000010010",
  36940=>"101001111",
  36941=>"000011101",
  36942=>"011000111",
  36943=>"011101101",
  36944=>"000101000",
  36945=>"001001001",
  36946=>"101110001",
  36947=>"110101000",
  36948=>"101011100",
  36949=>"111110001",
  36950=>"000000001",
  36951=>"101011001",
  36952=>"001111000",
  36953=>"000010111",
  36954=>"111011101",
  36955=>"101111111",
  36956=>"001010111",
  36957=>"000010100",
  36958=>"100101011",
  36959=>"000111101",
  36960=>"101001111",
  36961=>"100000000",
  36962=>"000011001",
  36963=>"111111110",
  36964=>"001000111",
  36965=>"011100111",
  36966=>"110100101",
  36967=>"000101110",
  36968=>"111101000",
  36969=>"000010110",
  36970=>"101010110",
  36971=>"101001100",
  36972=>"100110001",
  36973=>"111011110",
  36974=>"010111110",
  36975=>"010010000",
  36976=>"111110011",
  36977=>"111000110",
  36978=>"000000101",
  36979=>"010000101",
  36980=>"001101011",
  36981=>"111101011",
  36982=>"000101011",
  36983=>"010011001",
  36984=>"010100000",
  36985=>"000000001",
  36986=>"111110001",
  36987=>"110110110",
  36988=>"001001100",
  36989=>"111000110",
  36990=>"010011000",
  36991=>"110110001",
  36992=>"110111000",
  36993=>"101101011",
  36994=>"100001101",
  36995=>"011001001",
  36996=>"010010011",
  36997=>"000100011",
  36998=>"010110100",
  36999=>"001000011",
  37000=>"110001111",
  37001=>"101100010",
  37002=>"000110011",
  37003=>"010000011",
  37004=>"000000100",
  37005=>"100001001",
  37006=>"001011111",
  37007=>"001111001",
  37008=>"000010101",
  37009=>"101010111",
  37010=>"000001100",
  37011=>"101011001",
  37012=>"111101000",
  37013=>"100101011",
  37014=>"101010001",
  37015=>"110001011",
  37016=>"000100111",
  37017=>"110000110",
  37018=>"000010000",
  37019=>"110101110",
  37020=>"001100001",
  37021=>"111111011",
  37022=>"011110001",
  37023=>"100100001",
  37024=>"110101100",
  37025=>"001000101",
  37026=>"000000110",
  37027=>"001000001",
  37028=>"111100111",
  37029=>"101111001",
  37030=>"111110111",
  37031=>"101011011",
  37032=>"000101000",
  37033=>"010101001",
  37034=>"110010000",
  37035=>"111001111",
  37036=>"000011111",
  37037=>"001010101",
  37038=>"000101011",
  37039=>"111100111",
  37040=>"000000000",
  37041=>"101000110",
  37042=>"111011101",
  37043=>"100110101",
  37044=>"100110100",
  37045=>"010100001",
  37046=>"110110110",
  37047=>"011111110",
  37048=>"011010100",
  37049=>"111011001",
  37050=>"100101001",
  37051=>"100000110",
  37052=>"000111101",
  37053=>"001011010",
  37054=>"010110010",
  37055=>"111001111",
  37056=>"111001101",
  37057=>"111111111",
  37058=>"111011110",
  37059=>"111110110",
  37060=>"111110100",
  37061=>"001001100",
  37062=>"000110001",
  37063=>"001101000",
  37064=>"011101100",
  37065=>"100110010",
  37066=>"110000110",
  37067=>"011000010",
  37068=>"111100000",
  37069=>"000110100",
  37070=>"011111101",
  37071=>"001000001",
  37072=>"100110000",
  37073=>"000010100",
  37074=>"111011000",
  37075=>"000001011",
  37076=>"101001101",
  37077=>"010001101",
  37078=>"101010100",
  37079=>"110111101",
  37080=>"101100100",
  37081=>"011000011",
  37082=>"100001111",
  37083=>"111011101",
  37084=>"101010111",
  37085=>"111111010",
  37086=>"011110110",
  37087=>"011011110",
  37088=>"100000101",
  37089=>"000110100",
  37090=>"010001100",
  37091=>"110010001",
  37092=>"000011111",
  37093=>"110010000",
  37094=>"000000100",
  37095=>"100110001",
  37096=>"111111111",
  37097=>"110001111",
  37098=>"101001010",
  37099=>"110010000",
  37100=>"100000100",
  37101=>"011111111",
  37102=>"001101001",
  37103=>"100010001",
  37104=>"010111011",
  37105=>"000111110",
  37106=>"000010000",
  37107=>"100111001",
  37108=>"010011011",
  37109=>"000010110",
  37110=>"001001011",
  37111=>"011100011",
  37112=>"010011110",
  37113=>"000111010",
  37114=>"100001000",
  37115=>"110001001",
  37116=>"111001110",
  37117=>"000100111",
  37118=>"111101111",
  37119=>"001011100",
  37120=>"010110100",
  37121=>"001111111",
  37122=>"011101111",
  37123=>"101101100",
  37124=>"101000111",
  37125=>"011010111",
  37126=>"000100101",
  37127=>"111111111",
  37128=>"111100100",
  37129=>"101000001",
  37130=>"001101001",
  37131=>"110110010",
  37132=>"111101111",
  37133=>"010000111",
  37134=>"101000111",
  37135=>"000110010",
  37136=>"110101100",
  37137=>"001110110",
  37138=>"000010000",
  37139=>"010101111",
  37140=>"110110111",
  37141=>"011111110",
  37142=>"011000000",
  37143=>"001110110",
  37144=>"010100000",
  37145=>"000000111",
  37146=>"011000010",
  37147=>"110111011",
  37148=>"101111010",
  37149=>"110110100",
  37150=>"101111111",
  37151=>"101100001",
  37152=>"001100101",
  37153=>"111111110",
  37154=>"011011111",
  37155=>"011101110",
  37156=>"010100111",
  37157=>"111110100",
  37158=>"111000011",
  37159=>"100110000",
  37160=>"000011011",
  37161=>"001101101",
  37162=>"011110011",
  37163=>"110100111",
  37164=>"111000110",
  37165=>"111010011",
  37166=>"000110001",
  37167=>"001011110",
  37168=>"111101011",
  37169=>"010001010",
  37170=>"110101110",
  37171=>"100100101",
  37172=>"011001111",
  37173=>"011001110",
  37174=>"011110011",
  37175=>"011000000",
  37176=>"111111100",
  37177=>"110111011",
  37178=>"111011000",
  37179=>"000000010",
  37180=>"110101111",
  37181=>"100011001",
  37182=>"000000101",
  37183=>"000010010",
  37184=>"001101001",
  37185=>"001000010",
  37186=>"100100110",
  37187=>"110111111",
  37188=>"100001000",
  37189=>"101111010",
  37190=>"001110110",
  37191=>"100000001",
  37192=>"000011101",
  37193=>"111000100",
  37194=>"101010101",
  37195=>"010010001",
  37196=>"010111100",
  37197=>"100100110",
  37198=>"100000111",
  37199=>"100100101",
  37200=>"111111100",
  37201=>"010111100",
  37202=>"111110100",
  37203=>"100110101",
  37204=>"100011101",
  37205=>"001111010",
  37206=>"111111011",
  37207=>"001100100",
  37208=>"110100010",
  37209=>"000001001",
  37210=>"100001001",
  37211=>"101101111",
  37212=>"000100111",
  37213=>"110010111",
  37214=>"000110001",
  37215=>"000010111",
  37216=>"011001011",
  37217=>"100000011",
  37218=>"100100010",
  37219=>"001010010",
  37220=>"101011010",
  37221=>"011010101",
  37222=>"001010111",
  37223=>"011001000",
  37224=>"111101100",
  37225=>"101001111",
  37226=>"100110011",
  37227=>"111110110",
  37228=>"000100000",
  37229=>"101010001",
  37230=>"011100100",
  37231=>"001110100",
  37232=>"100011011",
  37233=>"110001000",
  37234=>"110110111",
  37235=>"100100110",
  37236=>"000011010",
  37237=>"011000100",
  37238=>"011011000",
  37239=>"111101101",
  37240=>"000110001",
  37241=>"001101000",
  37242=>"010100010",
  37243=>"111000100",
  37244=>"100000010",
  37245=>"101111101",
  37246=>"010100010",
  37247=>"001010110",
  37248=>"110011000",
  37249=>"100000110",
  37250=>"011001100",
  37251=>"101000010",
  37252=>"110110001",
  37253=>"010101000",
  37254=>"001110010",
  37255=>"101110010",
  37256=>"000100100",
  37257=>"110000100",
  37258=>"100001101",
  37259=>"000011010",
  37260=>"110110010",
  37261=>"010111010",
  37262=>"111010001",
  37263=>"101110010",
  37264=>"000101111",
  37265=>"110111001",
  37266=>"001011011",
  37267=>"000100101",
  37268=>"100110011",
  37269=>"001010001",
  37270=>"101011100",
  37271=>"111001001",
  37272=>"001001001",
  37273=>"001001100",
  37274=>"100010111",
  37275=>"100011011",
  37276=>"001101001",
  37277=>"101000101",
  37278=>"101110101",
  37279=>"111001100",
  37280=>"100101001",
  37281=>"100001010",
  37282=>"011100111",
  37283=>"101110011",
  37284=>"110100000",
  37285=>"111010011",
  37286=>"011000111",
  37287=>"010110111",
  37288=>"000110101",
  37289=>"001100111",
  37290=>"000110000",
  37291=>"100000110",
  37292=>"110111100",
  37293=>"010111000",
  37294=>"010100111",
  37295=>"010011111",
  37296=>"101001011",
  37297=>"111000111",
  37298=>"011100101",
  37299=>"100010010",
  37300=>"110011011",
  37301=>"111111001",
  37302=>"000110110",
  37303=>"001101111",
  37304=>"001010001",
  37305=>"101000101",
  37306=>"001001001",
  37307=>"011101100",
  37308=>"111010001",
  37309=>"010010001",
  37310=>"100101101",
  37311=>"100000000",
  37312=>"010100111",
  37313=>"011010000",
  37314=>"110111000",
  37315=>"000100101",
  37316=>"000011010",
  37317=>"111110010",
  37318=>"000000100",
  37319=>"111001010",
  37320=>"000101001",
  37321=>"000010111",
  37322=>"000010111",
  37323=>"100011000",
  37324=>"000110001",
  37325=>"111100011",
  37326=>"111010111",
  37327=>"011001100",
  37328=>"110110001",
  37329=>"010110110",
  37330=>"101101111",
  37331=>"010000001",
  37332=>"100000101",
  37333=>"110011001",
  37334=>"111110101",
  37335=>"111111111",
  37336=>"101011100",
  37337=>"100111000",
  37338=>"001110110",
  37339=>"001010000",
  37340=>"110001000",
  37341=>"001001001",
  37342=>"101110111",
  37343=>"100001100",
  37344=>"010111001",
  37345=>"110000001",
  37346=>"011001010",
  37347=>"101010100",
  37348=>"101010001",
  37349=>"001000101",
  37350=>"100101110",
  37351=>"000010110",
  37352=>"000111111",
  37353=>"101110001",
  37354=>"100110110",
  37355=>"100100001",
  37356=>"110011000",
  37357=>"101011010",
  37358=>"111100111",
  37359=>"011110011",
  37360=>"100110010",
  37361=>"011101001",
  37362=>"111000110",
  37363=>"011110100",
  37364=>"010011000",
  37365=>"010100110",
  37366=>"000000001",
  37367=>"000101111",
  37368=>"111111010",
  37369=>"001001110",
  37370=>"110010001",
  37371=>"000110111",
  37372=>"010001110",
  37373=>"100110001",
  37374=>"100010000",
  37375=>"010000100",
  37376=>"100100110",
  37377=>"001000011",
  37378=>"110100100",
  37379=>"111010000",
  37380=>"010000111",
  37381=>"100110110",
  37382=>"111001110",
  37383=>"101011110",
  37384=>"110100000",
  37385=>"000110101",
  37386=>"001100011",
  37387=>"101110011",
  37388=>"000110010",
  37389=>"110010001",
  37390=>"011000000",
  37391=>"101010100",
  37392=>"100111000",
  37393=>"111010110",
  37394=>"011100111",
  37395=>"110100110",
  37396=>"010100011",
  37397=>"101010001",
  37398=>"000000010",
  37399=>"010000111",
  37400=>"110001010",
  37401=>"011111100",
  37402=>"101110100",
  37403=>"111001000",
  37404=>"110111101",
  37405=>"111010001",
  37406=>"001101010",
  37407=>"010001001",
  37408=>"001011011",
  37409=>"000110100",
  37410=>"110111100",
  37411=>"111001011",
  37412=>"011110011",
  37413=>"010101111",
  37414=>"111101110",
  37415=>"101000100",
  37416=>"100111101",
  37417=>"101000111",
  37418=>"111101101",
  37419=>"000010010",
  37420=>"101111111",
  37421=>"111111011",
  37422=>"101101101",
  37423=>"110111111",
  37424=>"000011010",
  37425=>"111001100",
  37426=>"111000010",
  37427=>"101000001",
  37428=>"100001100",
  37429=>"100100111",
  37430=>"110011001",
  37431=>"000001100",
  37432=>"111101011",
  37433=>"000100000",
  37434=>"100100001",
  37435=>"100111001",
  37436=>"010011011",
  37437=>"001000001",
  37438=>"000110011",
  37439=>"101111111",
  37440=>"111000001",
  37441=>"100000100",
  37442=>"100100011",
  37443=>"000001111",
  37444=>"000010111",
  37445=>"001000110",
  37446=>"110001100",
  37447=>"001001011",
  37448=>"000001101",
  37449=>"110010001",
  37450=>"001011011",
  37451=>"000111000",
  37452=>"111011110",
  37453=>"101000011",
  37454=>"100101001",
  37455=>"001111101",
  37456=>"011111110",
  37457=>"101001110",
  37458=>"110111000",
  37459=>"001000111",
  37460=>"001101110",
  37461=>"001000110",
  37462=>"000100010",
  37463=>"000010011",
  37464=>"000111001",
  37465=>"111100011",
  37466=>"001011011",
  37467=>"110100111",
  37468=>"001001111",
  37469=>"101010000",
  37470=>"001001110",
  37471=>"001110100",
  37472=>"000011110",
  37473=>"010001110",
  37474=>"111111100",
  37475=>"101001011",
  37476=>"100011010",
  37477=>"010001010",
  37478=>"101001101",
  37479=>"000001000",
  37480=>"011100001",
  37481=>"111010110",
  37482=>"000010000",
  37483=>"111011100",
  37484=>"010011110",
  37485=>"001011110",
  37486=>"110001001",
  37487=>"000001110",
  37488=>"000001010",
  37489=>"110011101",
  37490=>"001000011",
  37491=>"000111101",
  37492=>"001100111",
  37493=>"001000010",
  37494=>"100001011",
  37495=>"100011100",
  37496=>"011100001",
  37497=>"100000101",
  37498=>"100011000",
  37499=>"101101100",
  37500=>"011100010",
  37501=>"110001010",
  37502=>"101101001",
  37503=>"111110111",
  37504=>"111000110",
  37505=>"001111100",
  37506=>"000011111",
  37507=>"001101110",
  37508=>"011010111",
  37509=>"111111110",
  37510=>"111111100",
  37511=>"011100000",
  37512=>"011010011",
  37513=>"111111101",
  37514=>"110110100",
  37515=>"100010110",
  37516=>"111100001",
  37517=>"111111100",
  37518=>"001100101",
  37519=>"011010001",
  37520=>"000011111",
  37521=>"001101001",
  37522=>"001000100",
  37523=>"100110110",
  37524=>"001000101",
  37525=>"001110101",
  37526=>"001000001",
  37527=>"101111101",
  37528=>"111100100",
  37529=>"110101001",
  37530=>"110010000",
  37531=>"000010000",
  37532=>"101010101",
  37533=>"010001000",
  37534=>"111111001",
  37535=>"100110010",
  37536=>"111000000",
  37537=>"101000111",
  37538=>"000000000",
  37539=>"100111111",
  37540=>"111010111",
  37541=>"110101000",
  37542=>"100111101",
  37543=>"000000001",
  37544=>"101100011",
  37545=>"101010000",
  37546=>"011101001",
  37547=>"011010110",
  37548=>"000010010",
  37549=>"101000100",
  37550=>"001100100",
  37551=>"101001011",
  37552=>"101111011",
  37553=>"001111000",
  37554=>"100110011",
  37555=>"001111000",
  37556=>"000111010",
  37557=>"100111000",
  37558=>"000110001",
  37559=>"110110100",
  37560=>"101101000",
  37561=>"111010101",
  37562=>"000011011",
  37563=>"101100000",
  37564=>"000101010",
  37565=>"001000000",
  37566=>"011100011",
  37567=>"001011100",
  37568=>"111010011",
  37569=>"000101011",
  37570=>"000100010",
  37571=>"011001010",
  37572=>"001110001",
  37573=>"000000111",
  37574=>"011100011",
  37575=>"100101001",
  37576=>"110000101",
  37577=>"000000111",
  37578=>"000110011",
  37579=>"000001001",
  37580=>"000000010",
  37581=>"010000100",
  37582=>"100110110",
  37583=>"011011000",
  37584=>"000011111",
  37585=>"000100111",
  37586=>"111011100",
  37587=>"101001011",
  37588=>"011011011",
  37589=>"001000010",
  37590=>"110011111",
  37591=>"111000101",
  37592=>"100001000",
  37593=>"111010011",
  37594=>"101101111",
  37595=>"101100111",
  37596=>"000111011",
  37597=>"100101111",
  37598=>"001110100",
  37599=>"010100110",
  37600=>"100001101",
  37601=>"011110111",
  37602=>"100010000",
  37603=>"100001000",
  37604=>"100100010",
  37605=>"001000111",
  37606=>"101010110",
  37607=>"001111111",
  37608=>"011100001",
  37609=>"111111111",
  37610=>"100111101",
  37611=>"000011001",
  37612=>"111101011",
  37613=>"100001100",
  37614=>"010110101",
  37615=>"101101111",
  37616=>"101110001",
  37617=>"110100011",
  37618=>"101111111",
  37619=>"111100010",
  37620=>"101010111",
  37621=>"110001011",
  37622=>"001100110",
  37623=>"010000001",
  37624=>"100010100",
  37625=>"010000101",
  37626=>"011010100",
  37627=>"101110101",
  37628=>"110001110",
  37629=>"100001110",
  37630=>"111001011",
  37631=>"010111000",
  37632=>"111100011",
  37633=>"110110010",
  37634=>"010100100",
  37635=>"100101100",
  37636=>"100001010",
  37637=>"010111110",
  37638=>"000000101",
  37639=>"101111100",
  37640=>"101101100",
  37641=>"100101110",
  37642=>"001111010",
  37643=>"111101010",
  37644=>"111001001",
  37645=>"100101000",
  37646=>"010011001",
  37647=>"111011011",
  37648=>"010110010",
  37649=>"000101011",
  37650=>"010010111",
  37651=>"001001001",
  37652=>"110111011",
  37653=>"010010011",
  37654=>"111101110",
  37655=>"000101000",
  37656=>"111011011",
  37657=>"000010100",
  37658=>"010000111",
  37659=>"100111111",
  37660=>"000110110",
  37661=>"011111101",
  37662=>"111001010",
  37663=>"001110101",
  37664=>"001100111",
  37665=>"001011001",
  37666=>"111110001",
  37667=>"100110001",
  37668=>"010100100",
  37669=>"101000000",
  37670=>"000001000",
  37671=>"011110110",
  37672=>"011010001",
  37673=>"101110111",
  37674=>"101101101",
  37675=>"100000011",
  37676=>"010001100",
  37677=>"010000001",
  37678=>"111011100",
  37679=>"101111110",
  37680=>"010110101",
  37681=>"001101011",
  37682=>"111111000",
  37683=>"011101010",
  37684=>"111010001",
  37685=>"010111100",
  37686=>"010010011",
  37687=>"111001100",
  37688=>"111010100",
  37689=>"001000001",
  37690=>"110111111",
  37691=>"111111100",
  37692=>"110000111",
  37693=>"100101110",
  37694=>"010000000",
  37695=>"000100011",
  37696=>"110001001",
  37697=>"101010010",
  37698=>"110101010",
  37699=>"101010111",
  37700=>"110110110",
  37701=>"101011010",
  37702=>"110000001",
  37703=>"111000101",
  37704=>"001010001",
  37705=>"010000000",
  37706=>"000001111",
  37707=>"110110100",
  37708=>"110101101",
  37709=>"011010000",
  37710=>"110001000",
  37711=>"001011111",
  37712=>"001100010",
  37713=>"100100010",
  37714=>"111111101",
  37715=>"110100101",
  37716=>"011001100",
  37717=>"101011010",
  37718=>"000011010",
  37719=>"100111101",
  37720=>"111011101",
  37721=>"000111010",
  37722=>"010011110",
  37723=>"110010010",
  37724=>"010101110",
  37725=>"101001001",
  37726=>"110000100",
  37727=>"010011000",
  37728=>"100010110",
  37729=>"101001000",
  37730=>"000101101",
  37731=>"111011011",
  37732=>"001101101",
  37733=>"110111001",
  37734=>"011101000",
  37735=>"001110110",
  37736=>"111011110",
  37737=>"101110101",
  37738=>"010011110",
  37739=>"011111010",
  37740=>"101000111",
  37741=>"000111111",
  37742=>"000111110",
  37743=>"010010011",
  37744=>"011001101",
  37745=>"100011111",
  37746=>"101001010",
  37747=>"100111001",
  37748=>"010110101",
  37749=>"101000111",
  37750=>"101110100",
  37751=>"110111101",
  37752=>"101011001",
  37753=>"000101001",
  37754=>"100111000",
  37755=>"110111110",
  37756=>"101011100",
  37757=>"111001000",
  37758=>"010011100",
  37759=>"111110111",
  37760=>"010101111",
  37761=>"010101000",
  37762=>"100110111",
  37763=>"011011011",
  37764=>"010110101",
  37765=>"011000111",
  37766=>"011110011",
  37767=>"011010110",
  37768=>"011111100",
  37769=>"001000101",
  37770=>"111110010",
  37771=>"001110000",
  37772=>"111111010",
  37773=>"000101000",
  37774=>"000111010",
  37775=>"101110001",
  37776=>"000011001",
  37777=>"110110101",
  37778=>"001011100",
  37779=>"011110011",
  37780=>"101100101",
  37781=>"100100001",
  37782=>"100001101",
  37783=>"100010010",
  37784=>"101101110",
  37785=>"110111000",
  37786=>"000111000",
  37787=>"010111101",
  37788=>"010111010",
  37789=>"111111000",
  37790=>"111001010",
  37791=>"111101011",
  37792=>"111110010",
  37793=>"111010011",
  37794=>"100011110",
  37795=>"010100001",
  37796=>"010000111",
  37797=>"110011111",
  37798=>"010001111",
  37799=>"110001101",
  37800=>"111111000",
  37801=>"000111000",
  37802=>"111111111",
  37803=>"010001001",
  37804=>"101100000",
  37805=>"001001010",
  37806=>"110101101",
  37807=>"100110111",
  37808=>"110000101",
  37809=>"001101001",
  37810=>"001010010",
  37811=>"000001001",
  37812=>"110001011",
  37813=>"101001001",
  37814=>"000111111",
  37815=>"101111100",
  37816=>"011011110",
  37817=>"110000101",
  37818=>"011101100",
  37819=>"101100111",
  37820=>"010100111",
  37821=>"001011110",
  37822=>"001101000",
  37823=>"110001111",
  37824=>"010111110",
  37825=>"110011001",
  37826=>"010101110",
  37827=>"010111001",
  37828=>"100000001",
  37829=>"110100100",
  37830=>"100101100",
  37831=>"100001010",
  37832=>"100110110",
  37833=>"111000011",
  37834=>"111000111",
  37835=>"000010100",
  37836=>"010011010",
  37837=>"000101100",
  37838=>"010101111",
  37839=>"100011111",
  37840=>"100110110",
  37841=>"001110110",
  37842=>"011011000",
  37843=>"110000111",
  37844=>"100010101",
  37845=>"010010101",
  37846=>"101001011",
  37847=>"101001000",
  37848=>"100100010",
  37849=>"000000011",
  37850=>"110101011",
  37851=>"011111001",
  37852=>"100101010",
  37853=>"110011100",
  37854=>"010111001",
  37855=>"100110010",
  37856=>"011100110",
  37857=>"100101101",
  37858=>"101100110",
  37859=>"001001011",
  37860=>"101110011",
  37861=>"101000000",
  37862=>"110010000",
  37863=>"100101010",
  37864=>"010011100",
  37865=>"110001001",
  37866=>"100011111",
  37867=>"001111110",
  37868=>"010111111",
  37869=>"100100101",
  37870=>"000001011",
  37871=>"110000111",
  37872=>"101101110",
  37873=>"111100011",
  37874=>"111011111",
  37875=>"010111100",
  37876=>"100101000",
  37877=>"101001000",
  37878=>"100001101",
  37879=>"011000010",
  37880=>"010000110",
  37881=>"001100101",
  37882=>"100001010",
  37883=>"000110101",
  37884=>"111010000",
  37885=>"110000111",
  37886=>"001100011",
  37887=>"001001110",
  37888=>"000011100",
  37889=>"011010111",
  37890=>"110101000",
  37891=>"101001010",
  37892=>"000000000",
  37893=>"001101011",
  37894=>"001000100",
  37895=>"111001101",
  37896=>"110110111",
  37897=>"100000001",
  37898=>"000110010",
  37899=>"001100010",
  37900=>"000010011",
  37901=>"110000010",
  37902=>"000001001",
  37903=>"001111111",
  37904=>"101011101",
  37905=>"111001010",
  37906=>"000100010",
  37907=>"110000011",
  37908=>"100101011",
  37909=>"011001100",
  37910=>"010001011",
  37911=>"011000010",
  37912=>"001100101",
  37913=>"010011100",
  37914=>"011001100",
  37915=>"011010010",
  37916=>"011110000",
  37917=>"100000000",
  37918=>"100100111",
  37919=>"110001111",
  37920=>"110010111",
  37921=>"101010111",
  37922=>"110010100",
  37923=>"010011010",
  37924=>"000100000",
  37925=>"100110100",
  37926=>"010101100",
  37927=>"001010000",
  37928=>"111111101",
  37929=>"001001010",
  37930=>"101101101",
  37931=>"110100011",
  37932=>"111111110",
  37933=>"001011110",
  37934=>"101010111",
  37935=>"011000000",
  37936=>"000010100",
  37937=>"111000110",
  37938=>"001000000",
  37939=>"001010110",
  37940=>"110111110",
  37941=>"111011110",
  37942=>"111111000",
  37943=>"100101100",
  37944=>"111000110",
  37945=>"101000011",
  37946=>"100000011",
  37947=>"111000001",
  37948=>"010010001",
  37949=>"101100100",
  37950=>"011111110",
  37951=>"111101110",
  37952=>"000000011",
  37953=>"010010001",
  37954=>"100000010",
  37955=>"010100000",
  37956=>"100000011",
  37957=>"111100011",
  37958=>"100001010",
  37959=>"000111000",
  37960=>"001000001",
  37961=>"110011111",
  37962=>"111101000",
  37963=>"111010011",
  37964=>"100001100",
  37965=>"110110001",
  37966=>"000101011",
  37967=>"011110111",
  37968=>"111010001",
  37969=>"000001101",
  37970=>"000110101",
  37971=>"100000101",
  37972=>"110111111",
  37973=>"000110010",
  37974=>"010111011",
  37975=>"110001010",
  37976=>"101110111",
  37977=>"110000111",
  37978=>"101011000",
  37979=>"010001000",
  37980=>"001001111",
  37981=>"011001111",
  37982=>"101111011",
  37983=>"001010001",
  37984=>"110010011",
  37985=>"011011100",
  37986=>"000100110",
  37987=>"001011111",
  37988=>"000010010",
  37989=>"110101010",
  37990=>"011111111",
  37991=>"010111010",
  37992=>"010001100",
  37993=>"000001000",
  37994=>"010110000",
  37995=>"100111000",
  37996=>"011011000",
  37997=>"100001111",
  37998=>"101110011",
  37999=>"110001001",
  38000=>"001000110",
  38001=>"000010010",
  38002=>"010010010",
  38003=>"000000111",
  38004=>"100010010",
  38005=>"110100111",
  38006=>"001001000",
  38007=>"000101100",
  38008=>"100000010",
  38009=>"110100000",
  38010=>"011111111",
  38011=>"011010010",
  38012=>"100010000",
  38013=>"011100010",
  38014=>"011011101",
  38015=>"010101011",
  38016=>"111001110",
  38017=>"000001011",
  38018=>"111010011",
  38019=>"111010010",
  38020=>"000000010",
  38021=>"001010100",
  38022=>"010110101",
  38023=>"100011000",
  38024=>"010000000",
  38025=>"010101111",
  38026=>"101000011",
  38027=>"001110110",
  38028=>"111101010",
  38029=>"011100111",
  38030=>"000001110",
  38031=>"110010100",
  38032=>"010011010",
  38033=>"001111010",
  38034=>"110001000",
  38035=>"111100010",
  38036=>"001111101",
  38037=>"010100110",
  38038=>"111001101",
  38039=>"001100001",
  38040=>"010101110",
  38041=>"011000001",
  38042=>"101100110",
  38043=>"110101011",
  38044=>"111010000",
  38045=>"000111100",
  38046=>"001001010",
  38047=>"101110010",
  38048=>"000100000",
  38049=>"101101001",
  38050=>"001111001",
  38051=>"111010111",
  38052=>"110011111",
  38053=>"010000100",
  38054=>"100101001",
  38055=>"111111111",
  38056=>"110011010",
  38057=>"110101110",
  38058=>"001011111",
  38059=>"110011000",
  38060=>"000101000",
  38061=>"001010000",
  38062=>"101000110",
  38063=>"100011010",
  38064=>"000001001",
  38065=>"000000111",
  38066=>"110011011",
  38067=>"100010001",
  38068=>"000101010",
  38069=>"011110011",
  38070=>"011110010",
  38071=>"110101001",
  38072=>"101010111",
  38073=>"110001010",
  38074=>"100100110",
  38075=>"010011110",
  38076=>"011101101",
  38077=>"101001001",
  38078=>"101001010",
  38079=>"000011001",
  38080=>"000101111",
  38081=>"000010011",
  38082=>"000010011",
  38083=>"100101101",
  38084=>"010001010",
  38085=>"110101000",
  38086=>"010000101",
  38087=>"011101010",
  38088=>"010100100",
  38089=>"111110111",
  38090=>"001101101",
  38091=>"100111010",
  38092=>"000111000",
  38093=>"001101100",
  38094=>"010101000",
  38095=>"001010010",
  38096=>"001101001",
  38097=>"001001100",
  38098=>"010001111",
  38099=>"100110011",
  38100=>"010110110",
  38101=>"001000011",
  38102=>"000001101",
  38103=>"110011001",
  38104=>"001100011",
  38105=>"101000000",
  38106=>"000111100",
  38107=>"100111110",
  38108=>"101011011",
  38109=>"010010110",
  38110=>"110111101",
  38111=>"111011001",
  38112=>"100010110",
  38113=>"011110111",
  38114=>"110111001",
  38115=>"000101111",
  38116=>"101100110",
  38117=>"111110100",
  38118=>"000001001",
  38119=>"110010010",
  38120=>"100001010",
  38121=>"100110111",
  38122=>"101011000",
  38123=>"101100100",
  38124=>"101111011",
  38125=>"110110100",
  38126=>"010101010",
  38127=>"010101001",
  38128=>"010111001",
  38129=>"101110111",
  38130=>"011100000",
  38131=>"111001100",
  38132=>"101011000",
  38133=>"000111001",
  38134=>"000101110",
  38135=>"010101101",
  38136=>"010101110",
  38137=>"010001000",
  38138=>"011001101",
  38139=>"010001110",
  38140=>"001001000",
  38141=>"010001111",
  38142=>"000100000",
  38143=>"101011100",
  38144=>"101100101",
  38145=>"100001101",
  38146=>"000100001",
  38147=>"001110010",
  38148=>"111101110",
  38149=>"000111111",
  38150=>"101110001",
  38151=>"011100001",
  38152=>"010010000",
  38153=>"011111100",
  38154=>"010110101",
  38155=>"110110101",
  38156=>"010011011",
  38157=>"110110011",
  38158=>"001000110",
  38159=>"111110100",
  38160=>"100100100",
  38161=>"001110010",
  38162=>"010111011",
  38163=>"000110100",
  38164=>"101101111",
  38165=>"011110011",
  38166=>"111011001",
  38167=>"000110110",
  38168=>"100001101",
  38169=>"001101110",
  38170=>"111111111",
  38171=>"110101110",
  38172=>"000100111",
  38173=>"001110101",
  38174=>"011001101",
  38175=>"000011010",
  38176=>"011110011",
  38177=>"100011101",
  38178=>"000110010",
  38179=>"001000000",
  38180=>"010000010",
  38181=>"101111011",
  38182=>"010011000",
  38183=>"011101101",
  38184=>"010111001",
  38185=>"000110000",
  38186=>"000100000",
  38187=>"011000111",
  38188=>"010110010",
  38189=>"010010110",
  38190=>"100000101",
  38191=>"110100110",
  38192=>"001000010",
  38193=>"110010111",
  38194=>"111100010",
  38195=>"000000010",
  38196=>"000011101",
  38197=>"000111110",
  38198=>"011100001",
  38199=>"110111011",
  38200=>"000000101",
  38201=>"110000001",
  38202=>"100011011",
  38203=>"011101100",
  38204=>"001110011",
  38205=>"110111100",
  38206=>"001000100",
  38207=>"110101110",
  38208=>"101111110",
  38209=>"100111110",
  38210=>"010000100",
  38211=>"010010100",
  38212=>"010101000",
  38213=>"110001001",
  38214=>"111101000",
  38215=>"000011011",
  38216=>"111111111",
  38217=>"110100100",
  38218=>"000001011",
  38219=>"010011101",
  38220=>"110100101",
  38221=>"111100001",
  38222=>"000101100",
  38223=>"000010100",
  38224=>"010110100",
  38225=>"010000100",
  38226=>"110011111",
  38227=>"111101010",
  38228=>"000001111",
  38229=>"100110000",
  38230=>"110000100",
  38231=>"100111101",
  38232=>"010011011",
  38233=>"001100001",
  38234=>"001111110",
  38235=>"000000110",
  38236=>"101001111",
  38237=>"100011111",
  38238=>"101100001",
  38239=>"011001011",
  38240=>"001101011",
  38241=>"110101110",
  38242=>"100110001",
  38243=>"010101101",
  38244=>"110011111",
  38245=>"001001100",
  38246=>"111010011",
  38247=>"100000100",
  38248=>"100100111",
  38249=>"111001000",
  38250=>"101000010",
  38251=>"010100111",
  38252=>"011100100",
  38253=>"011111111",
  38254=>"111010100",
  38255=>"010011110",
  38256=>"100010011",
  38257=>"111110001",
  38258=>"011101100",
  38259=>"101100001",
  38260=>"010001011",
  38261=>"000010110",
  38262=>"001011010",
  38263=>"000100100",
  38264=>"100100100",
  38265=>"100011111",
  38266=>"100100110",
  38267=>"110111110",
  38268=>"101100001",
  38269=>"011111011",
  38270=>"001011100",
  38271=>"011000000",
  38272=>"000010101",
  38273=>"010000001",
  38274=>"101010001",
  38275=>"010111111",
  38276=>"110101111",
  38277=>"100100000",
  38278=>"100101010",
  38279=>"000101011",
  38280=>"100101001",
  38281=>"110111000",
  38282=>"111011011",
  38283=>"111110011",
  38284=>"011010111",
  38285=>"000010011",
  38286=>"001100010",
  38287=>"111111101",
  38288=>"100110000",
  38289=>"010010000",
  38290=>"000010000",
  38291=>"101001111",
  38292=>"001001100",
  38293=>"101001000",
  38294=>"100100010",
  38295=>"010100011",
  38296=>"000001011",
  38297=>"000101100",
  38298=>"001011001",
  38299=>"111011100",
  38300=>"111101110",
  38301=>"010111101",
  38302=>"101110100",
  38303=>"101110000",
  38304=>"000010100",
  38305=>"010001001",
  38306=>"100011011",
  38307=>"111001100",
  38308=>"001111000",
  38309=>"011010000",
  38310=>"001101110",
  38311=>"101010001",
  38312=>"000110011",
  38313=>"100101101",
  38314=>"010100010",
  38315=>"010011000",
  38316=>"110100100",
  38317=>"010000010",
  38318=>"001011111",
  38319=>"001111111",
  38320=>"110001010",
  38321=>"001101000",
  38322=>"010100110",
  38323=>"111111111",
  38324=>"110000001",
  38325=>"111011000",
  38326=>"100111100",
  38327=>"011010001",
  38328=>"101001010",
  38329=>"100010001",
  38330=>"000011111",
  38331=>"001011000",
  38332=>"101101000",
  38333=>"110111110",
  38334=>"010100100",
  38335=>"001001001",
  38336=>"110100111",
  38337=>"001110011",
  38338=>"101001111",
  38339=>"011010100",
  38340=>"100111000",
  38341=>"111101000",
  38342=>"111101110",
  38343=>"000000001",
  38344=>"100001110",
  38345=>"000000010",
  38346=>"110111001",
  38347=>"111011111",
  38348=>"100111011",
  38349=>"010010110",
  38350=>"000000011",
  38351=>"101000110",
  38352=>"111001100",
  38353=>"011000000",
  38354=>"001011110",
  38355=>"110101111",
  38356=>"000000111",
  38357=>"110101001",
  38358=>"101110111",
  38359=>"100101011",
  38360=>"100000100",
  38361=>"111101001",
  38362=>"110111000",
  38363=>"111101001",
  38364=>"000101010",
  38365=>"100010111",
  38366=>"110101001",
  38367=>"101100110",
  38368=>"000100010",
  38369=>"001000011",
  38370=>"011000000",
  38371=>"001001001",
  38372=>"111111010",
  38373=>"011111110",
  38374=>"011100011",
  38375=>"101100010",
  38376=>"011011000",
  38377=>"100110100",
  38378=>"111000010",
  38379=>"100101100",
  38380=>"010101110",
  38381=>"100001001",
  38382=>"011101010",
  38383=>"001100100",
  38384=>"010011011",
  38385=>"110101110",
  38386=>"101101110",
  38387=>"110010011",
  38388=>"110110110",
  38389=>"111101000",
  38390=>"001000100",
  38391=>"110101111",
  38392=>"111101100",
  38393=>"111111110",
  38394=>"100010001",
  38395=>"010101100",
  38396=>"100011111",
  38397=>"000000110",
  38398=>"000101000",
  38399=>"011011011",
  38400=>"010001111",
  38401=>"011011100",
  38402=>"010111000",
  38403=>"011111100",
  38404=>"100001000",
  38405=>"111001000",
  38406=>"011010000",
  38407=>"000110101",
  38408=>"100000100",
  38409=>"111011000",
  38410=>"100100000",
  38411=>"111000000",
  38412=>"111001101",
  38413=>"010100001",
  38414=>"001101010",
  38415=>"001110110",
  38416=>"000100001",
  38417=>"001110101",
  38418=>"010100001",
  38419=>"011100100",
  38420=>"100100000",
  38421=>"101010100",
  38422=>"000010101",
  38423=>"101001110",
  38424=>"001011001",
  38425=>"010011011",
  38426=>"111010110",
  38427=>"101101100",
  38428=>"001111011",
  38429=>"001100111",
  38430=>"101000101",
  38431=>"110000101",
  38432=>"101011011",
  38433=>"110011011",
  38434=>"001001001",
  38435=>"100101011",
  38436=>"100111100",
  38437=>"011010001",
  38438=>"101110100",
  38439=>"001100110",
  38440=>"001110110",
  38441=>"010111111",
  38442=>"011010010",
  38443=>"110000110",
  38444=>"010010111",
  38445=>"000100110",
  38446=>"001110111",
  38447=>"000010100",
  38448=>"111110011",
  38449=>"001111001",
  38450=>"111010101",
  38451=>"110111101",
  38452=>"011111000",
  38453=>"001100000",
  38454=>"111101100",
  38455=>"001101110",
  38456=>"000111011",
  38457=>"111111000",
  38458=>"110010111",
  38459=>"100111010",
  38460=>"100110011",
  38461=>"101110000",
  38462=>"111000101",
  38463=>"010101011",
  38464=>"000100000",
  38465=>"110100001",
  38466=>"000010111",
  38467=>"010111001",
  38468=>"000010101",
  38469=>"010000011",
  38470=>"111110011",
  38471=>"010001011",
  38472=>"110111110",
  38473=>"101110010",
  38474=>"000000000",
  38475=>"111110110",
  38476=>"000100000",
  38477=>"100000001",
  38478=>"111100011",
  38479=>"001100001",
  38480=>"100000001",
  38481=>"100011110",
  38482=>"000000101",
  38483=>"101100100",
  38484=>"011101001",
  38485=>"000111101",
  38486=>"001100100",
  38487=>"010000000",
  38488=>"001111101",
  38489=>"010010010",
  38490=>"111110010",
  38491=>"010111010",
  38492=>"110010100",
  38493=>"101000010",
  38494=>"101001110",
  38495=>"110011111",
  38496=>"110001101",
  38497=>"001111000",
  38498=>"000111111",
  38499=>"100000101",
  38500=>"000010111",
  38501=>"101001010",
  38502=>"110000111",
  38503=>"100011011",
  38504=>"111010111",
  38505=>"010111110",
  38506=>"010011000",
  38507=>"111001010",
  38508=>"111011010",
  38509=>"000111010",
  38510=>"110110101",
  38511=>"110111111",
  38512=>"000011011",
  38513=>"010111010",
  38514=>"011101000",
  38515=>"000101011",
  38516=>"001001010",
  38517=>"100011101",
  38518=>"110010011",
  38519=>"000110111",
  38520=>"000111100",
  38521=>"001010010",
  38522=>"001101100",
  38523=>"010100010",
  38524=>"100100000",
  38525=>"100010000",
  38526=>"001101111",
  38527=>"010010111",
  38528=>"011111100",
  38529=>"110001011",
  38530=>"011011000",
  38531=>"100001011",
  38532=>"011110100",
  38533=>"100111111",
  38534=>"000110110",
  38535=>"110000111",
  38536=>"011001111",
  38537=>"001011000",
  38538=>"101001101",
  38539=>"001100111",
  38540=>"101010001",
  38541=>"110110010",
  38542=>"011011011",
  38543=>"011001011",
  38544=>"011010000",
  38545=>"110001111",
  38546=>"000000100",
  38547=>"011101001",
  38548=>"100101101",
  38549=>"100010110",
  38550=>"111000011",
  38551=>"101110110",
  38552=>"000000101",
  38553=>"111001101",
  38554=>"001101001",
  38555=>"111110110",
  38556=>"011011011",
  38557=>"001010001",
  38558=>"111101011",
  38559=>"101000010",
  38560=>"011100010",
  38561=>"011110011",
  38562=>"100111111",
  38563=>"011000001",
  38564=>"010110010",
  38565=>"001101111",
  38566=>"010000100",
  38567=>"000111011",
  38568=>"100101001",
  38569=>"010100010",
  38570=>"011011111",
  38571=>"101110011",
  38572=>"110010111",
  38573=>"011100100",
  38574=>"000110100",
  38575=>"111110110",
  38576=>"011101111",
  38577=>"111011111",
  38578=>"101101000",
  38579=>"001101001",
  38580=>"111010010",
  38581=>"101010000",
  38582=>"111100110",
  38583=>"101001010",
  38584=>"010011010",
  38585=>"011110100",
  38586=>"101011100",
  38587=>"000010111",
  38588=>"110000011",
  38589=>"100011101",
  38590=>"101111010",
  38591=>"000101111",
  38592=>"111001011",
  38593=>"001001111",
  38594=>"101001011",
  38595=>"000001110",
  38596=>"101010010",
  38597=>"010110111",
  38598=>"001000011",
  38599=>"001000011",
  38600=>"011101110",
  38601=>"000011011",
  38602=>"101010010",
  38603=>"001000100",
  38604=>"100001011",
  38605=>"110110011",
  38606=>"011101000",
  38607=>"100010011",
  38608=>"010100001",
  38609=>"100010001",
  38610=>"110100100",
  38611=>"110001101",
  38612=>"000010100",
  38613=>"001100100",
  38614=>"000000011",
  38615=>"101001111",
  38616=>"000110001",
  38617=>"101100111",
  38618=>"001000011",
  38619=>"010111100",
  38620=>"111100101",
  38621=>"100001001",
  38622=>"000001111",
  38623=>"010001000",
  38624=>"010000101",
  38625=>"000011111",
  38626=>"001001001",
  38627=>"010001101",
  38628=>"001010111",
  38629=>"001011000",
  38630=>"101110110",
  38631=>"111001010",
  38632=>"001011010",
  38633=>"010001000",
  38634=>"100111111",
  38635=>"011001010",
  38636=>"101101010",
  38637=>"101111011",
  38638=>"100111010",
  38639=>"110110111",
  38640=>"010100000",
  38641=>"001101111",
  38642=>"100000000",
  38643=>"111000001",
  38644=>"100100101",
  38645=>"111011111",
  38646=>"000011100",
  38647=>"011111110",
  38648=>"100010101",
  38649=>"111101100",
  38650=>"100100001",
  38651=>"001001111",
  38652=>"011001101",
  38653=>"110110111",
  38654=>"011101011",
  38655=>"010111110",
  38656=>"110100101",
  38657=>"000101100",
  38658=>"101010011",
  38659=>"011000111",
  38660=>"111101010",
  38661=>"100001100",
  38662=>"101100011",
  38663=>"111101101",
  38664=>"101000100",
  38665=>"010001001",
  38666=>"111011111",
  38667=>"000110100",
  38668=>"110110011",
  38669=>"101100101",
  38670=>"001111111",
  38671=>"101110010",
  38672=>"010000010",
  38673=>"010010010",
  38674=>"101000000",
  38675=>"001000111",
  38676=>"110001011",
  38677=>"110110100",
  38678=>"000001110",
  38679=>"011100101",
  38680=>"101101010",
  38681=>"100100011",
  38682=>"111101000",
  38683=>"100101010",
  38684=>"101111000",
  38685=>"001101010",
  38686=>"000011101",
  38687=>"111101001",
  38688=>"000000100",
  38689=>"100011101",
  38690=>"010011111",
  38691=>"010010001",
  38692=>"011111110",
  38693=>"000110001",
  38694=>"111101101",
  38695=>"000111000",
  38696=>"110110010",
  38697=>"010110110",
  38698=>"000100111",
  38699=>"011000000",
  38700=>"101001111",
  38701=>"001000011",
  38702=>"000001011",
  38703=>"101100100",
  38704=>"110100110",
  38705=>"101001110",
  38706=>"011001001",
  38707=>"010101111",
  38708=>"111011101",
  38709=>"110100010",
  38710=>"011000010",
  38711=>"000001100",
  38712=>"101110111",
  38713=>"110000100",
  38714=>"010010010",
  38715=>"011111001",
  38716=>"111010101",
  38717=>"100000111",
  38718=>"010010011",
  38719=>"001111000",
  38720=>"010010101",
  38721=>"000100100",
  38722=>"111001000",
  38723=>"111011100",
  38724=>"001000010",
  38725=>"011111001",
  38726=>"011000000",
  38727=>"101011100",
  38728=>"011101010",
  38729=>"100000010",
  38730=>"011111111",
  38731=>"011001011",
  38732=>"100010001",
  38733=>"100110101",
  38734=>"111011010",
  38735=>"111011111",
  38736=>"001001100",
  38737=>"110100111",
  38738=>"011011010",
  38739=>"010011111",
  38740=>"101011111",
  38741=>"010100111",
  38742=>"001011010",
  38743=>"011011011",
  38744=>"110110110",
  38745=>"011000101",
  38746=>"011001001",
  38747=>"100100011",
  38748=>"011010011",
  38749=>"011001111",
  38750=>"110011011",
  38751=>"010000001",
  38752=>"111011010",
  38753=>"111111111",
  38754=>"010100010",
  38755=>"001011111",
  38756=>"110110101",
  38757=>"000000010",
  38758=>"110011010",
  38759=>"110010000",
  38760=>"100011011",
  38761=>"001101001",
  38762=>"101011010",
  38763=>"001110011",
  38764=>"110101011",
  38765=>"111010111",
  38766=>"101111111",
  38767=>"110010100",
  38768=>"101001010",
  38769=>"010001011",
  38770=>"010100011",
  38771=>"001000011",
  38772=>"010001111",
  38773=>"101111101",
  38774=>"000010100",
  38775=>"111010001",
  38776=>"011001011",
  38777=>"100111010",
  38778=>"001000110",
  38779=>"001010110",
  38780=>"011011001",
  38781=>"101001111",
  38782=>"010000011",
  38783=>"001111100",
  38784=>"101001100",
  38785=>"000001000",
  38786=>"101110110",
  38787=>"010111000",
  38788=>"001101111",
  38789=>"100011110",
  38790=>"000000110",
  38791=>"000100101",
  38792=>"010011111",
  38793=>"110010101",
  38794=>"000001100",
  38795=>"010100000",
  38796=>"011110110",
  38797=>"010100111",
  38798=>"000010011",
  38799=>"101110000",
  38800=>"001000001",
  38801=>"101000100",
  38802=>"000001000",
  38803=>"001101001",
  38804=>"000100001",
  38805=>"101011110",
  38806=>"000111001",
  38807=>"011111111",
  38808=>"001110001",
  38809=>"101011101",
  38810=>"011110111",
  38811=>"000100100",
  38812=>"000000000",
  38813=>"011110010",
  38814=>"111010111",
  38815=>"001110000",
  38816=>"001001111",
  38817=>"010000111",
  38818=>"011110110",
  38819=>"101000111",
  38820=>"110010010",
  38821=>"110111011",
  38822=>"101001000",
  38823=>"101011010",
  38824=>"100000101",
  38825=>"010011000",
  38826=>"111011111",
  38827=>"110011000",
  38828=>"101010000",
  38829=>"011010110",
  38830=>"010100100",
  38831=>"010001110",
  38832=>"011101000",
  38833=>"000001100",
  38834=>"111000111",
  38835=>"010110010",
  38836=>"001111000",
  38837=>"111011111",
  38838=>"101100111",
  38839=>"001111011",
  38840=>"011010010",
  38841=>"111100011",
  38842=>"011010001",
  38843=>"110011100",
  38844=>"010011001",
  38845=>"011101000",
  38846=>"000000111",
  38847=>"100011011",
  38848=>"000101100",
  38849=>"011001100",
  38850=>"101100110",
  38851=>"100000100",
  38852=>"111100010",
  38853=>"001000001",
  38854=>"110010001",
  38855=>"101010100",
  38856=>"011110111",
  38857=>"100111001",
  38858=>"111000101",
  38859=>"000101110",
  38860=>"100100010",
  38861=>"110001000",
  38862=>"000101010",
  38863=>"100100111",
  38864=>"010010100",
  38865=>"001011110",
  38866=>"111000000",
  38867=>"100000111",
  38868=>"010001011",
  38869=>"100000101",
  38870=>"101001001",
  38871=>"010000110",
  38872=>"011100100",
  38873=>"101000001",
  38874=>"010001010",
  38875=>"111110110",
  38876=>"101001000",
  38877=>"111011110",
  38878=>"000011000",
  38879=>"111110001",
  38880=>"000100001",
  38881=>"011010001",
  38882=>"110010001",
  38883=>"110000110",
  38884=>"001111111",
  38885=>"101011100",
  38886=>"111101111",
  38887=>"001110111",
  38888=>"000110000",
  38889=>"001010111",
  38890=>"110010100",
  38891=>"001001111",
  38892=>"001001111",
  38893=>"011101101",
  38894=>"100100110",
  38895=>"010111101",
  38896=>"101100110",
  38897=>"101101100",
  38898=>"001111100",
  38899=>"001111000",
  38900=>"001100011",
  38901=>"110110101",
  38902=>"001100001",
  38903=>"000010001",
  38904=>"000001101",
  38905=>"101111000",
  38906=>"010010100",
  38907=>"101010101",
  38908=>"011011000",
  38909=>"011011111",
  38910=>"101000111",
  38911=>"000001001",
  38912=>"010000010",
  38913=>"000101010",
  38914=>"101010101",
  38915=>"101000000",
  38916=>"010111011",
  38917=>"001010011",
  38918=>"011100101",
  38919=>"010011011",
  38920=>"110111001",
  38921=>"000000100",
  38922=>"011110100",
  38923=>"001001111",
  38924=>"101110101",
  38925=>"111101001",
  38926=>"111100110",
  38927=>"110000001",
  38928=>"110011000",
  38929=>"010100101",
  38930=>"100000011",
  38931=>"101101101",
  38932=>"110111110",
  38933=>"101100010",
  38934=>"011011101",
  38935=>"110110101",
  38936=>"110011000",
  38937=>"001010110",
  38938=>"110100001",
  38939=>"010010100",
  38940=>"101100010",
  38941=>"001000101",
  38942=>"111001101",
  38943=>"001101100",
  38944=>"101110111",
  38945=>"000000100",
  38946=>"101011110",
  38947=>"100100110",
  38948=>"111111011",
  38949=>"010111011",
  38950=>"100000001",
  38951=>"110100000",
  38952=>"101111100",
  38953=>"001000000",
  38954=>"111000111",
  38955=>"111110101",
  38956=>"001000001",
  38957=>"111001111",
  38958=>"111000000",
  38959=>"111000010",
  38960=>"101010011",
  38961=>"111000110",
  38962=>"001001011",
  38963=>"011111111",
  38964=>"101100011",
  38965=>"000110011",
  38966=>"110100000",
  38967=>"010110001",
  38968=>"111010110",
  38969=>"111110001",
  38970=>"110001011",
  38971=>"101110111",
  38972=>"000000010",
  38973=>"101000000",
  38974=>"000110000",
  38975=>"110111101",
  38976=>"011101011",
  38977=>"001110001",
  38978=>"010101110",
  38979=>"011000111",
  38980=>"110101100",
  38981=>"100010100",
  38982=>"001110010",
  38983=>"110010110",
  38984=>"001101110",
  38985=>"011111010",
  38986=>"101101001",
  38987=>"001000100",
  38988=>"001100001",
  38989=>"100010010",
  38990=>"110011000",
  38991=>"010100010",
  38992=>"001001101",
  38993=>"111110011",
  38994=>"010101111",
  38995=>"001111100",
  38996=>"010000001",
  38997=>"010100110",
  38998=>"111111011",
  38999=>"001011111",
  39000=>"100011101",
  39001=>"010100010",
  39002=>"101100001",
  39003=>"101100100",
  39004=>"110000100",
  39005=>"101110110",
  39006=>"101111111",
  39007=>"100110101",
  39008=>"010100101",
  39009=>"111111000",
  39010=>"010000111",
  39011=>"001000101",
  39012=>"111110011",
  39013=>"100001011",
  39014=>"100010100",
  39015=>"011001100",
  39016=>"001100010",
  39017=>"110110110",
  39018=>"110001001",
  39019=>"101000001",
  39020=>"000100111",
  39021=>"101111000",
  39022=>"000010000",
  39023=>"101001001",
  39024=>"110101110",
  39025=>"010011100",
  39026=>"011001010",
  39027=>"100111111",
  39028=>"000110001",
  39029=>"110011100",
  39030=>"000001001",
  39031=>"010100000",
  39032=>"000100111",
  39033=>"000111000",
  39034=>"010100011",
  39035=>"111100110",
  39036=>"110111101",
  39037=>"011111011",
  39038=>"001001011",
  39039=>"011011000",
  39040=>"001110100",
  39041=>"000011010",
  39042=>"111000000",
  39043=>"000010110",
  39044=>"010001110",
  39045=>"110110111",
  39046=>"010001101",
  39047=>"000000110",
  39048=>"110000001",
  39049=>"110101111",
  39050=>"011100011",
  39051=>"111100101",
  39052=>"010110000",
  39053=>"111011001",
  39054=>"111000101",
  39055=>"100000001",
  39056=>"110101111",
  39057=>"010001110",
  39058=>"000000110",
  39059=>"110101110",
  39060=>"101011010",
  39061=>"011001110",
  39062=>"101101011",
  39063=>"111010111",
  39064=>"101110001",
  39065=>"010011011",
  39066=>"111011010",
  39067=>"010001110",
  39068=>"010000001",
  39069=>"111111010",
  39070=>"100011011",
  39071=>"100110010",
  39072=>"001100111",
  39073=>"001111110",
  39074=>"101010111",
  39075=>"001101000",
  39076=>"011001111",
  39077=>"111111100",
  39078=>"110111111",
  39079=>"011000000",
  39080=>"010101001",
  39081=>"001101010",
  39082=>"101011111",
  39083=>"111101010",
  39084=>"111111001",
  39085=>"101010011",
  39086=>"110000000",
  39087=>"100001110",
  39088=>"110011010",
  39089=>"010110010",
  39090=>"111111010",
  39091=>"111101011",
  39092=>"111111010",
  39093=>"010100001",
  39094=>"000001101",
  39095=>"000010111",
  39096=>"000100010",
  39097=>"001101000",
  39098=>"000001101",
  39099=>"110111001",
  39100=>"001100000",
  39101=>"011001111",
  39102=>"000100011",
  39103=>"001100110",
  39104=>"111001001",
  39105=>"100101000",
  39106=>"111111110",
  39107=>"110000010",
  39108=>"111111101",
  39109=>"100110111",
  39110=>"101100000",
  39111=>"001001110",
  39112=>"011110011",
  39113=>"000011111",
  39114=>"010011001",
  39115=>"111010110",
  39116=>"111111001",
  39117=>"110000000",
  39118=>"011000100",
  39119=>"000101001",
  39120=>"101101011",
  39121=>"100000100",
  39122=>"001010010",
  39123=>"000101101",
  39124=>"110100011",
  39125=>"001100000",
  39126=>"011111011",
  39127=>"010100001",
  39128=>"000011001",
  39129=>"000111011",
  39130=>"101000011",
  39131=>"101010010",
  39132=>"111100110",
  39133=>"101110000",
  39134=>"110100011",
  39135=>"001001111",
  39136=>"111111101",
  39137=>"101011000",
  39138=>"011000010",
  39139=>"101001100",
  39140=>"111111011",
  39141=>"010001010",
  39142=>"011000010",
  39143=>"110010011",
  39144=>"001100011",
  39145=>"001001010",
  39146=>"011011110",
  39147=>"000001100",
  39148=>"001100010",
  39149=>"010000001",
  39150=>"111011010",
  39151=>"011011011",
  39152=>"000110010",
  39153=>"000000100",
  39154=>"111010000",
  39155=>"100111010",
  39156=>"011011111",
  39157=>"011011011",
  39158=>"101010111",
  39159=>"011110000",
  39160=>"110010001",
  39161=>"100010000",
  39162=>"011000110",
  39163=>"001110000",
  39164=>"000111001",
  39165=>"111111100",
  39166=>"000100000",
  39167=>"110110110",
  39168=>"110011001",
  39169=>"001010000",
  39170=>"111110101",
  39171=>"100000100",
  39172=>"101001001",
  39173=>"110100100",
  39174=>"010111010",
  39175=>"111100110",
  39176=>"000010010",
  39177=>"110110001",
  39178=>"011011111",
  39179=>"101110111",
  39180=>"001110011",
  39181=>"011111110",
  39182=>"010100101",
  39183=>"111000000",
  39184=>"001100110",
  39185=>"010011011",
  39186=>"010000000",
  39187=>"101110101",
  39188=>"111101001",
  39189=>"100110101",
  39190=>"101011010",
  39191=>"000010010",
  39192=>"011000001",
  39193=>"001110101",
  39194=>"100111000",
  39195=>"010110101",
  39196=>"111111111",
  39197=>"110100000",
  39198=>"111010011",
  39199=>"010111001",
  39200=>"001100010",
  39201=>"000101001",
  39202=>"011001110",
  39203=>"010011011",
  39204=>"011101001",
  39205=>"100111111",
  39206=>"011000100",
  39207=>"001111101",
  39208=>"001100101",
  39209=>"111110000",
  39210=>"011000001",
  39211=>"111110110",
  39212=>"110100010",
  39213=>"000100111",
  39214=>"101111110",
  39215=>"100000110",
  39216=>"100010000",
  39217=>"101001000",
  39218=>"110000011",
  39219=>"100100000",
  39220=>"111110011",
  39221=>"100010101",
  39222=>"100001111",
  39223=>"000000101",
  39224=>"111101011",
  39225=>"001100010",
  39226=>"100101001",
  39227=>"000001110",
  39228=>"001011110",
  39229=>"011010110",
  39230=>"111001101",
  39231=>"000000100",
  39232=>"101001110",
  39233=>"100000100",
  39234=>"101110011",
  39235=>"010000001",
  39236=>"001100100",
  39237=>"010101101",
  39238=>"000011000",
  39239=>"100110000",
  39240=>"100000101",
  39241=>"110000010",
  39242=>"000111100",
  39243=>"011001010",
  39244=>"000010001",
  39245=>"000100100",
  39246=>"001101110",
  39247=>"010101011",
  39248=>"010111001",
  39249=>"101111110",
  39250=>"101101101",
  39251=>"000110000",
  39252=>"010100000",
  39253=>"011001010",
  39254=>"110101000",
  39255=>"101010001",
  39256=>"010100110",
  39257=>"010111010",
  39258=>"010011011",
  39259=>"001101011",
  39260=>"100110011",
  39261=>"010010000",
  39262=>"010101101",
  39263=>"010001101",
  39264=>"110110010",
  39265=>"000001100",
  39266=>"110101001",
  39267=>"000101011",
  39268=>"011001110",
  39269=>"010101100",
  39270=>"010011011",
  39271=>"111101000",
  39272=>"010001110",
  39273=>"110110000",
  39274=>"110100000",
  39275=>"000010010",
  39276=>"011000111",
  39277=>"010110111",
  39278=>"111110010",
  39279=>"000101011",
  39280=>"010010010",
  39281=>"101100110",
  39282=>"000000010",
  39283=>"101000100",
  39284=>"101101011",
  39285=>"101101010",
  39286=>"010100110",
  39287=>"111000110",
  39288=>"000001000",
  39289=>"000101101",
  39290=>"111100001",
  39291=>"010101111",
  39292=>"101000010",
  39293=>"000101010",
  39294=>"010100011",
  39295=>"011101111",
  39296=>"111011110",
  39297=>"111001101",
  39298=>"000101100",
  39299=>"001000010",
  39300=>"010111011",
  39301=>"100000101",
  39302=>"111111010",
  39303=>"110111100",
  39304=>"101101110",
  39305=>"000011110",
  39306=>"110111110",
  39307=>"100001100",
  39308=>"111100000",
  39309=>"101011100",
  39310=>"000101000",
  39311=>"000110010",
  39312=>"011111010",
  39313=>"011100100",
  39314=>"011100111",
  39315=>"101011100",
  39316=>"111000111",
  39317=>"011000011",
  39318=>"010010111",
  39319=>"011000000",
  39320=>"100000000",
  39321=>"001101100",
  39322=>"101001010",
  39323=>"111010100",
  39324=>"100111100",
  39325=>"000101110",
  39326=>"011001011",
  39327=>"001000001",
  39328=>"100010101",
  39329=>"010000011",
  39330=>"001010000",
  39331=>"001111010",
  39332=>"110010000",
  39333=>"110001010",
  39334=>"000010110",
  39335=>"110111011",
  39336=>"000101100",
  39337=>"111100100",
  39338=>"011011100",
  39339=>"111001111",
  39340=>"110111111",
  39341=>"101011101",
  39342=>"111001011",
  39343=>"010001011",
  39344=>"000001000",
  39345=>"000010001",
  39346=>"100110110",
  39347=>"000001110",
  39348=>"011111001",
  39349=>"111010101",
  39350=>"111011110",
  39351=>"111110011",
  39352=>"001110001",
  39353=>"011001110",
  39354=>"100111001",
  39355=>"010111110",
  39356=>"001010011",
  39357=>"111001101",
  39358=>"001000100",
  39359=>"000100101",
  39360=>"001001110",
  39361=>"100011111",
  39362=>"000110111",
  39363=>"101110011",
  39364=>"101110001",
  39365=>"100101110",
  39366=>"001000001",
  39367=>"000101100",
  39368=>"100000111",
  39369=>"001100111",
  39370=>"101110000",
  39371=>"111111011",
  39372=>"011111110",
  39373=>"100001010",
  39374=>"010111000",
  39375=>"101111011",
  39376=>"000011101",
  39377=>"011011110",
  39378=>"010011000",
  39379=>"111001000",
  39380=>"011100000",
  39381=>"011000111",
  39382=>"010000110",
  39383=>"001101001",
  39384=>"011010010",
  39385=>"001001010",
  39386=>"101110101",
  39387=>"011110101",
  39388=>"001010011",
  39389=>"000011010",
  39390=>"000110100",
  39391=>"100101011",
  39392=>"111011111",
  39393=>"101101000",
  39394=>"111111000",
  39395=>"011100010",
  39396=>"000110001",
  39397=>"010100011",
  39398=>"000001100",
  39399=>"001000001",
  39400=>"000010110",
  39401=>"001100011",
  39402=>"011000101",
  39403=>"011011110",
  39404=>"110110011",
  39405=>"010110100",
  39406=>"101101101",
  39407=>"011100111",
  39408=>"001111011",
  39409=>"101101111",
  39410=>"111111001",
  39411=>"000001000",
  39412=>"101000111",
  39413=>"100011001",
  39414=>"110111010",
  39415=>"000101111",
  39416=>"101011101",
  39417=>"110011101",
  39418=>"000010111",
  39419=>"101101001",
  39420=>"001110100",
  39421=>"110000010",
  39422=>"101100110",
  39423=>"011111111",
  39424=>"010000000",
  39425=>"101000010",
  39426=>"101111101",
  39427=>"100001001",
  39428=>"010110110",
  39429=>"001000001",
  39430=>"111101111",
  39431=>"110111100",
  39432=>"100000001",
  39433=>"111011101",
  39434=>"010000001",
  39435=>"110010010",
  39436=>"001100111",
  39437=>"111011100",
  39438=>"100000001",
  39439=>"101111110",
  39440=>"100111101",
  39441=>"111111000",
  39442=>"110111110",
  39443=>"101100110",
  39444=>"011000110",
  39445=>"100100011",
  39446=>"110001101",
  39447=>"010001001",
  39448=>"001000010",
  39449=>"101011000",
  39450=>"110000110",
  39451=>"010000111",
  39452=>"010001100",
  39453=>"110110111",
  39454=>"100010011",
  39455=>"110010100",
  39456=>"011101000",
  39457=>"101000111",
  39458=>"001010100",
  39459=>"010100110",
  39460=>"101011110",
  39461=>"000001001",
  39462=>"101101000",
  39463=>"010100101",
  39464=>"000010001",
  39465=>"111101011",
  39466=>"010001110",
  39467=>"110000110",
  39468=>"110010000",
  39469=>"110100100",
  39470=>"101111000",
  39471=>"101001110",
  39472=>"111010011",
  39473=>"111100100",
  39474=>"100110111",
  39475=>"001001100",
  39476=>"010000011",
  39477=>"111100000",
  39478=>"010111110",
  39479=>"000010000",
  39480=>"110111100",
  39481=>"110111010",
  39482=>"101000100",
  39483=>"100100011",
  39484=>"101110110",
  39485=>"101001001",
  39486=>"110101001",
  39487=>"000101100",
  39488=>"000001011",
  39489=>"010101001",
  39490=>"101100101",
  39491=>"010110000",
  39492=>"111111111",
  39493=>"110010011",
  39494=>"100010010",
  39495=>"111010011",
  39496=>"100100111",
  39497=>"110000100",
  39498=>"111101110",
  39499=>"111101111",
  39500=>"100110011",
  39501=>"110101001",
  39502=>"000011000",
  39503=>"101100001",
  39504=>"001001000",
  39505=>"011000110",
  39506=>"000101011",
  39507=>"100111001",
  39508=>"110010010",
  39509=>"001010110",
  39510=>"111100101",
  39511=>"000000010",
  39512=>"010101111",
  39513=>"111111100",
  39514=>"110010001",
  39515=>"110100111",
  39516=>"001000001",
  39517=>"101001011",
  39518=>"011100010",
  39519=>"110001101",
  39520=>"010000010",
  39521=>"101101001",
  39522=>"111000001",
  39523=>"000011000",
  39524=>"110011001",
  39525=>"110001011",
  39526=>"100010110",
  39527=>"000010011",
  39528=>"100111100",
  39529=>"000001010",
  39530=>"001010101",
  39531=>"001111011",
  39532=>"101001111",
  39533=>"011100110",
  39534=>"000110110",
  39535=>"110011001",
  39536=>"111101101",
  39537=>"111100000",
  39538=>"110110111",
  39539=>"101001110",
  39540=>"010101000",
  39541=>"100000010",
  39542=>"011010010",
  39543=>"100001000",
  39544=>"000110010",
  39545=>"000000000",
  39546=>"110011010",
  39547=>"000000110",
  39548=>"111000011",
  39549=>"000100001",
  39550=>"011111111",
  39551=>"111110111",
  39552=>"001100000",
  39553=>"011110101",
  39554=>"011111010",
  39555=>"100011110",
  39556=>"110011111",
  39557=>"101001001",
  39558=>"110000111",
  39559=>"110011111",
  39560=>"010101100",
  39561=>"101000100",
  39562=>"101110110",
  39563=>"100111011",
  39564=>"101000110",
  39565=>"100001011",
  39566=>"011111101",
  39567=>"100101011",
  39568=>"000010101",
  39569=>"000010100",
  39570=>"101001010",
  39571=>"111100111",
  39572=>"000110001",
  39573=>"100111111",
  39574=>"000100111",
  39575=>"100100000",
  39576=>"011001001",
  39577=>"110001111",
  39578=>"000101110",
  39579=>"001100101",
  39580=>"110010100",
  39581=>"111100110",
  39582=>"000010110",
  39583=>"011000110",
  39584=>"110100110",
  39585=>"111000000",
  39586=>"100111110",
  39587=>"000011111",
  39588=>"101101101",
  39589=>"010110001",
  39590=>"100000010",
  39591=>"101111111",
  39592=>"000110111",
  39593=>"000111011",
  39594=>"101101000",
  39595=>"110101010",
  39596=>"011101000",
  39597=>"100100010",
  39598=>"101010010",
  39599=>"110110110",
  39600=>"111110100",
  39601=>"101001101",
  39602=>"001111111",
  39603=>"110000011",
  39604=>"010000011",
  39605=>"011101001",
  39606=>"011111101",
  39607=>"101110111",
  39608=>"010100010",
  39609=>"111010100",
  39610=>"010010111",
  39611=>"100010001",
  39612=>"010100111",
  39613=>"011001001",
  39614=>"110011000",
  39615=>"101011100",
  39616=>"100011001",
  39617=>"100101111",
  39618=>"011100111",
  39619=>"110101110",
  39620=>"110111100",
  39621=>"011101100",
  39622=>"110001100",
  39623=>"001111000",
  39624=>"010000000",
  39625=>"010000011",
  39626=>"011001011",
  39627=>"001011001",
  39628=>"101101110",
  39629=>"000101111",
  39630=>"111000001",
  39631=>"111100111",
  39632=>"010110111",
  39633=>"000111111",
  39634=>"110011101",
  39635=>"001000110",
  39636=>"001111100",
  39637=>"010000011",
  39638=>"110010101",
  39639=>"011110010",
  39640=>"100010101",
  39641=>"111100011",
  39642=>"111111001",
  39643=>"000001110",
  39644=>"111101111",
  39645=>"011010110",
  39646=>"111000111",
  39647=>"010001010",
  39648=>"111111010",
  39649=>"111101010",
  39650=>"110011100",
  39651=>"001001010",
  39652=>"010001000",
  39653=>"011100101",
  39654=>"011100000",
  39655=>"111001000",
  39656=>"011111010",
  39657=>"011001111",
  39658=>"001000000",
  39659=>"111011010",
  39660=>"011111000",
  39661=>"101100110",
  39662=>"000101111",
  39663=>"010100101",
  39664=>"101000000",
  39665=>"101111010",
  39666=>"011111011",
  39667=>"000011001",
  39668=>"011000110",
  39669=>"000001111",
  39670=>"000011001",
  39671=>"101111100",
  39672=>"010110110",
  39673=>"000010000",
  39674=>"111101100",
  39675=>"010000001",
  39676=>"000001111",
  39677=>"011010001",
  39678=>"101001110",
  39679=>"110001111",
  39680=>"100000111",
  39681=>"011010101",
  39682=>"100100110",
  39683=>"011000100",
  39684=>"100010010",
  39685=>"000110011",
  39686=>"000100110",
  39687=>"101000001",
  39688=>"110010111",
  39689=>"010100011",
  39690=>"000111011",
  39691=>"000010100",
  39692=>"011001000",
  39693=>"110110010",
  39694=>"100101010",
  39695=>"101111111",
  39696=>"101101111",
  39697=>"010110011",
  39698=>"100010101",
  39699=>"001110100",
  39700=>"100110001",
  39701=>"011111011",
  39702=>"110110011",
  39703=>"010100101",
  39704=>"111111010",
  39705=>"010001010",
  39706=>"000111101",
  39707=>"011001001",
  39708=>"010001000",
  39709=>"000110111",
  39710=>"010111110",
  39711=>"001001010",
  39712=>"011000111",
  39713=>"111000010",
  39714=>"010100101",
  39715=>"000110010",
  39716=>"001111111",
  39717=>"111000000",
  39718=>"110001010",
  39719=>"111110011",
  39720=>"000110111",
  39721=>"101011100",
  39722=>"000101011",
  39723=>"001111111",
  39724=>"001100101",
  39725=>"111100111",
  39726=>"101110101",
  39727=>"010001001",
  39728=>"010010010",
  39729=>"100100001",
  39730=>"011101001",
  39731=>"011001101",
  39732=>"101100100",
  39733=>"011110110",
  39734=>"000001000",
  39735=>"110001000",
  39736=>"000100001",
  39737=>"000010001",
  39738=>"110100111",
  39739=>"010101010",
  39740=>"001010101",
  39741=>"000110001",
  39742=>"010101000",
  39743=>"101100000",
  39744=>"100001101",
  39745=>"111111110",
  39746=>"110100111",
  39747=>"110111000",
  39748=>"010111101",
  39749=>"011010001",
  39750=>"010010111",
  39751=>"001000010",
  39752=>"000010101",
  39753=>"000111101",
  39754=>"110101001",
  39755=>"111100111",
  39756=>"011110110",
  39757=>"100100110",
  39758=>"010100000",
  39759=>"100101101",
  39760=>"100111000",
  39761=>"111011110",
  39762=>"001111110",
  39763=>"110010110",
  39764=>"000011011",
  39765=>"111111111",
  39766=>"100111101",
  39767=>"000010101",
  39768=>"001000010",
  39769=>"011111100",
  39770=>"101000010",
  39771=>"110101000",
  39772=>"110101010",
  39773=>"111101000",
  39774=>"011101110",
  39775=>"100010000",
  39776=>"110111001",
  39777=>"000001110",
  39778=>"110110001",
  39779=>"110000001",
  39780=>"010110101",
  39781=>"111110111",
  39782=>"010001011",
  39783=>"110011011",
  39784=>"111001100",
  39785=>"101101101",
  39786=>"010000001",
  39787=>"010101100",
  39788=>"110011000",
  39789=>"011000010",
  39790=>"001101001",
  39791=>"001001110",
  39792=>"110100011",
  39793=>"010101001",
  39794=>"101110101",
  39795=>"001110010",
  39796=>"010010110",
  39797=>"111011001",
  39798=>"101001110",
  39799=>"111100010",
  39800=>"001011111",
  39801=>"100010111",
  39802=>"010100001",
  39803=>"000011000",
  39804=>"010000010",
  39805=>"100011101",
  39806=>"110110000",
  39807=>"110011000",
  39808=>"101010001",
  39809=>"011011101",
  39810=>"000001001",
  39811=>"011110010",
  39812=>"010000101",
  39813=>"110101010",
  39814=>"110100111",
  39815=>"001000101",
  39816=>"001001001",
  39817=>"000000110",
  39818=>"000100010",
  39819=>"110111111",
  39820=>"101010100",
  39821=>"011110111",
  39822=>"101101010",
  39823=>"010111100",
  39824=>"100100111",
  39825=>"011000110",
  39826=>"000011001",
  39827=>"010110111",
  39828=>"100101100",
  39829=>"100110011",
  39830=>"101111100",
  39831=>"011111000",
  39832=>"010000001",
  39833=>"111111000",
  39834=>"000100100",
  39835=>"100110101",
  39836=>"000001010",
  39837=>"000101000",
  39838=>"010011101",
  39839=>"001010011",
  39840=>"000000111",
  39841=>"111101110",
  39842=>"111111010",
  39843=>"101100011",
  39844=>"000010100",
  39845=>"111110101",
  39846=>"000001101",
  39847=>"001010110",
  39848=>"110001000",
  39849=>"111000100",
  39850=>"000110001",
  39851=>"011010101",
  39852=>"101011111",
  39853=>"110101100",
  39854=>"000000111",
  39855=>"110100111",
  39856=>"001101010",
  39857=>"110100001",
  39858=>"101101111",
  39859=>"100101001",
  39860=>"111101101",
  39861=>"000111101",
  39862=>"000000111",
  39863=>"100111101",
  39864=>"010010110",
  39865=>"010101001",
  39866=>"001100010",
  39867=>"000010010",
  39868=>"101101101",
  39869=>"000010000",
  39870=>"110110010",
  39871=>"000111101",
  39872=>"000110101",
  39873=>"000011010",
  39874=>"011001001",
  39875=>"110010100",
  39876=>"010010010",
  39877=>"001101010",
  39878=>"010101101",
  39879=>"000000111",
  39880=>"011000010",
  39881=>"100101001",
  39882=>"111000010",
  39883=>"110110010",
  39884=>"110110110",
  39885=>"111010001",
  39886=>"000100110",
  39887=>"100010000",
  39888=>"000101111",
  39889=>"011100110",
  39890=>"110011110",
  39891=>"111000000",
  39892=>"011111011",
  39893=>"001111011",
  39894=>"000000011",
  39895=>"111110100",
  39896=>"010000100",
  39897=>"111010001",
  39898=>"100110111",
  39899=>"011111111",
  39900=>"110101101",
  39901=>"011110000",
  39902=>"000001111",
  39903=>"100100101",
  39904=>"000001001",
  39905=>"110110000",
  39906=>"100001110",
  39907=>"000101110",
  39908=>"110001001",
  39909=>"100000001",
  39910=>"101100000",
  39911=>"101111001",
  39912=>"011000000",
  39913=>"111111000",
  39914=>"010110110",
  39915=>"010000100",
  39916=>"011000011",
  39917=>"110000111",
  39918=>"010110010",
  39919=>"011000001",
  39920=>"000110010",
  39921=>"000010001",
  39922=>"101000111",
  39923=>"010001001",
  39924=>"101011010",
  39925=>"001011000",
  39926=>"101001000",
  39927=>"011001100",
  39928=>"001010101",
  39929=>"100000100",
  39930=>"111001100",
  39931=>"111101100",
  39932=>"110101111",
  39933=>"100000010",
  39934=>"010001001",
  39935=>"010111011",
  39936=>"111111111",
  39937=>"001001011",
  39938=>"011011011",
  39939=>"010110000",
  39940=>"110010001",
  39941=>"110011001",
  39942=>"000111010",
  39943=>"000110000",
  39944=>"100001011",
  39945=>"100001101",
  39946=>"001111111",
  39947=>"111100000",
  39948=>"110010101",
  39949=>"010110001",
  39950=>"110011110",
  39951=>"111000001",
  39952=>"110011001",
  39953=>"010100001",
  39954=>"010010101",
  39955=>"010001011",
  39956=>"001110000",
  39957=>"011001101",
  39958=>"001100101",
  39959=>"010001100",
  39960=>"110001101",
  39961=>"111000111",
  39962=>"011111110",
  39963=>"011011111",
  39964=>"100011000",
  39965=>"001100110",
  39966=>"011001000",
  39967=>"101010000",
  39968=>"000000000",
  39969=>"010111000",
  39970=>"000011010",
  39971=>"001011110",
  39972=>"100000011",
  39973=>"001001111",
  39974=>"001101010",
  39975=>"000101011",
  39976=>"011001000",
  39977=>"000100101",
  39978=>"010100001",
  39979=>"100110100",
  39980=>"011100101",
  39981=>"011101001",
  39982=>"111101001",
  39983=>"010110100",
  39984=>"111010000",
  39985=>"011000100",
  39986=>"101111010",
  39987=>"011100010",
  39988=>"010100001",
  39989=>"011101010",
  39990=>"000001111",
  39991=>"010100001",
  39992=>"010101100",
  39993=>"110010001",
  39994=>"010000111",
  39995=>"101101000",
  39996=>"010001001",
  39997=>"111101011",
  39998=>"110010010",
  39999=>"100110111",
  40000=>"100111111",
  40001=>"011001101",
  40002=>"101000100",
  40003=>"000110110",
  40004=>"101101001",
  40005=>"010001111",
  40006=>"001000101",
  40007=>"100010101",
  40008=>"101011111",
  40009=>"010001001",
  40010=>"000000001",
  40011=>"101010001",
  40012=>"111101011",
  40013=>"110100100",
  40014=>"010100111",
  40015=>"100111110",
  40016=>"011111011",
  40017=>"000011000",
  40018=>"100110101",
  40019=>"111111110",
  40020=>"000111011",
  40021=>"100010010",
  40022=>"001000110",
  40023=>"001001111",
  40024=>"110011111",
  40025=>"010001101",
  40026=>"011010000",
  40027=>"001001110",
  40028=>"100100011",
  40029=>"000111101",
  40030=>"010011011",
  40031=>"010111111",
  40032=>"011110111",
  40033=>"110000001",
  40034=>"011001110",
  40035=>"001101101",
  40036=>"110000000",
  40037=>"010011011",
  40038=>"111000011",
  40039=>"100111110",
  40040=>"001111100",
  40041=>"111101011",
  40042=>"000000000",
  40043=>"011010001",
  40044=>"101100101",
  40045=>"000010101",
  40046=>"000001000",
  40047=>"000011000",
  40048=>"100011011",
  40049=>"111111100",
  40050=>"010001000",
  40051=>"101111010",
  40052=>"000110011",
  40053=>"010101110",
  40054=>"111011111",
  40055=>"111001111",
  40056=>"101100110",
  40057=>"101101000",
  40058=>"101011100",
  40059=>"001001010",
  40060=>"011100001",
  40061=>"011100100",
  40062=>"000011001",
  40063=>"001000110",
  40064=>"101001001",
  40065=>"000100110",
  40066=>"010010110",
  40067=>"110000111",
  40068=>"100110111",
  40069=>"010000000",
  40070=>"011000000",
  40071=>"111100011",
  40072=>"111111110",
  40073=>"000010011",
  40074=>"100101110",
  40075=>"101011000",
  40076=>"000001110",
  40077=>"100011010",
  40078=>"110000011",
  40079=>"100100011",
  40080=>"111001000",
  40081=>"010101111",
  40082=>"110101000",
  40083=>"101010111",
  40084=>"011111001",
  40085=>"111010110",
  40086=>"111111001",
  40087=>"101010011",
  40088=>"010001010",
  40089=>"110001101",
  40090=>"111110001",
  40091=>"011010011",
  40092=>"001110101",
  40093=>"101011010",
  40094=>"010111000",
  40095=>"111110001",
  40096=>"100110010",
  40097=>"001000100",
  40098=>"100101110",
  40099=>"111110001",
  40100=>"011111100",
  40101=>"000111010",
  40102=>"010110011",
  40103=>"111001011",
  40104=>"011010001",
  40105=>"111010001",
  40106=>"010100110",
  40107=>"000001011",
  40108=>"011111110",
  40109=>"111111010",
  40110=>"001011000",
  40111=>"000100001",
  40112=>"010110001",
  40113=>"001000110",
  40114=>"110100111",
  40115=>"101000110",
  40116=>"100111111",
  40117=>"110110010",
  40118=>"101000110",
  40119=>"000101110",
  40120=>"001000001",
  40121=>"101101100",
  40122=>"001100100",
  40123=>"010101100",
  40124=>"100101011",
  40125=>"001001101",
  40126=>"010010100",
  40127=>"111110110",
  40128=>"011001101",
  40129=>"100001111",
  40130=>"000100110",
  40131=>"101111101",
  40132=>"111011010",
  40133=>"011110010",
  40134=>"011110000",
  40135=>"100110001",
  40136=>"111111011",
  40137=>"111100111",
  40138=>"010111110",
  40139=>"001110100",
  40140=>"111001111",
  40141=>"111111000",
  40142=>"111010111",
  40143=>"011000111",
  40144=>"001000000",
  40145=>"010000110",
  40146=>"100101100",
  40147=>"000111000",
  40148=>"101001111",
  40149=>"000100101",
  40150=>"100011001",
  40151=>"001111010",
  40152=>"101010010",
  40153=>"100100001",
  40154=>"100010000",
  40155=>"000000000",
  40156=>"011110001",
  40157=>"001100011",
  40158=>"000001101",
  40159=>"000100100",
  40160=>"000001000",
  40161=>"010000011",
  40162=>"001010100",
  40163=>"001001110",
  40164=>"111000011",
  40165=>"010011001",
  40166=>"010111001",
  40167=>"010111111",
  40168=>"010100010",
  40169=>"000111011",
  40170=>"101011000",
  40171=>"101001100",
  40172=>"100101100",
  40173=>"100110100",
  40174=>"001011001",
  40175=>"001010110",
  40176=>"011011001",
  40177=>"110010100",
  40178=>"011001111",
  40179=>"000100011",
  40180=>"001100100",
  40181=>"010100001",
  40182=>"000101011",
  40183=>"101101110",
  40184=>"011001011",
  40185=>"111110111",
  40186=>"110000001",
  40187=>"011010110",
  40188=>"001111101",
  40189=>"110000000",
  40190=>"101001110",
  40191=>"101011111",
  40192=>"111011110",
  40193=>"100000111",
  40194=>"100000110",
  40195=>"110000000",
  40196=>"110100101",
  40197=>"001100101",
  40198=>"000010100",
  40199=>"000001010",
  40200=>"111011000",
  40201=>"000011010",
  40202=>"111110100",
  40203=>"100101001",
  40204=>"011100101",
  40205=>"011101010",
  40206=>"110100100",
  40207=>"011001001",
  40208=>"011000101",
  40209=>"110100001",
  40210=>"011101110",
  40211=>"010100101",
  40212=>"001110011",
  40213=>"101110101",
  40214=>"111111011",
  40215=>"000011111",
  40216=>"110001101",
  40217=>"100111111",
  40218=>"001110010",
  40219=>"011101110",
  40220=>"001001111",
  40221=>"000101000",
  40222=>"110111101",
  40223=>"000111001",
  40224=>"100011110",
  40225=>"100101110",
  40226=>"011000011",
  40227=>"001010101",
  40228=>"111101101",
  40229=>"101010001",
  40230=>"001101101",
  40231=>"101111000",
  40232=>"000111100",
  40233=>"001000110",
  40234=>"101001010",
  40235=>"001101100",
  40236=>"101001001",
  40237=>"101101111",
  40238=>"010001010",
  40239=>"111000111",
  40240=>"010001001",
  40241=>"110010100",
  40242=>"100111010",
  40243=>"000000110",
  40244=>"010100011",
  40245=>"001100111",
  40246=>"101100011",
  40247=>"100010111",
  40248=>"110100101",
  40249=>"111101101",
  40250=>"100101101",
  40251=>"000100011",
  40252=>"111001000",
  40253=>"001010100",
  40254=>"101001101",
  40255=>"111000011",
  40256=>"001101000",
  40257=>"111100010",
  40258=>"111100001",
  40259=>"011101111",
  40260=>"110000011",
  40261=>"000101011",
  40262=>"110000110",
  40263=>"110001001",
  40264=>"111000010",
  40265=>"001011001",
  40266=>"101010010",
  40267=>"001100111",
  40268=>"100110111",
  40269=>"010010110",
  40270=>"000001100",
  40271=>"000110111",
  40272=>"111100011",
  40273=>"011011110",
  40274=>"000110100",
  40275=>"000001110",
  40276=>"101101100",
  40277=>"000111011",
  40278=>"110010000",
  40279=>"110100101",
  40280=>"000111010",
  40281=>"000110011",
  40282=>"110011110",
  40283=>"011010010",
  40284=>"011111111",
  40285=>"100110100",
  40286=>"111001110",
  40287=>"100111101",
  40288=>"101001100",
  40289=>"010010001",
  40290=>"110010010",
  40291=>"010011111",
  40292=>"001111001",
  40293=>"011101010",
  40294=>"100001100",
  40295=>"000011000",
  40296=>"100100011",
  40297=>"111001001",
  40298=>"000101110",
  40299=>"000000010",
  40300=>"000111100",
  40301=>"111001110",
  40302=>"011000110",
  40303=>"110010100",
  40304=>"100111110",
  40305=>"001011001",
  40306=>"100001001",
  40307=>"010010011",
  40308=>"000001011",
  40309=>"101001100",
  40310=>"100111011",
  40311=>"100000111",
  40312=>"001010101",
  40313=>"001000001",
  40314=>"010111000",
  40315=>"111111011",
  40316=>"100001001",
  40317=>"010010111",
  40318=>"011001110",
  40319=>"101010100",
  40320=>"000001001",
  40321=>"010000100",
  40322=>"000111101",
  40323=>"101110110",
  40324=>"001001011",
  40325=>"001111011",
  40326=>"101100111",
  40327=>"011100101",
  40328=>"101001101",
  40329=>"000101111",
  40330=>"101110110",
  40331=>"000101111",
  40332=>"111101111",
  40333=>"001011101",
  40334=>"101001101",
  40335=>"111000000",
  40336=>"101000111",
  40337=>"000010100",
  40338=>"001010100",
  40339=>"001011000",
  40340=>"100011000",
  40341=>"001111001",
  40342=>"111010101",
  40343=>"101011100",
  40344=>"000111100",
  40345=>"110000000",
  40346=>"110100010",
  40347=>"100010101",
  40348=>"100100011",
  40349=>"001010111",
  40350=>"000001100",
  40351=>"111111110",
  40352=>"010100010",
  40353=>"011011001",
  40354=>"000111000",
  40355=>"011011001",
  40356=>"011110111",
  40357=>"000000100",
  40358=>"011000000",
  40359=>"001100010",
  40360=>"001001101",
  40361=>"010001111",
  40362=>"100100111",
  40363=>"011010100",
  40364=>"110111111",
  40365=>"010011110",
  40366=>"000000111",
  40367=>"100101011",
  40368=>"011110000",
  40369=>"001001100",
  40370=>"111110100",
  40371=>"101011110",
  40372=>"011001010",
  40373=>"001000001",
  40374=>"000100011",
  40375=>"110011101",
  40376=>"100100010",
  40377=>"100111101",
  40378=>"010101111",
  40379=>"100111110",
  40380=>"101101100",
  40381=>"001101111",
  40382=>"110101111",
  40383=>"110111011",
  40384=>"100100111",
  40385=>"010110010",
  40386=>"110000111",
  40387=>"001011001",
  40388=>"010100010",
  40389=>"001110010",
  40390=>"110010100",
  40391=>"101001001",
  40392=>"011111111",
  40393=>"111000011",
  40394=>"011000111",
  40395=>"110101111",
  40396=>"101000101",
  40397=>"110101100",
  40398=>"101000010",
  40399=>"110101001",
  40400=>"000010010",
  40401=>"001110000",
  40402=>"000101010",
  40403=>"111100000",
  40404=>"101011101",
  40405=>"101001000",
  40406=>"101101000",
  40407=>"101111010",
  40408=>"011000010",
  40409=>"000010011",
  40410=>"001011101",
  40411=>"101100001",
  40412=>"101100111",
  40413=>"011111001",
  40414=>"001110011",
  40415=>"001110100",
  40416=>"011101011",
  40417=>"011101010",
  40418=>"100100101",
  40419=>"011101101",
  40420=>"111010101",
  40421=>"111001011",
  40422=>"011001110",
  40423=>"110101000",
  40424=>"111000100",
  40425=>"010010011",
  40426=>"100001001",
  40427=>"001101010",
  40428=>"010101000",
  40429=>"010001000",
  40430=>"100111000",
  40431=>"011001001",
  40432=>"001100110",
  40433=>"001111000",
  40434=>"011011011",
  40435=>"101001011",
  40436=>"111001110",
  40437=>"010100100",
  40438=>"011000100",
  40439=>"111100000",
  40440=>"110010110",
  40441=>"011010011",
  40442=>"010111101",
  40443=>"110001011",
  40444=>"011010100",
  40445=>"000101101",
  40446=>"010001100",
  40447=>"111111000",
  40448=>"101111111",
  40449=>"100011010",
  40450=>"011000010",
  40451=>"100010100",
  40452=>"001000010",
  40453=>"101100100",
  40454=>"110100000",
  40455=>"100101101",
  40456=>"001001001",
  40457=>"110110011",
  40458=>"011010000",
  40459=>"111111000",
  40460=>"100111000",
  40461=>"001101110",
  40462=>"100000100",
  40463=>"111111110",
  40464=>"111000110",
  40465=>"111111010",
  40466=>"001100000",
  40467=>"101111111",
  40468=>"111100100",
  40469=>"000011011",
  40470=>"110010100",
  40471=>"010101000",
  40472=>"010100100",
  40473=>"011011011",
  40474=>"111111110",
  40475=>"000110100",
  40476=>"111110101",
  40477=>"111000111",
  40478=>"100110010",
  40479=>"000101001",
  40480=>"110001011",
  40481=>"010001101",
  40482=>"001011110",
  40483=>"000010001",
  40484=>"111100100",
  40485=>"110011110",
  40486=>"110010110",
  40487=>"100110000",
  40488=>"100000101",
  40489=>"111000011",
  40490=>"001111010",
  40491=>"101100000",
  40492=>"001010111",
  40493=>"100110000",
  40494=>"011110010",
  40495=>"110101000",
  40496=>"100000010",
  40497=>"000001001",
  40498=>"011110110",
  40499=>"011101000",
  40500=>"010001101",
  40501=>"111101100",
  40502=>"001011010",
  40503=>"011001101",
  40504=>"000010010",
  40505=>"001101011",
  40506=>"101100110",
  40507=>"101001111",
  40508=>"111100011",
  40509=>"000010010",
  40510=>"011100001",
  40511=>"010001001",
  40512=>"011110010",
  40513=>"111111101",
  40514=>"110001100",
  40515=>"101100010",
  40516=>"100101100",
  40517=>"011010000",
  40518=>"001111010",
  40519=>"100110011",
  40520=>"100010111",
  40521=>"010000000",
  40522=>"101010011",
  40523=>"011000100",
  40524=>"101001111",
  40525=>"011000010",
  40526=>"000011100",
  40527=>"011010000",
  40528=>"100110011",
  40529=>"111000001",
  40530=>"100101001",
  40531=>"001100101",
  40532=>"110110110",
  40533=>"100100101",
  40534=>"101010001",
  40535=>"100001100",
  40536=>"100101010",
  40537=>"110011000",
  40538=>"111000000",
  40539=>"001001100",
  40540=>"001011000",
  40541=>"011000011",
  40542=>"000011101",
  40543=>"111100100",
  40544=>"110001010",
  40545=>"011100001",
  40546=>"111101101",
  40547=>"100100000",
  40548=>"100010111",
  40549=>"010111100",
  40550=>"101010100",
  40551=>"011111101",
  40552=>"100010110",
  40553=>"001010101",
  40554=>"100011101",
  40555=>"110010100",
  40556=>"000001011",
  40557=>"010010111",
  40558=>"100011001",
  40559=>"111110001",
  40560=>"111010000",
  40561=>"110100100",
  40562=>"100100010",
  40563=>"010011111",
  40564=>"000001000",
  40565=>"110000100",
  40566=>"001011110",
  40567=>"110101101",
  40568=>"111111010",
  40569=>"000010000",
  40570=>"100001011",
  40571=>"110111000",
  40572=>"001000011",
  40573=>"100000000",
  40574=>"000110011",
  40575=>"101000101",
  40576=>"111111111",
  40577=>"111010110",
  40578=>"101101101",
  40579=>"010000100",
  40580=>"111111111",
  40581=>"101100110",
  40582=>"100110010",
  40583=>"010110011",
  40584=>"001000101",
  40585=>"101001100",
  40586=>"100110000",
  40587=>"001011010",
  40588=>"100001000",
  40589=>"111011010",
  40590=>"010101010",
  40591=>"000010011",
  40592=>"110100001",
  40593=>"110101010",
  40594=>"100000000",
  40595=>"101110100",
  40596=>"101010110",
  40597=>"100100101",
  40598=>"011110101",
  40599=>"001010000",
  40600=>"000110100",
  40601=>"011011010",
  40602=>"011111101",
  40603=>"011011110",
  40604=>"111000101",
  40605=>"101011110",
  40606=>"100100111",
  40607=>"001110010",
  40608=>"111100001",
  40609=>"100110111",
  40610=>"010111010",
  40611=>"010110001",
  40612=>"111001011",
  40613=>"000011101",
  40614=>"000110011",
  40615=>"000101001",
  40616=>"011111101",
  40617=>"101010001",
  40618=>"111001110",
  40619=>"001101010",
  40620=>"010111101",
  40621=>"101110001",
  40622=>"111011111",
  40623=>"101001101",
  40624=>"010110000",
  40625=>"000100010",
  40626=>"011101000",
  40627=>"010001010",
  40628=>"011110011",
  40629=>"000100110",
  40630=>"100000000",
  40631=>"011101011",
  40632=>"100010011",
  40633=>"011010111",
  40634=>"100111101",
  40635=>"111000110",
  40636=>"011010001",
  40637=>"010111100",
  40638=>"101000001",
  40639=>"000010000",
  40640=>"000010010",
  40641=>"111110111",
  40642=>"001000101",
  40643=>"010111001",
  40644=>"101101100",
  40645=>"011001010",
  40646=>"001010000",
  40647=>"101000110",
  40648=>"111111001",
  40649=>"001100001",
  40650=>"000011011",
  40651=>"011000011",
  40652=>"100111001",
  40653=>"110010101",
  40654=>"101001111",
  40655=>"110111101",
  40656=>"010101011",
  40657=>"011000000",
  40658=>"010011010",
  40659=>"111101110",
  40660=>"110101101",
  40661=>"111011000",
  40662=>"010111101",
  40663=>"001011101",
  40664=>"010000110",
  40665=>"101010001",
  40666=>"011101111",
  40667=>"000000111",
  40668=>"111101001",
  40669=>"111111001",
  40670=>"000101110",
  40671=>"111010000",
  40672=>"011110100",
  40673=>"101100001",
  40674=>"111010111",
  40675=>"100001000",
  40676=>"111111000",
  40677=>"010000100",
  40678=>"000000011",
  40679=>"011101111",
  40680=>"000010101",
  40681=>"110010111",
  40682=>"110111000",
  40683=>"010111011",
  40684=>"100000100",
  40685=>"000000001",
  40686=>"001010001",
  40687=>"101010100",
  40688=>"110110111",
  40689=>"000111110",
  40690=>"000000000",
  40691=>"001100011",
  40692=>"011101010",
  40693=>"011111100",
  40694=>"101001101",
  40695=>"101001100",
  40696=>"111000100",
  40697=>"111101101",
  40698=>"000011001",
  40699=>"000100010",
  40700=>"101000100",
  40701=>"010000110",
  40702=>"001001011",
  40703=>"000101001",
  40704=>"010001010",
  40705=>"000100111",
  40706=>"011001111",
  40707=>"011001001",
  40708=>"000010011",
  40709=>"100000110",
  40710=>"001000101",
  40711=>"110111110",
  40712=>"010010111",
  40713=>"100011011",
  40714=>"010100010",
  40715=>"111101110",
  40716=>"010011111",
  40717=>"000000100",
  40718=>"101010101",
  40719=>"000101100",
  40720=>"110000000",
  40721=>"000010101",
  40722=>"010111111",
  40723=>"110000000",
  40724=>"011010100",
  40725=>"110111011",
  40726=>"100001101",
  40727=>"100010100",
  40728=>"110011011",
  40729=>"000111001",
  40730=>"110111010",
  40731=>"011011111",
  40732=>"100100110",
  40733=>"010010000",
  40734=>"011000011",
  40735=>"110000011",
  40736=>"001111000",
  40737=>"001000000",
  40738=>"110001101",
  40739=>"000111101",
  40740=>"101010101",
  40741=>"010111111",
  40742=>"010111000",
  40743=>"111010111",
  40744=>"110111101",
  40745=>"101100011",
  40746=>"000111111",
  40747=>"100101111",
  40748=>"100010000",
  40749=>"010000000",
  40750=>"001100110",
  40751=>"111101110",
  40752=>"110000001",
  40753=>"101101111",
  40754=>"111011001",
  40755=>"011101011",
  40756=>"101101110",
  40757=>"110111010",
  40758=>"111100001",
  40759=>"110010000",
  40760=>"100010000",
  40761=>"111000101",
  40762=>"101001110",
  40763=>"110110100",
  40764=>"001001000",
  40765=>"000011000",
  40766=>"100010010",
  40767=>"010000010",
  40768=>"111101001",
  40769=>"111001000",
  40770=>"011011000",
  40771=>"101110111",
  40772=>"010111110",
  40773=>"101011010",
  40774=>"100010010",
  40775=>"100110000",
  40776=>"101110110",
  40777=>"010110101",
  40778=>"001101111",
  40779=>"010010010",
  40780=>"001101111",
  40781=>"011011111",
  40782=>"111000110",
  40783=>"111000110",
  40784=>"110010000",
  40785=>"011000111",
  40786=>"001101001",
  40787=>"101000001",
  40788=>"011010110",
  40789=>"011010101",
  40790=>"111100110",
  40791=>"000101111",
  40792=>"000001011",
  40793=>"000100100",
  40794=>"010100111",
  40795=>"100110011",
  40796=>"000011100",
  40797=>"100000000",
  40798=>"110001111",
  40799=>"110011001",
  40800=>"010000101",
  40801=>"100000010",
  40802=>"001101011",
  40803=>"111110100",
  40804=>"001001101",
  40805=>"111010001",
  40806=>"000101110",
  40807=>"111101011",
  40808=>"110101000",
  40809=>"101100110",
  40810=>"111111110",
  40811=>"111010001",
  40812=>"111110101",
  40813=>"001111101",
  40814=>"010000001",
  40815=>"110000111",
  40816=>"101010100",
  40817=>"111000010",
  40818=>"111011011",
  40819=>"111001011",
  40820=>"011101111",
  40821=>"110000111",
  40822=>"111001001",
  40823=>"000101000",
  40824=>"111001110",
  40825=>"000110011",
  40826=>"011110111",
  40827=>"010011001",
  40828=>"011011111",
  40829=>"001000000",
  40830=>"100101100",
  40831=>"001111011",
  40832=>"100100100",
  40833=>"111011011",
  40834=>"100000011",
  40835=>"111010101",
  40836=>"000010001",
  40837=>"001100010",
  40838=>"011001100",
  40839=>"101001110",
  40840=>"011100111",
  40841=>"000101111",
  40842=>"000000001",
  40843=>"000000000",
  40844=>"110100111",
  40845=>"101111110",
  40846=>"101111101",
  40847=>"111010110",
  40848=>"011100011",
  40849=>"111111011",
  40850=>"101000101",
  40851=>"101100100",
  40852=>"010001111",
  40853=>"101001100",
  40854=>"011011111",
  40855=>"000111101",
  40856=>"101001001",
  40857=>"000000100",
  40858=>"101000011",
  40859=>"010100110",
  40860=>"111000000",
  40861=>"101101110",
  40862=>"000000001",
  40863=>"111001011",
  40864=>"110110011",
  40865=>"111111011",
  40866=>"011011000",
  40867=>"101111111",
  40868=>"111001000",
  40869=>"010100111",
  40870=>"110111100",
  40871=>"110011010",
  40872=>"001110111",
  40873=>"000000111",
  40874=>"011111110",
  40875=>"111010100",
  40876=>"001010010",
  40877=>"000010101",
  40878=>"000010011",
  40879=>"111101100",
  40880=>"100010111",
  40881=>"110111100",
  40882=>"100100010",
  40883=>"100001011",
  40884=>"001000110",
  40885=>"101000010",
  40886=>"110100001",
  40887=>"010101101",
  40888=>"010111101",
  40889=>"110001010",
  40890=>"101001101",
  40891=>"110000101",
  40892=>"011100110",
  40893=>"110010011",
  40894=>"100000010",
  40895=>"010000011",
  40896=>"011011110",
  40897=>"001010011",
  40898=>"001000101",
  40899=>"111010111",
  40900=>"000011011",
  40901=>"010000011",
  40902=>"100001111",
  40903=>"101110111",
  40904=>"111000000",
  40905=>"000000110",
  40906=>"011101000",
  40907=>"111000101",
  40908=>"010101110",
  40909=>"000111011",
  40910=>"000111110",
  40911=>"011111011",
  40912=>"001110101",
  40913=>"010001010",
  40914=>"000110110",
  40915=>"001100101",
  40916=>"110100010",
  40917=>"000111101",
  40918=>"110100101",
  40919=>"111111101",
  40920=>"110011001",
  40921=>"010110110",
  40922=>"000111110",
  40923=>"001001110",
  40924=>"111111100",
  40925=>"010000000",
  40926=>"011100101",
  40927=>"010101001",
  40928=>"000100110",
  40929=>"100001001",
  40930=>"011001000",
  40931=>"011111000",
  40932=>"111111000",
  40933=>"000010111",
  40934=>"100101001",
  40935=>"010100111",
  40936=>"000100000",
  40937=>"110110100",
  40938=>"000010000",
  40939=>"010000100",
  40940=>"101101101",
  40941=>"010001010",
  40942=>"000000110",
  40943=>"001010011",
  40944=>"111111101",
  40945=>"100010001",
  40946=>"011101111",
  40947=>"110100100",
  40948=>"101111011",
  40949=>"000010011",
  40950=>"100011110",
  40951=>"001011100",
  40952=>"110101010",
  40953=>"101011001",
  40954=>"100101110",
  40955=>"011011110",
  40956=>"011010001",
  40957=>"010001101",
  40958=>"001000001",
  40959=>"110111100",
  40960=>"111100100",
  40961=>"010010101",
  40962=>"011010100",
  40963=>"101001111",
  40964=>"111101010",
  40965=>"011111100",
  40966=>"000111011",
  40967=>"001111011",
  40968=>"111100000",
  40969=>"100101000",
  40970=>"110111101",
  40971=>"010010111",
  40972=>"001011110",
  40973=>"010110011",
  40974=>"100010101",
  40975=>"000101111",
  40976=>"010100000",
  40977=>"000101011",
  40978=>"011110011",
  40979=>"000010110",
  40980=>"000001011",
  40981=>"010101100",
  40982=>"100010000",
  40983=>"101010110",
  40984=>"011011111",
  40985=>"101000110",
  40986=>"001000001",
  40987=>"111110110",
  40988=>"111010010",
  40989=>"011010110",
  40990=>"111111101",
  40991=>"111111000",
  40992=>"010111100",
  40993=>"000110111",
  40994=>"101111110",
  40995=>"100011001",
  40996=>"010000100",
  40997=>"111010010",
  40998=>"111001001",
  40999=>"111110101",
  41000=>"111011010",
  41001=>"100111111",
  41002=>"001111110",
  41003=>"001111101",
  41004=>"001110100",
  41005=>"110100110",
  41006=>"011011011",
  41007=>"101000111",
  41008=>"100111010",
  41009=>"000100010",
  41010=>"101111011",
  41011=>"111100100",
  41012=>"101110101",
  41013=>"011011000",
  41014=>"111001011",
  41015=>"001100111",
  41016=>"110010011",
  41017=>"010100100",
  41018=>"110101011",
  41019=>"111000001",
  41020=>"011010000",
  41021=>"100001110",
  41022=>"110011101",
  41023=>"000110010",
  41024=>"100101110",
  41025=>"001001000",
  41026=>"000101000",
  41027=>"000001110",
  41028=>"111111110",
  41029=>"001000001",
  41030=>"111000101",
  41031=>"100101010",
  41032=>"110010011",
  41033=>"000000010",
  41034=>"101010000",
  41035=>"000111101",
  41036=>"000000001",
  41037=>"110001000",
  41038=>"111100101",
  41039=>"100100001",
  41040=>"000010100",
  41041=>"101000110",
  41042=>"100100101",
  41043=>"000110110",
  41044=>"100001100",
  41045=>"111111100",
  41046=>"010101011",
  41047=>"101101101",
  41048=>"111011001",
  41049=>"110001001",
  41050=>"001000100",
  41051=>"011101110",
  41052=>"000100100",
  41053=>"100101101",
  41054=>"001100001",
  41055=>"110111110",
  41056=>"000000111",
  41057=>"101101110",
  41058=>"010100001",
  41059=>"011100000",
  41060=>"000001100",
  41061=>"011011110",
  41062=>"110100000",
  41063=>"101100000",
  41064=>"011000010",
  41065=>"100101010",
  41066=>"000011111",
  41067=>"100110000",
  41068=>"101100100",
  41069=>"100100100",
  41070=>"000001010",
  41071=>"010101101",
  41072=>"101110000",
  41073=>"001011000",
  41074=>"011100101",
  41075=>"000000011",
  41076=>"011110000",
  41077=>"010000010",
  41078=>"000001000",
  41079=>"111101011",
  41080=>"001101011",
  41081=>"011100010",
  41082=>"010001011",
  41083=>"100111000",
  41084=>"000010101",
  41085=>"011110110",
  41086=>"101001000",
  41087=>"111001000",
  41088=>"001000001",
  41089=>"011011011",
  41090=>"000010010",
  41091=>"101011101",
  41092=>"101001010",
  41093=>"010010000",
  41094=>"100001111",
  41095=>"011011000",
  41096=>"010010111",
  41097=>"000001000",
  41098=>"001010001",
  41099=>"000001111",
  41100=>"111111111",
  41101=>"101101001",
  41102=>"111100011",
  41103=>"011100111",
  41104=>"010100010",
  41105=>"000111110",
  41106=>"110111011",
  41107=>"011010100",
  41108=>"101000101",
  41109=>"111110100",
  41110=>"110011000",
  41111=>"011100110",
  41112=>"000000000",
  41113=>"110100111",
  41114=>"001001000",
  41115=>"010011001",
  41116=>"001001000",
  41117=>"010011011",
  41118=>"110001000",
  41119=>"011111110",
  41120=>"110010111",
  41121=>"011111011",
  41122=>"000001001",
  41123=>"110111000",
  41124=>"011011010",
  41125=>"010110000",
  41126=>"010100110",
  41127=>"000111110",
  41128=>"101111001",
  41129=>"011110101",
  41130=>"100000001",
  41131=>"111010000",
  41132=>"101011000",
  41133=>"010011110",
  41134=>"001000101",
  41135=>"010111110",
  41136=>"010000110",
  41137=>"001110000",
  41138=>"110100011",
  41139=>"101000001",
  41140=>"101111100",
  41141=>"111100100",
  41142=>"101111101",
  41143=>"001000011",
  41144=>"101000100",
  41145=>"110011011",
  41146=>"111000010",
  41147=>"100011101",
  41148=>"100010111",
  41149=>"010100111",
  41150=>"101110010",
  41151=>"111001111",
  41152=>"100010011",
  41153=>"101100000",
  41154=>"100011100",
  41155=>"011010101",
  41156=>"001011000",
  41157=>"000010101",
  41158=>"001001010",
  41159=>"010110000",
  41160=>"000011101",
  41161=>"010000010",
  41162=>"001111111",
  41163=>"001011010",
  41164=>"000110101",
  41165=>"000011001",
  41166=>"110101010",
  41167=>"000001110",
  41168=>"111010111",
  41169=>"101001011",
  41170=>"110001101",
  41171=>"110011110",
  41172=>"110010000",
  41173=>"100110010",
  41174=>"000101011",
  41175=>"101000110",
  41176=>"110000010",
  41177=>"100110001",
  41178=>"010111001",
  41179=>"110101110",
  41180=>"000010011",
  41181=>"110101111",
  41182=>"111000111",
  41183=>"010101101",
  41184=>"111011101",
  41185=>"110001101",
  41186=>"011111001",
  41187=>"000010100",
  41188=>"101010110",
  41189=>"010010010",
  41190=>"110100100",
  41191=>"011111011",
  41192=>"000000010",
  41193=>"011011110",
  41194=>"000011000",
  41195=>"100111101",
  41196=>"111110100",
  41197=>"010101110",
  41198=>"110001000",
  41199=>"000000111",
  41200=>"111101111",
  41201=>"000001100",
  41202=>"001111010",
  41203=>"100000101",
  41204=>"111010000",
  41205=>"001110011",
  41206=>"001010010",
  41207=>"111100001",
  41208=>"010100011",
  41209=>"000011010",
  41210=>"001101101",
  41211=>"100100100",
  41212=>"001010111",
  41213=>"011100011",
  41214=>"001100011",
  41215=>"011010011",
  41216=>"111110111",
  41217=>"110010000",
  41218=>"010100111",
  41219=>"101100010",
  41220=>"000100001",
  41221=>"101000011",
  41222=>"000001010",
  41223=>"101110111",
  41224=>"111101011",
  41225=>"010000011",
  41226=>"011111010",
  41227=>"101101111",
  41228=>"100010110",
  41229=>"000101000",
  41230=>"011000110",
  41231=>"001001000",
  41232=>"000101110",
  41233=>"101001010",
  41234=>"000010010",
  41235=>"000110001",
  41236=>"000101000",
  41237=>"010000001",
  41238=>"111111010",
  41239=>"110000111",
  41240=>"101101001",
  41241=>"010011100",
  41242=>"011001111",
  41243=>"111011011",
  41244=>"111011111",
  41245=>"111111000",
  41246=>"011110100",
  41247=>"001110000",
  41248=>"101111100",
  41249=>"111110111",
  41250=>"100000110",
  41251=>"000011010",
  41252=>"111000110",
  41253=>"110111110",
  41254=>"111100010",
  41255=>"111010001",
  41256=>"101010111",
  41257=>"101101011",
  41258=>"100001010",
  41259=>"010010010",
  41260=>"011000010",
  41261=>"000000001",
  41262=>"100010001",
  41263=>"101010011",
  41264=>"010011001",
  41265=>"101000110",
  41266=>"000110100",
  41267=>"100000100",
  41268=>"010001010",
  41269=>"011000000",
  41270=>"100000011",
  41271=>"111110101",
  41272=>"000001011",
  41273=>"001000101",
  41274=>"001111001",
  41275=>"000101110",
  41276=>"000000011",
  41277=>"111110111",
  41278=>"111011000",
  41279=>"010010111",
  41280=>"101000110",
  41281=>"100011001",
  41282=>"011011010",
  41283=>"100010000",
  41284=>"010111000",
  41285=>"011110111",
  41286=>"000111101",
  41287=>"001001110",
  41288=>"011000110",
  41289=>"110000010",
  41290=>"111101001",
  41291=>"111000000",
  41292=>"101000011",
  41293=>"010110001",
  41294=>"101111011",
  41295=>"110111001",
  41296=>"110110111",
  41297=>"110010001",
  41298=>"011010100",
  41299=>"101010111",
  41300=>"000110101",
  41301=>"000011111",
  41302=>"011011010",
  41303=>"010010110",
  41304=>"101100100",
  41305=>"101101011",
  41306=>"010101001",
  41307=>"010111101",
  41308=>"110100111",
  41309=>"000100111",
  41310=>"110100100",
  41311=>"111010011",
  41312=>"100110011",
  41313=>"111111000",
  41314=>"111000110",
  41315=>"000000000",
  41316=>"001010010",
  41317=>"000010110",
  41318=>"011011100",
  41319=>"101010101",
  41320=>"011011101",
  41321=>"011100000",
  41322=>"110110010",
  41323=>"000010000",
  41324=>"100010010",
  41325=>"100100101",
  41326=>"000001101",
  41327=>"111100011",
  41328=>"000001110",
  41329=>"110101001",
  41330=>"000101110",
  41331=>"100100010",
  41332=>"100000010",
  41333=>"010010000",
  41334=>"000011000",
  41335=>"110000110",
  41336=>"110000100",
  41337=>"011000111",
  41338=>"000100111",
  41339=>"100101101",
  41340=>"110101100",
  41341=>"100110011",
  41342=>"011011111",
  41343=>"001100000",
  41344=>"100000011",
  41345=>"010011111",
  41346=>"000111111",
  41347=>"000111111",
  41348=>"000010100",
  41349=>"000001000",
  41350=>"101101011",
  41351=>"111111010",
  41352=>"100110010",
  41353=>"100000111",
  41354=>"111001000",
  41355=>"100010110",
  41356=>"010010110",
  41357=>"110001110",
  41358=>"111101001",
  41359=>"100010110",
  41360=>"111000011",
  41361=>"000000001",
  41362=>"000000101",
  41363=>"011011100",
  41364=>"001110110",
  41365=>"010001011",
  41366=>"111110111",
  41367=>"010001010",
  41368=>"111011100",
  41369=>"100101011",
  41370=>"011010000",
  41371=>"111110101",
  41372=>"100111111",
  41373=>"111110010",
  41374=>"001011010",
  41375=>"000011001",
  41376=>"100000001",
  41377=>"001000001",
  41378=>"001100111",
  41379=>"000000000",
  41380=>"111101110",
  41381=>"101001000",
  41382=>"011001110",
  41383=>"001011111",
  41384=>"111011110",
  41385=>"100000100",
  41386=>"101110000",
  41387=>"010100000",
  41388=>"001010010",
  41389=>"111001001",
  41390=>"010011110",
  41391=>"000001010",
  41392=>"010000000",
  41393=>"011011000",
  41394=>"010100111",
  41395=>"010000111",
  41396=>"100111111",
  41397=>"001111010",
  41398=>"001011000",
  41399=>"001100011",
  41400=>"101110000",
  41401=>"101011100",
  41402=>"000000001",
  41403=>"101000001",
  41404=>"111011101",
  41405=>"000111001",
  41406=>"111101001",
  41407=>"010010101",
  41408=>"001110000",
  41409=>"101100011",
  41410=>"000110010",
  41411=>"111000101",
  41412=>"101100000",
  41413=>"000001100",
  41414=>"010001001",
  41415=>"100001000",
  41416=>"000100000",
  41417=>"000000100",
  41418=>"111110010",
  41419=>"110001101",
  41420=>"000010000",
  41421=>"101011110",
  41422=>"111011111",
  41423=>"100001001",
  41424=>"010100000",
  41425=>"101001100",
  41426=>"000000111",
  41427=>"111001110",
  41428=>"100001000",
  41429=>"100011000",
  41430=>"111000001",
  41431=>"011001100",
  41432=>"000000000",
  41433=>"110110001",
  41434=>"111110110",
  41435=>"001110001",
  41436=>"100010101",
  41437=>"110111010",
  41438=>"000110100",
  41439=>"100001111",
  41440=>"110101100",
  41441=>"110010000",
  41442=>"101010110",
  41443=>"001100000",
  41444=>"000110100",
  41445=>"001001101",
  41446=>"110001001",
  41447=>"001001010",
  41448=>"010010110",
  41449=>"000010110",
  41450=>"000000111",
  41451=>"100100000",
  41452=>"001010100",
  41453=>"111001000",
  41454=>"100011000",
  41455=>"001100110",
  41456=>"100100101",
  41457=>"111011101",
  41458=>"001110100",
  41459=>"010000001",
  41460=>"110001111",
  41461=>"001010110",
  41462=>"001110110",
  41463=>"001110001",
  41464=>"110110011",
  41465=>"110111000",
  41466=>"101010110",
  41467=>"100000111",
  41468=>"101010111",
  41469=>"100001000",
  41470=>"001001010",
  41471=>"110011010",
  41472=>"110111111",
  41473=>"100100111",
  41474=>"100111110",
  41475=>"010000000",
  41476=>"010010011",
  41477=>"110010001",
  41478=>"001100011",
  41479=>"001101110",
  41480=>"001110100",
  41481=>"110101111",
  41482=>"000010010",
  41483=>"111011001",
  41484=>"001000111",
  41485=>"000111010",
  41486=>"110100100",
  41487=>"000110100",
  41488=>"000101000",
  41489=>"000001001",
  41490=>"111101101",
  41491=>"011101110",
  41492=>"010100100",
  41493=>"111001011",
  41494=>"000110100",
  41495=>"111101000",
  41496=>"000110000",
  41497=>"001010010",
  41498=>"000100100",
  41499=>"000100010",
  41500=>"111110100",
  41501=>"011001011",
  41502=>"011111111",
  41503=>"010000000",
  41504=>"010011001",
  41505=>"101010100",
  41506=>"000101010",
  41507=>"010000000",
  41508=>"010001100",
  41509=>"100110110",
  41510=>"010001100",
  41511=>"110101000",
  41512=>"100010110",
  41513=>"111010011",
  41514=>"001001101",
  41515=>"100100000",
  41516=>"110111100",
  41517=>"010101010",
  41518=>"000100100",
  41519=>"000000001",
  41520=>"111000010",
  41521=>"000001000",
  41522=>"000101000",
  41523=>"101101101",
  41524=>"010100001",
  41525=>"110100010",
  41526=>"000101011",
  41527=>"100010110",
  41528=>"010000000",
  41529=>"100111001",
  41530=>"101100010",
  41531=>"111001010",
  41532=>"001111000",
  41533=>"110111011",
  41534=>"111100011",
  41535=>"111101011",
  41536=>"010011100",
  41537=>"001001011",
  41538=>"110001101",
  41539=>"011000010",
  41540=>"011000010",
  41541=>"101011100",
  41542=>"101000011",
  41543=>"100001010",
  41544=>"110110011",
  41545=>"101111001",
  41546=>"111001101",
  41547=>"010100110",
  41548=>"101111111",
  41549=>"111000110",
  41550=>"111000111",
  41551=>"011111000",
  41552=>"100010011",
  41553=>"010111001",
  41554=>"011101110",
  41555=>"000000100",
  41556=>"110000111",
  41557=>"100100100",
  41558=>"001011101",
  41559=>"111000010",
  41560=>"011000101",
  41561=>"000101111",
  41562=>"111101000",
  41563=>"010001000",
  41564=>"100001100",
  41565=>"100011000",
  41566=>"000000010",
  41567=>"111010001",
  41568=>"110010010",
  41569=>"111001001",
  41570=>"110010010",
  41571=>"010100011",
  41572=>"011110011",
  41573=>"000000111",
  41574=>"011010110",
  41575=>"001101101",
  41576=>"000110001",
  41577=>"110111011",
  41578=>"111111110",
  41579=>"110011111",
  41580=>"000000011",
  41581=>"011110111",
  41582=>"010000000",
  41583=>"011010110",
  41584=>"001001110",
  41585=>"001010100",
  41586=>"110010101",
  41587=>"111011011",
  41588=>"010000101",
  41589=>"011010110",
  41590=>"111110010",
  41591=>"100111010",
  41592=>"010110100",
  41593=>"010000100",
  41594=>"010000111",
  41595=>"000000101",
  41596=>"001001000",
  41597=>"000001010",
  41598=>"111100100",
  41599=>"101111110",
  41600=>"001001010",
  41601=>"011011001",
  41602=>"110111110",
  41603=>"000100001",
  41604=>"010000001",
  41605=>"001111000",
  41606=>"110000011",
  41607=>"101001001",
  41608=>"000111110",
  41609=>"000010100",
  41610=>"000111010",
  41611=>"000101001",
  41612=>"110010000",
  41613=>"101001000",
  41614=>"000011100",
  41615=>"111010110",
  41616=>"011001100",
  41617=>"110010001",
  41618=>"101010100",
  41619=>"110011001",
  41620=>"101110110",
  41621=>"001000100",
  41622=>"010011001",
  41623=>"001101101",
  41624=>"001101101",
  41625=>"100001101",
  41626=>"011110110",
  41627=>"000010101",
  41628=>"110010000",
  41629=>"011110110",
  41630=>"111100001",
  41631=>"111011101",
  41632=>"100001011",
  41633=>"100100110",
  41634=>"101111000",
  41635=>"001001001",
  41636=>"001110010",
  41637=>"110100110",
  41638=>"001001101",
  41639=>"110011110",
  41640=>"110000001",
  41641=>"100100101",
  41642=>"111100100",
  41643=>"111111110",
  41644=>"011101001",
  41645=>"010000110",
  41646=>"111100111",
  41647=>"011001001",
  41648=>"001011101",
  41649=>"101000111",
  41650=>"100010000",
  41651=>"110111100",
  41652=>"010011010",
  41653=>"010000111",
  41654=>"100000110",
  41655=>"011110010",
  41656=>"011101100",
  41657=>"011110100",
  41658=>"111000111",
  41659=>"101101101",
  41660=>"010010111",
  41661=>"111101100",
  41662=>"111111110",
  41663=>"110000011",
  41664=>"111001111",
  41665=>"110000001",
  41666=>"010010100",
  41667=>"101100000",
  41668=>"010101000",
  41669=>"001101010",
  41670=>"100101111",
  41671=>"000001100",
  41672=>"101100100",
  41673=>"110111011",
  41674=>"000000011",
  41675=>"001001000",
  41676=>"010110100",
  41677=>"010111000",
  41678=>"100111001",
  41679=>"011111100",
  41680=>"001100100",
  41681=>"110111111",
  41682=>"111110001",
  41683=>"010000111",
  41684=>"010001100",
  41685=>"000100000",
  41686=>"101001011",
  41687=>"111011000",
  41688=>"100010000",
  41689=>"100010101",
  41690=>"010001101",
  41691=>"110111010",
  41692=>"001101111",
  41693=>"111110100",
  41694=>"000010100",
  41695=>"001010000",
  41696=>"001000010",
  41697=>"100000110",
  41698=>"101000000",
  41699=>"111101000",
  41700=>"010010000",
  41701=>"011111000",
  41702=>"000100101",
  41703=>"111100010",
  41704=>"100000110",
  41705=>"100010111",
  41706=>"010000101",
  41707=>"010000111",
  41708=>"111101111",
  41709=>"000001100",
  41710=>"110000001",
  41711=>"000011110",
  41712=>"111111010",
  41713=>"000011111",
  41714=>"000110011",
  41715=>"011000011",
  41716=>"001000010",
  41717=>"110010111",
  41718=>"111110000",
  41719=>"000000011",
  41720=>"011110100",
  41721=>"010000110",
  41722=>"011110111",
  41723=>"011000010",
  41724=>"110011001",
  41725=>"111111111",
  41726=>"000000010",
  41727=>"100010000",
  41728=>"100001001",
  41729=>"110101000",
  41730=>"010110010",
  41731=>"010011101",
  41732=>"100111101",
  41733=>"000001001",
  41734=>"100110001",
  41735=>"111111101",
  41736=>"010000000",
  41737=>"001100010",
  41738=>"000010111",
  41739=>"110101100",
  41740=>"111110100",
  41741=>"010010100",
  41742=>"111110100",
  41743=>"111101100",
  41744=>"111110010",
  41745=>"000000000",
  41746=>"011110000",
  41747=>"100000100",
  41748=>"101100011",
  41749=>"111011000",
  41750=>"011100000",
  41751=>"000010011",
  41752=>"110001011",
  41753=>"110010010",
  41754=>"010011111",
  41755=>"000001110",
  41756=>"111110001",
  41757=>"101001010",
  41758=>"111000111",
  41759=>"110110011",
  41760=>"010010101",
  41761=>"100101110",
  41762=>"100010011",
  41763=>"010000000",
  41764=>"100110000",
  41765=>"110100010",
  41766=>"010101110",
  41767=>"010111101",
  41768=>"001101100",
  41769=>"000100100",
  41770=>"111101111",
  41771=>"011110110",
  41772=>"111111100",
  41773=>"000001000",
  41774=>"110011011",
  41775=>"010000011",
  41776=>"111111000",
  41777=>"101000001",
  41778=>"000101011",
  41779=>"001010000",
  41780=>"110010010",
  41781=>"101100001",
  41782=>"000100100",
  41783=>"111001000",
  41784=>"010101111",
  41785=>"111010101",
  41786=>"010010011",
  41787=>"101000000",
  41788=>"101111110",
  41789=>"011101110",
  41790=>"110111110",
  41791=>"000111011",
  41792=>"000101000",
  41793=>"110100011",
  41794=>"111111001",
  41795=>"111011100",
  41796=>"110100100",
  41797=>"001100111",
  41798=>"100111110",
  41799=>"000001110",
  41800=>"110011011",
  41801=>"111101111",
  41802=>"000111101",
  41803=>"101001011",
  41804=>"011101111",
  41805=>"000101011",
  41806=>"111011010",
  41807=>"011110011",
  41808=>"101101010",
  41809=>"001101010",
  41810=>"011111010",
  41811=>"100101110",
  41812=>"100100101",
  41813=>"000110001",
  41814=>"001001000",
  41815=>"110010000",
  41816=>"000111111",
  41817=>"100101011",
  41818=>"010111110",
  41819=>"111000110",
  41820=>"110100101",
  41821=>"000010111",
  41822=>"001110111",
  41823=>"010011000",
  41824=>"111000111",
  41825=>"111000110",
  41826=>"000111000",
  41827=>"011110000",
  41828=>"000000110",
  41829=>"000011001",
  41830=>"000100001",
  41831=>"000010001",
  41832=>"010011100",
  41833=>"010000011",
  41834=>"001010110",
  41835=>"010111001",
  41836=>"111011101",
  41837=>"110000010",
  41838=>"101101100",
  41839=>"001001111",
  41840=>"100111000",
  41841=>"000101100",
  41842=>"100100111",
  41843=>"000000100",
  41844=>"101100100",
  41845=>"011001110",
  41846=>"001100010",
  41847=>"101101111",
  41848=>"011000011",
  41849=>"010110111",
  41850=>"010111010",
  41851=>"101100010",
  41852=>"100000000",
  41853=>"000100010",
  41854=>"000001110",
  41855=>"011111110",
  41856=>"001011110",
  41857=>"111010110",
  41858=>"010010001",
  41859=>"100000011",
  41860=>"100111101",
  41861=>"111010100",
  41862=>"101000100",
  41863=>"011000000",
  41864=>"101100010",
  41865=>"101111011",
  41866=>"000000001",
  41867=>"010100011",
  41868=>"100110011",
  41869=>"011011111",
  41870=>"001000110",
  41871=>"000011011",
  41872=>"110101001",
  41873=>"010110100",
  41874=>"101101100",
  41875=>"011011001",
  41876=>"010001111",
  41877=>"111010111",
  41878=>"111110010",
  41879=>"100100100",
  41880=>"010011100",
  41881=>"100100111",
  41882=>"111111000",
  41883=>"000111111",
  41884=>"011101110",
  41885=>"000000101",
  41886=>"100110000",
  41887=>"001110011",
  41888=>"111111101",
  41889=>"111110110",
  41890=>"101110100",
  41891=>"111100110",
  41892=>"111110000",
  41893=>"111110101",
  41894=>"111011101",
  41895=>"001010000",
  41896=>"110110011",
  41897=>"001101100",
  41898=>"001000000",
  41899=>"000000101",
  41900=>"001111111",
  41901=>"001001000",
  41902=>"000010101",
  41903=>"111110001",
  41904=>"100111110",
  41905=>"111101001",
  41906=>"100100111",
  41907=>"000000110",
  41908=>"111101100",
  41909=>"011001011",
  41910=>"001000110",
  41911=>"010000000",
  41912=>"011000101",
  41913=>"111101011",
  41914=>"000011010",
  41915=>"011110000",
  41916=>"100011110",
  41917=>"111111110",
  41918=>"001111011",
  41919=>"111100011",
  41920=>"010110101",
  41921=>"011000010",
  41922=>"011000000",
  41923=>"111010111",
  41924=>"101100100",
  41925=>"100100111",
  41926=>"000011001",
  41927=>"110110000",
  41928=>"001010111",
  41929=>"010011101",
  41930=>"010000001",
  41931=>"000110110",
  41932=>"111101110",
  41933=>"100101100",
  41934=>"110001100",
  41935=>"100111101",
  41936=>"000100111",
  41937=>"110010011",
  41938=>"010000100",
  41939=>"010001111",
  41940=>"000000111",
  41941=>"110100110",
  41942=>"101111001",
  41943=>"001100011",
  41944=>"000100010",
  41945=>"000110110",
  41946=>"010100000",
  41947=>"100110111",
  41948=>"010000100",
  41949=>"111011111",
  41950=>"101001010",
  41951=>"110010000",
  41952=>"001100100",
  41953=>"100001010",
  41954=>"000111011",
  41955=>"001100010",
  41956=>"111000000",
  41957=>"000010111",
  41958=>"000010000",
  41959=>"110000000",
  41960=>"001010001",
  41961=>"101010010",
  41962=>"110110010",
  41963=>"010101010",
  41964=>"011001111",
  41965=>"100110110",
  41966=>"010111010",
  41967=>"110000100",
  41968=>"110010010",
  41969=>"101111100",
  41970=>"000100000",
  41971=>"000110110",
  41972=>"001010001",
  41973=>"111001111",
  41974=>"000100000",
  41975=>"000100111",
  41976=>"001111100",
  41977=>"010100100",
  41978=>"000101010",
  41979=>"111110110",
  41980=>"110010010",
  41981=>"000110011",
  41982=>"111100111",
  41983=>"111110011",
  41984=>"010101010",
  41985=>"100110111",
  41986=>"110101001",
  41987=>"111000111",
  41988=>"101001111",
  41989=>"110001000",
  41990=>"011100000",
  41991=>"100011101",
  41992=>"010110010",
  41993=>"001000000",
  41994=>"111010000",
  41995=>"110100001",
  41996=>"001110001",
  41997=>"110010000",
  41998=>"100100000",
  41999=>"101100001",
  42000=>"110111111",
  42001=>"001011010",
  42002=>"000111010",
  42003=>"100100111",
  42004=>"100001110",
  42005=>"110100000",
  42006=>"001000110",
  42007=>"111000101",
  42008=>"010000000",
  42009=>"000001100",
  42010=>"000011000",
  42011=>"100010001",
  42012=>"101001101",
  42013=>"100100110",
  42014=>"111101001",
  42015=>"011000000",
  42016=>"100010000",
  42017=>"110100000",
  42018=>"001001111",
  42019=>"010001010",
  42020=>"101110011",
  42021=>"011001001",
  42022=>"100001100",
  42023=>"010100000",
  42024=>"101101011",
  42025=>"010000011",
  42026=>"011011111",
  42027=>"101010100",
  42028=>"000111100",
  42029=>"011110100",
  42030=>"010010011",
  42031=>"010101111",
  42032=>"111111110",
  42033=>"011111101",
  42034=>"101110001",
  42035=>"100001001",
  42036=>"111000011",
  42037=>"000100100",
  42038=>"101110101",
  42039=>"101100000",
  42040=>"000011101",
  42041=>"101000111",
  42042=>"110100000",
  42043=>"001110001",
  42044=>"100101111",
  42045=>"100101100",
  42046=>"011100001",
  42047=>"000011110",
  42048=>"001001111",
  42049=>"011110000",
  42050=>"110001101",
  42051=>"000000111",
  42052=>"100110010",
  42053=>"000110000",
  42054=>"110011110",
  42055=>"111101111",
  42056=>"010000100",
  42057=>"100001100",
  42058=>"011010101",
  42059=>"101001101",
  42060=>"111010010",
  42061=>"001110000",
  42062=>"101011100",
  42063=>"110110011",
  42064=>"101101011",
  42065=>"111001101",
  42066=>"111111000",
  42067=>"010010101",
  42068=>"110110011",
  42069=>"011101111",
  42070=>"011101100",
  42071=>"001110001",
  42072=>"011010110",
  42073=>"100010000",
  42074=>"001010000",
  42075=>"000010111",
  42076=>"110000010",
  42077=>"011101110",
  42078=>"111111011",
  42079=>"011000011",
  42080=>"111101000",
  42081=>"111001100",
  42082=>"110111011",
  42083=>"100100111",
  42084=>"101100101",
  42085=>"000111000",
  42086=>"010100101",
  42087=>"010101011",
  42088=>"000010010",
  42089=>"111010101",
  42090=>"001101011",
  42091=>"101111111",
  42092=>"101010100",
  42093=>"011101110",
  42094=>"010000101",
  42095=>"111111111",
  42096=>"010001101",
  42097=>"101011010",
  42098=>"110110001",
  42099=>"001100111",
  42100=>"100100001",
  42101=>"101001010",
  42102=>"011011010",
  42103=>"111110100",
  42104=>"000000010",
  42105=>"111100010",
  42106=>"010101010",
  42107=>"110000101",
  42108=>"100000101",
  42109=>"010101011",
  42110=>"000100010",
  42111=>"011011111",
  42112=>"101110111",
  42113=>"111110000",
  42114=>"110001110",
  42115=>"010100010",
  42116=>"111000110",
  42117=>"101011011",
  42118=>"011010011",
  42119=>"111100010",
  42120=>"100101101",
  42121=>"000100111",
  42122=>"101110111",
  42123=>"101000110",
  42124=>"110010001",
  42125=>"001001011",
  42126=>"000001011",
  42127=>"011000001",
  42128=>"000001111",
  42129=>"111000101",
  42130=>"111110011",
  42131=>"010011100",
  42132=>"101010100",
  42133=>"000110000",
  42134=>"010001001",
  42135=>"001011101",
  42136=>"011101111",
  42137=>"010001011",
  42138=>"010011110",
  42139=>"011111101",
  42140=>"010000011",
  42141=>"110100100",
  42142=>"000011111",
  42143=>"001110010",
  42144=>"001111010",
  42145=>"001001000",
  42146=>"011110011",
  42147=>"111001111",
  42148=>"100001111",
  42149=>"001100110",
  42150=>"010101111",
  42151=>"011001000",
  42152=>"001010010",
  42153=>"110011011",
  42154=>"000001110",
  42155=>"101101111",
  42156=>"100011100",
  42157=>"111001100",
  42158=>"101010010",
  42159=>"010100010",
  42160=>"101100110",
  42161=>"110011111",
  42162=>"000100101",
  42163=>"001011010",
  42164=>"000101000",
  42165=>"000100011",
  42166=>"001111000",
  42167=>"000101101",
  42168=>"111111010",
  42169=>"011000101",
  42170=>"001111110",
  42171=>"101010010",
  42172=>"011000100",
  42173=>"000010110",
  42174=>"111001101",
  42175=>"010010111",
  42176=>"011100001",
  42177=>"001010101",
  42178=>"100001000",
  42179=>"100010101",
  42180=>"001011110",
  42181=>"010001011",
  42182=>"111101000",
  42183=>"100000111",
  42184=>"001100111",
  42185=>"011000000",
  42186=>"001100000",
  42187=>"100010101",
  42188=>"111100001",
  42189=>"011101110",
  42190=>"000110100",
  42191=>"011010101",
  42192=>"001110000",
  42193=>"010001111",
  42194=>"011001100",
  42195=>"001100101",
  42196=>"100010100",
  42197=>"110010000",
  42198=>"111011110",
  42199=>"001110001",
  42200=>"111101010",
  42201=>"010110110",
  42202=>"111011111",
  42203=>"101001001",
  42204=>"010010111",
  42205=>"101100100",
  42206=>"011001000",
  42207=>"111110000",
  42208=>"010011011",
  42209=>"000111000",
  42210=>"000100111",
  42211=>"111011110",
  42212=>"011001011",
  42213=>"001010100",
  42214=>"011111000",
  42215=>"100011110",
  42216=>"110011000",
  42217=>"001101101",
  42218=>"011000101",
  42219=>"101111001",
  42220=>"100010001",
  42221=>"111000010",
  42222=>"000001010",
  42223=>"111111111",
  42224=>"111111101",
  42225=>"001010110",
  42226=>"111011000",
  42227=>"100000100",
  42228=>"100010010",
  42229=>"010011011",
  42230=>"101110011",
  42231=>"000000111",
  42232=>"011010000",
  42233=>"001101111",
  42234=>"110110100",
  42235=>"100101001",
  42236=>"101110100",
  42237=>"011000000",
  42238=>"111011011",
  42239=>"000110101",
  42240=>"110110101",
  42241=>"111001100",
  42242=>"101011011",
  42243=>"101100100",
  42244=>"110111001",
  42245=>"010011110",
  42246=>"100100011",
  42247=>"011011001",
  42248=>"010010010",
  42249=>"010110111",
  42250=>"000110111",
  42251=>"100100000",
  42252=>"101001001",
  42253=>"110001100",
  42254=>"100000101",
  42255=>"111111110",
  42256=>"100110110",
  42257=>"011001111",
  42258=>"011100101",
  42259=>"011011001",
  42260=>"011110000",
  42261=>"010100011",
  42262=>"001001010",
  42263=>"000110010",
  42264=>"000010010",
  42265=>"110101010",
  42266=>"000001100",
  42267=>"110101111",
  42268=>"110100011",
  42269=>"011111111",
  42270=>"111100000",
  42271=>"001000101",
  42272=>"101000101",
  42273=>"101010001",
  42274=>"110111101",
  42275=>"111010001",
  42276=>"000010101",
  42277=>"000011001",
  42278=>"011111100",
  42279=>"011100100",
  42280=>"100010111",
  42281=>"000100100",
  42282=>"001001001",
  42283=>"011011111",
  42284=>"100100001",
  42285=>"000111001",
  42286=>"101100010",
  42287=>"101011101",
  42288=>"000010000",
  42289=>"110000101",
  42290=>"000101100",
  42291=>"101000001",
  42292=>"110111001",
  42293=>"101000100",
  42294=>"011001110",
  42295=>"110100101",
  42296=>"100110001",
  42297=>"011111000",
  42298=>"011011111",
  42299=>"110111110",
  42300=>"110001001",
  42301=>"111101100",
  42302=>"001010011",
  42303=>"111111001",
  42304=>"100000000",
  42305=>"110001100",
  42306=>"010011001",
  42307=>"111000110",
  42308=>"110100110",
  42309=>"111001110",
  42310=>"111010101",
  42311=>"110010011",
  42312=>"000101011",
  42313=>"000011101",
  42314=>"101001100",
  42315=>"111000110",
  42316=>"011111011",
  42317=>"000100110",
  42318=>"000110100",
  42319=>"110111110",
  42320=>"101101000",
  42321=>"111111000",
  42322=>"110011011",
  42323=>"101011101",
  42324=>"100111011",
  42325=>"100010111",
  42326=>"100001001",
  42327=>"110110110",
  42328=>"111011101",
  42329=>"111000110",
  42330=>"011111010",
  42331=>"001010000",
  42332=>"000101100",
  42333=>"100101000",
  42334=>"111110000",
  42335=>"100101000",
  42336=>"001011010",
  42337=>"001100101",
  42338=>"110100001",
  42339=>"110110001",
  42340=>"001011111",
  42341=>"100101110",
  42342=>"010110111",
  42343=>"001100100",
  42344=>"001010000",
  42345=>"000000100",
  42346=>"111000010",
  42347=>"111111110",
  42348=>"111101101",
  42349=>"100010100",
  42350=>"100001111",
  42351=>"001101010",
  42352=>"000001000",
  42353=>"001010100",
  42354=>"111000011",
  42355=>"111111110",
  42356=>"000101010",
  42357=>"000000010",
  42358=>"100010011",
  42359=>"011001010",
  42360=>"111100000",
  42361=>"010100111",
  42362=>"001001101",
  42363=>"110101110",
  42364=>"100010001",
  42365=>"010010100",
  42366=>"011001001",
  42367=>"011011110",
  42368=>"100010011",
  42369=>"111001100",
  42370=>"110110000",
  42371=>"011000111",
  42372=>"100110100",
  42373=>"011100000",
  42374=>"000010000",
  42375=>"100010110",
  42376=>"100000011",
  42377=>"001000110",
  42378=>"101111111",
  42379=>"101000100",
  42380=>"100000011",
  42381=>"111001111",
  42382=>"101000010",
  42383=>"101110011",
  42384=>"010001101",
  42385=>"101110001",
  42386=>"110101101",
  42387=>"101001011",
  42388=>"100101010",
  42389=>"100001110",
  42390=>"000000011",
  42391=>"010011111",
  42392=>"001111100",
  42393=>"110011101",
  42394=>"110010110",
  42395=>"001001001",
  42396=>"111001110",
  42397=>"000100010",
  42398=>"110011100",
  42399=>"101101111",
  42400=>"011011110",
  42401=>"001101101",
  42402=>"001001100",
  42403=>"100100000",
  42404=>"001000110",
  42405=>"110101011",
  42406=>"110110101",
  42407=>"010010011",
  42408=>"011111001",
  42409=>"111010001",
  42410=>"101100111",
  42411=>"101100010",
  42412=>"100110010",
  42413=>"100001110",
  42414=>"010000101",
  42415=>"011111110",
  42416=>"111100001",
  42417=>"001010011",
  42418=>"001011100",
  42419=>"001101001",
  42420=>"111011001",
  42421=>"010101100",
  42422=>"001110100",
  42423=>"110110101",
  42424=>"101000100",
  42425=>"001110111",
  42426=>"010100010",
  42427=>"110000111",
  42428=>"000111101",
  42429=>"101011011",
  42430=>"001000101",
  42431=>"000110001",
  42432=>"010110011",
  42433=>"110000001",
  42434=>"011011111",
  42435=>"110101111",
  42436=>"101010101",
  42437=>"011011100",
  42438=>"111011001",
  42439=>"011101011",
  42440=>"110001001",
  42441=>"101011010",
  42442=>"000001110",
  42443=>"100011100",
  42444=>"011111110",
  42445=>"010010110",
  42446=>"110100010",
  42447=>"000001100",
  42448=>"010100110",
  42449=>"101011011",
  42450=>"111111001",
  42451=>"010000100",
  42452=>"101111111",
  42453=>"101011111",
  42454=>"011010000",
  42455=>"011101011",
  42456=>"000010100",
  42457=>"011100001",
  42458=>"111000111",
  42459=>"110000101",
  42460=>"011000111",
  42461=>"101110111",
  42462=>"010110101",
  42463=>"011011111",
  42464=>"011001101",
  42465=>"011111010",
  42466=>"010100100",
  42467=>"001011111",
  42468=>"111110010",
  42469=>"101101001",
  42470=>"010010000",
  42471=>"101110000",
  42472=>"110000101",
  42473=>"001111001",
  42474=>"000001001",
  42475=>"110011010",
  42476=>"100111001",
  42477=>"100010001",
  42478=>"101100101",
  42479=>"110101010",
  42480=>"000001111",
  42481=>"111010100",
  42482=>"010011101",
  42483=>"001000100",
  42484=>"011000110",
  42485=>"110110001",
  42486=>"110110111",
  42487=>"000110111",
  42488=>"000001101",
  42489=>"111100100",
  42490=>"011100000",
  42491=>"110011111",
  42492=>"101100011",
  42493=>"111010011",
  42494=>"001110010",
  42495=>"101000011",
  42496=>"101000000",
  42497=>"111011011",
  42498=>"011010001",
  42499=>"100011111",
  42500=>"110111001",
  42501=>"000010111",
  42502=>"111110111",
  42503=>"101011110",
  42504=>"000011110",
  42505=>"110100111",
  42506=>"010100110",
  42507=>"001111111",
  42508=>"111111010",
  42509=>"000001001",
  42510=>"110000111",
  42511=>"101010111",
  42512=>"100101111",
  42513=>"010010010",
  42514=>"011010000",
  42515=>"010010101",
  42516=>"000000100",
  42517=>"101011100",
  42518=>"000010001",
  42519=>"100111000",
  42520=>"100111111",
  42521=>"011100100",
  42522=>"100111010",
  42523=>"011001001",
  42524=>"011101111",
  42525=>"100100000",
  42526=>"101011010",
  42527=>"000010000",
  42528=>"101010110",
  42529=>"111011101",
  42530=>"000111001",
  42531=>"001111001",
  42532=>"001101000",
  42533=>"001110010",
  42534=>"010100010",
  42535=>"001000100",
  42536=>"000100010",
  42537=>"011001011",
  42538=>"101111110",
  42539=>"110100111",
  42540=>"011010101",
  42541=>"100010011",
  42542=>"111001010",
  42543=>"011001000",
  42544=>"000111101",
  42545=>"101001000",
  42546=>"111001001",
  42547=>"110010000",
  42548=>"010011010",
  42549=>"000010010",
  42550=>"000011011",
  42551=>"111111010",
  42552=>"100010101",
  42553=>"111110011",
  42554=>"001110101",
  42555=>"101100101",
  42556=>"011010010",
  42557=>"011101110",
  42558=>"101100100",
  42559=>"101001000",
  42560=>"100100000",
  42561=>"011110010",
  42562=>"100111001",
  42563=>"100011011",
  42564=>"011111010",
  42565=>"111100001",
  42566=>"010100010",
  42567=>"110000110",
  42568=>"001111110",
  42569=>"100101000",
  42570=>"100100010",
  42571=>"000010000",
  42572=>"110110001",
  42573=>"010101100",
  42574=>"011111101",
  42575=>"001101000",
  42576=>"000110001",
  42577=>"010110001",
  42578=>"011011000",
  42579=>"000010110",
  42580=>"011010011",
  42581=>"111010000",
  42582=>"010011001",
  42583=>"101110110",
  42584=>"000100100",
  42585=>"101000000",
  42586=>"010011110",
  42587=>"101001101",
  42588=>"001010011",
  42589=>"100010011",
  42590=>"111101000",
  42591=>"101001011",
  42592=>"111010100",
  42593=>"101100001",
  42594=>"010000111",
  42595=>"110100111",
  42596=>"101110111",
  42597=>"001101111",
  42598=>"001101111",
  42599=>"100100100",
  42600=>"100000010",
  42601=>"011010001",
  42602=>"101101110",
  42603=>"000101110",
  42604=>"111000010",
  42605=>"000111001",
  42606=>"001110001",
  42607=>"110011110",
  42608=>"011001101",
  42609=>"110111000",
  42610=>"000100101",
  42611=>"100110010",
  42612=>"000001011",
  42613=>"011000110",
  42614=>"011101110",
  42615=>"101111111",
  42616=>"100100110",
  42617=>"100001100",
  42618=>"111110101",
  42619=>"001011111",
  42620=>"101001001",
  42621=>"011001000",
  42622=>"100101010",
  42623=>"000000100",
  42624=>"011100101",
  42625=>"110110001",
  42626=>"000010010",
  42627=>"000100100",
  42628=>"011001000",
  42629=>"001010110",
  42630=>"111000110",
  42631=>"011011011",
  42632=>"111011001",
  42633=>"000010000",
  42634=>"011010001",
  42635=>"110010111",
  42636=>"100000110",
  42637=>"001001100",
  42638=>"101110111",
  42639=>"011010000",
  42640=>"101001100",
  42641=>"000101110",
  42642=>"110110011",
  42643=>"100100100",
  42644=>"100111011",
  42645=>"100101111",
  42646=>"010110110",
  42647=>"001010101",
  42648=>"011100000",
  42649=>"100000001",
  42650=>"000101000",
  42651=>"001000001",
  42652=>"000000110",
  42653=>"100101011",
  42654=>"100010101",
  42655=>"100001011",
  42656=>"001100000",
  42657=>"010100100",
  42658=>"000110101",
  42659=>"000011011",
  42660=>"000001110",
  42661=>"011010000",
  42662=>"000101111",
  42663=>"000010001",
  42664=>"011000000",
  42665=>"000010101",
  42666=>"000100010",
  42667=>"100000111",
  42668=>"011010101",
  42669=>"010101000",
  42670=>"001111000",
  42671=>"101000010",
  42672=>"011001100",
  42673=>"000011000",
  42674=>"011011001",
  42675=>"111100100",
  42676=>"110111110",
  42677=>"011101101",
  42678=>"000011111",
  42679=>"111001110",
  42680=>"011101011",
  42681=>"010111101",
  42682=>"010001010",
  42683=>"001110100",
  42684=>"000011101",
  42685=>"011000001",
  42686=>"111001010",
  42687=>"111010001",
  42688=>"000001110",
  42689=>"010101010",
  42690=>"010111011",
  42691=>"100000111",
  42692=>"000111000",
  42693=>"011101111",
  42694=>"100110110",
  42695=>"111000001",
  42696=>"000110010",
  42697=>"011100110",
  42698=>"000010111",
  42699=>"100000111",
  42700=>"111111100",
  42701=>"000010110",
  42702=>"000100110",
  42703=>"001001011",
  42704=>"110111011",
  42705=>"110111100",
  42706=>"111010000",
  42707=>"001101001",
  42708=>"101110001",
  42709=>"010011111",
  42710=>"101100100",
  42711=>"101011110",
  42712=>"010010110",
  42713=>"010010111",
  42714=>"000011001",
  42715=>"100000100",
  42716=>"010001000",
  42717=>"001100011",
  42718=>"110010111",
  42719=>"011010010",
  42720=>"101001001",
  42721=>"001010110",
  42722=>"110101001",
  42723=>"011111011",
  42724=>"101000100",
  42725=>"001101110",
  42726=>"101110001",
  42727=>"101111000",
  42728=>"101111000",
  42729=>"101000110",
  42730=>"110101010",
  42731=>"001011000",
  42732=>"101001001",
  42733=>"010110100",
  42734=>"011111001",
  42735=>"001111011",
  42736=>"000001110",
  42737=>"111001100",
  42738=>"110011010",
  42739=>"001101110",
  42740=>"110010010",
  42741=>"011110100",
  42742=>"001100000",
  42743=>"000011000",
  42744=>"101011100",
  42745=>"000110000",
  42746=>"111001010",
  42747=>"000111110",
  42748=>"010010000",
  42749=>"010100100",
  42750=>"011111001",
  42751=>"011010100",
  42752=>"000010111",
  42753=>"100000100",
  42754=>"100110000",
  42755=>"110101000",
  42756=>"001000000",
  42757=>"100101010",
  42758=>"100000010",
  42759=>"111001110",
  42760=>"100011000",
  42761=>"111100000",
  42762=>"110110110",
  42763=>"000100011",
  42764=>"010000000",
  42765=>"111111010",
  42766=>"000111110",
  42767=>"111111010",
  42768=>"011101100",
  42769=>"001111110",
  42770=>"001001000",
  42771=>"100000111",
  42772=>"100111001",
  42773=>"010111011",
  42774=>"111010110",
  42775=>"010001001",
  42776=>"001000000",
  42777=>"100100110",
  42778=>"001100011",
  42779=>"011110011",
  42780=>"000001111",
  42781=>"001010111",
  42782=>"010101111",
  42783=>"100101110",
  42784=>"001001001",
  42785=>"011010110",
  42786=>"000000011",
  42787=>"010001000",
  42788=>"001110001",
  42789=>"111101001",
  42790=>"001011111",
  42791=>"110111111",
  42792=>"110100101",
  42793=>"000110101",
  42794=>"010100110",
  42795=>"110010101",
  42796=>"011100000",
  42797=>"110011101",
  42798=>"001010011",
  42799=>"110010110",
  42800=>"010001011",
  42801=>"010010110",
  42802=>"000001001",
  42803=>"010100100",
  42804=>"110011000",
  42805=>"110101101",
  42806=>"111001011",
  42807=>"000111101",
  42808=>"000010100",
  42809=>"001110010",
  42810=>"001000000",
  42811=>"010001010",
  42812=>"010010100",
  42813=>"001001000",
  42814=>"010010111",
  42815=>"111010001",
  42816=>"000100001",
  42817=>"110111010",
  42818=>"001111011",
  42819=>"011001111",
  42820=>"000010010",
  42821=>"111111111",
  42822=>"101010001",
  42823=>"011100000",
  42824=>"001000000",
  42825=>"100110001",
  42826=>"101001001",
  42827=>"010000011",
  42828=>"111011111",
  42829=>"111000010",
  42830=>"011110001",
  42831=>"110010100",
  42832=>"101000111",
  42833=>"100001001",
  42834=>"100010101",
  42835=>"011001011",
  42836=>"000001010",
  42837=>"000111111",
  42838=>"111111100",
  42839=>"011100001",
  42840=>"010010110",
  42841=>"110111001",
  42842=>"111101101",
  42843=>"110010101",
  42844=>"001000011",
  42845=>"010110110",
  42846=>"000101001",
  42847=>"000011111",
  42848=>"000110100",
  42849=>"001000000",
  42850=>"000101100",
  42851=>"000101000",
  42852=>"001001000",
  42853=>"010101010",
  42854=>"011010010",
  42855=>"011001101",
  42856=>"110100010",
  42857=>"000001111",
  42858=>"101000100",
  42859=>"111100100",
  42860=>"010111110",
  42861=>"111101010",
  42862=>"101001011",
  42863=>"110111010",
  42864=>"010011100",
  42865=>"110011101",
  42866=>"000011011",
  42867=>"000001101",
  42868=>"000110111",
  42869=>"011001000",
  42870=>"110010000",
  42871=>"110100010",
  42872=>"010101100",
  42873=>"100000011",
  42874=>"111111011",
  42875=>"101001001",
  42876=>"010000011",
  42877=>"001111110",
  42878=>"000000100",
  42879=>"011001110",
  42880=>"011100011",
  42881=>"101011010",
  42882=>"011101001",
  42883=>"111111111",
  42884=>"101110110",
  42885=>"001101011",
  42886=>"010010100",
  42887=>"101100000",
  42888=>"110110100",
  42889=>"010010011",
  42890=>"110111100",
  42891=>"111100111",
  42892=>"011101100",
  42893=>"111100111",
  42894=>"101101001",
  42895=>"000100110",
  42896=>"000000010",
  42897=>"110001000",
  42898=>"100010101",
  42899=>"001010110",
  42900=>"000111101",
  42901=>"101100011",
  42902=>"000101010",
  42903=>"000110110",
  42904=>"010001001",
  42905=>"001011001",
  42906=>"100011011",
  42907=>"101010111",
  42908=>"001010111",
  42909=>"101010100",
  42910=>"001010101",
  42911=>"001111110",
  42912=>"010000010",
  42913=>"100110010",
  42914=>"111010001",
  42915=>"111111111",
  42916=>"100110000",
  42917=>"011100111",
  42918=>"010010001",
  42919=>"010010100",
  42920=>"101100101",
  42921=>"011000000",
  42922=>"000111001",
  42923=>"101100000",
  42924=>"101100001",
  42925=>"101110110",
  42926=>"100011011",
  42927=>"100000111",
  42928=>"001100110",
  42929=>"111110111",
  42930=>"001010110",
  42931=>"010110000",
  42932=>"110101100",
  42933=>"111101111",
  42934=>"111110100",
  42935=>"000000110",
  42936=>"001001000",
  42937=>"011000111",
  42938=>"010011001",
  42939=>"110001110",
  42940=>"111101000",
  42941=>"100101100",
  42942=>"011111001",
  42943=>"000010100",
  42944=>"111101100",
  42945=>"111001110",
  42946=>"001101111",
  42947=>"001001100",
  42948=>"110100100",
  42949=>"000111001",
  42950=>"001101110",
  42951=>"010000100",
  42952=>"000000110",
  42953=>"000001100",
  42954=>"111100111",
  42955=>"110011001",
  42956=>"111001000",
  42957=>"010000101",
  42958=>"011100010",
  42959=>"101100101",
  42960=>"011011111",
  42961=>"001011110",
  42962=>"011101001",
  42963=>"111000110",
  42964=>"011010001",
  42965=>"001001100",
  42966=>"111100100",
  42967=>"000011101",
  42968=>"011001110",
  42969=>"111100001",
  42970=>"111010011",
  42971=>"011100000",
  42972=>"100001100",
  42973=>"010101001",
  42974=>"100100000",
  42975=>"110010010",
  42976=>"010011100",
  42977=>"010101010",
  42978=>"000000111",
  42979=>"011010000",
  42980=>"010000101",
  42981=>"101010100",
  42982=>"011101101",
  42983=>"010001110",
  42984=>"100111000",
  42985=>"000100100",
  42986=>"110010110",
  42987=>"000000110",
  42988=>"001111001",
  42989=>"101100010",
  42990=>"100011001",
  42991=>"111110001",
  42992=>"110101011",
  42993=>"100010011",
  42994=>"110111010",
  42995=>"011010010",
  42996=>"110110010",
  42997=>"001011001",
  42998=>"010101001",
  42999=>"010100000",
  43000=>"100110110",
  43001=>"100010000",
  43002=>"000101000",
  43003=>"100110101",
  43004=>"111100011",
  43005=>"010111111",
  43006=>"001110101",
  43007=>"010010011",
  43008=>"010000011",
  43009=>"111111101",
  43010=>"111001011",
  43011=>"010000000",
  43012=>"100110010",
  43013=>"001111001",
  43014=>"010101100",
  43015=>"100010100",
  43016=>"111110001",
  43017=>"110111001",
  43018=>"010001011",
  43019=>"010101100",
  43020=>"110011001",
  43021=>"010011110",
  43022=>"011001001",
  43023=>"111000011",
  43024=>"000001010",
  43025=>"000001110",
  43026=>"010010010",
  43027=>"100001100",
  43028=>"011111110",
  43029=>"011101101",
  43030=>"110000111",
  43031=>"000001111",
  43032=>"100010100",
  43033=>"101001110",
  43034=>"100111110",
  43035=>"010111011",
  43036=>"010100011",
  43037=>"101100111",
  43038=>"111001001",
  43039=>"000110101",
  43040=>"010011011",
  43041=>"101001001",
  43042=>"011100100",
  43043=>"001111100",
  43044=>"010101111",
  43045=>"011010111",
  43046=>"000000000",
  43047=>"111100011",
  43048=>"100010011",
  43049=>"010010001",
  43050=>"101111111",
  43051=>"111010011",
  43052=>"101001101",
  43053=>"111101011",
  43054=>"110100111",
  43055=>"101111001",
  43056=>"000110110",
  43057=>"110001111",
  43058=>"000110000",
  43059=>"110110010",
  43060=>"011000110",
  43061=>"011110001",
  43062=>"100100010",
  43063=>"001000001",
  43064=>"011000011",
  43065=>"100101001",
  43066=>"001001000",
  43067=>"011010010",
  43068=>"100010101",
  43069=>"001011101",
  43070=>"101101001",
  43071=>"011110000",
  43072=>"110001001",
  43073=>"000000000",
  43074=>"100110111",
  43075=>"000001100",
  43076=>"110011001",
  43077=>"101100110",
  43078=>"111110100",
  43079=>"111111101",
  43080=>"100110010",
  43081=>"010010000",
  43082=>"100101111",
  43083=>"010010000",
  43084=>"111110000",
  43085=>"111101000",
  43086=>"011001001",
  43087=>"101110010",
  43088=>"111000101",
  43089=>"100101111",
  43090=>"000010001",
  43091=>"000100001",
  43092=>"101111110",
  43093=>"001000000",
  43094=>"101011100",
  43095=>"100101111",
  43096=>"100111101",
  43097=>"111100011",
  43098=>"001111001",
  43099=>"111001101",
  43100=>"001100000",
  43101=>"110001011",
  43102=>"111110110",
  43103=>"010001110",
  43104=>"000100000",
  43105=>"111011101",
  43106=>"000110000",
  43107=>"000011111",
  43108=>"111000100",
  43109=>"001011010",
  43110=>"101001001",
  43111=>"100001100",
  43112=>"001111111",
  43113=>"000000100",
  43114=>"001000100",
  43115=>"101101111",
  43116=>"010100001",
  43117=>"001000010",
  43118=>"101011010",
  43119=>"001101110",
  43120=>"010101100",
  43121=>"111011101",
  43122=>"000001000",
  43123=>"000010111",
  43124=>"000000001",
  43125=>"110100110",
  43126=>"100001011",
  43127=>"000100110",
  43128=>"011011000",
  43129=>"001110000",
  43130=>"101101011",
  43131=>"110100101",
  43132=>"101110101",
  43133=>"101101110",
  43134=>"110101101",
  43135=>"000110001",
  43136=>"111010111",
  43137=>"100111100",
  43138=>"101101110",
  43139=>"101101110",
  43140=>"101000111",
  43141=>"101001110",
  43142=>"011110001",
  43143=>"010010000",
  43144=>"110011111",
  43145=>"001000001",
  43146=>"110011000",
  43147=>"000010001",
  43148=>"100111000",
  43149=>"110101110",
  43150=>"100111011",
  43151=>"100101010",
  43152=>"101100011",
  43153=>"010101000",
  43154=>"010001011",
  43155=>"101111011",
  43156=>"111100010",
  43157=>"100100011",
  43158=>"110111110",
  43159=>"010010000",
  43160=>"110110001",
  43161=>"001101011",
  43162=>"101010010",
  43163=>"000010001",
  43164=>"100111101",
  43165=>"001100001",
  43166=>"001001110",
  43167=>"101110011",
  43168=>"100100001",
  43169=>"111010101",
  43170=>"010111001",
  43171=>"100001010",
  43172=>"000101101",
  43173=>"001111111",
  43174=>"101011100",
  43175=>"111111110",
  43176=>"110010000",
  43177=>"111011100",
  43178=>"101111100",
  43179=>"101000011",
  43180=>"010111010",
  43181=>"011011100",
  43182=>"001000100",
  43183=>"000111100",
  43184=>"110010000",
  43185=>"101000010",
  43186=>"000001100",
  43187=>"001111001",
  43188=>"100100111",
  43189=>"100111001",
  43190=>"111011011",
  43191=>"101100010",
  43192=>"000001000",
  43193=>"001011001",
  43194=>"101100010",
  43195=>"110101010",
  43196=>"100000110",
  43197=>"011011001",
  43198=>"011101110",
  43199=>"111110000",
  43200=>"110001110",
  43201=>"110100010",
  43202=>"010001001",
  43203=>"100001001",
  43204=>"101010100",
  43205=>"111001011",
  43206=>"000000000",
  43207=>"111100011",
  43208=>"010111110",
  43209=>"011001001",
  43210=>"101010010",
  43211=>"011110001",
  43212=>"001000010",
  43213=>"111111111",
  43214=>"110000101",
  43215=>"000010111",
  43216=>"010111000",
  43217=>"110000000",
  43218=>"000001010",
  43219=>"101100111",
  43220=>"111000011",
  43221=>"010100010",
  43222=>"101001100",
  43223=>"101111110",
  43224=>"101001000",
  43225=>"001001110",
  43226=>"101101111",
  43227=>"100101110",
  43228=>"101100111",
  43229=>"110110010",
  43230=>"001110111",
  43231=>"010011000",
  43232=>"001101110",
  43233=>"001010010",
  43234=>"010100011",
  43235=>"100110101",
  43236=>"001001000",
  43237=>"011001101",
  43238=>"001100010",
  43239=>"001011100",
  43240=>"101100110",
  43241=>"111010110",
  43242=>"010000110",
  43243=>"110000101",
  43244=>"010101111",
  43245=>"100010011",
  43246=>"110111111",
  43247=>"010101010",
  43248=>"101000001",
  43249=>"110001000",
  43250=>"100110110",
  43251=>"001000111",
  43252=>"011101010",
  43253=>"100011000",
  43254=>"111101110",
  43255=>"101011000",
  43256=>"001000110",
  43257=>"011000011",
  43258=>"000001010",
  43259=>"010001001",
  43260=>"110101011",
  43261=>"000000010",
  43262=>"110111101",
  43263=>"000001010",
  43264=>"101110100",
  43265=>"110000011",
  43266=>"111110000",
  43267=>"011110001",
  43268=>"010101000",
  43269=>"001101100",
  43270=>"000001010",
  43271=>"010000011",
  43272=>"001000000",
  43273=>"111000101",
  43274=>"100111001",
  43275=>"111011111",
  43276=>"110010110",
  43277=>"100011011",
  43278=>"001100001",
  43279=>"110100010",
  43280=>"111100010",
  43281=>"000100101",
  43282=>"101101110",
  43283=>"011001010",
  43284=>"001000111",
  43285=>"111100010",
  43286=>"110111101",
  43287=>"101011010",
  43288=>"001000011",
  43289=>"010100100",
  43290=>"011000001",
  43291=>"101000110",
  43292=>"000101010",
  43293=>"110000010",
  43294=>"011111001",
  43295=>"110111010",
  43296=>"110010101",
  43297=>"100101100",
  43298=>"111110000",
  43299=>"000000111",
  43300=>"000010010",
  43301=>"101010011",
  43302=>"100100101",
  43303=>"000011001",
  43304=>"001101001",
  43305=>"101101110",
  43306=>"011110010",
  43307=>"100000111",
  43308=>"100101011",
  43309=>"000000100",
  43310=>"000010010",
  43311=>"110101111",
  43312=>"010011111",
  43313=>"010110100",
  43314=>"111011101",
  43315=>"000010111",
  43316=>"011001001",
  43317=>"001111000",
  43318=>"000110010",
  43319=>"011001110",
  43320=>"110001110",
  43321=>"011011100",
  43322=>"111110111",
  43323=>"111101000",
  43324=>"100001010",
  43325=>"001100000",
  43326=>"000100100",
  43327=>"001001010",
  43328=>"000101000",
  43329=>"001111101",
  43330=>"111010101",
  43331=>"100010101",
  43332=>"011011101",
  43333=>"101100100",
  43334=>"100010101",
  43335=>"110111001",
  43336=>"000110010",
  43337=>"100101010",
  43338=>"101100110",
  43339=>"010011001",
  43340=>"010101001",
  43341=>"111101001",
  43342=>"111110010",
  43343=>"111110011",
  43344=>"100101010",
  43345=>"000100001",
  43346=>"100101001",
  43347=>"100110111",
  43348=>"111111010",
  43349=>"100101010",
  43350=>"000100010",
  43351=>"010011111",
  43352=>"011111101",
  43353=>"111010110",
  43354=>"010000001",
  43355=>"010001011",
  43356=>"110101110",
  43357=>"101011100",
  43358=>"101001111",
  43359=>"010111010",
  43360=>"111010010",
  43361=>"100011110",
  43362=>"001101001",
  43363=>"100000111",
  43364=>"111111110",
  43365=>"000000001",
  43366=>"100111100",
  43367=>"111000100",
  43368=>"000100111",
  43369=>"011011011",
  43370=>"001001101",
  43371=>"101111101",
  43372=>"010101000",
  43373=>"011110010",
  43374=>"011001110",
  43375=>"110010101",
  43376=>"010001010",
  43377=>"100111111",
  43378=>"001110000",
  43379=>"111001011",
  43380=>"101010111",
  43381=>"000001111",
  43382=>"011001101",
  43383=>"010010111",
  43384=>"000101011",
  43385=>"011011100",
  43386=>"111000111",
  43387=>"000000000",
  43388=>"011100100",
  43389=>"000010100",
  43390=>"000101000",
  43391=>"110110111",
  43392=>"001110000",
  43393=>"001101011",
  43394=>"110111000",
  43395=>"110010011",
  43396=>"011101000",
  43397=>"101111111",
  43398=>"111001011",
  43399=>"000010011",
  43400=>"001000001",
  43401=>"001110111",
  43402=>"101011111",
  43403=>"001101100",
  43404=>"111010000",
  43405=>"100010011",
  43406=>"111001110",
  43407=>"001110110",
  43408=>"001010101",
  43409=>"100101111",
  43410=>"100110000",
  43411=>"100000111",
  43412=>"100101101",
  43413=>"011100001",
  43414=>"100011011",
  43415=>"010000001",
  43416=>"001101101",
  43417=>"101101001",
  43418=>"100111100",
  43419=>"001011010",
  43420=>"100101001",
  43421=>"101000011",
  43422=>"011100010",
  43423=>"101110101",
  43424=>"010000001",
  43425=>"011101100",
  43426=>"011001001",
  43427=>"110000011",
  43428=>"010001101",
  43429=>"011101000",
  43430=>"111010001",
  43431=>"111111111",
  43432=>"111101011",
  43433=>"000010111",
  43434=>"111110001",
  43435=>"100000000",
  43436=>"001011111",
  43437=>"010110001",
  43438=>"100010011",
  43439=>"001010101",
  43440=>"111010011",
  43441=>"000010010",
  43442=>"100010000",
  43443=>"110111111",
  43444=>"100111111",
  43445=>"000111010",
  43446=>"101111000",
  43447=>"000100000",
  43448=>"111111100",
  43449=>"001111010",
  43450=>"001000101",
  43451=>"001101010",
  43452=>"001111000",
  43453=>"100000111",
  43454=>"101110000",
  43455=>"111110011",
  43456=>"111001110",
  43457=>"001100110",
  43458=>"110010110",
  43459=>"011010101",
  43460=>"110110111",
  43461=>"100100101",
  43462=>"101101101",
  43463=>"100010100",
  43464=>"011100100",
  43465=>"110100001",
  43466=>"100001110",
  43467=>"100111101",
  43468=>"100111000",
  43469=>"110000101",
  43470=>"000011010",
  43471=>"001001001",
  43472=>"100111100",
  43473=>"111001101",
  43474=>"000011010",
  43475=>"000110010",
  43476=>"110100111",
  43477=>"101110111",
  43478=>"011001111",
  43479=>"000110110",
  43480=>"001101000",
  43481=>"100010000",
  43482=>"011100011",
  43483=>"001111100",
  43484=>"000011100",
  43485=>"110110100",
  43486=>"111110001",
  43487=>"110010100",
  43488=>"001010101",
  43489=>"100011110",
  43490=>"001100110",
  43491=>"011011100",
  43492=>"010000010",
  43493=>"111010110",
  43494=>"110001101",
  43495=>"000100101",
  43496=>"000001001",
  43497=>"010111010",
  43498=>"000010011",
  43499=>"011100011",
  43500=>"001111011",
  43501=>"011001001",
  43502=>"101010000",
  43503=>"110111110",
  43504=>"011111111",
  43505=>"001001110",
  43506=>"001011110",
  43507=>"101000110",
  43508=>"011100101",
  43509=>"000100100",
  43510=>"011111110",
  43511=>"111110111",
  43512=>"111001100",
  43513=>"110100111",
  43514=>"000000001",
  43515=>"010110001",
  43516=>"011001111",
  43517=>"101111000",
  43518=>"000001101",
  43519=>"001100101",
  43520=>"111100011",
  43521=>"000001011",
  43522=>"000010000",
  43523=>"000110011",
  43524=>"101001111",
  43525=>"000101110",
  43526=>"001001111",
  43527=>"001111010",
  43528=>"101111000",
  43529=>"000111001",
  43530=>"010000111",
  43531=>"011110010",
  43532=>"011100110",
  43533=>"010000000",
  43534=>"001111000",
  43535=>"110000011",
  43536=>"010100100",
  43537=>"101100100",
  43538=>"111000110",
  43539=>"100010011",
  43540=>"001110011",
  43541=>"111000111",
  43542=>"000100101",
  43543=>"010001011",
  43544=>"001110111",
  43545=>"010111100",
  43546=>"001001110",
  43547=>"110010001",
  43548=>"101000101",
  43549=>"110000101",
  43550=>"101111110",
  43551=>"101110000",
  43552=>"100100101",
  43553=>"101111110",
  43554=>"100001011",
  43555=>"000110111",
  43556=>"001101111",
  43557=>"000001001",
  43558=>"011101111",
  43559=>"010110011",
  43560=>"001001110",
  43561=>"011001011",
  43562=>"110101111",
  43563=>"000010101",
  43564=>"011100111",
  43565=>"001100111",
  43566=>"100111011",
  43567=>"101010000",
  43568=>"111110010",
  43569=>"010011101",
  43570=>"000001111",
  43571=>"000111001",
  43572=>"111100101",
  43573=>"011000100",
  43574=>"100000000",
  43575=>"001000111",
  43576=>"111001111",
  43577=>"010101100",
  43578=>"000011110",
  43579=>"001111010",
  43580=>"011100011",
  43581=>"100100010",
  43582=>"101101110",
  43583=>"100100100",
  43584=>"111111111",
  43585=>"011000000",
  43586=>"000010101",
  43587=>"011010001",
  43588=>"000000111",
  43589=>"000100011",
  43590=>"000011100",
  43591=>"001110111",
  43592=>"011011000",
  43593=>"111000000",
  43594=>"101001011",
  43595=>"000110110",
  43596=>"000011010",
  43597=>"010111000",
  43598=>"011000111",
  43599=>"011011100",
  43600=>"000110000",
  43601=>"111000100",
  43602=>"010101111",
  43603=>"001101010",
  43604=>"011010110",
  43605=>"010001011",
  43606=>"011111011",
  43607=>"011000100",
  43608=>"000110010",
  43609=>"100101110",
  43610=>"110111011",
  43611=>"111111010",
  43612=>"001110100",
  43613=>"000001010",
  43614=>"111100111",
  43615=>"111101111",
  43616=>"011010100",
  43617=>"101101100",
  43618=>"001011111",
  43619=>"001111100",
  43620=>"111011111",
  43621=>"111010110",
  43622=>"101110111",
  43623=>"001101011",
  43624=>"001000101",
  43625=>"001010011",
  43626=>"101000011",
  43627=>"000101011",
  43628=>"111110000",
  43629=>"001011001",
  43630=>"001111111",
  43631=>"001111100",
  43632=>"000011100",
  43633=>"000001100",
  43634=>"110100001",
  43635=>"111010110",
  43636=>"110111001",
  43637=>"110001000",
  43638=>"111011011",
  43639=>"101110000",
  43640=>"110000001",
  43641=>"010111100",
  43642=>"001010111",
  43643=>"000011100",
  43644=>"111001010",
  43645=>"000001000",
  43646=>"001011011",
  43647=>"010101010",
  43648=>"000001111",
  43649=>"111111010",
  43650=>"111011000",
  43651=>"011010101",
  43652=>"000010010",
  43653=>"101010010",
  43654=>"101010010",
  43655=>"011111011",
  43656=>"000010000",
  43657=>"100100000",
  43658=>"001111110",
  43659=>"010100000",
  43660=>"100000001",
  43661=>"001110110",
  43662=>"010100000",
  43663=>"111111110",
  43664=>"010111100",
  43665=>"101111111",
  43666=>"111000101",
  43667=>"000100111",
  43668=>"000100111",
  43669=>"101110000",
  43670=>"111001100",
  43671=>"100111110",
  43672=>"111100011",
  43673=>"100101000",
  43674=>"011011000",
  43675=>"010011000",
  43676=>"000000010",
  43677=>"000101011",
  43678=>"100101010",
  43679=>"101010010",
  43680=>"001010000",
  43681=>"110101110",
  43682=>"001110001",
  43683=>"000111010",
  43684=>"101011101",
  43685=>"001011011",
  43686=>"111000111",
  43687=>"001000010",
  43688=>"000010001",
  43689=>"010110110",
  43690=>"101110101",
  43691=>"111000001",
  43692=>"111000100",
  43693=>"000110110",
  43694=>"101110010",
  43695=>"001000111",
  43696=>"100001101",
  43697=>"111011111",
  43698=>"000101011",
  43699=>"000101111",
  43700=>"000011110",
  43701=>"100000111",
  43702=>"000001101",
  43703=>"010010000",
  43704=>"011111110",
  43705=>"010000000",
  43706=>"000111110",
  43707=>"100100001",
  43708=>"001101111",
  43709=>"100001100",
  43710=>"000101110",
  43711=>"010000110",
  43712=>"011011111",
  43713=>"110101011",
  43714=>"100111010",
  43715=>"111100001",
  43716=>"001110100",
  43717=>"100111111",
  43718=>"011111101",
  43719=>"010011100",
  43720=>"011100110",
  43721=>"101011011",
  43722=>"101111111",
  43723=>"011111001",
  43724=>"100110100",
  43725=>"011110111",
  43726=>"100000001",
  43727=>"100001010",
  43728=>"001110110",
  43729=>"101001100",
  43730=>"110111011",
  43731=>"101010110",
  43732=>"001011100",
  43733=>"111100101",
  43734=>"000000100",
  43735=>"010100000",
  43736=>"001111110",
  43737=>"100111111",
  43738=>"011101101",
  43739=>"010000001",
  43740=>"100000011",
  43741=>"010000010",
  43742=>"011111111",
  43743=>"010110010",
  43744=>"000010100",
  43745=>"100101100",
  43746=>"000000101",
  43747=>"111111110",
  43748=>"000011110",
  43749=>"110101011",
  43750=>"000001100",
  43751=>"100010100",
  43752=>"100111001",
  43753=>"110111111",
  43754=>"010101110",
  43755=>"101011010",
  43756=>"011100000",
  43757=>"111100011",
  43758=>"110011111",
  43759=>"000100101",
  43760=>"111111101",
  43761=>"001101010",
  43762=>"100010101",
  43763=>"011111000",
  43764=>"001101101",
  43765=>"001001011",
  43766=>"110111001",
  43767=>"100110011",
  43768=>"001001011",
  43769=>"111101110",
  43770=>"110011111",
  43771=>"110010111",
  43772=>"001000100",
  43773=>"101100011",
  43774=>"100000101",
  43775=>"101110111",
  43776=>"100010110",
  43777=>"010010010",
  43778=>"000001001",
  43779=>"110011110",
  43780=>"111010001",
  43781=>"001110001",
  43782=>"011001000",
  43783=>"101100110",
  43784=>"010101101",
  43785=>"110001001",
  43786=>"111000101",
  43787=>"000000100",
  43788=>"111011010",
  43789=>"000110101",
  43790=>"001101100",
  43791=>"110001000",
  43792=>"010010110",
  43793=>"000111000",
  43794=>"000000110",
  43795=>"100011101",
  43796=>"100000111",
  43797=>"100101010",
  43798=>"110000010",
  43799=>"001101011",
  43800=>"010010110",
  43801=>"000000111",
  43802=>"011001110",
  43803=>"001000011",
  43804=>"101010000",
  43805=>"101111011",
  43806=>"011010001",
  43807=>"011110000",
  43808=>"000001000",
  43809=>"111110110",
  43810=>"100100001",
  43811=>"010110110",
  43812=>"001111011",
  43813=>"000000011",
  43814=>"001011111",
  43815=>"000001101",
  43816=>"100000111",
  43817=>"111000111",
  43818=>"101011110",
  43819=>"110011011",
  43820=>"111101001",
  43821=>"010011110",
  43822=>"001011101",
  43823=>"000001011",
  43824=>"111101001",
  43825=>"100010000",
  43826=>"010101101",
  43827=>"111111101",
  43828=>"001101100",
  43829=>"000010010",
  43830=>"110101001",
  43831=>"011100100",
  43832=>"101001101",
  43833=>"100000101",
  43834=>"001011101",
  43835=>"000010000",
  43836=>"110101000",
  43837=>"000000111",
  43838=>"101100000",
  43839=>"001000100",
  43840=>"100011011",
  43841=>"101100000",
  43842=>"101000001",
  43843=>"001110111",
  43844=>"101001010",
  43845=>"000110011",
  43846=>"010000100",
  43847=>"100110100",
  43848=>"110110100",
  43849=>"000110111",
  43850=>"111001001",
  43851=>"001100011",
  43852=>"000100000",
  43853=>"010010011",
  43854=>"011101011",
  43855=>"110001010",
  43856=>"000011000",
  43857=>"100101100",
  43858=>"011101010",
  43859=>"100111010",
  43860=>"000111110",
  43861=>"100111110",
  43862=>"101000100",
  43863=>"000000110",
  43864=>"111110010",
  43865=>"111010110",
  43866=>"100001011",
  43867=>"101001001",
  43868=>"000101100",
  43869=>"001100111",
  43870=>"100100101",
  43871=>"001110100",
  43872=>"001001001",
  43873=>"000101011",
  43874=>"101011001",
  43875=>"011101011",
  43876=>"100111110",
  43877=>"101010101",
  43878=>"110010101",
  43879=>"100111100",
  43880=>"110011010",
  43881=>"010001110",
  43882=>"010110100",
  43883=>"011100000",
  43884=>"100001011",
  43885=>"000010100",
  43886=>"000100001",
  43887=>"111100100",
  43888=>"011010100",
  43889=>"111100001",
  43890=>"110001001",
  43891=>"100101110",
  43892=>"011011111",
  43893=>"010000011",
  43894=>"001111100",
  43895=>"100101110",
  43896=>"001101010",
  43897=>"010110110",
  43898=>"111001101",
  43899=>"010100111",
  43900=>"010100000",
  43901=>"110011101",
  43902=>"000011001",
  43903=>"011001101",
  43904=>"111001001",
  43905=>"111100100",
  43906=>"100010000",
  43907=>"011001000",
  43908=>"100100000",
  43909=>"111110011",
  43910=>"000010011",
  43911=>"110011101",
  43912=>"111001111",
  43913=>"110101100",
  43914=>"001001010",
  43915=>"100111001",
  43916=>"001111011",
  43917=>"110101111",
  43918=>"100101011",
  43919=>"001101011",
  43920=>"100010111",
  43921=>"110100110",
  43922=>"000100011",
  43923=>"011111100",
  43924=>"101000110",
  43925=>"010101100",
  43926=>"001111011",
  43927=>"100011101",
  43928=>"111011011",
  43929=>"100100100",
  43930=>"101000000",
  43931=>"100110110",
  43932=>"001101000",
  43933=>"111111110",
  43934=>"100010000",
  43935=>"100001110",
  43936=>"100000111",
  43937=>"000111111",
  43938=>"000100001",
  43939=>"001101100",
  43940=>"011001110",
  43941=>"111000111",
  43942=>"011011111",
  43943=>"111101100",
  43944=>"000111100",
  43945=>"111001001",
  43946=>"111010000",
  43947=>"111001011",
  43948=>"001001100",
  43949=>"110100011",
  43950=>"010100000",
  43951=>"010111111",
  43952=>"110111100",
  43953=>"000011110",
  43954=>"101000101",
  43955=>"010100011",
  43956=>"110011000",
  43957=>"010000101",
  43958=>"101001101",
  43959=>"101100111",
  43960=>"101000001",
  43961=>"100100110",
  43962=>"001101010",
  43963=>"011000000",
  43964=>"111111110",
  43965=>"111010100",
  43966=>"000111100",
  43967=>"111110010",
  43968=>"011100101",
  43969=>"111101100",
  43970=>"101100101",
  43971=>"001110100",
  43972=>"110010001",
  43973=>"101011110",
  43974=>"010111100",
  43975=>"011011100",
  43976=>"001001111",
  43977=>"110010000",
  43978=>"101001100",
  43979=>"001010000",
  43980=>"000100101",
  43981=>"100000011",
  43982=>"010100000",
  43983=>"000100100",
  43984=>"010011000",
  43985=>"110101110",
  43986=>"110101010",
  43987=>"110110011",
  43988=>"000101111",
  43989=>"110100110",
  43990=>"110101001",
  43991=>"011100010",
  43992=>"001000110",
  43993=>"110000100",
  43994=>"001001101",
  43995=>"000001001",
  43996=>"101000000",
  43997=>"101111100",
  43998=>"000000001",
  43999=>"010110011",
  44000=>"010000110",
  44001=>"110000100",
  44002=>"110000000",
  44003=>"111001001",
  44004=>"001010010",
  44005=>"111100001",
  44006=>"000101100",
  44007=>"010110100",
  44008=>"010110000",
  44009=>"001010000",
  44010=>"011000000",
  44011=>"011111010",
  44012=>"010000100",
  44013=>"111011110",
  44014=>"100001111",
  44015=>"011010101",
  44016=>"011010011",
  44017=>"010000100",
  44018=>"100001111",
  44019=>"101000110",
  44020=>"001110111",
  44021=>"001011010",
  44022=>"001101011",
  44023=>"010110011",
  44024=>"111110101",
  44025=>"111101111",
  44026=>"001110010",
  44027=>"001010001",
  44028=>"001011011",
  44029=>"100001101",
  44030=>"010001101",
  44031=>"100111111",
  44032=>"010111110",
  44033=>"011100000",
  44034=>"001100011",
  44035=>"111111111",
  44036=>"101000100",
  44037=>"111011101",
  44038=>"001000011",
  44039=>"011111110",
  44040=>"100001101",
  44041=>"101100000",
  44042=>"100100001",
  44043=>"010011101",
  44044=>"100000111",
  44045=>"100001111",
  44046=>"000110010",
  44047=>"110111011",
  44048=>"111110100",
  44049=>"110000100",
  44050=>"000101010",
  44051=>"100111000",
  44052=>"000110100",
  44053=>"100101111",
  44054=>"110110000",
  44055=>"110101000",
  44056=>"001010101",
  44057=>"000010011",
  44058=>"110101000",
  44059=>"101001110",
  44060=>"111101000",
  44061=>"011101101",
  44062=>"101000101",
  44063=>"010110000",
  44064=>"001000000",
  44065=>"101110010",
  44066=>"100001100",
  44067=>"100011110",
  44068=>"100010010",
  44069=>"000011100",
  44070=>"011010111",
  44071=>"101101011",
  44072=>"110100000",
  44073=>"111011101",
  44074=>"101101010",
  44075=>"001011011",
  44076=>"000111101",
  44077=>"010110010",
  44078=>"000001100",
  44079=>"010010010",
  44080=>"001001010",
  44081=>"110110000",
  44082=>"101001010",
  44083=>"000010111",
  44084=>"011111111",
  44085=>"011111010",
  44086=>"000001010",
  44087=>"110000101",
  44088=>"010100001",
  44089=>"101000111",
  44090=>"001111101",
  44091=>"000100000",
  44092=>"001001011",
  44093=>"001011011",
  44094=>"101110101",
  44095=>"110011101",
  44096=>"101000011",
  44097=>"110011010",
  44098=>"110010011",
  44099=>"100100011",
  44100=>"010000010",
  44101=>"111101011",
  44102=>"011011010",
  44103=>"011000101",
  44104=>"011010011",
  44105=>"110100010",
  44106=>"001011111",
  44107=>"010110001",
  44108=>"100000111",
  44109=>"000000100",
  44110=>"110011111",
  44111=>"111010000",
  44112=>"010000011",
  44113=>"110001001",
  44114=>"100010011",
  44115=>"000011111",
  44116=>"100100000",
  44117=>"001101011",
  44118=>"010011000",
  44119=>"000111000",
  44120=>"010111001",
  44121=>"110111101",
  44122=>"011111010",
  44123=>"111100011",
  44124=>"000111111",
  44125=>"010101111",
  44126=>"100000001",
  44127=>"100001100",
  44128=>"100000000",
  44129=>"010110010",
  44130=>"000001100",
  44131=>"110001010",
  44132=>"100101001",
  44133=>"110100001",
  44134=>"000000001",
  44135=>"010101100",
  44136=>"100011011",
  44137=>"100101100",
  44138=>"110000100",
  44139=>"100101001",
  44140=>"110100000",
  44141=>"011010110",
  44142=>"110000101",
  44143=>"100001100",
  44144=>"100010110",
  44145=>"000100101",
  44146=>"001011011",
  44147=>"100010000",
  44148=>"011101101",
  44149=>"111000011",
  44150=>"111011111",
  44151=>"001011010",
  44152=>"000010010",
  44153=>"001111100",
  44154=>"010010010",
  44155=>"111001001",
  44156=>"010010010",
  44157=>"011000011",
  44158=>"111111110",
  44159=>"101000110",
  44160=>"000110010",
  44161=>"001001101",
  44162=>"111101001",
  44163=>"101110001",
  44164=>"101100110",
  44165=>"011000101",
  44166=>"000001100",
  44167=>"000010101",
  44168=>"100010110",
  44169=>"001010010",
  44170=>"010001000",
  44171=>"111011100",
  44172=>"100000010",
  44173=>"100101000",
  44174=>"100110110",
  44175=>"010101100",
  44176=>"001011101",
  44177=>"000110111",
  44178=>"101110001",
  44179=>"101100011",
  44180=>"000010000",
  44181=>"110111010",
  44182=>"011001100",
  44183=>"001111011",
  44184=>"101011001",
  44185=>"110010000",
  44186=>"110100011",
  44187=>"011010011",
  44188=>"010111001",
  44189=>"000110111",
  44190=>"001011011",
  44191=>"011001010",
  44192=>"001111001",
  44193=>"011101011",
  44194=>"110100000",
  44195=>"100011100",
  44196=>"111111111",
  44197=>"110000110",
  44198=>"111011010",
  44199=>"111011110",
  44200=>"001110011",
  44201=>"000000000",
  44202=>"011111110",
  44203=>"000110100",
  44204=>"100001111",
  44205=>"000010001",
  44206=>"111000011",
  44207=>"000101110",
  44208=>"011000100",
  44209=>"101100011",
  44210=>"100001110",
  44211=>"010000010",
  44212=>"001101011",
  44213=>"111011110",
  44214=>"110111001",
  44215=>"010111011",
  44216=>"100110001",
  44217=>"011010000",
  44218=>"010000010",
  44219=>"011110011",
  44220=>"100001011",
  44221=>"101000100",
  44222=>"010000010",
  44223=>"001011000",
  44224=>"010110101",
  44225=>"010110000",
  44226=>"001000011",
  44227=>"101100100",
  44228=>"010110110",
  44229=>"110101110",
  44230=>"000110001",
  44231=>"111101011",
  44232=>"110011111",
  44233=>"010111010",
  44234=>"010000001",
  44235=>"110100101",
  44236=>"111000001",
  44237=>"101011010",
  44238=>"000110011",
  44239=>"001011100",
  44240=>"000001100",
  44241=>"010010110",
  44242=>"110101000",
  44243=>"000001111",
  44244=>"001011011",
  44245=>"110110010",
  44246=>"000000111",
  44247=>"000101110",
  44248=>"000111010",
  44249=>"000100101",
  44250=>"000000101",
  44251=>"010000000",
  44252=>"011011000",
  44253=>"101111110",
  44254=>"001011001",
  44255=>"111010010",
  44256=>"000000110",
  44257=>"000011000",
  44258=>"110001010",
  44259=>"000000100",
  44260=>"001100111",
  44261=>"011100011",
  44262=>"110001010",
  44263=>"110001001",
  44264=>"100110001",
  44265=>"111001011",
  44266=>"010000100",
  44267=>"001101010",
  44268=>"101000001",
  44269=>"010011110",
  44270=>"001100000",
  44271=>"100100001",
  44272=>"010001001",
  44273=>"100010001",
  44274=>"100101001",
  44275=>"000100000",
  44276=>"101100110",
  44277=>"010000101",
  44278=>"011010110",
  44279=>"110011100",
  44280=>"001011111",
  44281=>"101010010",
  44282=>"111001100",
  44283=>"101001101",
  44284=>"000001110",
  44285=>"010111000",
  44286=>"101011100",
  44287=>"110001001",
  44288=>"100010101",
  44289=>"111001111",
  44290=>"111101010",
  44291=>"011111101",
  44292=>"000001000",
  44293=>"001110111",
  44294=>"100110110",
  44295=>"101101101",
  44296=>"011010000",
  44297=>"000001100",
  44298=>"100011110",
  44299=>"001010011",
  44300=>"010000001",
  44301=>"111011111",
  44302=>"010001000",
  44303=>"001101111",
  44304=>"010010111",
  44305=>"111010101",
  44306=>"101111110",
  44307=>"011010000",
  44308=>"110001111",
  44309=>"011100011",
  44310=>"100101111",
  44311=>"001111010",
  44312=>"011011110",
  44313=>"011010111",
  44314=>"100010001",
  44315=>"111110110",
  44316=>"111101110",
  44317=>"100000000",
  44318=>"101000010",
  44319=>"000000011",
  44320=>"000000110",
  44321=>"000010001",
  44322=>"000111101",
  44323=>"011111000",
  44324=>"010000101",
  44325=>"001010101",
  44326=>"000011111",
  44327=>"111111011",
  44328=>"010111100",
  44329=>"101110110",
  44330=>"001000100",
  44331=>"000001001",
  44332=>"000010111",
  44333=>"100110000",
  44334=>"010001110",
  44335=>"001101111",
  44336=>"000111111",
  44337=>"101011110",
  44338=>"111011110",
  44339=>"010001000",
  44340=>"110110111",
  44341=>"011011111",
  44342=>"100010100",
  44343=>"110010010",
  44344=>"000010010",
  44345=>"110010010",
  44346=>"100101001",
  44347=>"011100011",
  44348=>"011101110",
  44349=>"000011011",
  44350=>"000011110",
  44351=>"011000111",
  44352=>"110011000",
  44353=>"110100001",
  44354=>"000010010",
  44355=>"110101101",
  44356=>"111111101",
  44357=>"000101000",
  44358=>"001010101",
  44359=>"000001010",
  44360=>"111111010",
  44361=>"101101101",
  44362=>"100011101",
  44363=>"001110010",
  44364=>"011000001",
  44365=>"100110110",
  44366=>"100110000",
  44367=>"110111000",
  44368=>"101001110",
  44369=>"010001101",
  44370=>"001101110",
  44371=>"000101111",
  44372=>"000100010",
  44373=>"111110000",
  44374=>"101010000",
  44375=>"001110010",
  44376=>"010111101",
  44377=>"100111110",
  44378=>"001001000",
  44379=>"000101101",
  44380=>"011110101",
  44381=>"110111100",
  44382=>"111011010",
  44383=>"001111100",
  44384=>"100110010",
  44385=>"011100000",
  44386=>"001000000",
  44387=>"000000110",
  44388=>"100101001",
  44389=>"100101011",
  44390=>"101011011",
  44391=>"101111010",
  44392=>"110111001",
  44393=>"001000000",
  44394=>"110000001",
  44395=>"110010101",
  44396=>"000100100",
  44397=>"110001010",
  44398=>"001010011",
  44399=>"100101101",
  44400=>"110010011",
  44401=>"110100101",
  44402=>"011100001",
  44403=>"000010001",
  44404=>"111101001",
  44405=>"011010011",
  44406=>"111101101",
  44407=>"010100100",
  44408=>"000111101",
  44409=>"010100110",
  44410=>"100011111",
  44411=>"101000000",
  44412=>"011111110",
  44413=>"011000011",
  44414=>"011011011",
  44415=>"111111011",
  44416=>"010011010",
  44417=>"000010010",
  44418=>"100110100",
  44419=>"011100000",
  44420=>"001100110",
  44421=>"011010101",
  44422=>"111000010",
  44423=>"001010000",
  44424=>"110100101",
  44425=>"101101000",
  44426=>"001111101",
  44427=>"100011010",
  44428=>"000011000",
  44429=>"101010001",
  44430=>"100100100",
  44431=>"100110001",
  44432=>"111001010",
  44433=>"001010000",
  44434=>"101011011",
  44435=>"000011101",
  44436=>"011011000",
  44437=>"011000000",
  44438=>"011101101",
  44439=>"100101011",
  44440=>"101001010",
  44441=>"001001000",
  44442=>"000011000",
  44443=>"011101110",
  44444=>"000000011",
  44445=>"111101101",
  44446=>"010011010",
  44447=>"111111110",
  44448=>"000111000",
  44449=>"010100010",
  44450=>"000101101",
  44451=>"010111100",
  44452=>"111101101",
  44453=>"100010001",
  44454=>"010101001",
  44455=>"100010100",
  44456=>"000000001",
  44457=>"110110101",
  44458=>"101101001",
  44459=>"010000101",
  44460=>"111110000",
  44461=>"011110000",
  44462=>"001111101",
  44463=>"010011110",
  44464=>"000110000",
  44465=>"000111100",
  44466=>"011101100",
  44467=>"101111010",
  44468=>"011000101",
  44469=>"110001010",
  44470=>"110101111",
  44471=>"111011111",
  44472=>"110110101",
  44473=>"100110010",
  44474=>"000101100",
  44475=>"000010001",
  44476=>"100001100",
  44477=>"110110001",
  44478=>"101011011",
  44479=>"001001101",
  44480=>"000111100",
  44481=>"011010010",
  44482=>"011101010",
  44483=>"001101011",
  44484=>"100110101",
  44485=>"100100101",
  44486=>"100000001",
  44487=>"100000101",
  44488=>"111100000",
  44489=>"001010101",
  44490=>"100101011",
  44491=>"011110101",
  44492=>"100110010",
  44493=>"000011001",
  44494=>"101000010",
  44495=>"101000010",
  44496=>"110100001",
  44497=>"101100011",
  44498=>"010101011",
  44499=>"001110111",
  44500=>"000101111",
  44501=>"000000111",
  44502=>"000010100",
  44503=>"010000100",
  44504=>"000101001",
  44505=>"101001010",
  44506=>"110000100",
  44507=>"011101111",
  44508=>"100010011",
  44509=>"101000110",
  44510=>"001111001",
  44511=>"101011101",
  44512=>"100011010",
  44513=>"011110001",
  44514=>"000000001",
  44515=>"101101011",
  44516=>"111100110",
  44517=>"100101101",
  44518=>"110110000",
  44519=>"000000000",
  44520=>"111111110",
  44521=>"000010010",
  44522=>"010001011",
  44523=>"110100111",
  44524=>"100000100",
  44525=>"111101000",
  44526=>"110100100",
  44527=>"100101101",
  44528=>"011011011",
  44529=>"101111110",
  44530=>"111111100",
  44531=>"001111100",
  44532=>"100000000",
  44533=>"111111010",
  44534=>"010001000",
  44535=>"011111110",
  44536=>"100000000",
  44537=>"100100000",
  44538=>"100000111",
  44539=>"000001101",
  44540=>"101110010",
  44541=>"001111001",
  44542=>"111001110",
  44543=>"010011001",
  44544=>"000110101",
  44545=>"011000000",
  44546=>"101100011",
  44547=>"110001111",
  44548=>"001111101",
  44549=>"001100000",
  44550=>"101001101",
  44551=>"000101010",
  44552=>"100011000",
  44553=>"010100010",
  44554=>"000110001",
  44555=>"010101111",
  44556=>"000001110",
  44557=>"011110111",
  44558=>"000100101",
  44559=>"110000111",
  44560=>"101100101",
  44561=>"101111000",
  44562=>"010110000",
  44563=>"111001101",
  44564=>"010111111",
  44565=>"010110101",
  44566=>"110001011",
  44567=>"001001101",
  44568=>"010001011",
  44569=>"010011011",
  44570=>"111101010",
  44571=>"110011101",
  44572=>"111000001",
  44573=>"111011101",
  44574=>"101100110",
  44575=>"110110011",
  44576=>"011011010",
  44577=>"111000100",
  44578=>"100101011",
  44579=>"011101110",
  44580=>"111101110",
  44581=>"100011011",
  44582=>"000110110",
  44583=>"001001001",
  44584=>"110100000",
  44585=>"111110111",
  44586=>"001010010",
  44587=>"100111110",
  44588=>"001000010",
  44589=>"001010110",
  44590=>"100000000",
  44591=>"010100010",
  44592=>"011000010",
  44593=>"010110111",
  44594=>"011101111",
  44595=>"110000111",
  44596=>"011000011",
  44597=>"110000110",
  44598=>"000000100",
  44599=>"000010110",
  44600=>"100110110",
  44601=>"111010011",
  44602=>"010000001",
  44603=>"111111010",
  44604=>"000000011",
  44605=>"010000011",
  44606=>"011001101",
  44607=>"000101100",
  44608=>"101111000",
  44609=>"101000101",
  44610=>"001001111",
  44611=>"000111001",
  44612=>"111010100",
  44613=>"011101111",
  44614=>"001110110",
  44615=>"110010011",
  44616=>"001110010",
  44617=>"101100110",
  44618=>"001001001",
  44619=>"100011011",
  44620=>"010111111",
  44621=>"100101101",
  44622=>"100011000",
  44623=>"001001000",
  44624=>"010010010",
  44625=>"001001101",
  44626=>"011100111",
  44627=>"000100001",
  44628=>"011000110",
  44629=>"101101011",
  44630=>"100110111",
  44631=>"110110110",
  44632=>"001000010",
  44633=>"110100011",
  44634=>"101000001",
  44635=>"010111100",
  44636=>"110011101",
  44637=>"100100000",
  44638=>"111001111",
  44639=>"110001011",
  44640=>"111111001",
  44641=>"000101111",
  44642=>"011001010",
  44643=>"001100110",
  44644=>"000110001",
  44645=>"101100000",
  44646=>"010110000",
  44647=>"110100001",
  44648=>"000100011",
  44649=>"110111100",
  44650=>"110000000",
  44651=>"111101011",
  44652=>"001000001",
  44653=>"101000100",
  44654=>"011110010",
  44655=>"000110111",
  44656=>"100011011",
  44657=>"000000001",
  44658=>"000101001",
  44659=>"000010100",
  44660=>"000111010",
  44661=>"000110001",
  44662=>"111011101",
  44663=>"011100011",
  44664=>"100101000",
  44665=>"001001011",
  44666=>"111111111",
  44667=>"111011101",
  44668=>"011100000",
  44669=>"101101001",
  44670=>"010110001",
  44671=>"010101110",
  44672=>"111111010",
  44673=>"000001100",
  44674=>"111111011",
  44675=>"001001101",
  44676=>"010010001",
  44677=>"010111000",
  44678=>"111110110",
  44679=>"101010010",
  44680=>"110011111",
  44681=>"001000111",
  44682=>"100011010",
  44683=>"100111001",
  44684=>"010000011",
  44685=>"001001001",
  44686=>"010010100",
  44687=>"000100001",
  44688=>"001111010",
  44689=>"000000011",
  44690=>"110001100",
  44691=>"010011110",
  44692=>"111100000",
  44693=>"011111000",
  44694=>"110101000",
  44695=>"101101100",
  44696=>"001011001",
  44697=>"011000001",
  44698=>"000110110",
  44699=>"110111100",
  44700=>"000100000",
  44701=>"110011011",
  44702=>"101010100",
  44703=>"000000011",
  44704=>"000101011",
  44705=>"000101100",
  44706=>"101111000",
  44707=>"101010100",
  44708=>"010010111",
  44709=>"000100101",
  44710=>"100111100",
  44711=>"000000000",
  44712=>"110100100",
  44713=>"100110100",
  44714=>"010110000",
  44715=>"000000001",
  44716=>"010110011",
  44717=>"000111100",
  44718=>"111010001",
  44719=>"111101000",
  44720=>"000011011",
  44721=>"100000011",
  44722=>"010110011",
  44723=>"111100001",
  44724=>"100001110",
  44725=>"111111111",
  44726=>"011101001",
  44727=>"000000011",
  44728=>"000011011",
  44729=>"001101100",
  44730=>"000000010",
  44731=>"110000010",
  44732=>"011110001",
  44733=>"001000011",
  44734=>"000000001",
  44735=>"011110001",
  44736=>"011001010",
  44737=>"011111100",
  44738=>"001010000",
  44739=>"010000110",
  44740=>"111011110",
  44741=>"100001101",
  44742=>"010100100",
  44743=>"001101000",
  44744=>"000001101",
  44745=>"100001110",
  44746=>"110001110",
  44747=>"100110011",
  44748=>"101001100",
  44749=>"100110011",
  44750=>"010001111",
  44751=>"110101011",
  44752=>"000000111",
  44753=>"111000101",
  44754=>"110110001",
  44755=>"101010000",
  44756=>"110100110",
  44757=>"100011111",
  44758=>"111000010",
  44759=>"010111000",
  44760=>"011010001",
  44761=>"110010011",
  44762=>"111100101",
  44763=>"001001010",
  44764=>"100010101",
  44765=>"100001110",
  44766=>"100000010",
  44767=>"100010010",
  44768=>"001010010",
  44769=>"001000001",
  44770=>"111011010",
  44771=>"101110111",
  44772=>"101011001",
  44773=>"010100001",
  44774=>"000001000",
  44775=>"010011110",
  44776=>"110101010",
  44777=>"001110110",
  44778=>"100011101",
  44779=>"101110011",
  44780=>"010000111",
  44781=>"100101010",
  44782=>"000110000",
  44783=>"111111111",
  44784=>"011101000",
  44785=>"101001111",
  44786=>"110000110",
  44787=>"110111011",
  44788=>"111010100",
  44789=>"110001011",
  44790=>"011000001",
  44791=>"111110110",
  44792=>"100000000",
  44793=>"010011111",
  44794=>"001000110",
  44795=>"010111111",
  44796=>"111001101",
  44797=>"011001101",
  44798=>"011011100",
  44799=>"011111101",
  44800=>"000110010",
  44801=>"100100111",
  44802=>"000110001",
  44803=>"010000001",
  44804=>"000111100",
  44805=>"000011010",
  44806=>"000000011",
  44807=>"101100001",
  44808=>"100000001",
  44809=>"101110100",
  44810=>"010100101",
  44811=>"101101100",
  44812=>"000001111",
  44813=>"111000011",
  44814=>"101100010",
  44815=>"111100100",
  44816=>"010010100",
  44817=>"011110101",
  44818=>"110010100",
  44819=>"100010101",
  44820=>"110101111",
  44821=>"000000100",
  44822=>"101101001",
  44823=>"001011111",
  44824=>"001010001",
  44825=>"001111010",
  44826=>"011111011",
  44827=>"010111011",
  44828=>"111001011",
  44829=>"001011111",
  44830=>"000100011",
  44831=>"101010010",
  44832=>"100101000",
  44833=>"011101101",
  44834=>"100111001",
  44835=>"000100010",
  44836=>"001101001",
  44837=>"101000100",
  44838=>"011100000",
  44839=>"100010100",
  44840=>"001000010",
  44841=>"111100111",
  44842=>"101100111",
  44843=>"111010001",
  44844=>"000001010",
  44845=>"000111110",
  44846=>"101100011",
  44847=>"110110111",
  44848=>"010100000",
  44849=>"000011001",
  44850=>"001000010",
  44851=>"101101010",
  44852=>"100000010",
  44853=>"111100001",
  44854=>"000011111",
  44855=>"101111010",
  44856=>"101111011",
  44857=>"011110010",
  44858=>"011011000",
  44859=>"011001011",
  44860=>"110010011",
  44861=>"001001011",
  44862=>"000101000",
  44863=>"001111000",
  44864=>"001101111",
  44865=>"111011110",
  44866=>"100101101",
  44867=>"000111101",
  44868=>"000000000",
  44869=>"000010111",
  44870=>"000101100",
  44871=>"011010000",
  44872=>"101100101",
  44873=>"010011000",
  44874=>"010001001",
  44875=>"001111010",
  44876=>"010001100",
  44877=>"101111110",
  44878=>"101101000",
  44879=>"010001101",
  44880=>"100011010",
  44881=>"100100101",
  44882=>"000000011",
  44883=>"101101101",
  44884=>"001000001",
  44885=>"110110100",
  44886=>"001010110",
  44887=>"101100011",
  44888=>"001110000",
  44889=>"011001110",
  44890=>"001001011",
  44891=>"101000010",
  44892=>"111011101",
  44893=>"110101111",
  44894=>"011011111",
  44895=>"000000001",
  44896=>"000010111",
  44897=>"001010101",
  44898=>"011100010",
  44899=>"111010000",
  44900=>"011000000",
  44901=>"100010001",
  44902=>"000010010",
  44903=>"110111000",
  44904=>"110000110",
  44905=>"111101100",
  44906=>"011000010",
  44907=>"011010101",
  44908=>"011110100",
  44909=>"101101111",
  44910=>"100000111",
  44911=>"010011110",
  44912=>"000100001",
  44913=>"010100110",
  44914=>"010011001",
  44915=>"110001011",
  44916=>"000111000",
  44917=>"111110100",
  44918=>"010010010",
  44919=>"000001001",
  44920=>"001001000",
  44921=>"001101110",
  44922=>"101000001",
  44923=>"011111000",
  44924=>"100010101",
  44925=>"001101000",
  44926=>"101001110",
  44927=>"100100100",
  44928=>"011101000",
  44929=>"001101111",
  44930=>"001011011",
  44931=>"010011010",
  44932=>"110001100",
  44933=>"011011101",
  44934=>"111100101",
  44935=>"100000111",
  44936=>"001111000",
  44937=>"000010000",
  44938=>"101111010",
  44939=>"100011001",
  44940=>"011111011",
  44941=>"000100100",
  44942=>"000001010",
  44943=>"100011001",
  44944=>"100111111",
  44945=>"011000111",
  44946=>"000110101",
  44947=>"100000110",
  44948=>"010011010",
  44949=>"101011100",
  44950=>"000001011",
  44951=>"111001110",
  44952=>"010100111",
  44953=>"001110100",
  44954=>"111110111",
  44955=>"000011100",
  44956=>"111000010",
  44957=>"111111100",
  44958=>"010110101",
  44959=>"110000110",
  44960=>"001011111",
  44961=>"100000000",
  44962=>"101101101",
  44963=>"101100101",
  44964=>"001000101",
  44965=>"001111000",
  44966=>"101111010",
  44967=>"011001111",
  44968=>"001100110",
  44969=>"100010100",
  44970=>"111111001",
  44971=>"000001011",
  44972=>"001000111",
  44973=>"010001001",
  44974=>"110110111",
  44975=>"010001110",
  44976=>"001100011",
  44977=>"111110011",
  44978=>"011100001",
  44979=>"000001001",
  44980=>"111010011",
  44981=>"011000010",
  44982=>"101111111",
  44983=>"000001110",
  44984=>"111000101",
  44985=>"000001110",
  44986=>"110011001",
  44987=>"111110101",
  44988=>"000111011",
  44989=>"110001001",
  44990=>"111001001",
  44991=>"100001010",
  44992=>"111101011",
  44993=>"010011000",
  44994=>"101101101",
  44995=>"011000000",
  44996=>"111101100",
  44997=>"101000110",
  44998=>"000000111",
  44999=>"010011100",
  45000=>"000111011",
  45001=>"010000000",
  45002=>"101011010",
  45003=>"000011100",
  45004=>"000010110",
  45005=>"101011010",
  45006=>"001000110",
  45007=>"001100111",
  45008=>"110000110",
  45009=>"000010011",
  45010=>"011111001",
  45011=>"000100100",
  45012=>"010011110",
  45013=>"011000110",
  45014=>"011101011",
  45015=>"011111100",
  45016=>"000000000",
  45017=>"110111011",
  45018=>"100010001",
  45019=>"010010100",
  45020=>"111001001",
  45021=>"010011101",
  45022=>"101010101",
  45023=>"011110011",
  45024=>"000100001",
  45025=>"100111001",
  45026=>"101001100",
  45027=>"011001000",
  45028=>"000000010",
  45029=>"000101110",
  45030=>"010110000",
  45031=>"000010111",
  45032=>"100011100",
  45033=>"000111101",
  45034=>"001000110",
  45035=>"000101100",
  45036=>"111001110",
  45037=>"111010001",
  45038=>"010111111",
  45039=>"010101010",
  45040=>"000010100",
  45041=>"000110011",
  45042=>"001011011",
  45043=>"010011101",
  45044=>"111110011",
  45045=>"001111111",
  45046=>"010110101",
  45047=>"011011101",
  45048=>"110001000",
  45049=>"011101010",
  45050=>"011000001",
  45051=>"000111010",
  45052=>"001011011",
  45053=>"101000111",
  45054=>"010010010",
  45055=>"001011011",
  45056=>"100111101",
  45057=>"111111011",
  45058=>"000101110",
  45059=>"010110000",
  45060=>"110110001",
  45061=>"001111011",
  45062=>"101110111",
  45063=>"000000111",
  45064=>"100111001",
  45065=>"100101111",
  45066=>"010011101",
  45067=>"101010101",
  45068=>"100011111",
  45069=>"001011101",
  45070=>"010010110",
  45071=>"010101011",
  45072=>"000011010",
  45073=>"101100101",
  45074=>"101100011",
  45075=>"100000011",
  45076=>"100000010",
  45077=>"001101011",
  45078=>"101010001",
  45079=>"101000001",
  45080=>"010101111",
  45081=>"101001001",
  45082=>"011100101",
  45083=>"001110110",
  45084=>"111001000",
  45085=>"110100011",
  45086=>"111010000",
  45087=>"000011100",
  45088=>"101100010",
  45089=>"100001001",
  45090=>"111100010",
  45091=>"000011101",
  45092=>"010111111",
  45093=>"110001011",
  45094=>"000000101",
  45095=>"000101010",
  45096=>"011100111",
  45097=>"010100101",
  45098=>"010100111",
  45099=>"100001101",
  45100=>"011000101",
  45101=>"011101011",
  45102=>"011110111",
  45103=>"101001011",
  45104=>"011001001",
  45105=>"000000000",
  45106=>"000110101",
  45107=>"001010001",
  45108=>"101001110",
  45109=>"100000000",
  45110=>"010111110",
  45111=>"010111101",
  45112=>"101101110",
  45113=>"100000000",
  45114=>"010010110",
  45115=>"100111111",
  45116=>"100000001",
  45117=>"111110000",
  45118=>"111110000",
  45119=>"100000000",
  45120=>"010100001",
  45121=>"001001000",
  45122=>"001010001",
  45123=>"100010011",
  45124=>"101111111",
  45125=>"001100110",
  45126=>"100111000",
  45127=>"010001011",
  45128=>"000001101",
  45129=>"001001011",
  45130=>"111000101",
  45131=>"000100011",
  45132=>"100000000",
  45133=>"010000010",
  45134=>"001111011",
  45135=>"111010101",
  45136=>"111001101",
  45137=>"100111110",
  45138=>"011110111",
  45139=>"011110111",
  45140=>"001110011",
  45141=>"100010001",
  45142=>"101111100",
  45143=>"010100010",
  45144=>"101000101",
  45145=>"000101000",
  45146=>"111111011",
  45147=>"001001011",
  45148=>"110111010",
  45149=>"000100000",
  45150=>"001110101",
  45151=>"011000000",
  45152=>"000010101",
  45153=>"010010010",
  45154=>"100000011",
  45155=>"001100111",
  45156=>"010101111",
  45157=>"011010100",
  45158=>"101001111",
  45159=>"000010010",
  45160=>"110010101",
  45161=>"011011110",
  45162=>"100101000",
  45163=>"010101001",
  45164=>"001001010",
  45165=>"100001010",
  45166=>"010110010",
  45167=>"111101101",
  45168=>"001101100",
  45169=>"111001111",
  45170=>"100010000",
  45171=>"100010101",
  45172=>"101101101",
  45173=>"001011001",
  45174=>"100111100",
  45175=>"001000000",
  45176=>"111101001",
  45177=>"011011011",
  45178=>"111010000",
  45179=>"100011100",
  45180=>"110001011",
  45181=>"110111101",
  45182=>"101101101",
  45183=>"100110000",
  45184=>"001001110",
  45185=>"000010010",
  45186=>"000000001",
  45187=>"000000010",
  45188=>"101011001",
  45189=>"110111111",
  45190=>"010001010",
  45191=>"011011011",
  45192=>"000110001",
  45193=>"011011011",
  45194=>"010001000",
  45195=>"010111111",
  45196=>"011100000",
  45197=>"101010101",
  45198=>"111010010",
  45199=>"101011001",
  45200=>"011110001",
  45201=>"100011011",
  45202=>"101101101",
  45203=>"000000011",
  45204=>"010110011",
  45205=>"001010110",
  45206=>"101110110",
  45207=>"000001001",
  45208=>"000011010",
  45209=>"001100011",
  45210=>"011110110",
  45211=>"100011110",
  45212=>"011100010",
  45213=>"110101101",
  45214=>"101001010",
  45215=>"010010010",
  45216=>"001111110",
  45217=>"011000100",
  45218=>"110100010",
  45219=>"010110100",
  45220=>"010101100",
  45221=>"110000000",
  45222=>"100011001",
  45223=>"001101110",
  45224=>"110110011",
  45225=>"100011000",
  45226=>"110001010",
  45227=>"110101011",
  45228=>"110000100",
  45229=>"000001110",
  45230=>"010111110",
  45231=>"110100010",
  45232=>"101110011",
  45233=>"110101110",
  45234=>"111000001",
  45235=>"001011001",
  45236=>"111100100",
  45237=>"001101001",
  45238=>"001001101",
  45239=>"100001110",
  45240=>"101011100",
  45241=>"000011100",
  45242=>"100011101",
  45243=>"001100001",
  45244=>"101010110",
  45245=>"010000110",
  45246=>"101011000",
  45247=>"000100100",
  45248=>"010001010",
  45249=>"111110101",
  45250=>"001100000",
  45251=>"101100000",
  45252=>"110100111",
  45253=>"101110111",
  45254=>"110111110",
  45255=>"110000001",
  45256=>"110010000",
  45257=>"101111010",
  45258=>"101101000",
  45259=>"110111101",
  45260=>"110000010",
  45261=>"110111101",
  45262=>"011101111",
  45263=>"101000001",
  45264=>"101101010",
  45265=>"101010001",
  45266=>"100010101",
  45267=>"111110010",
  45268=>"110100000",
  45269=>"110111111",
  45270=>"011111100",
  45271=>"101010011",
  45272=>"100101011",
  45273=>"101010111",
  45274=>"000011000",
  45275=>"100010011",
  45276=>"010111011",
  45277=>"101110100",
  45278=>"000111010",
  45279=>"100001000",
  45280=>"011110101",
  45281=>"001010011",
  45282=>"111011010",
  45283=>"111011100",
  45284=>"011111110",
  45285=>"010010011",
  45286=>"111010011",
  45287=>"111110011",
  45288=>"110000100",
  45289=>"001101110",
  45290=>"110101011",
  45291=>"111110000",
  45292=>"111111110",
  45293=>"011000000",
  45294=>"011011100",
  45295=>"001110110",
  45296=>"110101000",
  45297=>"111101100",
  45298=>"100111010",
  45299=>"101111011",
  45300=>"110010010",
  45301=>"101011111",
  45302=>"010110100",
  45303=>"000000010",
  45304=>"000011010",
  45305=>"001111100",
  45306=>"011010001",
  45307=>"000000010",
  45308=>"100001010",
  45309=>"110010000",
  45310=>"000010001",
  45311=>"011011111",
  45312=>"011110100",
  45313=>"101011011",
  45314=>"101100111",
  45315=>"000110011",
  45316=>"101000101",
  45317=>"111001000",
  45318=>"001010100",
  45319=>"100100100",
  45320=>"111100011",
  45321=>"100000111",
  45322=>"000101011",
  45323=>"100000111",
  45324=>"011010001",
  45325=>"011001001",
  45326=>"001111000",
  45327=>"001101000",
  45328=>"111101011",
  45329=>"000000100",
  45330=>"110110101",
  45331=>"110001110",
  45332=>"101100110",
  45333=>"001010011",
  45334=>"100011011",
  45335=>"011000010",
  45336=>"011110110",
  45337=>"101111111",
  45338=>"100100010",
  45339=>"110001000",
  45340=>"011010001",
  45341=>"011111000",
  45342=>"011101101",
  45343=>"001100010",
  45344=>"100000011",
  45345=>"110001111",
  45346=>"010001000",
  45347=>"110000111",
  45348=>"110110010",
  45349=>"110100010",
  45350=>"111010011",
  45351=>"100000000",
  45352=>"001111110",
  45353=>"111000110",
  45354=>"011100010",
  45355=>"011001001",
  45356=>"010010111",
  45357=>"010011011",
  45358=>"101111000",
  45359=>"000111011",
  45360=>"010000110",
  45361=>"010110111",
  45362=>"011110111",
  45363=>"111111010",
  45364=>"101110010",
  45365=>"001011011",
  45366=>"111110101",
  45367=>"111101001",
  45368=>"001110100",
  45369=>"100111011",
  45370=>"011111011",
  45371=>"111110010",
  45372=>"100100010",
  45373=>"111101110",
  45374=>"010110100",
  45375=>"011000000",
  45376=>"101001011",
  45377=>"001001000",
  45378=>"001100101",
  45379=>"010000011",
  45380=>"110101101",
  45381=>"110000100",
  45382=>"001100100",
  45383=>"011110001",
  45384=>"100111101",
  45385=>"100000110",
  45386=>"011101010",
  45387=>"101001111",
  45388=>"010000010",
  45389=>"110100110",
  45390=>"010110000",
  45391=>"110001110",
  45392=>"100011111",
  45393=>"100101000",
  45394=>"010100010",
  45395=>"000000000",
  45396=>"000110110",
  45397=>"000101001",
  45398=>"000101011",
  45399=>"100001001",
  45400=>"110100011",
  45401=>"110100001",
  45402=>"000011100",
  45403=>"010100000",
  45404=>"100000001",
  45405=>"100011011",
  45406=>"001010001",
  45407=>"001100000",
  45408=>"011101001",
  45409=>"101000011",
  45410=>"001111101",
  45411=>"110001110",
  45412=>"111111000",
  45413=>"001000100",
  45414=>"000010101",
  45415=>"100010100",
  45416=>"110111100",
  45417=>"010000100",
  45418=>"011101111",
  45419=>"010001001",
  45420=>"010010100",
  45421=>"011101010",
  45422=>"011111111",
  45423=>"101111111",
  45424=>"100010111",
  45425=>"000000000",
  45426=>"100111110",
  45427=>"011110110",
  45428=>"011100010",
  45429=>"111111110",
  45430=>"001000101",
  45431=>"011011011",
  45432=>"100110000",
  45433=>"111101101",
  45434=>"000011001",
  45435=>"011101001",
  45436=>"111101000",
  45437=>"101111100",
  45438=>"101110000",
  45439=>"011100111",
  45440=>"111100010",
  45441=>"001010000",
  45442=>"011110110",
  45443=>"101100101",
  45444=>"000101110",
  45445=>"011000110",
  45446=>"101000110",
  45447=>"000001100",
  45448=>"000110010",
  45449=>"010111011",
  45450=>"111101000",
  45451=>"101001011",
  45452=>"111110111",
  45453=>"001010000",
  45454=>"111011010",
  45455=>"011100110",
  45456=>"101110011",
  45457=>"100001100",
  45458=>"110111110",
  45459=>"111010001",
  45460=>"011101001",
  45461=>"100001011",
  45462=>"011010011",
  45463=>"011001100",
  45464=>"101110100",
  45465=>"110001010",
  45466=>"010100000",
  45467=>"000010110",
  45468=>"111000001",
  45469=>"101001001",
  45470=>"011011111",
  45471=>"100001101",
  45472=>"010101000",
  45473=>"000101110",
  45474=>"000000001",
  45475=>"100001100",
  45476=>"111111110",
  45477=>"100100011",
  45478=>"110101100",
  45479=>"111001110",
  45480=>"010100101",
  45481=>"001110110",
  45482=>"100000111",
  45483=>"010000000",
  45484=>"111100011",
  45485=>"111111010",
  45486=>"100000101",
  45487=>"100001000",
  45488=>"011001100",
  45489=>"011110011",
  45490=>"011000010",
  45491=>"011001000",
  45492=>"111001000",
  45493=>"111010111",
  45494=>"001001011",
  45495=>"011111011",
  45496=>"010001001",
  45497=>"100001011",
  45498=>"110110011",
  45499=>"101100101",
  45500=>"111010100",
  45501=>"001011101",
  45502=>"001101011",
  45503=>"111000000",
  45504=>"101111101",
  45505=>"111000110",
  45506=>"001100101",
  45507=>"010001100",
  45508=>"100010000",
  45509=>"010000000",
  45510=>"010001110",
  45511=>"100000000",
  45512=>"011111101",
  45513=>"001111111",
  45514=>"101100100",
  45515=>"000011001",
  45516=>"111111100",
  45517=>"000011110",
  45518=>"000111111",
  45519=>"111111011",
  45520=>"100011001",
  45521=>"000001011",
  45522=>"000001011",
  45523=>"100100000",
  45524=>"100110111",
  45525=>"110001000",
  45526=>"100101001",
  45527=>"001000110",
  45528=>"010111001",
  45529=>"001110111",
  45530=>"110101011",
  45531=>"000000101",
  45532=>"011110101",
  45533=>"000011100",
  45534=>"111001100",
  45535=>"000011001",
  45536=>"000100010",
  45537=>"011000100",
  45538=>"101011010",
  45539=>"111101100",
  45540=>"101000110",
  45541=>"101100101",
  45542=>"011011101",
  45543=>"111111010",
  45544=>"100000000",
  45545=>"111001111",
  45546=>"000111111",
  45547=>"101000011",
  45548=>"010101100",
  45549=>"111111011",
  45550=>"100110010",
  45551=>"110001100",
  45552=>"111110011",
  45553=>"110010101",
  45554=>"111000010",
  45555=>"011100001",
  45556=>"101000011",
  45557=>"001011101",
  45558=>"010110000",
  45559=>"100101101",
  45560=>"010011001",
  45561=>"101000101",
  45562=>"111101011",
  45563=>"101010110",
  45564=>"010100100",
  45565=>"010001000",
  45566=>"100101011",
  45567=>"000100000",
  45568=>"111100011",
  45569=>"101000011",
  45570=>"110010101",
  45571=>"000100000",
  45572=>"100001001",
  45573=>"100010001",
  45574=>"100001001",
  45575=>"001111000",
  45576=>"110000100",
  45577=>"011101110",
  45578=>"000011011",
  45579=>"011011100",
  45580=>"011011010",
  45581=>"010100110",
  45582=>"011001100",
  45583=>"011101111",
  45584=>"010110001",
  45585=>"100110111",
  45586=>"011101101",
  45587=>"010000100",
  45588=>"100010010",
  45589=>"101010011",
  45590=>"010111100",
  45591=>"110100010",
  45592=>"101000111",
  45593=>"111010000",
  45594=>"010011110",
  45595=>"100011111",
  45596=>"110110100",
  45597=>"100110100",
  45598=>"111111111",
  45599=>"111001100",
  45600=>"110101001",
  45601=>"001110010",
  45602=>"001100000",
  45603=>"001011010",
  45604=>"000111000",
  45605=>"101110110",
  45606=>"101001011",
  45607=>"101011011",
  45608=>"110011110",
  45609=>"100000100",
  45610=>"110011010",
  45611=>"101001101",
  45612=>"110011011",
  45613=>"000101011",
  45614=>"110011110",
  45615=>"111000110",
  45616=>"011100001",
  45617=>"000111010",
  45618=>"111000111",
  45619=>"000001000",
  45620=>"000010000",
  45621=>"000001000",
  45622=>"010100001",
  45623=>"011000001",
  45624=>"110111011",
  45625=>"011011110",
  45626=>"111100101",
  45627=>"110101001",
  45628=>"100101101",
  45629=>"000000101",
  45630=>"010111100",
  45631=>"000001010",
  45632=>"010011111",
  45633=>"111010001",
  45634=>"000001000",
  45635=>"010011000",
  45636=>"000110000",
  45637=>"111110010",
  45638=>"101000000",
  45639=>"010110111",
  45640=>"100111100",
  45641=>"101001110",
  45642=>"101001010",
  45643=>"101101101",
  45644=>"010010010",
  45645=>"010000110",
  45646=>"000010111",
  45647=>"001001010",
  45648=>"010011000",
  45649=>"000100110",
  45650=>"001011110",
  45651=>"010000000",
  45652=>"011101000",
  45653=>"000000100",
  45654=>"101111000",
  45655=>"110100000",
  45656=>"001111110",
  45657=>"000001001",
  45658=>"101100010",
  45659=>"000111101",
  45660=>"000001110",
  45661=>"010001001",
  45662=>"111000000",
  45663=>"111001110",
  45664=>"001111010",
  45665=>"000000010",
  45666=>"011110101",
  45667=>"011101111",
  45668=>"000001001",
  45669=>"001111110",
  45670=>"000111000",
  45671=>"011010100",
  45672=>"000011101",
  45673=>"000001110",
  45674=>"010000010",
  45675=>"010101000",
  45676=>"001101000",
  45677=>"101011001",
  45678=>"011000101",
  45679=>"110011011",
  45680=>"111110110",
  45681=>"001011101",
  45682=>"100001100",
  45683=>"001001001",
  45684=>"111100101",
  45685=>"000001011",
  45686=>"101010110",
  45687=>"010000101",
  45688=>"101100011",
  45689=>"101101100",
  45690=>"110111000",
  45691=>"100000001",
  45692=>"001101110",
  45693=>"011110100",
  45694=>"000010111",
  45695=>"001101000",
  45696=>"010001010",
  45697=>"111101010",
  45698=>"110010010",
  45699=>"011001111",
  45700=>"001110001",
  45701=>"100001111",
  45702=>"111011111",
  45703=>"001101000",
  45704=>"111010110",
  45705=>"001110110",
  45706=>"011110011",
  45707=>"100011101",
  45708=>"010101001",
  45709=>"111010010",
  45710=>"000000000",
  45711=>"100110110",
  45712=>"100000010",
  45713=>"101110110",
  45714=>"001001100",
  45715=>"100011000",
  45716=>"111111011",
  45717=>"110111001",
  45718=>"010010110",
  45719=>"000011101",
  45720=>"111000110",
  45721=>"000100100",
  45722=>"000000101",
  45723=>"111100010",
  45724=>"000000100",
  45725=>"010110100",
  45726=>"100010001",
  45727=>"000110101",
  45728=>"011000110",
  45729=>"101111001",
  45730=>"100010010",
  45731=>"000101010",
  45732=>"101001111",
  45733=>"101010001",
  45734=>"000111110",
  45735=>"100011111",
  45736=>"011001100",
  45737=>"111100001",
  45738=>"000011110",
  45739=>"011000000",
  45740=>"001011111",
  45741=>"110110001",
  45742=>"011101001",
  45743=>"010111101",
  45744=>"010000001",
  45745=>"110010000",
  45746=>"000010010",
  45747=>"110001110",
  45748=>"100100111",
  45749=>"001000100",
  45750=>"010011000",
  45751=>"010000010",
  45752=>"011110101",
  45753=>"000000011",
  45754=>"010001110",
  45755=>"011111110",
  45756=>"100001110",
  45757=>"111110100",
  45758=>"111101110",
  45759=>"111110000",
  45760=>"010011111",
  45761=>"001111010",
  45762=>"010100001",
  45763=>"111111111",
  45764=>"101000110",
  45765=>"101001011",
  45766=>"001010010",
  45767=>"101011011",
  45768=>"011000100",
  45769=>"101010101",
  45770=>"101101011",
  45771=>"100111011",
  45772=>"110001011",
  45773=>"001110100",
  45774=>"111011000",
  45775=>"110111110",
  45776=>"111010110",
  45777=>"101010011",
  45778=>"101001011",
  45779=>"010000000",
  45780=>"100100100",
  45781=>"110000001",
  45782=>"011011101",
  45783=>"100000010",
  45784=>"110101010",
  45785=>"101011010",
  45786=>"100001001",
  45787=>"101010001",
  45788=>"001111001",
  45789=>"010010100",
  45790=>"011001010",
  45791=>"110001111",
  45792=>"101000000",
  45793=>"100011100",
  45794=>"001111001",
  45795=>"100110100",
  45796=>"101100001",
  45797=>"101110000",
  45798=>"000101001",
  45799=>"111010010",
  45800=>"001001100",
  45801=>"011010111",
  45802=>"001010110",
  45803=>"000001000",
  45804=>"001100111",
  45805=>"100010011",
  45806=>"111111101",
  45807=>"110001101",
  45808=>"011111101",
  45809=>"000110111",
  45810=>"010000100",
  45811=>"010100011",
  45812=>"111011011",
  45813=>"000011100",
  45814=>"110111000",
  45815=>"010001101",
  45816=>"110010100",
  45817=>"110110110",
  45818=>"011110100",
  45819=>"111000000",
  45820=>"010000101",
  45821=>"100101011",
  45822=>"111001110",
  45823=>"000100011",
  45824=>"011001000",
  45825=>"000111110",
  45826=>"011000111",
  45827=>"111100000",
  45828=>"111111100",
  45829=>"100100100",
  45830=>"011011001",
  45831=>"110101001",
  45832=>"100010011",
  45833=>"010010001",
  45834=>"000111010",
  45835=>"010111111",
  45836=>"000001101",
  45837=>"100000000",
  45838=>"010110001",
  45839=>"111110111",
  45840=>"100101110",
  45841=>"000110000",
  45842=>"011011001",
  45843=>"101010011",
  45844=>"111001101",
  45845=>"100101111",
  45846=>"101011011",
  45847=>"000000000",
  45848=>"010110011",
  45849=>"101011000",
  45850=>"000110010",
  45851=>"101110100",
  45852=>"001100101",
  45853=>"010110110",
  45854=>"101000000",
  45855=>"110110010",
  45856=>"100010100",
  45857=>"001010001",
  45858=>"001101110",
  45859=>"001010111",
  45860=>"110000010",
  45861=>"100111001",
  45862=>"100100110",
  45863=>"100110100",
  45864=>"101100001",
  45865=>"000000001",
  45866=>"100101011",
  45867=>"001101000",
  45868=>"001000001",
  45869=>"110000000",
  45870=>"100011101",
  45871=>"110111001",
  45872=>"010000011",
  45873=>"010100111",
  45874=>"001000100",
  45875=>"000000001",
  45876=>"111101100",
  45877=>"000111101",
  45878=>"001010110",
  45879=>"001101101",
  45880=>"000100100",
  45881=>"010110101",
  45882=>"101011001",
  45883=>"101100100",
  45884=>"011001001",
  45885=>"101100110",
  45886=>"111001000",
  45887=>"010111011",
  45888=>"101000011",
  45889=>"111111110",
  45890=>"000111101",
  45891=>"010101011",
  45892=>"001010111",
  45893=>"001011110",
  45894=>"000101000",
  45895=>"010110110",
  45896=>"111010101",
  45897=>"111101110",
  45898=>"100101001",
  45899=>"111110110",
  45900=>"110000100",
  45901=>"110010010",
  45902=>"011000100",
  45903=>"100111000",
  45904=>"000000001",
  45905=>"110000000",
  45906=>"101110010",
  45907=>"010000111",
  45908=>"011011101",
  45909=>"000100101",
  45910=>"111011011",
  45911=>"110011010",
  45912=>"010011010",
  45913=>"000001000",
  45914=>"100101001",
  45915=>"001100011",
  45916=>"111001011",
  45917=>"011111101",
  45918=>"101000110",
  45919=>"011010011",
  45920=>"000010101",
  45921=>"000111101",
  45922=>"100000111",
  45923=>"011101000",
  45924=>"001110000",
  45925=>"100001100",
  45926=>"101100001",
  45927=>"001101000",
  45928=>"001001000",
  45929=>"100101011",
  45930=>"000100011",
  45931=>"000010101",
  45932=>"100100010",
  45933=>"100111011",
  45934=>"111011011",
  45935=>"101101101",
  45936=>"101000001",
  45937=>"110100000",
  45938=>"011111001",
  45939=>"011000100",
  45940=>"001000110",
  45941=>"001101100",
  45942=>"010111100",
  45943=>"000000111",
  45944=>"110001001",
  45945=>"111100110",
  45946=>"100100001",
  45947=>"100000110",
  45948=>"000000010",
  45949=>"110000011",
  45950=>"111110110",
  45951=>"011000110",
  45952=>"010001001",
  45953=>"111011000",
  45954=>"000100011",
  45955=>"001110001",
  45956=>"111100110",
  45957=>"010101110",
  45958=>"101010001",
  45959=>"111100111",
  45960=>"010011101",
  45961=>"111100000",
  45962=>"101100001",
  45963=>"111010101",
  45964=>"001011011",
  45965=>"100011001",
  45966=>"111010101",
  45967=>"110110001",
  45968=>"001100000",
  45969=>"001011110",
  45970=>"110001101",
  45971=>"001010100",
  45972=>"010111010",
  45973=>"100001111",
  45974=>"010111111",
  45975=>"100111001",
  45976=>"000100111",
  45977=>"110100001",
  45978=>"000110111",
  45979=>"101010110",
  45980=>"001101000",
  45981=>"000011111",
  45982=>"100100000",
  45983=>"001000100",
  45984=>"110111000",
  45985=>"110011111",
  45986=>"100011111",
  45987=>"010111111",
  45988=>"000100110",
  45989=>"100100001",
  45990=>"101101110",
  45991=>"110001010",
  45992=>"110001011",
  45993=>"010000000",
  45994=>"000111001",
  45995=>"101101010",
  45996=>"001001000",
  45997=>"011100001",
  45998=>"000011100",
  45999=>"001100101",
  46000=>"000011110",
  46001=>"100101000",
  46002=>"100010001",
  46003=>"010101000",
  46004=>"100001001",
  46005=>"000100101",
  46006=>"010111110",
  46007=>"111011110",
  46008=>"000101101",
  46009=>"010011010",
  46010=>"010000001",
  46011=>"111011010",
  46012=>"100111011",
  46013=>"110001101",
  46014=>"100100001",
  46015=>"010010001",
  46016=>"000001111",
  46017=>"100001110",
  46018=>"101100101",
  46019=>"010111111",
  46020=>"000111001",
  46021=>"111110000",
  46022=>"101111101",
  46023=>"010010011",
  46024=>"100110111",
  46025=>"101000100",
  46026=>"101010010",
  46027=>"111111111",
  46028=>"001000001",
  46029=>"101101010",
  46030=>"101111101",
  46031=>"100100001",
  46032=>"000001100",
  46033=>"000100100",
  46034=>"010111101",
  46035=>"010001000",
  46036=>"100011011",
  46037=>"000010101",
  46038=>"010000101",
  46039=>"111100110",
  46040=>"101100111",
  46041=>"100110100",
  46042=>"101110010",
  46043=>"000000010",
  46044=>"111000010",
  46045=>"010010100",
  46046=>"001101111",
  46047=>"101010010",
  46048=>"000111101",
  46049=>"001100110",
  46050=>"011011000",
  46051=>"111101100",
  46052=>"101011100",
  46053=>"000000001",
  46054=>"000111111",
  46055=>"010001010",
  46056=>"001010000",
  46057=>"101111101",
  46058=>"010111001",
  46059=>"101001110",
  46060=>"101011001",
  46061=>"001111001",
  46062=>"101100001",
  46063=>"000100010",
  46064=>"011100100",
  46065=>"101100010",
  46066=>"000000001",
  46067=>"100010110",
  46068=>"111001010",
  46069=>"001101000",
  46070=>"100011110",
  46071=>"010111000",
  46072=>"011011000",
  46073=>"011001111",
  46074=>"011101100",
  46075=>"011101001",
  46076=>"110101110",
  46077=>"000001001",
  46078=>"011101011",
  46079=>"101000000",
  46080=>"011000000",
  46081=>"101111011",
  46082=>"101111000",
  46083=>"111111100",
  46084=>"110111001",
  46085=>"011000100",
  46086=>"110001101",
  46087=>"011011111",
  46088=>"111110011",
  46089=>"111101111",
  46090=>"001111001",
  46091=>"100111001",
  46092=>"110001100",
  46093=>"001011001",
  46094=>"101110101",
  46095=>"010100000",
  46096=>"101011110",
  46097=>"111001010",
  46098=>"011010110",
  46099=>"100100110",
  46100=>"101000001",
  46101=>"111000000",
  46102=>"101010011",
  46103=>"110001111",
  46104=>"000000011",
  46105=>"100110110",
  46106=>"110101100",
  46107=>"101100010",
  46108=>"111001010",
  46109=>"100000011",
  46110=>"110000111",
  46111=>"100011110",
  46112=>"101000100",
  46113=>"100101101",
  46114=>"101101111",
  46115=>"101101100",
  46116=>"100001110",
  46117=>"000101101",
  46118=>"110011111",
  46119=>"100100011",
  46120=>"111110011",
  46121=>"100100010",
  46122=>"001010010",
  46123=>"111101001",
  46124=>"001100101",
  46125=>"011111011",
  46126=>"000111110",
  46127=>"000100101",
  46128=>"101100011",
  46129=>"011111011",
  46130=>"000000101",
  46131=>"010110011",
  46132=>"111010111",
  46133=>"010011001",
  46134=>"110110010",
  46135=>"111111001",
  46136=>"001000110",
  46137=>"000011011",
  46138=>"100101111",
  46139=>"111101111",
  46140=>"000100000",
  46141=>"101010011",
  46142=>"110010101",
  46143=>"010100101",
  46144=>"100000110",
  46145=>"011101000",
  46146=>"100010000",
  46147=>"101010101",
  46148=>"110110110",
  46149=>"011011000",
  46150=>"000100100",
  46151=>"101010110",
  46152=>"101001101",
  46153=>"010101110",
  46154=>"001001101",
  46155=>"000101000",
  46156=>"000110001",
  46157=>"011011100",
  46158=>"111010100",
  46159=>"111010111",
  46160=>"011001000",
  46161=>"001011000",
  46162=>"011100000",
  46163=>"001101110",
  46164=>"010100110",
  46165=>"010100010",
  46166=>"111101101",
  46167=>"110110000",
  46168=>"100110000",
  46169=>"110101100",
  46170=>"010110001",
  46171=>"000110111",
  46172=>"000011000",
  46173=>"000111111",
  46174=>"011000000",
  46175=>"101001100",
  46176=>"111100110",
  46177=>"111001100",
  46178=>"111111110",
  46179=>"011110011",
  46180=>"111000010",
  46181=>"100001000",
  46182=>"111111001",
  46183=>"000001100",
  46184=>"100001010",
  46185=>"001011001",
  46186=>"000100100",
  46187=>"100101000",
  46188=>"011010111",
  46189=>"110010000",
  46190=>"001100000",
  46191=>"100001011",
  46192=>"010000010",
  46193=>"101000011",
  46194=>"011010111",
  46195=>"010001000",
  46196=>"111001011",
  46197=>"111010000",
  46198=>"111000000",
  46199=>"001100001",
  46200=>"010011100",
  46201=>"011100000",
  46202=>"010101010",
  46203=>"100101111",
  46204=>"010110011",
  46205=>"011100111",
  46206=>"100101000",
  46207=>"000111001",
  46208=>"010010010",
  46209=>"111000000",
  46210=>"011111110",
  46211=>"111010100",
  46212=>"011000010",
  46213=>"001000011",
  46214=>"110011101",
  46215=>"001000001",
  46216=>"000011101",
  46217=>"001001110",
  46218=>"111011011",
  46219=>"001000010",
  46220=>"000101000",
  46221=>"001110011",
  46222=>"111001000",
  46223=>"111110001",
  46224=>"101101011",
  46225=>"111110011",
  46226=>"101000110",
  46227=>"011001100",
  46228=>"100010101",
  46229=>"100001001",
  46230=>"101110101",
  46231=>"111001011",
  46232=>"000100000",
  46233=>"111001101",
  46234=>"110011110",
  46235=>"011000000",
  46236=>"101110110",
  46237=>"011100100",
  46238=>"111001101",
  46239=>"011001100",
  46240=>"000000101",
  46241=>"000101001",
  46242=>"000101010",
  46243=>"010011100",
  46244=>"001000010",
  46245=>"001011100",
  46246=>"111110101",
  46247=>"100100110",
  46248=>"100011110",
  46249=>"111100010",
  46250=>"111101100",
  46251=>"010111110",
  46252=>"001101011",
  46253=>"010110101",
  46254=>"101101010",
  46255=>"001110000",
  46256=>"000110010",
  46257=>"100000010",
  46258=>"100011100",
  46259=>"110111001",
  46260=>"111100110",
  46261=>"010100101",
  46262=>"001010001",
  46263=>"000111011",
  46264=>"010111000",
  46265=>"101001111",
  46266=>"011100000",
  46267=>"110100011",
  46268=>"001101000",
  46269=>"001101101",
  46270=>"110101101",
  46271=>"111110000",
  46272=>"010101011",
  46273=>"110101011",
  46274=>"111111110",
  46275=>"000110010",
  46276=>"100100110",
  46277=>"011011010",
  46278=>"101111110",
  46279=>"010100100",
  46280=>"100010011",
  46281=>"110000110",
  46282=>"111010001",
  46283=>"100100000",
  46284=>"001111011",
  46285=>"111110110",
  46286=>"101110110",
  46287=>"010010010",
  46288=>"010110101",
  46289=>"011000001",
  46290=>"001011100",
  46291=>"111001100",
  46292=>"010001000",
  46293=>"011011100",
  46294=>"010011000",
  46295=>"101011001",
  46296=>"010111101",
  46297=>"000110010",
  46298=>"010010110",
  46299=>"001110110",
  46300=>"100110111",
  46301=>"111100100",
  46302=>"000101001",
  46303=>"100111001",
  46304=>"110110000",
  46305=>"001011100",
  46306=>"110100001",
  46307=>"010101000",
  46308=>"000100011",
  46309=>"001000111",
  46310=>"110111111",
  46311=>"100110000",
  46312=>"111010001",
  46313=>"110010010",
  46314=>"011101100",
  46315=>"001010001",
  46316=>"000011101",
  46317=>"110111111",
  46318=>"110011101",
  46319=>"010000000",
  46320=>"000111111",
  46321=>"111000000",
  46322=>"000001000",
  46323=>"111101101",
  46324=>"100111001",
  46325=>"100111000",
  46326=>"000010001",
  46327=>"101001111",
  46328=>"101010000",
  46329=>"110011110",
  46330=>"101000110",
  46331=>"110100110",
  46332=>"110011011",
  46333=>"011000000",
  46334=>"000011011",
  46335=>"101101000",
  46336=>"011110010",
  46337=>"101001001",
  46338=>"010110100",
  46339=>"010000111",
  46340=>"101011101",
  46341=>"111110011",
  46342=>"100010100",
  46343=>"110110010",
  46344=>"010001101",
  46345=>"000011101",
  46346=>"111001001",
  46347=>"011010110",
  46348=>"110001101",
  46349=>"011010111",
  46350=>"110101001",
  46351=>"001111101",
  46352=>"010101101",
  46353=>"110100100",
  46354=>"111101111",
  46355=>"111000000",
  46356=>"000011000",
  46357=>"101110011",
  46358=>"000010101",
  46359=>"111001101",
  46360=>"001100011",
  46361=>"101000100",
  46362=>"000110100",
  46363=>"100010010",
  46364=>"001111100",
  46365=>"001010110",
  46366=>"000100100",
  46367=>"001001111",
  46368=>"101110111",
  46369=>"111110110",
  46370=>"011010011",
  46371=>"110101000",
  46372=>"110011100",
  46373=>"000001111",
  46374=>"101100011",
  46375=>"000110101",
  46376=>"010110101",
  46377=>"111010110",
  46378=>"000110100",
  46379=>"110100100",
  46380=>"110110111",
  46381=>"100010010",
  46382=>"000100000",
  46383=>"010110111",
  46384=>"111100110",
  46385=>"011100101",
  46386=>"100011110",
  46387=>"100101100",
  46388=>"011000011",
  46389=>"111100100",
  46390=>"001100111",
  46391=>"111111110",
  46392=>"100111101",
  46393=>"010010010",
  46394=>"000001000",
  46395=>"000010001",
  46396=>"010111100",
  46397=>"000011101",
  46398=>"100011000",
  46399=>"110010000",
  46400=>"001110100",
  46401=>"101111111",
  46402=>"001110000",
  46403=>"101110011",
  46404=>"100000111",
  46405=>"111001111",
  46406=>"000000010",
  46407=>"001010010",
  46408=>"000011011",
  46409=>"011101011",
  46410=>"111101111",
  46411=>"001101111",
  46412=>"101110011",
  46413=>"011000100",
  46414=>"001110001",
  46415=>"101101011",
  46416=>"100000110",
  46417=>"011110101",
  46418=>"100100001",
  46419=>"001011101",
  46420=>"101101011",
  46421=>"010101110",
  46422=>"010101000",
  46423=>"001111000",
  46424=>"110011010",
  46425=>"001011110",
  46426=>"001111101",
  46427=>"111100000",
  46428=>"111010100",
  46429=>"101010111",
  46430=>"100000011",
  46431=>"111111110",
  46432=>"111011110",
  46433=>"011001110",
  46434=>"111011011",
  46435=>"000100001",
  46436=>"101100100",
  46437=>"111101010",
  46438=>"011101010",
  46439=>"000011010",
  46440=>"101100001",
  46441=>"100000100",
  46442=>"000100110",
  46443=>"010011111",
  46444=>"110110010",
  46445=>"000101101",
  46446=>"000000111",
  46447=>"110001101",
  46448=>"000111110",
  46449=>"001110011",
  46450=>"111110101",
  46451=>"111100100",
  46452=>"101010111",
  46453=>"010010100",
  46454=>"100011000",
  46455=>"100101101",
  46456=>"100000101",
  46457=>"101011011",
  46458=>"010000101",
  46459=>"011101000",
  46460=>"011111100",
  46461=>"111101100",
  46462=>"110000101",
  46463=>"101110000",
  46464=>"101011001",
  46465=>"101111000",
  46466=>"000111110",
  46467=>"001001101",
  46468=>"010100100",
  46469=>"000010110",
  46470=>"000101101",
  46471=>"000001100",
  46472=>"011000111",
  46473=>"011101000",
  46474=>"100000101",
  46475=>"101101011",
  46476=>"000000001",
  46477=>"001010101",
  46478=>"000010101",
  46479=>"110101011",
  46480=>"100000000",
  46481=>"111111011",
  46482=>"010100010",
  46483=>"110110100",
  46484=>"001011110",
  46485=>"011101111",
  46486=>"000010000",
  46487=>"000100101",
  46488=>"101110110",
  46489=>"101001000",
  46490=>"111100100",
  46491=>"011000101",
  46492=>"100010011",
  46493=>"100101110",
  46494=>"110011010",
  46495=>"010011110",
  46496=>"110001000",
  46497=>"010000011",
  46498=>"111100101",
  46499=>"000110100",
  46500=>"110111000",
  46501=>"010001000",
  46502=>"101110000",
  46503=>"001010110",
  46504=>"001110110",
  46505=>"100010000",
  46506=>"001110000",
  46507=>"010100001",
  46508=>"001101100",
  46509=>"010011000",
  46510=>"000000101",
  46511=>"110110100",
  46512=>"111010011",
  46513=>"000101001",
  46514=>"010011011",
  46515=>"000101000",
  46516=>"010110001",
  46517=>"101110110",
  46518=>"001000000",
  46519=>"001000001",
  46520=>"000011100",
  46521=>"010100011",
  46522=>"001000110",
  46523=>"001011011",
  46524=>"110000111",
  46525=>"011000110",
  46526=>"111010110",
  46527=>"101010010",
  46528=>"101111111",
  46529=>"110010010",
  46530=>"011101111",
  46531=>"011101100",
  46532=>"110101101",
  46533=>"011011001",
  46534=>"001101101",
  46535=>"111000011",
  46536=>"010001100",
  46537=>"001011100",
  46538=>"000111110",
  46539=>"000010110",
  46540=>"000010111",
  46541=>"110000100",
  46542=>"000100000",
  46543=>"010100111",
  46544=>"101000011",
  46545=>"100100111",
  46546=>"010101110",
  46547=>"101111101",
  46548=>"111101111",
  46549=>"011111101",
  46550=>"111110010",
  46551=>"101001011",
  46552=>"000011100",
  46553=>"101111010",
  46554=>"100110110",
  46555=>"001011101",
  46556=>"010100001",
  46557=>"101011011",
  46558=>"101000001",
  46559=>"001011010",
  46560=>"100101001",
  46561=>"010111110",
  46562=>"001011001",
  46563=>"111001111",
  46564=>"010010111",
  46565=>"010001011",
  46566=>"111111111",
  46567=>"001011000",
  46568=>"001111010",
  46569=>"011010001",
  46570=>"100000100",
  46571=>"011111010",
  46572=>"011111011",
  46573=>"101110101",
  46574=>"011000000",
  46575=>"100100111",
  46576=>"101111101",
  46577=>"101011101",
  46578=>"000000001",
  46579=>"101111111",
  46580=>"111110010",
  46581=>"101110000",
  46582=>"000011111",
  46583=>"001101100",
  46584=>"011110000",
  46585=>"000111010",
  46586=>"101010010",
  46587=>"001111010",
  46588=>"100001010",
  46589=>"001101010",
  46590=>"111100111",
  46591=>"000010011",
  46592=>"101101110",
  46593=>"001011001",
  46594=>"010101001",
  46595=>"110001001",
  46596=>"011011100",
  46597=>"101011101",
  46598=>"010001110",
  46599=>"110100001",
  46600=>"000010011",
  46601=>"000101010",
  46602=>"111111101",
  46603=>"000100000",
  46604=>"110110100",
  46605=>"111100001",
  46606=>"000100001",
  46607=>"100111110",
  46608=>"011101110",
  46609=>"001101101",
  46610=>"100000010",
  46611=>"010101000",
  46612=>"010010101",
  46613=>"000010000",
  46614=>"110010100",
  46615=>"110111110",
  46616=>"001110100",
  46617=>"011110001",
  46618=>"011000011",
  46619=>"001100100",
  46620=>"011000010",
  46621=>"010001100",
  46622=>"011001110",
  46623=>"011011111",
  46624=>"011101101",
  46625=>"100100100",
  46626=>"001100011",
  46627=>"111011100",
  46628=>"111001110",
  46629=>"000010001",
  46630=>"110001111",
  46631=>"100011001",
  46632=>"100111001",
  46633=>"110101010",
  46634=>"011100000",
  46635=>"100001101",
  46636=>"110111100",
  46637=>"101100101",
  46638=>"000001110",
  46639=>"000001010",
  46640=>"101001000",
  46641=>"110011101",
  46642=>"010000101",
  46643=>"001101000",
  46644=>"110101011",
  46645=>"000001011",
  46646=>"000110011",
  46647=>"000011111",
  46648=>"010001010",
  46649=>"001000000",
  46650=>"010011000",
  46651=>"100110000",
  46652=>"100010111",
  46653=>"011000101",
  46654=>"001001011",
  46655=>"101000101",
  46656=>"101110010",
  46657=>"100011111",
  46658=>"111000110",
  46659=>"101101010",
  46660=>"000101000",
  46661=>"010011110",
  46662=>"011010101",
  46663=>"100011001",
  46664=>"001011010",
  46665=>"010111010",
  46666=>"010010010",
  46667=>"000101100",
  46668=>"111110101",
  46669=>"111101001",
  46670=>"110111011",
  46671=>"010000001",
  46672=>"111010101",
  46673=>"111100010",
  46674=>"101000100",
  46675=>"011100000",
  46676=>"001110010",
  46677=>"110100110",
  46678=>"100000110",
  46679=>"000011101",
  46680=>"110011001",
  46681=>"000101000",
  46682=>"000100011",
  46683=>"000100111",
  46684=>"110101010",
  46685=>"101111101",
  46686=>"000111000",
  46687=>"001111000",
  46688=>"010000101",
  46689=>"000000101",
  46690=>"100010000",
  46691=>"111010011",
  46692=>"101011010",
  46693=>"100101001",
  46694=>"001000101",
  46695=>"010100011",
  46696=>"001000100",
  46697=>"001101010",
  46698=>"110010000",
  46699=>"110110101",
  46700=>"000000111",
  46701=>"000011100",
  46702=>"100011001",
  46703=>"101000001",
  46704=>"111101111",
  46705=>"001100110",
  46706=>"110010010",
  46707=>"101001011",
  46708=>"100110101",
  46709=>"010011001",
  46710=>"100000010",
  46711=>"110000101",
  46712=>"101001101",
  46713=>"111000010",
  46714=>"011111111",
  46715=>"100100011",
  46716=>"000001000",
  46717=>"001101010",
  46718=>"101101001",
  46719=>"111000110",
  46720=>"010001010",
  46721=>"100111110",
  46722=>"111101010",
  46723=>"101011101",
  46724=>"011101101",
  46725=>"000011101",
  46726=>"000001000",
  46727=>"111100111",
  46728=>"001100010",
  46729=>"110100011",
  46730=>"111001111",
  46731=>"011101101",
  46732=>"000010100",
  46733=>"001100111",
  46734=>"111011101",
  46735=>"100000100",
  46736=>"111000001",
  46737=>"110101001",
  46738=>"101110100",
  46739=>"111110111",
  46740=>"000111001",
  46741=>"010110000",
  46742=>"110111010",
  46743=>"100100100",
  46744=>"010010111",
  46745=>"101100101",
  46746=>"000100011",
  46747=>"100111101",
  46748=>"100000000",
  46749=>"000001011",
  46750=>"111100011",
  46751=>"111100001",
  46752=>"000010001",
  46753=>"111100000",
  46754=>"101001001",
  46755=>"110111111",
  46756=>"100100010",
  46757=>"101011100",
  46758=>"000011000",
  46759=>"111111001",
  46760=>"011000001",
  46761=>"001001001",
  46762=>"011110100",
  46763=>"001000011",
  46764=>"100101000",
  46765=>"011001101",
  46766=>"111010000",
  46767=>"101011101",
  46768=>"010101110",
  46769=>"100001011",
  46770=>"001111001",
  46771=>"110100101",
  46772=>"100111100",
  46773=>"101000001",
  46774=>"010110001",
  46775=>"010100000",
  46776=>"100110101",
  46777=>"001100101",
  46778=>"000110111",
  46779=>"010010111",
  46780=>"101100111",
  46781=>"101110101",
  46782=>"111010000",
  46783=>"111110101",
  46784=>"110011010",
  46785=>"000000110",
  46786=>"111100111",
  46787=>"100101001",
  46788=>"000010111",
  46789=>"000011100",
  46790=>"111111110",
  46791=>"000111101",
  46792=>"110011101",
  46793=>"110101111",
  46794=>"111100110",
  46795=>"110000110",
  46796=>"110101101",
  46797=>"011100110",
  46798=>"111110011",
  46799=>"010011010",
  46800=>"010001010",
  46801=>"111001100",
  46802=>"110011100",
  46803=>"100101111",
  46804=>"101100101",
  46805=>"011010111",
  46806=>"101110111",
  46807=>"100000000",
  46808=>"001111101",
  46809=>"010110000",
  46810=>"001110001",
  46811=>"100001000",
  46812=>"011100011",
  46813=>"100101100",
  46814=>"011010010",
  46815=>"101111011",
  46816=>"111101111",
  46817=>"110111110",
  46818=>"110011010",
  46819=>"101110010",
  46820=>"000111011",
  46821=>"110000011",
  46822=>"110111111",
  46823=>"100001101",
  46824=>"101000000",
  46825=>"110000101",
  46826=>"111011101",
  46827=>"000010010",
  46828=>"000111110",
  46829=>"110110010",
  46830=>"011011000",
  46831=>"101100001",
  46832=>"000010111",
  46833=>"011000100",
  46834=>"010001000",
  46835=>"000100010",
  46836=>"101001010",
  46837=>"010010010",
  46838=>"110010111",
  46839=>"010001001",
  46840=>"011010110",
  46841=>"100100000",
  46842=>"011111000",
  46843=>"010111001",
  46844=>"010111001",
  46845=>"000000011",
  46846=>"110111011",
  46847=>"001011000",
  46848=>"110111101",
  46849=>"101101011",
  46850=>"001110001",
  46851=>"000000010",
  46852=>"111111111",
  46853=>"011001111",
  46854=>"101111000",
  46855=>"010001001",
  46856=>"000101101",
  46857=>"011001101",
  46858=>"101100101",
  46859=>"111100011",
  46860=>"101000111",
  46861=>"111110000",
  46862=>"001101111",
  46863=>"011110000",
  46864=>"110110001",
  46865=>"111111111",
  46866=>"100010001",
  46867=>"011111011",
  46868=>"001011111",
  46869=>"111010001",
  46870=>"100011010",
  46871=>"111001011",
  46872=>"000011101",
  46873=>"110011100",
  46874=>"000101110",
  46875=>"101110110",
  46876=>"100101111",
  46877=>"101011011",
  46878=>"000001110",
  46879=>"010110100",
  46880=>"100001000",
  46881=>"011110011",
  46882=>"011110000",
  46883=>"101111111",
  46884=>"111100101",
  46885=>"000110011",
  46886=>"100110000",
  46887=>"101111111",
  46888=>"001110010",
  46889=>"110111110",
  46890=>"111111101",
  46891=>"000101100",
  46892=>"100001010",
  46893=>"110101000",
  46894=>"111001010",
  46895=>"100000000",
  46896=>"000000010",
  46897=>"101100110",
  46898=>"110111000",
  46899=>"010101010",
  46900=>"110100000",
  46901=>"111001100",
  46902=>"111100001",
  46903=>"010011010",
  46904=>"000100100",
  46905=>"001011001",
  46906=>"000100000",
  46907=>"011001111",
  46908=>"110011100",
  46909=>"100111101",
  46910=>"010000010",
  46911=>"101111110",
  46912=>"010001000",
  46913=>"001000111",
  46914=>"000011010",
  46915=>"000110001",
  46916=>"011011110",
  46917=>"001101001",
  46918=>"101000101",
  46919=>"111011000",
  46920=>"100000101",
  46921=>"100100011",
  46922=>"110111111",
  46923=>"010010111",
  46924=>"011110111",
  46925=>"001110101",
  46926=>"101101110",
  46927=>"001010110",
  46928=>"111000100",
  46929=>"010010101",
  46930=>"000111010",
  46931=>"111010001",
  46932=>"000001111",
  46933=>"000110011",
  46934=>"010010010",
  46935=>"110100101",
  46936=>"110100110",
  46937=>"001000110",
  46938=>"100101011",
  46939=>"010000000",
  46940=>"100110100",
  46941=>"110010010",
  46942=>"010000101",
  46943=>"100100111",
  46944=>"001111100",
  46945=>"110101110",
  46946=>"100011111",
  46947=>"000010000",
  46948=>"111000010",
  46949=>"001011101",
  46950=>"010011110",
  46951=>"010100011",
  46952=>"111001000",
  46953=>"001101010",
  46954=>"101010101",
  46955=>"111110001",
  46956=>"001111011",
  46957=>"110011100",
  46958=>"011011111",
  46959=>"011110101",
  46960=>"111011001",
  46961=>"101011111",
  46962=>"110111011",
  46963=>"000001000",
  46964=>"100010011",
  46965=>"011110100",
  46966=>"101110100",
  46967=>"010100000",
  46968=>"110100011",
  46969=>"001000001",
  46970=>"000011101",
  46971=>"101011001",
  46972=>"000000000",
  46973=>"011000011",
  46974=>"000101101",
  46975=>"110001001",
  46976=>"000010111",
  46977=>"100101000",
  46978=>"100010000",
  46979=>"111010001",
  46980=>"100001110",
  46981=>"100111001",
  46982=>"110111101",
  46983=>"001000010",
  46984=>"110010110",
  46985=>"001110100",
  46986=>"110001010",
  46987=>"111100010",
  46988=>"101111001",
  46989=>"010011101",
  46990=>"011001000",
  46991=>"100010100",
  46992=>"101111100",
  46993=>"110100000",
  46994=>"100001001",
  46995=>"100001011",
  46996=>"110011110",
  46997=>"101011100",
  46998=>"100001111",
  46999=>"011001010",
  47000=>"001011111",
  47001=>"111100000",
  47002=>"111111111",
  47003=>"110000010",
  47004=>"100101111",
  47005=>"010110001",
  47006=>"100001010",
  47007=>"001100100",
  47008=>"111101110",
  47009=>"011111110",
  47010=>"111100011",
  47011=>"011001111",
  47012=>"010010000",
  47013=>"110001110",
  47014=>"100001000",
  47015=>"100010110",
  47016=>"110010011",
  47017=>"100000011",
  47018=>"010001110",
  47019=>"100011011",
  47020=>"110011010",
  47021=>"101101100",
  47022=>"111010011",
  47023=>"010110000",
  47024=>"000000010",
  47025=>"011010011",
  47026=>"001101000",
  47027=>"101101111",
  47028=>"110011100",
  47029=>"000101001",
  47030=>"011000110",
  47031=>"000101001",
  47032=>"100001101",
  47033=>"010011101",
  47034=>"011010010",
  47035=>"001010011",
  47036=>"111110110",
  47037=>"010011111",
  47038=>"111001000",
  47039=>"010010101",
  47040=>"101111010",
  47041=>"011101111",
  47042=>"010100010",
  47043=>"011011100",
  47044=>"110101110",
  47045=>"101001100",
  47046=>"001110011",
  47047=>"111011011",
  47048=>"000010101",
  47049=>"001101100",
  47050=>"000101111",
  47051=>"000001101",
  47052=>"100010011",
  47053=>"001100110",
  47054=>"001111110",
  47055=>"100110110",
  47056=>"011010101",
  47057=>"000101010",
  47058=>"010010100",
  47059=>"101100000",
  47060=>"100000101",
  47061=>"111110001",
  47062=>"010111010",
  47063=>"101100010",
  47064=>"010101001",
  47065=>"111111111",
  47066=>"110110110",
  47067=>"000001000",
  47068=>"111010000",
  47069=>"001110000",
  47070=>"101000000",
  47071=>"001001010",
  47072=>"101001011",
  47073=>"000100001",
  47074=>"111010101",
  47075=>"001111101",
  47076=>"000000000",
  47077=>"111010011",
  47078=>"000011100",
  47079=>"100111010",
  47080=>"000111000",
  47081=>"001001010",
  47082=>"011001111",
  47083=>"001111001",
  47084=>"001011100",
  47085=>"010111100",
  47086=>"010100000",
  47087=>"000001111",
  47088=>"101100101",
  47089=>"111101100",
  47090=>"000010110",
  47091=>"111001000",
  47092=>"001011111",
  47093=>"111110100",
  47094=>"010010110",
  47095=>"011100100",
  47096=>"001010100",
  47097=>"000110011",
  47098=>"010101101",
  47099=>"111000101",
  47100=>"100111011",
  47101=>"010000101",
  47102=>"010010010",
  47103=>"011000111",
  47104=>"111000101",
  47105=>"101111111",
  47106=>"011110001",
  47107=>"111100001",
  47108=>"111011001",
  47109=>"010111101",
  47110=>"101111001",
  47111=>"110001111",
  47112=>"110111111",
  47113=>"101000010",
  47114=>"111101100",
  47115=>"101000110",
  47116=>"101110100",
  47117=>"010010100",
  47118=>"101111000",
  47119=>"100101100",
  47120=>"011100101",
  47121=>"110010101",
  47122=>"110101100",
  47123=>"000100110",
  47124=>"010100110",
  47125=>"001000001",
  47126=>"111011010",
  47127=>"010111011",
  47128=>"111111001",
  47129=>"101000100",
  47130=>"110000011",
  47131=>"101110010",
  47132=>"100111011",
  47133=>"110111011",
  47134=>"010011110",
  47135=>"011011100",
  47136=>"010001111",
  47137=>"000100001",
  47138=>"100000010",
  47139=>"101010000",
  47140=>"110110011",
  47141=>"000010100",
  47142=>"001000100",
  47143=>"001011111",
  47144=>"110010010",
  47145=>"000110100",
  47146=>"011110101",
  47147=>"110011101",
  47148=>"110101001",
  47149=>"011101110",
  47150=>"011101111",
  47151=>"101000101",
  47152=>"101010111",
  47153=>"010110111",
  47154=>"101101100",
  47155=>"010110010",
  47156=>"100111101",
  47157=>"010111011",
  47158=>"000010101",
  47159=>"000100111",
  47160=>"100111101",
  47161=>"000100111",
  47162=>"110111101",
  47163=>"000111011",
  47164=>"000100101",
  47165=>"011001011",
  47166=>"110000000",
  47167=>"111111110",
  47168=>"001110010",
  47169=>"001011000",
  47170=>"011110001",
  47171=>"001101000",
  47172=>"110000100",
  47173=>"110111110",
  47174=>"110111011",
  47175=>"010011110",
  47176=>"101111011",
  47177=>"101100110",
  47178=>"001001010",
  47179=>"001000100",
  47180=>"001001110",
  47181=>"111000100",
  47182=>"110111111",
  47183=>"000011101",
  47184=>"110111100",
  47185=>"110000001",
  47186=>"011010100",
  47187=>"010110010",
  47188=>"011111111",
  47189=>"001111111",
  47190=>"001111000",
  47191=>"010100001",
  47192=>"101100101",
  47193=>"001011111",
  47194=>"111101101",
  47195=>"110010101",
  47196=>"001100010",
  47197=>"011101101",
  47198=>"000010011",
  47199=>"110110011",
  47200=>"010000110",
  47201=>"010010101",
  47202=>"100100110",
  47203=>"101110001",
  47204=>"001000111",
  47205=>"101100111",
  47206=>"010011101",
  47207=>"001011110",
  47208=>"111100111",
  47209=>"110011101",
  47210=>"001110011",
  47211=>"101000110",
  47212=>"010110100",
  47213=>"110010011",
  47214=>"111010010",
  47215=>"010011000",
  47216=>"011010010",
  47217=>"101111001",
  47218=>"001010100",
  47219=>"101000101",
  47220=>"110000110",
  47221=>"111000001",
  47222=>"100110111",
  47223=>"100001100",
  47224=>"100000110",
  47225=>"111000011",
  47226=>"111100101",
  47227=>"111010010",
  47228=>"001101011",
  47229=>"001000011",
  47230=>"111101110",
  47231=>"001110101",
  47232=>"010101101",
  47233=>"101111010",
  47234=>"010010000",
  47235=>"101101001",
  47236=>"110110100",
  47237=>"011111111",
  47238=>"000100111",
  47239=>"011011010",
  47240=>"000111100",
  47241=>"010001001",
  47242=>"001001101",
  47243=>"111101001",
  47244=>"110000101",
  47245=>"010000001",
  47246=>"100111010",
  47247=>"110010100",
  47248=>"011000011",
  47249=>"011011001",
  47250=>"000010011",
  47251=>"111001010",
  47252=>"111001101",
  47253=>"000011010",
  47254=>"100001000",
  47255=>"011001101",
  47256=>"010011010",
  47257=>"110101110",
  47258=>"101000100",
  47259=>"101010011",
  47260=>"011000101",
  47261=>"000001001",
  47262=>"000100011",
  47263=>"100101001",
  47264=>"100000101",
  47265=>"001011000",
  47266=>"110100110",
  47267=>"101111100",
  47268=>"000111010",
  47269=>"001110111",
  47270=>"100010110",
  47271=>"101111000",
  47272=>"110010101",
  47273=>"000101001",
  47274=>"100111010",
  47275=>"110011001",
  47276=>"110001101",
  47277=>"001010001",
  47278=>"011110100",
  47279=>"110000100",
  47280=>"000110100",
  47281=>"110010101",
  47282=>"001010100",
  47283=>"101000001",
  47284=>"111101010",
  47285=>"011101111",
  47286=>"000110111",
  47287=>"001001010",
  47288=>"001111101",
  47289=>"100011011",
  47290=>"000011101",
  47291=>"001010011",
  47292=>"000111010",
  47293=>"110001111",
  47294=>"100111101",
  47295=>"110111010",
  47296=>"111111100",
  47297=>"001110011",
  47298=>"000111101",
  47299=>"000000011",
  47300=>"010010000",
  47301=>"011111110",
  47302=>"111000010",
  47303=>"010001001",
  47304=>"110110001",
  47305=>"101000000",
  47306=>"101111111",
  47307=>"000011001",
  47308=>"011010100",
  47309=>"001110101",
  47310=>"010100010",
  47311=>"010000011",
  47312=>"111010101",
  47313=>"111011110",
  47314=>"000000001",
  47315=>"110001001",
  47316=>"000111101",
  47317=>"011011111",
  47318=>"000110000",
  47319=>"001111001",
  47320=>"111101010",
  47321=>"100001101",
  47322=>"111000001",
  47323=>"000101100",
  47324=>"011111000",
  47325=>"101001001",
  47326=>"001011001",
  47327=>"001011110",
  47328=>"110010000",
  47329=>"111100001",
  47330=>"010010101",
  47331=>"000000101",
  47332=>"000001001",
  47333=>"110001101",
  47334=>"111101001",
  47335=>"000000011",
  47336=>"110101111",
  47337=>"000110110",
  47338=>"111111111",
  47339=>"010110101",
  47340=>"101101101",
  47341=>"000011000",
  47342=>"100101001",
  47343=>"100110011",
  47344=>"010110000",
  47345=>"100001101",
  47346=>"011000001",
  47347=>"011110010",
  47348=>"000011101",
  47349=>"011100101",
  47350=>"101110100",
  47351=>"000010000",
  47352=>"110110110",
  47353=>"110001000",
  47354=>"000101100",
  47355=>"010010110",
  47356=>"111010101",
  47357=>"000101011",
  47358=>"010111000",
  47359=>"011011001",
  47360=>"001010100",
  47361=>"110011101",
  47362=>"000110101",
  47363=>"000010111",
  47364=>"010000111",
  47365=>"100011000",
  47366=>"101110110",
  47367=>"110101010",
  47368=>"001010011",
  47369=>"100010000",
  47370=>"100101111",
  47371=>"100001101",
  47372=>"000100111",
  47373=>"010010110",
  47374=>"010010111",
  47375=>"001010011",
  47376=>"000011001",
  47377=>"100110010",
  47378=>"111110100",
  47379=>"001111101",
  47380=>"111000101",
  47381=>"001010000",
  47382=>"000001100",
  47383=>"110010000",
  47384=>"000000111",
  47385=>"010001110",
  47386=>"110010101",
  47387=>"101110100",
  47388=>"111010111",
  47389=>"011001100",
  47390=>"110101110",
  47391=>"111011000",
  47392=>"011111101",
  47393=>"001110011",
  47394=>"110110010",
  47395=>"000010111",
  47396=>"110000010",
  47397=>"110011100",
  47398=>"100111001",
  47399=>"000001110",
  47400=>"111011010",
  47401=>"000000101",
  47402=>"011110001",
  47403=>"010010111",
  47404=>"101100010",
  47405=>"000011101",
  47406=>"000110011",
  47407=>"111111001",
  47408=>"010011101",
  47409=>"100001001",
  47410=>"000000000",
  47411=>"110110010",
  47412=>"100010101",
  47413=>"000001111",
  47414=>"010011101",
  47415=>"000000000",
  47416=>"100111111",
  47417=>"000100111",
  47418=>"111011100",
  47419=>"100001111",
  47420=>"110110001",
  47421=>"001011000",
  47422=>"010011110",
  47423=>"110001000",
  47424=>"111101001",
  47425=>"111000010",
  47426=>"100101100",
  47427=>"111001011",
  47428=>"100100110",
  47429=>"101110000",
  47430=>"101000011",
  47431=>"000001000",
  47432=>"101101100",
  47433=>"100001100",
  47434=>"010100011",
  47435=>"001010110",
  47436=>"000000000",
  47437=>"101101001",
  47438=>"111011100",
  47439=>"110001111",
  47440=>"110011011",
  47441=>"101111010",
  47442=>"100000100",
  47443=>"111011101",
  47444=>"100110100",
  47445=>"011111100",
  47446=>"111000011",
  47447=>"101000110",
  47448=>"000010001",
  47449=>"011011110",
  47450=>"101110110",
  47451=>"000001110",
  47452=>"110110101",
  47453=>"111111111",
  47454=>"100000010",
  47455=>"101001001",
  47456=>"100011011",
  47457=>"100101101",
  47458=>"101101111",
  47459=>"010000011",
  47460=>"011111110",
  47461=>"011000110",
  47462=>"101111100",
  47463=>"111111011",
  47464=>"011000010",
  47465=>"011100111",
  47466=>"011010000",
  47467=>"111110000",
  47468=>"000100101",
  47469=>"111100110",
  47470=>"110111100",
  47471=>"110010011",
  47472=>"101100010",
  47473=>"110001000",
  47474=>"011010100",
  47475=>"011111100",
  47476=>"010110111",
  47477=>"001101000",
  47478=>"001000101",
  47479=>"100001001",
  47480=>"010001111",
  47481=>"100101010",
  47482=>"111011010",
  47483=>"010110010",
  47484=>"000100000",
  47485=>"110000111",
  47486=>"101101100",
  47487=>"011010111",
  47488=>"010010111",
  47489=>"000000011",
  47490=>"010111010",
  47491=>"100010001",
  47492=>"101011101",
  47493=>"010100110",
  47494=>"101111001",
  47495=>"000010001",
  47496=>"010010010",
  47497=>"101111011",
  47498=>"010001000",
  47499=>"001111110",
  47500=>"011010011",
  47501=>"001111111",
  47502=>"000111000",
  47503=>"100101011",
  47504=>"111011110",
  47505=>"110010110",
  47506=>"011011101",
  47507=>"011010100",
  47508=>"011110100",
  47509=>"011011100",
  47510=>"001010110",
  47511=>"000000111",
  47512=>"011001001",
  47513=>"001110011",
  47514=>"111101101",
  47515=>"101000011",
  47516=>"100100100",
  47517=>"110000110",
  47518=>"111110010",
  47519=>"100111010",
  47520=>"000001110",
  47521=>"010101110",
  47522=>"000100010",
  47523=>"101110011",
  47524=>"001010001",
  47525=>"000011011",
  47526=>"100110110",
  47527=>"100001010",
  47528=>"010011101",
  47529=>"011011101",
  47530=>"001101110",
  47531=>"001111101",
  47532=>"111111110",
  47533=>"000111001",
  47534=>"010011001",
  47535=>"111110100",
  47536=>"010000100",
  47537=>"110010001",
  47538=>"101101000",
  47539=>"011010001",
  47540=>"111000010",
  47541=>"111010101",
  47542=>"011110001",
  47543=>"010100110",
  47544=>"110110111",
  47545=>"110001111",
  47546=>"001000001",
  47547=>"000111100",
  47548=>"011111011",
  47549=>"010111000",
  47550=>"101111111",
  47551=>"101101100",
  47552=>"010110000",
  47553=>"110101100",
  47554=>"111111110",
  47555=>"101000011",
  47556=>"011111100",
  47557=>"010100000",
  47558=>"000010111",
  47559=>"100010000",
  47560=>"001010111",
  47561=>"111010011",
  47562=>"110011011",
  47563=>"100011111",
  47564=>"000101111",
  47565=>"101100010",
  47566=>"001110011",
  47567=>"010110011",
  47568=>"011111000",
  47569=>"101000101",
  47570=>"111011010",
  47571=>"010111000",
  47572=>"010011110",
  47573=>"010010010",
  47574=>"111010110",
  47575=>"001011010",
  47576=>"101111011",
  47577=>"111111111",
  47578=>"100001110",
  47579=>"100000101",
  47580=>"001101110",
  47581=>"010101000",
  47582=>"100010000",
  47583=>"110101010",
  47584=>"010010111",
  47585=>"010111011",
  47586=>"001101010",
  47587=>"101100110",
  47588=>"010000111",
  47589=>"111000010",
  47590=>"000010111",
  47591=>"110101110",
  47592=>"101101100",
  47593=>"110000010",
  47594=>"100010110",
  47595=>"110111111",
  47596=>"101010001",
  47597=>"101100000",
  47598=>"011001101",
  47599=>"000110110",
  47600=>"000011111",
  47601=>"111010000",
  47602=>"111001111",
  47603=>"010011100",
  47604=>"110111010",
  47605=>"010110101",
  47606=>"010111001",
  47607=>"011111101",
  47608=>"000000100",
  47609=>"010111111",
  47610=>"101001110",
  47611=>"110001100",
  47612=>"100101011",
  47613=>"011101101",
  47614=>"100100000",
  47615=>"111111010",
  47616=>"010110000",
  47617=>"011100000",
  47618=>"000000001",
  47619=>"011110011",
  47620=>"001111000",
  47621=>"001110001",
  47622=>"100000110",
  47623=>"011100111",
  47624=>"110001110",
  47625=>"000000001",
  47626=>"001101110",
  47627=>"111100001",
  47628=>"001101010",
  47629=>"100110111",
  47630=>"010111001",
  47631=>"110101000",
  47632=>"001000111",
  47633=>"010100010",
  47634=>"101100011",
  47635=>"101101110",
  47636=>"111110011",
  47637=>"111101001",
  47638=>"111001101",
  47639=>"100100111",
  47640=>"000110101",
  47641=>"010001111",
  47642=>"000000110",
  47643=>"110110000",
  47644=>"000010011",
  47645=>"110101101",
  47646=>"011010001",
  47647=>"101111110",
  47648=>"110001100",
  47649=>"000000111",
  47650=>"000010111",
  47651=>"000011010",
  47652=>"000010110",
  47653=>"010100001",
  47654=>"111111001",
  47655=>"110011001",
  47656=>"111010010",
  47657=>"010000000",
  47658=>"101000100",
  47659=>"110000101",
  47660=>"011011101",
  47661=>"001000111",
  47662=>"100100010",
  47663=>"011010100",
  47664=>"000001111",
  47665=>"000000101",
  47666=>"100010111",
  47667=>"100110010",
  47668=>"110010000",
  47669=>"000001100",
  47670=>"001110010",
  47671=>"001111001",
  47672=>"000101011",
  47673=>"000100000",
  47674=>"100110110",
  47675=>"000001001",
  47676=>"100111101",
  47677=>"010000000",
  47678=>"011001111",
  47679=>"111010111",
  47680=>"100000011",
  47681=>"010011111",
  47682=>"010000011",
  47683=>"010001010",
  47684=>"100101111",
  47685=>"111110100",
  47686=>"101110111",
  47687=>"000101101",
  47688=>"111010110",
  47689=>"110001110",
  47690=>"010000111",
  47691=>"011011110",
  47692=>"000001100",
  47693=>"000011110",
  47694=>"110100011",
  47695=>"111010010",
  47696=>"001010101",
  47697=>"111110101",
  47698=>"110110111",
  47699=>"101000000",
  47700=>"010000100",
  47701=>"010010111",
  47702=>"001101111",
  47703=>"100101011",
  47704=>"111111111",
  47705=>"100100001",
  47706=>"110110111",
  47707=>"010101011",
  47708=>"100000001",
  47709=>"000110001",
  47710=>"010001011",
  47711=>"000011111",
  47712=>"111000110",
  47713=>"000100110",
  47714=>"101111111",
  47715=>"000000010",
  47716=>"011011111",
  47717=>"111111101",
  47718=>"111100001",
  47719=>"001111011",
  47720=>"100111010",
  47721=>"000000010",
  47722=>"110101001",
  47723=>"100000100",
  47724=>"000011100",
  47725=>"111011011",
  47726=>"100101001",
  47727=>"001110011",
  47728=>"100100100",
  47729=>"001000000",
  47730=>"001111110",
  47731=>"111100000",
  47732=>"110111101",
  47733=>"011010111",
  47734=>"010111101",
  47735=>"010110101",
  47736=>"101000010",
  47737=>"001110100",
  47738=>"111100101",
  47739=>"010100001",
  47740=>"111011001",
  47741=>"000100010",
  47742=>"011110000",
  47743=>"101000000",
  47744=>"001110101",
  47745=>"100010111",
  47746=>"011110110",
  47747=>"010001011",
  47748=>"010011001",
  47749=>"010000100",
  47750=>"100000110",
  47751=>"110001100",
  47752=>"011100111",
  47753=>"001001100",
  47754=>"000011101",
  47755=>"011111000",
  47756=>"111010000",
  47757=>"011011001",
  47758=>"011110100",
  47759=>"011100101",
  47760=>"001111101",
  47761=>"111001010",
  47762=>"110101011",
  47763=>"110000001",
  47764=>"110001001",
  47765=>"111111111",
  47766=>"111100010",
  47767=>"000101100",
  47768=>"111100010",
  47769=>"111000001",
  47770=>"001001101",
  47771=>"101010100",
  47772=>"100001111",
  47773=>"011001110",
  47774=>"110101000",
  47775=>"000001100",
  47776=>"101001101",
  47777=>"101011110",
  47778=>"111011101",
  47779=>"010000001",
  47780=>"101100000",
  47781=>"011111011",
  47782=>"101101110",
  47783=>"000011001",
  47784=>"111110101",
  47785=>"001101111",
  47786=>"010010110",
  47787=>"101010010",
  47788=>"000011000",
  47789=>"011101101",
  47790=>"000111010",
  47791=>"110101010",
  47792=>"111100110",
  47793=>"101010101",
  47794=>"011101011",
  47795=>"011110111",
  47796=>"110101111",
  47797=>"011001101",
  47798=>"001010100",
  47799=>"001100110",
  47800=>"101011011",
  47801=>"111011110",
  47802=>"001010011",
  47803=>"001111011",
  47804=>"101011011",
  47805=>"010001011",
  47806=>"010111001",
  47807=>"011011100",
  47808=>"000000110",
  47809=>"101100100",
  47810=>"001011101",
  47811=>"111100011",
  47812=>"011001110",
  47813=>"010001111",
  47814=>"111001100",
  47815=>"001100111",
  47816=>"000000111",
  47817=>"010000000",
  47818=>"000011100",
  47819=>"111001110",
  47820=>"001110011",
  47821=>"001100001",
  47822=>"011111001",
  47823=>"000000010",
  47824=>"011001110",
  47825=>"100000011",
  47826=>"100101001",
  47827=>"111100101",
  47828=>"111111100",
  47829=>"100100010",
  47830=>"011001101",
  47831=>"011101001",
  47832=>"101010010",
  47833=>"110100111",
  47834=>"101001000",
  47835=>"101101001",
  47836=>"100000110",
  47837=>"111110110",
  47838=>"011110110",
  47839=>"001010100",
  47840=>"100001000",
  47841=>"110000100",
  47842=>"111001101",
  47843=>"111110101",
  47844=>"100000000",
  47845=>"100100000",
  47846=>"100010111",
  47847=>"110111010",
  47848=>"001100010",
  47849=>"001111101",
  47850=>"000001010",
  47851=>"011101110",
  47852=>"100111101",
  47853=>"000110110",
  47854=>"101011101",
  47855=>"111101101",
  47856=>"010000010",
  47857=>"111010001",
  47858=>"111110011",
  47859=>"000011000",
  47860=>"111011000",
  47861=>"001101110",
  47862=>"011110011",
  47863=>"000000001",
  47864=>"101000100",
  47865=>"010001100",
  47866=>"000100000",
  47867=>"001101100",
  47868=>"111011101",
  47869=>"000000101",
  47870=>"101000100",
  47871=>"111101111",
  47872=>"001001011",
  47873=>"111000010",
  47874=>"101011111",
  47875=>"110000100",
  47876=>"011011110",
  47877=>"001010001",
  47878=>"101110011",
  47879=>"110101101",
  47880=>"000001111",
  47881=>"111100101",
  47882=>"001111011",
  47883=>"000100011",
  47884=>"000100101",
  47885=>"111100100",
  47886=>"001001010",
  47887=>"001001010",
  47888=>"010110111",
  47889=>"101111010",
  47890=>"010000100",
  47891=>"110011110",
  47892=>"101000011",
  47893=>"000110110",
  47894=>"110101111",
  47895=>"000011101",
  47896=>"011111010",
  47897=>"000010110",
  47898=>"110000100",
  47899=>"101000100",
  47900=>"101001110",
  47901=>"110001101",
  47902=>"100000111",
  47903=>"011011010",
  47904=>"110001011",
  47905=>"110110011",
  47906=>"111110001",
  47907=>"001100111",
  47908=>"010011011",
  47909=>"011000000",
  47910=>"111011111",
  47911=>"100001000",
  47912=>"011101010",
  47913=>"100001111",
  47914=>"111010110",
  47915=>"001000011",
  47916=>"101101100",
  47917=>"001010101",
  47918=>"111011010",
  47919=>"111010110",
  47920=>"001011011",
  47921=>"110111001",
  47922=>"000011011",
  47923=>"110110100",
  47924=>"110001101",
  47925=>"101011100",
  47926=>"000111010",
  47927=>"001000101",
  47928=>"101000111",
  47929=>"011100100",
  47930=>"001111101",
  47931=>"100110001",
  47932=>"111100111",
  47933=>"100111110",
  47934=>"000101111",
  47935=>"101111011",
  47936=>"110111010",
  47937=>"101111011",
  47938=>"111111001",
  47939=>"100010111",
  47940=>"010001101",
  47941=>"111000101",
  47942=>"100000000",
  47943=>"011011100",
  47944=>"110100010",
  47945=>"110101111",
  47946=>"000001011",
  47947=>"110000110",
  47948=>"100011100",
  47949=>"000000011",
  47950=>"011010011",
  47951=>"001111101",
  47952=>"110010011",
  47953=>"100010010",
  47954=>"011010000",
  47955=>"000101011",
  47956=>"001011100",
  47957=>"101111111",
  47958=>"101011010",
  47959=>"010100000",
  47960=>"000101010",
  47961=>"010110111",
  47962=>"001000001",
  47963=>"100110000",
  47964=>"100001011",
  47965=>"000111011",
  47966=>"101011000",
  47967=>"011100010",
  47968=>"010101000",
  47969=>"001000011",
  47970=>"000110100",
  47971=>"110010011",
  47972=>"001001011",
  47973=>"000000001",
  47974=>"010110000",
  47975=>"011110110",
  47976=>"110000000",
  47977=>"111101100",
  47978=>"000011000",
  47979=>"000110110",
  47980=>"101000110",
  47981=>"010111100",
  47982=>"101010001",
  47983=>"101110000",
  47984=>"111100010",
  47985=>"010011010",
  47986=>"001011000",
  47987=>"011100011",
  47988=>"000010001",
  47989=>"100010100",
  47990=>"001110000",
  47991=>"110011110",
  47992=>"110011110",
  47993=>"010111011",
  47994=>"001111100",
  47995=>"000011001",
  47996=>"111000110",
  47997=>"000100110",
  47998=>"111111000",
  47999=>"101100001",
  48000=>"111101001",
  48001=>"001110010",
  48002=>"110011111",
  48003=>"010111000",
  48004=>"100101010",
  48005=>"100111000",
  48006=>"011010000",
  48007=>"111101010",
  48008=>"100000000",
  48009=>"100010000",
  48010=>"001110100",
  48011=>"010101010",
  48012=>"100100001",
  48013=>"001010110",
  48014=>"011101000",
  48015=>"000010010",
  48016=>"111010110",
  48017=>"010101110",
  48018=>"000001100",
  48019=>"111111100",
  48020=>"010110110",
  48021=>"111110010",
  48022=>"111100101",
  48023=>"111100000",
  48024=>"000001000",
  48025=>"001011010",
  48026=>"110010010",
  48027=>"111100100",
  48028=>"100111111",
  48029=>"010101101",
  48030=>"111101101",
  48031=>"110111001",
  48032=>"000011101",
  48033=>"100101000",
  48034=>"010100011",
  48035=>"100100110",
  48036=>"001010111",
  48037=>"101101000",
  48038=>"000100110",
  48039=>"010100000",
  48040=>"001111110",
  48041=>"010101100",
  48042=>"111000001",
  48043=>"110111101",
  48044=>"110100001",
  48045=>"001011101",
  48046=>"011001000",
  48047=>"001111011",
  48048=>"100000100",
  48049=>"000010010",
  48050=>"101111001",
  48051=>"110100110",
  48052=>"000011110",
  48053=>"110101100",
  48054=>"011111111",
  48055=>"000011110",
  48056=>"111100001",
  48057=>"111011100",
  48058=>"001010100",
  48059=>"101011011",
  48060=>"011011111",
  48061=>"100110100",
  48062=>"010000001",
  48063=>"111000001",
  48064=>"100010010",
  48065=>"100010011",
  48066=>"110111000",
  48067=>"000111100",
  48068=>"110111100",
  48069=>"011111111",
  48070=>"011001101",
  48071=>"001101100",
  48072=>"000000001",
  48073=>"001111000",
  48074=>"110100011",
  48075=>"011011101",
  48076=>"000111100",
  48077=>"101100100",
  48078=>"100000101",
  48079=>"110011110",
  48080=>"000000011",
  48081=>"000101011",
  48082=>"011001000",
  48083=>"100001011",
  48084=>"111100001",
  48085=>"000010000",
  48086=>"111010111",
  48087=>"011010111",
  48088=>"011101000",
  48089=>"011100111",
  48090=>"100010111",
  48091=>"010101000",
  48092=>"101010101",
  48093=>"010111110",
  48094=>"110110000",
  48095=>"010010100",
  48096=>"000100001",
  48097=>"001101110",
  48098=>"101000010",
  48099=>"111111010",
  48100=>"010000010",
  48101=>"101010111",
  48102=>"000011111",
  48103=>"100110100",
  48104=>"001101101",
  48105=>"001100110",
  48106=>"111101110",
  48107=>"110001110",
  48108=>"111111001",
  48109=>"000011001",
  48110=>"001101001",
  48111=>"010010111",
  48112=>"100000111",
  48113=>"011011111",
  48114=>"011011000",
  48115=>"101010010",
  48116=>"000111011",
  48117=>"010000000",
  48118=>"110100101",
  48119=>"111000010",
  48120=>"011011101",
  48121=>"100110010",
  48122=>"001001011",
  48123=>"111100110",
  48124=>"000000111",
  48125=>"100111100",
  48126=>"001011100",
  48127=>"001001011",
  48128=>"101111111",
  48129=>"100001101",
  48130=>"110110011",
  48131=>"100110010",
  48132=>"010011111",
  48133=>"110111101",
  48134=>"111011000",
  48135=>"100010011",
  48136=>"111101111",
  48137=>"000011111",
  48138=>"101101000",
  48139=>"010110001",
  48140=>"010000000",
  48141=>"000111011",
  48142=>"010110111",
  48143=>"111101101",
  48144=>"010011010",
  48145=>"011000010",
  48146=>"111011111",
  48147=>"110111001",
  48148=>"010110111",
  48149=>"000011101",
  48150=>"101011000",
  48151=>"011111001",
  48152=>"110011011",
  48153=>"111101101",
  48154=>"010101010",
  48155=>"100011110",
  48156=>"010010000",
  48157=>"011111011",
  48158=>"111111011",
  48159=>"101000100",
  48160=>"111000111",
  48161=>"110010111",
  48162=>"100010000",
  48163=>"101101001",
  48164=>"101111111",
  48165=>"100111111",
  48166=>"111010100",
  48167=>"011001110",
  48168=>"011100010",
  48169=>"111111111",
  48170=>"000101001",
  48171=>"001110110",
  48172=>"110001100",
  48173=>"011010000",
  48174=>"001011101",
  48175=>"110010011",
  48176=>"110000001",
  48177=>"010110010",
  48178=>"101001000",
  48179=>"100000000",
  48180=>"111111111",
  48181=>"101111011",
  48182=>"100010000",
  48183=>"101110011",
  48184=>"111111110",
  48185=>"000001000",
  48186=>"001011100",
  48187=>"110110011",
  48188=>"110001101",
  48189=>"001110011",
  48190=>"011100100",
  48191=>"111100000",
  48192=>"000100110",
  48193=>"000001000",
  48194=>"100110010",
  48195=>"111101110",
  48196=>"010110111",
  48197=>"100110010",
  48198=>"001101111",
  48199=>"001111100",
  48200=>"001011011",
  48201=>"011100000",
  48202=>"011000000",
  48203=>"111101101",
  48204=>"111110110",
  48205=>"111100111",
  48206=>"101110011",
  48207=>"001100011",
  48208=>"110100011",
  48209=>"000101001",
  48210=>"100010000",
  48211=>"011001100",
  48212=>"010011101",
  48213=>"011000110",
  48214=>"100010100",
  48215=>"000110111",
  48216=>"101111110",
  48217=>"110000110",
  48218=>"111100111",
  48219=>"110100001",
  48220=>"111000111",
  48221=>"000000100",
  48222=>"110110110",
  48223=>"100100010",
  48224=>"100100111",
  48225=>"011101000",
  48226=>"111010100",
  48227=>"010110100",
  48228=>"000101100",
  48229=>"110011101",
  48230=>"100000001",
  48231=>"100000000",
  48232=>"101111010",
  48233=>"011111011",
  48234=>"001000000",
  48235=>"010100100",
  48236=>"111110011",
  48237=>"111110110",
  48238=>"111000101",
  48239=>"110001010",
  48240=>"100101011",
  48241=>"010000011",
  48242=>"101001101",
  48243=>"111011001",
  48244=>"001010111",
  48245=>"111001011",
  48246=>"110111010",
  48247=>"101000000",
  48248=>"101110001",
  48249=>"001100011",
  48250=>"111011101",
  48251=>"100101111",
  48252=>"010100110",
  48253=>"000011010",
  48254=>"111111101",
  48255=>"011010010",
  48256=>"111011011",
  48257=>"001011100",
  48258=>"110100000",
  48259=>"011000000",
  48260=>"000111000",
  48261=>"000100010",
  48262=>"101101111",
  48263=>"100000001",
  48264=>"110011001",
  48265=>"000100101",
  48266=>"001000010",
  48267=>"101101000",
  48268=>"111011110",
  48269=>"000111010",
  48270=>"101010010",
  48271=>"110000001",
  48272=>"110110101",
  48273=>"000110100",
  48274=>"000001101",
  48275=>"010110001",
  48276=>"110101010",
  48277=>"111000011",
  48278=>"011011010",
  48279=>"000011101",
  48280=>"010111010",
  48281=>"100011011",
  48282=>"011100111",
  48283=>"000111011",
  48284=>"000000010",
  48285=>"000011100",
  48286=>"111111111",
  48287=>"110011000",
  48288=>"001101110",
  48289=>"110100000",
  48290=>"001110000",
  48291=>"100111100",
  48292=>"101010000",
  48293=>"110111000",
  48294=>"101000101",
  48295=>"010110111",
  48296=>"000011001",
  48297=>"011110010",
  48298=>"011000010",
  48299=>"111011001",
  48300=>"110101000",
  48301=>"111110000",
  48302=>"111100100",
  48303=>"100111100",
  48304=>"010101011",
  48305=>"101011111",
  48306=>"111101111",
  48307=>"100111000",
  48308=>"111101101",
  48309=>"101100111",
  48310=>"010010101",
  48311=>"000000010",
  48312=>"000010111",
  48313=>"010000101",
  48314=>"001011111",
  48315=>"101111011",
  48316=>"000010100",
  48317=>"001000010",
  48318=>"000011110",
  48319=>"011000101",
  48320=>"000000001",
  48321=>"000011110",
  48322=>"011101110",
  48323=>"100110111",
  48324=>"010011001",
  48325=>"001111011",
  48326=>"010000100",
  48327=>"001001011",
  48328=>"011100110",
  48329=>"011001001",
  48330=>"110001000",
  48331=>"011011011",
  48332=>"010010010",
  48333=>"101000010",
  48334=>"111100100",
  48335=>"100001111",
  48336=>"001010110",
  48337=>"001101001",
  48338=>"000111000",
  48339=>"001110111",
  48340=>"111011001",
  48341=>"110010110",
  48342=>"111111100",
  48343=>"100010011",
  48344=>"100111100",
  48345=>"000001000",
  48346=>"101001111",
  48347=>"111111011",
  48348=>"101001110",
  48349=>"011111011",
  48350=>"001100000",
  48351=>"101011111",
  48352=>"110101010",
  48353=>"010100011",
  48354=>"111011001",
  48355=>"110100001",
  48356=>"111011011",
  48357=>"111101000",
  48358=>"001001111",
  48359=>"101011000",
  48360=>"100101000",
  48361=>"010101111",
  48362=>"011011011",
  48363=>"111000000",
  48364=>"001101010",
  48365=>"100010001",
  48366=>"101100011",
  48367=>"000111101",
  48368=>"111101110",
  48369=>"000001110",
  48370=>"001010111",
  48371=>"000110100",
  48372=>"001100011",
  48373=>"100110100",
  48374=>"111100100",
  48375=>"010110011",
  48376=>"111010111",
  48377=>"000101101",
  48378=>"111010000",
  48379=>"010111110",
  48380=>"011010000",
  48381=>"101100100",
  48382=>"011111101",
  48383=>"010100100",
  48384=>"100000011",
  48385=>"110110000",
  48386=>"101011011",
  48387=>"111101011",
  48388=>"111000110",
  48389=>"101010000",
  48390=>"101110111",
  48391=>"010100010",
  48392=>"100101100",
  48393=>"100001101",
  48394=>"000110001",
  48395=>"011110010",
  48396=>"101101011",
  48397=>"011110011",
  48398=>"010000111",
  48399=>"100111110",
  48400=>"001000111",
  48401=>"011000001",
  48402=>"000000100",
  48403=>"001101011",
  48404=>"011010101",
  48405=>"011100101",
  48406=>"101000101",
  48407=>"100110000",
  48408=>"100001101",
  48409=>"010110011",
  48410=>"101000110",
  48411=>"001011000",
  48412=>"001011000",
  48413=>"001000111",
  48414=>"000110010",
  48415=>"100000001",
  48416=>"110101100",
  48417=>"000000111",
  48418=>"001011100",
  48419=>"000001110",
  48420=>"010011011",
  48421=>"001011111",
  48422=>"110001001",
  48423=>"011000010",
  48424=>"011000001",
  48425=>"011010010",
  48426=>"101101001",
  48427=>"101000000",
  48428=>"101001100",
  48429=>"010100101",
  48430=>"010000110",
  48431=>"010101000",
  48432=>"100101101",
  48433=>"011110100",
  48434=>"011001110",
  48435=>"000000101",
  48436=>"110001001",
  48437=>"101101101",
  48438=>"000100000",
  48439=>"110110101",
  48440=>"000010000",
  48441=>"001110010",
  48442=>"111111100",
  48443=>"010000100",
  48444=>"010011011",
  48445=>"001111011",
  48446=>"100101110",
  48447=>"111001101",
  48448=>"111110001",
  48449=>"000010111",
  48450=>"101101101",
  48451=>"110010000",
  48452=>"110101111",
  48453=>"000010111",
  48454=>"001111100",
  48455=>"000000110",
  48456=>"001100111",
  48457=>"100000000",
  48458=>"100011100",
  48459=>"011010001",
  48460=>"000101111",
  48461=>"110111001",
  48462=>"101100100",
  48463=>"110110110",
  48464=>"010011011",
  48465=>"011101001",
  48466=>"000001110",
  48467=>"010111111",
  48468=>"000001100",
  48469=>"001110100",
  48470=>"110011000",
  48471=>"001100100",
  48472=>"110101110",
  48473=>"110000010",
  48474=>"101001000",
  48475=>"010001101",
  48476=>"100110001",
  48477=>"101101000",
  48478=>"111110011",
  48479=>"110100100",
  48480=>"000000111",
  48481=>"100011010",
  48482=>"000011000",
  48483=>"000111101",
  48484=>"011100101",
  48485=>"111101111",
  48486=>"011101110",
  48487=>"001000100",
  48488=>"101111101",
  48489=>"111111011",
  48490=>"100011101",
  48491=>"000110110",
  48492=>"001000011",
  48493=>"111011111",
  48494=>"001111001",
  48495=>"000100110",
  48496=>"101111001",
  48497=>"110011011",
  48498=>"110110101",
  48499=>"101001000",
  48500=>"101010000",
  48501=>"000000011",
  48502=>"111111010",
  48503=>"100010000",
  48504=>"010000001",
  48505=>"010001110",
  48506=>"100010100",
  48507=>"101010000",
  48508=>"000111111",
  48509=>"111010011",
  48510=>"101101001",
  48511=>"111100101",
  48512=>"001110100",
  48513=>"001001111",
  48514=>"000111101",
  48515=>"000110100",
  48516=>"010001001",
  48517=>"001000001",
  48518=>"100100100",
  48519=>"010010100",
  48520=>"101111011",
  48521=>"110000010",
  48522=>"101100111",
  48523=>"011100001",
  48524=>"111100011",
  48525=>"001111011",
  48526=>"101010111",
  48527=>"111110000",
  48528=>"010100010",
  48529=>"000110110",
  48530=>"111010101",
  48531=>"001110110",
  48532=>"101000011",
  48533=>"111100010",
  48534=>"100011100",
  48535=>"111111111",
  48536=>"111111101",
  48537=>"000001111",
  48538=>"001001001",
  48539=>"000010111",
  48540=>"000010100",
  48541=>"111010101",
  48542=>"101110100",
  48543=>"110010000",
  48544=>"100011111",
  48545=>"011110101",
  48546=>"111100100",
  48547=>"000000001",
  48548=>"001100100",
  48549=>"100100000",
  48550=>"100101111",
  48551=>"111010000",
  48552=>"001100000",
  48553=>"011011100",
  48554=>"010000010",
  48555=>"001100101",
  48556=>"101000111",
  48557=>"100110011",
  48558=>"101001010",
  48559=>"101011100",
  48560=>"001010111",
  48561=>"001101100",
  48562=>"100110010",
  48563=>"111001110",
  48564=>"000110110",
  48565=>"101011010",
  48566=>"110011110",
  48567=>"001010001",
  48568=>"100001101",
  48569=>"000101101",
  48570=>"111011100",
  48571=>"011100010",
  48572=>"000111111",
  48573=>"101001101",
  48574=>"000100101",
  48575=>"101110001",
  48576=>"000101100",
  48577=>"100011101",
  48578=>"010111100",
  48579=>"111111011",
  48580=>"000001100",
  48581=>"001001100",
  48582=>"111011100",
  48583=>"101000111",
  48584=>"000110100",
  48585=>"011001110",
  48586=>"001010000",
  48587=>"101011100",
  48588=>"011110101",
  48589=>"010101010",
  48590=>"000100110",
  48591=>"010010010",
  48592=>"010110000",
  48593=>"011100010",
  48594=>"111111011",
  48595=>"000001101",
  48596=>"100011110",
  48597=>"010001110",
  48598=>"110000111",
  48599=>"101001011",
  48600=>"000001011",
  48601=>"001110110",
  48602=>"001100000",
  48603=>"010111110",
  48604=>"101000111",
  48605=>"011001000",
  48606=>"011010111",
  48607=>"010101111",
  48608=>"100111111",
  48609=>"001000000",
  48610=>"101011111",
  48611=>"001001100",
  48612=>"010100010",
  48613=>"000010011",
  48614=>"110100011",
  48615=>"000110000",
  48616=>"110110001",
  48617=>"101101001",
  48618=>"100000111",
  48619=>"111110010",
  48620=>"000001100",
  48621=>"001000011",
  48622=>"110111110",
  48623=>"010000000",
  48624=>"001000000",
  48625=>"011101111",
  48626=>"111010000",
  48627=>"111011011",
  48628=>"001001111",
  48629=>"101101001",
  48630=>"101001110",
  48631=>"110111111",
  48632=>"110111011",
  48633=>"000110110",
  48634=>"011100101",
  48635=>"011001110",
  48636=>"000000001",
  48637=>"100111101",
  48638=>"011111111",
  48639=>"001111010",
  48640=>"001010011",
  48641=>"101011010",
  48642=>"101111011",
  48643=>"000111010",
  48644=>"010011110",
  48645=>"111100011",
  48646=>"000100001",
  48647=>"110010010",
  48648=>"011100111",
  48649=>"110101010",
  48650=>"010001001",
  48651=>"011110001",
  48652=>"010010000",
  48653=>"100011011",
  48654=>"100001111",
  48655=>"010110111",
  48656=>"011110111",
  48657=>"001011000",
  48658=>"110011001",
  48659=>"001001101",
  48660=>"010011100",
  48661=>"111000010",
  48662=>"010001000",
  48663=>"000011111",
  48664=>"010011010",
  48665=>"110100010",
  48666=>"001010011",
  48667=>"111101100",
  48668=>"011011101",
  48669=>"111001011",
  48670=>"000011100",
  48671=>"011010001",
  48672=>"100111001",
  48673=>"000001101",
  48674=>"100001011",
  48675=>"111110010",
  48676=>"110110000",
  48677=>"101110011",
  48678=>"011100100",
  48679=>"000100010",
  48680=>"010110010",
  48681=>"010111010",
  48682=>"000101010",
  48683=>"001001100",
  48684=>"000111011",
  48685=>"010000000",
  48686=>"110010001",
  48687=>"101100101",
  48688=>"101001110",
  48689=>"011010100",
  48690=>"000011100",
  48691=>"010011111",
  48692=>"011111001",
  48693=>"011001001",
  48694=>"100100001",
  48695=>"100101111",
  48696=>"001001111",
  48697=>"010010111",
  48698=>"111010100",
  48699=>"110000001",
  48700=>"001110001",
  48701=>"000000101",
  48702=>"100010100",
  48703=>"011101001",
  48704=>"001010101",
  48705=>"100100100",
  48706=>"101001100",
  48707=>"111001011",
  48708=>"000000000",
  48709=>"101111101",
  48710=>"110111111",
  48711=>"000111110",
  48712=>"000011100",
  48713=>"010001000",
  48714=>"001110001",
  48715=>"001001101",
  48716=>"011101010",
  48717=>"000001100",
  48718=>"100100100",
  48719=>"010010111",
  48720=>"011111101",
  48721=>"011010101",
  48722=>"001011110",
  48723=>"010000110",
  48724=>"110101111",
  48725=>"110110100",
  48726=>"101101011",
  48727=>"011000111",
  48728=>"101001001",
  48729=>"101111110",
  48730=>"011010100",
  48731=>"000011100",
  48732=>"010011101",
  48733=>"100111001",
  48734=>"100000000",
  48735=>"000011011",
  48736=>"110010111",
  48737=>"011010010",
  48738=>"000001010",
  48739=>"000011001",
  48740=>"100010011",
  48741=>"001001001",
  48742=>"110000000",
  48743=>"100101110",
  48744=>"010100111",
  48745=>"111011011",
  48746=>"000101010",
  48747=>"110010111",
  48748=>"100010010",
  48749=>"101111101",
  48750=>"100100111",
  48751=>"010001011",
  48752=>"110011110",
  48753=>"000011110",
  48754=>"111011100",
  48755=>"111001111",
  48756=>"000010101",
  48757=>"100010110",
  48758=>"110100101",
  48759=>"010111001",
  48760=>"101011111",
  48761=>"100001110",
  48762=>"010111011",
  48763=>"100010001",
  48764=>"010000110",
  48765=>"110111001",
  48766=>"001101111",
  48767=>"101100010",
  48768=>"001100110",
  48769=>"100100010",
  48770=>"010010001",
  48771=>"110101110",
  48772=>"011001101",
  48773=>"111011011",
  48774=>"010010000",
  48775=>"011011100",
  48776=>"111101110",
  48777=>"001001100",
  48778=>"111111111",
  48779=>"111111011",
  48780=>"000010010",
  48781=>"000111011",
  48782=>"001111000",
  48783=>"101000101",
  48784=>"011000001",
  48785=>"101001100",
  48786=>"111100111",
  48787=>"110010000",
  48788=>"000000111",
  48789=>"001110000",
  48790=>"000100010",
  48791=>"110001010",
  48792=>"011101010",
  48793=>"101010010",
  48794=>"111111101",
  48795=>"111110010",
  48796=>"100000001",
  48797=>"010110101",
  48798=>"010011101",
  48799=>"101000010",
  48800=>"001001100",
  48801=>"110110111",
  48802=>"000000101",
  48803=>"011000010",
  48804=>"111001111",
  48805=>"010101110",
  48806=>"001001110",
  48807=>"001010000",
  48808=>"110011010",
  48809=>"111100111",
  48810=>"101111100",
  48811=>"001111011",
  48812=>"000010110",
  48813=>"001111111",
  48814=>"000100001",
  48815=>"001100010",
  48816=>"001110010",
  48817=>"000001010",
  48818=>"001011000",
  48819=>"101000110",
  48820=>"001011110",
  48821=>"110000100",
  48822=>"111110010",
  48823=>"100110111",
  48824=>"010000010",
  48825=>"100110011",
  48826=>"000011011",
  48827=>"001010011",
  48828=>"000011111",
  48829=>"000110011",
  48830=>"000111100",
  48831=>"100110000",
  48832=>"100001100",
  48833=>"110010011",
  48834=>"101011111",
  48835=>"111010000",
  48836=>"111101010",
  48837=>"111001011",
  48838=>"101010010",
  48839=>"001010000",
  48840=>"111011111",
  48841=>"100100010",
  48842=>"100010101",
  48843=>"110110011",
  48844=>"010111001",
  48845=>"110111110",
  48846=>"010100011",
  48847=>"101111100",
  48848=>"011001000",
  48849=>"101000001",
  48850=>"111010001",
  48851=>"110101101",
  48852=>"001001000",
  48853=>"110101111",
  48854=>"111100100",
  48855=>"010001101",
  48856=>"111001011",
  48857=>"011111001",
  48858=>"110100000",
  48859=>"101100000",
  48860=>"111011000",
  48861=>"111101101",
  48862=>"011000000",
  48863=>"011100110",
  48864=>"101010001",
  48865=>"100100110",
  48866=>"000101101",
  48867=>"001111001",
  48868=>"100000110",
  48869=>"011000001",
  48870=>"110100100",
  48871=>"010101001",
  48872=>"111101101",
  48873=>"110110110",
  48874=>"111011011",
  48875=>"010011111",
  48876=>"000000111",
  48877=>"100101101",
  48878=>"010000000",
  48879=>"101111000",
  48880=>"001010110",
  48881=>"111011111",
  48882=>"101000010",
  48883=>"100011000",
  48884=>"100101010",
  48885=>"001101101",
  48886=>"111011110",
  48887=>"000100100",
  48888=>"011100010",
  48889=>"001001101",
  48890=>"010010101",
  48891=>"100110000",
  48892=>"001110001",
  48893=>"111000100",
  48894=>"001100011",
  48895=>"111101111",
  48896=>"001110000",
  48897=>"110111010",
  48898=>"000000000",
  48899=>"000100000",
  48900=>"000100111",
  48901=>"001001100",
  48902=>"011110011",
  48903=>"001000110",
  48904=>"001000010",
  48905=>"111001000",
  48906=>"000001111",
  48907=>"100010110",
  48908=>"001110110",
  48909=>"000010010",
  48910=>"110100001",
  48911=>"101011101",
  48912=>"110011010",
  48913=>"100101011",
  48914=>"001100100",
  48915=>"001001001",
  48916=>"100011011",
  48917=>"011100100",
  48918=>"010011001",
  48919=>"101110101",
  48920=>"011011001",
  48921=>"011010100",
  48922=>"111111111",
  48923=>"111100011",
  48924=>"110110001",
  48925=>"110001100",
  48926=>"111000000",
  48927=>"110100001",
  48928=>"110100100",
  48929=>"101000111",
  48930=>"000110010",
  48931=>"000011011",
  48932=>"000100011",
  48933=>"111111111",
  48934=>"010000100",
  48935=>"011100011",
  48936=>"000010100",
  48937=>"001011001",
  48938=>"110010110",
  48939=>"110110000",
  48940=>"001010011",
  48941=>"010001001",
  48942=>"111110101",
  48943=>"111111000",
  48944=>"111011100",
  48945=>"000000010",
  48946=>"100111101",
  48947=>"001110010",
  48948=>"110111101",
  48949=>"110010001",
  48950=>"101001111",
  48951=>"111101111",
  48952=>"101001100",
  48953=>"111001000",
  48954=>"000010000",
  48955=>"100101011",
  48956=>"110010011",
  48957=>"101111110",
  48958=>"001100110",
  48959=>"001000001",
  48960=>"000101110",
  48961=>"001110010",
  48962=>"110110100",
  48963=>"000011010",
  48964=>"110100010",
  48965=>"001111110",
  48966=>"100001111",
  48967=>"111111101",
  48968=>"011111101",
  48969=>"010111010",
  48970=>"011100100",
  48971=>"010101100",
  48972=>"100000011",
  48973=>"110110111",
  48974=>"111010000",
  48975=>"000010110",
  48976=>"100111111",
  48977=>"101100001",
  48978=>"100000101",
  48979=>"101101011",
  48980=>"001000011",
  48981=>"110110100",
  48982=>"111101110",
  48983=>"001010000",
  48984=>"010001111",
  48985=>"010110101",
  48986=>"111110010",
  48987=>"101111111",
  48988=>"101000101",
  48989=>"001111011",
  48990=>"100111000",
  48991=>"101000111",
  48992=>"110010010",
  48993=>"101111010",
  48994=>"111011110",
  48995=>"010100010",
  48996=>"001111111",
  48997=>"100010101",
  48998=>"111100010",
  48999=>"000011001",
  49000=>"001101101",
  49001=>"011101001",
  49002=>"011100011",
  49003=>"000111001",
  49004=>"001001010",
  49005=>"101110111",
  49006=>"111111010",
  49007=>"101010000",
  49008=>"000000100",
  49009=>"000100011",
  49010=>"111100111",
  49011=>"100000011",
  49012=>"110100010",
  49013=>"000010110",
  49014=>"110110111",
  49015=>"001000011",
  49016=>"000011011",
  49017=>"111100001",
  49018=>"011001101",
  49019=>"101001011",
  49020=>"011010111",
  49021=>"011100000",
  49022=>"001110100",
  49023=>"110000100",
  49024=>"101001111",
  49025=>"000011101",
  49026=>"101011100",
  49027=>"111101111",
  49028=>"001010111",
  49029=>"110011111",
  49030=>"010110000",
  49031=>"000011001",
  49032=>"010100000",
  49033=>"101000001",
  49034=>"110000110",
  49035=>"010010110",
  49036=>"100000101",
  49037=>"010100010",
  49038=>"110011011",
  49039=>"101111000",
  49040=>"110111110",
  49041=>"010110110",
  49042=>"000011101",
  49043=>"111011011",
  49044=>"000000101",
  49045=>"110101110",
  49046=>"100101000",
  49047=>"011110011",
  49048=>"001000110",
  49049=>"000000111",
  49050=>"010001000",
  49051=>"000101100",
  49052=>"001000100",
  49053=>"001101010",
  49054=>"110001111",
  49055=>"110110000",
  49056=>"011001010",
  49057=>"011011001",
  49058=>"010100011",
  49059=>"001111111",
  49060=>"011011101",
  49061=>"111010010",
  49062=>"010101110",
  49063=>"111100110",
  49064=>"010111111",
  49065=>"010100110",
  49066=>"010101111",
  49067=>"001000001",
  49068=>"011110000",
  49069=>"001011011",
  49070=>"101101111",
  49071=>"111110010",
  49072=>"111111010",
  49073=>"110111111",
  49074=>"100001111",
  49075=>"000001000",
  49076=>"001001101",
  49077=>"010101010",
  49078=>"000100111",
  49079=>"001100101",
  49080=>"110110111",
  49081=>"110101011",
  49082=>"011101110",
  49083=>"011001010",
  49084=>"010100100",
  49085=>"100001101",
  49086=>"111001101",
  49087=>"001110011",
  49088=>"011110100",
  49089=>"001001001",
  49090=>"101110010",
  49091=>"011000010",
  49092=>"111010000",
  49093=>"001111100",
  49094=>"010001100",
  49095=>"011000100",
  49096=>"110001111",
  49097=>"111000001",
  49098=>"000001011",
  49099=>"011110010",
  49100=>"110000100",
  49101=>"011001000",
  49102=>"101111011",
  49103=>"111000010",
  49104=>"111100000",
  49105=>"000001011",
  49106=>"110010101",
  49107=>"011101001",
  49108=>"111000011",
  49109=>"111111101",
  49110=>"000100111",
  49111=>"000100001",
  49112=>"110000111",
  49113=>"011010110",
  49114=>"100100011",
  49115=>"101000111",
  49116=>"101000010",
  49117=>"001110100",
  49118=>"010001011",
  49119=>"000011100",
  49120=>"011101111",
  49121=>"110100001",
  49122=>"010111101",
  49123=>"001111001",
  49124=>"000100111",
  49125=>"010001101",
  49126=>"111011001",
  49127=>"111111011",
  49128=>"000010010",
  49129=>"010100111",
  49130=>"010011100",
  49131=>"111101011",
  49132=>"101000001",
  49133=>"000010010",
  49134=>"011100000",
  49135=>"000111010",
  49136=>"111110000",
  49137=>"011011100",
  49138=>"010011001",
  49139=>"111101001",
  49140=>"100101110",
  49141=>"011101000",
  49142=>"011101001",
  49143=>"011011000",
  49144=>"010000010",
  49145=>"101010011",
  49146=>"110001010",
  49147=>"001100110",
  49148=>"101010101",
  49149=>"000010000",
  49150=>"000100000",
  49151=>"010010010",
  49152=>"000100100",
  49153=>"010001110",
  49154=>"111101110",
  49155=>"010011111",
  49156=>"011011111",
  49157=>"101000000",
  49158=>"001010111",
  49159=>"111010000",
  49160=>"101101010",
  49161=>"111110101",
  49162=>"001010100",
  49163=>"010001101",
  49164=>"100001101",
  49165=>"000101110",
  49166=>"101001111",
  49167=>"011111111",
  49168=>"100110100",
  49169=>"100000101",
  49170=>"011110111",
  49171=>"010111100",
  49172=>"001001000",
  49173=>"100101001",
  49174=>"111010010",
  49175=>"010001011",
  49176=>"001001111",
  49177=>"011000100",
  49178=>"010000110",
  49179=>"010001011",
  49180=>"100100011",
  49181=>"110110001",
  49182=>"110110010",
  49183=>"101101010",
  49184=>"100001101",
  49185=>"000010111",
  49186=>"110011101",
  49187=>"101010000",
  49188=>"000010001",
  49189=>"011110010",
  49190=>"010100100",
  49191=>"100100011",
  49192=>"000010111",
  49193=>"001001111",
  49194=>"011001100",
  49195=>"100100110",
  49196=>"001111011",
  49197=>"011111101",
  49198=>"110010001",
  49199=>"100100101",
  49200=>"111000011",
  49201=>"111101000",
  49202=>"011000001",
  49203=>"000010110",
  49204=>"000001001",
  49205=>"100011000",
  49206=>"011101000",
  49207=>"000001001",
  49208=>"101110010",
  49209=>"011000001",
  49210=>"101100001",
  49211=>"101000001",
  49212=>"011111101",
  49213=>"001101111",
  49214=>"101011011",
  49215=>"000000011",
  49216=>"010100010",
  49217=>"111000001",
  49218=>"001001010",
  49219=>"110001100",
  49220=>"111010000",
  49221=>"111111011",
  49222=>"000110101",
  49223=>"110100101",
  49224=>"110101011",
  49225=>"101001111",
  49226=>"011010010",
  49227=>"000001100",
  49228=>"111001110",
  49229=>"110011001",
  49230=>"010100000",
  49231=>"101010111",
  49232=>"111100110",
  49233=>"110001011",
  49234=>"111111111",
  49235=>"010000101",
  49236=>"011011111",
  49237=>"001010110",
  49238=>"000111110",
  49239=>"010101011",
  49240=>"101001101",
  49241=>"110101110",
  49242=>"111110111",
  49243=>"100000100",
  49244=>"011111111",
  49245=>"011100100",
  49246=>"101011001",
  49247=>"110001011",
  49248=>"110101010",
  49249=>"100000110",
  49250=>"001001001",
  49251=>"011111001",
  49252=>"100000100",
  49253=>"000110011",
  49254=>"111100011",
  49255=>"010111111",
  49256=>"010110111",
  49257=>"001100110",
  49258=>"000111001",
  49259=>"101100100",
  49260=>"011110010",
  49261=>"111011000",
  49262=>"000000101",
  49263=>"010100100",
  49264=>"101000011",
  49265=>"111110101",
  49266=>"001001011",
  49267=>"001110001",
  49268=>"010001001",
  49269=>"000000110",
  49270=>"000011101",
  49271=>"111101011",
  49272=>"011100100",
  49273=>"100010011",
  49274=>"011011001",
  49275=>"101001101",
  49276=>"000101110",
  49277=>"100101101",
  49278=>"000000001",
  49279=>"100111101",
  49280=>"000100010",
  49281=>"001110111",
  49282=>"001111011",
  49283=>"000010110",
  49284=>"010101101",
  49285=>"010001101",
  49286=>"100110000",
  49287=>"101011111",
  49288=>"000111110",
  49289=>"100000000",
  49290=>"000001000",
  49291=>"111100111",
  49292=>"101111100",
  49293=>"000011101",
  49294=>"110010111",
  49295=>"101010010",
  49296=>"010111101",
  49297=>"101111101",
  49298=>"101010000",
  49299=>"000011000",
  49300=>"001111111",
  49301=>"000101101",
  49302=>"100001001",
  49303=>"110010000",
  49304=>"000011001",
  49305=>"100001101",
  49306=>"011010011",
  49307=>"101000101",
  49308=>"110100110",
  49309=>"100111110",
  49310=>"000100011",
  49311=>"100010001",
  49312=>"010101001",
  49313=>"000011110",
  49314=>"001110101",
  49315=>"010000110",
  49316=>"111000100",
  49317=>"001100101",
  49318=>"100111001",
  49319=>"001111011",
  49320=>"110001001",
  49321=>"010010010",
  49322=>"010010110",
  49323=>"111000111",
  49324=>"001011010",
  49325=>"000110010",
  49326=>"011010001",
  49327=>"101000001",
  49328=>"000100001",
  49329=>"001111011",
  49330=>"101100111",
  49331=>"100001000",
  49332=>"100100110",
  49333=>"001000000",
  49334=>"001100111",
  49335=>"100011111",
  49336=>"001010010",
  49337=>"111111111",
  49338=>"110111010",
  49339=>"110010001",
  49340=>"001111001",
  49341=>"110101001",
  49342=>"100111101",
  49343=>"001010101",
  49344=>"110111011",
  49345=>"000110010",
  49346=>"011101101",
  49347=>"000011010",
  49348=>"011010011",
  49349=>"011011101",
  49350=>"011010001",
  49351=>"100010011",
  49352=>"011000011",
  49353=>"110001001",
  49354=>"000100011",
  49355=>"011010001",
  49356=>"101010000",
  49357=>"011111011",
  49358=>"010100001",
  49359=>"000100001",
  49360=>"100101000",
  49361=>"101101111",
  49362=>"000101101",
  49363=>"010001000",
  49364=>"100111101",
  49365=>"101101100",
  49366=>"000000001",
  49367=>"111011101",
  49368=>"101000011",
  49369=>"101110010",
  49370=>"100001000",
  49371=>"000101111",
  49372=>"100001000",
  49373=>"110011101",
  49374=>"101000000",
  49375=>"000001110",
  49376=>"100101100",
  49377=>"111010111",
  49378=>"100011111",
  49379=>"111111001",
  49380=>"000111011",
  49381=>"000000100",
  49382=>"010100001",
  49383=>"100100101",
  49384=>"001010100",
  49385=>"000110100",
  49386=>"101100110",
  49387=>"011110010",
  49388=>"101111010",
  49389=>"000100001",
  49390=>"001101001",
  49391=>"101101010",
  49392=>"010011110",
  49393=>"011100111",
  49394=>"101100011",
  49395=>"011110111",
  49396=>"000110110",
  49397=>"101101111",
  49398=>"000001110",
  49399=>"100000001",
  49400=>"010011011",
  49401=>"101001111",
  49402=>"001111101",
  49403=>"000001010",
  49404=>"100010010",
  49405=>"100110001",
  49406=>"111110110",
  49407=>"100000110",
  49408=>"111000001",
  49409=>"101000000",
  49410=>"000111100",
  49411=>"010010010",
  49412=>"000111111",
  49413=>"010110100",
  49414=>"101100010",
  49415=>"111001010",
  49416=>"100100111",
  49417=>"111101010",
  49418=>"000000100",
  49419=>"001100101",
  49420=>"011110011",
  49421=>"110111111",
  49422=>"101000010",
  49423=>"010010000",
  49424=>"111001110",
  49425=>"111011011",
  49426=>"010000101",
  49427=>"110111111",
  49428=>"101101000",
  49429=>"000101010",
  49430=>"100100101",
  49431=>"101111111",
  49432=>"000001010",
  49433=>"000101110",
  49434=>"110111010",
  49435=>"111111000",
  49436=>"111101111",
  49437=>"001000110",
  49438=>"011010011",
  49439=>"011010101",
  49440=>"101000011",
  49441=>"010110000",
  49442=>"111001111",
  49443=>"011110101",
  49444=>"001000100",
  49445=>"111011011",
  49446=>"111000111",
  49447=>"111011000",
  49448=>"010011101",
  49449=>"001110110",
  49450=>"110001110",
  49451=>"111100000",
  49452=>"100000000",
  49453=>"010101101",
  49454=>"000100000",
  49455=>"101101011",
  49456=>"011100111",
  49457=>"000010001",
  49458=>"111101101",
  49459=>"101110000",
  49460=>"101110111",
  49461=>"100011110",
  49462=>"001111011",
  49463=>"001001000",
  49464=>"100111011",
  49465=>"100011110",
  49466=>"011001111",
  49467=>"111101111",
  49468=>"110011010",
  49469=>"111001101",
  49470=>"110100010",
  49471=>"110000101",
  49472=>"111111111",
  49473=>"111000101",
  49474=>"000001100",
  49475=>"111100001",
  49476=>"101000001",
  49477=>"100010111",
  49478=>"101001000",
  49479=>"100111100",
  49480=>"011011010",
  49481=>"110010000",
  49482=>"100010011",
  49483=>"000000000",
  49484=>"110101100",
  49485=>"001101101",
  49486=>"010001010",
  49487=>"011010011",
  49488=>"111010100",
  49489=>"011011010",
  49490=>"101001100",
  49491=>"110001100",
  49492=>"000001111",
  49493=>"110111011",
  49494=>"011100101",
  49495=>"001100101",
  49496=>"110000110",
  49497=>"111101110",
  49498=>"011111110",
  49499=>"100000100",
  49500=>"010110011",
  49501=>"011010101",
  49502=>"000110011",
  49503=>"000011011",
  49504=>"110010001",
  49505=>"010000000",
  49506=>"001100011",
  49507=>"111101110",
  49508=>"000110011",
  49509=>"000100001",
  49510=>"000000100",
  49511=>"001000100",
  49512=>"001010001",
  49513=>"111110010",
  49514=>"010101000",
  49515=>"111111101",
  49516=>"101110001",
  49517=>"111111001",
  49518=>"010001011",
  49519=>"101111001",
  49520=>"010111000",
  49521=>"100010100",
  49522=>"000101110",
  49523=>"100001110",
  49524=>"100111100",
  49525=>"101001011",
  49526=>"101111110",
  49527=>"111100111",
  49528=>"000100101",
  49529=>"000000101",
  49530=>"101110000",
  49531=>"000011101",
  49532=>"000111100",
  49533=>"110100011",
  49534=>"100011011",
  49535=>"110010010",
  49536=>"000001010",
  49537=>"001011111",
  49538=>"010101101",
  49539=>"010010111",
  49540=>"011101000",
  49541=>"011001101",
  49542=>"100100111",
  49543=>"101001111",
  49544=>"010110001",
  49545=>"001001010",
  49546=>"101111000",
  49547=>"001000010",
  49548=>"101001101",
  49549=>"011111011",
  49550=>"001001100",
  49551=>"010000101",
  49552=>"100111011",
  49553=>"110000101",
  49554=>"001001111",
  49555=>"110111111",
  49556=>"111001001",
  49557=>"100010001",
  49558=>"100100011",
  49559=>"111001001",
  49560=>"011100100",
  49561=>"001001100",
  49562=>"101111101",
  49563=>"000001001",
  49564=>"101101110",
  49565=>"110100100",
  49566=>"011100101",
  49567=>"001110011",
  49568=>"000010111",
  49569=>"101001101",
  49570=>"111110001",
  49571=>"000011000",
  49572=>"001010110",
  49573=>"001000001",
  49574=>"011101100",
  49575=>"010101101",
  49576=>"010101011",
  49577=>"110000000",
  49578=>"111011111",
  49579=>"101111111",
  49580=>"001000101",
  49581=>"110011110",
  49582=>"000110001",
  49583=>"101011001",
  49584=>"011000101",
  49585=>"100101001",
  49586=>"000010110",
  49587=>"110001010",
  49588=>"000111111",
  49589=>"111011001",
  49590=>"010110100",
  49591=>"001000100",
  49592=>"101101011",
  49593=>"011100011",
  49594=>"000100011",
  49595=>"101111111",
  49596=>"011001010",
  49597=>"101000101",
  49598=>"000011110",
  49599=>"101111111",
  49600=>"001011001",
  49601=>"001001110",
  49602=>"011010011",
  49603=>"110100100",
  49604=>"010000101",
  49605=>"100100101",
  49606=>"110010110",
  49607=>"000011111",
  49608=>"011001101",
  49609=>"011110100",
  49610=>"101001010",
  49611=>"010111010",
  49612=>"010110010",
  49613=>"101111000",
  49614=>"010110010",
  49615=>"000000111",
  49616=>"111011101",
  49617=>"010101110",
  49618=>"000000100",
  49619=>"111111111",
  49620=>"101001100",
  49621=>"110100000",
  49622=>"101110011",
  49623=>"100010001",
  49624=>"111101100",
  49625=>"101111001",
  49626=>"011011101",
  49627=>"110101110",
  49628=>"000010010",
  49629=>"001011111",
  49630=>"100111110",
  49631=>"101111101",
  49632=>"100110111",
  49633=>"111011001",
  49634=>"010011100",
  49635=>"100011111",
  49636=>"100111111",
  49637=>"011001110",
  49638=>"000100110",
  49639=>"001101001",
  49640=>"110010001",
  49641=>"101010001",
  49642=>"010001100",
  49643=>"100111011",
  49644=>"001100100",
  49645=>"110000011",
  49646=>"110101001",
  49647=>"101101011",
  49648=>"100101011",
  49649=>"010011000",
  49650=>"100101010",
  49651=>"011000000",
  49652=>"100011011",
  49653=>"000101010",
  49654=>"001011000",
  49655=>"001100111",
  49656=>"101011110",
  49657=>"000000010",
  49658=>"001100010",
  49659=>"110000101",
  49660=>"110101011",
  49661=>"111001101",
  49662=>"001010101",
  49663=>"110110110",
  49664=>"111001100",
  49665=>"000011000",
  49666=>"111000010",
  49667=>"001000001",
  49668=>"000011000",
  49669=>"100010100",
  49670=>"110111001",
  49671=>"111011001",
  49672=>"011001111",
  49673=>"110001111",
  49674=>"000011101",
  49675=>"001010001",
  49676=>"001011001",
  49677=>"011100100",
  49678=>"100010011",
  49679=>"100110100",
  49680=>"111000000",
  49681=>"111100010",
  49682=>"000101010",
  49683=>"000011001",
  49684=>"101011000",
  49685=>"100101001",
  49686=>"110111011",
  49687=>"111101110",
  49688=>"101110011",
  49689=>"010001100",
  49690=>"000001110",
  49691=>"100000100",
  49692=>"011100101",
  49693=>"101100010",
  49694=>"000101001",
  49695=>"001000000",
  49696=>"011001000",
  49697=>"110101010",
  49698=>"111101111",
  49699=>"110000101",
  49700=>"110110010",
  49701=>"110110001",
  49702=>"000101100",
  49703=>"000011011",
  49704=>"010111001",
  49705=>"010100000",
  49706=>"001010110",
  49707=>"011001100",
  49708=>"101011011",
  49709=>"010101000",
  49710=>"101111010",
  49711=>"001110010",
  49712=>"001111111",
  49713=>"100110000",
  49714=>"001110000",
  49715=>"001000010",
  49716=>"010000010",
  49717=>"100010100",
  49718=>"011001011",
  49719=>"001100101",
  49720=>"001101000",
  49721=>"001000000",
  49722=>"111011000",
  49723=>"101011101",
  49724=>"011001100",
  49725=>"110000100",
  49726=>"101000010",
  49727=>"101100110",
  49728=>"101100000",
  49729=>"100000011",
  49730=>"100100101",
  49731=>"110011000",
  49732=>"100111001",
  49733=>"100001100",
  49734=>"010000011",
  49735=>"100110010",
  49736=>"110000111",
  49737=>"111110101",
  49738=>"100000100",
  49739=>"001001110",
  49740=>"110001110",
  49741=>"011000001",
  49742=>"111101101",
  49743=>"111001000",
  49744=>"011100111",
  49745=>"011111011",
  49746=>"010000100",
  49747=>"011001110",
  49748=>"111111010",
  49749=>"001100011",
  49750=>"110111111",
  49751=>"001000110",
  49752=>"111100110",
  49753=>"001000000",
  49754=>"010001100",
  49755=>"111111111",
  49756=>"101011011",
  49757=>"010001101",
  49758=>"011101100",
  49759=>"110101111",
  49760=>"110100100",
  49761=>"110100111",
  49762=>"111001001",
  49763=>"010101010",
  49764=>"110100010",
  49765=>"100101100",
  49766=>"010001101",
  49767=>"101111111",
  49768=>"000000100",
  49769=>"010100000",
  49770=>"010001000",
  49771=>"101101010",
  49772=>"011011101",
  49773=>"001010111",
  49774=>"010000100",
  49775=>"101000110",
  49776=>"111010101",
  49777=>"111010011",
  49778=>"011101000",
  49779=>"011011100",
  49780=>"101101010",
  49781=>"010101110",
  49782=>"100100110",
  49783=>"001101111",
  49784=>"010110110",
  49785=>"100010100",
  49786=>"001001111",
  49787=>"101110000",
  49788=>"001010000",
  49789=>"111101100",
  49790=>"111010011",
  49791=>"010110101",
  49792=>"110000000",
  49793=>"100000110",
  49794=>"111100011",
  49795=>"000110111",
  49796=>"000001101",
  49797=>"000000000",
  49798=>"001001011",
  49799=>"010010001",
  49800=>"101000100",
  49801=>"100000111",
  49802=>"111101111",
  49803=>"000000010",
  49804=>"010110010",
  49805=>"111101010",
  49806=>"001000000",
  49807=>"000100101",
  49808=>"101100011",
  49809=>"101001100",
  49810=>"011100010",
  49811=>"000011001",
  49812=>"001101000",
  49813=>"101000110",
  49814=>"110111010",
  49815=>"110101001",
  49816=>"000010100",
  49817=>"110100100",
  49818=>"110110101",
  49819=>"111011001",
  49820=>"111011010",
  49821=>"001101010",
  49822=>"110000010",
  49823=>"111101100",
  49824=>"011110010",
  49825=>"101111001",
  49826=>"101100000",
  49827=>"111110010",
  49828=>"001100111",
  49829=>"100000001",
  49830=>"001110011",
  49831=>"001001001",
  49832=>"011011000",
  49833=>"000001101",
  49834=>"010001000",
  49835=>"111111011",
  49836=>"011001100",
  49837=>"101101011",
  49838=>"110011101",
  49839=>"101101010",
  49840=>"011011000",
  49841=>"000100001",
  49842=>"001000111",
  49843=>"000001000",
  49844=>"011011010",
  49845=>"011011100",
  49846=>"011101110",
  49847=>"111010101",
  49848=>"100111101",
  49849=>"111111111",
  49850=>"001001100",
  49851=>"100011101",
  49852=>"101011001",
  49853=>"011111101",
  49854=>"000110100",
  49855=>"111101110",
  49856=>"001000100",
  49857=>"011001101",
  49858=>"001001110",
  49859=>"101000101",
  49860=>"001001001",
  49861=>"111001001",
  49862=>"111110110",
  49863=>"111111100",
  49864=>"001000111",
  49865=>"011101000",
  49866=>"011010100",
  49867=>"000011001",
  49868=>"110101110",
  49869=>"010011000",
  49870=>"101111101",
  49871=>"000011010",
  49872=>"000100010",
  49873=>"000100000",
  49874=>"000001011",
  49875=>"000011000",
  49876=>"111101001",
  49877=>"110100000",
  49878=>"101001100",
  49879=>"000010000",
  49880=>"000100011",
  49881=>"001000000",
  49882=>"101001110",
  49883=>"000101101",
  49884=>"111011001",
  49885=>"000100000",
  49886=>"000000011",
  49887=>"111000100",
  49888=>"110100100",
  49889=>"101011011",
  49890=>"101011111",
  49891=>"110110001",
  49892=>"010011011",
  49893=>"101101100",
  49894=>"101010011",
  49895=>"001101010",
  49896=>"010011101",
  49897=>"110010010",
  49898=>"110000000",
  49899=>"100101001",
  49900=>"000111100",
  49901=>"011011010",
  49902=>"000100101",
  49903=>"010011111",
  49904=>"011011010",
  49905=>"011000110",
  49906=>"001111010",
  49907=>"000001111",
  49908=>"000000010",
  49909=>"000100101",
  49910=>"101010011",
  49911=>"010110101",
  49912=>"100110101",
  49913=>"011110101",
  49914=>"101000110",
  49915=>"010101000",
  49916=>"111011011",
  49917=>"011101110",
  49918=>"110011000",
  49919=>"000010000",
  49920=>"100101000",
  49921=>"011010010",
  49922=>"001100110",
  49923=>"000000100",
  49924=>"011111000",
  49925=>"010010101",
  49926=>"100110011",
  49927=>"100011000",
  49928=>"110001001",
  49929=>"100100000",
  49930=>"001010000",
  49931=>"101000101",
  49932=>"111011100",
  49933=>"010011010",
  49934=>"001011100",
  49935=>"010000001",
  49936=>"010011001",
  49937=>"001111000",
  49938=>"001001110",
  49939=>"100100010",
  49940=>"100011001",
  49941=>"111110110",
  49942=>"010000101",
  49943=>"101000000",
  49944=>"011001001",
  49945=>"000111100",
  49946=>"000110011",
  49947=>"110011101",
  49948=>"100111110",
  49949=>"001110100",
  49950=>"010000000",
  49951=>"001001001",
  49952=>"110001110",
  49953=>"000010110",
  49954=>"001101101",
  49955=>"111101101",
  49956=>"001010101",
  49957=>"110001101",
  49958=>"100001111",
  49959=>"000001000",
  49960=>"101011111",
  49961=>"010000101",
  49962=>"110111111",
  49963=>"000101110",
  49964=>"010001010",
  49965=>"101100001",
  49966=>"001010110",
  49967=>"000001110",
  49968=>"101000001",
  49969=>"001010100",
  49970=>"111000011",
  49971=>"011010110",
  49972=>"011101000",
  49973=>"100000110",
  49974=>"010111111",
  49975=>"000010011",
  49976=>"101100100",
  49977=>"101000000",
  49978=>"011101101",
  49979=>"110000010",
  49980=>"111001110",
  49981=>"010010000",
  49982=>"111010011",
  49983=>"110001110",
  49984=>"101111110",
  49985=>"101011100",
  49986=>"101010111",
  49987=>"010000010",
  49988=>"001001001",
  49989=>"001001101",
  49990=>"001000010",
  49991=>"101100111",
  49992=>"100010010",
  49993=>"001101010",
  49994=>"000101010",
  49995=>"110100111",
  49996=>"010111000",
  49997=>"010100100",
  49998=>"110111100",
  49999=>"001011100",
  50000=>"011110100",
  50001=>"000110111",
  50002=>"010111100",
  50003=>"110010000",
  50004=>"111110110",
  50005=>"101011111",
  50006=>"001110010",
  50007=>"011010101",
  50008=>"011011111",
  50009=>"111000111",
  50010=>"100100110",
  50011=>"110010110",
  50012=>"111111011",
  50013=>"111101101",
  50014=>"011000111",
  50015=>"001001000",
  50016=>"001111000",
  50017=>"010010101",
  50018=>"101110101",
  50019=>"001111101",
  50020=>"111111011",
  50021=>"000000101",
  50022=>"011000101",
  50023=>"100011011",
  50024=>"101000001",
  50025=>"100111110",
  50026=>"111111111",
  50027=>"011111110",
  50028=>"100101100",
  50029=>"101110001",
  50030=>"000000110",
  50031=>"001001111",
  50032=>"101001110",
  50033=>"100011001",
  50034=>"101101011",
  50035=>"011001110",
  50036=>"100110000",
  50037=>"011100001",
  50038=>"111101111",
  50039=>"111000010",
  50040=>"000010101",
  50041=>"001100111",
  50042=>"110001011",
  50043=>"011001110",
  50044=>"001000100",
  50045=>"000011001",
  50046=>"100100011",
  50047=>"100111110",
  50048=>"110011100",
  50049=>"100100011",
  50050=>"000111011",
  50051=>"100101011",
  50052=>"101010010",
  50053=>"010101000",
  50054=>"101000101",
  50055=>"010101100",
  50056=>"111011010",
  50057=>"011011011",
  50058=>"011100111",
  50059=>"011000000",
  50060=>"011111010",
  50061=>"111111111",
  50062=>"001110101",
  50063=>"110010100",
  50064=>"001101100",
  50065=>"000001010",
  50066=>"100111001",
  50067=>"101110111",
  50068=>"000010010",
  50069=>"010010110",
  50070=>"100000000",
  50071=>"110011111",
  50072=>"100000010",
  50073=>"000010101",
  50074=>"010001100",
  50075=>"110110011",
  50076=>"110101010",
  50077=>"001001010",
  50078=>"100010111",
  50079=>"011101001",
  50080=>"111111011",
  50081=>"111110010",
  50082=>"011111011",
  50083=>"011110101",
  50084=>"100101110",
  50085=>"100111111",
  50086=>"101000010",
  50087=>"001010010",
  50088=>"000000110",
  50089=>"101010011",
  50090=>"010001101",
  50091=>"111011001",
  50092=>"000111011",
  50093=>"010000000",
  50094=>"001100001",
  50095=>"000010100",
  50096=>"001000011",
  50097=>"010110001",
  50098=>"111110111",
  50099=>"010001001",
  50100=>"110101000",
  50101=>"110001011",
  50102=>"011110100",
  50103=>"010010001",
  50104=>"101110001",
  50105=>"101100010",
  50106=>"011000100",
  50107=>"011111111",
  50108=>"101001100",
  50109=>"111010100",
  50110=>"111000110",
  50111=>"111001000",
  50112=>"000010111",
  50113=>"001111111",
  50114=>"111100101",
  50115=>"111111110",
  50116=>"110010100",
  50117=>"111010111",
  50118=>"000111111",
  50119=>"101011001",
  50120=>"100111000",
  50121=>"111000011",
  50122=>"011101011",
  50123=>"101110111",
  50124=>"101011000",
  50125=>"011010101",
  50126=>"111001011",
  50127=>"000001001",
  50128=>"001000011",
  50129=>"100111001",
  50130=>"001100000",
  50131=>"010001100",
  50132=>"010001010",
  50133=>"011100110",
  50134=>"101011100",
  50135=>"101000001",
  50136=>"110010010",
  50137=>"001100000",
  50138=>"100010010",
  50139=>"101010001",
  50140=>"001011001",
  50141=>"000000100",
  50142=>"011000000",
  50143=>"110111000",
  50144=>"111111100",
  50145=>"000000011",
  50146=>"000111111",
  50147=>"011010000",
  50148=>"001001001",
  50149=>"011010000",
  50150=>"111000000",
  50151=>"100100011",
  50152=>"110101101",
  50153=>"100111011",
  50154=>"101100000",
  50155=>"111011010",
  50156=>"101101111",
  50157=>"000000001",
  50158=>"100111111",
  50159=>"100011111",
  50160=>"100111111",
  50161=>"101100011",
  50162=>"011001101",
  50163=>"000101011",
  50164=>"100101011",
  50165=>"001000100",
  50166=>"111011111",
  50167=>"000111001",
  50168=>"111101001",
  50169=>"001110010",
  50170=>"110110111",
  50171=>"110111001",
  50172=>"000000111",
  50173=>"001010000",
  50174=>"100010101",
  50175=>"101111010",
  50176=>"000000011",
  50177=>"000101111",
  50178=>"011110001",
  50179=>"011011010",
  50180=>"100000100",
  50181=>"100001100",
  50182=>"001000111",
  50183=>"001111101",
  50184=>"111010000",
  50185=>"010001100",
  50186=>"010000110",
  50187=>"111001011",
  50188=>"001101001",
  50189=>"000000100",
  50190=>"100001100",
  50191=>"111011000",
  50192=>"010111000",
  50193=>"011111010",
  50194=>"011011011",
  50195=>"011010110",
  50196=>"010101000",
  50197=>"001000010",
  50198=>"111110101",
  50199=>"010000000",
  50200=>"100101111",
  50201=>"000100000",
  50202=>"000100001",
  50203=>"011001100",
  50204=>"011011110",
  50205=>"110111101",
  50206=>"010111000",
  50207=>"010000000",
  50208=>"101010001",
  50209=>"100101100",
  50210=>"000110000",
  50211=>"101111011",
  50212=>"001100101",
  50213=>"011100101",
  50214=>"001011001",
  50215=>"011110111",
  50216=>"111101011",
  50217=>"010110101",
  50218=>"000011000",
  50219=>"010111101",
  50220=>"000000010",
  50221=>"000011101",
  50222=>"001111110",
  50223=>"101000111",
  50224=>"111101111",
  50225=>"101010011",
  50226=>"100001010",
  50227=>"001011110",
  50228=>"101000111",
  50229=>"010111011",
  50230=>"011001001",
  50231=>"010001001",
  50232=>"000011000",
  50233=>"000000110",
  50234=>"111011101",
  50235=>"000111011",
  50236=>"000100010",
  50237=>"001101011",
  50238=>"001000000",
  50239=>"010100001",
  50240=>"000111100",
  50241=>"010110110",
  50242=>"110111100",
  50243=>"001101010",
  50244=>"100000000",
  50245=>"101101111",
  50246=>"111011101",
  50247=>"100101000",
  50248=>"110101101",
  50249=>"101100001",
  50250=>"001110000",
  50251=>"011000111",
  50252=>"000000100",
  50253=>"011111110",
  50254=>"111001001",
  50255=>"111100000",
  50256=>"001000001",
  50257=>"111010101",
  50258=>"111011101",
  50259=>"100110001",
  50260=>"000000101",
  50261=>"001010101",
  50262=>"000101010",
  50263=>"100101100",
  50264=>"111011001",
  50265=>"111110110",
  50266=>"000000100",
  50267=>"110110000",
  50268=>"011100101",
  50269=>"110100010",
  50270=>"110100111",
  50271=>"101000111",
  50272=>"110100100",
  50273=>"110001100",
  50274=>"010110100",
  50275=>"010011000",
  50276=>"000100011",
  50277=>"110010000",
  50278=>"000011001",
  50279=>"000011101",
  50280=>"111100101",
  50281=>"010011001",
  50282=>"010110011",
  50283=>"110001110",
  50284=>"001010110",
  50285=>"111010010",
  50286=>"110001010",
  50287=>"010011000",
  50288=>"000101001",
  50289=>"011100111",
  50290=>"110000000",
  50291=>"011100110",
  50292=>"111110001",
  50293=>"110000100",
  50294=>"111100110",
  50295=>"110011011",
  50296=>"111000001",
  50297=>"100100010",
  50298=>"100100110",
  50299=>"111000011",
  50300=>"101000000",
  50301=>"110000110",
  50302=>"110100010",
  50303=>"100010001",
  50304=>"010101110",
  50305=>"010111111",
  50306=>"100000000",
  50307=>"000111010",
  50308=>"000010001",
  50309=>"000000010",
  50310=>"101101101",
  50311=>"100100001",
  50312=>"110011101",
  50313=>"100000001",
  50314=>"001110110",
  50315=>"001000011",
  50316=>"111110111",
  50317=>"001101001",
  50318=>"110000101",
  50319=>"010100111",
  50320=>"111010000",
  50321=>"011110010",
  50322=>"000000000",
  50323=>"000010001",
  50324=>"110100111",
  50325=>"100011110",
  50326=>"001100010",
  50327=>"000110010",
  50328=>"000000011",
  50329=>"001100100",
  50330=>"000100000",
  50331=>"001010010",
  50332=>"101100101",
  50333=>"110000000",
  50334=>"101100111",
  50335=>"000011000",
  50336=>"100100111",
  50337=>"111011001",
  50338=>"001001101",
  50339=>"011000110",
  50340=>"011100010",
  50341=>"001100111",
  50342=>"001100000",
  50343=>"100101110",
  50344=>"100101001",
  50345=>"111101010",
  50346=>"100110001",
  50347=>"111111000",
  50348=>"111110000",
  50349=>"111000001",
  50350=>"100011100",
  50351=>"011001110",
  50352=>"000010010",
  50353=>"001100000",
  50354=>"101010100",
  50355=>"010000100",
  50356=>"010010010",
  50357=>"011011111",
  50358=>"111011101",
  50359=>"110011000",
  50360=>"100010001",
  50361=>"011110000",
  50362=>"010110100",
  50363=>"111100011",
  50364=>"001001111",
  50365=>"101101011",
  50366=>"001110010",
  50367=>"010001000",
  50368=>"101011011",
  50369=>"011000010",
  50370=>"000101011",
  50371=>"110000111",
  50372=>"111010010",
  50373=>"011101100",
  50374=>"101100101",
  50375=>"000101001",
  50376=>"011001011",
  50377=>"011110011",
  50378=>"100010100",
  50379=>"111111001",
  50380=>"111001010",
  50381=>"001010011",
  50382=>"111011000",
  50383=>"101100000",
  50384=>"010100001",
  50385=>"111000011",
  50386=>"000100000",
  50387=>"111101011",
  50388=>"000110111",
  50389=>"010101100",
  50390=>"000010010",
  50391=>"111110011",
  50392=>"011011011",
  50393=>"011010000",
  50394=>"011011111",
  50395=>"101010100",
  50396=>"001010000",
  50397=>"001111101",
  50398=>"011001111",
  50399=>"011010101",
  50400=>"001001000",
  50401=>"011100101",
  50402=>"000001111",
  50403=>"101110001",
  50404=>"010111011",
  50405=>"000110110",
  50406=>"101100111",
  50407=>"100001011",
  50408=>"010000001",
  50409=>"001010010",
  50410=>"000010100",
  50411=>"110000000",
  50412=>"100101010",
  50413=>"000110001",
  50414=>"011101101",
  50415=>"111000101",
  50416=>"000011010",
  50417=>"111000111",
  50418=>"110011010",
  50419=>"110001100",
  50420=>"000101000",
  50421=>"101111100",
  50422=>"110001010",
  50423=>"010101101",
  50424=>"101100111",
  50425=>"010000001",
  50426=>"010010101",
  50427=>"001010000",
  50428=>"000001010",
  50429=>"000000111",
  50430=>"110010001",
  50431=>"010111011",
  50432=>"100011010",
  50433=>"001001011",
  50434=>"011000111",
  50435=>"010011110",
  50436=>"001010011",
  50437=>"100000010",
  50438=>"010110000",
  50439=>"110000000",
  50440=>"000000010",
  50441=>"110000010",
  50442=>"100110110",
  50443=>"011100101",
  50444=>"111011111",
  50445=>"100101111",
  50446=>"110001111",
  50447=>"100010001",
  50448=>"111110000",
  50449=>"100001100",
  50450=>"011000011",
  50451=>"100111111",
  50452=>"101101101",
  50453=>"100001110",
  50454=>"100100110",
  50455=>"101000101",
  50456=>"101101100",
  50457=>"010110000",
  50458=>"100001101",
  50459=>"001110000",
  50460=>"100011011",
  50461=>"010100100",
  50462=>"001011000",
  50463=>"010001110",
  50464=>"001011010",
  50465=>"000111010",
  50466=>"001101010",
  50467=>"101010010",
  50468=>"010001100",
  50469=>"010000111",
  50470=>"100011000",
  50471=>"110010000",
  50472=>"110000010",
  50473=>"010010110",
  50474=>"011110110",
  50475=>"100000101",
  50476=>"001110111",
  50477=>"001010100",
  50478=>"001011001",
  50479=>"100100110",
  50480=>"111100001",
  50481=>"101101111",
  50482=>"110110101",
  50483=>"010010000",
  50484=>"111011010",
  50485=>"001000000",
  50486=>"011100000",
  50487=>"011101011",
  50488=>"010000100",
  50489=>"101011011",
  50490=>"110101000",
  50491=>"111011000",
  50492=>"001100010",
  50493=>"101111110",
  50494=>"110101101",
  50495=>"011100111",
  50496=>"101101111",
  50497=>"001011010",
  50498=>"000100100",
  50499=>"000001101",
  50500=>"010001011",
  50501=>"100101000",
  50502=>"001000100",
  50503=>"000010010",
  50504=>"011111100",
  50505=>"111111000",
  50506=>"001110011",
  50507=>"001101101",
  50508=>"101010110",
  50509=>"011100101",
  50510=>"000011010",
  50511=>"011101110",
  50512=>"101011110",
  50513=>"100111001",
  50514=>"100010001",
  50515=>"010010110",
  50516=>"001001110",
  50517=>"111110001",
  50518=>"111110101",
  50519=>"001110000",
  50520=>"100011011",
  50521=>"001110110",
  50522=>"100110010",
  50523=>"110110100",
  50524=>"110010010",
  50525=>"001100001",
  50526=>"111111010",
  50527=>"101000010",
  50528=>"111101101",
  50529=>"111100010",
  50530=>"110011011",
  50531=>"100110110",
  50532=>"001001001",
  50533=>"101001110",
  50534=>"010010100",
  50535=>"111000111",
  50536=>"101100010",
  50537=>"001101000",
  50538=>"011110111",
  50539=>"011100110",
  50540=>"100010001",
  50541=>"100011101",
  50542=>"000001000",
  50543=>"011110110",
  50544=>"110011000",
  50545=>"110101011",
  50546=>"011011000",
  50547=>"100110100",
  50548=>"110011010",
  50549=>"000101111",
  50550=>"110000011",
  50551=>"110111101",
  50552=>"111111010",
  50553=>"010001000",
  50554=>"010000001",
  50555=>"000001101",
  50556=>"100011011",
  50557=>"000111110",
  50558=>"101111101",
  50559=>"101100010",
  50560=>"111110001",
  50561=>"101011111",
  50562=>"011011001",
  50563=>"000101011",
  50564=>"110010110",
  50565=>"111000010",
  50566=>"000101011",
  50567=>"000100101",
  50568=>"001011100",
  50569=>"110101101",
  50570=>"000101001",
  50571=>"010000000",
  50572=>"100010000",
  50573=>"010001111",
  50574=>"011101000",
  50575=>"110110111",
  50576=>"001111011",
  50577=>"001000000",
  50578=>"011000001",
  50579=>"101111100",
  50580=>"010011100",
  50581=>"001100000",
  50582=>"111111000",
  50583=>"111110000",
  50584=>"110101010",
  50585=>"101001010",
  50586=>"110001101",
  50587=>"101011110",
  50588=>"001110101",
  50589=>"000001100",
  50590=>"100110101",
  50591=>"111111000",
  50592=>"111000011",
  50593=>"010000100",
  50594=>"010001111",
  50595=>"000000100",
  50596=>"010101100",
  50597=>"111101011",
  50598=>"111000100",
  50599=>"001101111",
  50600=>"111011110",
  50601=>"011011000",
  50602=>"000100011",
  50603=>"011100100",
  50604=>"111101100",
  50605=>"001101001",
  50606=>"101110001",
  50607=>"101101010",
  50608=>"010001010",
  50609=>"111101110",
  50610=>"110111111",
  50611=>"011100010",
  50612=>"110001110",
  50613=>"001001110",
  50614=>"000101011",
  50615=>"110100100",
  50616=>"101101100",
  50617=>"110000101",
  50618=>"101000111",
  50619=>"110001000",
  50620=>"010000000",
  50621=>"000111011",
  50622=>"111000100",
  50623=>"010100000",
  50624=>"011010111",
  50625=>"101010100",
  50626=>"011100101",
  50627=>"001111111",
  50628=>"110000010",
  50629=>"011110001",
  50630=>"001000011",
  50631=>"101100011",
  50632=>"110001101",
  50633=>"110100100",
  50634=>"101100010",
  50635=>"110010110",
  50636=>"001000001",
  50637=>"110010111",
  50638=>"111011010",
  50639=>"100010101",
  50640=>"011101110",
  50641=>"001001010",
  50642=>"010001101",
  50643=>"101100001",
  50644=>"000111010",
  50645=>"101001011",
  50646=>"100000000",
  50647=>"110011000",
  50648=>"010001011",
  50649=>"111110000",
  50650=>"110101111",
  50651=>"101000011",
  50652=>"101101110",
  50653=>"111101010",
  50654=>"011110111",
  50655=>"011011111",
  50656=>"011110001",
  50657=>"011011110",
  50658=>"000100111",
  50659=>"100000011",
  50660=>"001000000",
  50661=>"101001100",
  50662=>"001001000",
  50663=>"101001000",
  50664=>"010010011",
  50665=>"101010010",
  50666=>"101000100",
  50667=>"101100010",
  50668=>"110010000",
  50669=>"100001000",
  50670=>"000110110",
  50671=>"010000011",
  50672=>"110010110",
  50673=>"010111000",
  50674=>"110100001",
  50675=>"011011010",
  50676=>"011111100",
  50677=>"000100101",
  50678=>"001100110",
  50679=>"010011000",
  50680=>"100111000",
  50681=>"001001000",
  50682=>"111010000",
  50683=>"001010111",
  50684=>"110001100",
  50685=>"010010010",
  50686=>"010111100",
  50687=>"101111101",
  50688=>"000111000",
  50689=>"001111111",
  50690=>"011101011",
  50691=>"011100110",
  50692=>"111011001",
  50693=>"001110000",
  50694=>"010010100",
  50695=>"001000110",
  50696=>"111110111",
  50697=>"001101110",
  50698=>"110011101",
  50699=>"011111000",
  50700=>"100010011",
  50701=>"111111011",
  50702=>"111000000",
  50703=>"110010111",
  50704=>"001011111",
  50705=>"110000110",
  50706=>"011011100",
  50707=>"000000100",
  50708=>"101011100",
  50709=>"101001100",
  50710=>"001001110",
  50711=>"101011100",
  50712=>"111111110",
  50713=>"110000011",
  50714=>"000000010",
  50715=>"110000101",
  50716=>"001000101",
  50717=>"011100101",
  50718=>"000000100",
  50719=>"101101011",
  50720=>"100101001",
  50721=>"110101000",
  50722=>"001101010",
  50723=>"111010100",
  50724=>"111101001",
  50725=>"000010101",
  50726=>"100110011",
  50727=>"000110011",
  50728=>"111110101",
  50729=>"001010011",
  50730=>"111001001",
  50731=>"010110101",
  50732=>"100110010",
  50733=>"011001110",
  50734=>"111000101",
  50735=>"100110111",
  50736=>"010100111",
  50737=>"011100011",
  50738=>"000000010",
  50739=>"000001110",
  50740=>"001111100",
  50741=>"011100010",
  50742=>"000001011",
  50743=>"111011111",
  50744=>"100110110",
  50745=>"110010000",
  50746=>"000001000",
  50747=>"101110101",
  50748=>"100011010",
  50749=>"000111001",
  50750=>"000100110",
  50751=>"111100110",
  50752=>"010101000",
  50753=>"100101101",
  50754=>"101110011",
  50755=>"100010110",
  50756=>"011111001",
  50757=>"011111011",
  50758=>"101110001",
  50759=>"100010100",
  50760=>"111011010",
  50761=>"000000111",
  50762=>"110111010",
  50763=>"101000101",
  50764=>"010111111",
  50765=>"100110111",
  50766=>"101110000",
  50767=>"110111010",
  50768=>"101110110",
  50769=>"001011101",
  50770=>"111001000",
  50771=>"000010000",
  50772=>"111000100",
  50773=>"101100000",
  50774=>"111001010",
  50775=>"100010011",
  50776=>"010111000",
  50777=>"011111001",
  50778=>"110011100",
  50779=>"000010000",
  50780=>"000100000",
  50781=>"100100010",
  50782=>"000111010",
  50783=>"101110111",
  50784=>"111110001",
  50785=>"100001010",
  50786=>"100101111",
  50787=>"001001000",
  50788=>"111000010",
  50789=>"010101001",
  50790=>"101110110",
  50791=>"000111110",
  50792=>"001011100",
  50793=>"000001100",
  50794=>"010011010",
  50795=>"101000111",
  50796=>"010001000",
  50797=>"100001001",
  50798=>"110111110",
  50799=>"110101101",
  50800=>"001000000",
  50801=>"001101000",
  50802=>"111110100",
  50803=>"111000000",
  50804=>"011101110",
  50805=>"010111010",
  50806=>"011110000",
  50807=>"001001101",
  50808=>"111100011",
  50809=>"100011101",
  50810=>"101011000",
  50811=>"110110010",
  50812=>"010001000",
  50813=>"010010111",
  50814=>"111111101",
  50815=>"010101010",
  50816=>"000010110",
  50817=>"010101101",
  50818=>"100011011",
  50819=>"101000011",
  50820=>"001000000",
  50821=>"000111101",
  50822=>"101100001",
  50823=>"010001101",
  50824=>"110000100",
  50825=>"000100001",
  50826=>"110010010",
  50827=>"111011111",
  50828=>"111101000",
  50829=>"111100100",
  50830=>"001011000",
  50831=>"010110111",
  50832=>"011010010",
  50833=>"000011011",
  50834=>"110110011",
  50835=>"100000110",
  50836=>"011001100",
  50837=>"110111110",
  50838=>"110010110",
  50839=>"010000110",
  50840=>"110001011",
  50841=>"000111101",
  50842=>"100000000",
  50843=>"100011011",
  50844=>"000101111",
  50845=>"110000100",
  50846=>"011011010",
  50847=>"001101000",
  50848=>"000010101",
  50849=>"110010001",
  50850=>"011111110",
  50851=>"000110100",
  50852=>"010111001",
  50853=>"000010000",
  50854=>"101100101",
  50855=>"100111111",
  50856=>"111100101",
  50857=>"000000111",
  50858=>"101100110",
  50859=>"110010000",
  50860=>"001011000",
  50861=>"101000000",
  50862=>"100100101",
  50863=>"110001011",
  50864=>"111100111",
  50865=>"100010110",
  50866=>"111111001",
  50867=>"001011010",
  50868=>"100100110",
  50869=>"010001001",
  50870=>"011111000",
  50871=>"010011111",
  50872=>"101010011",
  50873=>"001100000",
  50874=>"100000110",
  50875=>"100101010",
  50876=>"010010111",
  50877=>"001000101",
  50878=>"000011010",
  50879=>"001001001",
  50880=>"101110011",
  50881=>"110110011",
  50882=>"100001011",
  50883=>"000011100",
  50884=>"110001111",
  50885=>"010010100",
  50886=>"110110110",
  50887=>"000000111",
  50888=>"111011101",
  50889=>"011100010",
  50890=>"001001111",
  50891=>"001100010",
  50892=>"011110110",
  50893=>"101001000",
  50894=>"100001101",
  50895=>"010011011",
  50896=>"001001000",
  50897=>"000010000",
  50898=>"000100000",
  50899=>"001011100",
  50900=>"101101101",
  50901=>"011110000",
  50902=>"011010011",
  50903=>"000011110",
  50904=>"100110001",
  50905=>"111110101",
  50906=>"111100110",
  50907=>"001100010",
  50908=>"101001101",
  50909=>"110100011",
  50910=>"110101110",
  50911=>"101111000",
  50912=>"011011000",
  50913=>"110001010",
  50914=>"101100101",
  50915=>"101111111",
  50916=>"110111100",
  50917=>"000100101",
  50918=>"111000001",
  50919=>"100010010",
  50920=>"100011000",
  50921=>"111110010",
  50922=>"001101001",
  50923=>"110110010",
  50924=>"110110000",
  50925=>"000111010",
  50926=>"011100111",
  50927=>"000010111",
  50928=>"110000010",
  50929=>"000000101",
  50930=>"101101101",
  50931=>"110111111",
  50932=>"011011101",
  50933=>"100000110",
  50934=>"001001010",
  50935=>"001000110",
  50936=>"000001011",
  50937=>"111100100",
  50938=>"001100001",
  50939=>"000111111",
  50940=>"100111011",
  50941=>"010010000",
  50942=>"010000011",
  50943=>"011100011",
  50944=>"111110100",
  50945=>"001111111",
  50946=>"000111101",
  50947=>"100110000",
  50948=>"100101100",
  50949=>"000000100",
  50950=>"100101010",
  50951=>"000011010",
  50952=>"001001000",
  50953=>"110101000",
  50954=>"101001111",
  50955=>"001000000",
  50956=>"111111100",
  50957=>"110111111",
  50958=>"001001000",
  50959=>"101010111",
  50960=>"110111001",
  50961=>"110000011",
  50962=>"101111001",
  50963=>"101110011",
  50964=>"000001110",
  50965=>"110010010",
  50966=>"001001110",
  50967=>"011110101",
  50968=>"110100101",
  50969=>"010100001",
  50970=>"000000000",
  50971=>"101101101",
  50972=>"001101011",
  50973=>"000101011",
  50974=>"110011001",
  50975=>"110010011",
  50976=>"110001011",
  50977=>"000110000",
  50978=>"101110101",
  50979=>"000110100",
  50980=>"010110010",
  50981=>"110100100",
  50982=>"000001010",
  50983=>"111100101",
  50984=>"000011001",
  50985=>"000010011",
  50986=>"101010111",
  50987=>"110011111",
  50988=>"001011000",
  50989=>"000001101",
  50990=>"010000011",
  50991=>"101011010",
  50992=>"000001000",
  50993=>"000000011",
  50994=>"111010001",
  50995=>"101001101",
  50996=>"110111011",
  50997=>"001011110",
  50998=>"110100011",
  50999=>"101001010",
  51000=>"101010110",
  51001=>"000100100",
  51002=>"010001001",
  51003=>"001101110",
  51004=>"101110000",
  51005=>"000010100",
  51006=>"011100110",
  51007=>"000011101",
  51008=>"011111001",
  51009=>"011001000",
  51010=>"011010100",
  51011=>"101100111",
  51012=>"011101110",
  51013=>"110101001",
  51014=>"100100111",
  51015=>"000000010",
  51016=>"011000111",
  51017=>"001010011",
  51018=>"000111000",
  51019=>"000011101",
  51020=>"001111101",
  51021=>"101111001",
  51022=>"101100110",
  51023=>"111010010",
  51024=>"110100011",
  51025=>"010111100",
  51026=>"001111001",
  51027=>"101100110",
  51028=>"100111111",
  51029=>"001010011",
  51030=>"100001011",
  51031=>"010101000",
  51032=>"011101011",
  51033=>"111110110",
  51034=>"011100001",
  51035=>"001001110",
  51036=>"101011000",
  51037=>"101101101",
  51038=>"000110111",
  51039=>"100000000",
  51040=>"011001010",
  51041=>"110110111",
  51042=>"011101010",
  51043=>"100001110",
  51044=>"111101010",
  51045=>"000010011",
  51046=>"010111010",
  51047=>"001011011",
  51048=>"011101011",
  51049=>"111010101",
  51050=>"110100000",
  51051=>"111111100",
  51052=>"001011100",
  51053=>"010100000",
  51054=>"110110101",
  51055=>"110111101",
  51056=>"001101111",
  51057=>"011001100",
  51058=>"101111010",
  51059=>"011101111",
  51060=>"011111110",
  51061=>"001001001",
  51062=>"111110001",
  51063=>"101110110",
  51064=>"000011000",
  51065=>"011100110",
  51066=>"011011101",
  51067=>"010001110",
  51068=>"001000100",
  51069=>"011001000",
  51070=>"100101110",
  51071=>"010100100",
  51072=>"100010010",
  51073=>"100010001",
  51074=>"000110101",
  51075=>"100101000",
  51076=>"000000110",
  51077=>"001011100",
  51078=>"100001110",
  51079=>"101000011",
  51080=>"111111111",
  51081=>"110000111",
  51082=>"100101111",
  51083=>"011010110",
  51084=>"100011000",
  51085=>"111001011",
  51086=>"100110000",
  51087=>"110000011",
  51088=>"011011111",
  51089=>"101100110",
  51090=>"000100100",
  51091=>"011011110",
  51092=>"101110010",
  51093=>"010111110",
  51094=>"000010111",
  51095=>"111100100",
  51096=>"111000011",
  51097=>"001011111",
  51098=>"010101100",
  51099=>"101100100",
  51100=>"100100010",
  51101=>"000101000",
  51102=>"000001001",
  51103=>"011110101",
  51104=>"011000001",
  51105=>"000110011",
  51106=>"011001001",
  51107=>"100100100",
  51108=>"110101110",
  51109=>"010100100",
  51110=>"110010011",
  51111=>"010111000",
  51112=>"101101000",
  51113=>"001111001",
  51114=>"111010110",
  51115=>"010000001",
  51116=>"100010000",
  51117=>"101100010",
  51118=>"101011001",
  51119=>"100101100",
  51120=>"011101000",
  51121=>"011111011",
  51122=>"111110111",
  51123=>"011110011",
  51124=>"001110001",
  51125=>"000100100",
  51126=>"111000000",
  51127=>"111011100",
  51128=>"001101010",
  51129=>"010100011",
  51130=>"101010010",
  51131=>"110010111",
  51132=>"101100001",
  51133=>"011001100",
  51134=>"110100010",
  51135=>"111001000",
  51136=>"100110010",
  51137=>"011100001",
  51138=>"101100111",
  51139=>"100001010",
  51140=>"111010010",
  51141=>"000011011",
  51142=>"001011010",
  51143=>"000111100",
  51144=>"100011100",
  51145=>"001000011",
  51146=>"000001011",
  51147=>"111100111",
  51148=>"001111110",
  51149=>"000100011",
  51150=>"000100110",
  51151=>"110000001",
  51152=>"101001000",
  51153=>"000000101",
  51154=>"111000000",
  51155=>"011001011",
  51156=>"101010111",
  51157=>"111001101",
  51158=>"010100001",
  51159=>"111101111",
  51160=>"010101110",
  51161=>"110010100",
  51162=>"101001101",
  51163=>"001101010",
  51164=>"000011100",
  51165=>"110011100",
  51166=>"101011110",
  51167=>"001000001",
  51168=>"100001101",
  51169=>"101011111",
  51170=>"010000001",
  51171=>"010010000",
  51172=>"001110011",
  51173=>"011011000",
  51174=>"000110100",
  51175=>"000100000",
  51176=>"110000000",
  51177=>"111011110",
  51178=>"001001100",
  51179=>"111000010",
  51180=>"101001001",
  51181=>"110011100",
  51182=>"110000101",
  51183=>"010101011",
  51184=>"110010100",
  51185=>"110110101",
  51186=>"101000111",
  51187=>"110010100",
  51188=>"010000101",
  51189=>"110110000",
  51190=>"000110111",
  51191=>"100100111",
  51192=>"011111000",
  51193=>"001111100",
  51194=>"011010011",
  51195=>"011110111",
  51196=>"111000110",
  51197=>"111111110",
  51198=>"001101000",
  51199=>"001010001",
  51200=>"110110010",
  51201=>"010110111",
  51202=>"000010110",
  51203=>"110110000",
  51204=>"011110101",
  51205=>"001101100",
  51206=>"000111111",
  51207=>"011010101",
  51208=>"000000100",
  51209=>"011100011",
  51210=>"101010101",
  51211=>"100100001",
  51212=>"111001100",
  51213=>"101000000",
  51214=>"100000100",
  51215=>"001111111",
  51216=>"011110000",
  51217=>"001101001",
  51218=>"111010101",
  51219=>"001111101",
  51220=>"100111110",
  51221=>"010001011",
  51222=>"000010011",
  51223=>"101100100",
  51224=>"011001010",
  51225=>"011010001",
  51226=>"100111101",
  51227=>"101001011",
  51228=>"111110001",
  51229=>"100010110",
  51230=>"001100100",
  51231=>"101000010",
  51232=>"001101111",
  51233=>"110001011",
  51234=>"011100010",
  51235=>"100011101",
  51236=>"110010010",
  51237=>"000101010",
  51238=>"100000001",
  51239=>"110111010",
  51240=>"100100101",
  51241=>"101000000",
  51242=>"110110101",
  51243=>"000110001",
  51244=>"100110110",
  51245=>"101110010",
  51246=>"001010111",
  51247=>"100010110",
  51248=>"100010111",
  51249=>"010000100",
  51250=>"111101111",
  51251=>"000000100",
  51252=>"110000100",
  51253=>"100110111",
  51254=>"110111100",
  51255=>"010010110",
  51256=>"001101001",
  51257=>"000111011",
  51258=>"001110111",
  51259=>"101010100",
  51260=>"111011001",
  51261=>"111001100",
  51262=>"000011010",
  51263=>"001110000",
  51264=>"010001001",
  51265=>"000010100",
  51266=>"000111011",
  51267=>"101000001",
  51268=>"110011000",
  51269=>"011100101",
  51270=>"011010111",
  51271=>"000010111",
  51272=>"010101010",
  51273=>"100110101",
  51274=>"110000011",
  51275=>"000000101",
  51276=>"000110010",
  51277=>"000010010",
  51278=>"100110001",
  51279=>"010000111",
  51280=>"100101000",
  51281=>"010010000",
  51282=>"110000100",
  51283=>"110000001",
  51284=>"100011001",
  51285=>"101100000",
  51286=>"100101010",
  51287=>"011010011",
  51288=>"001100001",
  51289=>"111101101",
  51290=>"001110010",
  51291=>"010110101",
  51292=>"011101100",
  51293=>"010001101",
  51294=>"011000001",
  51295=>"110011110",
  51296=>"111110011",
  51297=>"000001011",
  51298=>"101011000",
  51299=>"001010010",
  51300=>"010101100",
  51301=>"110000000",
  51302=>"111101111",
  51303=>"011110100",
  51304=>"011000011",
  51305=>"111001100",
  51306=>"111000111",
  51307=>"000101100",
  51308=>"010100101",
  51309=>"111101011",
  51310=>"101110110",
  51311=>"101010000",
  51312=>"101011111",
  51313=>"101011011",
  51314=>"010011101",
  51315=>"110000110",
  51316=>"111101011",
  51317=>"010110000",
  51318=>"010110111",
  51319=>"000001010",
  51320=>"001011100",
  51321=>"010010111",
  51322=>"101001011",
  51323=>"001000001",
  51324=>"110011100",
  51325=>"111101110",
  51326=>"001011000",
  51327=>"000100001",
  51328=>"101000101",
  51329=>"000111111",
  51330=>"111011011",
  51331=>"010111010",
  51332=>"100101000",
  51333=>"110011011",
  51334=>"100110100",
  51335=>"111000100",
  51336=>"100000010",
  51337=>"111010000",
  51338=>"000100111",
  51339=>"011100000",
  51340=>"001100001",
  51341=>"010101001",
  51342=>"011010110",
  51343=>"111001000",
  51344=>"011110001",
  51345=>"011110010",
  51346=>"011111011",
  51347=>"000000101",
  51348=>"001111100",
  51349=>"000011000",
  51350=>"011110100",
  51351=>"110001000",
  51352=>"100011001",
  51353=>"110111101",
  51354=>"101001011",
  51355=>"000101100",
  51356=>"101100100",
  51357=>"111100011",
  51358=>"010000001",
  51359=>"001000010",
  51360=>"110101110",
  51361=>"001101100",
  51362=>"011110100",
  51363=>"100110111",
  51364=>"101011000",
  51365=>"010000100",
  51366=>"100011110",
  51367=>"111000111",
  51368=>"001101000",
  51369=>"100110100",
  51370=>"010000011",
  51371=>"011000110",
  51372=>"111101011",
  51373=>"101111101",
  51374=>"100111110",
  51375=>"111101100",
  51376=>"001101010",
  51377=>"100001100",
  51378=>"110110110",
  51379=>"001001001",
  51380=>"111101010",
  51381=>"011101000",
  51382=>"011110111",
  51383=>"011000101",
  51384=>"010011101",
  51385=>"001001011",
  51386=>"011111101",
  51387=>"011100011",
  51388=>"111110101",
  51389=>"001011001",
  51390=>"001001101",
  51391=>"100100001",
  51392=>"011001100",
  51393=>"101111111",
  51394=>"010011111",
  51395=>"101110001",
  51396=>"000110010",
  51397=>"100111000",
  51398=>"100010110",
  51399=>"000000101",
  51400=>"100001000",
  51401=>"101011001",
  51402=>"110100010",
  51403=>"100000001",
  51404=>"000100010",
  51405=>"010000101",
  51406=>"001010110",
  51407=>"000001010",
  51408=>"101011110",
  51409=>"100110100",
  51410=>"111110011",
  51411=>"000101100",
  51412=>"011110110",
  51413=>"001000000",
  51414=>"110010010",
  51415=>"101110110",
  51416=>"001011101",
  51417=>"111100100",
  51418=>"111111011",
  51419=>"101000011",
  51420=>"100011110",
  51421=>"000100010",
  51422=>"011111111",
  51423=>"101101101",
  51424=>"111111100",
  51425=>"011011001",
  51426=>"100101011",
  51427=>"011101001",
  51428=>"111010101",
  51429=>"000011001",
  51430=>"000010101",
  51431=>"101011001",
  51432=>"001100001",
  51433=>"000101000",
  51434=>"000100000",
  51435=>"000100111",
  51436=>"110101011",
  51437=>"001101110",
  51438=>"100110010",
  51439=>"100001101",
  51440=>"001101100",
  51441=>"110110010",
  51442=>"001110011",
  51443=>"111110101",
  51444=>"101101101",
  51445=>"100110110",
  51446=>"111110111",
  51447=>"100001101",
  51448=>"101010001",
  51449=>"110010101",
  51450=>"100101111",
  51451=>"000110001",
  51452=>"111100100",
  51453=>"101100010",
  51454=>"101100110",
  51455=>"101111000",
  51456=>"101001011",
  51457=>"001100110",
  51458=>"110010100",
  51459=>"111111010",
  51460=>"000010100",
  51461=>"010111111",
  51462=>"101001110",
  51463=>"100110111",
  51464=>"000011001",
  51465=>"000001001",
  51466=>"101110111",
  51467=>"110110010",
  51468=>"011101011",
  51469=>"001010100",
  51470=>"011110010",
  51471=>"001011101",
  51472=>"101010011",
  51473=>"011000000",
  51474=>"001011000",
  51475=>"010001010",
  51476=>"010111001",
  51477=>"001010000",
  51478=>"010000101",
  51479=>"100001000",
  51480=>"011111100",
  51481=>"100111101",
  51482=>"000001100",
  51483=>"111110000",
  51484=>"110001001",
  51485=>"000001111",
  51486=>"111111101",
  51487=>"000001000",
  51488=>"111001101",
  51489=>"001111111",
  51490=>"001000011",
  51491=>"011100011",
  51492=>"000100101",
  51493=>"100001000",
  51494=>"111111111",
  51495=>"010101100",
  51496=>"011101001",
  51497=>"000101111",
  51498=>"100111111",
  51499=>"011010110",
  51500=>"111110000",
  51501=>"010100010",
  51502=>"010110010",
  51503=>"001100111",
  51504=>"010111110",
  51505=>"000101011",
  51506=>"001010010",
  51507=>"010011111",
  51508=>"000111111",
  51509=>"011010101",
  51510=>"000101010",
  51511=>"101010100",
  51512=>"001010000",
  51513=>"100000101",
  51514=>"001010101",
  51515=>"100011111",
  51516=>"010001111",
  51517=>"101101101",
  51518=>"100101110",
  51519=>"011010100",
  51520=>"110011011",
  51521=>"001001010",
  51522=>"111010100",
  51523=>"100011101",
  51524=>"110001001",
  51525=>"010111011",
  51526=>"100100010",
  51527=>"010100010",
  51528=>"101000111",
  51529=>"000101101",
  51530=>"001011111",
  51531=>"111001110",
  51532=>"010101001",
  51533=>"110100100",
  51534=>"111110101",
  51535=>"110010110",
  51536=>"110010000",
  51537=>"111011110",
  51538=>"111000100",
  51539=>"110100001",
  51540=>"010110010",
  51541=>"001100010",
  51542=>"101001001",
  51543=>"000010111",
  51544=>"110011110",
  51545=>"011100100",
  51546=>"011000100",
  51547=>"101010000",
  51548=>"111001010",
  51549=>"011111001",
  51550=>"010110100",
  51551=>"000001000",
  51552=>"000011001",
  51553=>"011101100",
  51554=>"111111101",
  51555=>"100010000",
  51556=>"111011010",
  51557=>"000001101",
  51558=>"101001000",
  51559=>"101111101",
  51560=>"111010001",
  51561=>"010111011",
  51562=>"001100100",
  51563=>"000010011",
  51564=>"010110111",
  51565=>"010001010",
  51566=>"000011001",
  51567=>"000011011",
  51568=>"010100010",
  51569=>"011000110",
  51570=>"110011001",
  51571=>"000010010",
  51572=>"001011011",
  51573=>"000101101",
  51574=>"111000001",
  51575=>"101111111",
  51576=>"111000110",
  51577=>"011111111",
  51578=>"000010011",
  51579=>"001101101",
  51580=>"111010111",
  51581=>"101000111",
  51582=>"111110100",
  51583=>"010000110",
  51584=>"000001011",
  51585=>"000011111",
  51586=>"001011011",
  51587=>"000111101",
  51588=>"100000000",
  51589=>"000101010",
  51590=>"010101010",
  51591=>"111101001",
  51592=>"110010111",
  51593=>"001110001",
  51594=>"111010101",
  51595=>"010011101",
  51596=>"010011111",
  51597=>"010100011",
  51598=>"100000000",
  51599=>"010100101",
  51600=>"010001111",
  51601=>"101000110",
  51602=>"110111011",
  51603=>"111011111",
  51604=>"001000100",
  51605=>"101011110",
  51606=>"100011000",
  51607=>"011100100",
  51608=>"011011001",
  51609=>"000011011",
  51610=>"001101001",
  51611=>"000101011",
  51612=>"111110111",
  51613=>"011001010",
  51614=>"110100110",
  51615=>"110111100",
  51616=>"101011010",
  51617=>"111011010",
  51618=>"111001001",
  51619=>"011111101",
  51620=>"000001000",
  51621=>"000011100",
  51622=>"110001110",
  51623=>"100011001",
  51624=>"011110110",
  51625=>"110001000",
  51626=>"001100100",
  51627=>"000110100",
  51628=>"000011101",
  51629=>"011111111",
  51630=>"110001110",
  51631=>"011011001",
  51632=>"011101000",
  51633=>"001111111",
  51634=>"101110111",
  51635=>"001001001",
  51636=>"010010000",
  51637=>"100011110",
  51638=>"100111111",
  51639=>"010011100",
  51640=>"101011101",
  51641=>"010110001",
  51642=>"000110110",
  51643=>"101101001",
  51644=>"011111100",
  51645=>"001100011",
  51646=>"110101001",
  51647=>"010110100",
  51648=>"001000011",
  51649=>"000110001",
  51650=>"001000001",
  51651=>"100110011",
  51652=>"111011110",
  51653=>"110001010",
  51654=>"001111110",
  51655=>"000101001",
  51656=>"001000111",
  51657=>"011011111",
  51658=>"011110110",
  51659=>"101101010",
  51660=>"101000001",
  51661=>"111111001",
  51662=>"001111100",
  51663=>"111101001",
  51664=>"000001100",
  51665=>"111011001",
  51666=>"001010000",
  51667=>"111110000",
  51668=>"011011100",
  51669=>"000001110",
  51670=>"011011011",
  51671=>"001001000",
  51672=>"101000101",
  51673=>"101111010",
  51674=>"010100000",
  51675=>"001000100",
  51676=>"101011010",
  51677=>"001111100",
  51678=>"010011000",
  51679=>"010111000",
  51680=>"101111110",
  51681=>"111110010",
  51682=>"000000010",
  51683=>"000111011",
  51684=>"010001000",
  51685=>"010110101",
  51686=>"011011111",
  51687=>"001100111",
  51688=>"110101011",
  51689=>"011010000",
  51690=>"011100010",
  51691=>"010100001",
  51692=>"110101011",
  51693=>"010100100",
  51694=>"110011110",
  51695=>"011100110",
  51696=>"111101010",
  51697=>"000001001",
  51698=>"010100010",
  51699=>"010100100",
  51700=>"100111111",
  51701=>"100011101",
  51702=>"011000011",
  51703=>"100001110",
  51704=>"100001100",
  51705=>"111101001",
  51706=>"000001110",
  51707=>"111001111",
  51708=>"011100111",
  51709=>"001110001",
  51710=>"011000010",
  51711=>"000000011",
  51712=>"100011000",
  51713=>"000000111",
  51714=>"110010011",
  51715=>"111010111",
  51716=>"011100111",
  51717=>"100101100",
  51718=>"010110111",
  51719=>"111001011",
  51720=>"111011000",
  51721=>"001100101",
  51722=>"111100010",
  51723=>"110101000",
  51724=>"000000000",
  51725=>"011110100",
  51726=>"110001011",
  51727=>"000001110",
  51728=>"000100101",
  51729=>"110011001",
  51730=>"001001010",
  51731=>"100011000",
  51732=>"110110001",
  51733=>"111110011",
  51734=>"000011000",
  51735=>"111001110",
  51736=>"010111001",
  51737=>"110000010",
  51738=>"010011011",
  51739=>"101001011",
  51740=>"000100010",
  51741=>"000100111",
  51742=>"011110111",
  51743=>"011001010",
  51744=>"101011000",
  51745=>"011010001",
  51746=>"000100001",
  51747=>"111001000",
  51748=>"010000011",
  51749=>"001000101",
  51750=>"010111000",
  51751=>"101010001",
  51752=>"001000011",
  51753=>"110111110",
  51754=>"110111011",
  51755=>"101111100",
  51756=>"110101011",
  51757=>"110000100",
  51758=>"001000111",
  51759=>"001100101",
  51760=>"101100101",
  51761=>"011000000",
  51762=>"000001000",
  51763=>"011001111",
  51764=>"110100101",
  51765=>"000100001",
  51766=>"101110010",
  51767=>"110110000",
  51768=>"011100100",
  51769=>"101100011",
  51770=>"001100010",
  51771=>"010101110",
  51772=>"101001101",
  51773=>"100110100",
  51774=>"011011111",
  51775=>"010111111",
  51776=>"010000100",
  51777=>"011110100",
  51778=>"011111011",
  51779=>"111101000",
  51780=>"101101110",
  51781=>"100000100",
  51782=>"101100001",
  51783=>"000110011",
  51784=>"100000101",
  51785=>"011000001",
  51786=>"111010010",
  51787=>"011010010",
  51788=>"110000000",
  51789=>"011101101",
  51790=>"101011111",
  51791=>"100010001",
  51792=>"001101101",
  51793=>"011010011",
  51794=>"010110000",
  51795=>"000110101",
  51796=>"010010001",
  51797=>"011111001",
  51798=>"001110111",
  51799=>"011101000",
  51800=>"011011000",
  51801=>"101100010",
  51802=>"100010011",
  51803=>"000001010",
  51804=>"001000111",
  51805=>"000000100",
  51806=>"101100101",
  51807=>"001101101",
  51808=>"111000010",
  51809=>"100000011",
  51810=>"100000000",
  51811=>"010000111",
  51812=>"000001101",
  51813=>"011001010",
  51814=>"100001100",
  51815=>"001010111",
  51816=>"011001110",
  51817=>"011100101",
  51818=>"010100011",
  51819=>"101001111",
  51820=>"000100111",
  51821=>"110010000",
  51822=>"110110111",
  51823=>"010101010",
  51824=>"000001110",
  51825=>"001100011",
  51826=>"010010010",
  51827=>"010011011",
  51828=>"001111011",
  51829=>"111000101",
  51830=>"000010101",
  51831=>"011010111",
  51832=>"111000110",
  51833=>"011110101",
  51834=>"010011101",
  51835=>"001011111",
  51836=>"011010110",
  51837=>"000011011",
  51838=>"010010111",
  51839=>"011011111",
  51840=>"111110101",
  51841=>"100100101",
  51842=>"001100011",
  51843=>"011101011",
  51844=>"011100001",
  51845=>"000000111",
  51846=>"000001101",
  51847=>"101110111",
  51848=>"001001000",
  51849=>"001000011",
  51850=>"010011101",
  51851=>"100000001",
  51852=>"000011000",
  51853=>"001011010",
  51854=>"100001101",
  51855=>"010101101",
  51856=>"111111111",
  51857=>"001011001",
  51858=>"001000011",
  51859=>"011000001",
  51860=>"011111011",
  51861=>"100100010",
  51862=>"010111100",
  51863=>"110111100",
  51864=>"100000111",
  51865=>"101010010",
  51866=>"001100100",
  51867=>"110001010",
  51868=>"000100010",
  51869=>"101100100",
  51870=>"010000111",
  51871=>"101001001",
  51872=>"100100101",
  51873=>"111001011",
  51874=>"001001111",
  51875=>"001100110",
  51876=>"011101011",
  51877=>"110101000",
  51878=>"000010100",
  51879=>"111111001",
  51880=>"010010000",
  51881=>"010010111",
  51882=>"010101110",
  51883=>"110101100",
  51884=>"001110000",
  51885=>"100000110",
  51886=>"011111101",
  51887=>"100101111",
  51888=>"111001010",
  51889=>"010100011",
  51890=>"100111011",
  51891=>"101001000",
  51892=>"010010000",
  51893=>"111111111",
  51894=>"011111001",
  51895=>"010111110",
  51896=>"101010100",
  51897=>"100000001",
  51898=>"110110101",
  51899=>"001110001",
  51900=>"110010001",
  51901=>"110101110",
  51902=>"000011111",
  51903=>"101100100",
  51904=>"010011001",
  51905=>"101100001",
  51906=>"000100000",
  51907=>"100100001",
  51908=>"101101010",
  51909=>"011001000",
  51910=>"100010111",
  51911=>"100001011",
  51912=>"001011110",
  51913=>"001101101",
  51914=>"011111010",
  51915=>"111110001",
  51916=>"010000010",
  51917=>"011111111",
  51918=>"110100010",
  51919=>"000000010",
  51920=>"100001100",
  51921=>"010101100",
  51922=>"110000001",
  51923=>"000101101",
  51924=>"101001000",
  51925=>"010011011",
  51926=>"100011001",
  51927=>"100011000",
  51928=>"001011011",
  51929=>"010101010",
  51930=>"101010100",
  51931=>"110111000",
  51932=>"001001100",
  51933=>"110100110",
  51934=>"110100000",
  51935=>"100100101",
  51936=>"110101000",
  51937=>"001111110",
  51938=>"010001000",
  51939=>"100110011",
  51940=>"011101111",
  51941=>"000000011",
  51942=>"110000000",
  51943=>"011110000",
  51944=>"101011111",
  51945=>"101000000",
  51946=>"100110001",
  51947=>"111011010",
  51948=>"111001001",
  51949=>"011010101",
  51950=>"010111010",
  51951=>"001010100",
  51952=>"101111100",
  51953=>"101101100",
  51954=>"111010011",
  51955=>"011010001",
  51956=>"100001011",
  51957=>"110101111",
  51958=>"111111000",
  51959=>"111001111",
  51960=>"011110001",
  51961=>"100001101",
  51962=>"011100011",
  51963=>"000010111",
  51964=>"010011111",
  51965=>"010000001",
  51966=>"111010111",
  51967=>"011010001",
  51968=>"110100000",
  51969=>"011000111",
  51970=>"011110010",
  51971=>"101011010",
  51972=>"111000101",
  51973=>"000100001",
  51974=>"010101011",
  51975=>"000011101",
  51976=>"000100001",
  51977=>"010011100",
  51978=>"001101001",
  51979=>"000001000",
  51980=>"100010011",
  51981=>"001110011",
  51982=>"000001101",
  51983=>"010001110",
  51984=>"100111111",
  51985=>"001001011",
  51986=>"001100111",
  51987=>"100101111",
  51988=>"101000111",
  51989=>"000101101",
  51990=>"100110101",
  51991=>"000001000",
  51992=>"001111110",
  51993=>"110111000",
  51994=>"111100000",
  51995=>"001001000",
  51996=>"111100000",
  51997=>"010100001",
  51998=>"111110000",
  51999=>"001110011",
  52000=>"100111110",
  52001=>"110000110",
  52002=>"100110000",
  52003=>"000100100",
  52004=>"011000101",
  52005=>"000101100",
  52006=>"001100011",
  52007=>"000111001",
  52008=>"010100010",
  52009=>"111010111",
  52010=>"010001010",
  52011=>"101100100",
  52012=>"110011111",
  52013=>"110000100",
  52014=>"000100001",
  52015=>"110011010",
  52016=>"000101111",
  52017=>"100011001",
  52018=>"111001110",
  52019=>"001100110",
  52020=>"101000001",
  52021=>"111100111",
  52022=>"000111111",
  52023=>"000111101",
  52024=>"100001000",
  52025=>"110100100",
  52026=>"111001110",
  52027=>"001001010",
  52028=>"111100100",
  52029=>"001110001",
  52030=>"010100001",
  52031=>"111100000",
  52032=>"111100110",
  52033=>"000110110",
  52034=>"100010001",
  52035=>"000000001",
  52036=>"001100001",
  52037=>"010001110",
  52038=>"001100010",
  52039=>"011101100",
  52040=>"100100000",
  52041=>"010010111",
  52042=>"000100001",
  52043=>"011011101",
  52044=>"000100010",
  52045=>"101011100",
  52046=>"110110000",
  52047=>"011101000",
  52048=>"001000100",
  52049=>"100010110",
  52050=>"111000101",
  52051=>"001100100",
  52052=>"000000000",
  52053=>"000111001",
  52054=>"011001101",
  52055=>"100001001",
  52056=>"000000111",
  52057=>"001011110",
  52058=>"011001001",
  52059=>"100111111",
  52060=>"111100101",
  52061=>"111101111",
  52062=>"111011001",
  52063=>"001001101",
  52064=>"011101001",
  52065=>"111001001",
  52066=>"010010110",
  52067=>"010010011",
  52068=>"110011110",
  52069=>"010000001",
  52070=>"100010101",
  52071=>"100110101",
  52072=>"011101011",
  52073=>"000111111",
  52074=>"110101110",
  52075=>"010000010",
  52076=>"111110111",
  52077=>"101110011",
  52078=>"111110000",
  52079=>"000011011",
  52080=>"111001011",
  52081=>"000001010",
  52082=>"101101111",
  52083=>"110011101",
  52084=>"001010010",
  52085=>"000000110",
  52086=>"010100010",
  52087=>"101100100",
  52088=>"110101011",
  52089=>"001101100",
  52090=>"001101101",
  52091=>"011010110",
  52092=>"011010001",
  52093=>"101010111",
  52094=>"011011000",
  52095=>"111000010",
  52096=>"011010010",
  52097=>"111001000",
  52098=>"100110100",
  52099=>"010101101",
  52100=>"100110110",
  52101=>"101011011",
  52102=>"011110110",
  52103=>"101011101",
  52104=>"111111110",
  52105=>"110101101",
  52106=>"010110111",
  52107=>"000011000",
  52108=>"011111100",
  52109=>"000110111",
  52110=>"000100111",
  52111=>"000110101",
  52112=>"011010011",
  52113=>"111010000",
  52114=>"101010000",
  52115=>"101100010",
  52116=>"110111010",
  52117=>"000111001",
  52118=>"111011010",
  52119=>"101010100",
  52120=>"000000111",
  52121=>"110100001",
  52122=>"010110100",
  52123=>"010011000",
  52124=>"111110100",
  52125=>"101110010",
  52126=>"010010110",
  52127=>"000100101",
  52128=>"100001001",
  52129=>"110111011",
  52130=>"000011100",
  52131=>"101011100",
  52132=>"100011111",
  52133=>"011100010",
  52134=>"011111001",
  52135=>"011011111",
  52136=>"110000111",
  52137=>"111010101",
  52138=>"001001010",
  52139=>"101111001",
  52140=>"111111000",
  52141=>"110101110",
  52142=>"110110110",
  52143=>"100100010",
  52144=>"001110110",
  52145=>"101100100",
  52146=>"011110000",
  52147=>"100010100",
  52148=>"000000001",
  52149=>"111100000",
  52150=>"000000010",
  52151=>"000111111",
  52152=>"011101000",
  52153=>"101111010",
  52154=>"001011110",
  52155=>"100110110",
  52156=>"101111111",
  52157=>"001111010",
  52158=>"111010000",
  52159=>"101011011",
  52160=>"001111000",
  52161=>"100011101",
  52162=>"010001100",
  52163=>"110100000",
  52164=>"100110110",
  52165=>"111110101",
  52166=>"001111100",
  52167=>"000111111",
  52168=>"100001111",
  52169=>"001110101",
  52170=>"001000111",
  52171=>"100000100",
  52172=>"100001010",
  52173=>"000011101",
  52174=>"000111111",
  52175=>"110000011",
  52176=>"111001101",
  52177=>"001001101",
  52178=>"010101101",
  52179=>"000000100",
  52180=>"100000110",
  52181=>"001101001",
  52182=>"100101110",
  52183=>"111011100",
  52184=>"111110011",
  52185=>"111001110",
  52186=>"111111010",
  52187=>"000010011",
  52188=>"010101010",
  52189=>"011001010",
  52190=>"100001000",
  52191=>"010111001",
  52192=>"011100101",
  52193=>"111000100",
  52194=>"011111111",
  52195=>"001111011",
  52196=>"100111010",
  52197=>"011110100",
  52198=>"000110101",
  52199=>"000000010",
  52200=>"000011110",
  52201=>"111011010",
  52202=>"000011001",
  52203=>"101010011",
  52204=>"000001100",
  52205=>"100011110",
  52206=>"010011010",
  52207=>"001100011",
  52208=>"101000101",
  52209=>"010100001",
  52210=>"111010011",
  52211=>"110001101",
  52212=>"110110100",
  52213=>"001000111",
  52214=>"011100001",
  52215=>"000000110",
  52216=>"100010111",
  52217=>"010111010",
  52218=>"110111001",
  52219=>"101001011",
  52220=>"000101000",
  52221=>"010010101",
  52222=>"000100011",
  52223=>"010101101",
  52224=>"000001010",
  52225=>"110010010",
  52226=>"110100010",
  52227=>"100001000",
  52228=>"011100000",
  52229=>"010110000",
  52230=>"001110000",
  52231=>"111110100",
  52232=>"011000110",
  52233=>"110001110",
  52234=>"010110110",
  52235=>"101011001",
  52236=>"000110110",
  52237=>"010100001",
  52238=>"011111011",
  52239=>"000110000",
  52240=>"100110100",
  52241=>"000010110",
  52242=>"111001100",
  52243=>"100101010",
  52244=>"011010100",
  52245=>"111001110",
  52246=>"000111010",
  52247=>"111000000",
  52248=>"101100000",
  52249=>"101110100",
  52250=>"101001001",
  52251=>"110000000",
  52252=>"011100011",
  52253=>"110111011",
  52254=>"011101010",
  52255=>"000000100",
  52256=>"000001000",
  52257=>"011110101",
  52258=>"110111011",
  52259=>"011001000",
  52260=>"010110011",
  52261=>"110000010",
  52262=>"110010000",
  52263=>"111101111",
  52264=>"000111001",
  52265=>"000000010",
  52266=>"001111001",
  52267=>"101000101",
  52268=>"000000101",
  52269=>"000000010",
  52270=>"110010011",
  52271=>"101110110",
  52272=>"111001100",
  52273=>"011101010",
  52274=>"100011101",
  52275=>"101100010",
  52276=>"011000110",
  52277=>"110101000",
  52278=>"101010110",
  52279=>"001000011",
  52280=>"110000000",
  52281=>"111111111",
  52282=>"110110111",
  52283=>"010110110",
  52284=>"111010100",
  52285=>"010100111",
  52286=>"000100001",
  52287=>"010010001",
  52288=>"010101011",
  52289=>"011011110",
  52290=>"010000000",
  52291=>"100110111",
  52292=>"100010111",
  52293=>"111000100",
  52294=>"011100000",
  52295=>"101011100",
  52296=>"100100000",
  52297=>"000000010",
  52298=>"101110010",
  52299=>"010001100",
  52300=>"101000111",
  52301=>"101011110",
  52302=>"010011000",
  52303=>"110010001",
  52304=>"011111011",
  52305=>"111010010",
  52306=>"100100001",
  52307=>"010001101",
  52308=>"100000011",
  52309=>"010101111",
  52310=>"000001010",
  52311=>"100000001",
  52312=>"000111011",
  52313=>"111011010",
  52314=>"011010111",
  52315=>"010110100",
  52316=>"001011100",
  52317=>"000101101",
  52318=>"000101110",
  52319=>"010111111",
  52320=>"011101101",
  52321=>"010011010",
  52322=>"111111000",
  52323=>"110100000",
  52324=>"001010010",
  52325=>"010010000",
  52326=>"111011101",
  52327=>"110011000",
  52328=>"010101100",
  52329=>"010011000",
  52330=>"111111000",
  52331=>"101110100",
  52332=>"101001010",
  52333=>"010010000",
  52334=>"111001101",
  52335=>"101011000",
  52336=>"111111011",
  52337=>"010001111",
  52338=>"101101101",
  52339=>"000001011",
  52340=>"000101110",
  52341=>"101010100",
  52342=>"111000010",
  52343=>"010100011",
  52344=>"010100000",
  52345=>"100110000",
  52346=>"000110110",
  52347=>"011111011",
  52348=>"011100101",
  52349=>"011100110",
  52350=>"111000010",
  52351=>"100010001",
  52352=>"011001011",
  52353=>"001111011",
  52354=>"011101110",
  52355=>"100000010",
  52356=>"010001100",
  52357=>"101000000",
  52358=>"011110001",
  52359=>"010110110",
  52360=>"010110111",
  52361=>"000110001",
  52362=>"000111001",
  52363=>"011111111",
  52364=>"111000101",
  52365=>"110100101",
  52366=>"001011101",
  52367=>"000000010",
  52368=>"001001011",
  52369=>"100110000",
  52370=>"001101011",
  52371=>"010101110",
  52372=>"111101111",
  52373=>"001011110",
  52374=>"010001100",
  52375=>"111100001",
  52376=>"011110111",
  52377=>"000110110",
  52378=>"110001110",
  52379=>"000000001",
  52380=>"011100001",
  52381=>"001000001",
  52382=>"000110011",
  52383=>"011001100",
  52384=>"101101011",
  52385=>"100010100",
  52386=>"011101110",
  52387=>"100100001",
  52388=>"011011010",
  52389=>"101101111",
  52390=>"100110010",
  52391=>"100001000",
  52392=>"111010100",
  52393=>"101010110",
  52394=>"011010010",
  52395=>"011011010",
  52396=>"111101111",
  52397=>"001110111",
  52398=>"001101111",
  52399=>"100010110",
  52400=>"100010000",
  52401=>"110100011",
  52402=>"011100001",
  52403=>"001111011",
  52404=>"101100110",
  52405=>"000000101",
  52406=>"000010101",
  52407=>"111001011",
  52408=>"110001001",
  52409=>"010110100",
  52410=>"001010100",
  52411=>"110000100",
  52412=>"011001000",
  52413=>"101101001",
  52414=>"110001000",
  52415=>"101001001",
  52416=>"111010110",
  52417=>"101001000",
  52418=>"010111111",
  52419=>"010111110",
  52420=>"100000001",
  52421=>"001011101",
  52422=>"001101000",
  52423=>"011110100",
  52424=>"011111111",
  52425=>"100000101",
  52426=>"001001001",
  52427=>"000101100",
  52428=>"110000011",
  52429=>"100011110",
  52430=>"000001001",
  52431=>"000010000",
  52432=>"100000101",
  52433=>"001011100",
  52434=>"011010101",
  52435=>"101100010",
  52436=>"011000010",
  52437=>"000110111",
  52438=>"100010011",
  52439=>"011101111",
  52440=>"100100001",
  52441=>"011000000",
  52442=>"111101101",
  52443=>"010001100",
  52444=>"100101101",
  52445=>"110101101",
  52446=>"111001110",
  52447=>"010000101",
  52448=>"010011001",
  52449=>"100111101",
  52450=>"010001110",
  52451=>"000100111",
  52452=>"110110100",
  52453=>"100010100",
  52454=>"110111010",
  52455=>"000001010",
  52456=>"011001000",
  52457=>"110100111",
  52458=>"110111000",
  52459=>"001001011",
  52460=>"000010110",
  52461=>"111101011",
  52462=>"110011010",
  52463=>"111110100",
  52464=>"111010010",
  52465=>"110111011",
  52466=>"110100100",
  52467=>"110110100",
  52468=>"001011000",
  52469=>"000101100",
  52470=>"110110110",
  52471=>"000100110",
  52472=>"011100010",
  52473=>"010010101",
  52474=>"010011010",
  52475=>"101001000",
  52476=>"000001101",
  52477=>"010110001",
  52478=>"000000011",
  52479=>"111111110",
  52480=>"110000001",
  52481=>"111010101",
  52482=>"000111101",
  52483=>"111011010",
  52484=>"100010010",
  52485=>"111011001",
  52486=>"011010110",
  52487=>"001011100",
  52488=>"100001100",
  52489=>"011001100",
  52490=>"010001011",
  52491=>"100001001",
  52492=>"100010010",
  52493=>"111001110",
  52494=>"111000101",
  52495=>"011011011",
  52496=>"111010001",
  52497=>"100110101",
  52498=>"100101100",
  52499=>"110111011",
  52500=>"101101001",
  52501=>"010110110",
  52502=>"100100110",
  52503=>"110111010",
  52504=>"010110011",
  52505=>"110001100",
  52506=>"111011001",
  52507=>"000001101",
  52508=>"111110000",
  52509=>"100000111",
  52510=>"111100110",
  52511=>"101101000",
  52512=>"011001100",
  52513=>"101001011",
  52514=>"111001110",
  52515=>"001101010",
  52516=>"101001111",
  52517=>"001010110",
  52518=>"110010111",
  52519=>"010011011",
  52520=>"111101110",
  52521=>"110011110",
  52522=>"000101011",
  52523=>"011000101",
  52524=>"011100101",
  52525=>"001101101",
  52526=>"110000001",
  52527=>"100110001",
  52528=>"110100011",
  52529=>"111001011",
  52530=>"000010001",
  52531=>"000110010",
  52532=>"110111100",
  52533=>"101011111",
  52534=>"010000000",
  52535=>"000111011",
  52536=>"100000111",
  52537=>"101101011",
  52538=>"111111111",
  52539=>"111111011",
  52540=>"000100011",
  52541=>"111010011",
  52542=>"001100101",
  52543=>"011111100",
  52544=>"010111010",
  52545=>"001000001",
  52546=>"111110110",
  52547=>"101000001",
  52548=>"011001000",
  52549=>"000110101",
  52550=>"000000001",
  52551=>"111111101",
  52552=>"101110101",
  52553=>"100110001",
  52554=>"100011001",
  52555=>"111001011",
  52556=>"010111010",
  52557=>"110100110",
  52558=>"100000000",
  52559=>"111111101",
  52560=>"111101100",
  52561=>"000010100",
  52562=>"000100111",
  52563=>"010101100",
  52564=>"010100111",
  52565=>"000010101",
  52566=>"001100101",
  52567=>"011111101",
  52568=>"110110000",
  52569=>"001001100",
  52570=>"010100001",
  52571=>"111111001",
  52572=>"101110000",
  52573=>"000000111",
  52574=>"001101110",
  52575=>"001011001",
  52576=>"010110101",
  52577=>"010110111",
  52578=>"000011110",
  52579=>"111111100",
  52580=>"001001101",
  52581=>"110001010",
  52582=>"000100110",
  52583=>"011111110",
  52584=>"000000011",
  52585=>"010001111",
  52586=>"101011111",
  52587=>"100111111",
  52588=>"010110000",
  52589=>"101000001",
  52590=>"010100100",
  52591=>"010010010",
  52592=>"110101111",
  52593=>"011001000",
  52594=>"001011001",
  52595=>"110000001",
  52596=>"101101100",
  52597=>"010111111",
  52598=>"001100011",
  52599=>"011000000",
  52600=>"111100000",
  52601=>"010011110",
  52602=>"011001010",
  52603=>"010000001",
  52604=>"000110011",
  52605=>"111100101",
  52606=>"000001110",
  52607=>"110111101",
  52608=>"000000101",
  52609=>"111110100",
  52610=>"100100101",
  52611=>"100011110",
  52612=>"100000010",
  52613=>"010101111",
  52614=>"010001010",
  52615=>"001100101",
  52616=>"010010000",
  52617=>"001101101",
  52618=>"000010010",
  52619=>"111011110",
  52620=>"000000111",
  52621=>"011110000",
  52622=>"011001010",
  52623=>"111110010",
  52624=>"000100100",
  52625=>"100000000",
  52626=>"110001001",
  52627=>"000101000",
  52628=>"011110100",
  52629=>"000110110",
  52630=>"010101100",
  52631=>"100110000",
  52632=>"001111000",
  52633=>"010100010",
  52634=>"110101001",
  52635=>"001010101",
  52636=>"111011001",
  52637=>"010000100",
  52638=>"000101101",
  52639=>"000001101",
  52640=>"100011110",
  52641=>"001011110",
  52642=>"110000000",
  52643=>"100010000",
  52644=>"100001010",
  52645=>"000111011",
  52646=>"111011001",
  52647=>"111111010",
  52648=>"101100101",
  52649=>"111000001",
  52650=>"000110111",
  52651=>"010100001",
  52652=>"111110011",
  52653=>"000000101",
  52654=>"110110101",
  52655=>"011001010",
  52656=>"010100110",
  52657=>"110110101",
  52658=>"001100111",
  52659=>"100000001",
  52660=>"101000001",
  52661=>"011110110",
  52662=>"000100101",
  52663=>"010110111",
  52664=>"110101001",
  52665=>"110001011",
  52666=>"010111100",
  52667=>"001011011",
  52668=>"100110110",
  52669=>"100101110",
  52670=>"111111011",
  52671=>"010011010",
  52672=>"010000000",
  52673=>"010001101",
  52674=>"010011010",
  52675=>"101111110",
  52676=>"100010011",
  52677=>"001110011",
  52678=>"101111100",
  52679=>"000001000",
  52680=>"101000100",
  52681=>"001010101",
  52682=>"000110000",
  52683=>"111000011",
  52684=>"011011010",
  52685=>"010001010",
  52686=>"010010101",
  52687=>"100011010",
  52688=>"100101001",
  52689=>"010100000",
  52690=>"000110100",
  52691=>"000100101",
  52692=>"010111000",
  52693=>"101001101",
  52694=>"001010000",
  52695=>"000001101",
  52696=>"110101000",
  52697=>"110101001",
  52698=>"100110101",
  52699=>"110011110",
  52700=>"001111101",
  52701=>"111000010",
  52702=>"110011111",
  52703=>"001111001",
  52704=>"101001010",
  52705=>"100111100",
  52706=>"110001110",
  52707=>"000111001",
  52708=>"010010010",
  52709=>"101001100",
  52710=>"101001111",
  52711=>"010110000",
  52712=>"101001100",
  52713=>"100100101",
  52714=>"011001110",
  52715=>"001011110",
  52716=>"111110000",
  52717=>"111000110",
  52718=>"110101011",
  52719=>"000000001",
  52720=>"000011110",
  52721=>"010111001",
  52722=>"110111001",
  52723=>"001010001",
  52724=>"011001010",
  52725=>"010000001",
  52726=>"110001000",
  52727=>"010000100",
  52728=>"100000001",
  52729=>"110101110",
  52730=>"001101001",
  52731=>"000110111",
  52732=>"000100011",
  52733=>"011001010",
  52734=>"100100000",
  52735=>"000000100",
  52736=>"010011111",
  52737=>"101010001",
  52738=>"110001000",
  52739=>"101010111",
  52740=>"001001001",
  52741=>"010011000",
  52742=>"011001111",
  52743=>"010001011",
  52744=>"010000000",
  52745=>"010011101",
  52746=>"100000010",
  52747=>"111110011",
  52748=>"100111001",
  52749=>"101101100",
  52750=>"111010110",
  52751=>"000011011",
  52752=>"111111101",
  52753=>"010110011",
  52754=>"100010110",
  52755=>"101001110",
  52756=>"100100110",
  52757=>"100101011",
  52758=>"111101111",
  52759=>"001001100",
  52760=>"100001111",
  52761=>"010100010",
  52762=>"001000100",
  52763=>"101011011",
  52764=>"000110001",
  52765=>"000101000",
  52766=>"101010111",
  52767=>"101100001",
  52768=>"010010010",
  52769=>"011110111",
  52770=>"111000000",
  52771=>"001100000",
  52772=>"101011000",
  52773=>"010110111",
  52774=>"110001100",
  52775=>"100011100",
  52776=>"000100101",
  52777=>"011111011",
  52778=>"100000100",
  52779=>"100101001",
  52780=>"101000011",
  52781=>"100101101",
  52782=>"011000101",
  52783=>"001110101",
  52784=>"001101011",
  52785=>"100101110",
  52786=>"101011011",
  52787=>"010010101",
  52788=>"010011001",
  52789=>"001010000",
  52790=>"001110011",
  52791=>"100010011",
  52792=>"100101110",
  52793=>"111101101",
  52794=>"000111010",
  52795=>"000010011",
  52796=>"001001001",
  52797=>"001001100",
  52798=>"100011010",
  52799=>"000101111",
  52800=>"010110100",
  52801=>"000001101",
  52802=>"010010111",
  52803=>"000010011",
  52804=>"000000101",
  52805=>"011011100",
  52806=>"000100001",
  52807=>"000000110",
  52808=>"000010010",
  52809=>"110011111",
  52810=>"001110110",
  52811=>"110110101",
  52812=>"101110000",
  52813=>"100100101",
  52814=>"111001000",
  52815=>"011101101",
  52816=>"111010000",
  52817=>"101100011",
  52818=>"010110011",
  52819=>"100000101",
  52820=>"101011101",
  52821=>"010010000",
  52822=>"001000000",
  52823=>"100101001",
  52824=>"100110011",
  52825=>"100111111",
  52826=>"100110000",
  52827=>"110101100",
  52828=>"100100000",
  52829=>"100110110",
  52830=>"000001111",
  52831=>"110100101",
  52832=>"001101111",
  52833=>"010011001",
  52834=>"111100101",
  52835=>"001000100",
  52836=>"101010010",
  52837=>"000010011",
  52838=>"000011110",
  52839=>"110110101",
  52840=>"011101001",
  52841=>"100001000",
  52842=>"011000101",
  52843=>"101111101",
  52844=>"011010111",
  52845=>"001010000",
  52846=>"111011011",
  52847=>"011101100",
  52848=>"010100110",
  52849=>"100010100",
  52850=>"110011001",
  52851=>"000000000",
  52852=>"110010111",
  52853=>"000001010",
  52854=>"101101000",
  52855=>"010000001",
  52856=>"010001110",
  52857=>"011111011",
  52858=>"010001001",
  52859=>"110001001",
  52860=>"101101110",
  52861=>"000000010",
  52862=>"001010011",
  52863=>"001011110",
  52864=>"010100110",
  52865=>"110011011",
  52866=>"000101110",
  52867=>"111010010",
  52868=>"100011011",
  52869=>"110100101",
  52870=>"110111111",
  52871=>"010111111",
  52872=>"011100001",
  52873=>"010010100",
  52874=>"000100000",
  52875=>"000011110",
  52876=>"111001111",
  52877=>"001000100",
  52878=>"011110101",
  52879=>"000000110",
  52880=>"110011010",
  52881=>"000110100",
  52882=>"110001110",
  52883=>"001101100",
  52884=>"110110000",
  52885=>"010000111",
  52886=>"000001111",
  52887=>"010001001",
  52888=>"111110000",
  52889=>"111011010",
  52890=>"000111000",
  52891=>"001110000",
  52892=>"100011110",
  52893=>"100101101",
  52894=>"111011111",
  52895=>"101010000",
  52896=>"010011000",
  52897=>"000000100",
  52898=>"111010010",
  52899=>"100010011",
  52900=>"000000100",
  52901=>"001010100",
  52902=>"100100101",
  52903=>"111011011",
  52904=>"110010100",
  52905=>"010000000",
  52906=>"010011000",
  52907=>"110111110",
  52908=>"000001000",
  52909=>"110000111",
  52910=>"110011000",
  52911=>"000011011",
  52912=>"000000111",
  52913=>"000000010",
  52914=>"001001011",
  52915=>"110101011",
  52916=>"000101101",
  52917=>"010010100",
  52918=>"111111101",
  52919=>"000011101",
  52920=>"010000001",
  52921=>"101100101",
  52922=>"001110101",
  52923=>"010010111",
  52924=>"100100001",
  52925=>"110010010",
  52926=>"000111001",
  52927=>"111110100",
  52928=>"110010001",
  52929=>"100011011",
  52930=>"101001110",
  52931=>"101000001",
  52932=>"100111010",
  52933=>"100000011",
  52934=>"110010110",
  52935=>"001011001",
  52936=>"101001010",
  52937=>"110011110",
  52938=>"111011101",
  52939=>"101100000",
  52940=>"010001111",
  52941=>"001011111",
  52942=>"110011010",
  52943=>"010100110",
  52944=>"101101000",
  52945=>"001111001",
  52946=>"000001001",
  52947=>"010011101",
  52948=>"100010000",
  52949=>"100010001",
  52950=>"001001111",
  52951=>"000001110",
  52952=>"011000110",
  52953=>"001011110",
  52954=>"111110000",
  52955=>"011101010",
  52956=>"000101100",
  52957=>"111001100",
  52958=>"011010011",
  52959=>"000101111",
  52960=>"010011111",
  52961=>"010011101",
  52962=>"010110101",
  52963=>"010100000",
  52964=>"101110110",
  52965=>"010111011",
  52966=>"011001100",
  52967=>"000001111",
  52968=>"000000100",
  52969=>"001001111",
  52970=>"100100000",
  52971=>"010110000",
  52972=>"111001000",
  52973=>"100110111",
  52974=>"100101000",
  52975=>"000110110",
  52976=>"101011010",
  52977=>"110110110",
  52978=>"101100000",
  52979=>"011111011",
  52980=>"000001011",
  52981=>"011101100",
  52982=>"010000011",
  52983=>"110101001",
  52984=>"111111011",
  52985=>"010011110",
  52986=>"111010011",
  52987=>"110100000",
  52988=>"111111101",
  52989=>"110100010",
  52990=>"111111100",
  52991=>"011100010",
  52992=>"000101000",
  52993=>"100011011",
  52994=>"101100001",
  52995=>"000101001",
  52996=>"010001001",
  52997=>"000000011",
  52998=>"001011110",
  52999=>"011010101",
  53000=>"011100000",
  53001=>"100111110",
  53002=>"000101011",
  53003=>"000110110",
  53004=>"000011110",
  53005=>"000011010",
  53006=>"101011110",
  53007=>"111110110",
  53008=>"001110010",
  53009=>"110110100",
  53010=>"001010011",
  53011=>"001100011",
  53012=>"111110100",
  53013=>"001101110",
  53014=>"110000010",
  53015=>"110000001",
  53016=>"000111011",
  53017=>"011100011",
  53018=>"010101010",
  53019=>"001011011",
  53020=>"001010001",
  53021=>"111111001",
  53022=>"011111000",
  53023=>"000100101",
  53024=>"010000101",
  53025=>"000010101",
  53026=>"110010001",
  53027=>"110001100",
  53028=>"100100010",
  53029=>"001010011",
  53030=>"110001010",
  53031=>"011101110",
  53032=>"001001101",
  53033=>"101001011",
  53034=>"000101010",
  53035=>"110110010",
  53036=>"001110101",
  53037=>"010000110",
  53038=>"100001011",
  53039=>"001101011",
  53040=>"000101010",
  53041=>"011011011",
  53042=>"001011101",
  53043=>"011001000",
  53044=>"000000011",
  53045=>"001001000",
  53046=>"001011111",
  53047=>"001010010",
  53048=>"110101000",
  53049=>"000111111",
  53050=>"111001001",
  53051=>"011111101",
  53052=>"010000001",
  53053=>"000100000",
  53054=>"111001010",
  53055=>"110100111",
  53056=>"001101010",
  53057=>"100011100",
  53058=>"101101110",
  53059=>"010100111",
  53060=>"000010110",
  53061=>"110100100",
  53062=>"101100001",
  53063=>"000001111",
  53064=>"011011110",
  53065=>"111001000",
  53066=>"000111001",
  53067=>"011111100",
  53068=>"001110010",
  53069=>"011011001",
  53070=>"101101001",
  53071=>"000000000",
  53072=>"111111011",
  53073=>"011110100",
  53074=>"010011000",
  53075=>"000101010",
  53076=>"100001001",
  53077=>"001011001",
  53078=>"110001101",
  53079=>"001001010",
  53080=>"010111100",
  53081=>"101001100",
  53082=>"010001111",
  53083=>"111110001",
  53084=>"101010010",
  53085=>"101111010",
  53086=>"000000101",
  53087=>"100000101",
  53088=>"101000011",
  53089=>"110000110",
  53090=>"000101010",
  53091=>"100001011",
  53092=>"010010111",
  53093=>"010111010",
  53094=>"000010111",
  53095=>"001110110",
  53096=>"011110000",
  53097=>"100100111",
  53098=>"001001110",
  53099=>"110011001",
  53100=>"111000001",
  53101=>"101011110",
  53102=>"111011110",
  53103=>"011100000",
  53104=>"111101011",
  53105=>"010011110",
  53106=>"100101100",
  53107=>"101000101",
  53108=>"100001000",
  53109=>"110010111",
  53110=>"000011110",
  53111=>"010001010",
  53112=>"011100110",
  53113=>"100000111",
  53114=>"101011010",
  53115=>"011010001",
  53116=>"000100110",
  53117=>"110101100",
  53118=>"011011001",
  53119=>"100011110",
  53120=>"001101101",
  53121=>"000101111",
  53122=>"011000011",
  53123=>"111011000",
  53124=>"101011110",
  53125=>"101001000",
  53126=>"010111011",
  53127=>"000110011",
  53128=>"011001010",
  53129=>"011111111",
  53130=>"101001010",
  53131=>"000001001",
  53132=>"011111001",
  53133=>"011101010",
  53134=>"101111010",
  53135=>"111110011",
  53136=>"110101111",
  53137=>"100100100",
  53138=>"001000010",
  53139=>"000010001",
  53140=>"000101001",
  53141=>"111100010",
  53142=>"010100000",
  53143=>"111011001",
  53144=>"111100111",
  53145=>"100110100",
  53146=>"010011001",
  53147=>"000111011",
  53148=>"100010010",
  53149=>"001111100",
  53150=>"100001011",
  53151=>"101110011",
  53152=>"001000100",
  53153=>"000110011",
  53154=>"101001000",
  53155=>"010000101",
  53156=>"000010111",
  53157=>"011001101",
  53158=>"111110101",
  53159=>"101100111",
  53160=>"100110111",
  53161=>"010011011",
  53162=>"001101100",
  53163=>"000010110",
  53164=>"101010001",
  53165=>"001000111",
  53166=>"110010010",
  53167=>"001101001",
  53168=>"101101100",
  53169=>"001110100",
  53170=>"101110100",
  53171=>"111011010",
  53172=>"011111001",
  53173=>"101101000",
  53174=>"110111111",
  53175=>"010011100",
  53176=>"111001000",
  53177=>"110001100",
  53178=>"111001111",
  53179=>"111000110",
  53180=>"111110001",
  53181=>"110000110",
  53182=>"111001111",
  53183=>"100000001",
  53184=>"100001100",
  53185=>"101011010",
  53186=>"111110011",
  53187=>"001010000",
  53188=>"001101001",
  53189=>"000010110",
  53190=>"110100010",
  53191=>"010101010",
  53192=>"001100001",
  53193=>"001100111",
  53194=>"111101010",
  53195=>"111110011",
  53196=>"011010100",
  53197=>"001101101",
  53198=>"011101011",
  53199=>"010100101",
  53200=>"100101111",
  53201=>"101000010",
  53202=>"000110000",
  53203=>"001111010",
  53204=>"011100111",
  53205=>"111101010",
  53206=>"011011110",
  53207=>"100101100",
  53208=>"111001101",
  53209=>"101101011",
  53210=>"111111101",
  53211=>"010110101",
  53212=>"011000001",
  53213=>"010101011",
  53214=>"000010101",
  53215=>"001111100",
  53216=>"100101111",
  53217=>"100101011",
  53218=>"000000001",
  53219=>"010000110",
  53220=>"100000010",
  53221=>"100001010",
  53222=>"010001100",
  53223=>"100010101",
  53224=>"000000111",
  53225=>"111111011",
  53226=>"000000000",
  53227=>"100110011",
  53228=>"110010010",
  53229=>"111010000",
  53230=>"110100000",
  53231=>"001010000",
  53232=>"000101111",
  53233=>"100011110",
  53234=>"110100110",
  53235=>"000000101",
  53236=>"010010100",
  53237=>"001101000",
  53238=>"101100110",
  53239=>"001110000",
  53240=>"110101101",
  53241=>"011100111",
  53242=>"110001101",
  53243=>"001011100",
  53244=>"110001010",
  53245=>"001101001",
  53246=>"101000011",
  53247=>"011000101",
  53248=>"101000000",
  53249=>"000011001",
  53250=>"011110101",
  53251=>"010001100",
  53252=>"111110001",
  53253=>"101110100",
  53254=>"100110101",
  53255=>"111010111",
  53256=>"001101100",
  53257=>"111010001",
  53258=>"101111010",
  53259=>"010110010",
  53260=>"000111001",
  53261=>"111101111",
  53262=>"001000100",
  53263=>"101011101",
  53264=>"111000001",
  53265=>"100010001",
  53266=>"000001010",
  53267=>"000010000",
  53268=>"111101011",
  53269=>"010001011",
  53270=>"110100000",
  53271=>"111101100",
  53272=>"001111111",
  53273=>"000000100",
  53274=>"001110000",
  53275=>"011010000",
  53276=>"111100111",
  53277=>"011111010",
  53278=>"110001100",
  53279=>"010000010",
  53280=>"011010100",
  53281=>"111101101",
  53282=>"100101010",
  53283=>"110100001",
  53284=>"000010000",
  53285=>"001011011",
  53286=>"111010110",
  53287=>"010000000",
  53288=>"111101000",
  53289=>"110110011",
  53290=>"100111010",
  53291=>"100010010",
  53292=>"001000000",
  53293=>"110010011",
  53294=>"001101101",
  53295=>"010011011",
  53296=>"111000001",
  53297=>"001011101",
  53298=>"000111001",
  53299=>"110110011",
  53300=>"011011110",
  53301=>"000001100",
  53302=>"000101111",
  53303=>"100000100",
  53304=>"000110100",
  53305=>"101010111",
  53306=>"111111111",
  53307=>"000100110",
  53308=>"110011011",
  53309=>"100011101",
  53310=>"111100101",
  53311=>"011001000",
  53312=>"000111110",
  53313=>"101100011",
  53314=>"000010000",
  53315=>"010100010",
  53316=>"110011001",
  53317=>"011101011",
  53318=>"111000010",
  53319=>"000101101",
  53320=>"111110000",
  53321=>"000000001",
  53322=>"011011001",
  53323=>"000010011",
  53324=>"010111011",
  53325=>"110011100",
  53326=>"001101100",
  53327=>"011010000",
  53328=>"010001011",
  53329=>"011110011",
  53330=>"101000100",
  53331=>"111100000",
  53332=>"001100101",
  53333=>"000001010",
  53334=>"011111011",
  53335=>"001000001",
  53336=>"000011111",
  53337=>"011101100",
  53338=>"000000001",
  53339=>"110010101",
  53340=>"011101110",
  53341=>"010111111",
  53342=>"010101101",
  53343=>"111101101",
  53344=>"011001111",
  53345=>"111111101",
  53346=>"100100111",
  53347=>"000000110",
  53348=>"010110110",
  53349=>"010111011",
  53350=>"100111011",
  53351=>"010111001",
  53352=>"010111111",
  53353=>"110001001",
  53354=>"111110111",
  53355=>"111100110",
  53356=>"111001110",
  53357=>"011000000",
  53358=>"011001001",
  53359=>"000110111",
  53360=>"001010001",
  53361=>"001111110",
  53362=>"010011100",
  53363=>"011100010",
  53364=>"100110100",
  53365=>"111011100",
  53366=>"011001011",
  53367=>"101111100",
  53368=>"000001111",
  53369=>"001001011",
  53370=>"011001110",
  53371=>"011110100",
  53372=>"100111100",
  53373=>"000001010",
  53374=>"101010000",
  53375=>"000101001",
  53376=>"011100110",
  53377=>"101100111",
  53378=>"010101000",
  53379=>"000111000",
  53380=>"000110111",
  53381=>"110110100",
  53382=>"100101100",
  53383=>"111100000",
  53384=>"111011011",
  53385=>"011110101",
  53386=>"000111001",
  53387=>"000100111",
  53388=>"111001000",
  53389=>"001011111",
  53390=>"010001100",
  53391=>"011011011",
  53392=>"110001111",
  53393=>"111011010",
  53394=>"010100001",
  53395=>"001101001",
  53396=>"101000011",
  53397=>"101110000",
  53398=>"111111001",
  53399=>"100000000",
  53400=>"001010001",
  53401=>"101110001",
  53402=>"110000111",
  53403=>"100111100",
  53404=>"000110110",
  53405=>"100101110",
  53406=>"000100000",
  53407=>"011101111",
  53408=>"010011100",
  53409=>"010100101",
  53410=>"001101111",
  53411=>"011010001",
  53412=>"000011000",
  53413=>"100010000",
  53414=>"001110110",
  53415=>"000101111",
  53416=>"100011001",
  53417=>"111010101",
  53418=>"101000000",
  53419=>"100100100",
  53420=>"101100100",
  53421=>"001101100",
  53422=>"101001011",
  53423=>"111000000",
  53424=>"000000001",
  53425=>"011100000",
  53426=>"100001010",
  53427=>"010100001",
  53428=>"011110111",
  53429=>"101000011",
  53430=>"011001100",
  53431=>"011010110",
  53432=>"001100100",
  53433=>"010000101",
  53434=>"001010010",
  53435=>"010001100",
  53436=>"011001101",
  53437=>"111111111",
  53438=>"110000000",
  53439=>"001001011",
  53440=>"100100000",
  53441=>"110100110",
  53442=>"001100111",
  53443=>"000010010",
  53444=>"001100011",
  53445=>"010011010",
  53446=>"100010000",
  53447=>"001001001",
  53448=>"101100011",
  53449=>"100111101",
  53450=>"010010101",
  53451=>"111110010",
  53452=>"100010110",
  53453=>"110010010",
  53454=>"011000001",
  53455=>"111001001",
  53456=>"000011101",
  53457=>"000011000",
  53458=>"111100100",
  53459=>"101001101",
  53460=>"111000111",
  53461=>"011110001",
  53462=>"101011101",
  53463=>"111100110",
  53464=>"000001001",
  53465=>"101000001",
  53466=>"001101000",
  53467=>"111101110",
  53468=>"100011100",
  53469=>"000101100",
  53470=>"000001110",
  53471=>"111011111",
  53472=>"010010111",
  53473=>"100110001",
  53474=>"100111111",
  53475=>"001000001",
  53476=>"100011010",
  53477=>"110110110",
  53478=>"100110000",
  53479=>"100000000",
  53480=>"011111100",
  53481=>"001100111",
  53482=>"000100111",
  53483=>"000000011",
  53484=>"010000010",
  53485=>"011000110",
  53486=>"111110100",
  53487=>"000001011",
  53488=>"101111111",
  53489=>"100000011",
  53490=>"000010001",
  53491=>"011001110",
  53492=>"010001111",
  53493=>"011101101",
  53494=>"011000000",
  53495=>"110001000",
  53496=>"101100100",
  53497=>"101111011",
  53498=>"000110011",
  53499=>"100101000",
  53500=>"110011100",
  53501=>"000110111",
  53502=>"001010001",
  53503=>"011011010",
  53504=>"110001000",
  53505=>"011000000",
  53506=>"111010100",
  53507=>"111001000",
  53508=>"010100000",
  53509=>"111101111",
  53510=>"000010011",
  53511=>"100000100",
  53512=>"100001001",
  53513=>"010010011",
  53514=>"011010010",
  53515=>"000001101",
  53516=>"101111100",
  53517=>"000011101",
  53518=>"111000111",
  53519=>"000000011",
  53520=>"111111110",
  53521=>"110011010",
  53522=>"001000100",
  53523=>"000111111",
  53524=>"100000011",
  53525=>"010000000",
  53526=>"100111001",
  53527=>"110001110",
  53528=>"001101011",
  53529=>"000110001",
  53530=>"101001111",
  53531=>"110111001",
  53532=>"010001010",
  53533=>"110111110",
  53534=>"010101011",
  53535=>"110010010",
  53536=>"100101000",
  53537=>"101100101",
  53538=>"110011101",
  53539=>"001101101",
  53540=>"100010101",
  53541=>"100010101",
  53542=>"111000101",
  53543=>"101100000",
  53544=>"001001101",
  53545=>"000001000",
  53546=>"111000110",
  53547=>"110101011",
  53548=>"000010000",
  53549=>"001110011",
  53550=>"110010110",
  53551=>"001100011",
  53552=>"011110100",
  53553=>"110001111",
  53554=>"010100101",
  53555=>"110111101",
  53556=>"101001010",
  53557=>"000111100",
  53558=>"100010110",
  53559=>"101001000",
  53560=>"101101000",
  53561=>"111111001",
  53562=>"100110010",
  53563=>"010001000",
  53564=>"100100101",
  53565=>"001010101",
  53566=>"100010101",
  53567=>"000010111",
  53568=>"100111100",
  53569=>"010011111",
  53570=>"101001001",
  53571=>"101101110",
  53572=>"000000101",
  53573=>"011011011",
  53574=>"001110011",
  53575=>"000001100",
  53576=>"101111100",
  53577=>"000000011",
  53578=>"001101010",
  53579=>"001001111",
  53580=>"011111101",
  53581=>"101100000",
  53582=>"101110110",
  53583=>"010101111",
  53584=>"001011010",
  53585=>"000100100",
  53586=>"101000000",
  53587=>"010110110",
  53588=>"111100011",
  53589=>"100000100",
  53590=>"000100111",
  53591=>"000010111",
  53592=>"100000001",
  53593=>"001110001",
  53594=>"100100000",
  53595=>"110010100",
  53596=>"101011110",
  53597=>"111111110",
  53598=>"100100101",
  53599=>"001100000",
  53600=>"001000100",
  53601=>"110111000",
  53602=>"000011000",
  53603=>"111100100",
  53604=>"101110001",
  53605=>"010101100",
  53606=>"110100111",
  53607=>"110100100",
  53608=>"101111000",
  53609=>"111000101",
  53610=>"010110111",
  53611=>"111111010",
  53612=>"110110011",
  53613=>"101011101",
  53614=>"000100100",
  53615=>"011011101",
  53616=>"110000001",
  53617=>"010100110",
  53618=>"110110010",
  53619=>"011011101",
  53620=>"111110100",
  53621=>"000011010",
  53622=>"111100001",
  53623=>"111110001",
  53624=>"010110000",
  53625=>"000101001",
  53626=>"011011111",
  53627=>"001011111",
  53628=>"011010110",
  53629=>"001110111",
  53630=>"101111000",
  53631=>"010001111",
  53632=>"100101000",
  53633=>"100011110",
  53634=>"101110010",
  53635=>"001000100",
  53636=>"011101100",
  53637=>"001111011",
  53638=>"110010011",
  53639=>"011001011",
  53640=>"111100011",
  53641=>"101110010",
  53642=>"010101001",
  53643=>"110000101",
  53644=>"010010110",
  53645=>"100010000",
  53646=>"100110110",
  53647=>"010101111",
  53648=>"001001000",
  53649=>"010101010",
  53650=>"011101110",
  53651=>"101000110",
  53652=>"111100011",
  53653=>"111101111",
  53654=>"000000001",
  53655=>"010110010",
  53656=>"110001110",
  53657=>"101011010",
  53658=>"111000011",
  53659=>"000010101",
  53660=>"100100101",
  53661=>"100000000",
  53662=>"000010101",
  53663=>"010110011",
  53664=>"001111101",
  53665=>"111010011",
  53666=>"011111010",
  53667=>"011111111",
  53668=>"000101011",
  53669=>"000000011",
  53670=>"000100000",
  53671=>"011010000",
  53672=>"010101100",
  53673=>"000101010",
  53674=>"101101111",
  53675=>"111010000",
  53676=>"001001100",
  53677=>"010000101",
  53678=>"100010101",
  53679=>"000111111",
  53680=>"100101111",
  53681=>"011111011",
  53682=>"001010011",
  53683=>"000011011",
  53684=>"011001001",
  53685=>"001100011",
  53686=>"011000101",
  53687=>"011010010",
  53688=>"101101001",
  53689=>"000000000",
  53690=>"000000111",
  53691=>"001111110",
  53692=>"010000111",
  53693=>"011111111",
  53694=>"111011101",
  53695=>"100011100",
  53696=>"100010110",
  53697=>"011000011",
  53698=>"010110111",
  53699=>"110100111",
  53700=>"100111111",
  53701=>"100100101",
  53702=>"001110111",
  53703=>"001100111",
  53704=>"010010110",
  53705=>"111011110",
  53706=>"010111111",
  53707=>"111011000",
  53708=>"010111110",
  53709=>"010111100",
  53710=>"110010011",
  53711=>"010110111",
  53712=>"101000010",
  53713=>"111000011",
  53714=>"000001111",
  53715=>"010010110",
  53716=>"010111110",
  53717=>"001010000",
  53718=>"010000011",
  53719=>"111100100",
  53720=>"100011001",
  53721=>"001000011",
  53722=>"111000100",
  53723=>"010110010",
  53724=>"110101010",
  53725=>"010000001",
  53726=>"101011011",
  53727=>"100010101",
  53728=>"110110000",
  53729=>"111101111",
  53730=>"011101101",
  53731=>"110111111",
  53732=>"111110000",
  53733=>"001011010",
  53734=>"100100111",
  53735=>"000000011",
  53736=>"001110110",
  53737=>"000110000",
  53738=>"100100001",
  53739=>"001111001",
  53740=>"101011011",
  53741=>"110010101",
  53742=>"101100011",
  53743=>"110101100",
  53744=>"111111000",
  53745=>"000000010",
  53746=>"010011001",
  53747=>"100011111",
  53748=>"111100111",
  53749=>"100000000",
  53750=>"011101010",
  53751=>"111010000",
  53752=>"000101001",
  53753=>"110111010",
  53754=>"011010000",
  53755=>"101000000",
  53756=>"000100101",
  53757=>"111111100",
  53758=>"000010001",
  53759=>"011111111",
  53760=>"111100001",
  53761=>"111010000",
  53762=>"100001000",
  53763=>"110111010",
  53764=>"010011011",
  53765=>"111100111",
  53766=>"111101010",
  53767=>"111001011",
  53768=>"000110101",
  53769=>"110001101",
  53770=>"101001101",
  53771=>"100011000",
  53772=>"010101010",
  53773=>"110100000",
  53774=>"001110111",
  53775=>"000000111",
  53776=>"100111100",
  53777=>"111010110",
  53778=>"010010001",
  53779=>"001101011",
  53780=>"010000100",
  53781=>"001100100",
  53782=>"000110110",
  53783=>"000001011",
  53784=>"000010000",
  53785=>"011110010",
  53786=>"000001101",
  53787=>"000001010",
  53788=>"110001101",
  53789=>"011010100",
  53790=>"011101000",
  53791=>"111001010",
  53792=>"101000010",
  53793=>"111011111",
  53794=>"011111100",
  53795=>"111111000",
  53796=>"111001101",
  53797=>"000110010",
  53798=>"110101001",
  53799=>"111100010",
  53800=>"000101001",
  53801=>"100101001",
  53802=>"011110111",
  53803=>"100000101",
  53804=>"000001100",
  53805=>"000111111",
  53806=>"010000111",
  53807=>"110010000",
  53808=>"011010001",
  53809=>"001101000",
  53810=>"111111101",
  53811=>"001000110",
  53812=>"101001000",
  53813=>"010010010",
  53814=>"100010011",
  53815=>"110110111",
  53816=>"011011100",
  53817=>"011001110",
  53818=>"111111111",
  53819=>"011100010",
  53820=>"010010000",
  53821=>"110111111",
  53822=>"000101110",
  53823=>"100011111",
  53824=>"111000010",
  53825=>"011110110",
  53826=>"100111110",
  53827=>"110001001",
  53828=>"110011101",
  53829=>"111001111",
  53830=>"001000001",
  53831=>"101000101",
  53832=>"010010011",
  53833=>"100101011",
  53834=>"101000001",
  53835=>"001011101",
  53836=>"101001110",
  53837=>"000011001",
  53838=>"000110101",
  53839=>"010100011",
  53840=>"001001111",
  53841=>"011101011",
  53842=>"011010100",
  53843=>"110010101",
  53844=>"011110010",
  53845=>"010101010",
  53846=>"110001111",
  53847=>"001000100",
  53848=>"110011010",
  53849=>"011111101",
  53850=>"011111010",
  53851=>"111001001",
  53852=>"010011001",
  53853=>"110101001",
  53854=>"111001011",
  53855=>"010000001",
  53856=>"100100100",
  53857=>"101100111",
  53858=>"110101000",
  53859=>"000001000",
  53860=>"100010111",
  53861=>"100010010",
  53862=>"011110111",
  53863=>"101110111",
  53864=>"010111111",
  53865=>"100001000",
  53866=>"110000000",
  53867=>"000111100",
  53868=>"001100101",
  53869=>"011111001",
  53870=>"101100000",
  53871=>"111111001",
  53872=>"110001011",
  53873=>"001110010",
  53874=>"001110011",
  53875=>"000001011",
  53876=>"001000111",
  53877=>"001111011",
  53878=>"100001101",
  53879=>"111001000",
  53880=>"011000010",
  53881=>"001110000",
  53882=>"110101001",
  53883=>"010011011",
  53884=>"101101110",
  53885=>"011010000",
  53886=>"000101110",
  53887=>"110010110",
  53888=>"000100011",
  53889=>"100001011",
  53890=>"111000111",
  53891=>"100011010",
  53892=>"000011001",
  53893=>"010100011",
  53894=>"100100000",
  53895=>"001011011",
  53896=>"000101010",
  53897=>"110010111",
  53898=>"111101100",
  53899=>"100101110",
  53900=>"000111101",
  53901=>"001001001",
  53902=>"111010000",
  53903=>"000110101",
  53904=>"100110011",
  53905=>"111001110",
  53906=>"010000001",
  53907=>"110110100",
  53908=>"011101000",
  53909=>"001001111",
  53910=>"101101000",
  53911=>"101100100",
  53912=>"010111010",
  53913=>"101100001",
  53914=>"000100001",
  53915=>"011000011",
  53916=>"101000010",
  53917=>"001010000",
  53918=>"000110000",
  53919=>"110111111",
  53920=>"110101100",
  53921=>"100011111",
  53922=>"100101110",
  53923=>"001001101",
  53924=>"001000100",
  53925=>"100001011",
  53926=>"011101110",
  53927=>"011111101",
  53928=>"000000110",
  53929=>"101101011",
  53930=>"001000000",
  53931=>"101101000",
  53932=>"000000000",
  53933=>"111101000",
  53934=>"110000001",
  53935=>"100001010",
  53936=>"011110001",
  53937=>"000111111",
  53938=>"011110011",
  53939=>"110000111",
  53940=>"000111100",
  53941=>"010000011",
  53942=>"011111011",
  53943=>"000011000",
  53944=>"010000100",
  53945=>"000010011",
  53946=>"111110001",
  53947=>"001000010",
  53948=>"100111000",
  53949=>"010111111",
  53950=>"111011101",
  53951=>"011110000",
  53952=>"001000101",
  53953=>"010000000",
  53954=>"100100000",
  53955=>"101100011",
  53956=>"110101000",
  53957=>"001100110",
  53958=>"101111110",
  53959=>"100001101",
  53960=>"110101110",
  53961=>"111011001",
  53962=>"100001011",
  53963=>"100101001",
  53964=>"111111010",
  53965=>"010111010",
  53966=>"110111010",
  53967=>"100111100",
  53968=>"111000000",
  53969=>"001101110",
  53970=>"110111010",
  53971=>"100000101",
  53972=>"100100110",
  53973=>"110100001",
  53974=>"100000010",
  53975=>"000001000",
  53976=>"100001101",
  53977=>"111110111",
  53978=>"111101010",
  53979=>"000000111",
  53980=>"100110101",
  53981=>"001110011",
  53982=>"101100000",
  53983=>"111110110",
  53984=>"101100001",
  53985=>"101111111",
  53986=>"110100111",
  53987=>"110100001",
  53988=>"010000000",
  53989=>"110101000",
  53990=>"001100001",
  53991=>"011111110",
  53992=>"010110111",
  53993=>"010001001",
  53994=>"000101100",
  53995=>"001111111",
  53996=>"011000111",
  53997=>"011001001",
  53998=>"010001010",
  53999=>"000010001",
  54000=>"001111011",
  54001=>"111110101",
  54002=>"000101001",
  54003=>"101100111",
  54004=>"011000010",
  54005=>"000111100",
  54006=>"101101001",
  54007=>"000010100",
  54008=>"010000111",
  54009=>"110111001",
  54010=>"001110000",
  54011=>"010100111",
  54012=>"100110001",
  54013=>"111110110",
  54014=>"110100010",
  54015=>"101000101",
  54016=>"100010000",
  54017=>"011011111",
  54018=>"101111100",
  54019=>"110110000",
  54020=>"111111111",
  54021=>"000010110",
  54022=>"100100001",
  54023=>"111110010",
  54024=>"001101110",
  54025=>"011101100",
  54026=>"000011001",
  54027=>"010111010",
  54028=>"001100110",
  54029=>"010111010",
  54030=>"000010101",
  54031=>"010111000",
  54032=>"010111101",
  54033=>"111111100",
  54034=>"110111011",
  54035=>"001111000",
  54036=>"000111011",
  54037=>"011011100",
  54038=>"011000111",
  54039=>"001011110",
  54040=>"100000011",
  54041=>"000010011",
  54042=>"010111101",
  54043=>"010111001",
  54044=>"000110011",
  54045=>"111001111",
  54046=>"101110000",
  54047=>"110011010",
  54048=>"100110000",
  54049=>"010100000",
  54050=>"000001001",
  54051=>"001111110",
  54052=>"111100001",
  54053=>"111011100",
  54054=>"111011101",
  54055=>"110110000",
  54056=>"010110010",
  54057=>"000010101",
  54058=>"111000010",
  54059=>"001110001",
  54060=>"110111001",
  54061=>"001011111",
  54062=>"101110001",
  54063=>"001110000",
  54064=>"010101101",
  54065=>"011111100",
  54066=>"101111111",
  54067=>"010110010",
  54068=>"110000001",
  54069=>"111010111",
  54070=>"100110100",
  54071=>"100000111",
  54072=>"011011110",
  54073=>"100110101",
  54074=>"011010010",
  54075=>"000110011",
  54076=>"100000000",
  54077=>"000000000",
  54078=>"100101110",
  54079=>"110101110",
  54080=>"100110011",
  54081=>"111000010",
  54082=>"110011011",
  54083=>"111101011",
  54084=>"000000000",
  54085=>"000000000",
  54086=>"100110010",
  54087=>"000100011",
  54088=>"011110100",
  54089=>"010011001",
  54090=>"110111010",
  54091=>"001001101",
  54092=>"001001100",
  54093=>"011000000",
  54094=>"000010001",
  54095=>"000100110",
  54096=>"001110011",
  54097=>"101010000",
  54098=>"101011101",
  54099=>"101011110",
  54100=>"000010010",
  54101=>"100010100",
  54102=>"001010100",
  54103=>"000100010",
  54104=>"001001010",
  54105=>"111011101",
  54106=>"110100100",
  54107=>"000101000",
  54108=>"001110111",
  54109=>"001001001",
  54110=>"011100101",
  54111=>"111111101",
  54112=>"010000011",
  54113=>"111110101",
  54114=>"010010001",
  54115=>"100001101",
  54116=>"100011111",
  54117=>"000000010",
  54118=>"111001001",
  54119=>"010000010",
  54120=>"011101111",
  54121=>"000110101",
  54122=>"011010001",
  54123=>"111001101",
  54124=>"111001000",
  54125=>"011000110",
  54126=>"101110010",
  54127=>"010110010",
  54128=>"100011110",
  54129=>"111001101",
  54130=>"111010111",
  54131=>"101000001",
  54132=>"011010001",
  54133=>"110010010",
  54134=>"100101001",
  54135=>"110100001",
  54136=>"000001101",
  54137=>"000010100",
  54138=>"011001101",
  54139=>"110011100",
  54140=>"010100010",
  54141=>"001111100",
  54142=>"010011001",
  54143=>"111001100",
  54144=>"001010001",
  54145=>"000011010",
  54146=>"011110010",
  54147=>"100111101",
  54148=>"110110111",
  54149=>"101000110",
  54150=>"100011100",
  54151=>"011100101",
  54152=>"011011100",
  54153=>"010011100",
  54154=>"110100101",
  54155=>"101001111",
  54156=>"101011010",
  54157=>"110101010",
  54158=>"100010000",
  54159=>"000100101",
  54160=>"111101101",
  54161=>"110001011",
  54162=>"101011000",
  54163=>"100001100",
  54164=>"011110010",
  54165=>"000110011",
  54166=>"111001100",
  54167=>"000100000",
  54168=>"000011000",
  54169=>"111010110",
  54170=>"111011111",
  54171=>"011010001",
  54172=>"000000100",
  54173=>"100101010",
  54174=>"001110010",
  54175=>"010111010",
  54176=>"101110111",
  54177=>"011111010",
  54178=>"100101101",
  54179=>"110000100",
  54180=>"011100110",
  54181=>"011101010",
  54182=>"010010011",
  54183=>"110110010",
  54184=>"111111111",
  54185=>"011011110",
  54186=>"001101010",
  54187=>"010001100",
  54188=>"011100110",
  54189=>"000001001",
  54190=>"101001000",
  54191=>"101001100",
  54192=>"100001011",
  54193=>"100000101",
  54194=>"111000100",
  54195=>"101101000",
  54196=>"110101111",
  54197=>"011110010",
  54198=>"010111101",
  54199=>"110011000",
  54200=>"001010100",
  54201=>"010000101",
  54202=>"110111110",
  54203=>"101000011",
  54204=>"110111010",
  54205=>"010101101",
  54206=>"000100000",
  54207=>"101010111",
  54208=>"111111111",
  54209=>"110000010",
  54210=>"100111001",
  54211=>"111100000",
  54212=>"101111010",
  54213=>"000110001",
  54214=>"010101101",
  54215=>"100000000",
  54216=>"000011000",
  54217=>"110111110",
  54218=>"000001000",
  54219=>"110101001",
  54220=>"110001101",
  54221=>"110101011",
  54222=>"000111111",
  54223=>"101001110",
  54224=>"000010111",
  54225=>"001001101",
  54226=>"000011011",
  54227=>"000101011",
  54228=>"111111110",
  54229=>"101011010",
  54230=>"110010101",
  54231=>"101110111",
  54232=>"000101110",
  54233=>"110101110",
  54234=>"010111111",
  54235=>"000001111",
  54236=>"111100101",
  54237=>"111100011",
  54238=>"000010111",
  54239=>"101000011",
  54240=>"111111011",
  54241=>"001100010",
  54242=>"010011101",
  54243=>"011001111",
  54244=>"111000011",
  54245=>"000010010",
  54246=>"110100000",
  54247=>"010000110",
  54248=>"000000111",
  54249=>"101010001",
  54250=>"100001001",
  54251=>"000101100",
  54252=>"011110000",
  54253=>"011101000",
  54254=>"111000100",
  54255=>"011101011",
  54256=>"101000001",
  54257=>"100010001",
  54258=>"001001011",
  54259=>"101101000",
  54260=>"110011010",
  54261=>"001010100",
  54262=>"111001110",
  54263=>"111000100",
  54264=>"010101100",
  54265=>"101000101",
  54266=>"100101001",
  54267=>"010111110",
  54268=>"101101101",
  54269=>"110101011",
  54270=>"000000100",
  54271=>"000100101",
  54272=>"101101101",
  54273=>"011001010",
  54274=>"100011101",
  54275=>"010110000",
  54276=>"001111011",
  54277=>"011001010",
  54278=>"100100100",
  54279=>"010101100",
  54280=>"011001110",
  54281=>"100110001",
  54282=>"101110001",
  54283=>"100101110",
  54284=>"100110111",
  54285=>"010111110",
  54286=>"110110111",
  54287=>"111011011",
  54288=>"111011110",
  54289=>"011000100",
  54290=>"011110011",
  54291=>"011110001",
  54292=>"111101000",
  54293=>"100100010",
  54294=>"001001010",
  54295=>"010100110",
  54296=>"000111001",
  54297=>"010001011",
  54298=>"011011011",
  54299=>"101111010",
  54300=>"111101011",
  54301=>"100100011",
  54302=>"101111111",
  54303=>"001111111",
  54304=>"011111001",
  54305=>"111001001",
  54306=>"110010000",
  54307=>"011010111",
  54308=>"000011100",
  54309=>"101000101",
  54310=>"101110110",
  54311=>"011011001",
  54312=>"101010010",
  54313=>"101111111",
  54314=>"110111111",
  54315=>"100110001",
  54316=>"001101001",
  54317=>"111011110",
  54318=>"110010000",
  54319=>"111101001",
  54320=>"001000001",
  54321=>"101110000",
  54322=>"111001101",
  54323=>"101100010",
  54324=>"011001101",
  54325=>"011100011",
  54326=>"101100111",
  54327=>"101000111",
  54328=>"001101100",
  54329=>"101100110",
  54330=>"110100011",
  54331=>"100011000",
  54332=>"110010101",
  54333=>"001101010",
  54334=>"100101000",
  54335=>"111011010",
  54336=>"010100110",
  54337=>"000011101",
  54338=>"100000001",
  54339=>"111000010",
  54340=>"010010100",
  54341=>"101100110",
  54342=>"111001001",
  54343=>"111000101",
  54344=>"011001110",
  54345=>"000001000",
  54346=>"010000000",
  54347=>"011010100",
  54348=>"101000010",
  54349=>"001101011",
  54350=>"010100110",
  54351=>"010011111",
  54352=>"000010001",
  54353=>"100110101",
  54354=>"110111001",
  54355=>"100000100",
  54356=>"000100010",
  54357=>"100000100",
  54358=>"100000100",
  54359=>"101110001",
  54360=>"110100010",
  54361=>"001111111",
  54362=>"000100101",
  54363=>"001111111",
  54364=>"000010000",
  54365=>"101110101",
  54366=>"001000010",
  54367=>"111010100",
  54368=>"000001010",
  54369=>"010100101",
  54370=>"100100010",
  54371=>"101110011",
  54372=>"011101011",
  54373=>"110011110",
  54374=>"111111111",
  54375=>"111010100",
  54376=>"010111000",
  54377=>"111111101",
  54378=>"110100010",
  54379=>"111111010",
  54380=>"010000000",
  54381=>"000100011",
  54382=>"010000001",
  54383=>"110010111",
  54384=>"110100000",
  54385=>"100000111",
  54386=>"100111111",
  54387=>"110100100",
  54388=>"000000101",
  54389=>"101011001",
  54390=>"001110011",
  54391=>"001000100",
  54392=>"000010100",
  54393=>"111011011",
  54394=>"010110000",
  54395=>"011001101",
  54396=>"011011000",
  54397=>"101100100",
  54398=>"010000010",
  54399=>"011111111",
  54400=>"011111100",
  54401=>"000101010",
  54402=>"111111011",
  54403=>"010101000",
  54404=>"001001000",
  54405=>"111000110",
  54406=>"100000001",
  54407=>"000100101",
  54408=>"001000001",
  54409=>"010000111",
  54410=>"001100111",
  54411=>"001111001",
  54412=>"101111000",
  54413=>"101001000",
  54414=>"100000010",
  54415=>"100001000",
  54416=>"000010011",
  54417=>"000100001",
  54418=>"110001000",
  54419=>"111101011",
  54420=>"101010100",
  54421=>"011011111",
  54422=>"111010111",
  54423=>"101111111",
  54424=>"100001110",
  54425=>"011001001",
  54426=>"111111110",
  54427=>"101101101",
  54428=>"100100111",
  54429=>"110000111",
  54430=>"000101100",
  54431=>"110110011",
  54432=>"000111101",
  54433=>"001010110",
  54434=>"100100000",
  54435=>"010101101",
  54436=>"100101000",
  54437=>"110011101",
  54438=>"001011111",
  54439=>"101001110",
  54440=>"000110110",
  54441=>"011011001",
  54442=>"110111001",
  54443=>"111101011",
  54444=>"101110100",
  54445=>"100101111",
  54446=>"101111111",
  54447=>"000111100",
  54448=>"111101011",
  54449=>"100000000",
  54450=>"111100001",
  54451=>"110001110",
  54452=>"111010101",
  54453=>"000101000",
  54454=>"000001111",
  54455=>"100111100",
  54456=>"001111100",
  54457=>"110101111",
  54458=>"110011101",
  54459=>"100110000",
  54460=>"000110111",
  54461=>"111001110",
  54462=>"101010111",
  54463=>"110100110",
  54464=>"111110101",
  54465=>"110001111",
  54466=>"000100000",
  54467=>"010011011",
  54468=>"001011110",
  54469=>"110000001",
  54470=>"101010010",
  54471=>"001100111",
  54472=>"001111100",
  54473=>"010111011",
  54474=>"101101110",
  54475=>"001110110",
  54476=>"000000111",
  54477=>"000000000",
  54478=>"100000010",
  54479=>"001011000",
  54480=>"000101011",
  54481=>"111110111",
  54482=>"000011100",
  54483=>"101101100",
  54484=>"101011111",
  54485=>"011111000",
  54486=>"100010001",
  54487=>"010010000",
  54488=>"111000001",
  54489=>"101001011",
  54490=>"100001111",
  54491=>"111001110",
  54492=>"010011010",
  54493=>"001110000",
  54494=>"000100100",
  54495=>"101100000",
  54496=>"100100100",
  54497=>"100000001",
  54498=>"100010111",
  54499=>"000001001",
  54500=>"011110001",
  54501=>"011001001",
  54502=>"110111000",
  54503=>"000010010",
  54504=>"110101000",
  54505=>"100000001",
  54506=>"101000110",
  54507=>"100011011",
  54508=>"011100101",
  54509=>"111110110",
  54510=>"100000100",
  54511=>"010001000",
  54512=>"111010000",
  54513=>"101010010",
  54514=>"011101110",
  54515=>"110110001",
  54516=>"110111111",
  54517=>"000100101",
  54518=>"110100010",
  54519=>"000000101",
  54520=>"101001000",
  54521=>"111110001",
  54522=>"011001100",
  54523=>"000110011",
  54524=>"001100011",
  54525=>"110001111",
  54526=>"110011010",
  54527=>"100110010",
  54528=>"100000110",
  54529=>"100001101",
  54530=>"010011001",
  54531=>"111001111",
  54532=>"110001001",
  54533=>"010000001",
  54534=>"010010101",
  54535=>"011010101",
  54536=>"010000100",
  54537=>"111001010",
  54538=>"100110101",
  54539=>"001001011",
  54540=>"001111001",
  54541=>"110111111",
  54542=>"101111110",
  54543=>"010101011",
  54544=>"111000101",
  54545=>"100001111",
  54546=>"100011001",
  54547=>"000100011",
  54548=>"101101000",
  54549=>"001110001",
  54550=>"111011111",
  54551=>"101101011",
  54552=>"001001101",
  54553=>"011001001",
  54554=>"010110101",
  54555=>"000100000",
  54556=>"000101101",
  54557=>"010110011",
  54558=>"100110000",
  54559=>"111111100",
  54560=>"110000011",
  54561=>"000001010",
  54562=>"110101100",
  54563=>"001100010",
  54564=>"010000001",
  54565=>"010000100",
  54566=>"011100010",
  54567=>"001110011",
  54568=>"001001011",
  54569=>"101111101",
  54570=>"101100011",
  54571=>"111000000",
  54572=>"010100100",
  54573=>"111111101",
  54574=>"111011001",
  54575=>"010110110",
  54576=>"111000110",
  54577=>"100101101",
  54578=>"011010110",
  54579=>"101010001",
  54580=>"001001011",
  54581=>"010110000",
  54582=>"111111111",
  54583=>"001100010",
  54584=>"000001100",
  54585=>"101000111",
  54586=>"111111100",
  54587=>"111000001",
  54588=>"101000100",
  54589=>"100111010",
  54590=>"001001001",
  54591=>"010100100",
  54592=>"101001011",
  54593=>"110011101",
  54594=>"111010001",
  54595=>"101000100",
  54596=>"101001101",
  54597=>"011000110",
  54598=>"100011000",
  54599=>"000011001",
  54600=>"101011010",
  54601=>"001101001",
  54602=>"101001011",
  54603=>"010000111",
  54604=>"110001101",
  54605=>"110110011",
  54606=>"100001100",
  54607=>"001001101",
  54608=>"100101110",
  54609=>"101101110",
  54610=>"110001110",
  54611=>"111011101",
  54612=>"000000111",
  54613=>"011111010",
  54614=>"001000100",
  54615=>"010101011",
  54616=>"100110001",
  54617=>"110011101",
  54618=>"010001100",
  54619=>"111000111",
  54620=>"110011011",
  54621=>"111111100",
  54622=>"111100110",
  54623=>"101111011",
  54624=>"101100110",
  54625=>"110110000",
  54626=>"011110011",
  54627=>"011111101",
  54628=>"111100011",
  54629=>"001011001",
  54630=>"000010111",
  54631=>"001000001",
  54632=>"101001011",
  54633=>"101110000",
  54634=>"010101100",
  54635=>"100011001",
  54636=>"001000000",
  54637=>"100100001",
  54638=>"000110100",
  54639=>"000001010",
  54640=>"101111001",
  54641=>"110000000",
  54642=>"100111111",
  54643=>"000111011",
  54644=>"101111111",
  54645=>"000101100",
  54646=>"110011111",
  54647=>"110010001",
  54648=>"100011100",
  54649=>"010001101",
  54650=>"111100101",
  54651=>"100000100",
  54652=>"100111000",
  54653=>"110000110",
  54654=>"001011001",
  54655=>"100011010",
  54656=>"010000000",
  54657=>"011111001",
  54658=>"011101001",
  54659=>"100000111",
  54660=>"101001100",
  54661=>"001100100",
  54662=>"001100001",
  54663=>"011111101",
  54664=>"010100110",
  54665=>"011101100",
  54666=>"110010111",
  54667=>"001011010",
  54668=>"101011111",
  54669=>"000111101",
  54670=>"100101111",
  54671=>"000111010",
  54672=>"100110100",
  54673=>"010010001",
  54674=>"111001100",
  54675=>"000010010",
  54676=>"000100010",
  54677=>"101111101",
  54678=>"110100100",
  54679=>"011000110",
  54680=>"001000101",
  54681=>"011011110",
  54682=>"111100110",
  54683=>"000111111",
  54684=>"111000000",
  54685=>"110101001",
  54686=>"110101110",
  54687=>"000011101",
  54688=>"000101100",
  54689=>"011001110",
  54690=>"010100100",
  54691=>"100011011",
  54692=>"001010110",
  54693=>"000111000",
  54694=>"100110111",
  54695=>"001100111",
  54696=>"100001000",
  54697=>"011000101",
  54698=>"001101100",
  54699=>"110011110",
  54700=>"011100101",
  54701=>"010010111",
  54702=>"111101010",
  54703=>"110010110",
  54704=>"111110110",
  54705=>"010011011",
  54706=>"111010011",
  54707=>"011101010",
  54708=>"000010010",
  54709=>"011010110",
  54710=>"101101000",
  54711=>"001001110",
  54712=>"000000111",
  54713=>"000011010",
  54714=>"000000111",
  54715=>"111000101",
  54716=>"000001011",
  54717=>"100101001",
  54718=>"001010110",
  54719=>"001111000",
  54720=>"001000100",
  54721=>"001110011",
  54722=>"011111011",
  54723=>"101010111",
  54724=>"000001000",
  54725=>"100010101",
  54726=>"011101000",
  54727=>"100001101",
  54728=>"111010111",
  54729=>"100111011",
  54730=>"000101000",
  54731=>"100011010",
  54732=>"000011000",
  54733=>"110111001",
  54734=>"000100010",
  54735=>"011000100",
  54736=>"011100000",
  54737=>"101110011",
  54738=>"100101110",
  54739=>"101010101",
  54740=>"010110000",
  54741=>"110010010",
  54742=>"001000101",
  54743=>"000011010",
  54744=>"100011000",
  54745=>"001110100",
  54746=>"101010011",
  54747=>"001011011",
  54748=>"101010001",
  54749=>"011101000",
  54750=>"111010111",
  54751=>"101001000",
  54752=>"001101001",
  54753=>"010000011",
  54754=>"011001111",
  54755=>"110010001",
  54756=>"011010001",
  54757=>"000010011",
  54758=>"010011011",
  54759=>"000001101",
  54760=>"001010001",
  54761=>"101100001",
  54762=>"100011100",
  54763=>"110000000",
  54764=>"010000101",
  54765=>"101110000",
  54766=>"000010000",
  54767=>"001011011",
  54768=>"011111101",
  54769=>"110010000",
  54770=>"100010010",
  54771=>"010001010",
  54772=>"111110110",
  54773=>"001010001",
  54774=>"100111001",
  54775=>"101010111",
  54776=>"010110100",
  54777=>"110011011",
  54778=>"000111111",
  54779=>"010111001",
  54780=>"110111010",
  54781=>"111011010",
  54782=>"001100000",
  54783=>"001001010",
  54784=>"100001011",
  54785=>"011000011",
  54786=>"100001011",
  54787=>"011010111",
  54788=>"000000000",
  54789=>"010000111",
  54790=>"111100111",
  54791=>"111001110",
  54792=>"111000111",
  54793=>"100100010",
  54794=>"001101110",
  54795=>"101100101",
  54796=>"010110000",
  54797=>"100010111",
  54798=>"101111010",
  54799=>"101101000",
  54800=>"011010011",
  54801=>"000100011",
  54802=>"100111000",
  54803=>"000010111",
  54804=>"100100101",
  54805=>"010100000",
  54806=>"011010101",
  54807=>"111011000",
  54808=>"100000101",
  54809=>"111011100",
  54810=>"010110010",
  54811=>"001010000",
  54812=>"111010011",
  54813=>"010111010",
  54814=>"000110110",
  54815=>"100000011",
  54816=>"101110100",
  54817=>"111000000",
  54818=>"001100010",
  54819=>"000010111",
  54820=>"000101000",
  54821=>"100110111",
  54822=>"110000000",
  54823=>"000111001",
  54824=>"111100000",
  54825=>"011111011",
  54826=>"000100011",
  54827=>"111010011",
  54828=>"111011010",
  54829=>"111100100",
  54830=>"101111101",
  54831=>"010111111",
  54832=>"110101100",
  54833=>"110010010",
  54834=>"111000001",
  54835=>"000100101",
  54836=>"101101101",
  54837=>"000100011",
  54838=>"001000101",
  54839=>"101011111",
  54840=>"010000011",
  54841=>"111111110",
  54842=>"000101110",
  54843=>"110001100",
  54844=>"111110000",
  54845=>"100000111",
  54846=>"110001111",
  54847=>"000001010",
  54848=>"001101100",
  54849=>"010111101",
  54850=>"100101101",
  54851=>"110111001",
  54852=>"001011000",
  54853=>"000111001",
  54854=>"000011101",
  54855=>"010111100",
  54856=>"001101100",
  54857=>"111100001",
  54858=>"001111000",
  54859=>"001001110",
  54860=>"110001100",
  54861=>"101000001",
  54862=>"010010100",
  54863=>"101010111",
  54864=>"110110111",
  54865=>"001011000",
  54866=>"001110110",
  54867=>"111100111",
  54868=>"001110101",
  54869=>"001001001",
  54870=>"111110111",
  54871=>"010111111",
  54872=>"101110000",
  54873=>"001001101",
  54874=>"011100010",
  54875=>"011010101",
  54876=>"010101111",
  54877=>"101011001",
  54878=>"111111110",
  54879=>"011011011",
  54880=>"110101110",
  54881=>"111101111",
  54882=>"010010011",
  54883=>"000000011",
  54884=>"110100010",
  54885=>"000111001",
  54886=>"000110011",
  54887=>"101110011",
  54888=>"011100111",
  54889=>"010111011",
  54890=>"000000000",
  54891=>"101011101",
  54892=>"111100010",
  54893=>"100010111",
  54894=>"101000100",
  54895=>"110011101",
  54896=>"001000001",
  54897=>"101010000",
  54898=>"100110000",
  54899=>"100101110",
  54900=>"111001011",
  54901=>"001011110",
  54902=>"011011110",
  54903=>"100011111",
  54904=>"011011101",
  54905=>"111000101",
  54906=>"000001000",
  54907=>"000011110",
  54908=>"111100001",
  54909=>"010001111",
  54910=>"000000010",
  54911=>"011111001",
  54912=>"000101110",
  54913=>"000010110",
  54914=>"001001010",
  54915=>"110101100",
  54916=>"111100010",
  54917=>"100110011",
  54918=>"000000110",
  54919=>"000100111",
  54920=>"001110101",
  54921=>"101111000",
  54922=>"001110010",
  54923=>"110110001",
  54924=>"010011101",
  54925=>"110111101",
  54926=>"100001110",
  54927=>"101110101",
  54928=>"100110111",
  54929=>"010111011",
  54930=>"111001100",
  54931=>"001000011",
  54932=>"110100001",
  54933=>"101111101",
  54934=>"000111111",
  54935=>"110011100",
  54936=>"100100100",
  54937=>"010110011",
  54938=>"000101000",
  54939=>"001010011",
  54940=>"011000100",
  54941=>"101110110",
  54942=>"001101101",
  54943=>"001110001",
  54944=>"110111101",
  54945=>"111001111",
  54946=>"101011000",
  54947=>"010100101",
  54948=>"010110010",
  54949=>"100010000",
  54950=>"100110001",
  54951=>"010000110",
  54952=>"011110111",
  54953=>"010011100",
  54954=>"100010100",
  54955=>"010000011",
  54956=>"010000001",
  54957=>"000001101",
  54958=>"101010000",
  54959=>"101000100",
  54960=>"001011001",
  54961=>"010111000",
  54962=>"110000101",
  54963=>"101101100",
  54964=>"110110111",
  54965=>"110111111",
  54966=>"000110110",
  54967=>"000100010",
  54968=>"001011010",
  54969=>"011110111",
  54970=>"100010100",
  54971=>"111000000",
  54972=>"111011010",
  54973=>"001100100",
  54974=>"101010100",
  54975=>"001010000",
  54976=>"100000001",
  54977=>"110110010",
  54978=>"000110000",
  54979=>"110000011",
  54980=>"101110111",
  54981=>"110101110",
  54982=>"011110111",
  54983=>"010101010",
  54984=>"100111010",
  54985=>"011101101",
  54986=>"010110011",
  54987=>"100011011",
  54988=>"010010000",
  54989=>"001100011",
  54990=>"010110010",
  54991=>"001101011",
  54992=>"011101110",
  54993=>"111001010",
  54994=>"100100100",
  54995=>"100110110",
  54996=>"111100101",
  54997=>"101010010",
  54998=>"000011010",
  54999=>"001001000",
  55000=>"010011111",
  55001=>"010000101",
  55002=>"111110100",
  55003=>"010010101",
  55004=>"111101111",
  55005=>"000011101",
  55006=>"110011101",
  55007=>"110100000",
  55008=>"111111011",
  55009=>"111111100",
  55010=>"111100101",
  55011=>"100111100",
  55012=>"000000101",
  55013=>"111010101",
  55014=>"001000011",
  55015=>"000111111",
  55016=>"111111111",
  55017=>"011100110",
  55018=>"000111101",
  55019=>"001000010",
  55020=>"100010001",
  55021=>"001111101",
  55022=>"011101001",
  55023=>"001110001",
  55024=>"100111101",
  55025=>"101011110",
  55026=>"101101001",
  55027=>"111010001",
  55028=>"000010000",
  55029=>"110110001",
  55030=>"010111101",
  55031=>"111000010",
  55032=>"110100101",
  55033=>"011110100",
  55034=>"110001000",
  55035=>"001101110",
  55036=>"111110100",
  55037=>"101010000",
  55038=>"100111111",
  55039=>"100000110",
  55040=>"001001100",
  55041=>"111111011",
  55042=>"100001101",
  55043=>"101011110",
  55044=>"000000011",
  55045=>"110110010",
  55046=>"111010111",
  55047=>"000101011",
  55048=>"011111110",
  55049=>"011100101",
  55050=>"110101011",
  55051=>"111101111",
  55052=>"110111011",
  55053=>"000001110",
  55054=>"010110110",
  55055=>"100011011",
  55056=>"100100100",
  55057=>"110110110",
  55058=>"011010011",
  55059=>"111011110",
  55060=>"101001101",
  55061=>"001000001",
  55062=>"000000111",
  55063=>"100111111",
  55064=>"011101001",
  55065=>"111100011",
  55066=>"010001000",
  55067=>"000111110",
  55068=>"001000011",
  55069=>"110001000",
  55070=>"010011011",
  55071=>"000011111",
  55072=>"001111011",
  55073=>"010001000",
  55074=>"010110010",
  55075=>"111110111",
  55076=>"010010000",
  55077=>"100001001",
  55078=>"111110100",
  55079=>"111101101",
  55080=>"101100011",
  55081=>"001100000",
  55082=>"110010010",
  55083=>"100111001",
  55084=>"111011011",
  55085=>"101111010",
  55086=>"011111011",
  55087=>"100110011",
  55088=>"000111101",
  55089=>"001101100",
  55090=>"101100101",
  55091=>"101101000",
  55092=>"010101010",
  55093=>"110001011",
  55094=>"111010101",
  55095=>"110111001",
  55096=>"001100001",
  55097=>"111101101",
  55098=>"010101100",
  55099=>"100100010",
  55100=>"011110101",
  55101=>"001101100",
  55102=>"011011011",
  55103=>"110110111",
  55104=>"000000001",
  55105=>"001001000",
  55106=>"011101101",
  55107=>"000111010",
  55108=>"110010001",
  55109=>"111001011",
  55110=>"110110111",
  55111=>"011110110",
  55112=>"111110010",
  55113=>"100000111",
  55114=>"001110011",
  55115=>"000000000",
  55116=>"000100010",
  55117=>"001001100",
  55118=>"000101010",
  55119=>"110000000",
  55120=>"000100101",
  55121=>"000111011",
  55122=>"111111110",
  55123=>"000110101",
  55124=>"110001000",
  55125=>"101100101",
  55126=>"011001000",
  55127=>"100110001",
  55128=>"011110000",
  55129=>"110110001",
  55130=>"001001100",
  55131=>"111011100",
  55132=>"010001000",
  55133=>"101110011",
  55134=>"111001101",
  55135=>"101001010",
  55136=>"000100111",
  55137=>"110000110",
  55138=>"110011001",
  55139=>"111101000",
  55140=>"011001110",
  55141=>"010101111",
  55142=>"101001001",
  55143=>"000011010",
  55144=>"111100001",
  55145=>"111001010",
  55146=>"010110101",
  55147=>"101111011",
  55148=>"110111001",
  55149=>"011010110",
  55150=>"101101111",
  55151=>"001101000",
  55152=>"011000100",
  55153=>"000011001",
  55154=>"111111110",
  55155=>"101001101",
  55156=>"110000110",
  55157=>"000100000",
  55158=>"000100000",
  55159=>"100100010",
  55160=>"011011110",
  55161=>"010001011",
  55162=>"100110011",
  55163=>"111010010",
  55164=>"100111001",
  55165=>"101101111",
  55166=>"000111101",
  55167=>"100111110",
  55168=>"000001111",
  55169=>"011011011",
  55170=>"101100111",
  55171=>"011101011",
  55172=>"110100100",
  55173=>"110100011",
  55174=>"000010111",
  55175=>"111110011",
  55176=>"101110100",
  55177=>"010101001",
  55178=>"000010100",
  55179=>"011101011",
  55180=>"100011111",
  55181=>"010001111",
  55182=>"000011001",
  55183=>"010110111",
  55184=>"111000101",
  55185=>"000111110",
  55186=>"000000101",
  55187=>"111100011",
  55188=>"011010111",
  55189=>"001011100",
  55190=>"110101000",
  55191=>"100000010",
  55192=>"001000101",
  55193=>"101101110",
  55194=>"100000001",
  55195=>"111111011",
  55196=>"111111101",
  55197=>"111111011",
  55198=>"010001001",
  55199=>"011010101",
  55200=>"010011100",
  55201=>"011001010",
  55202=>"001111001",
  55203=>"101101100",
  55204=>"100110110",
  55205=>"100100111",
  55206=>"100110001",
  55207=>"101110010",
  55208=>"000100100",
  55209=>"010100101",
  55210=>"011111111",
  55211=>"110001010",
  55212=>"000100100",
  55213=>"101100111",
  55214=>"101001101",
  55215=>"100110001",
  55216=>"010110000",
  55217=>"010110110",
  55218=>"011100000",
  55219=>"100010000",
  55220=>"110110110",
  55221=>"011111011",
  55222=>"110010110",
  55223=>"110100000",
  55224=>"111101110",
  55225=>"010011110",
  55226=>"110111111",
  55227=>"111111110",
  55228=>"010011001",
  55229=>"000100001",
  55230=>"110000000",
  55231=>"011000010",
  55232=>"100101000",
  55233=>"001001110",
  55234=>"100100110",
  55235=>"110010000",
  55236=>"001000010",
  55237=>"100100101",
  55238=>"010110111",
  55239=>"101000001",
  55240=>"101010000",
  55241=>"101111010",
  55242=>"000101110",
  55243=>"110100001",
  55244=>"110111010",
  55245=>"111111011",
  55246=>"100100111",
  55247=>"001011000",
  55248=>"101010010",
  55249=>"000101001",
  55250=>"001101100",
  55251=>"000101101",
  55252=>"011000101",
  55253=>"111011111",
  55254=>"100010111",
  55255=>"101000111",
  55256=>"010100101",
  55257=>"000010100",
  55258=>"111100011",
  55259=>"001000100",
  55260=>"111101111",
  55261=>"101101111",
  55262=>"100101110",
  55263=>"100000110",
  55264=>"110101010",
  55265=>"111001101",
  55266=>"110111011",
  55267=>"010101110",
  55268=>"000110101",
  55269=>"000111100",
  55270=>"110011010",
  55271=>"011110101",
  55272=>"010010001",
  55273=>"100111011",
  55274=>"100111101",
  55275=>"111101100",
  55276=>"101110111",
  55277=>"111110100",
  55278=>"100110010",
  55279=>"101011011",
  55280=>"000000010",
  55281=>"110011101",
  55282=>"000000010",
  55283=>"111010100",
  55284=>"100111101",
  55285=>"011101011",
  55286=>"111101111",
  55287=>"101001000",
  55288=>"010110111",
  55289=>"010001110",
  55290=>"001101000",
  55291=>"110001101",
  55292=>"110001101",
  55293=>"001101100",
  55294=>"100100100",
  55295=>"100100110",
  55296=>"100110111",
  55297=>"011001110",
  55298=>"111011001",
  55299=>"000010101",
  55300=>"101101011",
  55301=>"000000111",
  55302=>"111000001",
  55303=>"101001010",
  55304=>"101101010",
  55305=>"001101111",
  55306=>"110110011",
  55307=>"100000111",
  55308=>"010110010",
  55309=>"100101110",
  55310=>"000000100",
  55311=>"100011001",
  55312=>"110101101",
  55313=>"111111000",
  55314=>"110010001",
  55315=>"001000101",
  55316=>"111101000",
  55317=>"000010010",
  55318=>"100111010",
  55319=>"100111100",
  55320=>"000110010",
  55321=>"100100111",
  55322=>"000101110",
  55323=>"000110101",
  55324=>"101010000",
  55325=>"100010101",
  55326=>"111110111",
  55327=>"101001011",
  55328=>"111100011",
  55329=>"100010010",
  55330=>"010111111",
  55331=>"110000011",
  55332=>"000011101",
  55333=>"101100000",
  55334=>"111010110",
  55335=>"110100110",
  55336=>"110101110",
  55337=>"011010111",
  55338=>"101100111",
  55339=>"010000001",
  55340=>"001000010",
  55341=>"110100000",
  55342=>"100011010",
  55343=>"000100100",
  55344=>"111111011",
  55345=>"110000010",
  55346=>"001011000",
  55347=>"110110110",
  55348=>"011001000",
  55349=>"100100000",
  55350=>"110110101",
  55351=>"000100111",
  55352=>"010111011",
  55353=>"101110101",
  55354=>"010000111",
  55355=>"101000100",
  55356=>"001111000",
  55357=>"101101111",
  55358=>"110011000",
  55359=>"010010000",
  55360=>"011001100",
  55361=>"001011101",
  55362=>"010010100",
  55363=>"111111100",
  55364=>"101111111",
  55365=>"100100110",
  55366=>"110000011",
  55367=>"011100001",
  55368=>"010000001",
  55369=>"010111010",
  55370=>"010101111",
  55371=>"001111111",
  55372=>"011100010",
  55373=>"010000011",
  55374=>"110111010",
  55375=>"100010011",
  55376=>"011000000",
  55377=>"100000100",
  55378=>"101100010",
  55379=>"111001101",
  55380=>"010101110",
  55381=>"110000101",
  55382=>"010000010",
  55383=>"011100000",
  55384=>"111100101",
  55385=>"000011100",
  55386=>"100010110",
  55387=>"100100100",
  55388=>"001100001",
  55389=>"001110111",
  55390=>"010101000",
  55391=>"010110011",
  55392=>"010010110",
  55393=>"010011001",
  55394=>"001010100",
  55395=>"011111001",
  55396=>"100001000",
  55397=>"011100001",
  55398=>"101001101",
  55399=>"000101101",
  55400=>"100100110",
  55401=>"100000001",
  55402=>"001100001",
  55403=>"100110010",
  55404=>"000011111",
  55405=>"010000001",
  55406=>"001000000",
  55407=>"101110011",
  55408=>"110010000",
  55409=>"101000010",
  55410=>"111100101",
  55411=>"001101000",
  55412=>"100010101",
  55413=>"110000000",
  55414=>"001000010",
  55415=>"001111001",
  55416=>"001010100",
  55417=>"101011011",
  55418=>"010001100",
  55419=>"001101011",
  55420=>"001100000",
  55421=>"011101010",
  55422=>"101100011",
  55423=>"101010000",
  55424=>"101100101",
  55425=>"000100111",
  55426=>"010101010",
  55427=>"010100101",
  55428=>"111000101",
  55429=>"001100011",
  55430=>"100010011",
  55431=>"101001000",
  55432=>"111111011",
  55433=>"000101101",
  55434=>"010101100",
  55435=>"010010001",
  55436=>"100001001",
  55437=>"110101111",
  55438=>"100010111",
  55439=>"101100011",
  55440=>"111101101",
  55441=>"000011001",
  55442=>"010001000",
  55443=>"001100111",
  55444=>"011101001",
  55445=>"011001100",
  55446=>"100100011",
  55447=>"010000000",
  55448=>"111101101",
  55449=>"001011100",
  55450=>"011111000",
  55451=>"000101111",
  55452=>"110110111",
  55453=>"100001111",
  55454=>"001100100",
  55455=>"100111111",
  55456=>"000110010",
  55457=>"110110001",
  55458=>"100110101",
  55459=>"000001000",
  55460=>"000110001",
  55461=>"110000100",
  55462=>"101110010",
  55463=>"101011101",
  55464=>"010101010",
  55465=>"000100001",
  55466=>"101111110",
  55467=>"011111011",
  55468=>"111111110",
  55469=>"010000100",
  55470=>"101000000",
  55471=>"101110010",
  55472=>"001011100",
  55473=>"100110101",
  55474=>"001010100",
  55475=>"001001010",
  55476=>"101101001",
  55477=>"011001001",
  55478=>"000100010",
  55479=>"011110000",
  55480=>"100000100",
  55481=>"110101110",
  55482=>"001000010",
  55483=>"111111110",
  55484=>"110010100",
  55485=>"001001010",
  55486=>"101110101",
  55487=>"001000101",
  55488=>"010010001",
  55489=>"001001111",
  55490=>"111011001",
  55491=>"001001000",
  55492=>"100000100",
  55493=>"111111001",
  55494=>"101111111",
  55495=>"000101111",
  55496=>"000101001",
  55497=>"110000001",
  55498=>"111100100",
  55499=>"001010000",
  55500=>"001000000",
  55501=>"011001001",
  55502=>"111001000",
  55503=>"000010100",
  55504=>"100001100",
  55505=>"000000100",
  55506=>"101100110",
  55507=>"000000011",
  55508=>"101010101",
  55509=>"100011000",
  55510=>"000011010",
  55511=>"111111001",
  55512=>"000110001",
  55513=>"000110100",
  55514=>"110100011",
  55515=>"001000000",
  55516=>"010111110",
  55517=>"000101111",
  55518=>"001110011",
  55519=>"000000100",
  55520=>"101010000",
  55521=>"010000100",
  55522=>"010010111",
  55523=>"100100001",
  55524=>"110011010",
  55525=>"111010100",
  55526=>"100101100",
  55527=>"111111111",
  55528=>"110110010",
  55529=>"100001001",
  55530=>"010011100",
  55531=>"001101010",
  55532=>"100111110",
  55533=>"100101111",
  55534=>"101110110",
  55535=>"010100000",
  55536=>"110110101",
  55537=>"110011000",
  55538=>"001111001",
  55539=>"000100110",
  55540=>"011101000",
  55541=>"111011110",
  55542=>"001011010",
  55543=>"001001101",
  55544=>"000101001",
  55545=>"100111111",
  55546=>"100100111",
  55547=>"011000111",
  55548=>"010000001",
  55549=>"101100101",
  55550=>"010111000",
  55551=>"000100100",
  55552=>"001000000",
  55553=>"010000011",
  55554=>"010011001",
  55555=>"101110001",
  55556=>"100010110",
  55557=>"000011000",
  55558=>"011100100",
  55559=>"000101100",
  55560=>"111001011",
  55561=>"001000011",
  55562=>"111110010",
  55563=>"001001100",
  55564=>"101001010",
  55565=>"010011100",
  55566=>"110001110",
  55567=>"110100100",
  55568=>"001111111",
  55569=>"000100100",
  55570=>"101111111",
  55571=>"000001001",
  55572=>"111110100",
  55573=>"011001001",
  55574=>"101100101",
  55575=>"111011110",
  55576=>"110010101",
  55577=>"010100100",
  55578=>"000111110",
  55579=>"110011011",
  55580=>"111111001",
  55581=>"101000111",
  55582=>"000100101",
  55583=>"111111011",
  55584=>"110100110",
  55585=>"100010111",
  55586=>"011001010",
  55587=>"100111100",
  55588=>"101010011",
  55589=>"110011010",
  55590=>"011110101",
  55591=>"100110000",
  55592=>"100101000",
  55593=>"100000001",
  55594=>"001011011",
  55595=>"100010001",
  55596=>"110010111",
  55597=>"111101101",
  55598=>"110010110",
  55599=>"010110101",
  55600=>"001011111",
  55601=>"110100111",
  55602=>"101111101",
  55603=>"101011011",
  55604=>"110111100",
  55605=>"111111110",
  55606=>"000111000",
  55607=>"010101010",
  55608=>"111111110",
  55609=>"111100010",
  55610=>"001111111",
  55611=>"111001110",
  55612=>"001001110",
  55613=>"100111001",
  55614=>"110110000",
  55615=>"100000110",
  55616=>"000111110",
  55617=>"010110000",
  55618=>"011110111",
  55619=>"110011100",
  55620=>"011111111",
  55621=>"101010000",
  55622=>"011100001",
  55623=>"100101110",
  55624=>"111111111",
  55625=>"001000001",
  55626=>"011001000",
  55627=>"000011000",
  55628=>"100101000",
  55629=>"110111010",
  55630=>"111000001",
  55631=>"110011001",
  55632=>"000001001",
  55633=>"000100100",
  55634=>"101101000",
  55635=>"101101110",
  55636=>"000000001",
  55637=>"010111100",
  55638=>"100000111",
  55639=>"000100101",
  55640=>"010000001",
  55641=>"000011101",
  55642=>"010101010",
  55643=>"110100100",
  55644=>"011100100",
  55645=>"010011110",
  55646=>"100111000",
  55647=>"001101101",
  55648=>"111101001",
  55649=>"000010000",
  55650=>"000011000",
  55651=>"100110111",
  55652=>"101100101",
  55653=>"011010101",
  55654=>"010100110",
  55655=>"100000010",
  55656=>"011110101",
  55657=>"001110001",
  55658=>"001010100",
  55659=>"010011010",
  55660=>"001101000",
  55661=>"101111101",
  55662=>"101100101",
  55663=>"101011111",
  55664=>"101110111",
  55665=>"000100000",
  55666=>"001010110",
  55667=>"101011011",
  55668=>"000001011",
  55669=>"101011110",
  55670=>"010101010",
  55671=>"011100010",
  55672=>"111100111",
  55673=>"010110111",
  55674=>"010100011",
  55675=>"101101110",
  55676=>"101010110",
  55677=>"001111001",
  55678=>"111001101",
  55679=>"111111001",
  55680=>"010101110",
  55681=>"000010110",
  55682=>"011001100",
  55683=>"110000110",
  55684=>"110010010",
  55685=>"101011100",
  55686=>"000011001",
  55687=>"001100111",
  55688=>"011000011",
  55689=>"100001011",
  55690=>"001111101",
  55691=>"101101101",
  55692=>"111101010",
  55693=>"100000000",
  55694=>"110110000",
  55695=>"001010111",
  55696=>"111110100",
  55697=>"111111100",
  55698=>"100010110",
  55699=>"011010101",
  55700=>"011110000",
  55701=>"010101100",
  55702=>"000011111",
  55703=>"101011000",
  55704=>"100111000",
  55705=>"111000011",
  55706=>"000111100",
  55707=>"000011111",
  55708=>"010111110",
  55709=>"111100111",
  55710=>"010110000",
  55711=>"000000101",
  55712=>"111111001",
  55713=>"000011001",
  55714=>"101000000",
  55715=>"011000110",
  55716=>"001100010",
  55717=>"000101000",
  55718=>"100001000",
  55719=>"000000001",
  55720=>"001001101",
  55721=>"110111100",
  55722=>"101111000",
  55723=>"000111000",
  55724=>"100011011",
  55725=>"101100101",
  55726=>"101110010",
  55727=>"010001001",
  55728=>"011110111",
  55729=>"101010001",
  55730=>"010111010",
  55731=>"100110011",
  55732=>"000110001",
  55733=>"110101110",
  55734=>"110110001",
  55735=>"010001110",
  55736=>"001101010",
  55737=>"001011111",
  55738=>"110100010",
  55739=>"110010010",
  55740=>"010011000",
  55741=>"010111010",
  55742=>"110111111",
  55743=>"000111011",
  55744=>"111001001",
  55745=>"000011101",
  55746=>"100101110",
  55747=>"011101101",
  55748=>"111110001",
  55749=>"010110000",
  55750=>"100010000",
  55751=>"101111110",
  55752=>"110110001",
  55753=>"100100011",
  55754=>"010110001",
  55755=>"010010011",
  55756=>"111101100",
  55757=>"001100111",
  55758=>"110110010",
  55759=>"001010100",
  55760=>"000001000",
  55761=>"000000100",
  55762=>"001010101",
  55763=>"010001101",
  55764=>"110101110",
  55765=>"000001001",
  55766=>"000001111",
  55767=>"000001110",
  55768=>"001111000",
  55769=>"011001001",
  55770=>"001010000",
  55771=>"000111011",
  55772=>"110011110",
  55773=>"101100000",
  55774=>"111101001",
  55775=>"110011011",
  55776=>"000001101",
  55777=>"100111011",
  55778=>"000101011",
  55779=>"110001000",
  55780=>"100101001",
  55781=>"000110111",
  55782=>"011001111",
  55783=>"100100000",
  55784=>"101000001",
  55785=>"111011000",
  55786=>"110110101",
  55787=>"011100011",
  55788=>"000011100",
  55789=>"000100101",
  55790=>"010001100",
  55791=>"000110100",
  55792=>"001010100",
  55793=>"101010111",
  55794=>"011000001",
  55795=>"001111100",
  55796=>"111010101",
  55797=>"111101001",
  55798=>"011010011",
  55799=>"101111100",
  55800=>"110110100",
  55801=>"000100101",
  55802=>"100001001",
  55803=>"001110101",
  55804=>"010010111",
  55805=>"100100011",
  55806=>"101111001",
  55807=>"100100101",
  55808=>"011110000",
  55809=>"000101110",
  55810=>"000010101",
  55811=>"101001010",
  55812=>"001101111",
  55813=>"000111100",
  55814=>"011101010",
  55815=>"000010010",
  55816=>"010001011",
  55817=>"001011000",
  55818=>"011011001",
  55819=>"001111111",
  55820=>"101000011",
  55821=>"100100100",
  55822=>"100001011",
  55823=>"111110011",
  55824=>"110111111",
  55825=>"111101011",
  55826=>"010110000",
  55827=>"010100010",
  55828=>"111001000",
  55829=>"111011110",
  55830=>"010100001",
  55831=>"001000001",
  55832=>"000010101",
  55833=>"100111111",
  55834=>"011010100",
  55835=>"111110011",
  55836=>"010000010",
  55837=>"011010100",
  55838=>"011000101",
  55839=>"100110110",
  55840=>"011011011",
  55841=>"111100001",
  55842=>"101011010",
  55843=>"000110000",
  55844=>"000110110",
  55845=>"010001000",
  55846=>"010001111",
  55847=>"001110011",
  55848=>"001111011",
  55849=>"110010000",
  55850=>"011110110",
  55851=>"111111000",
  55852=>"101101100",
  55853=>"110010011",
  55854=>"111100001",
  55855=>"010111000",
  55856=>"100101001",
  55857=>"110111111",
  55858=>"011111000",
  55859=>"111011111",
  55860=>"001110000",
  55861=>"101001000",
  55862=>"111010000",
  55863=>"011100111",
  55864=>"011010000",
  55865=>"001101101",
  55866=>"111111111",
  55867=>"111111000",
  55868=>"110011011",
  55869=>"000110110",
  55870=>"001001110",
  55871=>"010011111",
  55872=>"110111111",
  55873=>"000000010",
  55874=>"100110001",
  55875=>"111111000",
  55876=>"101011011",
  55877=>"100001011",
  55878=>"011011010",
  55879=>"111011110",
  55880=>"111001011",
  55881=>"101011001",
  55882=>"000101000",
  55883=>"101111110",
  55884=>"110110110",
  55885=>"101101001",
  55886=>"000100111",
  55887=>"001001011",
  55888=>"001011100",
  55889=>"000111111",
  55890=>"101111100",
  55891=>"011010111",
  55892=>"111010001",
  55893=>"111000101",
  55894=>"111110100",
  55895=>"010111110",
  55896=>"100110000",
  55897=>"011010110",
  55898=>"001000001",
  55899=>"111111000",
  55900=>"111100000",
  55901=>"000001110",
  55902=>"100100011",
  55903=>"000010011",
  55904=>"111001011",
  55905=>"011011101",
  55906=>"111110000",
  55907=>"010001110",
  55908=>"110011100",
  55909=>"111110000",
  55910=>"111000000",
  55911=>"001011101",
  55912=>"101010110",
  55913=>"001011001",
  55914=>"010110110",
  55915=>"000100000",
  55916=>"111011001",
  55917=>"100111100",
  55918=>"100100001",
  55919=>"001101101",
  55920=>"111100110",
  55921=>"011111110",
  55922=>"010101101",
  55923=>"000111110",
  55924=>"000011101",
  55925=>"100101100",
  55926=>"011001011",
  55927=>"001010011",
  55928=>"110011001",
  55929=>"010111011",
  55930=>"001101100",
  55931=>"100101100",
  55932=>"000000001",
  55933=>"011001111",
  55934=>"000000110",
  55935=>"111100111",
  55936=>"110010010",
  55937=>"110111101",
  55938=>"011111011",
  55939=>"011000110",
  55940=>"011110000",
  55941=>"110010111",
  55942=>"010110000",
  55943=>"100000101",
  55944=>"100110001",
  55945=>"110111111",
  55946=>"011010010",
  55947=>"111001110",
  55948=>"000110000",
  55949=>"111111110",
  55950=>"101011101",
  55951=>"001101101",
  55952=>"101000111",
  55953=>"011101101",
  55954=>"111101000",
  55955=>"110000101",
  55956=>"001011100",
  55957=>"000000011",
  55958=>"011001000",
  55959=>"101011111",
  55960=>"101110000",
  55961=>"100000001",
  55962=>"010001110",
  55963=>"100101011",
  55964=>"001100011",
  55965=>"001000001",
  55966=>"000101011",
  55967=>"011100110",
  55968=>"010000000",
  55969=>"111001100",
  55970=>"110111110",
  55971=>"010111110",
  55972=>"111101111",
  55973=>"110101100",
  55974=>"111110100",
  55975=>"111011100",
  55976=>"000011000",
  55977=>"100000011",
  55978=>"110110101",
  55979=>"110000001",
  55980=>"000101111",
  55981=>"001001010",
  55982=>"011110110",
  55983=>"001011000",
  55984=>"000100000",
  55985=>"000111010",
  55986=>"010110011",
  55987=>"001010110",
  55988=>"110001011",
  55989=>"010101111",
  55990=>"001000001",
  55991=>"010010110",
  55992=>"101011001",
  55993=>"001111111",
  55994=>"110010000",
  55995=>"110101110",
  55996=>"000000101",
  55997=>"001110001",
  55998=>"001001110",
  55999=>"001001010",
  56000=>"000100000",
  56001=>"000001011",
  56002=>"100111010",
  56003=>"001000111",
  56004=>"011001100",
  56005=>"101000000",
  56006=>"110010010",
  56007=>"001011100",
  56008=>"010101110",
  56009=>"010011010",
  56010=>"000011111",
  56011=>"001101010",
  56012=>"100011011",
  56013=>"101001010",
  56014=>"101110011",
  56015=>"100001010",
  56016=>"011110110",
  56017=>"010010110",
  56018=>"000011110",
  56019=>"011110111",
  56020=>"111110101",
  56021=>"001001111",
  56022=>"001111011",
  56023=>"001011111",
  56024=>"110110000",
  56025=>"011100011",
  56026=>"101011011",
  56027=>"000110011",
  56028=>"000000000",
  56029=>"111001000",
  56030=>"101001101",
  56031=>"000101011",
  56032=>"001001111",
  56033=>"001010000",
  56034=>"011010111",
  56035=>"000011111",
  56036=>"000111100",
  56037=>"100010010",
  56038=>"000000001",
  56039=>"001011111",
  56040=>"001001001",
  56041=>"010110101",
  56042=>"111110010",
  56043=>"011111011",
  56044=>"011100110",
  56045=>"110110100",
  56046=>"110011000",
  56047=>"111111100",
  56048=>"100001110",
  56049=>"101001010",
  56050=>"101000100",
  56051=>"101010000",
  56052=>"010111011",
  56053=>"000101000",
  56054=>"101111111",
  56055=>"101111000",
  56056=>"110010100",
  56057=>"101111010",
  56058=>"000101000",
  56059=>"000011100",
  56060=>"000110000",
  56061=>"110011111",
  56062=>"000110100",
  56063=>"010100110",
  56064=>"000100000",
  56065=>"100110111",
  56066=>"000011100",
  56067=>"000010110",
  56068=>"011110111",
  56069=>"000001010",
  56070=>"001000011",
  56071=>"001111010",
  56072=>"101100011",
  56073=>"101000011",
  56074=>"000011111",
  56075=>"100011000",
  56076=>"001000101",
  56077=>"100011100",
  56078=>"100010111",
  56079=>"111000000",
  56080=>"001110001",
  56081=>"110010011",
  56082=>"000100100",
  56083=>"100011100",
  56084=>"101111100",
  56085=>"101101000",
  56086=>"010010110",
  56087=>"000000000",
  56088=>"000010011",
  56089=>"010010111",
  56090=>"111010001",
  56091=>"110010000",
  56092=>"100100101",
  56093=>"110110111",
  56094=>"100111011",
  56095=>"000010111",
  56096=>"100100011",
  56097=>"001101011",
  56098=>"011001001",
  56099=>"100010111",
  56100=>"110110010",
  56101=>"010000100",
  56102=>"000111011",
  56103=>"101011000",
  56104=>"001111011",
  56105=>"001111011",
  56106=>"110010010",
  56107=>"100111111",
  56108=>"111000010",
  56109=>"011001100",
  56110=>"010010111",
  56111=>"001010101",
  56112=>"000001010",
  56113=>"011111110",
  56114=>"101000100",
  56115=>"001010000",
  56116=>"010011001",
  56117=>"110101000",
  56118=>"011111000",
  56119=>"010101000",
  56120=>"011110000",
  56121=>"010101111",
  56122=>"100111011",
  56123=>"100000101",
  56124=>"010000010",
  56125=>"000011010",
  56126=>"010000101",
  56127=>"100110000",
  56128=>"011101001",
  56129=>"111001000",
  56130=>"101001110",
  56131=>"100100100",
  56132=>"111101001",
  56133=>"111010100",
  56134=>"110110111",
  56135=>"101010111",
  56136=>"010110111",
  56137=>"101011011",
  56138=>"000110110",
  56139=>"111100000",
  56140=>"101010010",
  56141=>"110100111",
  56142=>"001111010",
  56143=>"100110000",
  56144=>"111111111",
  56145=>"011011011",
  56146=>"100110001",
  56147=>"011010010",
  56148=>"000010110",
  56149=>"010110000",
  56150=>"010110100",
  56151=>"000110111",
  56152=>"001110110",
  56153=>"011010110",
  56154=>"100111100",
  56155=>"100110000",
  56156=>"011111001",
  56157=>"010001000",
  56158=>"001110111",
  56159=>"001010011",
  56160=>"011110101",
  56161=>"000011011",
  56162=>"000100010",
  56163=>"010111010",
  56164=>"000000000",
  56165=>"101011000",
  56166=>"111010011",
  56167=>"000111000",
  56168=>"000001000",
  56169=>"111111001",
  56170=>"010110100",
  56171=>"000001011",
  56172=>"101010001",
  56173=>"100001111",
  56174=>"010001100",
  56175=>"100100001",
  56176=>"011011010",
  56177=>"001001110",
  56178=>"101111001",
  56179=>"110111000",
  56180=>"111110101",
  56181=>"010100010",
  56182=>"101100100",
  56183=>"000001010",
  56184=>"011100100",
  56185=>"001001011",
  56186=>"110101010",
  56187=>"100011100",
  56188=>"000101000",
  56189=>"010001101",
  56190=>"100101111",
  56191=>"000011110",
  56192=>"101101110",
  56193=>"101111100",
  56194=>"111000111",
  56195=>"110100111",
  56196=>"000100010",
  56197=>"001000011",
  56198=>"000101011",
  56199=>"101000100",
  56200=>"001010110",
  56201=>"011100110",
  56202=>"111101010",
  56203=>"000001010",
  56204=>"011011101",
  56205=>"111100000",
  56206=>"111110111",
  56207=>"010011000",
  56208=>"011100101",
  56209=>"010100110",
  56210=>"100001101",
  56211=>"001111110",
  56212=>"001110000",
  56213=>"011000110",
  56214=>"001010001",
  56215=>"001011100",
  56216=>"101000010",
  56217=>"001110111",
  56218=>"110101000",
  56219=>"001100100",
  56220=>"011010110",
  56221=>"001101011",
  56222=>"100100000",
  56223=>"111100100",
  56224=>"000000000",
  56225=>"100110111",
  56226=>"000111110",
  56227=>"100000011",
  56228=>"111010000",
  56229=>"010010010",
  56230=>"001010000",
  56231=>"010100101",
  56232=>"010011111",
  56233=>"100100000",
  56234=>"000101011",
  56235=>"010011101",
  56236=>"001001011",
  56237=>"000010010",
  56238=>"010000001",
  56239=>"000111111",
  56240=>"011000101",
  56241=>"111001101",
  56242=>"100111110",
  56243=>"001101101",
  56244=>"110110000",
  56245=>"111100001",
  56246=>"110100111",
  56247=>"001001111",
  56248=>"110010001",
  56249=>"001101011",
  56250=>"011100100",
  56251=>"011111000",
  56252=>"000010110",
  56253=>"010000100",
  56254=>"000000000",
  56255=>"011100100",
  56256=>"001111000",
  56257=>"100001100",
  56258=>"011010000",
  56259=>"001100001",
  56260=>"010000101",
  56261=>"000101011",
  56262=>"110000110",
  56263=>"101100100",
  56264=>"001101100",
  56265=>"000010010",
  56266=>"010110001",
  56267=>"101101100",
  56268=>"010111111",
  56269=>"111010100",
  56270=>"011111010",
  56271=>"001011110",
  56272=>"011010100",
  56273=>"111011111",
  56274=>"011101011",
  56275=>"110000101",
  56276=>"011110011",
  56277=>"100101010",
  56278=>"111111111",
  56279=>"111000011",
  56280=>"111011000",
  56281=>"001001010",
  56282=>"110111000",
  56283=>"101111000",
  56284=>"001110010",
  56285=>"000000011",
  56286=>"001011011",
  56287=>"110010001",
  56288=>"111000100",
  56289=>"110000100",
  56290=>"101100100",
  56291=>"000000000",
  56292=>"010111001",
  56293=>"100111110",
  56294=>"000111111",
  56295=>"000000111",
  56296=>"001101000",
  56297=>"100001001",
  56298=>"001101010",
  56299=>"000110111",
  56300=>"010010011",
  56301=>"000010111",
  56302=>"110111100",
  56303=>"100110111",
  56304=>"101110111",
  56305=>"011100011",
  56306=>"111101110",
  56307=>"001001010",
  56308=>"011010110",
  56309=>"010011111",
  56310=>"000011011",
  56311=>"111111110",
  56312=>"101011011",
  56313=>"000011111",
  56314=>"010000101",
  56315=>"000011000",
  56316=>"110001111",
  56317=>"011100001",
  56318=>"110010100",
  56319=>"001111111",
  56320=>"000000100",
  56321=>"011001111",
  56322=>"101010110",
  56323=>"111010111",
  56324=>"111010101",
  56325=>"111011110",
  56326=>"000000010",
  56327=>"000001001",
  56328=>"101010000",
  56329=>"001001010",
  56330=>"001111110",
  56331=>"011001101",
  56332=>"010010000",
  56333=>"000010001",
  56334=>"010001100",
  56335=>"100110101",
  56336=>"110000001",
  56337=>"110011011",
  56338=>"000000110",
  56339=>"101100001",
  56340=>"110011010",
  56341=>"001010000",
  56342=>"101110010",
  56343=>"101001010",
  56344=>"111100101",
  56345=>"011001001",
  56346=>"101111110",
  56347=>"101011010",
  56348=>"010111100",
  56349=>"100100100",
  56350=>"010100111",
  56351=>"111100100",
  56352=>"110101101",
  56353=>"010011010",
  56354=>"110111010",
  56355=>"110100001",
  56356=>"111110000",
  56357=>"011000000",
  56358=>"011101101",
  56359=>"101001001",
  56360=>"101100100",
  56361=>"111000011",
  56362=>"101101000",
  56363=>"000110100",
  56364=>"011110101",
  56365=>"000011001",
  56366=>"010000000",
  56367=>"010100010",
  56368=>"110100110",
  56369=>"001011011",
  56370=>"101111001",
  56371=>"101100111",
  56372=>"110101100",
  56373=>"001100110",
  56374=>"011001100",
  56375=>"000001001",
  56376=>"110011111",
  56377=>"001101010",
  56378=>"100010011",
  56379=>"011111011",
  56380=>"110110001",
  56381=>"000000100",
  56382=>"011111110",
  56383=>"010011010",
  56384=>"101011100",
  56385=>"000000000",
  56386=>"101011010",
  56387=>"000111000",
  56388=>"011011110",
  56389=>"110111110",
  56390=>"010111100",
  56391=>"000111111",
  56392=>"011101100",
  56393=>"110110011",
  56394=>"110101100",
  56395=>"110010001",
  56396=>"101110110",
  56397=>"111010000",
  56398=>"100111001",
  56399=>"110001010",
  56400=>"010100011",
  56401=>"011111111",
  56402=>"110001110",
  56403=>"010011000",
  56404=>"111011100",
  56405=>"100010100",
  56406=>"111111101",
  56407=>"111100111",
  56408=>"100011100",
  56409=>"101111110",
  56410=>"000010110",
  56411=>"111101111",
  56412=>"001110011",
  56413=>"010000100",
  56414=>"001010011",
  56415=>"100111111",
  56416=>"110011001",
  56417=>"101101010",
  56418=>"111010100",
  56419=>"110101010",
  56420=>"101111001",
  56421=>"110110101",
  56422=>"110001010",
  56423=>"101001111",
  56424=>"001011110",
  56425=>"110000000",
  56426=>"010100010",
  56427=>"000110100",
  56428=>"110001010",
  56429=>"101111001",
  56430=>"001111001",
  56431=>"001000011",
  56432=>"101111111",
  56433=>"001010101",
  56434=>"001110111",
  56435=>"101011011",
  56436=>"001101000",
  56437=>"000101101",
  56438=>"110101000",
  56439=>"001100111",
  56440=>"100100000",
  56441=>"100000111",
  56442=>"101010000",
  56443=>"011110100",
  56444=>"111000101",
  56445=>"001111100",
  56446=>"101110111",
  56447=>"100001111",
  56448=>"011011111",
  56449=>"111100001",
  56450=>"100001000",
  56451=>"000011111",
  56452=>"110101000",
  56453=>"110101110",
  56454=>"111010011",
  56455=>"011100111",
  56456=>"111101110",
  56457=>"011000110",
  56458=>"001101111",
  56459=>"010110101",
  56460=>"011000001",
  56461=>"101101101",
  56462=>"000010100",
  56463=>"100111001",
  56464=>"000001110",
  56465=>"010001000",
  56466=>"110011010",
  56467=>"011010010",
  56468=>"010000100",
  56469=>"111100010",
  56470=>"111011010",
  56471=>"000110111",
  56472=>"111001010",
  56473=>"111010000",
  56474=>"100001100",
  56475=>"111011011",
  56476=>"100000100",
  56477=>"000001000",
  56478=>"110000111",
  56479=>"011010110",
  56480=>"111011111",
  56481=>"000001100",
  56482=>"100111101",
  56483=>"111110011",
  56484=>"101110110",
  56485=>"000101111",
  56486=>"101110001",
  56487=>"111110101",
  56488=>"100011111",
  56489=>"111001110",
  56490=>"101100110",
  56491=>"110001100",
  56492=>"001010111",
  56493=>"001101101",
  56494=>"111011100",
  56495=>"010100001",
  56496=>"011000110",
  56497=>"101001010",
  56498=>"010010000",
  56499=>"110100001",
  56500=>"011100010",
  56501=>"011011101",
  56502=>"110101001",
  56503=>"111111000",
  56504=>"011001101",
  56505=>"101100101",
  56506=>"101100001",
  56507=>"011001000",
  56508=>"011010110",
  56509=>"001001110",
  56510=>"000101001",
  56511=>"111011110",
  56512=>"010101101",
  56513=>"110011101",
  56514=>"110100100",
  56515=>"110010001",
  56516=>"101100001",
  56517=>"100101011",
  56518=>"101100000",
  56519=>"000000000",
  56520=>"000000010",
  56521=>"000111011",
  56522=>"101110011",
  56523=>"111001000",
  56524=>"111010000",
  56525=>"000010111",
  56526=>"000110100",
  56527=>"111111111",
  56528=>"100000000",
  56529=>"000010010",
  56530=>"111010010",
  56531=>"100000001",
  56532=>"000110111",
  56533=>"101011001",
  56534=>"000101000",
  56535=>"110011010",
  56536=>"101100000",
  56537=>"000101001",
  56538=>"111011000",
  56539=>"001000010",
  56540=>"000001101",
  56541=>"011000001",
  56542=>"011110001",
  56543=>"111111100",
  56544=>"110101100",
  56545=>"000010001",
  56546=>"111010101",
  56547=>"000011101",
  56548=>"010000101",
  56549=>"010100101",
  56550=>"001001010",
  56551=>"001001011",
  56552=>"111110111",
  56553=>"001001010",
  56554=>"000101110",
  56555=>"111000111",
  56556=>"011110101",
  56557=>"111100100",
  56558=>"100111100",
  56559=>"100101010",
  56560=>"100011000",
  56561=>"000100100",
  56562=>"110110011",
  56563=>"101111101",
  56564=>"101110100",
  56565=>"001010111",
  56566=>"011111000",
  56567=>"001000001",
  56568=>"101000110",
  56569=>"011011101",
  56570=>"000100000",
  56571=>"011001010",
  56572=>"110111110",
  56573=>"011010010",
  56574=>"011000001",
  56575=>"011100111",
  56576=>"001100000",
  56577=>"010101001",
  56578=>"010111001",
  56579=>"111011001",
  56580=>"111110111",
  56581=>"010001001",
  56582=>"011001000",
  56583=>"010001111",
  56584=>"110110110",
  56585=>"101101101",
  56586=>"010011111",
  56587=>"001100100",
  56588=>"101111010",
  56589=>"110010101",
  56590=>"111110000",
  56591=>"001001010",
  56592=>"101111101",
  56593=>"111101010",
  56594=>"001111000",
  56595=>"011101111",
  56596=>"000000001",
  56597=>"100011100",
  56598=>"111000110",
  56599=>"111100111",
  56600=>"001000001",
  56601=>"100011111",
  56602=>"111010111",
  56603=>"000110000",
  56604=>"001001001",
  56605=>"101001101",
  56606=>"000111001",
  56607=>"111000100",
  56608=>"000001010",
  56609=>"110010011",
  56610=>"100111110",
  56611=>"111100111",
  56612=>"110110010",
  56613=>"101111111",
  56614=>"101110011",
  56615=>"010100001",
  56616=>"001000010",
  56617=>"110010110",
  56618=>"100110101",
  56619=>"011000111",
  56620=>"001111110",
  56621=>"000100011",
  56622=>"110011011",
  56623=>"110000011",
  56624=>"110101011",
  56625=>"001010001",
  56626=>"111100011",
  56627=>"110000000",
  56628=>"100111001",
  56629=>"001000110",
  56630=>"000110001",
  56631=>"000001011",
  56632=>"100011101",
  56633=>"011110101",
  56634=>"101100110",
  56635=>"000110110",
  56636=>"010010001",
  56637=>"001101110",
  56638=>"101111011",
  56639=>"001000110",
  56640=>"010001011",
  56641=>"110001101",
  56642=>"100011000",
  56643=>"001101011",
  56644=>"110010110",
  56645=>"111110010",
  56646=>"110101011",
  56647=>"111010110",
  56648=>"011111110",
  56649=>"110000010",
  56650=>"000000111",
  56651=>"111111110",
  56652=>"101100101",
  56653=>"010111010",
  56654=>"010111001",
  56655=>"101011001",
  56656=>"001101011",
  56657=>"110001010",
  56658=>"011011010",
  56659=>"010100111",
  56660=>"010111001",
  56661=>"000000101",
  56662=>"010100110",
  56663=>"110101001",
  56664=>"101010111",
  56665=>"010100000",
  56666=>"110100100",
  56667=>"111101111",
  56668=>"110110110",
  56669=>"011100000",
  56670=>"011110011",
  56671=>"110000101",
  56672=>"001010101",
  56673=>"001011101",
  56674=>"001001000",
  56675=>"111010111",
  56676=>"010110100",
  56677=>"100000011",
  56678=>"000101110",
  56679=>"100001001",
  56680=>"101011100",
  56681=>"100000100",
  56682=>"011100110",
  56683=>"111001101",
  56684=>"111110000",
  56685=>"010101010",
  56686=>"000110001",
  56687=>"010010011",
  56688=>"011010101",
  56689=>"110011011",
  56690=>"001111010",
  56691=>"000001010",
  56692=>"111100010",
  56693=>"001100101",
  56694=>"111101100",
  56695=>"101001111",
  56696=>"010010011",
  56697=>"000111011",
  56698=>"011000111",
  56699=>"100000000",
  56700=>"111110100",
  56701=>"110001110",
  56702=>"011111000",
  56703=>"011010001",
  56704=>"010100100",
  56705=>"001111111",
  56706=>"001010011",
  56707=>"000001100",
  56708=>"110001000",
  56709=>"011000111",
  56710=>"001011000",
  56711=>"111010101",
  56712=>"111110011",
  56713=>"111101011",
  56714=>"000010100",
  56715=>"100001001",
  56716=>"001011100",
  56717=>"111110001",
  56718=>"011110001",
  56719=>"100100111",
  56720=>"000101111",
  56721=>"111000110",
  56722=>"110011110",
  56723=>"001010000",
  56724=>"101111111",
  56725=>"000000000",
  56726=>"110101001",
  56727=>"110001101",
  56728=>"110011101",
  56729=>"000101000",
  56730=>"111110111",
  56731=>"011100110",
  56732=>"111000010",
  56733=>"001011100",
  56734=>"011010111",
  56735=>"000110000",
  56736=>"000110000",
  56737=>"101110110",
  56738=>"011110010",
  56739=>"000001100",
  56740=>"111001101",
  56741=>"000001101",
  56742=>"110110101",
  56743=>"111110011",
  56744=>"011101110",
  56745=>"000101010",
  56746=>"011000100",
  56747=>"111000011",
  56748=>"100110011",
  56749=>"110110010",
  56750=>"100001110",
  56751=>"001110011",
  56752=>"111000100",
  56753=>"110111110",
  56754=>"111111011",
  56755=>"010100110",
  56756=>"001101111",
  56757=>"111001110",
  56758=>"100001100",
  56759=>"101000000",
  56760=>"010111110",
  56761=>"001101110",
  56762=>"000010011",
  56763=>"001101111",
  56764=>"101110111",
  56765=>"011101011",
  56766=>"111001011",
  56767=>"011000100",
  56768=>"011100010",
  56769=>"001101001",
  56770=>"001110011",
  56771=>"101101001",
  56772=>"100110110",
  56773=>"001001100",
  56774=>"010011000",
  56775=>"111101111",
  56776=>"010010001",
  56777=>"101001110",
  56778=>"010001100",
  56779=>"100001001",
  56780=>"111001010",
  56781=>"101010000",
  56782=>"010100110",
  56783=>"001010111",
  56784=>"101110100",
  56785=>"010010011",
  56786=>"100011010",
  56787=>"000100010",
  56788=>"111110110",
  56789=>"101001001",
  56790=>"110000010",
  56791=>"000111000",
  56792=>"000000010",
  56793=>"011100011",
  56794=>"101100110",
  56795=>"000111101",
  56796=>"001000001",
  56797=>"111001010",
  56798=>"101110011",
  56799=>"100101010",
  56800=>"001110100",
  56801=>"111101111",
  56802=>"110111010",
  56803=>"010000101",
  56804=>"000111010",
  56805=>"111111100",
  56806=>"001101111",
  56807=>"111111110",
  56808=>"110110101",
  56809=>"000100010",
  56810=>"101010000",
  56811=>"010100001",
  56812=>"010000010",
  56813=>"000001010",
  56814=>"110011011",
  56815=>"101011010",
  56816=>"011100000",
  56817=>"111000010",
  56818=>"000110110",
  56819=>"101111100",
  56820=>"100100101",
  56821=>"010010110",
  56822=>"010000001",
  56823=>"010000001",
  56824=>"000001111",
  56825=>"010111000",
  56826=>"110110111",
  56827=>"100010101",
  56828=>"010100000",
  56829=>"010110100",
  56830=>"101011001",
  56831=>"011101111",
  56832=>"000101010",
  56833=>"111110100",
  56834=>"000000000",
  56835=>"010110011",
  56836=>"011100000",
  56837=>"101011101",
  56838=>"001000000",
  56839=>"111111000",
  56840=>"100010100",
  56841=>"100000011",
  56842=>"000111100",
  56843=>"000001011",
  56844=>"110100011",
  56845=>"100001100",
  56846=>"111100110",
  56847=>"111011000",
  56848=>"101011101",
  56849=>"001110000",
  56850=>"000011000",
  56851=>"100111100",
  56852=>"101001100",
  56853=>"011110110",
  56854=>"110010010",
  56855=>"001001000",
  56856=>"000100111",
  56857=>"101101100",
  56858=>"011110001",
  56859=>"111000111",
  56860=>"100010000",
  56861=>"101111110",
  56862=>"001100101",
  56863=>"010100110",
  56864=>"010101001",
  56865=>"101110100",
  56866=>"010100100",
  56867=>"000011000",
  56868=>"111110111",
  56869=>"000100110",
  56870=>"011000001",
  56871=>"010100111",
  56872=>"100111111",
  56873=>"111111101",
  56874=>"010001001",
  56875=>"111010100",
  56876=>"000011110",
  56877=>"101010011",
  56878=>"100010000",
  56879=>"111010001",
  56880=>"001011110",
  56881=>"011111001",
  56882=>"111110110",
  56883=>"101111011",
  56884=>"011111110",
  56885=>"100011010",
  56886=>"100001101",
  56887=>"101100101",
  56888=>"111111101",
  56889=>"100001001",
  56890=>"000011110",
  56891=>"100111001",
  56892=>"001100100",
  56893=>"010011010",
  56894=>"100101111",
  56895=>"100000000",
  56896=>"011000101",
  56897=>"000001110",
  56898=>"100000011",
  56899=>"111011101",
  56900=>"001010110",
  56901=>"111100010",
  56902=>"010011111",
  56903=>"010100101",
  56904=>"110101000",
  56905=>"101011111",
  56906=>"110000101",
  56907=>"111010000",
  56908=>"011111001",
  56909=>"011111001",
  56910=>"110001110",
  56911=>"001001110",
  56912=>"100110000",
  56913=>"010010010",
  56914=>"010010000",
  56915=>"010111000",
  56916=>"111111010",
  56917=>"000100111",
  56918=>"110100111",
  56919=>"001111101",
  56920=>"100011001",
  56921=>"111010001",
  56922=>"100010010",
  56923=>"111000101",
  56924=>"011001011",
  56925=>"011101001",
  56926=>"111100011",
  56927=>"011001111",
  56928=>"010100001",
  56929=>"110001110",
  56930=>"001110111",
  56931=>"000011101",
  56932=>"001110110",
  56933=>"110110010",
  56934=>"111001010",
  56935=>"011110101",
  56936=>"010001000",
  56937=>"100001001",
  56938=>"111110111",
  56939=>"111011100",
  56940=>"010101010",
  56941=>"111101111",
  56942=>"111010000",
  56943=>"110011110",
  56944=>"110111010",
  56945=>"110001110",
  56946=>"011010110",
  56947=>"110011011",
  56948=>"000000011",
  56949=>"011010100",
  56950=>"010001000",
  56951=>"110000010",
  56952=>"101011110",
  56953=>"001000111",
  56954=>"000000100",
  56955=>"010000001",
  56956=>"001000011",
  56957=>"001000010",
  56958=>"010111100",
  56959=>"010011101",
  56960=>"100011010",
  56961=>"010001100",
  56962=>"110010100",
  56963=>"110011100",
  56964=>"101011010",
  56965=>"111000110",
  56966=>"011000011",
  56967=>"010001000",
  56968=>"010101000",
  56969=>"001101010",
  56970=>"011011000",
  56971=>"100010001",
  56972=>"010010100",
  56973=>"110100100",
  56974=>"010011011",
  56975=>"001001000",
  56976=>"001011011",
  56977=>"000010111",
  56978=>"011101111",
  56979=>"011101101",
  56980=>"000110010",
  56981=>"001111110",
  56982=>"011000110",
  56983=>"100100100",
  56984=>"100001000",
  56985=>"010101101",
  56986=>"001101011",
  56987=>"010101011",
  56988=>"000111000",
  56989=>"010110100",
  56990=>"000010010",
  56991=>"100100001",
  56992=>"000001001",
  56993=>"010011001",
  56994=>"110010011",
  56995=>"111111111",
  56996=>"101101111",
  56997=>"011010010",
  56998=>"111001110",
  56999=>"000000010",
  57000=>"110100001",
  57001=>"101010100",
  57002=>"010101000",
  57003=>"000111001",
  57004=>"101000000",
  57005=>"100011000",
  57006=>"110100110",
  57007=>"101110111",
  57008=>"111001010",
  57009=>"001011001",
  57010=>"101011001",
  57011=>"010101000",
  57012=>"010110101",
  57013=>"010110001",
  57014=>"001110111",
  57015=>"101101011",
  57016=>"111110100",
  57017=>"110111110",
  57018=>"100110111",
  57019=>"000111101",
  57020=>"010011101",
  57021=>"011111101",
  57022=>"111011110",
  57023=>"000000001",
  57024=>"001000110",
  57025=>"110100010",
  57026=>"101010110",
  57027=>"101001010",
  57028=>"100001000",
  57029=>"001101111",
  57030=>"110001010",
  57031=>"001000000",
  57032=>"011111000",
  57033=>"011110010",
  57034=>"110110100",
  57035=>"111010001",
  57036=>"111110110",
  57037=>"101010010",
  57038=>"100100011",
  57039=>"100011011",
  57040=>"111111110",
  57041=>"000010000",
  57042=>"000110000",
  57043=>"110101000",
  57044=>"010100110",
  57045=>"111011111",
  57046=>"011011110",
  57047=>"100000111",
  57048=>"000000111",
  57049=>"001011101",
  57050=>"101111001",
  57051=>"110100000",
  57052=>"010001100",
  57053=>"100010101",
  57054=>"001011011",
  57055=>"110001100",
  57056=>"000000000",
  57057=>"001110110",
  57058=>"000000010",
  57059=>"111000110",
  57060=>"111111001",
  57061=>"100000010",
  57062=>"000111000",
  57063=>"000110000",
  57064=>"001110100",
  57065=>"111100011",
  57066=>"000010001",
  57067=>"100000100",
  57068=>"010001001",
  57069=>"111000011",
  57070=>"100110111",
  57071=>"111010001",
  57072=>"001010001",
  57073=>"000000010",
  57074=>"110001001",
  57075=>"101010010",
  57076=>"000111010",
  57077=>"111100011",
  57078=>"000100111",
  57079=>"011001100",
  57080=>"100110011",
  57081=>"111000010",
  57082=>"111001101",
  57083=>"101000101",
  57084=>"001111111",
  57085=>"101011111",
  57086=>"110010001",
  57087=>"001001001",
  57088=>"111111110",
  57089=>"010000010",
  57090=>"010010100",
  57091=>"100000110",
  57092=>"110001100",
  57093=>"011001001",
  57094=>"011101010",
  57095=>"110101010",
  57096=>"110010000",
  57097=>"100011010",
  57098=>"001010011",
  57099=>"010010001",
  57100=>"100110100",
  57101=>"100100100",
  57102=>"010111001",
  57103=>"111101111",
  57104=>"111001100",
  57105=>"110110110",
  57106=>"100111001",
  57107=>"011010101",
  57108=>"111100000",
  57109=>"011111100",
  57110=>"011001001",
  57111=>"111110011",
  57112=>"111000110",
  57113=>"110000010",
  57114=>"001100111",
  57115=>"000110110",
  57116=>"010110101",
  57117=>"111011111",
  57118=>"111111010",
  57119=>"010100110",
  57120=>"000101001",
  57121=>"011000101",
  57122=>"101011100",
  57123=>"101000000",
  57124=>"011010111",
  57125=>"110000110",
  57126=>"100100101",
  57127=>"011110000",
  57128=>"010000010",
  57129=>"110001001",
  57130=>"100001011",
  57131=>"101110111",
  57132=>"100000101",
  57133=>"001000000",
  57134=>"100100011",
  57135=>"100010101",
  57136=>"110001001",
  57137=>"110110100",
  57138=>"001101110",
  57139=>"100001001",
  57140=>"000010111",
  57141=>"101100100",
  57142=>"011011000",
  57143=>"001111110",
  57144=>"001011010",
  57145=>"001100000",
  57146=>"110001000",
  57147=>"101110011",
  57148=>"010100010",
  57149=>"001000101",
  57150=>"100111010",
  57151=>"010001111",
  57152=>"111001001",
  57153=>"101111111",
  57154=>"100110110",
  57155=>"111111111",
  57156=>"001011101",
  57157=>"000100011",
  57158=>"011010001",
  57159=>"111001000",
  57160=>"011100100",
  57161=>"100000011",
  57162=>"010001110",
  57163=>"011011111",
  57164=>"000010001",
  57165=>"001010001",
  57166=>"011000100",
  57167=>"001000011",
  57168=>"110000000",
  57169=>"111011001",
  57170=>"010100101",
  57171=>"110100110",
  57172=>"111001110",
  57173=>"010100000",
  57174=>"111011101",
  57175=>"101001001",
  57176=>"101000101",
  57177=>"111101001",
  57178=>"100111101",
  57179=>"000000111",
  57180=>"110010111",
  57181=>"101001001",
  57182=>"010111000",
  57183=>"111000101",
  57184=>"101110101",
  57185=>"111011011",
  57186=>"111101111",
  57187=>"001101111",
  57188=>"111101010",
  57189=>"011011010",
  57190=>"111110010",
  57191=>"001001110",
  57192=>"001001010",
  57193=>"101000011",
  57194=>"010101001",
  57195=>"001100010",
  57196=>"000001001",
  57197=>"100100010",
  57198=>"101111101",
  57199=>"111111001",
  57200=>"101010010",
  57201=>"010111010",
  57202=>"100110110",
  57203=>"011011011",
  57204=>"000010100",
  57205=>"000111110",
  57206=>"000000111",
  57207=>"010011100",
  57208=>"100101110",
  57209=>"011010001",
  57210=>"110000110",
  57211=>"000001010",
  57212=>"001011010",
  57213=>"001010001",
  57214=>"001111001",
  57215=>"101110111",
  57216=>"011100000",
  57217=>"111101010",
  57218=>"011110111",
  57219=>"100101101",
  57220=>"101000011",
  57221=>"010100001",
  57222=>"110011001",
  57223=>"000100100",
  57224=>"010100010",
  57225=>"100010001",
  57226=>"111111111",
  57227=>"110010010",
  57228=>"100110100",
  57229=>"100111001",
  57230=>"110111010",
  57231=>"000010101",
  57232=>"110010000",
  57233=>"010110101",
  57234=>"111110001",
  57235=>"111011000",
  57236=>"011010111",
  57237=>"010001101",
  57238=>"000110100",
  57239=>"000111001",
  57240=>"101100001",
  57241=>"101000100",
  57242=>"010110010",
  57243=>"111111010",
  57244=>"010000001",
  57245=>"010001101",
  57246=>"000000010",
  57247=>"101011101",
  57248=>"000111000",
  57249=>"110000101",
  57250=>"011001001",
  57251=>"101000001",
  57252=>"000010100",
  57253=>"101011011",
  57254=>"011101111",
  57255=>"111011101",
  57256=>"101110101",
  57257=>"000000101",
  57258=>"011100010",
  57259=>"011101101",
  57260=>"101100000",
  57261=>"001000101",
  57262=>"011010011",
  57263=>"101111000",
  57264=>"100010111",
  57265=>"000111001",
  57266=>"101001011",
  57267=>"000011111",
  57268=>"010001001",
  57269=>"111011001",
  57270=>"001111011",
  57271=>"111010111",
  57272=>"010000111",
  57273=>"111000001",
  57274=>"000101011",
  57275=>"100101100",
  57276=>"100010000",
  57277=>"010111000",
  57278=>"111000010",
  57279=>"000111001",
  57280=>"000001000",
  57281=>"101101100",
  57282=>"111100000",
  57283=>"101111000",
  57284=>"000100000",
  57285=>"111111100",
  57286=>"010011110",
  57287=>"100101101",
  57288=>"000100101",
  57289=>"100101110",
  57290=>"000001110",
  57291=>"011001010",
  57292=>"010101011",
  57293=>"000111000",
  57294=>"101010011",
  57295=>"000100000",
  57296=>"111100010",
  57297=>"000011010",
  57298=>"000010001",
  57299=>"010101101",
  57300=>"001011111",
  57301=>"011111011",
  57302=>"111111100",
  57303=>"000001111",
  57304=>"000111010",
  57305=>"101111100",
  57306=>"010011101",
  57307=>"111110011",
  57308=>"110111100",
  57309=>"010010000",
  57310=>"110110001",
  57311=>"000000101",
  57312=>"011111001",
  57313=>"101101110",
  57314=>"001001011",
  57315=>"110001011",
  57316=>"100011101",
  57317=>"000111010",
  57318=>"111100011",
  57319=>"100100000",
  57320=>"010101010",
  57321=>"011011010",
  57322=>"110110001",
  57323=>"010110010",
  57324=>"101101101",
  57325=>"001010010",
  57326=>"100000100",
  57327=>"101000100",
  57328=>"101010000",
  57329=>"101001110",
  57330=>"110011111",
  57331=>"011000010",
  57332=>"010011010",
  57333=>"101000000",
  57334=>"101100110",
  57335=>"000000110",
  57336=>"011010001",
  57337=>"100111010",
  57338=>"000000001",
  57339=>"100111111",
  57340=>"011001001",
  57341=>"000100001",
  57342=>"000100011",
  57343=>"000111010",
  57344=>"010101001",
  57345=>"100001000",
  57346=>"011110101",
  57347=>"110110010",
  57348=>"110100001",
  57349=>"100111110",
  57350=>"001100110",
  57351=>"100000001",
  57352=>"101010010",
  57353=>"101001101",
  57354=>"111010010",
  57355=>"100010010",
  57356=>"001100011",
  57357=>"110100101",
  57358=>"110000011",
  57359=>"001100111",
  57360=>"110111001",
  57361=>"001110011",
  57362=>"000011001",
  57363=>"001000011",
  57364=>"101101111",
  57365=>"010101001",
  57366=>"110100010",
  57367=>"011010100",
  57368=>"000100001",
  57369=>"000001000",
  57370=>"101100111",
  57371=>"011110001",
  57372=>"011100101",
  57373=>"100011100",
  57374=>"101101010",
  57375=>"111000000",
  57376=>"000011110",
  57377=>"111111111",
  57378=>"111111011",
  57379=>"101010110",
  57380=>"010001010",
  57381=>"111101010",
  57382=>"000100101",
  57383=>"001010000",
  57384=>"100110100",
  57385=>"111111110",
  57386=>"011010111",
  57387=>"010011010",
  57388=>"000010010",
  57389=>"110100101",
  57390=>"101001100",
  57391=>"000001111",
  57392=>"000010100",
  57393=>"100100101",
  57394=>"001101110",
  57395=>"001101010",
  57396=>"000010100",
  57397=>"110010011",
  57398=>"000011110",
  57399=>"010001100",
  57400=>"110110000",
  57401=>"111000001",
  57402=>"101110100",
  57403=>"111110000",
  57404=>"000010000",
  57405=>"001000110",
  57406=>"111101000",
  57407=>"000011111",
  57408=>"001001010",
  57409=>"010011110",
  57410=>"010101010",
  57411=>"000101111",
  57412=>"011110010",
  57413=>"011001110",
  57414=>"001101000",
  57415=>"000011101",
  57416=>"000000110",
  57417=>"000010110",
  57418=>"110001111",
  57419=>"000110111",
  57420=>"000001011",
  57421=>"110101001",
  57422=>"010011001",
  57423=>"100101110",
  57424=>"111100100",
  57425=>"000010000",
  57426=>"010101001",
  57427=>"100110001",
  57428=>"101010100",
  57429=>"011010011",
  57430=>"101101001",
  57431=>"110000000",
  57432=>"000111001",
  57433=>"111101101",
  57434=>"001101111",
  57435=>"011000011",
  57436=>"001110101",
  57437=>"011010000",
  57438=>"011010011",
  57439=>"000111111",
  57440=>"000001100",
  57441=>"001110001",
  57442=>"101000101",
  57443=>"100000000",
  57444=>"001010010",
  57445=>"010001001",
  57446=>"001110101",
  57447=>"010110101",
  57448=>"000010111",
  57449=>"010000010",
  57450=>"111110111",
  57451=>"000100010",
  57452=>"111001001",
  57453=>"111011101",
  57454=>"100100101",
  57455=>"000000010",
  57456=>"000001011",
  57457=>"101000111",
  57458=>"101000101",
  57459=>"011001001",
  57460=>"000101111",
  57461=>"000100100",
  57462=>"001011111",
  57463=>"000011010",
  57464=>"011111011",
  57465=>"000111111",
  57466=>"000001000",
  57467=>"011110010",
  57468=>"001011110",
  57469=>"101011000",
  57470=>"010000010",
  57471=>"011010101",
  57472=>"110001110",
  57473=>"101111001",
  57474=>"111010110",
  57475=>"010110011",
  57476=>"111110101",
  57477=>"111100100",
  57478=>"100001101",
  57479=>"111100001",
  57480=>"110011111",
  57481=>"010000101",
  57482=>"000111001",
  57483=>"110100100",
  57484=>"001011011",
  57485=>"001010111",
  57486=>"100110000",
  57487=>"111111111",
  57488=>"100000010",
  57489=>"011010110",
  57490=>"010100000",
  57491=>"000000000",
  57492=>"000010011",
  57493=>"101110111",
  57494=>"001000011",
  57495=>"101000010",
  57496=>"000011000",
  57497=>"000100101",
  57498=>"010000001",
  57499=>"101111110",
  57500=>"000100011",
  57501=>"000101111",
  57502=>"000011101",
  57503=>"000011111",
  57504=>"010000000",
  57505=>"110000001",
  57506=>"111101110",
  57507=>"000001000",
  57508=>"111100110",
  57509=>"011110001",
  57510=>"010001101",
  57511=>"100110111",
  57512=>"000101001",
  57513=>"111011001",
  57514=>"011000010",
  57515=>"010101010",
  57516=>"001100100",
  57517=>"010010111",
  57518=>"000110000",
  57519=>"110011111",
  57520=>"000011011",
  57521=>"000010000",
  57522=>"100000101",
  57523=>"100001000",
  57524=>"010101101",
  57525=>"011010101",
  57526=>"111110000",
  57527=>"111100001",
  57528=>"000011110",
  57529=>"101001101",
  57530=>"000101111",
  57531=>"011010010",
  57532=>"001101000",
  57533=>"111101101",
  57534=>"010010110",
  57535=>"001000010",
  57536=>"101101010",
  57537=>"000101001",
  57538=>"101001000",
  57539=>"011101001",
  57540=>"010010001",
  57541=>"110111011",
  57542=>"000011001",
  57543=>"010001010",
  57544=>"101111000",
  57545=>"111010001",
  57546=>"000110000",
  57547=>"111011101",
  57548=>"000001100",
  57549=>"011010011",
  57550=>"111011110",
  57551=>"010101111",
  57552=>"100001101",
  57553=>"111101111",
  57554=>"100111100",
  57555=>"110101100",
  57556=>"101001001",
  57557=>"101010101",
  57558=>"000001010",
  57559=>"110011000",
  57560=>"101101010",
  57561=>"000011001",
  57562=>"010001110",
  57563=>"000100000",
  57564=>"001010011",
  57565=>"000101011",
  57566=>"001100001",
  57567=>"011110111",
  57568=>"111111101",
  57569=>"000010100",
  57570=>"011110100",
  57571=>"111110110",
  57572=>"001000010",
  57573=>"001100100",
  57574=>"011011010",
  57575=>"001111000",
  57576=>"101010111",
  57577=>"001111111",
  57578=>"110100110",
  57579=>"001111001",
  57580=>"101011000",
  57581=>"110001101",
  57582=>"100011101",
  57583=>"010011100",
  57584=>"100001000",
  57585=>"111111001",
  57586=>"001101000",
  57587=>"100100001",
  57588=>"001001010",
  57589=>"010000010",
  57590=>"111010010",
  57591=>"110001000",
  57592=>"100000001",
  57593=>"000101101",
  57594=>"110111001",
  57595=>"000001111",
  57596=>"111110111",
  57597=>"000110011",
  57598=>"111010100",
  57599=>"010011000",
  57600=>"110010000",
  57601=>"000000010",
  57602=>"011001011",
  57603=>"111001110",
  57604=>"100111001",
  57605=>"001000001",
  57606=>"100011100",
  57607=>"101100001",
  57608=>"101110100",
  57609=>"101001001",
  57610=>"001010010",
  57611=>"010111101",
  57612=>"100001101",
  57613=>"011110110",
  57614=>"101111000",
  57615=>"000000101",
  57616=>"110011000",
  57617=>"000011010",
  57618=>"100100001",
  57619=>"001011010",
  57620=>"010101111",
  57621=>"011111101",
  57622=>"110101110",
  57623=>"100001110",
  57624=>"111001010",
  57625=>"011101101",
  57626=>"010011010",
  57627=>"001011000",
  57628=>"011011001",
  57629=>"101111000",
  57630=>"111110100",
  57631=>"110111100",
  57632=>"100000100",
  57633=>"010001000",
  57634=>"101110110",
  57635=>"110001010",
  57636=>"100100101",
  57637=>"111111111",
  57638=>"011000111",
  57639=>"010011001",
  57640=>"110011011",
  57641=>"000011110",
  57642=>"101111100",
  57643=>"010000010",
  57644=>"111111111",
  57645=>"100100000",
  57646=>"011000100",
  57647=>"011111001",
  57648=>"000100001",
  57649=>"011011100",
  57650=>"111110101",
  57651=>"000111111",
  57652=>"011010010",
  57653=>"011011000",
  57654=>"110101110",
  57655=>"000010101",
  57656=>"001011111",
  57657=>"100110010",
  57658=>"010010110",
  57659=>"110110110",
  57660=>"110111001",
  57661=>"010110100",
  57662=>"011010110",
  57663=>"010110101",
  57664=>"000111101",
  57665=>"011010100",
  57666=>"110101100",
  57667=>"101111100",
  57668=>"001100100",
  57669=>"011111111",
  57670=>"100000001",
  57671=>"011000001",
  57672=>"111111111",
  57673=>"000001000",
  57674=>"100100000",
  57675=>"000010010",
  57676=>"100011100",
  57677=>"010101000",
  57678=>"000100010",
  57679=>"001011101",
  57680=>"111100001",
  57681=>"111000011",
  57682=>"110010001",
  57683=>"010111000",
  57684=>"101000010",
  57685=>"110011011",
  57686=>"111101000",
  57687=>"001001000",
  57688=>"000000000",
  57689=>"001000001",
  57690=>"011101011",
  57691=>"011010100",
  57692=>"011000000",
  57693=>"111111110",
  57694=>"111001011",
  57695=>"111111000",
  57696=>"100111001",
  57697=>"010010000",
  57698=>"100000001",
  57699=>"001110110",
  57700=>"001011100",
  57701=>"000010101",
  57702=>"101110110",
  57703=>"101010100",
  57704=>"010110100",
  57705=>"000100110",
  57706=>"010011010",
  57707=>"011111101",
  57708=>"011111011",
  57709=>"101100000",
  57710=>"001010000",
  57711=>"100010000",
  57712=>"001001100",
  57713=>"001011001",
  57714=>"100000110",
  57715=>"111110111",
  57716=>"011100011",
  57717=>"101010000",
  57718=>"110111001",
  57719=>"000110100",
  57720=>"100000010",
  57721=>"000100100",
  57722=>"111011110",
  57723=>"011100111",
  57724=>"110101100",
  57725=>"000101001",
  57726=>"101100000",
  57727=>"011101000",
  57728=>"111100010",
  57729=>"101001011",
  57730=>"000110010",
  57731=>"011111011",
  57732=>"010010100",
  57733=>"100000010",
  57734=>"100010110",
  57735=>"111111111",
  57736=>"001101000",
  57737=>"100110010",
  57738=>"100000110",
  57739=>"001111110",
  57740=>"000001011",
  57741=>"000101001",
  57742=>"101111010",
  57743=>"001000110",
  57744=>"011110111",
  57745=>"011001000",
  57746=>"000010111",
  57747=>"000010001",
  57748=>"100010101",
  57749=>"101000011",
  57750=>"110000000",
  57751=>"110000101",
  57752=>"001000011",
  57753=>"000100010",
  57754=>"100100011",
  57755=>"000000000",
  57756=>"000011111",
  57757=>"011101001",
  57758=>"000011110",
  57759=>"100011110",
  57760=>"001000011",
  57761=>"101101011",
  57762=>"011001010",
  57763=>"101110100",
  57764=>"001111001",
  57765=>"001100000",
  57766=>"100011000",
  57767=>"000101001",
  57768=>"011110101",
  57769=>"101001001",
  57770=>"101001100",
  57771=>"111011011",
  57772=>"000011001",
  57773=>"100101000",
  57774=>"000111000",
  57775=>"001110010",
  57776=>"111111000",
  57777=>"011011011",
  57778=>"101001001",
  57779=>"100100100",
  57780=>"101100101",
  57781=>"000100011",
  57782=>"000100001",
  57783=>"001110010",
  57784=>"000111100",
  57785=>"101001010",
  57786=>"011001011",
  57787=>"001100101",
  57788=>"100100111",
  57789=>"110010101",
  57790=>"000001010",
  57791=>"011111001",
  57792=>"101011110",
  57793=>"011100110",
  57794=>"011110011",
  57795=>"110110010",
  57796=>"001110010",
  57797=>"110101110",
  57798=>"010100011",
  57799=>"111100111",
  57800=>"101011011",
  57801=>"011111111",
  57802=>"101011100",
  57803=>"100110000",
  57804=>"111111010",
  57805=>"111100111",
  57806=>"000100100",
  57807=>"101110100",
  57808=>"011000010",
  57809=>"001000001",
  57810=>"110101001",
  57811=>"100011101",
  57812=>"101001100",
  57813=>"010100101",
  57814=>"110000000",
  57815=>"010000111",
  57816=>"100101010",
  57817=>"010101111",
  57818=>"111111011",
  57819=>"000101110",
  57820=>"100111111",
  57821=>"010011111",
  57822=>"010001111",
  57823=>"101111101",
  57824=>"100011111",
  57825=>"110001110",
  57826=>"111000100",
  57827=>"100101110",
  57828=>"011110110",
  57829=>"101001111",
  57830=>"000000000",
  57831=>"010010010",
  57832=>"011001010",
  57833=>"111111010",
  57834=>"100000001",
  57835=>"101000101",
  57836=>"110111110",
  57837=>"110000111",
  57838=>"100110110",
  57839=>"111111101",
  57840=>"000011100",
  57841=>"001011011",
  57842=>"000010001",
  57843=>"010110111",
  57844=>"000010000",
  57845=>"000000110",
  57846=>"100101100",
  57847=>"010001010",
  57848=>"101110101",
  57849=>"010010011",
  57850=>"101011010",
  57851=>"010100000",
  57852=>"011110110",
  57853=>"000110101",
  57854=>"110110101",
  57855=>"111110110",
  57856=>"111111011",
  57857=>"111101010",
  57858=>"000101001",
  57859=>"110101111",
  57860=>"011000001",
  57861=>"101100101",
  57862=>"000111100",
  57863=>"111101100",
  57864=>"010001000",
  57865=>"011111111",
  57866=>"111100010",
  57867=>"011010011",
  57868=>"010000001",
  57869=>"100101010",
  57870=>"111010000",
  57871=>"111001111",
  57872=>"100101111",
  57873=>"111110010",
  57874=>"011001011",
  57875=>"001011101",
  57876=>"000100100",
  57877=>"010011000",
  57878=>"111110001",
  57879=>"110010010",
  57880=>"100110110",
  57881=>"010101101",
  57882=>"011001111",
  57883=>"010001110",
  57884=>"011010101",
  57885=>"001111101",
  57886=>"000001111",
  57887=>"001100001",
  57888=>"001001101",
  57889=>"010111011",
  57890=>"111101110",
  57891=>"100111010",
  57892=>"010101001",
  57893=>"101000000",
  57894=>"010000111",
  57895=>"001001011",
  57896=>"001110000",
  57897=>"000110111",
  57898=>"100100101",
  57899=>"011111111",
  57900=>"101110011",
  57901=>"000101011",
  57902=>"101010010",
  57903=>"000000000",
  57904=>"111000110",
  57905=>"100001101",
  57906=>"011010001",
  57907=>"111010100",
  57908=>"010011011",
  57909=>"011010111",
  57910=>"101010010",
  57911=>"011110100",
  57912=>"101110011",
  57913=>"101001011",
  57914=>"110000110",
  57915=>"100111100",
  57916=>"110101011",
  57917=>"000010110",
  57918=>"101100000",
  57919=>"110011010",
  57920=>"101101011",
  57921=>"000001000",
  57922=>"000000100",
  57923=>"111111111",
  57924=>"001011001",
  57925=>"000011101",
  57926=>"101000010",
  57927=>"100111010",
  57928=>"100101110",
  57929=>"010110010",
  57930=>"110110110",
  57931=>"111010111",
  57932=>"111010101",
  57933=>"111100010",
  57934=>"011011111",
  57935=>"111101000",
  57936=>"010010001",
  57937=>"000010101",
  57938=>"011000001",
  57939=>"010001110",
  57940=>"010101011",
  57941=>"111010011",
  57942=>"100000111",
  57943=>"011110101",
  57944=>"110001101",
  57945=>"011101011",
  57946=>"101001111",
  57947=>"111010110",
  57948=>"111000000",
  57949=>"000110111",
  57950=>"000100011",
  57951=>"101011101",
  57952=>"001100000",
  57953=>"111010110",
  57954=>"100010000",
  57955=>"110101110",
  57956=>"101111101",
  57957=>"100000110",
  57958=>"110000100",
  57959=>"111000001",
  57960=>"011010100",
  57961=>"110010010",
  57962=>"101100111",
  57963=>"110101111",
  57964=>"101001100",
  57965=>"111010001",
  57966=>"110110101",
  57967=>"010001100",
  57968=>"111111100",
  57969=>"111111000",
  57970=>"001110011",
  57971=>"110000111",
  57972=>"111111101",
  57973=>"000000100",
  57974=>"000101010",
  57975=>"000100001",
  57976=>"011010100",
  57977=>"111111010",
  57978=>"001000010",
  57979=>"000111101",
  57980=>"101011011",
  57981=>"011001101",
  57982=>"101001011",
  57983=>"001001110",
  57984=>"010101011",
  57985=>"010111011",
  57986=>"000001000",
  57987=>"001110110",
  57988=>"101001110",
  57989=>"100100011",
  57990=>"000001010",
  57991=>"100110000",
  57992=>"001011001",
  57993=>"111111100",
  57994=>"001110111",
  57995=>"101001110",
  57996=>"101010011",
  57997=>"001010001",
  57998=>"010011000",
  57999=>"111001101",
  58000=>"010011001",
  58001=>"001111010",
  58002=>"110110101",
  58003=>"001100001",
  58004=>"000100100",
  58005=>"001111010",
  58006=>"000011011",
  58007=>"000000101",
  58008=>"101101101",
  58009=>"000111001",
  58010=>"101111110",
  58011=>"001101100",
  58012=>"110001101",
  58013=>"111000001",
  58014=>"011000100",
  58015=>"010010110",
  58016=>"000011000",
  58017=>"100000011",
  58018=>"000010111",
  58019=>"110101000",
  58020=>"011100111",
  58021=>"010111011",
  58022=>"000101001",
  58023=>"100100101",
  58024=>"101110000",
  58025=>"000101001",
  58026=>"111110000",
  58027=>"110110100",
  58028=>"010101000",
  58029=>"101100101",
  58030=>"010000101",
  58031=>"101101010",
  58032=>"110100001",
  58033=>"101101100",
  58034=>"110110000",
  58035=>"011000111",
  58036=>"001110100",
  58037=>"000100001",
  58038=>"110111001",
  58039=>"011111111",
  58040=>"101000001",
  58041=>"101010011",
  58042=>"111111010",
  58043=>"111010001",
  58044=>"101011111",
  58045=>"000111111",
  58046=>"001000011",
  58047=>"110111010",
  58048=>"001011001",
  58049=>"000100011",
  58050=>"110000111",
  58051=>"001000010",
  58052=>"000011010",
  58053=>"101010100",
  58054=>"000110000",
  58055=>"110111110",
  58056=>"101110011",
  58057=>"100000000",
  58058=>"110001001",
  58059=>"111001011",
  58060=>"000110001",
  58061=>"101110110",
  58062=>"100010101",
  58063=>"100000100",
  58064=>"111101111",
  58065=>"011010010",
  58066=>"111011110",
  58067=>"010111000",
  58068=>"101001000",
  58069=>"010111111",
  58070=>"100111000",
  58071=>"011000001",
  58072=>"100000011",
  58073=>"001100111",
  58074=>"100101101",
  58075=>"101001000",
  58076=>"111110000",
  58077=>"000000111",
  58078=>"001110100",
  58079=>"011101001",
  58080=>"111111001",
  58081=>"101111101",
  58082=>"110011101",
  58083=>"100111111",
  58084=>"000010101",
  58085=>"011001000",
  58086=>"001011111",
  58087=>"111011100",
  58088=>"111101110",
  58089=>"010101100",
  58090=>"001000110",
  58091=>"010110000",
  58092=>"010000100",
  58093=>"111110100",
  58094=>"011010110",
  58095=>"101011111",
  58096=>"101111111",
  58097=>"101111111",
  58098=>"010000001",
  58099=>"011010000",
  58100=>"101111011",
  58101=>"111011000",
  58102=>"000111010",
  58103=>"111111100",
  58104=>"100000001",
  58105=>"100101011",
  58106=>"100011111",
  58107=>"101010010",
  58108=>"100011111",
  58109=>"010010010",
  58110=>"111110011",
  58111=>"001010001",
  58112=>"010100000",
  58113=>"110001110",
  58114=>"011101101",
  58115=>"111101100",
  58116=>"010001000",
  58117=>"000101000",
  58118=>"111111011",
  58119=>"001000111",
  58120=>"100000000",
  58121=>"000100111",
  58122=>"000010001",
  58123=>"111011000",
  58124=>"001111100",
  58125=>"100110111",
  58126=>"011101001",
  58127=>"010001110",
  58128=>"110100001",
  58129=>"111001000",
  58130=>"001011011",
  58131=>"100000101",
  58132=>"100110101",
  58133=>"011010101",
  58134=>"101000111",
  58135=>"001000011",
  58136=>"101010110",
  58137=>"010011110",
  58138=>"010110100",
  58139=>"110001000",
  58140=>"100100111",
  58141=>"100000001",
  58142=>"010101111",
  58143=>"010100101",
  58144=>"011111101",
  58145=>"000010101",
  58146=>"101001000",
  58147=>"110000001",
  58148=>"110100010",
  58149=>"000111000",
  58150=>"000000000",
  58151=>"101111110",
  58152=>"100001111",
  58153=>"001100101",
  58154=>"111010100",
  58155=>"110010010",
  58156=>"000100011",
  58157=>"100000000",
  58158=>"001000101",
  58159=>"011011110",
  58160=>"100110101",
  58161=>"100111011",
  58162=>"100100010",
  58163=>"101001001",
  58164=>"111010110",
  58165=>"101110110",
  58166=>"000010000",
  58167=>"110000110",
  58168=>"001011011",
  58169=>"101100101",
  58170=>"001011000",
  58171=>"101101011",
  58172=>"100001010",
  58173=>"001000000",
  58174=>"101011001",
  58175=>"110100111",
  58176=>"110101111",
  58177=>"011110010",
  58178=>"111100111",
  58179=>"111011010",
  58180=>"000001011",
  58181=>"011110110",
  58182=>"001000000",
  58183=>"111101111",
  58184=>"111010000",
  58185=>"011111010",
  58186=>"000011001",
  58187=>"010011101",
  58188=>"000000011",
  58189=>"001001100",
  58190=>"011001000",
  58191=>"000011000",
  58192=>"000001001",
  58193=>"101100111",
  58194=>"110110011",
  58195=>"001000011",
  58196=>"111101010",
  58197=>"010001110",
  58198=>"000100110",
  58199=>"001001011",
  58200=>"010100010",
  58201=>"100100001",
  58202=>"100100101",
  58203=>"000100011",
  58204=>"010001100",
  58205=>"010101011",
  58206=>"100010110",
  58207=>"110000010",
  58208=>"100101101",
  58209=>"111100010",
  58210=>"011001001",
  58211=>"011111100",
  58212=>"010011000",
  58213=>"111111011",
  58214=>"011100001",
  58215=>"010001110",
  58216=>"011000111",
  58217=>"001111111",
  58218=>"011101010",
  58219=>"111101001",
  58220=>"101100001",
  58221=>"101001001",
  58222=>"001000100",
  58223=>"011011000",
  58224=>"000000011",
  58225=>"101110111",
  58226=>"111011110",
  58227=>"111101110",
  58228=>"000000101",
  58229=>"010100101",
  58230=>"100111101",
  58231=>"001000110",
  58232=>"111111101",
  58233=>"011001000",
  58234=>"111101010",
  58235=>"001001010",
  58236=>"111001000",
  58237=>"111011100",
  58238=>"111110111",
  58239=>"000110001",
  58240=>"100100001",
  58241=>"001010101",
  58242=>"001011101",
  58243=>"111010100",
  58244=>"011111100",
  58245=>"000101100",
  58246=>"101110111",
  58247=>"110110010",
  58248=>"001101001",
  58249=>"110110000",
  58250=>"111100000",
  58251=>"001011110",
  58252=>"010110101",
  58253=>"101001111",
  58254=>"111001111",
  58255=>"110100111",
  58256=>"101000100",
  58257=>"001011011",
  58258=>"101001001",
  58259=>"111000101",
  58260=>"011000001",
  58261=>"100001001",
  58262=>"011011100",
  58263=>"010001000",
  58264=>"000001101",
  58265=>"111101001",
  58266=>"111001001",
  58267=>"011001111",
  58268=>"000001000",
  58269=>"101110000",
  58270=>"000100110",
  58271=>"001111100",
  58272=>"110011111",
  58273=>"111101001",
  58274=>"010101000",
  58275=>"011111110",
  58276=>"111110111",
  58277=>"001111000",
  58278=>"101010100",
  58279=>"000011110",
  58280=>"000000001",
  58281=>"111000111",
  58282=>"000100111",
  58283=>"010101100",
  58284=>"100000001",
  58285=>"010000111",
  58286=>"011010110",
  58287=>"001011101",
  58288=>"110111110",
  58289=>"010111111",
  58290=>"100110010",
  58291=>"011000011",
  58292=>"011110110",
  58293=>"011010000",
  58294=>"010101000",
  58295=>"110001110",
  58296=>"001011010",
  58297=>"111101010",
  58298=>"100100010",
  58299=>"101010001",
  58300=>"110000101",
  58301=>"100111011",
  58302=>"000011001",
  58303=>"011111010",
  58304=>"010110110",
  58305=>"111111011",
  58306=>"010110010",
  58307=>"100110011",
  58308=>"010011000",
  58309=>"100100110",
  58310=>"001101100",
  58311=>"000000010",
  58312=>"001000000",
  58313=>"101101001",
  58314=>"011101000",
  58315=>"111010011",
  58316=>"010101011",
  58317=>"100110010",
  58318=>"100111100",
  58319=>"000011000",
  58320=>"100111101",
  58321=>"100000001",
  58322=>"011111111",
  58323=>"000000010",
  58324=>"000010010",
  58325=>"011100011",
  58326=>"011101011",
  58327=>"101001011",
  58328=>"000111000",
  58329=>"011001011",
  58330=>"110111110",
  58331=>"100001000",
  58332=>"100110110",
  58333=>"110011111",
  58334=>"111001001",
  58335=>"110000101",
  58336=>"100011001",
  58337=>"001100001",
  58338=>"110111110",
  58339=>"001100110",
  58340=>"100000010",
  58341=>"010010001",
  58342=>"011100011",
  58343=>"111111100",
  58344=>"101111000",
  58345=>"110110100",
  58346=>"111100101",
  58347=>"001100100",
  58348=>"000100111",
  58349=>"101110011",
  58350=>"111001010",
  58351=>"110111101",
  58352=>"000001000",
  58353=>"000000111",
  58354=>"111111101",
  58355=>"011011110",
  58356=>"000111100",
  58357=>"011001110",
  58358=>"000010111",
  58359=>"111110010",
  58360=>"010011100",
  58361=>"011001111",
  58362=>"110101111",
  58363=>"110100011",
  58364=>"000001110",
  58365=>"110011100",
  58366=>"111010000",
  58367=>"011011000",
  58368=>"010111111",
  58369=>"011001010",
  58370=>"001101000",
  58371=>"011010000",
  58372=>"000101110",
  58373=>"010000010",
  58374=>"100001111",
  58375=>"110110011",
  58376=>"001000000",
  58377=>"110000001",
  58378=>"101100100",
  58379=>"011111100",
  58380=>"111100000",
  58381=>"001001110",
  58382=>"111010110",
  58383=>"100100000",
  58384=>"001110011",
  58385=>"000100110",
  58386=>"001010111",
  58387=>"011101100",
  58388=>"110010011",
  58389=>"010100110",
  58390=>"111011110",
  58391=>"000001001",
  58392=>"111100011",
  58393=>"000100010",
  58394=>"001000100",
  58395=>"110111111",
  58396=>"111000000",
  58397=>"011000110",
  58398=>"010011011",
  58399=>"000000010",
  58400=>"111100100",
  58401=>"100001011",
  58402=>"000001101",
  58403=>"111011111",
  58404=>"110000011",
  58405=>"010100000",
  58406=>"111011010",
  58407=>"011010001",
  58408=>"000110010",
  58409=>"000111000",
  58410=>"110001001",
  58411=>"111000011",
  58412=>"001000010",
  58413=>"001011111",
  58414=>"010001001",
  58415=>"011001110",
  58416=>"111101011",
  58417=>"000000001",
  58418=>"010111100",
  58419=>"110110000",
  58420=>"010110111",
  58421=>"100101101",
  58422=>"011100010",
  58423=>"111110110",
  58424=>"100010101",
  58425=>"001011100",
  58426=>"011010111",
  58427=>"011001011",
  58428=>"000010110",
  58429=>"110100110",
  58430=>"101110110",
  58431=>"110000100",
  58432=>"100001001",
  58433=>"010011011",
  58434=>"110111100",
  58435=>"010111110",
  58436=>"011001010",
  58437=>"111001100",
  58438=>"001011011",
  58439=>"101011111",
  58440=>"110100101",
  58441=>"001101000",
  58442=>"010010011",
  58443=>"011100010",
  58444=>"110111001",
  58445=>"011101111",
  58446=>"000000100",
  58447=>"100011000",
  58448=>"111011011",
  58449=>"000000101",
  58450=>"101000001",
  58451=>"011100110",
  58452=>"001010001",
  58453=>"111110110",
  58454=>"100011000",
  58455=>"000000101",
  58456=>"111011001",
  58457=>"001111110",
  58458=>"111011010",
  58459=>"001000000",
  58460=>"100010000",
  58461=>"100011010",
  58462=>"001110010",
  58463=>"110101000",
  58464=>"100001001",
  58465=>"011101110",
  58466=>"000111111",
  58467=>"011111001",
  58468=>"100001000",
  58469=>"100100110",
  58470=>"101001111",
  58471=>"100100101",
  58472=>"110100000",
  58473=>"001101100",
  58474=>"100000110",
  58475=>"011001010",
  58476=>"000111101",
  58477=>"000110100",
  58478=>"100001000",
  58479=>"111100011",
  58480=>"101001110",
  58481=>"101001000",
  58482=>"001101011",
  58483=>"101010000",
  58484=>"110010101",
  58485=>"101110111",
  58486=>"100011101",
  58487=>"001001001",
  58488=>"001100101",
  58489=>"011101000",
  58490=>"101001011",
  58491=>"111111111",
  58492=>"001001111",
  58493=>"001111000",
  58494=>"000001111",
  58495=>"100110000",
  58496=>"001111101",
  58497=>"111111111",
  58498=>"111101110",
  58499=>"101001010",
  58500=>"000010100",
  58501=>"100001111",
  58502=>"001101000",
  58503=>"111100011",
  58504=>"111011001",
  58505=>"110101001",
  58506=>"101110011",
  58507=>"110111011",
  58508=>"100110110",
  58509=>"000011100",
  58510=>"010111101",
  58511=>"101111100",
  58512=>"101011111",
  58513=>"010110101",
  58514=>"000001011",
  58515=>"101001100",
  58516=>"111110101",
  58517=>"011100110",
  58518=>"010110101",
  58519=>"011110000",
  58520=>"101100101",
  58521=>"001101100",
  58522=>"010100000",
  58523=>"101011010",
  58524=>"100110001",
  58525=>"100011100",
  58526=>"110111010",
  58527=>"010001011",
  58528=>"101101110",
  58529=>"111110010",
  58530=>"101000000",
  58531=>"010001101",
  58532=>"110110001",
  58533=>"110111101",
  58534=>"011100110",
  58535=>"110010011",
  58536=>"000011111",
  58537=>"001011100",
  58538=>"011110100",
  58539=>"111011101",
  58540=>"010010101",
  58541=>"101111001",
  58542=>"110011101",
  58543=>"111100001",
  58544=>"010000001",
  58545=>"010011011",
  58546=>"111010100",
  58547=>"100100101",
  58548=>"010100010",
  58549=>"111111111",
  58550=>"011110101",
  58551=>"010000000",
  58552=>"001111000",
  58553=>"001111100",
  58554=>"000110110",
  58555=>"110000010",
  58556=>"101010100",
  58557=>"000001110",
  58558=>"111010001",
  58559=>"101001100",
  58560=>"000011000",
  58561=>"000101111",
  58562=>"111010110",
  58563=>"000001101",
  58564=>"100110001",
  58565=>"110101111",
  58566=>"000000011",
  58567=>"100100111",
  58568=>"001110000",
  58569=>"110000011",
  58570=>"110110101",
  58571=>"100100100",
  58572=>"101001001",
  58573=>"101000111",
  58574=>"100000100",
  58575=>"010101111",
  58576=>"101001111",
  58577=>"001101100",
  58578=>"100011100",
  58579=>"100111001",
  58580=>"001001101",
  58581=>"100101001",
  58582=>"000110100",
  58583=>"100011011",
  58584=>"001110010",
  58585=>"001101011",
  58586=>"001100011",
  58587=>"101001111",
  58588=>"101111010",
  58589=>"010101010",
  58590=>"101111000",
  58591=>"000010110",
  58592=>"100100110",
  58593=>"100100110",
  58594=>"110110100",
  58595=>"000011111",
  58596=>"011100110",
  58597=>"010101111",
  58598=>"011011111",
  58599=>"110111110",
  58600=>"110101001",
  58601=>"101001000",
  58602=>"001100011",
  58603=>"001011010",
  58604=>"100111100",
  58605=>"001000000",
  58606=>"110010010",
  58607=>"110110010",
  58608=>"101101110",
  58609=>"101010101",
  58610=>"101001111",
  58611=>"101000101",
  58612=>"111100111",
  58613=>"000010100",
  58614=>"010100100",
  58615=>"100100101",
  58616=>"111101111",
  58617=>"001010101",
  58618=>"001110010",
  58619=>"000000110",
  58620=>"000100010",
  58621=>"111001011",
  58622=>"100111101",
  58623=>"101111111",
  58624=>"000011101",
  58625=>"001110011",
  58626=>"100110101",
  58627=>"000101110",
  58628=>"111101001",
  58629=>"101001111",
  58630=>"111011100",
  58631=>"000101010",
  58632=>"110011101",
  58633=>"101000101",
  58634=>"100100010",
  58635=>"100001001",
  58636=>"000100001",
  58637=>"100010011",
  58638=>"000000010",
  58639=>"000111011",
  58640=>"110100111",
  58641=>"110001100",
  58642=>"010101011",
  58643=>"110001010",
  58644=>"101101010",
  58645=>"101111111",
  58646=>"000010000",
  58647=>"011110101",
  58648=>"000001010",
  58649=>"101001000",
  58650=>"010000011",
  58651=>"101101011",
  58652=>"111011000",
  58653=>"101001111",
  58654=>"100000101",
  58655=>"101100010",
  58656=>"110011101",
  58657=>"011001010",
  58658=>"011100000",
  58659=>"101101000",
  58660=>"100110001",
  58661=>"010010111",
  58662=>"001111101",
  58663=>"010000001",
  58664=>"110111001",
  58665=>"000101010",
  58666=>"101110111",
  58667=>"101101110",
  58668=>"110001111",
  58669=>"111110111",
  58670=>"000101100",
  58671=>"001001001",
  58672=>"101110101",
  58673=>"110111010",
  58674=>"011011001",
  58675=>"100111111",
  58676=>"101010100",
  58677=>"000001000",
  58678=>"110110100",
  58679=>"001111101",
  58680=>"101000000",
  58681=>"101111000",
  58682=>"101111111",
  58683=>"100100111",
  58684=>"110000010",
  58685=>"111000101",
  58686=>"100000111",
  58687=>"100011010",
  58688=>"101111001",
  58689=>"000010100",
  58690=>"011111001",
  58691=>"101001001",
  58692=>"111111101",
  58693=>"010011011",
  58694=>"011010100",
  58695=>"100110011",
  58696=>"110111101",
  58697=>"110001001",
  58698=>"011000100",
  58699=>"100101101",
  58700=>"010101011",
  58701=>"011111101",
  58702=>"110011010",
  58703=>"000010010",
  58704=>"010011011",
  58705=>"101101101",
  58706=>"110010000",
  58707=>"001111011",
  58708=>"101111111",
  58709=>"000101101",
  58710=>"011000010",
  58711=>"100010111",
  58712=>"000001100",
  58713=>"010000000",
  58714=>"111101101",
  58715=>"111101000",
  58716=>"011000100",
  58717=>"111101101",
  58718=>"011010001",
  58719=>"011110110",
  58720=>"000100010",
  58721=>"000110111",
  58722=>"010011100",
  58723=>"010101001",
  58724=>"101101001",
  58725=>"010000001",
  58726=>"010010100",
  58727=>"000011101",
  58728=>"011011101",
  58729=>"100110011",
  58730=>"010011100",
  58731=>"110101101",
  58732=>"101000001",
  58733=>"101000010",
  58734=>"110101110",
  58735=>"111100001",
  58736=>"011000010",
  58737=>"100111100",
  58738=>"100001001",
  58739=>"010000101",
  58740=>"010111000",
  58741=>"101000001",
  58742=>"000110000",
  58743=>"000000110",
  58744=>"001100000",
  58745=>"011110010",
  58746=>"010100000",
  58747=>"111111011",
  58748=>"010101110",
  58749=>"001111011",
  58750=>"110010001",
  58751=>"010110110",
  58752=>"101110100",
  58753=>"010000011",
  58754=>"100101101",
  58755=>"110001101",
  58756=>"010001110",
  58757=>"000010001",
  58758=>"101001101",
  58759=>"110100100",
  58760=>"010010100",
  58761=>"101001101",
  58762=>"010011100",
  58763=>"111110110",
  58764=>"000100110",
  58765=>"110101110",
  58766=>"000101111",
  58767=>"111101001",
  58768=>"111100111",
  58769=>"100111101",
  58770=>"011011111",
  58771=>"111000000",
  58772=>"010110001",
  58773=>"111000000",
  58774=>"110101010",
  58775=>"010100001",
  58776=>"010100100",
  58777=>"000101110",
  58778=>"101111111",
  58779=>"110011111",
  58780=>"011010010",
  58781=>"100101110",
  58782=>"010010001",
  58783=>"111001000",
  58784=>"110111101",
  58785=>"011100000",
  58786=>"000010100",
  58787=>"011100101",
  58788=>"011001000",
  58789=>"000001000",
  58790=>"001000101",
  58791=>"111101100",
  58792=>"110101101",
  58793=>"010010001",
  58794=>"001101000",
  58795=>"101011101",
  58796=>"000110001",
  58797=>"001110100",
  58798=>"101100011",
  58799=>"010101001",
  58800=>"101000001",
  58801=>"100110101",
  58802=>"000100000",
  58803=>"100101011",
  58804=>"010001000",
  58805=>"110011000",
  58806=>"001100110",
  58807=>"010000100",
  58808=>"110000001",
  58809=>"010111001",
  58810=>"000110001",
  58811=>"010011110",
  58812=>"001111001",
  58813=>"000010000",
  58814=>"000010001",
  58815=>"010100010",
  58816=>"001101011",
  58817=>"110001101",
  58818=>"011101011",
  58819=>"101001101",
  58820=>"111011111",
  58821=>"101011011",
  58822=>"110111111",
  58823=>"101110000",
  58824=>"110001111",
  58825=>"111001010",
  58826=>"110010000",
  58827=>"010001100",
  58828=>"101111101",
  58829=>"101100000",
  58830=>"000000010",
  58831=>"001010011",
  58832=>"111101001",
  58833=>"111111011",
  58834=>"010001011",
  58835=>"010010001",
  58836=>"110001110",
  58837=>"011001011",
  58838=>"000110110",
  58839=>"100110110",
  58840=>"010000000",
  58841=>"111011111",
  58842=>"111111001",
  58843=>"001111000",
  58844=>"101110111",
  58845=>"000010111",
  58846=>"010011000",
  58847=>"111001100",
  58848=>"111011111",
  58849=>"100111001",
  58850=>"000110111",
  58851=>"111111000",
  58852=>"110010010",
  58853=>"000101111",
  58854=>"111100001",
  58855=>"010000001",
  58856=>"101011000",
  58857=>"111110100",
  58858=>"100110100",
  58859=>"111110110",
  58860=>"000110001",
  58861=>"000101010",
  58862=>"101000001",
  58863=>"101110001",
  58864=>"011001011",
  58865=>"101010011",
  58866=>"011000001",
  58867=>"000000100",
  58868=>"100100010",
  58869=>"010001010",
  58870=>"010101001",
  58871=>"000001111",
  58872=>"010100101",
  58873=>"000100000",
  58874=>"101100010",
  58875=>"101011000",
  58876=>"100111010",
  58877=>"010111100",
  58878=>"111001111",
  58879=>"010000000",
  58880=>"101011010",
  58881=>"001000000",
  58882=>"000111000",
  58883=>"101000001",
  58884=>"111111011",
  58885=>"111111111",
  58886=>"111010000",
  58887=>"100001011",
  58888=>"011100010",
  58889=>"010110101",
  58890=>"110000011",
  58891=>"010001010",
  58892=>"010111000",
  58893=>"001010010",
  58894=>"000000000",
  58895=>"111111101",
  58896=>"000101010",
  58897=>"010101110",
  58898=>"111001011",
  58899=>"100100000",
  58900=>"011101000",
  58901=>"111010011",
  58902=>"111111100",
  58903=>"001000001",
  58904=>"001001000",
  58905=>"111100100",
  58906=>"111100010",
  58907=>"110101011",
  58908=>"000110101",
  58909=>"001001110",
  58910=>"101010001",
  58911=>"111111001",
  58912=>"110111011",
  58913=>"011001001",
  58914=>"010010111",
  58915=>"000111111",
  58916=>"110010000",
  58917=>"000101011",
  58918=>"011001111",
  58919=>"110001011",
  58920=>"110010011",
  58921=>"001100010",
  58922=>"100101101",
  58923=>"111101101",
  58924=>"000101000",
  58925=>"101000000",
  58926=>"110111101",
  58927=>"000000100",
  58928=>"010111010",
  58929=>"110101001",
  58930=>"001000010",
  58931=>"110111111",
  58932=>"011011111",
  58933=>"001110100",
  58934=>"100011011",
  58935=>"010010001",
  58936=>"101011000",
  58937=>"111100101",
  58938=>"010010000",
  58939=>"011101110",
  58940=>"010101100",
  58941=>"011000100",
  58942=>"000110010",
  58943=>"000110111",
  58944=>"000100000",
  58945=>"000011000",
  58946=>"111000010",
  58947=>"111010111",
  58948=>"101010010",
  58949=>"111111101",
  58950=>"010000011",
  58951=>"101010101",
  58952=>"001110001",
  58953=>"011101111",
  58954=>"110100110",
  58955=>"111010011",
  58956=>"011001101",
  58957=>"111111000",
  58958=>"111010111",
  58959=>"110100010",
  58960=>"011110111",
  58961=>"010001000",
  58962=>"001011101",
  58963=>"110001011",
  58964=>"000010000",
  58965=>"111011100",
  58966=>"111111001",
  58967=>"011011011",
  58968=>"001100101",
  58969=>"000100110",
  58970=>"000001001",
  58971=>"010101110",
  58972=>"001011100",
  58973=>"000110000",
  58974=>"011100001",
  58975=>"110010101",
  58976=>"100011001",
  58977=>"001101001",
  58978=>"001010110",
  58979=>"111000011",
  58980=>"010110111",
  58981=>"011101010",
  58982=>"101000111",
  58983=>"111110110",
  58984=>"011011111",
  58985=>"111010110",
  58986=>"011001101",
  58987=>"110111011",
  58988=>"110110001",
  58989=>"000101000",
  58990=>"010100011",
  58991=>"001111010",
  58992=>"000111001",
  58993=>"100011000",
  58994=>"011011011",
  58995=>"010010101",
  58996=>"110011010",
  58997=>"111100110",
  58998=>"101001000",
  58999=>"101010111",
  59000=>"010010001",
  59001=>"101101111",
  59002=>"111011001",
  59003=>"010000110",
  59004=>"001010000",
  59005=>"111111110",
  59006=>"110110001",
  59007=>"110100100",
  59008=>"001011100",
  59009=>"001111000",
  59010=>"110100000",
  59011=>"101111110",
  59012=>"100110000",
  59013=>"001011010",
  59014=>"100111110",
  59015=>"111110100",
  59016=>"011010001",
  59017=>"000001001",
  59018=>"110010101",
  59019=>"001100000",
  59020=>"000001010",
  59021=>"100101001",
  59022=>"101000001",
  59023=>"101111010",
  59024=>"011010000",
  59025=>"111001010",
  59026=>"111001001",
  59027=>"111110110",
  59028=>"101001010",
  59029=>"011001010",
  59030=>"010101001",
  59031=>"110010100",
  59032=>"001001010",
  59033=>"000001100",
  59034=>"101001101",
  59035=>"011111011",
  59036=>"001101110",
  59037=>"010101111",
  59038=>"110011101",
  59039=>"110110101",
  59040=>"010111010",
  59041=>"110111100",
  59042=>"010111110",
  59043=>"010111101",
  59044=>"100000110",
  59045=>"010000000",
  59046=>"001101110",
  59047=>"000001000",
  59048=>"011111000",
  59049=>"010010100",
  59050=>"010011101",
  59051=>"000100110",
  59052=>"000100011",
  59053=>"001101011",
  59054=>"001100010",
  59055=>"010101010",
  59056=>"010001000",
  59057=>"001100111",
  59058=>"110000100",
  59059=>"010111100",
  59060=>"100001111",
  59061=>"000000011",
  59062=>"001100110",
  59063=>"011101010",
  59064=>"100110011",
  59065=>"001010101",
  59066=>"001110011",
  59067=>"101101001",
  59068=>"101110010",
  59069=>"011000101",
  59070=>"000010100",
  59071=>"101100111",
  59072=>"011001001",
  59073=>"010010111",
  59074=>"110000000",
  59075=>"010011001",
  59076=>"101111011",
  59077=>"010110111",
  59078=>"011100100",
  59079=>"100000010",
  59080=>"010101011",
  59081=>"100000000",
  59082=>"111111110",
  59083=>"000001001",
  59084=>"001100111",
  59085=>"101011110",
  59086=>"000111100",
  59087=>"110111011",
  59088=>"000101001",
  59089=>"110101010",
  59090=>"101100100",
  59091=>"110101000",
  59092=>"010100010",
  59093=>"010011001",
  59094=>"000000110",
  59095=>"100100100",
  59096=>"110011010",
  59097=>"111100100",
  59098=>"000110110",
  59099=>"101101110",
  59100=>"100000010",
  59101=>"011011010",
  59102=>"111100001",
  59103=>"101111001",
  59104=>"000111010",
  59105=>"000111100",
  59106=>"110101000",
  59107=>"101110101",
  59108=>"110111000",
  59109=>"111111011",
  59110=>"111011100",
  59111=>"001110011",
  59112=>"110011101",
  59113=>"010101000",
  59114=>"001011100",
  59115=>"010011010",
  59116=>"011010001",
  59117=>"110101000",
  59118=>"111011010",
  59119=>"111110110",
  59120=>"111011001",
  59121=>"000101000",
  59122=>"000010100",
  59123=>"001010100",
  59124=>"000010101",
  59125=>"111111000",
  59126=>"101110110",
  59127=>"010001110",
  59128=>"111001001",
  59129=>"011100101",
  59130=>"110111000",
  59131=>"010110000",
  59132=>"011110010",
  59133=>"001100010",
  59134=>"001001000",
  59135=>"111010111",
  59136=>"111000101",
  59137=>"000001010",
  59138=>"000000100",
  59139=>"001111101",
  59140=>"011010001",
  59141=>"000111010",
  59142=>"111000110",
  59143=>"100110100",
  59144=>"000100010",
  59145=>"110001110",
  59146=>"011100101",
  59147=>"000001111",
  59148=>"011111110",
  59149=>"100111000",
  59150=>"101100110",
  59151=>"000001010",
  59152=>"000111100",
  59153=>"110111010",
  59154=>"101011001",
  59155=>"000110100",
  59156=>"010100000",
  59157=>"011000101",
  59158=>"111000101",
  59159=>"000011000",
  59160=>"001000000",
  59161=>"001101111",
  59162=>"100111100",
  59163=>"111000101",
  59164=>"101010100",
  59165=>"101000110",
  59166=>"010101000",
  59167=>"001001001",
  59168=>"100111101",
  59169=>"010011000",
  59170=>"000100001",
  59171=>"001011111",
  59172=>"101000110",
  59173=>"110110011",
  59174=>"110101100",
  59175=>"010000110",
  59176=>"111001000",
  59177=>"111001110",
  59178=>"100110010",
  59179=>"111110000",
  59180=>"111000110",
  59181=>"110110010",
  59182=>"000101010",
  59183=>"100000101",
  59184=>"111011000",
  59185=>"101000000",
  59186=>"100101101",
  59187=>"000110001",
  59188=>"111111010",
  59189=>"100111011",
  59190=>"110010110",
  59191=>"110100111",
  59192=>"101111011",
  59193=>"011000101",
  59194=>"010010010",
  59195=>"000110111",
  59196=>"001000011",
  59197=>"111111101",
  59198=>"101001000",
  59199=>"000000100",
  59200=>"010101110",
  59201=>"100000001",
  59202=>"110010100",
  59203=>"011101110",
  59204=>"111001111",
  59205=>"011010001",
  59206=>"101101111",
  59207=>"101000011",
  59208=>"001011110",
  59209=>"111111101",
  59210=>"001000000",
  59211=>"101000001",
  59212=>"110010001",
  59213=>"100100011",
  59214=>"111111100",
  59215=>"001100010",
  59216=>"111111001",
  59217=>"000000111",
  59218=>"110111110",
  59219=>"111111000",
  59220=>"100101001",
  59221=>"111000001",
  59222=>"110100100",
  59223=>"001000110",
  59224=>"000000111",
  59225=>"001000111",
  59226=>"010001010",
  59227=>"111111011",
  59228=>"010111000",
  59229=>"010000110",
  59230=>"110010000",
  59231=>"000010100",
  59232=>"000100011",
  59233=>"110110111",
  59234=>"000110000",
  59235=>"000100000",
  59236=>"111001111",
  59237=>"100100110",
  59238=>"001001101",
  59239=>"011000000",
  59240=>"100010000",
  59241=>"100000010",
  59242=>"010010001",
  59243=>"000100010",
  59244=>"001110001",
  59245=>"101100011",
  59246=>"100010000",
  59247=>"100011110",
  59248=>"011001100",
  59249=>"100110101",
  59250=>"010111010",
  59251=>"111011100",
  59252=>"101010010",
  59253=>"000010001",
  59254=>"111010010",
  59255=>"110010100",
  59256=>"100011010",
  59257=>"100101001",
  59258=>"111101010",
  59259=>"100101110",
  59260=>"100111111",
  59261=>"101000001",
  59262=>"111000101",
  59263=>"000110101",
  59264=>"000101110",
  59265=>"011010011",
  59266=>"101011011",
  59267=>"111010111",
  59268=>"110100101",
  59269=>"000110111",
  59270=>"111110100",
  59271=>"001001100",
  59272=>"100000100",
  59273=>"010111001",
  59274=>"101001010",
  59275=>"001000111",
  59276=>"011011101",
  59277=>"010100111",
  59278=>"100001111",
  59279=>"000111000",
  59280=>"011001111",
  59281=>"110100101",
  59282=>"000001000",
  59283=>"010011101",
  59284=>"010010100",
  59285=>"001111000",
  59286=>"110010110",
  59287=>"000111001",
  59288=>"101101001",
  59289=>"101000011",
  59290=>"000001001",
  59291=>"101111100",
  59292=>"000101110",
  59293=>"111101000",
  59294=>"000101100",
  59295=>"101110001",
  59296=>"010010000",
  59297=>"011011111",
  59298=>"001001100",
  59299=>"001010100",
  59300=>"101011101",
  59301=>"010101101",
  59302=>"101000100",
  59303=>"111010010",
  59304=>"100000100",
  59305=>"011101110",
  59306=>"010000011",
  59307=>"011001101",
  59308=>"110001110",
  59309=>"110001110",
  59310=>"111001010",
  59311=>"100100100",
  59312=>"100011011",
  59313=>"000100000",
  59314=>"011010101",
  59315=>"111101011",
  59316=>"111100010",
  59317=>"000100011",
  59318=>"110011011",
  59319=>"010101001",
  59320=>"111101010",
  59321=>"010110011",
  59322=>"010010001",
  59323=>"010101110",
  59324=>"100101001",
  59325=>"001000101",
  59326=>"110000001",
  59327=>"001011010",
  59328=>"101010010",
  59329=>"100000111",
  59330=>"100011000",
  59331=>"111011111",
  59332=>"100011100",
  59333=>"011101011",
  59334=>"111110111",
  59335=>"111011101",
  59336=>"101101001",
  59337=>"001111011",
  59338=>"111010001",
  59339=>"110100011",
  59340=>"101001000",
  59341=>"110000111",
  59342=>"011011010",
  59343=>"011110011",
  59344=>"000101100",
  59345=>"100100101",
  59346=>"111101101",
  59347=>"100001001",
  59348=>"010011111",
  59349=>"000110101",
  59350=>"011100101",
  59351=>"001010010",
  59352=>"001110001",
  59353=>"110011101",
  59354=>"000000010",
  59355=>"100000000",
  59356=>"010010011",
  59357=>"101101100",
  59358=>"011100111",
  59359=>"110010010",
  59360=>"110101101",
  59361=>"110001100",
  59362=>"111010111",
  59363=>"101001111",
  59364=>"001001010",
  59365=>"111110111",
  59366=>"010001111",
  59367=>"111000001",
  59368=>"000111100",
  59369=>"101110111",
  59370=>"011000110",
  59371=>"110110100",
  59372=>"100000110",
  59373=>"010001100",
  59374=>"010111000",
  59375=>"110011110",
  59376=>"110001100",
  59377=>"101010000",
  59378=>"110010111",
  59379=>"101100011",
  59380=>"111011111",
  59381=>"010010111",
  59382=>"101100000",
  59383=>"100001000",
  59384=>"101101010",
  59385=>"000001111",
  59386=>"001000100",
  59387=>"101011010",
  59388=>"111000000",
  59389=>"100010001",
  59390=>"110110010",
  59391=>"001101001",
  59392=>"000111000",
  59393=>"110000011",
  59394=>"001011011",
  59395=>"000010010",
  59396=>"111100000",
  59397=>"000110001",
  59398=>"011001101",
  59399=>"110011110",
  59400=>"011110100",
  59401=>"011110011",
  59402=>"001101110",
  59403=>"111010100",
  59404=>"001100010",
  59405=>"100011000",
  59406=>"101000000",
  59407=>"001101011",
  59408=>"101110111",
  59409=>"011010010",
  59410=>"111001110",
  59411=>"000011000",
  59412=>"000000011",
  59413=>"011111011",
  59414=>"001111100",
  59415=>"001111111",
  59416=>"010110001",
  59417=>"111101011",
  59418=>"101010111",
  59419=>"000000000",
  59420=>"011011101",
  59421=>"110011111",
  59422=>"010101110",
  59423=>"100010100",
  59424=>"101010010",
  59425=>"011110111",
  59426=>"000101001",
  59427=>"111101111",
  59428=>"001001010",
  59429=>"110000010",
  59430=>"100010011",
  59431=>"001101001",
  59432=>"101001101",
  59433=>"000101000",
  59434=>"110110011",
  59435=>"100111101",
  59436=>"011100011",
  59437=>"000010110",
  59438=>"111111111",
  59439=>"000100100",
  59440=>"000110000",
  59441=>"111111101",
  59442=>"111101100",
  59443=>"011100111",
  59444=>"001000011",
  59445=>"110110001",
  59446=>"011111001",
  59447=>"011010100",
  59448=>"000000001",
  59449=>"100011100",
  59450=>"100010010",
  59451=>"110011001",
  59452=>"001000000",
  59453=>"011100011",
  59454=>"001000100",
  59455=>"000011000",
  59456=>"001010110",
  59457=>"000100101",
  59458=>"101010100",
  59459=>"100101001",
  59460=>"110011001",
  59461=>"111111101",
  59462=>"101111111",
  59463=>"101010011",
  59464=>"000000111",
  59465=>"001001011",
  59466=>"110000010",
  59467=>"001010010",
  59468=>"001010000",
  59469=>"101001000",
  59470=>"111100001",
  59471=>"100111111",
  59472=>"010100000",
  59473=>"010001001",
  59474=>"010001110",
  59475=>"100010101",
  59476=>"110011000",
  59477=>"100011001",
  59478=>"001011101",
  59479=>"000000000",
  59480=>"010011100",
  59481=>"001001011",
  59482=>"101100001",
  59483=>"101111011",
  59484=>"111110101",
  59485=>"101000010",
  59486=>"001101000",
  59487=>"001111111",
  59488=>"100110001",
  59489=>"001001101",
  59490=>"101010100",
  59491=>"100110000",
  59492=>"011011100",
  59493=>"100101111",
  59494=>"111010000",
  59495=>"100110100",
  59496=>"001101010",
  59497=>"111011011",
  59498=>"000011011",
  59499=>"100110110",
  59500=>"110110011",
  59501=>"101111000",
  59502=>"001110011",
  59503=>"000110101",
  59504=>"011110001",
  59505=>"010010010",
  59506=>"011000111",
  59507=>"110111001",
  59508=>"011111100",
  59509=>"000111101",
  59510=>"111111100",
  59511=>"101000000",
  59512=>"100011011",
  59513=>"001001110",
  59514=>"011100011",
  59515=>"110011111",
  59516=>"101001011",
  59517=>"010110111",
  59518=>"111001110",
  59519=>"100100011",
  59520=>"001100000",
  59521=>"001000111",
  59522=>"111011001",
  59523=>"111111111",
  59524=>"101010111",
  59525=>"011000110",
  59526=>"101100001",
  59527=>"110111101",
  59528=>"001011010",
  59529=>"110001101",
  59530=>"000100000",
  59531=>"010000111",
  59532=>"111111111",
  59533=>"000011101",
  59534=>"100100000",
  59535=>"100111100",
  59536=>"101110010",
  59537=>"101101100",
  59538=>"100011110",
  59539=>"110110111",
  59540=>"001010100",
  59541=>"110111000",
  59542=>"111101001",
  59543=>"111100101",
  59544=>"101011111",
  59545=>"111010011",
  59546=>"001111001",
  59547=>"100011000",
  59548=>"100001011",
  59549=>"111011110",
  59550=>"111010010",
  59551=>"110010011",
  59552=>"010100001",
  59553=>"101011100",
  59554=>"111111110",
  59555=>"011101000",
  59556=>"001001101",
  59557=>"001000000",
  59558=>"101101101",
  59559=>"111110010",
  59560=>"000111100",
  59561=>"010000101",
  59562=>"101010110",
  59563=>"011000000",
  59564=>"011001010",
  59565=>"100000000",
  59566=>"101101111",
  59567=>"011011101",
  59568=>"000111101",
  59569=>"000010000",
  59570=>"000000011",
  59571=>"101100010",
  59572=>"000101000",
  59573=>"000010011",
  59574=>"011010010",
  59575=>"001111010",
  59576=>"110000000",
  59577=>"111110001",
  59578=>"000011110",
  59579=>"111111011",
  59580=>"101110000",
  59581=>"100101110",
  59582=>"100001011",
  59583=>"110111100",
  59584=>"111000101",
  59585=>"000010011",
  59586=>"000110001",
  59587=>"111011011",
  59588=>"001101111",
  59589=>"001111110",
  59590=>"001101100",
  59591=>"000010001",
  59592=>"001100101",
  59593=>"001101101",
  59594=>"110100110",
  59595=>"110110011",
  59596=>"110010111",
  59597=>"101001010",
  59598=>"100000010",
  59599=>"100011100",
  59600=>"000110111",
  59601=>"011111000",
  59602=>"100001010",
  59603=>"000100111",
  59604=>"011101000",
  59605=>"010111111",
  59606=>"000001101",
  59607=>"011010110",
  59608=>"001111001",
  59609=>"011001000",
  59610=>"100100110",
  59611=>"100000010",
  59612=>"000110010",
  59613=>"011110011",
  59614=>"100011101",
  59615=>"101100001",
  59616=>"111110110",
  59617=>"001100100",
  59618=>"110111111",
  59619=>"000011010",
  59620=>"110010100",
  59621=>"101101010",
  59622=>"101110110",
  59623=>"000101000",
  59624=>"001000100",
  59625=>"110100111",
  59626=>"101010010",
  59627=>"111000000",
  59628=>"000111101",
  59629=>"000111111",
  59630=>"100011100",
  59631=>"100011100",
  59632=>"000000100",
  59633=>"110000000",
  59634=>"100110011",
  59635=>"110010000",
  59636=>"101000010",
  59637=>"101111001",
  59638=>"111111111",
  59639=>"000101000",
  59640=>"000100011",
  59641=>"000111000",
  59642=>"001000010",
  59643=>"010101111",
  59644=>"001101110",
  59645=>"101101100",
  59646=>"111011000",
  59647=>"001101000",
  59648=>"000110010",
  59649=>"101000000",
  59650=>"111010111",
  59651=>"101000011",
  59652=>"000111011",
  59653=>"000111010",
  59654=>"011110010",
  59655=>"111001110",
  59656=>"010000011",
  59657=>"001110111",
  59658=>"100110100",
  59659=>"001010101",
  59660=>"011000011",
  59661=>"100000000",
  59662=>"110100101",
  59663=>"000000100",
  59664=>"000001011",
  59665=>"101111111",
  59666=>"001000001",
  59667=>"100000001",
  59668=>"011010001",
  59669=>"101011111",
  59670=>"100110101",
  59671=>"110111000",
  59672=>"001000011",
  59673=>"101101101",
  59674=>"001110110",
  59675=>"110001110",
  59676=>"011110000",
  59677=>"101101001",
  59678=>"101111010",
  59679=>"011011111",
  59680=>"011010001",
  59681=>"001110011",
  59682=>"011010000",
  59683=>"101000000",
  59684=>"111001001",
  59685=>"100100000",
  59686=>"101100010",
  59687=>"101010101",
  59688=>"000001111",
  59689=>"111110010",
  59690=>"001111110",
  59691=>"000000100",
  59692=>"001111110",
  59693=>"101011111",
  59694=>"101000110",
  59695=>"101010101",
  59696=>"001100001",
  59697=>"101001101",
  59698=>"000001000",
  59699=>"001101101",
  59700=>"010000100",
  59701=>"001101010",
  59702=>"101001100",
  59703=>"100001011",
  59704=>"100100001",
  59705=>"011010111",
  59706=>"001000010",
  59707=>"000010011",
  59708=>"111100101",
  59709=>"000100011",
  59710=>"101111100",
  59711=>"010111001",
  59712=>"000100001",
  59713=>"111111001",
  59714=>"011110111",
  59715=>"100001110",
  59716=>"010000100",
  59717=>"110010010",
  59718=>"001010101",
  59719=>"100001101",
  59720=>"010010011",
  59721=>"000011000",
  59722=>"011001000",
  59723=>"001000001",
  59724=>"001110001",
  59725=>"101001100",
  59726=>"100101001",
  59727=>"110111101",
  59728=>"111101101",
  59729=>"001100000",
  59730=>"111100100",
  59731=>"000000010",
  59732=>"101110011",
  59733=>"011101000",
  59734=>"110001100",
  59735=>"110001111",
  59736=>"010101110",
  59737=>"000000101",
  59738=>"000111011",
  59739=>"011100011",
  59740=>"100110000",
  59741=>"011001011",
  59742=>"000100100",
  59743=>"000101010",
  59744=>"000110110",
  59745=>"000100001",
  59746=>"110010000",
  59747=>"100011010",
  59748=>"100110110",
  59749=>"000010011",
  59750=>"100011000",
  59751=>"000010000",
  59752=>"100100110",
  59753=>"110100100",
  59754=>"010111100",
  59755=>"111101001",
  59756=>"001101111",
  59757=>"110011001",
  59758=>"101000000",
  59759=>"010001001",
  59760=>"100001000",
  59761=>"110010011",
  59762=>"110100000",
  59763=>"011010000",
  59764=>"011010011",
  59765=>"101011111",
  59766=>"000000001",
  59767=>"011011000",
  59768=>"110111010",
  59769=>"010010001",
  59770=>"000001111",
  59771=>"110101010",
  59772=>"110001001",
  59773=>"111101101",
  59774=>"101010011",
  59775=>"000011101",
  59776=>"000001101",
  59777=>"010100010",
  59778=>"001111001",
  59779=>"111110010",
  59780=>"111000011",
  59781=>"101110001",
  59782=>"011100000",
  59783=>"110000110",
  59784=>"000000011",
  59785=>"001110000",
  59786=>"111001011",
  59787=>"100011001",
  59788=>"100101000",
  59789=>"011111110",
  59790=>"001100000",
  59791=>"001000010",
  59792=>"001111100",
  59793=>"010001001",
  59794=>"100111011",
  59795=>"101010100",
  59796=>"011101001",
  59797=>"110101000",
  59798=>"110101100",
  59799=>"101011011",
  59800=>"100100000",
  59801=>"111000110",
  59802=>"001100100",
  59803=>"011100001",
  59804=>"001000100",
  59805=>"101000001",
  59806=>"100111000",
  59807=>"001100010",
  59808=>"101100101",
  59809=>"001111111",
  59810=>"001101100",
  59811=>"111000001",
  59812=>"000100111",
  59813=>"100011010",
  59814=>"011011100",
  59815=>"001111111",
  59816=>"111011111",
  59817=>"001001000",
  59818=>"100011000",
  59819=>"010001011",
  59820=>"011011001",
  59821=>"100101000",
  59822=>"110110111",
  59823=>"100011100",
  59824=>"000001001",
  59825=>"101100010",
  59826=>"011100000",
  59827=>"000001110",
  59828=>"110111010",
  59829=>"010111010",
  59830=>"111110111",
  59831=>"111110100",
  59832=>"111110010",
  59833=>"101011000",
  59834=>"000000010",
  59835=>"010000001",
  59836=>"111101110",
  59837=>"011101011",
  59838=>"001010001",
  59839=>"000111000",
  59840=>"101111011",
  59841=>"010111101",
  59842=>"101100001",
  59843=>"011101001",
  59844=>"110110011",
  59845=>"000100101",
  59846=>"001101010",
  59847=>"000110010",
  59848=>"001000101",
  59849=>"111001000",
  59850=>"000010110",
  59851=>"110110111",
  59852=>"001101000",
  59853=>"010111100",
  59854=>"000000000",
  59855=>"101001010",
  59856=>"110101011",
  59857=>"111011010",
  59858=>"100001001",
  59859=>"001101111",
  59860=>"111100011",
  59861=>"001010110",
  59862=>"001010100",
  59863=>"001000010",
  59864=>"001100100",
  59865=>"100011110",
  59866=>"101000110",
  59867=>"110101100",
  59868=>"111010000",
  59869=>"100101101",
  59870=>"111111101",
  59871=>"010011011",
  59872=>"011100100",
  59873=>"001000010",
  59874=>"010100001",
  59875=>"101001011",
  59876=>"010000000",
  59877=>"111110110",
  59878=>"110011010",
  59879=>"101101011",
  59880=>"111101110",
  59881=>"000000101",
  59882=>"000101100",
  59883=>"000010110",
  59884=>"010110101",
  59885=>"110011000",
  59886=>"111000100",
  59887=>"101101100",
  59888=>"110000011",
  59889=>"011111011",
  59890=>"101110010",
  59891=>"010001101",
  59892=>"110011000",
  59893=>"110011101",
  59894=>"000110101",
  59895=>"010111001",
  59896=>"101010000",
  59897=>"110010100",
  59898=>"000110010",
  59899=>"110111010",
  59900=>"101100000",
  59901=>"001000001",
  59902=>"111100111",
  59903=>"001111011",
  59904=>"111101110",
  59905=>"010001110",
  59906=>"111111111",
  59907=>"001010100",
  59908=>"010001000",
  59909=>"111011100",
  59910=>"110110001",
  59911=>"011111111",
  59912=>"111111111",
  59913=>"010111100",
  59914=>"110000010",
  59915=>"111010001",
  59916=>"100100101",
  59917=>"010111011",
  59918=>"101111000",
  59919=>"111000111",
  59920=>"101101100",
  59921=>"010100110",
  59922=>"010001011",
  59923=>"000101100",
  59924=>"000100100",
  59925=>"011000001",
  59926=>"010010010",
  59927=>"000010111",
  59928=>"110110010",
  59929=>"111110101",
  59930=>"010011101",
  59931=>"011000000",
  59932=>"110101010",
  59933=>"000000101",
  59934=>"010101000",
  59935=>"010001100",
  59936=>"011110001",
  59937=>"101111101",
  59938=>"000111001",
  59939=>"000100001",
  59940=>"111010101",
  59941=>"100010000",
  59942=>"010010001",
  59943=>"010000001",
  59944=>"000010001",
  59945=>"110111011",
  59946=>"110100110",
  59947=>"011010010",
  59948=>"111010001",
  59949=>"001010001",
  59950=>"000101101",
  59951=>"111001100",
  59952=>"110000101",
  59953=>"011101110",
  59954=>"111001011",
  59955=>"100010000",
  59956=>"001001011",
  59957=>"010010001",
  59958=>"110101011",
  59959=>"111001010",
  59960=>"111011100",
  59961=>"110010010",
  59962=>"110011000",
  59963=>"001001000",
  59964=>"111000101",
  59965=>"110010000",
  59966=>"000111011",
  59967=>"101001100",
  59968=>"111110010",
  59969=>"000111100",
  59970=>"000001011",
  59971=>"101101010",
  59972=>"100100011",
  59973=>"101001100",
  59974=>"001110100",
  59975=>"110100011",
  59976=>"010010010",
  59977=>"100111110",
  59978=>"111100011",
  59979=>"010000000",
  59980=>"101101010",
  59981=>"100110100",
  59982=>"011101001",
  59983=>"010001001",
  59984=>"000011011",
  59985=>"110110000",
  59986=>"101111100",
  59987=>"010011101",
  59988=>"011010101",
  59989=>"100001010",
  59990=>"111001101",
  59991=>"111000001",
  59992=>"001010100",
  59993=>"001001001",
  59994=>"101011000",
  59995=>"001011000",
  59996=>"000101000",
  59997=>"010111110",
  59998=>"101011001",
  59999=>"111111110",
  60000=>"000111100",
  60001=>"000110001",
  60002=>"101010010",
  60003=>"000110101",
  60004=>"100110101",
  60005=>"101101100",
  60006=>"010110111",
  60007=>"001001010",
  60008=>"001010101",
  60009=>"101110100",
  60010=>"011100100",
  60011=>"000111110",
  60012=>"101101100",
  60013=>"100100001",
  60014=>"001111101",
  60015=>"001000010",
  60016=>"000010011",
  60017=>"000100101",
  60018=>"110001111",
  60019=>"001001111",
  60020=>"000000000",
  60021=>"010110010",
  60022=>"110010100",
  60023=>"111001101",
  60024=>"001001101",
  60025=>"100001000",
  60026=>"001110000",
  60027=>"001100110",
  60028=>"001000100",
  60029=>"111010110",
  60030=>"000101000",
  60031=>"111100101",
  60032=>"111011010",
  60033=>"001011100",
  60034=>"010101000",
  60035=>"110010011",
  60036=>"111001111",
  60037=>"100110100",
  60038=>"111111000",
  60039=>"110100000",
  60040=>"111010100",
  60041=>"101001100",
  60042=>"000111101",
  60043=>"111001110",
  60044=>"011010000",
  60045=>"101001001",
  60046=>"011111110",
  60047=>"010101111",
  60048=>"101011100",
  60049=>"010010010",
  60050=>"101111100",
  60051=>"111111111",
  60052=>"001001110",
  60053=>"010010111",
  60054=>"110011100",
  60055=>"100111100",
  60056=>"000100101",
  60057=>"101000001",
  60058=>"001000010",
  60059=>"011111111",
  60060=>"001011110",
  60061=>"001101111",
  60062=>"010100111",
  60063=>"010111000",
  60064=>"000000100",
  60065=>"111101001",
  60066=>"100100000",
  60067=>"110010111",
  60068=>"111011101",
  60069=>"010100001",
  60070=>"001000101",
  60071=>"111010100",
  60072=>"000010001",
  60073=>"001111011",
  60074=>"100110100",
  60075=>"010000111",
  60076=>"110000001",
  60077=>"011111001",
  60078=>"101101100",
  60079=>"101111110",
  60080=>"011011110",
  60081=>"011001011",
  60082=>"100001010",
  60083=>"111011110",
  60084=>"111101100",
  60085=>"111010110",
  60086=>"010011001",
  60087=>"101110110",
  60088=>"100111100",
  60089=>"110011001",
  60090=>"011101000",
  60091=>"100010010",
  60092=>"110011011",
  60093=>"110101000",
  60094=>"000101111",
  60095=>"111110110",
  60096=>"111111000",
  60097=>"010011100",
  60098=>"011110001",
  60099=>"000100100",
  60100=>"000100100",
  60101=>"100100001",
  60102=>"110001111",
  60103=>"010000010",
  60104=>"000100010",
  60105=>"001011001",
  60106=>"111111011",
  60107=>"001110011",
  60108=>"011111111",
  60109=>"001000100",
  60110=>"101000100",
  60111=>"001011000",
  60112=>"010100000",
  60113=>"101111110",
  60114=>"110001000",
  60115=>"110000010",
  60116=>"101011100",
  60117=>"000100000",
  60118=>"100000100",
  60119=>"100101010",
  60120=>"000001110",
  60121=>"010011111",
  60122=>"001100111",
  60123=>"010111011",
  60124=>"010010101",
  60125=>"010001011",
  60126=>"110000110",
  60127=>"011100011",
  60128=>"001011111",
  60129=>"101110000",
  60130=>"010010010",
  60131=>"011100101",
  60132=>"001011111",
  60133=>"000111101",
  60134=>"100001001",
  60135=>"010001101",
  60136=>"100111100",
  60137=>"101000001",
  60138=>"010001000",
  60139=>"001110101",
  60140=>"000110010",
  60141=>"110101101",
  60142=>"111110011",
  60143=>"000000011",
  60144=>"110010001",
  60145=>"111100100",
  60146=>"110001101",
  60147=>"111110101",
  60148=>"000110010",
  60149=>"001111101",
  60150=>"011011101",
  60151=>"110101110",
  60152=>"110100010",
  60153=>"111100101",
  60154=>"010001100",
  60155=>"001100110",
  60156=>"000011111",
  60157=>"000001010",
  60158=>"010001101",
  60159=>"010100110",
  60160=>"101110010",
  60161=>"100011011",
  60162=>"011111010",
  60163=>"111000000",
  60164=>"000100101",
  60165=>"010010111",
  60166=>"101111000",
  60167=>"001110100",
  60168=>"101110010",
  60169=>"010000110",
  60170=>"100011111",
  60171=>"101000011",
  60172=>"010110100",
  60173=>"010001100",
  60174=>"100000010",
  60175=>"011001111",
  60176=>"111011000",
  60177=>"000111111",
  60178=>"101010010",
  60179=>"100010010",
  60180=>"101111001",
  60181=>"000111110",
  60182=>"111011100",
  60183=>"100001100",
  60184=>"000100001",
  60185=>"100110001",
  60186=>"100000011",
  60187=>"001011100",
  60188=>"111101011",
  60189=>"001000010",
  60190=>"101000000",
  60191=>"101110000",
  60192=>"010111101",
  60193=>"001010001",
  60194=>"100000010",
  60195=>"011100010",
  60196=>"111111010",
  60197=>"100011010",
  60198=>"011001011",
  60199=>"000111111",
  60200=>"001111001",
  60201=>"111110001",
  60202=>"101011101",
  60203=>"111000110",
  60204=>"100000111",
  60205=>"011101010",
  60206=>"010000000",
  60207=>"101110000",
  60208=>"010101110",
  60209=>"101001000",
  60210=>"100011010",
  60211=>"011011111",
  60212=>"001001000",
  60213=>"110011110",
  60214=>"001111001",
  60215=>"110001100",
  60216=>"000100000",
  60217=>"110011000",
  60218=>"110111101",
  60219=>"100111110",
  60220=>"010011011",
  60221=>"000110001",
  60222=>"101101001",
  60223=>"100010000",
  60224=>"001110010",
  60225=>"011111111",
  60226=>"110011110",
  60227=>"100110111",
  60228=>"110010111",
  60229=>"001010010",
  60230=>"011100000",
  60231=>"001001101",
  60232=>"110001010",
  60233=>"100101100",
  60234=>"000010011",
  60235=>"101110110",
  60236=>"010100000",
  60237=>"111101000",
  60238=>"111000111",
  60239=>"001010111",
  60240=>"110001100",
  60241=>"110101100",
  60242=>"111110000",
  60243=>"111110011",
  60244=>"110100110",
  60245=>"111111111",
  60246=>"100010101",
  60247=>"010110100",
  60248=>"010011001",
  60249=>"111111110",
  60250=>"111011110",
  60251=>"110100001",
  60252=>"000100111",
  60253=>"101111111",
  60254=>"001111110",
  60255=>"000000111",
  60256=>"110110110",
  60257=>"001111001",
  60258=>"000010000",
  60259=>"000110001",
  60260=>"100001100",
  60261=>"000110011",
  60262=>"110011010",
  60263=>"111010111",
  60264=>"001111110",
  60265=>"010111010",
  60266=>"101111101",
  60267=>"101111001",
  60268=>"110100111",
  60269=>"000010011",
  60270=>"100010000",
  60271=>"001101011",
  60272=>"011101111",
  60273=>"010010000",
  60274=>"101101101",
  60275=>"001101101",
  60276=>"100000001",
  60277=>"001110010",
  60278=>"000011110",
  60279=>"000010111",
  60280=>"001110100",
  60281=>"110011111",
  60282=>"010101111",
  60283=>"001111110",
  60284=>"000100001",
  60285=>"100010100",
  60286=>"101000101",
  60287=>"000111001",
  60288=>"000000001",
  60289=>"100110110",
  60290=>"000111000",
  60291=>"000111010",
  60292=>"000010010",
  60293=>"101100000",
  60294=>"111010011",
  60295=>"111001001",
  60296=>"110111110",
  60297=>"011110010",
  60298=>"101101000",
  60299=>"011111100",
  60300=>"110101011",
  60301=>"011110000",
  60302=>"001001000",
  60303=>"110000000",
  60304=>"001001100",
  60305=>"001011010",
  60306=>"110110010",
  60307=>"101101000",
  60308=>"001100010",
  60309=>"111101100",
  60310=>"110000101",
  60311=>"111000011",
  60312=>"111010001",
  60313=>"110010001",
  60314=>"100010010",
  60315=>"100001100",
  60316=>"111011110",
  60317=>"101001000",
  60318=>"110101001",
  60319=>"000111111",
  60320=>"000001011",
  60321=>"110101001",
  60322=>"100000110",
  60323=>"111000000",
  60324=>"000100110",
  60325=>"000011000",
  60326=>"101111100",
  60327=>"001010111",
  60328=>"110111000",
  60329=>"000010000",
  60330=>"110011011",
  60331=>"100001101",
  60332=>"000011100",
  60333=>"010110001",
  60334=>"001100101",
  60335=>"111010100",
  60336=>"010100111",
  60337=>"010111111",
  60338=>"100001001",
  60339=>"011111011",
  60340=>"011011011",
  60341=>"000001010",
  60342=>"010101111",
  60343=>"111101010",
  60344=>"000101011",
  60345=>"010011000",
  60346=>"001001010",
  60347=>"111010010",
  60348=>"111101100",
  60349=>"111100100",
  60350=>"110001101",
  60351=>"000000100",
  60352=>"001011011",
  60353=>"110010010",
  60354=>"011011110",
  60355=>"110110110",
  60356=>"110110010",
  60357=>"110111011",
  60358=>"110110100",
  60359=>"010110001",
  60360=>"010011100",
  60361=>"101000111",
  60362=>"110100101",
  60363=>"000111111",
  60364=>"010101001",
  60365=>"000010101",
  60366=>"101101001",
  60367=>"111110110",
  60368=>"001111010",
  60369=>"110001101",
  60370=>"101110000",
  60371=>"010000011",
  60372=>"001010111",
  60373=>"000001010",
  60374=>"110000100",
  60375=>"101110101",
  60376=>"011111011",
  60377=>"001000101",
  60378=>"001100111",
  60379=>"111011110",
  60380=>"110110000",
  60381=>"111101010",
  60382=>"101111000",
  60383=>"001111101",
  60384=>"010101111",
  60385=>"111101111",
  60386=>"001110111",
  60387=>"000011011",
  60388=>"010100000",
  60389=>"110001001",
  60390=>"010001011",
  60391=>"001100001",
  60392=>"001011000",
  60393=>"110100001",
  60394=>"110111111",
  60395=>"101110000",
  60396=>"000100000",
  60397=>"101000011",
  60398=>"100100111",
  60399=>"000000111",
  60400=>"101010110",
  60401=>"100101010",
  60402=>"010010000",
  60403=>"111111100",
  60404=>"100110010",
  60405=>"100011011",
  60406=>"101000011",
  60407=>"000000000",
  60408=>"001100001",
  60409=>"001010110",
  60410=>"000001101",
  60411=>"011001011",
  60412=>"000010011",
  60413=>"000011111",
  60414=>"000011100",
  60415=>"101101100",
  60416=>"010011110",
  60417=>"000011010",
  60418=>"010011111",
  60419=>"101010010",
  60420=>"101111111",
  60421=>"000000100",
  60422=>"101000001",
  60423=>"101011111",
  60424=>"111011001",
  60425=>"111011101",
  60426=>"011010100",
  60427=>"111000110",
  60428=>"111001100",
  60429=>"110010111",
  60430=>"101101100",
  60431=>"111101110",
  60432=>"011100111",
  60433=>"100110100",
  60434=>"000010000",
  60435=>"111100111",
  60436=>"111111100",
  60437=>"111100001",
  60438=>"010000000",
  60439=>"111010110",
  60440=>"000100010",
  60441=>"000000011",
  60442=>"001011101",
  60443=>"011001010",
  60444=>"001011010",
  60445=>"000111110",
  60446=>"101001111",
  60447=>"111000011",
  60448=>"001100000",
  60449=>"011100100",
  60450=>"010001010",
  60451=>"000010111",
  60452=>"001101011",
  60453=>"001100101",
  60454=>"101010011",
  60455=>"111111001",
  60456=>"110011011",
  60457=>"100101000",
  60458=>"011000100",
  60459=>"110010001",
  60460=>"000111101",
  60461=>"001010011",
  60462=>"000010111",
  60463=>"100100000",
  60464=>"000101010",
  60465=>"111000110",
  60466=>"110110111",
  60467=>"011011100",
  60468=>"100101110",
  60469=>"000011011",
  60470=>"110000010",
  60471=>"001000000",
  60472=>"110110100",
  60473=>"101010100",
  60474=>"100001101",
  60475=>"010001000",
  60476=>"001111001",
  60477=>"010111100",
  60478=>"110110100",
  60479=>"101001101",
  60480=>"101011011",
  60481=>"001001111",
  60482=>"111000100",
  60483=>"010011001",
  60484=>"010111100",
  60485=>"110001011",
  60486=>"100010101",
  60487=>"101111110",
  60488=>"100011000",
  60489=>"100111101",
  60490=>"101110000",
  60491=>"001010000",
  60492=>"100101010",
  60493=>"011110100",
  60494=>"010101001",
  60495=>"011111101",
  60496=>"101000000",
  60497=>"000010101",
  60498=>"001111000",
  60499=>"100111011",
  60500=>"111001100",
  60501=>"001110101",
  60502=>"110010000",
  60503=>"100100111",
  60504=>"111101100",
  60505=>"111110111",
  60506=>"000010011",
  60507=>"111101111",
  60508=>"001101110",
  60509=>"100110010",
  60510=>"001000110",
  60511=>"000110111",
  60512=>"000111010",
  60513=>"110100101",
  60514=>"110000001",
  60515=>"100111111",
  60516=>"010100100",
  60517=>"101110011",
  60518=>"100110011",
  60519=>"111111001",
  60520=>"110010110",
  60521=>"000110110",
  60522=>"101000011",
  60523=>"001100110",
  60524=>"110110110",
  60525=>"001000101",
  60526=>"011111000",
  60527=>"010000100",
  60528=>"000101010",
  60529=>"101100001",
  60530=>"010000101",
  60531=>"011111101",
  60532=>"000100000",
  60533=>"010110001",
  60534=>"000100111",
  60535=>"111101110",
  60536=>"101100100",
  60537=>"011111010",
  60538=>"100101111",
  60539=>"101011100",
  60540=>"000000000",
  60541=>"101100111",
  60542=>"101101000",
  60543=>"100000111",
  60544=>"110010001",
  60545=>"111001011",
  60546=>"111111110",
  60547=>"001011010",
  60548=>"001010001",
  60549=>"000001011",
  60550=>"010111000",
  60551=>"001010000",
  60552=>"000101010",
  60553=>"110001111",
  60554=>"111100001",
  60555=>"000111011",
  60556=>"110111100",
  60557=>"111000001",
  60558=>"110000100",
  60559=>"000000000",
  60560=>"000010101",
  60561=>"110000011",
  60562=>"100010101",
  60563=>"001001011",
  60564=>"111000111",
  60565=>"100000010",
  60566=>"100000001",
  60567=>"101111000",
  60568=>"111110000",
  60569=>"111000111",
  60570=>"000000110",
  60571=>"010010000",
  60572=>"010101110",
  60573=>"100010110",
  60574=>"000001101",
  60575=>"010000000",
  60576=>"111010001",
  60577=>"001110101",
  60578=>"000110111",
  60579=>"101000000",
  60580=>"001010001",
  60581=>"001010000",
  60582=>"000101001",
  60583=>"111011110",
  60584=>"101111011",
  60585=>"101000000",
  60586=>"111000100",
  60587=>"001100111",
  60588=>"011111110",
  60589=>"001110110",
  60590=>"011100000",
  60591=>"011001001",
  60592=>"010000010",
  60593=>"000100110",
  60594=>"100000100",
  60595=>"010010101",
  60596=>"010111000",
  60597=>"000010111",
  60598=>"010111111",
  60599=>"110001110",
  60600=>"011101111",
  60601=>"001110111",
  60602=>"110101110",
  60603=>"111001101",
  60604=>"100001100",
  60605=>"011000101",
  60606=>"100110111",
  60607=>"111101110",
  60608=>"110100111",
  60609=>"010110110",
  60610=>"110101010",
  60611=>"010011011",
  60612=>"111011010",
  60613=>"000101110",
  60614=>"000100101",
  60615=>"010001011",
  60616=>"010111001",
  60617=>"001011000",
  60618=>"101101010",
  60619=>"001111000",
  60620=>"111101001",
  60621=>"001101110",
  60622=>"101100111",
  60623=>"010110000",
  60624=>"001110011",
  60625=>"100110000",
  60626=>"110110100",
  60627=>"011110111",
  60628=>"100010001",
  60629=>"110101011",
  60630=>"010101011",
  60631=>"100001110",
  60632=>"011001000",
  60633=>"001111001",
  60634=>"111101011",
  60635=>"000010001",
  60636=>"110111110",
  60637=>"110111011",
  60638=>"110111001",
  60639=>"010010110",
  60640=>"010100100",
  60641=>"101101011",
  60642=>"001101000",
  60643=>"100001000",
  60644=>"100101010",
  60645=>"111011001",
  60646=>"000001100",
  60647=>"010001011",
  60648=>"010010100",
  60649=>"111010000",
  60650=>"000010000",
  60651=>"011111001",
  60652=>"110101010",
  60653=>"001100000",
  60654=>"000000001",
  60655=>"001101100",
  60656=>"111011100",
  60657=>"111011101",
  60658=>"011111100",
  60659=>"000011011",
  60660=>"100001111",
  60661=>"010000101",
  60662=>"110001100",
  60663=>"000011010",
  60664=>"111011111",
  60665=>"111100010",
  60666=>"100011000",
  60667=>"000111000",
  60668=>"011111000",
  60669=>"101000000",
  60670=>"010001110",
  60671=>"001001011",
  60672=>"100011101",
  60673=>"010011100",
  60674=>"011111001",
  60675=>"000101101",
  60676=>"001010010",
  60677=>"100111000",
  60678=>"100011110",
  60679=>"111000111",
  60680=>"111010001",
  60681=>"010111011",
  60682=>"011000000",
  60683=>"000100110",
  60684=>"111110111",
  60685=>"010000110",
  60686=>"010111010",
  60687=>"111010101",
  60688=>"110100110",
  60689=>"111011111",
  60690=>"111110111",
  60691=>"110100001",
  60692=>"110111101",
  60693=>"000000101",
  60694=>"000101111",
  60695=>"100000100",
  60696=>"101011011",
  60697=>"010110010",
  60698=>"000000010",
  60699=>"100001110",
  60700=>"110100101",
  60701=>"101000001",
  60702=>"111001100",
  60703=>"101001111",
  60704=>"000000111",
  60705=>"111110001",
  60706=>"111001101",
  60707=>"010001010",
  60708=>"011001100",
  60709=>"001100011",
  60710=>"001010100",
  60711=>"100011011",
  60712=>"011100011",
  60713=>"100001101",
  60714=>"101000101",
  60715=>"011100100",
  60716=>"010010000",
  60717=>"011111110",
  60718=>"100000001",
  60719=>"100010011",
  60720=>"001111110",
  60721=>"110011110",
  60722=>"011001010",
  60723=>"110101011",
  60724=>"001000101",
  60725=>"000001000",
  60726=>"110000110",
  60727=>"001000110",
  60728=>"011111100",
  60729=>"110000101",
  60730=>"111101111",
  60731=>"001101001",
  60732=>"110011111",
  60733=>"111000001",
  60734=>"100001010",
  60735=>"000000000",
  60736=>"100100101",
  60737=>"000011110",
  60738=>"011100100",
  60739=>"100001010",
  60740=>"100101010",
  60741=>"100110100",
  60742=>"100001000",
  60743=>"010100001",
  60744=>"110001000",
  60745=>"111110100",
  60746=>"000110111",
  60747=>"111010001",
  60748=>"011010011",
  60749=>"001100001",
  60750=>"111111101",
  60751=>"111010100",
  60752=>"001111000",
  60753=>"011000110",
  60754=>"101010010",
  60755=>"110111000",
  60756=>"001110001",
  60757=>"111111111",
  60758=>"000010011",
  60759=>"100101001",
  60760=>"111001110",
  60761=>"111010010",
  60762=>"101101000",
  60763=>"000100010",
  60764=>"110101100",
  60765=>"010000100",
  60766=>"111000101",
  60767=>"110001001",
  60768=>"000000101",
  60769=>"000111000",
  60770=>"110000011",
  60771=>"101101011",
  60772=>"010000100",
  60773=>"010100001",
  60774=>"000100101",
  60775=>"001010001",
  60776=>"110101010",
  60777=>"010100001",
  60778=>"111111000",
  60779=>"010100001",
  60780=>"001001001",
  60781=>"111111100",
  60782=>"110011110",
  60783=>"011011110",
  60784=>"000110010",
  60785=>"101000110",
  60786=>"001111011",
  60787=>"011011100",
  60788=>"110011111",
  60789=>"001000001",
  60790=>"000111101",
  60791=>"101000010",
  60792=>"001011000",
  60793=>"011100001",
  60794=>"001101101",
  60795=>"100100101",
  60796=>"000101001",
  60797=>"111110011",
  60798=>"100101111",
  60799=>"000000011",
  60800=>"000010001",
  60801=>"011011011",
  60802=>"101011001",
  60803=>"111111011",
  60804=>"000001101",
  60805=>"111001010",
  60806=>"101110011",
  60807=>"011111010",
  60808=>"001100001",
  60809=>"010111001",
  60810=>"001000001",
  60811=>"100000000",
  60812=>"101010111",
  60813=>"001000000",
  60814=>"000001110",
  60815=>"100111001",
  60816=>"110000001",
  60817=>"000101000",
  60818=>"110101000",
  60819=>"100100100",
  60820=>"111000010",
  60821=>"111000001",
  60822=>"110111111",
  60823=>"110001110",
  60824=>"001101100",
  60825=>"111111100",
  60826=>"111110111",
  60827=>"101110110",
  60828=>"010101110",
  60829=>"110000101",
  60830=>"010000101",
  60831=>"101100011",
  60832=>"100101010",
  60833=>"010000110",
  60834=>"101101101",
  60835=>"010101110",
  60836=>"010001111",
  60837=>"100000101",
  60838=>"100100001",
  60839=>"110000011",
  60840=>"000111000",
  60841=>"100111101",
  60842=>"100000000",
  60843=>"010011111",
  60844=>"101010101",
  60845=>"011010001",
  60846=>"100101011",
  60847=>"011111111",
  60848=>"111011011",
  60849=>"101010000",
  60850=>"000100111",
  60851=>"100101100",
  60852=>"000101001",
  60853=>"001011001",
  60854=>"101010100",
  60855=>"011110000",
  60856=>"001001101",
  60857=>"111001000",
  60858=>"011101010",
  60859=>"001101011",
  60860=>"010101101",
  60861=>"011111101",
  60862=>"011001001",
  60863=>"110101100",
  60864=>"011100100",
  60865=>"011000110",
  60866=>"010000010",
  60867=>"110100000",
  60868=>"000110110",
  60869=>"101001100",
  60870=>"010001111",
  60871=>"100100001",
  60872=>"000000001",
  60873=>"011101100",
  60874=>"000011011",
  60875=>"111110001",
  60876=>"111011000",
  60877=>"000001110",
  60878=>"111010010",
  60879=>"010011011",
  60880=>"101001100",
  60881=>"111111101",
  60882=>"101011001",
  60883=>"111111001",
  60884=>"100110001",
  60885=>"010010010",
  60886=>"000001011",
  60887=>"001100001",
  60888=>"000000010",
  60889=>"110010110",
  60890=>"000100101",
  60891=>"000110101",
  60892=>"010011011",
  60893=>"000111111",
  60894=>"001100000",
  60895=>"100001111",
  60896=>"011001110",
  60897=>"001110101",
  60898=>"111100010",
  60899=>"000101001",
  60900=>"101110101",
  60901=>"100011010",
  60902=>"000100111",
  60903=>"011001100",
  60904=>"100110100",
  60905=>"100010001",
  60906=>"010000011",
  60907=>"100001100",
  60908=>"110000001",
  60909=>"101011001",
  60910=>"100101010",
  60911=>"110111110",
  60912=>"000110111",
  60913=>"000001100",
  60914=>"110111011",
  60915=>"011111011",
  60916=>"000000111",
  60917=>"001001100",
  60918=>"000001010",
  60919=>"101001100",
  60920=>"111000000",
  60921=>"111001010",
  60922=>"100000111",
  60923=>"000001000",
  60924=>"111010111",
  60925=>"010111000",
  60926=>"111001010",
  60927=>"001010111",
  60928=>"000110000",
  60929=>"010111010",
  60930=>"010001111",
  60931=>"000101010",
  60932=>"001110000",
  60933=>"001101100",
  60934=>"000101101",
  60935=>"011111011",
  60936=>"001000000",
  60937=>"101110101",
  60938=>"001010100",
  60939=>"111001110",
  60940=>"101011001",
  60941=>"000010110",
  60942=>"000100000",
  60943=>"111001111",
  60944=>"101001000",
  60945=>"100110010",
  60946=>"001010001",
  60947=>"010110011",
  60948=>"000101011",
  60949=>"000010000",
  60950=>"100000001",
  60951=>"111101011",
  60952=>"111110101",
  60953=>"001110000",
  60954=>"000110110",
  60955=>"011010000",
  60956=>"011000010",
  60957=>"010001000",
  60958=>"001111100",
  60959=>"000100011",
  60960=>"111110011",
  60961=>"110000001",
  60962=>"000111101",
  60963=>"000000010",
  60964=>"111011101",
  60965=>"010010001",
  60966=>"001010010",
  60967=>"111101011",
  60968=>"111111011",
  60969=>"110000110",
  60970=>"000001000",
  60971=>"101001001",
  60972=>"000110101",
  60973=>"100100111",
  60974=>"000101110",
  60975=>"000100000",
  60976=>"000000000",
  60977=>"111000101",
  60978=>"001111010",
  60979=>"100110011",
  60980=>"101011010",
  60981=>"000011111",
  60982=>"111001001",
  60983=>"110101000",
  60984=>"001010100",
  60985=>"101010011",
  60986=>"100000111",
  60987=>"010111101",
  60988=>"111011111",
  60989=>"110111101",
  60990=>"001000000",
  60991=>"111011010",
  60992=>"110101111",
  60993=>"100100011",
  60994=>"110111110",
  60995=>"110101110",
  60996=>"111010010",
  60997=>"100110010",
  60998=>"101010001",
  60999=>"011001011",
  61000=>"111111000",
  61001=>"111100011",
  61002=>"100101101",
  61003=>"000011110",
  61004=>"011000001",
  61005=>"000101110",
  61006=>"111001011",
  61007=>"000110101",
  61008=>"101100001",
  61009=>"100000101",
  61010=>"110001101",
  61011=>"001000011",
  61012=>"011110010",
  61013=>"011101010",
  61014=>"111101101",
  61015=>"100110001",
  61016=>"110010110",
  61017=>"110110000",
  61018=>"111100111",
  61019=>"100111110",
  61020=>"010101101",
  61021=>"100000110",
  61022=>"111111100",
  61023=>"101000011",
  61024=>"011000010",
  61025=>"001100000",
  61026=>"001011110",
  61027=>"000111110",
  61028=>"110101110",
  61029=>"010010111",
  61030=>"011110111",
  61031=>"000100111",
  61032=>"000000000",
  61033=>"100111000",
  61034=>"111000110",
  61035=>"101011011",
  61036=>"100001010",
  61037=>"111001011",
  61038=>"000011100",
  61039=>"010001000",
  61040=>"001000111",
  61041=>"000110010",
  61042=>"000100011",
  61043=>"110101100",
  61044=>"001110111",
  61045=>"010001100",
  61046=>"111101110",
  61047=>"111111010",
  61048=>"011110001",
  61049=>"101010100",
  61050=>"111100010",
  61051=>"000001001",
  61052=>"000100001",
  61053=>"101100101",
  61054=>"001011010",
  61055=>"010100100",
  61056=>"111110010",
  61057=>"101101010",
  61058=>"001000000",
  61059=>"011111100",
  61060=>"011001100",
  61061=>"101001000",
  61062=>"110001111",
  61063=>"001111100",
  61064=>"010111010",
  61065=>"011001011",
  61066=>"010101111",
  61067=>"001111000",
  61068=>"011010001",
  61069=>"111000000",
  61070=>"000010110",
  61071=>"111110100",
  61072=>"000110010",
  61073=>"000111110",
  61074=>"001010111",
  61075=>"010010111",
  61076=>"000011110",
  61077=>"011010101",
  61078=>"001001011",
  61079=>"000001110",
  61080=>"110011001",
  61081=>"001000010",
  61082=>"111000000",
  61083=>"000111011",
  61084=>"111101101",
  61085=>"100000100",
  61086=>"011101111",
  61087=>"110011101",
  61088=>"000111111",
  61089=>"010010000",
  61090=>"001011010",
  61091=>"010001110",
  61092=>"010010101",
  61093=>"100011101",
  61094=>"100110011",
  61095=>"000111101",
  61096=>"111110010",
  61097=>"110101010",
  61098=>"000101011",
  61099=>"000100011",
  61100=>"100110000",
  61101=>"100001010",
  61102=>"001101011",
  61103=>"110000010",
  61104=>"011110010",
  61105=>"100101111",
  61106=>"011100110",
  61107=>"011101101",
  61108=>"110100110",
  61109=>"000010101",
  61110=>"100000010",
  61111=>"101001111",
  61112=>"111000101",
  61113=>"010100001",
  61114=>"000101011",
  61115=>"000000101",
  61116=>"010011011",
  61117=>"010101010",
  61118=>"000111010",
  61119=>"000110111",
  61120=>"111110100",
  61121=>"100000100",
  61122=>"001101000",
  61123=>"001010101",
  61124=>"011000101",
  61125=>"111000001",
  61126=>"101001111",
  61127=>"101101010",
  61128=>"100000001",
  61129=>"101000110",
  61130=>"110110100",
  61131=>"010110101",
  61132=>"000111010",
  61133=>"111000010",
  61134=>"000010001",
  61135=>"100000100",
  61136=>"001011111",
  61137=>"101100010",
  61138=>"011111100",
  61139=>"011101111",
  61140=>"100100111",
  61141=>"000010001",
  61142=>"101101010",
  61143=>"000110010",
  61144=>"110101011",
  61145=>"001011011",
  61146=>"000011101",
  61147=>"111110100",
  61148=>"011110010",
  61149=>"000001100",
  61150=>"001100011",
  61151=>"001110010",
  61152=>"100000110",
  61153=>"101001101",
  61154=>"000001000",
  61155=>"010101110",
  61156=>"110111110",
  61157=>"010111010",
  61158=>"110001010",
  61159=>"001111100",
  61160=>"011101100",
  61161=>"100110100",
  61162=>"011010011",
  61163=>"010000010",
  61164=>"111001010",
  61165=>"011110000",
  61166=>"110011100",
  61167=>"000100010",
  61168=>"110001111",
  61169=>"000011101",
  61170=>"010001000",
  61171=>"000110000",
  61172=>"010100110",
  61173=>"111100111",
  61174=>"001110100",
  61175=>"110011010",
  61176=>"111000111",
  61177=>"011110010",
  61178=>"110111101",
  61179=>"100100000",
  61180=>"011110110",
  61181=>"100110111",
  61182=>"101110000",
  61183=>"001101101",
  61184=>"111011100",
  61185=>"101111111",
  61186=>"101001111",
  61187=>"001001010",
  61188=>"100000110",
  61189=>"101000000",
  61190=>"100001010",
  61191=>"101100000",
  61192=>"000010000",
  61193=>"100101000",
  61194=>"011010000",
  61195=>"000000110",
  61196=>"111001111",
  61197=>"000101100",
  61198=>"010011000",
  61199=>"110011101",
  61200=>"010000111",
  61201=>"100101000",
  61202=>"101010000",
  61203=>"000000011",
  61204=>"010000000",
  61205=>"010110010",
  61206=>"010101000",
  61207=>"010001100",
  61208=>"111100001",
  61209=>"111100001",
  61210=>"101001010",
  61211=>"101011101",
  61212=>"111100011",
  61213=>"001100100",
  61214=>"110011110",
  61215=>"100011111",
  61216=>"001000000",
  61217=>"011110001",
  61218=>"010101111",
  61219=>"110101001",
  61220=>"011101111",
  61221=>"101101000",
  61222=>"100111110",
  61223=>"110000100",
  61224=>"000000011",
  61225=>"101101101",
  61226=>"100100011",
  61227=>"100110110",
  61228=>"110010000",
  61229=>"000101111",
  61230=>"000010110",
  61231=>"001101110",
  61232=>"011111111",
  61233=>"011100000",
  61234=>"101011101",
  61235=>"000100111",
  61236=>"100101000",
  61237=>"110110010",
  61238=>"111000111",
  61239=>"110101011",
  61240=>"010001001",
  61241=>"101010001",
  61242=>"010001000",
  61243=>"110111011",
  61244=>"000110000",
  61245=>"101000101",
  61246=>"010111101",
  61247=>"100100100",
  61248=>"011100100",
  61249=>"001100000",
  61250=>"001010001",
  61251=>"110011100",
  61252=>"001101110",
  61253=>"100101111",
  61254=>"010001000",
  61255=>"001011111",
  61256=>"011001001",
  61257=>"110000000",
  61258=>"111000110",
  61259=>"001100001",
  61260=>"001111011",
  61261=>"110001010",
  61262=>"011010011",
  61263=>"001000100",
  61264=>"011000111",
  61265=>"010111001",
  61266=>"000011010",
  61267=>"011100100",
  61268=>"000101011",
  61269=>"001011111",
  61270=>"000000000",
  61271=>"000110111",
  61272=>"110001100",
  61273=>"111101001",
  61274=>"001000011",
  61275=>"000101110",
  61276=>"001101001",
  61277=>"001001100",
  61278=>"100011010",
  61279=>"000011110",
  61280=>"011010100",
  61281=>"110101110",
  61282=>"100000110",
  61283=>"111111001",
  61284=>"010110111",
  61285=>"100000000",
  61286=>"001010100",
  61287=>"010110010",
  61288=>"001100001",
  61289=>"110000000",
  61290=>"101100010",
  61291=>"011000100",
  61292=>"001111111",
  61293=>"110100100",
  61294=>"100100110",
  61295=>"111011010",
  61296=>"000010001",
  61297=>"001000010",
  61298=>"100000110",
  61299=>"101000111",
  61300=>"010101111",
  61301=>"101111111",
  61302=>"001011010",
  61303=>"110010001",
  61304=>"000000110",
  61305=>"011011100",
  61306=>"110100001",
  61307=>"110101001",
  61308=>"101010110",
  61309=>"011100011",
  61310=>"001000011",
  61311=>"110111010",
  61312=>"000011111",
  61313=>"001010010",
  61314=>"101111110",
  61315=>"011100100",
  61316=>"101010000",
  61317=>"101111101",
  61318=>"000110000",
  61319=>"100111111",
  61320=>"011101001",
  61321=>"010100001",
  61322=>"000000110",
  61323=>"000000100",
  61324=>"010011010",
  61325=>"110111111",
  61326=>"100110010",
  61327=>"010101011",
  61328=>"100110001",
  61329=>"011110110",
  61330=>"010001010",
  61331=>"101100101",
  61332=>"101101000",
  61333=>"010101110",
  61334=>"001010000",
  61335=>"000000011",
  61336=>"111001010",
  61337=>"001001011",
  61338=>"000111111",
  61339=>"110110000",
  61340=>"010010101",
  61341=>"111101010",
  61342=>"100000111",
  61343=>"110011111",
  61344=>"010111111",
  61345=>"101011001",
  61346=>"001000001",
  61347=>"001101001",
  61348=>"111101001",
  61349=>"100110100",
  61350=>"001011110",
  61351=>"110111000",
  61352=>"000101001",
  61353=>"111010101",
  61354=>"110110100",
  61355=>"111110110",
  61356=>"111011110",
  61357=>"111111100",
  61358=>"010000000",
  61359=>"001111001",
  61360=>"110111000",
  61361=>"100100111",
  61362=>"101011011",
  61363=>"001010100",
  61364=>"011100101",
  61365=>"111110111",
  61366=>"010110100",
  61367=>"001110101",
  61368=>"101100011",
  61369=>"001000111",
  61370=>"100110100",
  61371=>"010111111",
  61372=>"111101001",
  61373=>"011000101",
  61374=>"101001101",
  61375=>"010000101",
  61376=>"101010011",
  61377=>"001100110",
  61378=>"110000100",
  61379=>"101111100",
  61380=>"000010011",
  61381=>"000100001",
  61382=>"010001001",
  61383=>"110111100",
  61384=>"100010101",
  61385=>"010110000",
  61386=>"010001000",
  61387=>"101011001",
  61388=>"000100111",
  61389=>"000000011",
  61390=>"101100100",
  61391=>"010010001",
  61392=>"001100011",
  61393=>"111101101",
  61394=>"001011111",
  61395=>"000011101",
  61396=>"100010111",
  61397=>"010110101",
  61398=>"011000100",
  61399=>"000111000",
  61400=>"001100100",
  61401=>"010000001",
  61402=>"110110010",
  61403=>"100000111",
  61404=>"000111000",
  61405=>"110100100",
  61406=>"100110000",
  61407=>"101001101",
  61408=>"110101010",
  61409=>"000100100",
  61410=>"000000110",
  61411=>"101100111",
  61412=>"001010001",
  61413=>"101110110",
  61414=>"101000000",
  61415=>"110010001",
  61416=>"000010111",
  61417=>"101000111",
  61418=>"001110100",
  61419=>"000111011",
  61420=>"110011011",
  61421=>"011001110",
  61422=>"011110111",
  61423=>"111111110",
  61424=>"000000100",
  61425=>"000001011",
  61426=>"010100111",
  61427=>"011101000",
  61428=>"011101011",
  61429=>"101010101",
  61430=>"011010010",
  61431=>"100000101",
  61432=>"000001110",
  61433=>"110111011",
  61434=>"010010101",
  61435=>"111100000",
  61436=>"101010000",
  61437=>"111011001",
  61438=>"101001001",
  61439=>"000101110",
  61440=>"110110110",
  61441=>"101001010",
  61442=>"110101100",
  61443=>"011101010",
  61444=>"110101010",
  61445=>"111001100",
  61446=>"110101010",
  61447=>"001111111",
  61448=>"010011010",
  61449=>"101011101",
  61450=>"011000011",
  61451=>"100101110",
  61452=>"011011011",
  61453=>"001001011",
  61454=>"010110001",
  61455=>"101010110",
  61456=>"101010110",
  61457=>"010010111",
  61458=>"010010110",
  61459=>"011000101",
  61460=>"000110110",
  61461=>"100111011",
  61462=>"001010011",
  61463=>"110111001",
  61464=>"001100110",
  61465=>"101100000",
  61466=>"111001101",
  61467=>"110100010",
  61468=>"110101110",
  61469=>"000011010",
  61470=>"010101001",
  61471=>"001101001",
  61472=>"111101011",
  61473=>"110000100",
  61474=>"000011000",
  61475=>"100100100",
  61476=>"101001111",
  61477=>"101011100",
  61478=>"010111110",
  61479=>"100001111",
  61480=>"010101110",
  61481=>"010001101",
  61482=>"110111010",
  61483=>"101110111",
  61484=>"001111100",
  61485=>"110010101",
  61486=>"001000011",
  61487=>"111001010",
  61488=>"000000111",
  61489=>"000111101",
  61490=>"111101001",
  61491=>"011010100",
  61492=>"000100100",
  61493=>"010011010",
  61494=>"101100000",
  61495=>"011111010",
  61496=>"000110000",
  61497=>"100000111",
  61498=>"001001001",
  61499=>"000011011",
  61500=>"111111011",
  61501=>"000111100",
  61502=>"011000010",
  61503=>"011001110",
  61504=>"111011110",
  61505=>"001110110",
  61506=>"010011001",
  61507=>"111001010",
  61508=>"000101010",
  61509=>"110011111",
  61510=>"001001001",
  61511=>"100011101",
  61512=>"011110001",
  61513=>"011100110",
  61514=>"110000010",
  61515=>"001111111",
  61516=>"101110000",
  61517=>"101110001",
  61518=>"110111011",
  61519=>"000010010",
  61520=>"101010010",
  61521=>"110000110",
  61522=>"111000001",
  61523=>"101001001",
  61524=>"000110000",
  61525=>"010010010",
  61526=>"000001101",
  61527=>"010010111",
  61528=>"101011010",
  61529=>"000000100",
  61530=>"101011000",
  61531=>"111011110",
  61532=>"000010000",
  61533=>"111011111",
  61534=>"001100000",
  61535=>"001110001",
  61536=>"111001001",
  61537=>"011101001",
  61538=>"110100101",
  61539=>"101001011",
  61540=>"111110011",
  61541=>"001011111",
  61542=>"101100110",
  61543=>"010000010",
  61544=>"101011011",
  61545=>"100100101",
  61546=>"000110100",
  61547=>"110101110",
  61548=>"100001111",
  61549=>"110110101",
  61550=>"101011111",
  61551=>"011101101",
  61552=>"001100110",
  61553=>"000000110",
  61554=>"001000100",
  61555=>"111110110",
  61556=>"010010011",
  61557=>"010100110",
  61558=>"010101101",
  61559=>"111110110",
  61560=>"000000100",
  61561=>"111011001",
  61562=>"011101100",
  61563=>"100110011",
  61564=>"001100101",
  61565=>"110111110",
  61566=>"100101001",
  61567=>"000101010",
  61568=>"101000110",
  61569=>"010000101",
  61570=>"100001101",
  61571=>"111101000",
  61572=>"110111000",
  61573=>"000100001",
  61574=>"011101100",
  61575=>"110100100",
  61576=>"000011001",
  61577=>"110010011",
  61578=>"011010111",
  61579=>"101110011",
  61580=>"010001011",
  61581=>"001100110",
  61582=>"111011000",
  61583=>"010101101",
  61584=>"110110011",
  61585=>"001100010",
  61586=>"111011011",
  61587=>"100001111",
  61588=>"000111101",
  61589=>"010010011",
  61590=>"110111011",
  61591=>"101000100",
  61592=>"110001000",
  61593=>"010100001",
  61594=>"100101111",
  61595=>"100101011",
  61596=>"010111011",
  61597=>"011110010",
  61598=>"101000000",
  61599=>"011000100",
  61600=>"101101101",
  61601=>"100111001",
  61602=>"010100100",
  61603=>"110000101",
  61604=>"101001011",
  61605=>"101110100",
  61606=>"101010001",
  61607=>"101010010",
  61608=>"110110101",
  61609=>"111101010",
  61610=>"111001010",
  61611=>"011111100",
  61612=>"111111010",
  61613=>"111010111",
  61614=>"011000011",
  61615=>"010101000",
  61616=>"000010111",
  61617=>"011011101",
  61618=>"101100111",
  61619=>"001100111",
  61620=>"111110010",
  61621=>"100100000",
  61622=>"100011101",
  61623=>"001100111",
  61624=>"101100110",
  61625=>"001110001",
  61626=>"001101000",
  61627=>"011001001",
  61628=>"011101001",
  61629=>"111011001",
  61630=>"111101100",
  61631=>"100110001",
  61632=>"011100000",
  61633=>"101000001",
  61634=>"101110001",
  61635=>"010011010",
  61636=>"110111000",
  61637=>"101010010",
  61638=>"111110110",
  61639=>"111100000",
  61640=>"010000110",
  61641=>"011111001",
  61642=>"110101101",
  61643=>"101100111",
  61644=>"000100111",
  61645=>"011101100",
  61646=>"100001000",
  61647=>"000011100",
  61648=>"111101010",
  61649=>"011010010",
  61650=>"010000111",
  61651=>"100101110",
  61652=>"101101000",
  61653=>"110110011",
  61654=>"110100110",
  61655=>"100110110",
  61656=>"101110011",
  61657=>"001110011",
  61658=>"010101101",
  61659=>"001011111",
  61660=>"010000100",
  61661=>"000111010",
  61662=>"010111000",
  61663=>"000000100",
  61664=>"010100100",
  61665=>"000000100",
  61666=>"010110110",
  61667=>"111011001",
  61668=>"001111010",
  61669=>"011010111",
  61670=>"100001101",
  61671=>"000100100",
  61672=>"001111011",
  61673=>"100001100",
  61674=>"111001110",
  61675=>"000010111",
  61676=>"001111101",
  61677=>"100010100",
  61678=>"100010000",
  61679=>"110010101",
  61680=>"100000101",
  61681=>"100011010",
  61682=>"001111110",
  61683=>"011101000",
  61684=>"010010110",
  61685=>"010110101",
  61686=>"101100101",
  61687=>"001001111",
  61688=>"000000011",
  61689=>"100011111",
  61690=>"000000010",
  61691=>"011110010",
  61692=>"100110110",
  61693=>"011000000",
  61694=>"110111110",
  61695=>"100000011",
  61696=>"111100101",
  61697=>"011100100",
  61698=>"111001011",
  61699=>"111000111",
  61700=>"010111001",
  61701=>"001111110",
  61702=>"001011001",
  61703=>"111100110",
  61704=>"010000100",
  61705=>"110101111",
  61706=>"001111111",
  61707=>"000010110",
  61708=>"010100000",
  61709=>"111010010",
  61710=>"101100001",
  61711=>"101000111",
  61712=>"010011001",
  61713=>"010101000",
  61714=>"011011110",
  61715=>"010010001",
  61716=>"110001110",
  61717=>"111100001",
  61718=>"000001001",
  61719=>"011110110",
  61720=>"011000001",
  61721=>"110010101",
  61722=>"010111111",
  61723=>"101110110",
  61724=>"010100011",
  61725=>"001111011",
  61726=>"111111010",
  61727=>"000111000",
  61728=>"011011010",
  61729=>"111000010",
  61730=>"011101010",
  61731=>"110100100",
  61732=>"011001001",
  61733=>"101111001",
  61734=>"000100100",
  61735=>"011100111",
  61736=>"111000001",
  61737=>"100011110",
  61738=>"111001111",
  61739=>"010100111",
  61740=>"110111111",
  61741=>"001101000",
  61742=>"110001111",
  61743=>"111000111",
  61744=>"111001111",
  61745=>"111101111",
  61746=>"011010111",
  61747=>"011000111",
  61748=>"100110101",
  61749=>"010000011",
  61750=>"110000101",
  61751=>"000101010",
  61752=>"101011101",
  61753=>"100010100",
  61754=>"011110100",
  61755=>"000010001",
  61756=>"000000110",
  61757=>"111110001",
  61758=>"100111111",
  61759=>"011001011",
  61760=>"111100011",
  61761=>"000010011",
  61762=>"001011010",
  61763=>"011100100",
  61764=>"110100100",
  61765=>"011100110",
  61766=>"111111111",
  61767=>"000111101",
  61768=>"000101100",
  61769=>"100011110",
  61770=>"001011101",
  61771=>"010000011",
  61772=>"001101101",
  61773=>"010101100",
  61774=>"110000100",
  61775=>"111011001",
  61776=>"001011010",
  61777=>"101011001",
  61778=>"110111001",
  61779=>"000110110",
  61780=>"101100000",
  61781=>"010100011",
  61782=>"100101111",
  61783=>"011011011",
  61784=>"000101100",
  61785=>"001011011",
  61786=>"111011100",
  61787=>"111110110",
  61788=>"100110110",
  61789=>"011010010",
  61790=>"011110100",
  61791=>"011110111",
  61792=>"000000001",
  61793=>"111010101",
  61794=>"111101101",
  61795=>"101000110",
  61796=>"001000100",
  61797=>"000000101",
  61798=>"111110011",
  61799=>"011011110",
  61800=>"110011011",
  61801=>"110011000",
  61802=>"100001111",
  61803=>"001000000",
  61804=>"111111100",
  61805=>"110011010",
  61806=>"011110000",
  61807=>"011011011",
  61808=>"101001110",
  61809=>"010111011",
  61810=>"110010011",
  61811=>"010111110",
  61812=>"011000011",
  61813=>"000100001",
  61814=>"011110000",
  61815=>"110101000",
  61816=>"111010110",
  61817=>"111110111",
  61818=>"110101100",
  61819=>"110110101",
  61820=>"110001101",
  61821=>"010001010",
  61822=>"011000100",
  61823=>"110010111",
  61824=>"001011010",
  61825=>"010001000",
  61826=>"000111010",
  61827=>"001100100",
  61828=>"011001010",
  61829=>"011111000",
  61830=>"100111101",
  61831=>"011001011",
  61832=>"000000010",
  61833=>"011000010",
  61834=>"101001010",
  61835=>"011100000",
  61836=>"110110000",
  61837=>"010111000",
  61838=>"010010010",
  61839=>"001110010",
  61840=>"010100010",
  61841=>"011110101",
  61842=>"110010110",
  61843=>"101111011",
  61844=>"011001110",
  61845=>"101100110",
  61846=>"001111110",
  61847=>"111001001",
  61848=>"001110011",
  61849=>"001010011",
  61850=>"100000110",
  61851=>"001001111",
  61852=>"111010100",
  61853=>"011100010",
  61854=>"000000101",
  61855=>"110001001",
  61856=>"100101001",
  61857=>"111111101",
  61858=>"001011101",
  61859=>"000011001",
  61860=>"100000010",
  61861=>"111100101",
  61862=>"000000000",
  61863=>"101110100",
  61864=>"010100010",
  61865=>"011011000",
  61866=>"110111001",
  61867=>"010001110",
  61868=>"100101110",
  61869=>"100111110",
  61870=>"010000010",
  61871=>"000011010",
  61872=>"110000110",
  61873=>"110000100",
  61874=>"010110001",
  61875=>"111000010",
  61876=>"111111011",
  61877=>"010010110",
  61878=>"100101001",
  61879=>"101110111",
  61880=>"111000110",
  61881=>"100010000",
  61882=>"110101101",
  61883=>"101110111",
  61884=>"100100001",
  61885=>"010010101",
  61886=>"110010101",
  61887=>"011100101",
  61888=>"100101000",
  61889=>"111101100",
  61890=>"001000100",
  61891=>"011111011",
  61892=>"010110000",
  61893=>"010110011",
  61894=>"011110001",
  61895=>"011010010",
  61896=>"101001010",
  61897=>"001000111",
  61898=>"100100001",
  61899=>"100110011",
  61900=>"101000111",
  61901=>"001001000",
  61902=>"111111001",
  61903=>"101001100",
  61904=>"001010010",
  61905=>"000110100",
  61906=>"100011111",
  61907=>"010101110",
  61908=>"001110001",
  61909=>"101100001",
  61910=>"101111011",
  61911=>"000011010",
  61912=>"001101101",
  61913=>"100101000",
  61914=>"100100110",
  61915=>"110000100",
  61916=>"111110010",
  61917=>"110011101",
  61918=>"001011011",
  61919=>"000100101",
  61920=>"101110000",
  61921=>"101101111",
  61922=>"000000001",
  61923=>"001010110",
  61924=>"000010111",
  61925=>"100000011",
  61926=>"110001011",
  61927=>"000000110",
  61928=>"010110001",
  61929=>"001110111",
  61930=>"010101011",
  61931=>"000110111",
  61932=>"010010110",
  61933=>"011101100",
  61934=>"001000111",
  61935=>"010000001",
  61936=>"111111111",
  61937=>"100111111",
  61938=>"101011111",
  61939=>"000010101",
  61940=>"101011100",
  61941=>"000000000",
  61942=>"011101001",
  61943=>"000010001",
  61944=>"100010001",
  61945=>"100001000",
  61946=>"001101101",
  61947=>"100110111",
  61948=>"001000000",
  61949=>"011010100",
  61950=>"111011000",
  61951=>"100010011",
  61952=>"010111100",
  61953=>"100011100",
  61954=>"111000011",
  61955=>"011111011",
  61956=>"001011111",
  61957=>"010100110",
  61958=>"111111111",
  61959=>"010100110",
  61960=>"010101010",
  61961=>"101001000",
  61962=>"101001101",
  61963=>"111100100",
  61964=>"110111110",
  61965=>"111001100",
  61966=>"000000000",
  61967=>"111001001",
  61968=>"000111010",
  61969=>"010000100",
  61970=>"011100100",
  61971=>"010011100",
  61972=>"110110011",
  61973=>"111110010",
  61974=>"101110101",
  61975=>"110001111",
  61976=>"100000010",
  61977=>"011111011",
  61978=>"011010001",
  61979=>"010111010",
  61980=>"001010010",
  61981=>"000110011",
  61982=>"000111010",
  61983=>"010000010",
  61984=>"101001010",
  61985=>"010100000",
  61986=>"111001011",
  61987=>"111111111",
  61988=>"111000001",
  61989=>"100010010",
  61990=>"101101011",
  61991=>"010110010",
  61992=>"101001111",
  61993=>"111111111",
  61994=>"111010110",
  61995=>"011110010",
  61996=>"111000111",
  61997=>"110000011",
  61998=>"101011000",
  61999=>"010111011",
  62000=>"110010101",
  62001=>"110101000",
  62002=>"111110101",
  62003=>"001010001",
  62004=>"110011111",
  62005=>"011110111",
  62006=>"001000100",
  62007=>"010010110",
  62008=>"011111110",
  62009=>"101010000",
  62010=>"010100111",
  62011=>"001000000",
  62012=>"011101001",
  62013=>"001111101",
  62014=>"101011101",
  62015=>"000011111",
  62016=>"110101011",
  62017=>"111110101",
  62018=>"000001000",
  62019=>"101001111",
  62020=>"011111111",
  62021=>"110110100",
  62022=>"000011001",
  62023=>"000100100",
  62024=>"011010000",
  62025=>"001101011",
  62026=>"100101001",
  62027=>"111011000",
  62028=>"101011000",
  62029=>"001000000",
  62030=>"000110100",
  62031=>"101111000",
  62032=>"100000100",
  62033=>"011010010",
  62034=>"000010101",
  62035=>"100100101",
  62036=>"001101111",
  62037=>"010100110",
  62038=>"111100111",
  62039=>"010100111",
  62040=>"010100011",
  62041=>"110011001",
  62042=>"000110100",
  62043=>"010000101",
  62044=>"101010101",
  62045=>"100001000",
  62046=>"000100111",
  62047=>"101111001",
  62048=>"100010101",
  62049=>"000010100",
  62050=>"001011101",
  62051=>"111100011",
  62052=>"000000010",
  62053=>"101111111",
  62054=>"010011001",
  62055=>"000010000",
  62056=>"111010111",
  62057=>"101110111",
  62058=>"010010010",
  62059=>"001100111",
  62060=>"001001111",
  62061=>"110101111",
  62062=>"111101100",
  62063=>"101100001",
  62064=>"111010010",
  62065=>"011101000",
  62066=>"010100011",
  62067=>"101010000",
  62068=>"101000001",
  62069=>"101010001",
  62070=>"111001101",
  62071=>"011110100",
  62072=>"001100100",
  62073=>"001101000",
  62074=>"000110010",
  62075=>"000110101",
  62076=>"101001111",
  62077=>"010111110",
  62078=>"111100101",
  62079=>"010110110",
  62080=>"100110100",
  62081=>"100110110",
  62082=>"110110101",
  62083=>"100100010",
  62084=>"100110011",
  62085=>"001100000",
  62086=>"101111111",
  62087=>"011100101",
  62088=>"000101011",
  62089=>"010000010",
  62090=>"101111000",
  62091=>"001000000",
  62092=>"010111000",
  62093=>"001010010",
  62094=>"011100100",
  62095=>"110010111",
  62096=>"011000010",
  62097=>"000110110",
  62098=>"101000110",
  62099=>"100000010",
  62100=>"100111011",
  62101=>"100001111",
  62102=>"010100101",
  62103=>"101001111",
  62104=>"010100011",
  62105=>"111011110",
  62106=>"100101111",
  62107=>"101010011",
  62108=>"111010010",
  62109=>"101000001",
  62110=>"101001111",
  62111=>"001010101",
  62112=>"101000001",
  62113=>"000000111",
  62114=>"111001101",
  62115=>"011010010",
  62116=>"010100100",
  62117=>"000111100",
  62118=>"010100011",
  62119=>"011010011",
  62120=>"010111110",
  62121=>"100000010",
  62122=>"011010110",
  62123=>"110111101",
  62124=>"000000001",
  62125=>"100111111",
  62126=>"010000010",
  62127=>"011101011",
  62128=>"011010111",
  62129=>"001100111",
  62130=>"101001001",
  62131=>"100110110",
  62132=>"100110101",
  62133=>"010010101",
  62134=>"101001010",
  62135=>"010110111",
  62136=>"001101000",
  62137=>"101011100",
  62138=>"000111100",
  62139=>"001110000",
  62140=>"001010010",
  62141=>"010000000",
  62142=>"101001001",
  62143=>"001100000",
  62144=>"100100110",
  62145=>"010010110",
  62146=>"101100011",
  62147=>"111000111",
  62148=>"000111110",
  62149=>"010110001",
  62150=>"001000110",
  62151=>"110100100",
  62152=>"101101010",
  62153=>"100111110",
  62154=>"010010001",
  62155=>"111101101",
  62156=>"001100001",
  62157=>"101100000",
  62158=>"011110111",
  62159=>"011010111",
  62160=>"010100100",
  62161=>"111011110",
  62162=>"001110010",
  62163=>"111110011",
  62164=>"000011001",
  62165=>"111111111",
  62166=>"100010110",
  62167=>"001010000",
  62168=>"100010101",
  62169=>"111111100",
  62170=>"110100100",
  62171=>"000001110",
  62172=>"110110010",
  62173=>"111011011",
  62174=>"101101010",
  62175=>"001100011",
  62176=>"101110001",
  62177=>"101100000",
  62178=>"100011001",
  62179=>"011101001",
  62180=>"111110111",
  62181=>"101011100",
  62182=>"101001001",
  62183=>"011001101",
  62184=>"001110010",
  62185=>"000110001",
  62186=>"000110010",
  62187=>"010011010",
  62188=>"001101111",
  62189=>"001100011",
  62190=>"000011101",
  62191=>"000110100",
  62192=>"110010111",
  62193=>"111101101",
  62194=>"111010111",
  62195=>"011101110",
  62196=>"000101011",
  62197=>"010001111",
  62198=>"000100100",
  62199=>"110101111",
  62200=>"101101101",
  62201=>"100011101",
  62202=>"101011111",
  62203=>"000000111",
  62204=>"011000011",
  62205=>"110110101",
  62206=>"010111011",
  62207=>"000010001",
  62208=>"100001011",
  62209=>"000000001",
  62210=>"000001101",
  62211=>"101010100",
  62212=>"100011010",
  62213=>"011111001",
  62214=>"110111001",
  62215=>"001110001",
  62216=>"101111111",
  62217=>"010010000",
  62218=>"010100110",
  62219=>"011100111",
  62220=>"100011111",
  62221=>"110011011",
  62222=>"111110110",
  62223=>"111101100",
  62224=>"110111110",
  62225=>"010011110",
  62226=>"000011111",
  62227=>"001101110",
  62228=>"001111111",
  62229=>"110010010",
  62230=>"101010001",
  62231=>"110001011",
  62232=>"010001000",
  62233=>"010100010",
  62234=>"100000000",
  62235=>"011111001",
  62236=>"000001011",
  62237=>"001001000",
  62238=>"010001110",
  62239=>"011110011",
  62240=>"100101001",
  62241=>"010001101",
  62242=>"111010110",
  62243=>"111011100",
  62244=>"110100111",
  62245=>"101110010",
  62246=>"111011100",
  62247=>"111110001",
  62248=>"010000100",
  62249=>"000000001",
  62250=>"111001100",
  62251=>"001011000",
  62252=>"110100011",
  62253=>"001101111",
  62254=>"001011111",
  62255=>"001011010",
  62256=>"111000010",
  62257=>"111000100",
  62258=>"000000001",
  62259=>"110110100",
  62260=>"000001000",
  62261=>"101111101",
  62262=>"100100001",
  62263=>"001100010",
  62264=>"001011011",
  62265=>"111111110",
  62266=>"010111101",
  62267=>"000001101",
  62268=>"100010101",
  62269=>"101100000",
  62270=>"001000000",
  62271=>"000100111",
  62272=>"000001111",
  62273=>"100110111",
  62274=>"100101011",
  62275=>"010001001",
  62276=>"111111100",
  62277=>"000010011",
  62278=>"110100001",
  62279=>"111001100",
  62280=>"001111111",
  62281=>"111111011",
  62282=>"010111111",
  62283=>"010100011",
  62284=>"000101011",
  62285=>"010100001",
  62286=>"111101111",
  62287=>"100011100",
  62288=>"111111110",
  62289=>"010000010",
  62290=>"111100010",
  62291=>"100101100",
  62292=>"101111101",
  62293=>"000001010",
  62294=>"110011111",
  62295=>"100001011",
  62296=>"111011101",
  62297=>"101010011",
  62298=>"101101100",
  62299=>"111100010",
  62300=>"000000000",
  62301=>"111110100",
  62302=>"110111000",
  62303=>"111111110",
  62304=>"001100001",
  62305=>"011101010",
  62306=>"011000110",
  62307=>"101110001",
  62308=>"001111111",
  62309=>"010110001",
  62310=>"110111100",
  62311=>"000110010",
  62312=>"101100010",
  62313=>"010110101",
  62314=>"101100010",
  62315=>"101100010",
  62316=>"111101110",
  62317=>"111001000",
  62318=>"101010011",
  62319=>"000000001",
  62320=>"111011100",
  62321=>"010111101",
  62322=>"100001110",
  62323=>"010110101",
  62324=>"000011111",
  62325=>"101000000",
  62326=>"111010001",
  62327=>"000000000",
  62328=>"001011101",
  62329=>"100001101",
  62330=>"010100000",
  62331=>"001011110",
  62332=>"000110010",
  62333=>"011101101",
  62334=>"101000110",
  62335=>"011001000",
  62336=>"000110100",
  62337=>"011011010",
  62338=>"000101010",
  62339=>"010101010",
  62340=>"001110110",
  62341=>"001010000",
  62342=>"010110100",
  62343=>"111000101",
  62344=>"011011100",
  62345=>"111001110",
  62346=>"110101001",
  62347=>"101000110",
  62348=>"001100011",
  62349=>"100011010",
  62350=>"011010000",
  62351=>"001110001",
  62352=>"110011010",
  62353=>"001011010",
  62354=>"000000011",
  62355=>"000111010",
  62356=>"100100101",
  62357=>"110010100",
  62358=>"101110111",
  62359=>"011110011",
  62360=>"001001100",
  62361=>"111111100",
  62362=>"110100100",
  62363=>"000000011",
  62364=>"111101001",
  62365=>"011100101",
  62366=>"111001111",
  62367=>"110000000",
  62368=>"000000001",
  62369=>"100011100",
  62370=>"110011101",
  62371=>"111010111",
  62372=>"111101101",
  62373=>"000000100",
  62374=>"101010010",
  62375=>"101100110",
  62376=>"000011000",
  62377=>"101111100",
  62378=>"100000111",
  62379=>"010101111",
  62380=>"001010111",
  62381=>"011100110",
  62382=>"001011101",
  62383=>"111001011",
  62384=>"000011100",
  62385=>"001001011",
  62386=>"000101010",
  62387=>"011111011",
  62388=>"000010000",
  62389=>"000101110",
  62390=>"111111110",
  62391=>"001110101",
  62392=>"100011101",
  62393=>"100110110",
  62394=>"111000110",
  62395=>"010011000",
  62396=>"010010110",
  62397=>"001001001",
  62398=>"100100000",
  62399=>"111111110",
  62400=>"111001010",
  62401=>"010100001",
  62402=>"000111111",
  62403=>"001010101",
  62404=>"111110011",
  62405=>"111100100",
  62406=>"011110010",
  62407=>"100100011",
  62408=>"101010000",
  62409=>"011010000",
  62410=>"110111000",
  62411=>"010000101",
  62412=>"010101011",
  62413=>"101011000",
  62414=>"011000011",
  62415=>"101000000",
  62416=>"000100000",
  62417=>"011110100",
  62418=>"001010001",
  62419=>"111010001",
  62420=>"110001111",
  62421=>"001000000",
  62422=>"111000111",
  62423=>"000100000",
  62424=>"000100100",
  62425=>"110001100",
  62426=>"101100000",
  62427=>"001001001",
  62428=>"010010010",
  62429=>"011011001",
  62430=>"000110001",
  62431=>"001010110",
  62432=>"010001000",
  62433=>"000111000",
  62434=>"010111100",
  62435=>"111011000",
  62436=>"111111011",
  62437=>"111001000",
  62438=>"010110010",
  62439=>"111110000",
  62440=>"011111011",
  62441=>"110011001",
  62442=>"100110101",
  62443=>"000001100",
  62444=>"100001000",
  62445=>"111011111",
  62446=>"100100101",
  62447=>"100010001",
  62448=>"010111111",
  62449=>"100001011",
  62450=>"100101101",
  62451=>"011111110",
  62452=>"100010110",
  62453=>"000011010",
  62454=>"101100100",
  62455=>"100110110",
  62456=>"000100100",
  62457=>"111101010",
  62458=>"110010010",
  62459=>"111101111",
  62460=>"110001100",
  62461=>"010010101",
  62462=>"010000001",
  62463=>"100110110",
  62464=>"001111101",
  62465=>"000101010",
  62466=>"101001111",
  62467=>"011000100",
  62468=>"111101100",
  62469=>"110100110",
  62470=>"000111010",
  62471=>"110100111",
  62472=>"011101101",
  62473=>"010101100",
  62474=>"111100001",
  62475=>"101010000",
  62476=>"000000110",
  62477=>"110101100",
  62478=>"011001101",
  62479=>"101001000",
  62480=>"100101010",
  62481=>"111010010",
  62482=>"000101101",
  62483=>"110001001",
  62484=>"001100011",
  62485=>"011000010",
  62486=>"011100001",
  62487=>"001010010",
  62488=>"001010110",
  62489=>"101001100",
  62490=>"010010001",
  62491=>"100111111",
  62492=>"110010111",
  62493=>"111100000",
  62494=>"001111000",
  62495=>"101000001",
  62496=>"100000010",
  62497=>"111110011",
  62498=>"000010011",
  62499=>"101110000",
  62500=>"101111101",
  62501=>"000011001",
  62502=>"100010100",
  62503=>"010000001",
  62504=>"010101111",
  62505=>"001100001",
  62506=>"101100011",
  62507=>"000000011",
  62508=>"000010111",
  62509=>"101111010",
  62510=>"110010000",
  62511=>"110111011",
  62512=>"111001100",
  62513=>"110001011",
  62514=>"001110110",
  62515=>"111011110",
  62516=>"011110111",
  62517=>"010000111",
  62518=>"111111011",
  62519=>"111111000",
  62520=>"001101110",
  62521=>"000011100",
  62522=>"101011010",
  62523=>"101001000",
  62524=>"010001000",
  62525=>"010011001",
  62526=>"100100111",
  62527=>"111111001",
  62528=>"101100001",
  62529=>"000000101",
  62530=>"110100011",
  62531=>"010101001",
  62532=>"100100001",
  62533=>"010010001",
  62534=>"010011111",
  62535=>"001000100",
  62536=>"000100011",
  62537=>"000110100",
  62538=>"011010110",
  62539=>"101101000",
  62540=>"000011110",
  62541=>"100101111",
  62542=>"010101000",
  62543=>"000001010",
  62544=>"100110010",
  62545=>"111110101",
  62546=>"011111110",
  62547=>"110110110",
  62548=>"010011111",
  62549=>"011101011",
  62550=>"011011100",
  62551=>"110110011",
  62552=>"111010001",
  62553=>"100111110",
  62554=>"000001111",
  62555=>"001110000",
  62556=>"000000001",
  62557=>"010111001",
  62558=>"001101001",
  62559=>"000111000",
  62560=>"111000100",
  62561=>"100000101",
  62562=>"001000001",
  62563=>"000000000",
  62564=>"011000110",
  62565=>"001110101",
  62566=>"110101110",
  62567=>"110010000",
  62568=>"000101101",
  62569=>"011011001",
  62570=>"000001111",
  62571=>"111001100",
  62572=>"011110100",
  62573=>"000101110",
  62574=>"100010000",
  62575=>"011010000",
  62576=>"010011110",
  62577=>"100011000",
  62578=>"111110001",
  62579=>"000011101",
  62580=>"110111000",
  62581=>"001111001",
  62582=>"011011000",
  62583=>"000100010",
  62584=>"100001110",
  62585=>"000111111",
  62586=>"011111001",
  62587=>"001000100",
  62588=>"010000100",
  62589=>"111000110",
  62590=>"100100100",
  62591=>"111010100",
  62592=>"000000000",
  62593=>"101101001",
  62594=>"010111001",
  62595=>"110101011",
  62596=>"010000100",
  62597=>"010010011",
  62598=>"011011010",
  62599=>"011011011",
  62600=>"101010110",
  62601=>"101101101",
  62602=>"010110001",
  62603=>"001110111",
  62604=>"101000011",
  62605=>"110000010",
  62606=>"000010111",
  62607=>"001101000",
  62608=>"111101001",
  62609=>"011000011",
  62610=>"001011101",
  62611=>"110111101",
  62612=>"000000111",
  62613=>"110100010",
  62614=>"000100000",
  62615=>"101011110",
  62616=>"000000000",
  62617=>"101100000",
  62618=>"101001100",
  62619=>"011000000",
  62620=>"010011000",
  62621=>"001101001",
  62622=>"110000101",
  62623=>"110011101",
  62624=>"010010100",
  62625=>"110010111",
  62626=>"101011010",
  62627=>"001100111",
  62628=>"001011100",
  62629=>"110000011",
  62630=>"100011101",
  62631=>"100001011",
  62632=>"010011111",
  62633=>"100111110",
  62634=>"111111110",
  62635=>"101101101",
  62636=>"001000100",
  62637=>"011001100",
  62638=>"101010011",
  62639=>"010000010",
  62640=>"001000010",
  62641=>"100111111",
  62642=>"010100111",
  62643=>"110100000",
  62644=>"111011100",
  62645=>"101101101",
  62646=>"011000000",
  62647=>"000011001",
  62648=>"110000111",
  62649=>"111111010",
  62650=>"101011011",
  62651=>"011111111",
  62652=>"011100100",
  62653=>"000111101",
  62654=>"000000101",
  62655=>"011011110",
  62656=>"110110000",
  62657=>"101011010",
  62658=>"000010011",
  62659=>"111100011",
  62660=>"110010111",
  62661=>"011100010",
  62662=>"100010110",
  62663=>"010101001",
  62664=>"010000001",
  62665=>"010101111",
  62666=>"111011111",
  62667=>"010100101",
  62668=>"000111110",
  62669=>"011000110",
  62670=>"011011000",
  62671=>"111010000",
  62672=>"000001010",
  62673=>"010000101",
  62674=>"011100101",
  62675=>"110000011",
  62676=>"111010010",
  62677=>"001010010",
  62678=>"001011001",
  62679=>"101100011",
  62680=>"100111001",
  62681=>"100000100",
  62682=>"010010001",
  62683=>"111001000",
  62684=>"000100101",
  62685=>"000010001",
  62686=>"100011010",
  62687=>"110101011",
  62688=>"011110011",
  62689=>"111010111",
  62690=>"001000101",
  62691=>"101001100",
  62692=>"010110111",
  62693=>"101101011",
  62694=>"111010010",
  62695=>"111110011",
  62696=>"001001000",
  62697=>"100101111",
  62698=>"110000010",
  62699=>"001010111",
  62700=>"111010110",
  62701=>"001100010",
  62702=>"110110111",
  62703=>"011111010",
  62704=>"100111101",
  62705=>"110001001",
  62706=>"000000010",
  62707=>"101010011",
  62708=>"100001100",
  62709=>"101001101",
  62710=>"010001011",
  62711=>"001101100",
  62712=>"110001100",
  62713=>"001000100",
  62714=>"100100000",
  62715=>"000000101",
  62716=>"000100011",
  62717=>"001100001",
  62718=>"010111001",
  62719=>"001010000",
  62720=>"110111110",
  62721=>"110000110",
  62722=>"001111110",
  62723=>"100010010",
  62724=>"001001011",
  62725=>"101000110",
  62726=>"111100000",
  62727=>"010100001",
  62728=>"010110000",
  62729=>"010101111",
  62730=>"100010101",
  62731=>"111011010",
  62732=>"111011000",
  62733=>"000000111",
  62734=>"100001000",
  62735=>"011111010",
  62736=>"111101100",
  62737=>"011011001",
  62738=>"110010101",
  62739=>"111111111",
  62740=>"101111010",
  62741=>"100110101",
  62742=>"000110010",
  62743=>"111000011",
  62744=>"101011111",
  62745=>"111110111",
  62746=>"011110010",
  62747=>"000010111",
  62748=>"111010001",
  62749=>"000111100",
  62750=>"101100101",
  62751=>"101110100",
  62752=>"101101000",
  62753=>"010011011",
  62754=>"101001101",
  62755=>"011000100",
  62756=>"101110011",
  62757=>"100111000",
  62758=>"010000101",
  62759=>"010100001",
  62760=>"001000010",
  62761=>"100110000",
  62762=>"101100010",
  62763=>"001010000",
  62764=>"100100101",
  62765=>"110001100",
  62766=>"000000010",
  62767=>"110000011",
  62768=>"010110010",
  62769=>"101010111",
  62770=>"010110111",
  62771=>"011110001",
  62772=>"000101111",
  62773=>"101010011",
  62774=>"100000011",
  62775=>"101111101",
  62776=>"000011110",
  62777=>"001000011",
  62778=>"111001110",
  62779=>"100110011",
  62780=>"110000001",
  62781=>"010100000",
  62782=>"000010001",
  62783=>"111111111",
  62784=>"101010111",
  62785=>"100111010",
  62786=>"001000010",
  62787=>"101010000",
  62788=>"001111010",
  62789=>"110101001",
  62790=>"010100010",
  62791=>"101101100",
  62792=>"100011001",
  62793=>"100111000",
  62794=>"101000000",
  62795=>"110101001",
  62796=>"011110000",
  62797=>"110110100",
  62798=>"101000110",
  62799=>"110000011",
  62800=>"100010001",
  62801=>"100100010",
  62802=>"001110001",
  62803=>"001011111",
  62804=>"100110110",
  62805=>"001110011",
  62806=>"100111001",
  62807=>"110010110",
  62808=>"101010101",
  62809=>"100100110",
  62810=>"000110101",
  62811=>"010000011",
  62812=>"110011101",
  62813=>"001111001",
  62814=>"000100011",
  62815=>"000010111",
  62816=>"110101110",
  62817=>"111101100",
  62818=>"100100001",
  62819=>"000110000",
  62820=>"000101111",
  62821=>"001100100",
  62822=>"101000000",
  62823=>"001010110",
  62824=>"000011010",
  62825=>"001101000",
  62826=>"011001011",
  62827=>"000001111",
  62828=>"110001001",
  62829=>"111110111",
  62830=>"101010000",
  62831=>"010001110",
  62832=>"000010101",
  62833=>"001011110",
  62834=>"001110111",
  62835=>"000101101",
  62836=>"001010111",
  62837=>"011011100",
  62838=>"001110010",
  62839=>"011110011",
  62840=>"101001111",
  62841=>"111011010",
  62842=>"010000011",
  62843=>"000010011",
  62844=>"110010011",
  62845=>"111011001",
  62846=>"100011000",
  62847=>"111110011",
  62848=>"111111011",
  62849=>"111010111",
  62850=>"000111110",
  62851=>"001110101",
  62852=>"101111000",
  62853=>"001001011",
  62854=>"011011110",
  62855=>"010011111",
  62856=>"000100111",
  62857=>"111101001",
  62858=>"100001110",
  62859=>"100100111",
  62860=>"100010100",
  62861=>"001101100",
  62862=>"101010010",
  62863=>"100100110",
  62864=>"000111001",
  62865=>"100011111",
  62866=>"001010000",
  62867=>"111111100",
  62868=>"001001010",
  62869=>"100010100",
  62870=>"011010101",
  62871=>"000111101",
  62872=>"000101001",
  62873=>"101001100",
  62874=>"000111000",
  62875=>"001101100",
  62876=>"110010110",
  62877=>"001101100",
  62878=>"111011100",
  62879=>"111100111",
  62880=>"000111000",
  62881=>"000101000",
  62882=>"001111011",
  62883=>"000000100",
  62884=>"100100001",
  62885=>"000100000",
  62886=>"111000111",
  62887=>"110010111",
  62888=>"011101101",
  62889=>"010010001",
  62890=>"000010100",
  62891=>"000110100",
  62892=>"100010000",
  62893=>"100011111",
  62894=>"011010111",
  62895=>"000011110",
  62896=>"000010111",
  62897=>"001100100",
  62898=>"101000011",
  62899=>"111010011",
  62900=>"100011000",
  62901=>"101111000",
  62902=>"010001010",
  62903=>"010011110",
  62904=>"001110001",
  62905=>"011000001",
  62906=>"001111111",
  62907=>"101111111",
  62908=>"110111001",
  62909=>"100100010",
  62910=>"001000011",
  62911=>"011100010",
  62912=>"100111000",
  62913=>"010000010",
  62914=>"001001101",
  62915=>"001100110",
  62916=>"111001001",
  62917=>"111101111",
  62918=>"010010000",
  62919=>"000001101",
  62920=>"110010000",
  62921=>"100101111",
  62922=>"010001001",
  62923=>"000010101",
  62924=>"000000101",
  62925=>"100000111",
  62926=>"001100011",
  62927=>"001100011",
  62928=>"011001111",
  62929=>"001110111",
  62930=>"110111111",
  62931=>"111101000",
  62932=>"111100010",
  62933=>"111101110",
  62934=>"000000010",
  62935=>"111110101",
  62936=>"001010000",
  62937=>"000011000",
  62938=>"011101000",
  62939=>"011111000",
  62940=>"001111110",
  62941=>"001010011",
  62942=>"100001111",
  62943=>"001001111",
  62944=>"011001111",
  62945=>"110110000",
  62946=>"110010111",
  62947=>"111001001",
  62948=>"000100011",
  62949=>"010011111",
  62950=>"110100111",
  62951=>"011110100",
  62952=>"001001000",
  62953=>"111110010",
  62954=>"000101101",
  62955=>"111100101",
  62956=>"100010110",
  62957=>"001000000",
  62958=>"010000010",
  62959=>"110001101",
  62960=>"100100111",
  62961=>"101000100",
  62962=>"001110000",
  62963=>"011010010",
  62964=>"100101011",
  62965=>"101000110",
  62966=>"010110111",
  62967=>"001100111",
  62968=>"000011001",
  62969=>"001001110",
  62970=>"101110100",
  62971=>"100110000",
  62972=>"111111101",
  62973=>"010110011",
  62974=>"000000110",
  62975=>"001110111",
  62976=>"000100011",
  62977=>"000001111",
  62978=>"011111001",
  62979=>"011001010",
  62980=>"100010111",
  62981=>"101100000",
  62982=>"000011110",
  62983=>"001110001",
  62984=>"010001110",
  62985=>"010011010",
  62986=>"011000010",
  62987=>"000100000",
  62988=>"101101011",
  62989=>"110101111",
  62990=>"111100001",
  62991=>"000100000",
  62992=>"000110110",
  62993=>"101111110",
  62994=>"010001010",
  62995=>"101001011",
  62996=>"010010000",
  62997=>"010100010",
  62998=>"110000001",
  62999=>"001010011",
  63000=>"111110101",
  63001=>"100001000",
  63002=>"010100000",
  63003=>"111000110",
  63004=>"000000111",
  63005=>"110101000",
  63006=>"100111100",
  63007=>"111101010",
  63008=>"110100100",
  63009=>"101111011",
  63010=>"001000000",
  63011=>"001111100",
  63012=>"100001011",
  63013=>"011111001",
  63014=>"111110111",
  63015=>"001110010",
  63016=>"100011110",
  63017=>"000001100",
  63018=>"000011100",
  63019=>"000001011",
  63020=>"100000110",
  63021=>"000110010",
  63022=>"111011001",
  63023=>"000100110",
  63024=>"001110010",
  63025=>"110100000",
  63026=>"010101010",
  63027=>"111111000",
  63028=>"011000101",
  63029=>"100101001",
  63030=>"001000010",
  63031=>"000111100",
  63032=>"010111101",
  63033=>"110111101",
  63034=>"110010001",
  63035=>"001000101",
  63036=>"011100000",
  63037=>"111000111",
  63038=>"100001010",
  63039=>"011010111",
  63040=>"100100011",
  63041=>"001000111",
  63042=>"011100001",
  63043=>"110011110",
  63044=>"011100011",
  63045=>"000011110",
  63046=>"000100100",
  63047=>"100100111",
  63048=>"000110110",
  63049=>"111110000",
  63050=>"001001000",
  63051=>"100001010",
  63052=>"110001000",
  63053=>"001010001",
  63054=>"001111111",
  63055=>"001000000",
  63056=>"011111101",
  63057=>"111011101",
  63058=>"111100010",
  63059=>"011100010",
  63060=>"001110001",
  63061=>"000111001",
  63062=>"000110100",
  63063=>"010000011",
  63064=>"000000001",
  63065=>"001110010",
  63066=>"001101011",
  63067=>"000000001",
  63068=>"010010010",
  63069=>"100110011",
  63070=>"110110001",
  63071=>"110110111",
  63072=>"011101011",
  63073=>"111110000",
  63074=>"100101011",
  63075=>"010010100",
  63076=>"111111101",
  63077=>"000000101",
  63078=>"000011011",
  63079=>"001001010",
  63080=>"111001000",
  63081=>"001011100",
  63082=>"011010111",
  63083=>"100000100",
  63084=>"010001001",
  63085=>"111000000",
  63086=>"111101000",
  63087=>"001011101",
  63088=>"000000011",
  63089=>"111100110",
  63090=>"101101100",
  63091=>"000111001",
  63092=>"001000010",
  63093=>"110001101",
  63094=>"010000101",
  63095=>"000000110",
  63096=>"100000100",
  63097=>"101101011",
  63098=>"101111111",
  63099=>"001000101",
  63100=>"101000110",
  63101=>"000110011",
  63102=>"001001011",
  63103=>"010110111",
  63104=>"110001101",
  63105=>"110111001",
  63106=>"001101000",
  63107=>"000010100",
  63108=>"010101001",
  63109=>"000000110",
  63110=>"000111101",
  63111=>"111010000",
  63112=>"000101010",
  63113=>"000010100",
  63114=>"010110111",
  63115=>"101110010",
  63116=>"010010001",
  63117=>"111001011",
  63118=>"111001001",
  63119=>"001101100",
  63120=>"111110110",
  63121=>"011110011",
  63122=>"011101110",
  63123=>"111010101",
  63124=>"111100010",
  63125=>"001101000",
  63126=>"000111010",
  63127=>"010010110",
  63128=>"110010111",
  63129=>"110100010",
  63130=>"110001001",
  63131=>"110111111",
  63132=>"011110000",
  63133=>"010001000",
  63134=>"010100000",
  63135=>"100000101",
  63136=>"100011000",
  63137=>"000010101",
  63138=>"010000111",
  63139=>"100000000",
  63140=>"010001111",
  63141=>"101110101",
  63142=>"011111010",
  63143=>"001001001",
  63144=>"011111100",
  63145=>"001100001",
  63146=>"001011110",
  63147=>"001001100",
  63148=>"101000111",
  63149=>"000101001",
  63150=>"000110001",
  63151=>"100000001",
  63152=>"100101101",
  63153=>"000011101",
  63154=>"111111011",
  63155=>"000101010",
  63156=>"100100010",
  63157=>"100001010",
  63158=>"110100011",
  63159=>"101110010",
  63160=>"100110000",
  63161=>"100001010",
  63162=>"101111011",
  63163=>"011011111",
  63164=>"000100100",
  63165=>"000000010",
  63166=>"111011000",
  63167=>"100101111",
  63168=>"001110100",
  63169=>"110011101",
  63170=>"110011101",
  63171=>"011011001",
  63172=>"111110010",
  63173=>"101000101",
  63174=>"010110000",
  63175=>"011101111",
  63176=>"100000110",
  63177=>"001111001",
  63178=>"100101110",
  63179=>"000010000",
  63180=>"001000110",
  63181=>"111111001",
  63182=>"011011111",
  63183=>"110010110",
  63184=>"001101111",
  63185=>"110011011",
  63186=>"010011011",
  63187=>"111010000",
  63188=>"101010101",
  63189=>"001011010",
  63190=>"000110000",
  63191=>"001111101",
  63192=>"111110011",
  63193=>"001000000",
  63194=>"110100011",
  63195=>"010101011",
  63196=>"011011100",
  63197=>"111000001",
  63198=>"000011000",
  63199=>"000111110",
  63200=>"011110111",
  63201=>"001110010",
  63202=>"100101100",
  63203=>"010100001",
  63204=>"011011100",
  63205=>"000000101",
  63206=>"101011001",
  63207=>"101001100",
  63208=>"101110101",
  63209=>"011100101",
  63210=>"010100011",
  63211=>"011000011",
  63212=>"011001010",
  63213=>"110010111",
  63214=>"100101011",
  63215=>"010001111",
  63216=>"101110100",
  63217=>"011000001",
  63218=>"010100100",
  63219=>"001110011",
  63220=>"011001100",
  63221=>"110111101",
  63222=>"010010011",
  63223=>"011001011",
  63224=>"100101011",
  63225=>"001101011",
  63226=>"010110000",
  63227=>"100110110",
  63228=>"111010111",
  63229=>"111010110",
  63230=>"010110100",
  63231=>"001111110",
  63232=>"010101101",
  63233=>"000110011",
  63234=>"110110111",
  63235=>"001100000",
  63236=>"011111000",
  63237=>"101001001",
  63238=>"010001000",
  63239=>"111101010",
  63240=>"111000000",
  63241=>"111000111",
  63242=>"001110101",
  63243=>"010110110",
  63244=>"110011101",
  63245=>"011100111",
  63246=>"000001100",
  63247=>"011001000",
  63248=>"100100110",
  63249=>"101001110",
  63250=>"101111110",
  63251=>"011101001",
  63252=>"011011000",
  63253=>"010000100",
  63254=>"111000101",
  63255=>"000111010",
  63256=>"001000000",
  63257=>"000000111",
  63258=>"010010000",
  63259=>"011000100",
  63260=>"111110111",
  63261=>"011011001",
  63262=>"100100110",
  63263=>"111100110",
  63264=>"110001101",
  63265=>"101000111",
  63266=>"100010100",
  63267=>"110010000",
  63268=>"110000010",
  63269=>"110001000",
  63270=>"111011010",
  63271=>"010110101",
  63272=>"111101101",
  63273=>"100001101",
  63274=>"111100110",
  63275=>"110011011",
  63276=>"001100000",
  63277=>"101110010",
  63278=>"000001100",
  63279=>"000011011",
  63280=>"011111001",
  63281=>"001010000",
  63282=>"010001110",
  63283=>"010001100",
  63284=>"011010111",
  63285=>"010010100",
  63286=>"110110100",
  63287=>"111010110",
  63288=>"111101110",
  63289=>"100000111",
  63290=>"110101000",
  63291=>"101000011",
  63292=>"111000011",
  63293=>"000100101",
  63294=>"010100001",
  63295=>"100000101",
  63296=>"011110000",
  63297=>"110000010",
  63298=>"101010110",
  63299=>"011000110",
  63300=>"111001101",
  63301=>"110011110",
  63302=>"110000100",
  63303=>"010011111",
  63304=>"000000101",
  63305=>"111111001",
  63306=>"101001111",
  63307=>"000001110",
  63308=>"110010010",
  63309=>"100011011",
  63310=>"000010101",
  63311=>"110111101",
  63312=>"001011100",
  63313=>"000101011",
  63314=>"111111001",
  63315=>"001101111",
  63316=>"000111010",
  63317=>"110001000",
  63318=>"000100011",
  63319=>"000001100",
  63320=>"110101111",
  63321=>"100100000",
  63322=>"111011100",
  63323=>"011111111",
  63324=>"010001110",
  63325=>"000010110",
  63326=>"100000111",
  63327=>"000001111",
  63328=>"001101000",
  63329=>"001101100",
  63330=>"101011100",
  63331=>"000111101",
  63332=>"100001000",
  63333=>"000001101",
  63334=>"111001000",
  63335=>"110111010",
  63336=>"111001100",
  63337=>"101101101",
  63338=>"011010100",
  63339=>"101101001",
  63340=>"001010000",
  63341=>"111000110",
  63342=>"111000101",
  63343=>"100010001",
  63344=>"111111110",
  63345=>"101000001",
  63346=>"001011010",
  63347=>"101001001",
  63348=>"000000111",
  63349=>"100000100",
  63350=>"100010001",
  63351=>"001100001",
  63352=>"101101010",
  63353=>"001101101",
  63354=>"100001000",
  63355=>"100011011",
  63356=>"010000000",
  63357=>"011111000",
  63358=>"101111101",
  63359=>"000000010",
  63360=>"010100100",
  63361=>"010111000",
  63362=>"000110010",
  63363=>"001110001",
  63364=>"100011010",
  63365=>"111000000",
  63366=>"000010110",
  63367=>"001100100",
  63368=>"011100001",
  63369=>"110101111",
  63370=>"000011101",
  63371=>"111000001",
  63372=>"000010111",
  63373=>"001100001",
  63374=>"000000010",
  63375=>"111101000",
  63376=>"111000110",
  63377=>"010101101",
  63378=>"101001111",
  63379=>"000110110",
  63380=>"110010111",
  63381=>"011010110",
  63382=>"100010100",
  63383=>"001101000",
  63384=>"010001000",
  63385=>"001110001",
  63386=>"110111001",
  63387=>"000010100",
  63388=>"111100111",
  63389=>"101111000",
  63390=>"111110100",
  63391=>"100011001",
  63392=>"011111000",
  63393=>"001000010",
  63394=>"111011010",
  63395=>"010110101",
  63396=>"000001110",
  63397=>"110111010",
  63398=>"000100100",
  63399=>"011101000",
  63400=>"001011000",
  63401=>"010110100",
  63402=>"101101100",
  63403=>"001000011",
  63404=>"111000000",
  63405=>"010100101",
  63406=>"011000111",
  63407=>"101111111",
  63408=>"000101110",
  63409=>"100100110",
  63410=>"011011101",
  63411=>"011101101",
  63412=>"001100000",
  63413=>"000001011",
  63414=>"001101011",
  63415=>"111100100",
  63416=>"011011011",
  63417=>"011110110",
  63418=>"110110111",
  63419=>"000111101",
  63420=>"011110001",
  63421=>"100000111",
  63422=>"101010110",
  63423=>"000110111",
  63424=>"001011100",
  63425=>"011000010",
  63426=>"110010110",
  63427=>"001010100",
  63428=>"101101100",
  63429=>"010000010",
  63430=>"101010000",
  63431=>"101100101",
  63432=>"111100101",
  63433=>"000001000",
  63434=>"111100110",
  63435=>"100000000",
  63436=>"101110101",
  63437=>"110011011",
  63438=>"010100110",
  63439=>"010001110",
  63440=>"111100101",
  63441=>"010001110",
  63442=>"110011111",
  63443=>"011011100",
  63444=>"011100101",
  63445=>"100011001",
  63446=>"010010101",
  63447=>"100001001",
  63448=>"000110000",
  63449=>"110010111",
  63450=>"100110100",
  63451=>"100110000",
  63452=>"011101011",
  63453=>"010001001",
  63454=>"000110010",
  63455=>"111000011",
  63456=>"001000001",
  63457=>"001111111",
  63458=>"011111011",
  63459=>"100101011",
  63460=>"111010000",
  63461=>"001010100",
  63462=>"011100000",
  63463=>"111101000",
  63464=>"000000010",
  63465=>"110100111",
  63466=>"001100100",
  63467=>"110100000",
  63468=>"111101011",
  63469=>"000001101",
  63470=>"100111111",
  63471=>"000100110",
  63472=>"001100010",
  63473=>"111101001",
  63474=>"111000100",
  63475=>"010110001",
  63476=>"001000100",
  63477=>"000000001",
  63478=>"111110101",
  63479=>"000101010",
  63480=>"111101011",
  63481=>"000011111",
  63482=>"011010100",
  63483=>"010100011",
  63484=>"110100000",
  63485=>"001100110",
  63486=>"100010000",
  63487=>"001101001",
  63488=>"000010000",
  63489=>"000000100",
  63490=>"110100101",
  63491=>"000100101",
  63492=>"001100110",
  63493=>"010000100",
  63494=>"001100001",
  63495=>"101110001",
  63496=>"001010110",
  63497=>"001001000",
  63498=>"011111110",
  63499=>"010001010",
  63500=>"000011001",
  63501=>"110011100",
  63502=>"000111100",
  63503=>"101110011",
  63504=>"010111110",
  63505=>"111000001",
  63506=>"100100100",
  63507=>"100010000",
  63508=>"100001001",
  63509=>"000101101",
  63510=>"011100111",
  63511=>"011010010",
  63512=>"010110010",
  63513=>"110011001",
  63514=>"000100111",
  63515=>"101000010",
  63516=>"111111110",
  63517=>"001000001",
  63518=>"110111111",
  63519=>"100100101",
  63520=>"101111010",
  63521=>"010100001",
  63522=>"111010110",
  63523=>"100111100",
  63524=>"111101100",
  63525=>"101100001",
  63526=>"110010101",
  63527=>"010001011",
  63528=>"110011001",
  63529=>"001001000",
  63530=>"111110101",
  63531=>"101101100",
  63532=>"010000010",
  63533=>"001110001",
  63534=>"101010000",
  63535=>"100001111",
  63536=>"110010010",
  63537=>"111011001",
  63538=>"010110010",
  63539=>"000001011",
  63540=>"100000011",
  63541=>"000111100",
  63542=>"110111111",
  63543=>"111101010",
  63544=>"000010011",
  63545=>"110011000",
  63546=>"100101110",
  63547=>"111010000",
  63548=>"011100001",
  63549=>"010010110",
  63550=>"010001011",
  63551=>"101100101",
  63552=>"110100110",
  63553=>"101011000",
  63554=>"001001000",
  63555=>"011011001",
  63556=>"001001011",
  63557=>"111100101",
  63558=>"111010111",
  63559=>"000010110",
  63560=>"101011011",
  63561=>"000100100",
  63562=>"010100101",
  63563=>"011101001",
  63564=>"011100110",
  63565=>"000110100",
  63566=>"001110100",
  63567=>"010011011",
  63568=>"011001111",
  63569=>"011010111",
  63570=>"000111101",
  63571=>"100000010",
  63572=>"110101110",
  63573=>"110111101",
  63574=>"001110011",
  63575=>"001101111",
  63576=>"000001111",
  63577=>"100100000",
  63578=>"011000011",
  63579=>"000011011",
  63580=>"000011010",
  63581=>"001000001",
  63582=>"111101000",
  63583=>"010101101",
  63584=>"000111000",
  63585=>"110001010",
  63586=>"100100100",
  63587=>"101000110",
  63588=>"101010110",
  63589=>"000001011",
  63590=>"011100011",
  63591=>"111111011",
  63592=>"111111010",
  63593=>"101100111",
  63594=>"100101111",
  63595=>"101010110",
  63596=>"111100100",
  63597=>"110010010",
  63598=>"000001100",
  63599=>"000111000",
  63600=>"101010100",
  63601=>"111000100",
  63602=>"111111101",
  63603=>"111011111",
  63604=>"000010101",
  63605=>"001011100",
  63606=>"110100011",
  63607=>"111111110",
  63608=>"110111001",
  63609=>"011111100",
  63610=>"000110010",
  63611=>"100101011",
  63612=>"001111110",
  63613=>"000111101",
  63614=>"010000001",
  63615=>"101101000",
  63616=>"000010110",
  63617=>"111100111",
  63618=>"100010001",
  63619=>"011011000",
  63620=>"000011001",
  63621=>"101100010",
  63622=>"110110101",
  63623=>"001000111",
  63624=>"000111001",
  63625=>"010010101",
  63626=>"110110101",
  63627=>"001011101",
  63628=>"011110001",
  63629=>"011001011",
  63630=>"100011000",
  63631=>"111000110",
  63632=>"000100111",
  63633=>"111001101",
  63634=>"101011101",
  63635=>"011011110",
  63636=>"101001100",
  63637=>"100100101",
  63638=>"000000100",
  63639=>"110101001",
  63640=>"000000100",
  63641=>"011101010",
  63642=>"111010000",
  63643=>"101100011",
  63644=>"001011111",
  63645=>"110111100",
  63646=>"101001010",
  63647=>"100011000",
  63648=>"100110111",
  63649=>"000100111",
  63650=>"000100110",
  63651=>"111001100",
  63652=>"100011100",
  63653=>"111101001",
  63654=>"100111000",
  63655=>"110000101",
  63656=>"111101110",
  63657=>"011101101",
  63658=>"111110011",
  63659=>"011101110",
  63660=>"111111000",
  63661=>"100100011",
  63662=>"011100100",
  63663=>"010101110",
  63664=>"001000110",
  63665=>"100001010",
  63666=>"000101010",
  63667=>"100000110",
  63668=>"001000010",
  63669=>"010001101",
  63670=>"100101010",
  63671=>"111111111",
  63672=>"101010001",
  63673=>"111110000",
  63674=>"100111000",
  63675=>"010000001",
  63676=>"110001101",
  63677=>"000110111",
  63678=>"010001000",
  63679=>"101110100",
  63680=>"100100110",
  63681=>"101101111",
  63682=>"111111111",
  63683=>"100111101",
  63684=>"101001110",
  63685=>"011101101",
  63686=>"010100010",
  63687=>"101100010",
  63688=>"001000000",
  63689=>"100010001",
  63690=>"111000001",
  63691=>"010011001",
  63692=>"101011001",
  63693=>"000101110",
  63694=>"100011001",
  63695=>"001011101",
  63696=>"000101101",
  63697=>"110101011",
  63698=>"001110110",
  63699=>"000101000",
  63700=>"101111110",
  63701=>"111000011",
  63702=>"100000111",
  63703=>"100010100",
  63704=>"000100110",
  63705=>"011000001",
  63706=>"101111101",
  63707=>"010111110",
  63708=>"110101101",
  63709=>"010100110",
  63710=>"011110000",
  63711=>"001011010",
  63712=>"111100011",
  63713=>"111110010",
  63714=>"001101001",
  63715=>"010010011",
  63716=>"101010111",
  63717=>"001010110",
  63718=>"110110010",
  63719=>"110001101",
  63720=>"111111111",
  63721=>"110111001",
  63722=>"100001000",
  63723=>"010111000",
  63724=>"100010111",
  63725=>"101110000",
  63726=>"110010100",
  63727=>"011101111",
  63728=>"100101101",
  63729=>"001101001",
  63730=>"111100010",
  63731=>"010111010",
  63732=>"011111101",
  63733=>"000111100",
  63734=>"010110010",
  63735=>"101101000",
  63736=>"110101111",
  63737=>"110111001",
  63738=>"000001101",
  63739=>"110101101",
  63740=>"011000011",
  63741=>"010101111",
  63742=>"000100000",
  63743=>"111100101",
  63744=>"110111011",
  63745=>"100101100",
  63746=>"000101110",
  63747=>"100001101",
  63748=>"100101000",
  63749=>"111111101",
  63750=>"111010001",
  63751=>"000001101",
  63752=>"000011110",
  63753=>"010010100",
  63754=>"011101110",
  63755=>"000010110",
  63756=>"001100011",
  63757=>"110110001",
  63758=>"000100110",
  63759=>"000000001",
  63760=>"111000111",
  63761=>"101001010",
  63762=>"111010011",
  63763=>"111101111",
  63764=>"010010100",
  63765=>"100111100",
  63766=>"010110111",
  63767=>"110001001",
  63768=>"101000001",
  63769=>"000100010",
  63770=>"101001111",
  63771=>"000011111",
  63772=>"001011110",
  63773=>"011100010",
  63774=>"110111010",
  63775=>"001100001",
  63776=>"000000010",
  63777=>"101000011",
  63778=>"111101100",
  63779=>"010100011",
  63780=>"101110101",
  63781=>"011001100",
  63782=>"000001100",
  63783=>"000100000",
  63784=>"110010101",
  63785=>"011111101",
  63786=>"110000011",
  63787=>"101011111",
  63788=>"111110000",
  63789=>"000000001",
  63790=>"111111010",
  63791=>"110111101",
  63792=>"000101000",
  63793=>"011101001",
  63794=>"101001010",
  63795=>"010110010",
  63796=>"101111011",
  63797=>"011110000",
  63798=>"010011011",
  63799=>"101010101",
  63800=>"001101101",
  63801=>"011100000",
  63802=>"001100101",
  63803=>"000000000",
  63804=>"110000110",
  63805=>"011001000",
  63806=>"010001011",
  63807=>"111111001",
  63808=>"100100100",
  63809=>"000000011",
  63810=>"110111111",
  63811=>"011101101",
  63812=>"000111100",
  63813=>"111100111",
  63814=>"000100100",
  63815=>"000001111",
  63816=>"010010100",
  63817=>"010011110",
  63818=>"100001011",
  63819=>"000000101",
  63820=>"100001011",
  63821=>"000111111",
  63822=>"010011100",
  63823=>"111011110",
  63824=>"101111111",
  63825=>"001010111",
  63826=>"000010101",
  63827=>"000000000",
  63828=>"100010001",
  63829=>"011010010",
  63830=>"000000011",
  63831=>"100100110",
  63832=>"110100101",
  63833=>"111111110",
  63834=>"001101011",
  63835=>"101100010",
  63836=>"101100010",
  63837=>"101010010",
  63838=>"110111011",
  63839=>"111000110",
  63840=>"001000010",
  63841=>"001100000",
  63842=>"101100101",
  63843=>"101001001",
  63844=>"100111000",
  63845=>"000010100",
  63846=>"001001001",
  63847=>"010000010",
  63848=>"111100111",
  63849=>"010100110",
  63850=>"010010010",
  63851=>"100110011",
  63852=>"111101011",
  63853=>"110110101",
  63854=>"101100100",
  63855=>"111001001",
  63856=>"010110001",
  63857=>"011010011",
  63858=>"010011001",
  63859=>"100010011",
  63860=>"010010001",
  63861=>"100001001",
  63862=>"110101010",
  63863=>"011001101",
  63864=>"000001111",
  63865=>"100001101",
  63866=>"101100110",
  63867=>"101011100",
  63868=>"010110001",
  63869=>"111110111",
  63870=>"110010100",
  63871=>"000110001",
  63872=>"110001000",
  63873=>"010110000",
  63874=>"101111011",
  63875=>"110101110",
  63876=>"011111011",
  63877=>"111111011",
  63878=>"010111000",
  63879=>"111000011",
  63880=>"111100010",
  63881=>"011111010",
  63882=>"110011111",
  63883=>"111110010",
  63884=>"010011010",
  63885=>"001000111",
  63886=>"100010011",
  63887=>"010100001",
  63888=>"110001111",
  63889=>"100010000",
  63890=>"101011111",
  63891=>"110001101",
  63892=>"101100110",
  63893=>"000001011",
  63894=>"100001110",
  63895=>"111100010",
  63896=>"010001111",
  63897=>"101000001",
  63898=>"000011001",
  63899=>"101001011",
  63900=>"110101101",
  63901=>"000010000",
  63902=>"010100101",
  63903=>"000100000",
  63904=>"111010111",
  63905=>"000110101",
  63906=>"000001000",
  63907=>"110110011",
  63908=>"101110001",
  63909=>"100011000",
  63910=>"001000101",
  63911=>"010001000",
  63912=>"011010101",
  63913=>"011110101",
  63914=>"001000111",
  63915=>"011001000",
  63916=>"001010110",
  63917=>"011101100",
  63918=>"010101110",
  63919=>"001110000",
  63920=>"000100000",
  63921=>"010111111",
  63922=>"001110000",
  63923=>"011100000",
  63924=>"010100110",
  63925=>"101111100",
  63926=>"101111101",
  63927=>"101001101",
  63928=>"010111110",
  63929=>"000100111",
  63930=>"011100110",
  63931=>"011110001",
  63932=>"110010000",
  63933=>"100011010",
  63934=>"110111011",
  63935=>"111011100",
  63936=>"011110001",
  63937=>"000011100",
  63938=>"010110100",
  63939=>"110000011",
  63940=>"000110011",
  63941=>"100101000",
  63942=>"010110010",
  63943=>"010010000",
  63944=>"111110001",
  63945=>"100001110",
  63946=>"010110111",
  63947=>"110110101",
  63948=>"011000010",
  63949=>"010110101",
  63950=>"001100111",
  63951=>"111011010",
  63952=>"110011111",
  63953=>"111010100",
  63954=>"010111010",
  63955=>"100001001",
  63956=>"011110111",
  63957=>"100010001",
  63958=>"111100100",
  63959=>"111110000",
  63960=>"100001101",
  63961=>"110001010",
  63962=>"111000001",
  63963=>"110001011",
  63964=>"000010000",
  63965=>"010000101",
  63966=>"000000101",
  63967=>"110011010",
  63968=>"110111100",
  63969=>"100101011",
  63970=>"011000000",
  63971=>"011101110",
  63972=>"110110001",
  63973=>"101011001",
  63974=>"111100111",
  63975=>"000101000",
  63976=>"000101111",
  63977=>"000101001",
  63978=>"111010111",
  63979=>"011010110",
  63980=>"001000100",
  63981=>"010001011",
  63982=>"101101111",
  63983=>"100101111",
  63984=>"110100011",
  63985=>"010000101",
  63986=>"010101000",
  63987=>"111110010",
  63988=>"010100100",
  63989=>"000010011",
  63990=>"111111110",
  63991=>"000100100",
  63992=>"000011011",
  63993=>"010100110",
  63994=>"100000011",
  63995=>"011010101",
  63996=>"000010011",
  63997=>"111001000",
  63998=>"010011101",
  63999=>"010001000",
  64000=>"111110001",
  64001=>"011000000",
  64002=>"000001110",
  64003=>"110010100",
  64004=>"010110000",
  64005=>"111101000",
  64006=>"011010110",
  64007=>"011000101",
  64008=>"100001100",
  64009=>"101101011",
  64010=>"111110000",
  64011=>"000011001",
  64012=>"011011100",
  64013=>"111000010",
  64014=>"000000000",
  64015=>"010110100",
  64016=>"010000000",
  64017=>"100011010",
  64018=>"010101011",
  64019=>"011001010",
  64020=>"011101010",
  64021=>"000000111",
  64022=>"110111100",
  64023=>"000010110",
  64024=>"100100001",
  64025=>"010000000",
  64026=>"000000000",
  64027=>"001010010",
  64028=>"011100001",
  64029=>"101010011",
  64030=>"101110100",
  64031=>"101101111",
  64032=>"110011010",
  64033=>"100111001",
  64034=>"101101100",
  64035=>"111001010",
  64036=>"000100111",
  64037=>"000010111",
  64038=>"101110111",
  64039=>"101000110",
  64040=>"100000100",
  64041=>"010000001",
  64042=>"010000011",
  64043=>"001100111",
  64044=>"001000111",
  64045=>"010101000",
  64046=>"010010111",
  64047=>"000100011",
  64048=>"100011110",
  64049=>"011010100",
  64050=>"111101110",
  64051=>"000111000",
  64052=>"000010110",
  64053=>"000110110",
  64054=>"011111111",
  64055=>"011001100",
  64056=>"000011001",
  64057=>"010000000",
  64058=>"111101111",
  64059=>"110111010",
  64060=>"001100001",
  64061=>"011011110",
  64062=>"110011010",
  64063=>"101001110",
  64064=>"000100100",
  64065=>"110011001",
  64066=>"110010000",
  64067=>"101101000",
  64068=>"101110110",
  64069=>"010010100",
  64070=>"111001010",
  64071=>"000000000",
  64072=>"010000001",
  64073=>"110110010",
  64074=>"010111010",
  64075=>"110111110",
  64076=>"010000011",
  64077=>"001000100",
  64078=>"000001100",
  64079=>"001001101",
  64080=>"101101000",
  64081=>"000000101",
  64082=>"110110001",
  64083=>"100101110",
  64084=>"000111000",
  64085=>"110001111",
  64086=>"001000010",
  64087=>"010111100",
  64088=>"010001110",
  64089=>"011110100",
  64090=>"100011101",
  64091=>"110111010",
  64092=>"100001101",
  64093=>"001001110",
  64094=>"111110001",
  64095=>"001010011",
  64096=>"010011111",
  64097=>"010000000",
  64098=>"001000000",
  64099=>"011010011",
  64100=>"111110110",
  64101=>"010111111",
  64102=>"010011101",
  64103=>"011011100",
  64104=>"001111010",
  64105=>"001110010",
  64106=>"011101100",
  64107=>"010100000",
  64108=>"011110101",
  64109=>"001101101",
  64110=>"000011000",
  64111=>"100011100",
  64112=>"011101100",
  64113=>"111111110",
  64114=>"100101100",
  64115=>"111101011",
  64116=>"110001100",
  64117=>"010101111",
  64118=>"111001111",
  64119=>"011010111",
  64120=>"111110001",
  64121=>"100100000",
  64122=>"000111111",
  64123=>"101110111",
  64124=>"000111001",
  64125=>"011110111",
  64126=>"101101010",
  64127=>"010010110",
  64128=>"001110100",
  64129=>"100110010",
  64130=>"010111101",
  64131=>"111101100",
  64132=>"011010010",
  64133=>"101000010",
  64134=>"001100001",
  64135=>"111110000",
  64136=>"111111110",
  64137=>"001000011",
  64138=>"111000100",
  64139=>"000110011",
  64140=>"001111001",
  64141=>"100010000",
  64142=>"011000010",
  64143=>"001010000",
  64144=>"110101100",
  64145=>"011110010",
  64146=>"100100111",
  64147=>"011010100",
  64148=>"110001101",
  64149=>"011110100",
  64150=>"101000101",
  64151=>"100000010",
  64152=>"010110111",
  64153=>"001111000",
  64154=>"101111110",
  64155=>"101000111",
  64156=>"101110001",
  64157=>"111111011",
  64158=>"001001110",
  64159=>"111110100",
  64160=>"111101110",
  64161=>"011000101",
  64162=>"110101100",
  64163=>"011010100",
  64164=>"110110000",
  64165=>"110010110",
  64166=>"010110001",
  64167=>"001110100",
  64168=>"111111010",
  64169=>"001111111",
  64170=>"100010000",
  64171=>"100100000",
  64172=>"001100110",
  64173=>"001100100",
  64174=>"000000110",
  64175=>"001001000",
  64176=>"110010011",
  64177=>"011110100",
  64178=>"000110001",
  64179=>"010101100",
  64180=>"001110101",
  64181=>"000101010",
  64182=>"010001010",
  64183=>"001111100",
  64184=>"001001001",
  64185=>"100110000",
  64186=>"101110001",
  64187=>"000000000",
  64188=>"100101100",
  64189=>"000001110",
  64190=>"010101001",
  64191=>"111101001",
  64192=>"111010100",
  64193=>"000100010",
  64194=>"100100101",
  64195=>"011000010",
  64196=>"011101100",
  64197=>"100000101",
  64198=>"110101000",
  64199=>"100010010",
  64200=>"100001000",
  64201=>"000010000",
  64202=>"001100000",
  64203=>"111110011",
  64204=>"011001000",
  64205=>"100011111",
  64206=>"100111111",
  64207=>"100001100",
  64208=>"110011010",
  64209=>"100101100",
  64210=>"110000000",
  64211=>"001011000",
  64212=>"100011101",
  64213=>"000110011",
  64214=>"001101011",
  64215=>"001110110",
  64216=>"010000110",
  64217=>"000000100",
  64218=>"111110111",
  64219=>"111100001",
  64220=>"110010011",
  64221=>"000101110",
  64222=>"110001000",
  64223=>"001101000",
  64224=>"110101111",
  64225=>"101111101",
  64226=>"101110111",
  64227=>"010110100",
  64228=>"101100000",
  64229=>"000010010",
  64230=>"100110101",
  64231=>"111101111",
  64232=>"101111001",
  64233=>"111101010",
  64234=>"101000000",
  64235=>"101011000",
  64236=>"111001111",
  64237=>"001100011",
  64238=>"011001011",
  64239=>"100011110",
  64240=>"110111001",
  64241=>"010110101",
  64242=>"001001011",
  64243=>"000000111",
  64244=>"010001011",
  64245=>"010010110",
  64246=>"101000110",
  64247=>"010000010",
  64248=>"010001000",
  64249=>"010001111",
  64250=>"111011111",
  64251=>"000100111",
  64252=>"001101011",
  64253=>"101100110",
  64254=>"000100001",
  64255=>"101011110",
  64256=>"001010010",
  64257=>"110110011",
  64258=>"110111110",
  64259=>"000010000",
  64260=>"100001001",
  64261=>"000010000",
  64262=>"110011001",
  64263=>"111110100",
  64264=>"010100110",
  64265=>"110111101",
  64266=>"001101110",
  64267=>"101010101",
  64268=>"000101000",
  64269=>"001111111",
  64270=>"000000001",
  64271=>"110000001",
  64272=>"000101100",
  64273=>"010101100",
  64274=>"001010101",
  64275=>"100000101",
  64276=>"000111011",
  64277=>"010111001",
  64278=>"111110101",
  64279=>"010001001",
  64280=>"110111101",
  64281=>"000000000",
  64282=>"000010101",
  64283=>"001011110",
  64284=>"001111100",
  64285=>"001010000",
  64286=>"110011110",
  64287=>"000110000",
  64288=>"011111100",
  64289=>"000010111",
  64290=>"010100101",
  64291=>"110100011",
  64292=>"000101011",
  64293=>"110100000",
  64294=>"111001110",
  64295=>"110001111",
  64296=>"011110100",
  64297=>"000110011",
  64298=>"000000011",
  64299=>"001001010",
  64300=>"010011110",
  64301=>"000011111",
  64302=>"100000001",
  64303=>"001000010",
  64304=>"010010011",
  64305=>"101000000",
  64306=>"111111001",
  64307=>"100010011",
  64308=>"100111011",
  64309=>"010111001",
  64310=>"011110011",
  64311=>"101010101",
  64312=>"001000100",
  64313=>"001000101",
  64314=>"011001001",
  64315=>"101001000",
  64316=>"010101000",
  64317=>"001011110",
  64318=>"101011000",
  64319=>"111001001",
  64320=>"000001000",
  64321=>"110100110",
  64322=>"010111010",
  64323=>"110101011",
  64324=>"110011110",
  64325=>"101010101",
  64326=>"000000110",
  64327=>"001001101",
  64328=>"000101000",
  64329=>"010111101",
  64330=>"111000010",
  64331=>"101011111",
  64332=>"111111111",
  64333=>"111001000",
  64334=>"101100010",
  64335=>"111110100",
  64336=>"111000101",
  64337=>"100101100",
  64338=>"011101011",
  64339=>"011001001",
  64340=>"000010111",
  64341=>"110110101",
  64342=>"101110100",
  64343=>"001101000",
  64344=>"000001011",
  64345=>"110001000",
  64346=>"011100010",
  64347=>"100000010",
  64348=>"010000110",
  64349=>"010100011",
  64350=>"110110111",
  64351=>"101010001",
  64352=>"010100011",
  64353=>"100010111",
  64354=>"001101101",
  64355=>"111010110",
  64356=>"010111110",
  64357=>"000100100",
  64358=>"101010100",
  64359=>"001111111",
  64360=>"000111101",
  64361=>"010111010",
  64362=>"011111001",
  64363=>"100001101",
  64364=>"010110000",
  64365=>"100001001",
  64366=>"111011000",
  64367=>"100100001",
  64368=>"000100011",
  64369=>"101010011",
  64370=>"001001000",
  64371=>"111110000",
  64372=>"010111110",
  64373=>"010100100",
  64374=>"111110001",
  64375=>"011100100",
  64376=>"111111101",
  64377=>"100110011",
  64378=>"001011111",
  64379=>"011110001",
  64380=>"000110000",
  64381=>"000011101",
  64382=>"101000101",
  64383=>"110110111",
  64384=>"011100001",
  64385=>"101111010",
  64386=>"000010101",
  64387=>"000000000",
  64388=>"000100100",
  64389=>"101111101",
  64390=>"010100111",
  64391=>"111000111",
  64392=>"101110100",
  64393=>"100101101",
  64394=>"101000000",
  64395=>"101110001",
  64396=>"111111100",
  64397=>"000111101",
  64398=>"101110101",
  64399=>"101111110",
  64400=>"101110001",
  64401=>"000001011",
  64402=>"011110110",
  64403=>"101101011",
  64404=>"010000010",
  64405=>"110000101",
  64406=>"110101111",
  64407=>"011011010",
  64408=>"100010100",
  64409=>"000010110",
  64410=>"100110100",
  64411=>"110010010",
  64412=>"000010100",
  64413=>"100010111",
  64414=>"101000001",
  64415=>"001111111",
  64416=>"011101010",
  64417=>"000100000",
  64418=>"111111000",
  64419=>"100001101",
  64420=>"111010000",
  64421=>"001011111",
  64422=>"000001101",
  64423=>"011011010",
  64424=>"000110110",
  64425=>"111111101",
  64426=>"000011001",
  64427=>"101111000",
  64428=>"110101011",
  64429=>"010011011",
  64430=>"011101000",
  64431=>"010100110",
  64432=>"110101010",
  64433=>"000010110",
  64434=>"111101011",
  64435=>"010010001",
  64436=>"000100011",
  64437=>"111111111",
  64438=>"110000000",
  64439=>"111001101",
  64440=>"111000010",
  64441=>"110011101",
  64442=>"100000010",
  64443=>"011011100",
  64444=>"111111001",
  64445=>"010010000",
  64446=>"110010001",
  64447=>"110100100",
  64448=>"011011110",
  64449=>"101000100",
  64450=>"110100101",
  64451=>"101111010",
  64452=>"111001011",
  64453=>"100101011",
  64454=>"111110101",
  64455=>"111100111",
  64456=>"011000010",
  64457=>"101111110",
  64458=>"110001100",
  64459=>"001111001",
  64460=>"111011011",
  64461=>"100111100",
  64462=>"101101111",
  64463=>"101100101",
  64464=>"000111111",
  64465=>"101001110",
  64466=>"101000110",
  64467=>"100000110",
  64468=>"100101111",
  64469=>"000001001",
  64470=>"011111101",
  64471=>"111110101",
  64472=>"010100010",
  64473=>"111101010",
  64474=>"000010111",
  64475=>"100101110",
  64476=>"001101010",
  64477=>"001011110",
  64478=>"000001011",
  64479=>"001000000",
  64480=>"110101110",
  64481=>"001111111",
  64482=>"101111110",
  64483=>"110010110",
  64484=>"011011000",
  64485=>"000000001",
  64486=>"101000100",
  64487=>"001010000",
  64488=>"101000011",
  64489=>"000100000",
  64490=>"110100101",
  64491=>"000000000",
  64492=>"111010110",
  64493=>"100010010",
  64494=>"111110100",
  64495=>"011101000",
  64496=>"111101011",
  64497=>"100000110",
  64498=>"010100000",
  64499=>"111110000",
  64500=>"010010001",
  64501=>"000100100",
  64502=>"111111000",
  64503=>"111101101",
  64504=>"010011111",
  64505=>"100111100",
  64506=>"011011011",
  64507=>"100011010",
  64508=>"100000010",
  64509=>"001100010",
  64510=>"000111111",
  64511=>"111000001",
  64512=>"110001100",
  64513=>"110010100",
  64514=>"111111100",
  64515=>"000111110",
  64516=>"110111001",
  64517=>"100110111",
  64518=>"001000111",
  64519=>"011110100",
  64520=>"110000000",
  64521=>"111110101",
  64522=>"100100001",
  64523=>"100101000",
  64524=>"110000100",
  64525=>"010110100",
  64526=>"011101101",
  64527=>"101001100",
  64528=>"001000000",
  64529=>"101000010",
  64530=>"010110000",
  64531=>"011000100",
  64532=>"011011101",
  64533=>"111001111",
  64534=>"001001011",
  64535=>"010111000",
  64536=>"001011001",
  64537=>"110101000",
  64538=>"111100110",
  64539=>"011111101",
  64540=>"001011101",
  64541=>"010011001",
  64542=>"001000100",
  64543=>"010100100",
  64544=>"011111001",
  64545=>"000010111",
  64546=>"100110010",
  64547=>"001000110",
  64548=>"110111010",
  64549=>"011000100",
  64550=>"111110101",
  64551=>"111010101",
  64552=>"001011001",
  64553=>"111101100",
  64554=>"110111000",
  64555=>"111110011",
  64556=>"101010001",
  64557=>"110111011",
  64558=>"001010000",
  64559=>"010000111",
  64560=>"100010010",
  64561=>"010110100",
  64562=>"000000001",
  64563=>"111111001",
  64564=>"100111100",
  64565=>"001001110",
  64566=>"101000000",
  64567=>"100001010",
  64568=>"111011100",
  64569=>"011000000",
  64570=>"000001101",
  64571=>"001101010",
  64572=>"001010000",
  64573=>"000011101",
  64574=>"111100100",
  64575=>"010001100",
  64576=>"001010000",
  64577=>"000010010",
  64578=>"011111011",
  64579=>"111010011",
  64580=>"101101101",
  64581=>"111010110",
  64582=>"000001001",
  64583=>"001011001",
  64584=>"000101001",
  64585=>"101111111",
  64586=>"110001101",
  64587=>"111011010",
  64588=>"000010111",
  64589=>"111010110",
  64590=>"011100111",
  64591=>"100101110",
  64592=>"000000100",
  64593=>"000110000",
  64594=>"101011100",
  64595=>"000111011",
  64596=>"010110001",
  64597=>"010000001",
  64598=>"110000101",
  64599=>"001000000",
  64600=>"011110011",
  64601=>"011110000",
  64602=>"010011110",
  64603=>"000001100",
  64604=>"100010110",
  64605=>"100011011",
  64606=>"110111001",
  64607=>"001000111",
  64608=>"001100000",
  64609=>"011111011",
  64610=>"011010001",
  64611=>"011101100",
  64612=>"011011011",
  64613=>"110100100",
  64614=>"001010010",
  64615=>"101010010",
  64616=>"111111001",
  64617=>"010100010",
  64618=>"100111111",
  64619=>"010110000",
  64620=>"101110101",
  64621=>"010111010",
  64622=>"100110011",
  64623=>"000101010",
  64624=>"100011100",
  64625=>"000000111",
  64626=>"011000100",
  64627=>"011100111",
  64628=>"100000011",
  64629=>"101111000",
  64630=>"100101100",
  64631=>"001111100",
  64632=>"000000110",
  64633=>"001011010",
  64634=>"010011000",
  64635=>"000111111",
  64636=>"010110010",
  64637=>"000011100",
  64638=>"001000100",
  64639=>"011111010",
  64640=>"110100000",
  64641=>"100001111",
  64642=>"001000000",
  64643=>"001011111",
  64644=>"011001010",
  64645=>"001110010",
  64646=>"011101101",
  64647=>"001000101",
  64648=>"100001010",
  64649=>"010101010",
  64650=>"001011100",
  64651=>"110100011",
  64652=>"000000011",
  64653=>"001110011",
  64654=>"100100101",
  64655=>"111011111",
  64656=>"001110000",
  64657=>"111100101",
  64658=>"100000111",
  64659=>"001011000",
  64660=>"011100011",
  64661=>"110100111",
  64662=>"011001110",
  64663=>"111001010",
  64664=>"100111110",
  64665=>"110111000",
  64666=>"101010001",
  64667=>"010010010",
  64668=>"011110100",
  64669=>"100001111",
  64670=>"101101101",
  64671=>"110001010",
  64672=>"010111010",
  64673=>"111011011",
  64674=>"010110011",
  64675=>"111000110",
  64676=>"100111000",
  64677=>"011001101",
  64678=>"101000100",
  64679=>"000010001",
  64680=>"010010001",
  64681=>"111111000",
  64682=>"111111011",
  64683=>"001001001",
  64684=>"111001110",
  64685=>"100010100",
  64686=>"110000001",
  64687=>"110011000",
  64688=>"110000000",
  64689=>"101101001",
  64690=>"001100100",
  64691=>"111111111",
  64692=>"010001001",
  64693=>"100001001",
  64694=>"000100011",
  64695=>"011010001",
  64696=>"001000101",
  64697=>"000000001",
  64698=>"101110010",
  64699=>"100011111",
  64700=>"011010010",
  64701=>"001110000",
  64702=>"100000100",
  64703=>"000001100",
  64704=>"110000110",
  64705=>"100001101",
  64706=>"011001001",
  64707=>"000010100",
  64708=>"000000110",
  64709=>"001000010",
  64710=>"001000010",
  64711=>"100011011",
  64712=>"000110011",
  64713=>"111011011",
  64714=>"001010011",
  64715=>"111000001",
  64716=>"111000111",
  64717=>"110010011",
  64718=>"001011000",
  64719=>"000001110",
  64720=>"101010001",
  64721=>"001011001",
  64722=>"101110010",
  64723=>"101000100",
  64724=>"110100010",
  64725=>"000101000",
  64726=>"100101001",
  64727=>"111111101",
  64728=>"010101010",
  64729=>"101001111",
  64730=>"001111110",
  64731=>"001010010",
  64732=>"111111010",
  64733=>"110110110",
  64734=>"001100011",
  64735=>"101100001",
  64736=>"101011010",
  64737=>"001001110",
  64738=>"000000111",
  64739=>"111011011",
  64740=>"111001011",
  64741=>"011111110",
  64742=>"101101010",
  64743=>"000000101",
  64744=>"011010101",
  64745=>"101000011",
  64746=>"100010111",
  64747=>"110111100",
  64748=>"001100100",
  64749=>"101010101",
  64750=>"011110000",
  64751=>"100000011",
  64752=>"001011001",
  64753=>"000001101",
  64754=>"000001101",
  64755=>"010110000",
  64756=>"001011010",
  64757=>"001100100",
  64758=>"011001000",
  64759=>"000110010",
  64760=>"001100110",
  64761=>"110010000",
  64762=>"111100001",
  64763=>"111101110",
  64764=>"000001101",
  64765=>"001110010",
  64766=>"110011010",
  64767=>"101010000",
  64768=>"001101111",
  64769=>"110000100",
  64770=>"001100011",
  64771=>"010110010",
  64772=>"000100001",
  64773=>"111101011",
  64774=>"100111111",
  64775=>"000100101",
  64776=>"001111101",
  64777=>"011100011",
  64778=>"111011010",
  64779=>"100011100",
  64780=>"000001001",
  64781=>"000000110",
  64782=>"111111111",
  64783=>"010001010",
  64784=>"000011011",
  64785=>"011001110",
  64786=>"111000011",
  64787=>"011011110",
  64788=>"000011110",
  64789=>"010000011",
  64790=>"010101101",
  64791=>"010000000",
  64792=>"001000011",
  64793=>"100000000",
  64794=>"010100100",
  64795=>"011101100",
  64796=>"000110111",
  64797=>"011001100",
  64798=>"101111101",
  64799=>"110010010",
  64800=>"000110101",
  64801=>"000010001",
  64802=>"101011111",
  64803=>"100101101",
  64804=>"011101101",
  64805=>"010100100",
  64806=>"110110111",
  64807=>"101011111",
  64808=>"100001101",
  64809=>"100010001",
  64810=>"001111101",
  64811=>"010010100",
  64812=>"011011010",
  64813=>"101001001",
  64814=>"011101111",
  64815=>"001011111",
  64816=>"001001110",
  64817=>"111111000",
  64818=>"111111001",
  64819=>"011001111",
  64820=>"100000111",
  64821=>"010000010",
  64822=>"000100000",
  64823=>"011000110",
  64824=>"001001100",
  64825=>"110001011",
  64826=>"000000100",
  64827=>"111010100",
  64828=>"000100100",
  64829=>"000011100",
  64830=>"110010110",
  64831=>"110001111",
  64832=>"111010101",
  64833=>"011011111",
  64834=>"000010001",
  64835=>"111010010",
  64836=>"001011110",
  64837=>"110010110",
  64838=>"000100011",
  64839=>"101000101",
  64840=>"011101100",
  64841=>"111010011",
  64842=>"110011010",
  64843=>"001010100",
  64844=>"010000010",
  64845=>"101010100",
  64846=>"100111100",
  64847=>"111100111",
  64848=>"000011100",
  64849=>"100111011",
  64850=>"101011010",
  64851=>"000011010",
  64852=>"111101001",
  64853=>"000100100",
  64854=>"100111010",
  64855=>"000100000",
  64856=>"000111011",
  64857=>"100001011",
  64858=>"111001010",
  64859=>"000000001",
  64860=>"101110000",
  64861=>"100100000",
  64862=>"001001100",
  64863=>"100100100",
  64864=>"000101111",
  64865=>"111101110",
  64866=>"100101001",
  64867=>"001101110",
  64868=>"010110000",
  64869=>"001001100",
  64870=>"100010001",
  64871=>"111111111",
  64872=>"011111001",
  64873=>"001000111",
  64874=>"001001111",
  64875=>"000010110",
  64876=>"001010000",
  64877=>"011011101",
  64878=>"000000100",
  64879=>"000110110",
  64880=>"010100100",
  64881=>"001001110",
  64882=>"001110001",
  64883=>"111100111",
  64884=>"100011101",
  64885=>"111011010",
  64886=>"000100010",
  64887=>"110111011",
  64888=>"100110010",
  64889=>"001100001",
  64890=>"111110101",
  64891=>"111010101",
  64892=>"011000110",
  64893=>"011000110",
  64894=>"110001100",
  64895=>"001001011",
  64896=>"000010000",
  64897=>"110000111",
  64898=>"110010101",
  64899=>"000001011",
  64900=>"101100101",
  64901=>"111110110",
  64902=>"100111101",
  64903=>"111000010",
  64904=>"010110001",
  64905=>"111101011",
  64906=>"111101001",
  64907=>"011011100",
  64908=>"011000101",
  64909=>"101111100",
  64910=>"000001000",
  64911=>"110011000",
  64912=>"100111110",
  64913=>"000000001",
  64914=>"010001001",
  64915=>"000000110",
  64916=>"001011010",
  64917=>"100010101",
  64918=>"000000000",
  64919=>"010110000",
  64920=>"000000100",
  64921=>"000000001",
  64922=>"110000110",
  64923=>"010011001",
  64924=>"101001110",
  64925=>"101100101",
  64926=>"111111001",
  64927=>"111101010",
  64928=>"110001110",
  64929=>"111101010",
  64930=>"011011010",
  64931=>"001011111",
  64932=>"010111001",
  64933=>"111001100",
  64934=>"111011100",
  64935=>"010010101",
  64936=>"010010100",
  64937=>"101110101",
  64938=>"001100000",
  64939=>"001101011",
  64940=>"001111001",
  64941=>"100110000",
  64942=>"100001001",
  64943=>"111011001",
  64944=>"010000010",
  64945=>"000101000",
  64946=>"111111111",
  64947=>"101010011",
  64948=>"101101001",
  64949=>"000010001",
  64950=>"010001010",
  64951=>"001001100",
  64952=>"111010111",
  64953=>"101001010",
  64954=>"100100111",
  64955=>"100011100",
  64956=>"110100111",
  64957=>"011111111",
  64958=>"000011101",
  64959=>"010110111",
  64960=>"001111000",
  64961=>"100010010",
  64962=>"100000010",
  64963=>"111110101",
  64964=>"010110111",
  64965=>"011010110",
  64966=>"000011010",
  64967=>"111011000",
  64968=>"011011001",
  64969=>"000100110",
  64970=>"100010100",
  64971=>"110111101",
  64972=>"001100000",
  64973=>"001010001",
  64974=>"101010001",
  64975=>"101010011",
  64976=>"011101101",
  64977=>"011011101",
  64978=>"110111101",
  64979=>"000110100",
  64980=>"010000010",
  64981=>"010100001",
  64982=>"101000111",
  64983=>"110111010",
  64984=>"101100011",
  64985=>"110010001",
  64986=>"111110101",
  64987=>"101101011",
  64988=>"111101000",
  64989=>"111000111",
  64990=>"010101101",
  64991=>"111111011",
  64992=>"010001110",
  64993=>"011010011",
  64994=>"111111000",
  64995=>"111110101",
  64996=>"101010110",
  64997=>"011111101",
  64998=>"000000101",
  64999=>"001001100",
  65000=>"100111111",
  65001=>"001100001",
  65002=>"000010000",
  65003=>"001101010",
  65004=>"000111011",
  65005=>"110000000",
  65006=>"111001101",
  65007=>"101101111",
  65008=>"000010000",
  65009=>"110100011",
  65010=>"011001010",
  65011=>"000110100",
  65012=>"101000011",
  65013=>"101101011",
  65014=>"010101101",
  65015=>"001010100",
  65016=>"011000000",
  65017=>"110010101",
  65018=>"011011001",
  65019=>"001101111",
  65020=>"010101111",
  65021=>"001011111",
  65022=>"100000111",
  65023=>"110001010",
  65024=>"011000001",
  65025=>"101111100",
  65026=>"101100100",
  65027=>"110101100",
  65028=>"100001010",
  65029=>"010001101",
  65030=>"100011010",
  65031=>"011000110",
  65032=>"000001100",
  65033=>"010010010",
  65034=>"001010111",
  65035=>"100010010",
  65036=>"101010010",
  65037=>"100000001",
  65038=>"111010011",
  65039=>"111010000",
  65040=>"110110011",
  65041=>"110001000",
  65042=>"011011101",
  65043=>"101011110",
  65044=>"111001000",
  65045=>"010010001",
  65046=>"001100110",
  65047=>"101100111",
  65048=>"010001101",
  65049=>"111110110",
  65050=>"100011000",
  65051=>"101101111",
  65052=>"110001010",
  65053=>"010101110",
  65054=>"100100011",
  65055=>"011100100",
  65056=>"001111000",
  65057=>"101010010",
  65058=>"000001101",
  65059=>"000111011",
  65060=>"011000010",
  65061=>"010100111",
  65062=>"110110011",
  65063=>"011100111",
  65064=>"010000000",
  65065=>"100011010",
  65066=>"111011010",
  65067=>"110110111",
  65068=>"001111101",
  65069=>"000100101",
  65070=>"001000111",
  65071=>"011011001",
  65072=>"010110000",
  65073=>"001010110",
  65074=>"110101011",
  65075=>"010111001",
  65076=>"110010111",
  65077=>"001001100",
  65078=>"011010010",
  65079=>"110100111",
  65080=>"011011000",
  65081=>"100101100",
  65082=>"001001010",
  65083=>"010001101",
  65084=>"001100100",
  65085=>"010100101",
  65086=>"011101101",
  65087=>"100000101",
  65088=>"011001101",
  65089=>"011000000",
  65090=>"101101100",
  65091=>"001111111",
  65092=>"000011001",
  65093=>"001110100",
  65094=>"010111010",
  65095=>"100111100",
  65096=>"111001001",
  65097=>"111111100",
  65098=>"010111111",
  65099=>"100101110",
  65100=>"010000001",
  65101=>"111001000",
  65102=>"000011000",
  65103=>"011010111",
  65104=>"110011100",
  65105=>"110010001",
  65106=>"000010110",
  65107=>"001010000",
  65108=>"000011101",
  65109=>"001010011",
  65110=>"101111001",
  65111=>"111010001",
  65112=>"111100101",
  65113=>"101110000",
  65114=>"011010010",
  65115=>"010111111",
  65116=>"101101010",
  65117=>"110100000",
  65118=>"001101101",
  65119=>"110011100",
  65120=>"001011101",
  65121=>"011001010",
  65122=>"011000110",
  65123=>"011011001",
  65124=>"100011000",
  65125=>"001011011",
  65126=>"010101111",
  65127=>"100001000",
  65128=>"000001011",
  65129=>"111001101",
  65130=>"011001110",
  65131=>"001001100",
  65132=>"110010001",
  65133=>"111101000",
  65134=>"001001010",
  65135=>"001001110",
  65136=>"001110000",
  65137=>"001010010",
  65138=>"000001010",
  65139=>"011110111",
  65140=>"100001010",
  65141=>"010010000",
  65142=>"110100100",
  65143=>"111001110",
  65144=>"111010000",
  65145=>"011110001",
  65146=>"111011100",
  65147=>"111110111",
  65148=>"011001010",
  65149=>"101001010",
  65150=>"101100001",
  65151=>"110010000",
  65152=>"000101111",
  65153=>"000101011",
  65154=>"000011101",
  65155=>"111101010",
  65156=>"100110010",
  65157=>"100100010",
  65158=>"110000000",
  65159=>"110001111",
  65160=>"010011110",
  65161=>"110111000",
  65162=>"000001010",
  65163=>"110100101",
  65164=>"011100100",
  65165=>"000000111",
  65166=>"101010000",
  65167=>"000010100",
  65168=>"011001110",
  65169=>"011001111",
  65170=>"110001100",
  65171=>"100010110",
  65172=>"101110111",
  65173=>"110110010",
  65174=>"101001000",
  65175=>"101110110",
  65176=>"101100010",
  65177=>"110011111",
  65178=>"101011110",
  65179=>"001000011",
  65180=>"111110100",
  65181=>"111110101",
  65182=>"000101101",
  65183=>"000111111",
  65184=>"011011011",
  65185=>"001011100",
  65186=>"000100010",
  65187=>"011001011",
  65188=>"110101101",
  65189=>"011101110",
  65190=>"011101101",
  65191=>"000100111",
  65192=>"001111111",
  65193=>"100110100",
  65194=>"000001111",
  65195=>"111000100",
  65196=>"011010000",
  65197=>"101011110",
  65198=>"000001000",
  65199=>"000010111",
  65200=>"000010110",
  65201=>"101000010",
  65202=>"010011100",
  65203=>"011001001",
  65204=>"100100101",
  65205=>"110011111",
  65206=>"111111111",
  65207=>"000110110",
  65208=>"101000000",
  65209=>"011110101",
  65210=>"101111111",
  65211=>"010110011",
  65212=>"101001000",
  65213=>"011001101",
  65214=>"011011010",
  65215=>"100111001",
  65216=>"001101000",
  65217=>"000110110",
  65218=>"000000010",
  65219=>"111100010",
  65220=>"000100101",
  65221=>"101110100",
  65222=>"011111001",
  65223=>"101111000",
  65224=>"110000000",
  65225=>"010000011",
  65226=>"000000110",
  65227=>"101010001",
  65228=>"100000110",
  65229=>"000101111",
  65230=>"001011001",
  65231=>"011001010",
  65232=>"110100000",
  65233=>"101000010",
  65234=>"100010011",
  65235=>"000111110",
  65236=>"011111100",
  65237=>"100000011",
  65238=>"001000011",
  65239=>"111011110",
  65240=>"101100000",
  65241=>"010000101",
  65242=>"111110010",
  65243=>"011011010",
  65244=>"010000101",
  65245=>"111111010",
  65246=>"000001100",
  65247=>"100111001",
  65248=>"100001001",
  65249=>"010010000",
  65250=>"111010110",
  65251=>"000010000",
  65252=>"010011000",
  65253=>"111101110",
  65254=>"001010100",
  65255=>"000110111",
  65256=>"000011110",
  65257=>"000101110",
  65258=>"110111111",
  65259=>"001001000",
  65260=>"111000001",
  65261=>"101010101",
  65262=>"001000100",
  65263=>"010001111",
  65264=>"010111010",
  65265=>"101111010",
  65266=>"001001010",
  65267=>"011011110",
  65268=>"001110001",
  65269=>"001000110",
  65270=>"010101100",
  65271=>"100110101",
  65272=>"111110011",
  65273=>"000110110",
  65274=>"011110101",
  65275=>"110101011",
  65276=>"100101111",
  65277=>"000111101",
  65278=>"101101110",
  65279=>"100000010",
  65280=>"010101010",
  65281=>"111010010",
  65282=>"000000111",
  65283=>"001100101",
  65284=>"101000010",
  65285=>"000001000",
  65286=>"011101010",
  65287=>"111100001",
  65288=>"000001000",
  65289=>"010010000",
  65290=>"010111000",
  65291=>"111010001",
  65292=>"011110010",
  65293=>"010100010",
  65294=>"100011101",
  65295=>"000111100",
  65296=>"000011111",
  65297=>"000000011",
  65298=>"010011111",
  65299=>"110010100",
  65300=>"001101110",
  65301=>"101101011",
  65302=>"001110100",
  65303=>"111111100",
  65304=>"001001000",
  65305=>"001100100",
  65306=>"100011101",
  65307=>"110110101",
  65308=>"001100100",
  65309=>"110110111",
  65310=>"110001001",
  65311=>"100110001",
  65312=>"110110001",
  65313=>"100110111",
  65314=>"100001100",
  65315=>"100100111",
  65316=>"100110011",
  65317=>"101010011",
  65318=>"001010110",
  65319=>"010101001",
  65320=>"000010010",
  65321=>"111000110",
  65322=>"011110001",
  65323=>"111010111",
  65324=>"000011010",
  65325=>"001000001",
  65326=>"000001000",
  65327=>"100000101",
  65328=>"000001010",
  65329=>"101110100",
  65330=>"011101111",
  65331=>"110100111",
  65332=>"001101110",
  65333=>"101110001",
  65334=>"000110100",
  65335=>"000111101",
  65336=>"010101001",
  65337=>"111011001",
  65338=>"000100101",
  65339=>"111011000",
  65340=>"011101111",
  65341=>"111000010",
  65342=>"111001001",
  65343=>"000001101",
  65344=>"100011000",
  65345=>"010110111",
  65346=>"100000011",
  65347=>"000100110",
  65348=>"111100001",
  65349=>"011101111",
  65350=>"011000000",
  65351=>"000110011",
  65352=>"111011110",
  65353=>"001001111",
  65354=>"100001011",
  65355=>"110000000",
  65356=>"001010011",
  65357=>"100110100",
  65358=>"110010010",
  65359=>"101000111",
  65360=>"001101011",
  65361=>"111100000",
  65362=>"000000001",
  65363=>"101101001",
  65364=>"001111110",
  65365=>"011111101",
  65366=>"010110001",
  65367=>"011010011",
  65368=>"010100010",
  65369=>"110110110",
  65370=>"000100000",
  65371=>"010001110",
  65372=>"010110011",
  65373=>"100111000",
  65374=>"111000011",
  65375=>"000000000",
  65376=>"110110000",
  65377=>"011010111",
  65378=>"010001111",
  65379=>"100001000",
  65380=>"101001110",
  65381=>"110110010",
  65382=>"101100110",
  65383=>"100101100",
  65384=>"001111111",
  65385=>"110111011",
  65386=>"100100010",
  65387=>"011111110",
  65388=>"101010111",
  65389=>"110100000",
  65390=>"010111100",
  65391=>"110010010",
  65392=>"111001000",
  65393=>"100011011",
  65394=>"010000001",
  65395=>"101110101",
  65396=>"001000101",
  65397=>"111110001",
  65398=>"010000100",
  65399=>"010101111",
  65400=>"110100001",
  65401=>"000100001",
  65402=>"101101001",
  65403=>"001100001",
  65404=>"001011000",
  65405=>"110001000",
  65406=>"111110011",
  65407=>"111000000",
  65408=>"111111000",
  65409=>"001010010",
  65410=>"111001111",
  65411=>"010010000",
  65412=>"110100110",
  65413=>"100110100",
  65414=>"010001110",
  65415=>"111101000",
  65416=>"011011101",
  65417=>"011000101",
  65418=>"010110110",
  65419=>"111101110",
  65420=>"110110000",
  65421=>"010000111",
  65422=>"111010100",
  65423=>"000001100",
  65424=>"101001111",
  65425=>"101100000",
  65426=>"101111001",
  65427=>"111111001",
  65428=>"110111001",
  65429=>"111001101",
  65430=>"101111001",
  65431=>"111000011",
  65432=>"100101001",
  65433=>"111000011",
  65434=>"010011010",
  65435=>"000010100",
  65436=>"010000001",
  65437=>"000000000",
  65438=>"001010001",
  65439=>"110001100",
  65440=>"001111010",
  65441=>"101111101",
  65442=>"111101111",
  65443=>"101000110",
  65444=>"101010100",
  65445=>"001110111",
  65446=>"010110100",
  65447=>"100010010",
  65448=>"011100100",
  65449=>"011011101",
  65450=>"111011101",
  65451=>"100100000",
  65452=>"110011101",
  65453=>"000100000",
  65454=>"110010100",
  65455=>"100010000",
  65456=>"011101010",
  65457=>"001001010",
  65458=>"001101001",
  65459=>"111111011",
  65460=>"011100000",
  65461=>"111000010",
  65462=>"101110000",
  65463=>"011101111",
  65464=>"000001000",
  65465=>"001000101",
  65466=>"000010000",
  65467=>"100100110",
  65468=>"111110110",
  65469=>"100111010",
  65470=>"111110000",
  65471=>"000010010",
  65472=>"000011111",
  65473=>"011110110",
  65474=>"111001011",
  65475=>"000110011",
  65476=>"000101011",
  65477=>"110100010",
  65478=>"010110010",
  65479=>"000101111",
  65480=>"001010111",
  65481=>"100000010",
  65482=>"100100000",
  65483=>"000100111",
  65484=>"011011110",
  65485=>"110000000",
  65486=>"011111110",
  65487=>"100001000",
  65488=>"001000001",
  65489=>"100111101",
  65490=>"010001010",
  65491=>"001111110",
  65492=>"010100000",
  65493=>"110010101",
  65494=>"010001010",
  65495=>"000001001",
  65496=>"100001111",
  65497=>"111010101",
  65498=>"111111000",
  65499=>"111111110",
  65500=>"000101101",
  65501=>"010100001",
  65502=>"110001010",
  65503=>"000110100",
  65504=>"100100010",
  65505=>"010011010",
  65506=>"101010001",
  65507=>"001101011",
  65508=>"111010010",
  65509=>"000010000",
  65510=>"100001001",
  65511=>"110000100",
  65512=>"011000000",
  65513=>"100010001",
  65514=>"110101011",
  65515=>"000011001",
  65516=>"111111101",
  65517=>"100111111",
  65518=>"100111101",
  65519=>"111111101",
  65520=>"011010000",
  65521=>"101110101",
  65522=>"101001010",
  65523=>"010101101",
  65524=>"000000010",
  65525=>"011001101",
  65526=>"100100100",
  65527=>"110000110",
  65528=>"010001101",
  65529=>"101010101",
  65530=>"001111001",
  65531=>"010100101",
  65532=>"001010101",
  65533=>"000100000",
  65534=>"001000000",
  65535=>"111100001");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;