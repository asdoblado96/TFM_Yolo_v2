LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_8_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_8_BNROM;

ARCHITECTURE RTL OF L8_8_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0000111011010101"&"0010011011010110",
  1=>"0000101100110101"&"0010100000101011",
  2=>"0001100011111111"&"0010010001100000",
  3=>"0001101100011010"&"0010010110110101",
  4=>"0001000101000000"&"0010000110100011",
  5=>"0001101110100101"&"0010010001101010",
  6=>"0000101001111011"&"0010001110111010",
  7=>"1111111100001000"&"0010001100101110",
  8=>"0010001001010111"&"0010001110010011",
  9=>"0000010110001101"&"0010000110011001",
  10=>"0001100101100010"&"0010011100111011",
  11=>"0000100000111110"&"0010000010110001",
  12=>"1110101110011011"&"0001100000110101",
  13=>"0010000100100001"&"0001111001110101",
  14=>"0000101110101110"&"0001110101110011",
  15=>"1111111111101101"&"0001111000110101",
  16=>"1111001011011111"&"0010000101110000",
  17=>"0001101111011000"&"0010001000110111",
  18=>"0010110001000000"&"0010000011010010",
  19=>"0001101000111011"&"0010010111001111",
  20=>"0000111011010010"&"0001111010000101",
  21=>"0001001110100011"&"0010010110010000",
  22=>"0000010000000100"&"0010010110100100",
  23=>"0000101011100000"&"0010011111011100",
  24=>"0001001010111011"&"0001101110001010",
  25=>"0000010111100110"&"0010001100011011",
  26=>"1111110111000000"&"0001100110001001",
  27=>"0000011011010011"&"0001111111001111",
  28=>"0001000001111011"&"0010011111011010",
  29=>"0001100100000001"&"0010010101001010",
  30=>"0000011101101010"&"0010001011011100",
  31=>"0000001101011010"&"0010100000101111",
  32=>"0001011100011101"&"0010001100001000",
  33=>"0001101100110001"&"0010010000010101",
  34=>"0001001001110100"&"0001111111011001",
  35=>"0000110111011101"&"0001011011100111",
  36=>"0000001001100001"&"0001011100010000",
  37=>"0000011110100010"&"0010001101100100",
  38=>"1111010001111000"&"0010000000010100",
  39=>"0011000011011101"&"0001110111001000",
  40=>"0000111101011010"&"0010001101000000",
  41=>"0000011000001011"&"0001111001111000",
  42=>"0000010110000111"&"0001110111101011",
  43=>"0001100010000010"&"0010011010010001",
  44=>"0000010100000100"&"0001101010110001",
  45=>"0000100011111100"&"0010011010001100",
  46=>"0010001110101110"&"0010010000101010",
  47=>"0001010000010100"&"0010010001000110",
  48=>"0001111111110010"&"0001111111100010",
  49=>"0001110011110000"&"0010011001110111",
  50=>"0001100010010101"&"0010000011100011",
  51=>"0001110100000001"&"0010001101111110",
  52=>"0001100001110100"&"0010001101111111",
  53=>"0001110101000110"&"0010001001110101",
  54=>"0000110111100101"&"0010001011011000",
  55=>"0000111101000011"&"0010000001110010",
  56=>"0010000001111011"&"0010010000101010",
  57=>"0001100101011001"&"0010011000011100",
  58=>"0000100100011110"&"0001111110001101",
  59=>"0001001011100000"&"0010001011011010",
  60=>"0001000111000101"&"0001110110110010",
  61=>"0001110101100001"&"0010010110110010",
  62=>"0001000011001101"&"0010010111100100",
  63=>"0001110011001100"&"0010000100000001");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;