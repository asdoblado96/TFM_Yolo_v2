LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_11_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_11_WROM;

ARCHITECTURE RTL OF L8_11_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"101011101",
  1=>"110000010",
  2=>"100110000",
  3=>"000100111",
  4=>"010000001",
  5=>"111001111",
  6=>"100101010",
  7=>"011010111",
  8=>"101000101",
  9=>"111011111",
  10=>"011000110",
  11=>"000100111",
  12=>"011101011",
  13=>"000010111",
  14=>"000011101",
  15=>"000100100",
  16=>"010001100",
  17=>"001111100",
  18=>"011001110",
  19=>"101001101",
  20=>"000101010",
  21=>"000000000",
  22=>"100001111",
  23=>"000000010",
  24=>"010010101",
  25=>"100001111",
  26=>"001100110",
  27=>"011010000",
  28=>"011011000",
  29=>"111111011",
  30=>"000110100",
  31=>"011001001",
  32=>"011010110",
  33=>"001000100",
  34=>"111111011",
  35=>"010101000",
  36=>"100100101",
  37=>"110101011",
  38=>"001000011",
  39=>"000111011",
  40=>"111000000",
  41=>"011010111",
  42=>"000000100",
  43=>"011011101",
  44=>"101100100",
  45=>"100000111",
  46=>"110111101",
  47=>"100111010",
  48=>"111011001",
  49=>"011000000",
  50=>"100010100",
  51=>"110111000",
  52=>"001010111",
  53=>"100110000",
  54=>"111101010",
  55=>"001100001",
  56=>"111011001",
  57=>"010100000",
  58=>"000100001",
  59=>"110001011",
  60=>"010001000",
  61=>"010111010",
  62=>"000001010",
  63=>"000000001",
  64=>"000011001",
  65=>"111100010",
  66=>"000000101",
  67=>"011010010",
  68=>"001111010",
  69=>"001001100",
  70=>"111001000",
  71=>"100100100",
  72=>"110110010",
  73=>"001100111",
  74=>"011100110",
  75=>"100000011",
  76=>"011011000",
  77=>"101001011",
  78=>"011000011",
  79=>"111010100",
  80=>"101101100",
  81=>"000001100",
  82=>"011011100",
  83=>"011000110",
  84=>"111110111",
  85=>"110011001",
  86=>"100000010",
  87=>"111000111",
  88=>"011110010",
  89=>"101011001",
  90=>"001111011",
  91=>"001001000",
  92=>"100100100",
  93=>"010011111",
  94=>"000011000",
  95=>"001100011",
  96=>"100101011",
  97=>"001111101",
  98=>"011110111",
  99=>"010100000",
  100=>"100111010",
  101=>"010100000",
  102=>"011111010",
  103=>"110011111",
  104=>"100011100",
  105=>"100100111",
  106=>"001000100",
  107=>"001000100",
  108=>"010111101",
  109=>"101101000",
  110=>"111000110",
  111=>"111100100",
  112=>"011011110",
  113=>"101000101",
  114=>"000110010",
  115=>"000010000",
  116=>"011010110",
  117=>"011011001",
  118=>"000100111",
  119=>"111011001",
  120=>"000111011",
  121=>"010101000",
  122=>"010010000",
  123=>"100011101",
  124=>"110010001",
  125=>"110011011",
  126=>"111110001",
  127=>"000110000",
  128=>"000011000",
  129=>"010010110",
  130=>"011101001",
  131=>"001010000",
  132=>"010100000",
  133=>"110110011",
  134=>"001110110",
  135=>"001100110",
  136=>"010000110",
  137=>"000010111",
  138=>"000000011",
  139=>"110100101",
  140=>"001010011",
  141=>"001111000",
  142=>"110001101",
  143=>"000100111",
  144=>"111010111",
  145=>"101111011",
  146=>"100110101",
  147=>"011100110",
  148=>"011001011",
  149=>"100101010",
  150=>"011111110",
  151=>"001011001",
  152=>"100001100",
  153=>"100010111",
  154=>"011011011",
  155=>"111111001",
  156=>"011001101",
  157=>"101100000",
  158=>"011010000",
  159=>"101001110",
  160=>"111000111",
  161=>"000110011",
  162=>"110101110",
  163=>"111111111",
  164=>"011111011",
  165=>"100111110",
  166=>"000111100",
  167=>"100101001",
  168=>"011101001",
  169=>"111110100",
  170=>"110111001",
  171=>"010111001",
  172=>"011001100",
  173=>"001010011",
  174=>"011110010",
  175=>"101100100",
  176=>"001001001",
  177=>"100000001",
  178=>"100011110",
  179=>"101000001",
  180=>"000100000",
  181=>"010111010",
  182=>"010001111",
  183=>"110111111",
  184=>"010110011",
  185=>"101100011",
  186=>"100100110",
  187=>"111000001",
  188=>"101101011",
  189=>"010110010",
  190=>"010101010",
  191=>"111001111",
  192=>"111001011",
  193=>"000111101",
  194=>"110100010",
  195=>"100011001",
  196=>"001010001",
  197=>"100011000",
  198=>"001100110",
  199=>"101101000",
  200=>"001011111",
  201=>"001110100",
  202=>"000110000",
  203=>"000111100",
  204=>"110010101",
  205=>"001001101",
  206=>"111010110",
  207=>"000101101",
  208=>"101000000",
  209=>"011110100",
  210=>"010111101",
  211=>"101010110",
  212=>"011101000",
  213=>"110000010",
  214=>"110000001",
  215=>"101101011",
  216=>"001011111",
  217=>"101110101",
  218=>"010101111",
  219=>"001100011",
  220=>"011011101",
  221=>"010011100",
  222=>"011010111",
  223=>"110111100",
  224=>"001000000",
  225=>"111111101",
  226=>"100011001",
  227=>"001001000",
  228=>"111111111",
  229=>"111001111",
  230=>"100100010",
  231=>"011011010",
  232=>"110010100",
  233=>"100000111",
  234=>"100101111",
  235=>"000110101",
  236=>"011111010",
  237=>"001101101",
  238=>"100100011",
  239=>"111111110",
  240=>"100100011",
  241=>"011001010",
  242=>"101011011",
  243=>"101111000",
  244=>"111100101",
  245=>"110111100",
  246=>"001110011",
  247=>"010001010",
  248=>"110000111",
  249=>"100010100",
  250=>"101101111",
  251=>"110011010",
  252=>"000001000",
  253=>"000001110",
  254=>"010110110",
  255=>"100011001",
  256=>"100000111",
  257=>"001100110",
  258=>"010110111",
  259=>"100000101",
  260=>"010100011",
  261=>"110110101",
  262=>"001011001",
  263=>"101001010",
  264=>"100011111",
  265=>"100100000",
  266=>"101000000",
  267=>"010000001",
  268=>"010110100",
  269=>"001100010",
  270=>"010111000",
  271=>"000000001",
  272=>"000000000",
  273=>"010001011",
  274=>"011000100",
  275=>"101110111",
  276=>"101101100",
  277=>"110100100",
  278=>"111111000",
  279=>"110010000",
  280=>"101011001",
  281=>"110101101",
  282=>"001110100",
  283=>"000101110",
  284=>"001011010",
  285=>"000000000",
  286=>"000101000",
  287=>"000001010",
  288=>"110110001",
  289=>"100100010",
  290=>"001001110",
  291=>"011110100",
  292=>"110101101",
  293=>"001000110",
  294=>"000110001",
  295=>"110111110",
  296=>"000010100",
  297=>"101011101",
  298=>"111111110",
  299=>"011000101",
  300=>"001000111",
  301=>"100011000",
  302=>"101001111",
  303=>"100110010",
  304=>"001001011",
  305=>"110010011",
  306=>"101001110",
  307=>"000111010",
  308=>"011011000",
  309=>"111001111",
  310=>"111011100",
  311=>"011111001",
  312=>"100100111",
  313=>"000101001",
  314=>"101000010",
  315=>"010111111",
  316=>"000111011",
  317=>"010110111",
  318=>"111010010",
  319=>"101010111",
  320=>"110011111",
  321=>"110010011",
  322=>"001010000",
  323=>"000011001",
  324=>"010110001",
  325=>"001011101",
  326=>"000001001",
  327=>"110001011",
  328=>"000001110",
  329=>"001001000",
  330=>"001111111",
  331=>"111001101",
  332=>"011101010",
  333=>"001101000",
  334=>"000100010",
  335=>"011011110",
  336=>"111101110",
  337=>"000100101",
  338=>"010101011",
  339=>"101000011",
  340=>"100000101",
  341=>"001101111",
  342=>"010000000",
  343=>"111011001",
  344=>"101101000",
  345=>"111010111",
  346=>"101101100",
  347=>"011101010",
  348=>"110111011",
  349=>"100001001",
  350=>"110001100",
  351=>"110001110",
  352=>"100011110",
  353=>"010010011",
  354=>"011000111",
  355=>"010111000",
  356=>"011001101",
  357=>"011100010",
  358=>"100000100",
  359=>"110010010",
  360=>"100000101",
  361=>"001111110",
  362=>"101001000",
  363=>"000000111",
  364=>"001010100",
  365=>"011111011",
  366=>"100010001",
  367=>"101010011",
  368=>"100011111",
  369=>"100101101",
  370=>"110001010",
  371=>"001011011",
  372=>"000000101",
  373=>"100110000",
  374=>"110110001",
  375=>"011100101",
  376=>"001011100",
  377=>"100001011",
  378=>"010000110",
  379=>"110000110",
  380=>"000001101",
  381=>"011001001",
  382=>"111111111",
  383=>"010011101",
  384=>"111100000",
  385=>"001111000",
  386=>"100111111",
  387=>"011011101",
  388=>"111111110",
  389=>"001000111",
  390=>"010000001",
  391=>"100011011",
  392=>"110011001",
  393=>"011101001",
  394=>"001000001",
  395=>"000001011",
  396=>"011100110",
  397=>"010101011",
  398=>"100011011",
  399=>"001100100",
  400=>"010110011",
  401=>"000000010",
  402=>"101111110",
  403=>"100000010",
  404=>"101001100",
  405=>"100001100",
  406=>"111111011",
  407=>"110110010",
  408=>"100001000",
  409=>"011001000",
  410=>"000100111",
  411=>"111001100",
  412=>"110101001",
  413=>"010011101",
  414=>"011010101",
  415=>"011100001",
  416=>"111010001",
  417=>"001101111",
  418=>"101110010",
  419=>"100010000",
  420=>"010100100",
  421=>"110110000",
  422=>"110000010",
  423=>"010100110",
  424=>"111010111",
  425=>"100011010",
  426=>"110100111",
  427=>"100101011",
  428=>"001001101",
  429=>"011101101",
  430=>"011001010",
  431=>"011000100",
  432=>"001001000",
  433=>"000101000",
  434=>"010011011",
  435=>"111111101",
  436=>"000100111",
  437=>"101000011",
  438=>"011101100",
  439=>"110101001",
  440=>"001011100",
  441=>"000001101",
  442=>"111100110",
  443=>"100010010",
  444=>"010010001",
  445=>"111011100",
  446=>"100111000",
  447=>"000100100",
  448=>"010000001",
  449=>"101101010",
  450=>"001111000",
  451=>"001110110",
  452=>"111110010",
  453=>"101000011",
  454=>"100000110",
  455=>"010000000",
  456=>"101001011",
  457=>"111101110",
  458=>"100101010",
  459=>"000110011",
  460=>"000011100",
  461=>"111010101",
  462=>"000011100",
  463=>"010110111",
  464=>"111111110",
  465=>"100011101",
  466=>"100101111",
  467=>"010010111",
  468=>"101101001",
  469=>"001011010",
  470=>"110111111",
  471=>"010100011",
  472=>"000110010",
  473=>"011110100",
  474=>"101011001",
  475=>"111010111",
  476=>"000010001",
  477=>"110001010",
  478=>"100010000",
  479=>"011100011",
  480=>"000110011",
  481=>"100110000",
  482=>"000010000",
  483=>"000000000",
  484=>"100000001",
  485=>"101100111",
  486=>"110110101",
  487=>"010001010",
  488=>"010100101",
  489=>"100100110",
  490=>"010000001",
  491=>"001011001",
  492=>"100001111",
  493=>"011011111",
  494=>"110111101",
  495=>"000000001",
  496=>"000101111",
  497=>"111110001",
  498=>"111100000",
  499=>"110010110",
  500=>"010001100",
  501=>"100111000",
  502=>"001111101",
  503=>"110100100",
  504=>"111000111",
  505=>"011100101",
  506=>"100011101",
  507=>"001111010",
  508=>"111101111",
  509=>"011001000",
  510=>"011011011",
  511=>"110110100",
  512=>"010100100",
  513=>"101010010",
  514=>"111010110",
  515=>"000000100",
  516=>"111011100",
  517=>"000001011",
  518=>"101101010",
  519=>"011111011",
  520=>"011000100",
  521=>"100001110",
  522=>"100111011",
  523=>"000110100",
  524=>"101010000",
  525=>"010001011",
  526=>"000100111",
  527=>"110010011",
  528=>"001111011",
  529=>"101011001",
  530=>"010110011",
  531=>"011000101",
  532=>"101001100",
  533=>"001101100",
  534=>"100101000",
  535=>"000110010",
  536=>"000001010",
  537=>"000010001",
  538=>"000000010",
  539=>"010101111",
  540=>"111101011",
  541=>"001010101",
  542=>"110000011",
  543=>"110100010",
  544=>"010011011",
  545=>"000101000",
  546=>"011000011",
  547=>"001000000",
  548=>"111010011",
  549=>"010011011",
  550=>"110000010",
  551=>"101111110",
  552=>"101101111",
  553=>"110000110",
  554=>"101000000",
  555=>"110110111",
  556=>"100000100",
  557=>"110010000",
  558=>"111101101",
  559=>"000111000",
  560=>"011111001",
  561=>"011100011",
  562=>"011010111",
  563=>"001001101",
  564=>"001110100",
  565=>"000101101",
  566=>"111101110",
  567=>"100000000",
  568=>"011110010",
  569=>"000000110",
  570=>"111110010",
  571=>"101011111",
  572=>"010111111",
  573=>"000100111",
  574=>"000110011",
  575=>"011100100",
  576=>"000011110",
  577=>"001000101",
  578=>"100110000",
  579=>"100110010",
  580=>"001001000",
  581=>"010110010",
  582=>"101011110",
  583=>"100100100",
  584=>"111110010",
  585=>"001000110",
  586=>"101010010",
  587=>"111000101",
  588=>"001111011",
  589=>"110000000",
  590=>"101010110",
  591=>"011000110",
  592=>"101111000",
  593=>"001101101",
  594=>"000100111",
  595=>"101101110",
  596=>"010101111",
  597=>"000010011",
  598=>"100000001",
  599=>"100110110",
  600=>"100011001",
  601=>"111001010",
  602=>"111111100",
  603=>"101010000",
  604=>"010001110",
  605=>"110000111",
  606=>"011110110",
  607=>"100100000",
  608=>"000011110",
  609=>"010000011",
  610=>"011000100",
  611=>"110010000",
  612=>"010001101",
  613=>"111111100",
  614=>"011100100",
  615=>"011010001",
  616=>"000010110",
  617=>"000110110",
  618=>"011111011",
  619=>"101001001",
  620=>"000110010",
  621=>"001100111",
  622=>"011101001",
  623=>"000100111",
  624=>"110100011",
  625=>"100100000",
  626=>"001100110",
  627=>"000110000",
  628=>"101010100",
  629=>"110011111",
  630=>"010110011",
  631=>"011101010",
  632=>"101001010",
  633=>"001011010",
  634=>"011010100",
  635=>"010101000",
  636=>"110001010",
  637=>"111100111",
  638=>"110011001",
  639=>"110010001",
  640=>"100000100",
  641=>"110101101",
  642=>"010011111",
  643=>"001001000",
  644=>"110111001",
  645=>"100001101",
  646=>"000000101",
  647=>"101110000",
  648=>"110111100",
  649=>"110001111",
  650=>"111100001",
  651=>"100111001",
  652=>"101110011",
  653=>"100101111",
  654=>"101010111",
  655=>"110010110",
  656=>"010000001",
  657=>"111100110",
  658=>"111111110",
  659=>"011000001",
  660=>"001110101",
  661=>"011010111",
  662=>"110110110",
  663=>"100000001",
  664=>"100100011",
  665=>"101010110",
  666=>"101010101",
  667=>"010001001",
  668=>"000011111",
  669=>"010000001",
  670=>"110011110",
  671=>"010101010",
  672=>"100011011",
  673=>"110101110",
  674=>"101000001",
  675=>"000001010",
  676=>"101001111",
  677=>"111111011",
  678=>"100001100",
  679=>"111100000",
  680=>"010000111",
  681=>"000000000",
  682=>"000010010",
  683=>"100001001",
  684=>"000001010",
  685=>"001010001",
  686=>"000101110",
  687=>"100111010",
  688=>"000011110",
  689=>"110100011",
  690=>"100100110",
  691=>"011011100",
  692=>"010010000",
  693=>"011110000",
  694=>"111001011",
  695=>"001000100",
  696=>"110111110",
  697=>"111001111",
  698=>"101001111",
  699=>"000000101",
  700=>"010110111",
  701=>"011001010",
  702=>"101000101",
  703=>"001111010",
  704=>"000110111",
  705=>"010110111",
  706=>"100011001",
  707=>"100001100",
  708=>"011101111",
  709=>"010111100",
  710=>"001001010",
  711=>"000011011",
  712=>"000000001",
  713=>"111010110",
  714=>"001000111",
  715=>"010000111",
  716=>"001100100",
  717=>"000011010",
  718=>"111101110",
  719=>"010110011",
  720=>"111110000",
  721=>"001111101",
  722=>"101110000",
  723=>"111010010",
  724=>"110101101",
  725=>"010100001",
  726=>"100110000",
  727=>"100011101",
  728=>"010110011",
  729=>"001000111",
  730=>"010000110",
  731=>"000110110",
  732=>"101110010",
  733=>"010001011",
  734=>"011101100",
  735=>"111011101",
  736=>"101011000",
  737=>"101111011",
  738=>"000001101",
  739=>"100110101",
  740=>"001010001",
  741=>"111101101",
  742=>"000100010",
  743=>"000011001",
  744=>"000010000",
  745=>"001001000",
  746=>"111011000",
  747=>"001111011",
  748=>"100111111",
  749=>"111101100",
  750=>"001100001",
  751=>"111010001",
  752=>"001010000",
  753=>"011100101",
  754=>"111101000",
  755=>"010100100",
  756=>"101010110",
  757=>"011100111",
  758=>"011010110",
  759=>"001010110",
  760=>"011110000",
  761=>"110011111",
  762=>"000100000",
  763=>"001001000",
  764=>"111100100",
  765=>"101111101",
  766=>"111101101",
  767=>"000001000",
  768=>"010000000",
  769=>"100110111",
  770=>"010110011",
  771=>"011001010",
  772=>"100001111",
  773=>"100001111",
  774=>"100101000",
  775=>"010110011",
  776=>"101101110",
  777=>"100000110",
  778=>"101111111",
  779=>"001111000",
  780=>"010001000",
  781=>"001110100",
  782=>"001001100",
  783=>"000001000",
  784=>"001011011",
  785=>"011110010",
  786=>"110111011",
  787=>"011011111",
  788=>"100000000",
  789=>"010111110",
  790=>"111111100",
  791=>"100111001",
  792=>"010010011",
  793=>"011100010",
  794=>"110010110",
  795=>"100111001",
  796=>"010011100",
  797=>"101001010",
  798=>"000010111",
  799=>"111110100",
  800=>"110000100",
  801=>"001101001",
  802=>"001010010",
  803=>"100101000",
  804=>"101101001",
  805=>"010001110",
  806=>"011110110",
  807=>"111001000",
  808=>"111000101",
  809=>"100101111",
  810=>"111010001",
  811=>"101001001",
  812=>"111011000",
  813=>"010100001",
  814=>"101000110",
  815=>"001110110",
  816=>"111101100",
  817=>"101101100",
  818=>"010010001",
  819=>"100111111",
  820=>"011000001",
  821=>"001001010",
  822=>"111000000",
  823=>"111100010",
  824=>"110111101",
  825=>"011100111",
  826=>"000010001",
  827=>"110110111",
  828=>"010001010",
  829=>"000010110",
  830=>"011101111",
  831=>"110101011",
  832=>"111000010",
  833=>"111011000",
  834=>"110010111",
  835=>"111011011",
  836=>"101100110",
  837=>"010110110",
  838=>"011101001",
  839=>"111101100",
  840=>"110101000",
  841=>"001000010",
  842=>"101110111",
  843=>"101111010",
  844=>"010101001",
  845=>"011011111",
  846=>"010010000",
  847=>"010000110",
  848=>"001000100",
  849=>"111101100",
  850=>"001111011",
  851=>"000001100",
  852=>"101010101",
  853=>"001110011",
  854=>"110101111",
  855=>"000100111",
  856=>"011110010",
  857=>"100010000",
  858=>"101110111",
  859=>"000001001",
  860=>"110100000",
  861=>"111110100",
  862=>"111001110",
  863=>"001110001",
  864=>"100010011",
  865=>"000010000",
  866=>"111110111",
  867=>"101101000",
  868=>"001010010",
  869=>"011010100",
  870=>"101110010",
  871=>"111010001",
  872=>"101100011",
  873=>"010010001",
  874=>"010110101",
  875=>"101010111",
  876=>"001010101",
  877=>"101110010",
  878=>"000011011",
  879=>"010001110",
  880=>"011001101",
  881=>"100110011",
  882=>"011101000",
  883=>"101100001",
  884=>"011111110",
  885=>"010010111",
  886=>"010110000",
  887=>"101001101",
  888=>"000000000",
  889=>"101010111",
  890=>"100010101",
  891=>"101001010",
  892=>"000000000",
  893=>"100110110",
  894=>"000101101",
  895=>"010100010",
  896=>"100010001",
  897=>"110111110",
  898=>"111110011",
  899=>"010101110",
  900=>"100110001",
  901=>"101110001",
  902=>"110000111",
  903=>"010010100",
  904=>"100101100",
  905=>"110011110",
  906=>"001110000",
  907=>"101110011",
  908=>"101001110",
  909=>"010111010",
  910=>"011000011",
  911=>"001111100",
  912=>"011100110",
  913=>"001010011",
  914=>"000000111",
  915=>"011111010",
  916=>"110101100",
  917=>"000100001",
  918=>"110001011",
  919=>"010001101",
  920=>"000100110",
  921=>"010100111",
  922=>"000001000",
  923=>"001011000",
  924=>"000111111",
  925=>"010100011",
  926=>"010100111",
  927=>"110000101",
  928=>"111001001",
  929=>"000101000",
  930=>"000110000",
  931=>"111101011",
  932=>"001001000",
  933=>"100100010",
  934=>"010111010",
  935=>"111001101",
  936=>"010110111",
  937=>"010111101",
  938=>"101011111",
  939=>"010010001",
  940=>"100110000",
  941=>"000111010",
  942=>"100000011",
  943=>"111011100",
  944=>"110100011",
  945=>"101011101",
  946=>"100011100",
  947=>"101011110",
  948=>"100000101",
  949=>"111110010",
  950=>"111001011",
  951=>"111001001",
  952=>"110100100",
  953=>"001101000",
  954=>"011011111",
  955=>"101110111",
  956=>"001000010",
  957=>"001010010",
  958=>"110001110",
  959=>"010110100",
  960=>"100111010",
  961=>"000010110",
  962=>"110001001",
  963=>"010011010",
  964=>"010110111",
  965=>"001101010",
  966=>"010100001",
  967=>"111000001",
  968=>"001000001",
  969=>"010011110",
  970=>"111100111",
  971=>"111001000",
  972=>"101110110",
  973=>"000100010",
  974=>"101000000",
  975=>"110000101",
  976=>"011110110",
  977=>"100011101",
  978=>"111110110",
  979=>"011100010",
  980=>"011111101",
  981=>"011010111",
  982=>"110010110",
  983=>"111001101",
  984=>"010000111",
  985=>"001110010",
  986=>"000000101",
  987=>"000111110",
  988=>"111011111",
  989=>"011000100",
  990=>"001010011",
  991=>"000001010",
  992=>"010111001",
  993=>"010000111",
  994=>"110111000",
  995=>"110111111",
  996=>"001011000",
  997=>"111111011",
  998=>"111111001",
  999=>"110101101",
  1000=>"011000000",
  1001=>"100101101",
  1002=>"001111000",
  1003=>"100000111",
  1004=>"000000010",
  1005=>"000111100",
  1006=>"000100001",
  1007=>"101110111",
  1008=>"001000001",
  1009=>"110011001",
  1010=>"110101111",
  1011=>"100001010",
  1012=>"010000001",
  1013=>"111000100",
  1014=>"011100010",
  1015=>"111000011",
  1016=>"011000111",
  1017=>"011100111",
  1018=>"100000101",
  1019=>"000010110",
  1020=>"010111101",
  1021=>"100001101",
  1022=>"101000000",
  1023=>"011011010",
  1024=>"000111110",
  1025=>"010001010",
  1026=>"111110110",
  1027=>"111011111",
  1028=>"000001010",
  1029=>"110001000",
  1030=>"100111010",
  1031=>"001111011",
  1032=>"010000111",
  1033=>"001110101",
  1034=>"000111001",
  1035=>"010111000",
  1036=>"011101111",
  1037=>"111111100",
  1038=>"111000011",
  1039=>"001001101",
  1040=>"110011001",
  1041=>"100011110",
  1042=>"100100000",
  1043=>"100100110",
  1044=>"101001101",
  1045=>"100110111",
  1046=>"111010100",
  1047=>"001001011",
  1048=>"100010110",
  1049=>"001100000",
  1050=>"110110100",
  1051=>"111100110",
  1052=>"001011101",
  1053=>"001001001",
  1054=>"011010000",
  1055=>"100100001",
  1056=>"000101101",
  1057=>"100011111",
  1058=>"001110100",
  1059=>"011001100",
  1060=>"101111110",
  1061=>"110110100",
  1062=>"101101110",
  1063=>"101001010",
  1064=>"010111101",
  1065=>"000000100",
  1066=>"101011111",
  1067=>"101011110",
  1068=>"010010001",
  1069=>"110100110",
  1070=>"011000101",
  1071=>"010100001",
  1072=>"101100010",
  1073=>"001110110",
  1074=>"010001110",
  1075=>"100101111",
  1076=>"111110110",
  1077=>"001111111",
  1078=>"111101110",
  1079=>"011001001",
  1080=>"001000000",
  1081=>"110100001",
  1082=>"000011010",
  1083=>"010100101",
  1084=>"010010000",
  1085=>"100010101",
  1086=>"101001001",
  1087=>"000001000",
  1088=>"100101010",
  1089=>"001010010",
  1090=>"101110001",
  1091=>"101010111",
  1092=>"010100010",
  1093=>"010110100",
  1094=>"000100110",
  1095=>"011101111",
  1096=>"101110001",
  1097=>"001010000",
  1098=>"011111111",
  1099=>"000001110",
  1100=>"111100111",
  1101=>"110010100",
  1102=>"011010100",
  1103=>"110010100",
  1104=>"011001110",
  1105=>"110100100",
  1106=>"000110111",
  1107=>"111001000",
  1108=>"010011110",
  1109=>"000000110",
  1110=>"001011011",
  1111=>"000001000",
  1112=>"000101111",
  1113=>"011101101",
  1114=>"001001001",
  1115=>"011100010",
  1116=>"111101110",
  1117=>"101111100",
  1118=>"001110101",
  1119=>"000101110",
  1120=>"001101000",
  1121=>"010011110",
  1122=>"011110000",
  1123=>"101100110",
  1124=>"011100000",
  1125=>"100111101",
  1126=>"101100100",
  1127=>"100001110",
  1128=>"111011010",
  1129=>"101011010",
  1130=>"000101101",
  1131=>"101001110",
  1132=>"010111001",
  1133=>"000111001",
  1134=>"101100111",
  1135=>"100001101",
  1136=>"000101011",
  1137=>"010011111",
  1138=>"100101111",
  1139=>"000001101",
  1140=>"101111100",
  1141=>"000001111",
  1142=>"100110110",
  1143=>"101101011",
  1144=>"101001000",
  1145=>"111111100",
  1146=>"000010111",
  1147=>"011101110",
  1148=>"101100010",
  1149=>"111011010",
  1150=>"110101110",
  1151=>"001100010",
  1152=>"011110001",
  1153=>"101010000",
  1154=>"010000010",
  1155=>"100110100",
  1156=>"111110111",
  1157=>"000110001",
  1158=>"000101110",
  1159=>"000000100",
  1160=>"110101110",
  1161=>"000111011",
  1162=>"101100111",
  1163=>"101111011",
  1164=>"111111010",
  1165=>"101110111",
  1166=>"100110110",
  1167=>"011101100",
  1168=>"001101111",
  1169=>"101001011",
  1170=>"001111101",
  1171=>"111001001",
  1172=>"011101110",
  1173=>"111000110",
  1174=>"001100001",
  1175=>"001001100",
  1176=>"111101111",
  1177=>"000101011",
  1178=>"101110111",
  1179=>"011000001",
  1180=>"100000110",
  1181=>"101111000",
  1182=>"011100111",
  1183=>"100000000",
  1184=>"110000110",
  1185=>"100000000",
  1186=>"111000010",
  1187=>"101011110",
  1188=>"111111110",
  1189=>"110000011",
  1190=>"101011101",
  1191=>"000100100",
  1192=>"111111110",
  1193=>"101101001",
  1194=>"101010111",
  1195=>"001011010",
  1196=>"110111111",
  1197=>"010111111",
  1198=>"100000010",
  1199=>"011001100",
  1200=>"011101100",
  1201=>"011110101",
  1202=>"010110001",
  1203=>"100010010",
  1204=>"100010101",
  1205=>"100001110",
  1206=>"111111101",
  1207=>"100111010",
  1208=>"011000110",
  1209=>"000110001",
  1210=>"011101001",
  1211=>"101010001",
  1212=>"111101111",
  1213=>"110111110",
  1214=>"010011101",
  1215=>"000010100",
  1216=>"100110110",
  1217=>"111000110",
  1218=>"100111110",
  1219=>"010111110",
  1220=>"110000100",
  1221=>"011010011",
  1222=>"111001111",
  1223=>"110010011",
  1224=>"101011000",
  1225=>"010001011",
  1226=>"111001000",
  1227=>"101110000",
  1228=>"000110001",
  1229=>"000011111",
  1230=>"000001011",
  1231=>"001100001",
  1232=>"101001001",
  1233=>"011101010",
  1234=>"010101000",
  1235=>"100100110",
  1236=>"011011111",
  1237=>"100100101",
  1238=>"000001000",
  1239=>"111001101",
  1240=>"100011110",
  1241=>"100011001",
  1242=>"110101110",
  1243=>"000111111",
  1244=>"000001010",
  1245=>"010111100",
  1246=>"111000111",
  1247=>"001010000",
  1248=>"100010000",
  1249=>"001011111",
  1250=>"101111011",
  1251=>"111101000",
  1252=>"010110010",
  1253=>"011010110",
  1254=>"110111111",
  1255=>"100111001",
  1256=>"111100100",
  1257=>"001111100",
  1258=>"011000100",
  1259=>"000100000",
  1260=>"110100110",
  1261=>"110000110",
  1262=>"001011111",
  1263=>"011111110",
  1264=>"100101000",
  1265=>"010100100",
  1266=>"011111110",
  1267=>"101100111",
  1268=>"101010000",
  1269=>"101101100",
  1270=>"100101111",
  1271=>"010100010",
  1272=>"011010100",
  1273=>"101010110",
  1274=>"000000001",
  1275=>"000110011",
  1276=>"010100100",
  1277=>"000100110",
  1278=>"001101111",
  1279=>"011111010",
  1280=>"110000111",
  1281=>"111111001",
  1282=>"001100110",
  1283=>"011001000",
  1284=>"001101011",
  1285=>"101000101",
  1286=>"000010011",
  1287=>"010011010",
  1288=>"110010010",
  1289=>"111110000",
  1290=>"000101010",
  1291=>"011011010",
  1292=>"001010110",
  1293=>"010011011",
  1294=>"101000001",
  1295=>"010001101",
  1296=>"000101100",
  1297=>"110100011",
  1298=>"110101100",
  1299=>"000111101",
  1300=>"000011100",
  1301=>"100000000",
  1302=>"010010111",
  1303=>"000100001",
  1304=>"110000011",
  1305=>"111011101",
  1306=>"110110110",
  1307=>"100110101",
  1308=>"010111111",
  1309=>"110011111",
  1310=>"101111111",
  1311=>"001010010",
  1312=>"000010011",
  1313=>"100110010",
  1314=>"100111111",
  1315=>"000001100",
  1316=>"010011001",
  1317=>"100011110",
  1318=>"000010011",
  1319=>"010011111",
  1320=>"001000000",
  1321=>"011000100",
  1322=>"011111001",
  1323=>"011101111",
  1324=>"110110100",
  1325=>"001000100",
  1326=>"100010111",
  1327=>"111111101",
  1328=>"000000010",
  1329=>"101101000",
  1330=>"001010101",
  1331=>"010010111",
  1332=>"110011011",
  1333=>"110100100",
  1334=>"000100110",
  1335=>"100110001",
  1336=>"101011010",
  1337=>"101100110",
  1338=>"110110100",
  1339=>"100111010",
  1340=>"101111000",
  1341=>"101101101",
  1342=>"010100001",
  1343=>"111001001",
  1344=>"010001101",
  1345=>"010001010",
  1346=>"100010000",
  1347=>"000101100",
  1348=>"100110100",
  1349=>"010000010",
  1350=>"010011010",
  1351=>"010101111",
  1352=>"100000010",
  1353=>"110100000",
  1354=>"011010101",
  1355=>"100010111",
  1356=>"100010010",
  1357=>"001000000",
  1358=>"101011100",
  1359=>"000110010",
  1360=>"000110000",
  1361=>"011101011",
  1362=>"001000001",
  1363=>"001000001",
  1364=>"100011001",
  1365=>"011111100",
  1366=>"110110101",
  1367=>"011010001",
  1368=>"001001100",
  1369=>"000000111",
  1370=>"000110111",
  1371=>"101001011",
  1372=>"111001010",
  1373=>"101111101",
  1374=>"101011000",
  1375=>"000111111",
  1376=>"111110011",
  1377=>"000111010",
  1378=>"010011110",
  1379=>"000101000",
  1380=>"101010000",
  1381=>"000000110",
  1382=>"101011110",
  1383=>"010111110",
  1384=>"110101000",
  1385=>"000000001",
  1386=>"110010111",
  1387=>"000010100",
  1388=>"101011010",
  1389=>"010010100",
  1390=>"100110000",
  1391=>"010011110",
  1392=>"110100000",
  1393=>"000101010",
  1394=>"110100000",
  1395=>"001101100",
  1396=>"001011000",
  1397=>"001001001",
  1398=>"110110110",
  1399=>"110111101",
  1400=>"001000011",
  1401=>"010111101",
  1402=>"000101111",
  1403=>"001110100",
  1404=>"001000000",
  1405=>"000001110",
  1406=>"110000000",
  1407=>"010101110",
  1408=>"100110001",
  1409=>"010110100",
  1410=>"000010011",
  1411=>"010011110",
  1412=>"011100010",
  1413=>"100100010",
  1414=>"011111010",
  1415=>"101010111",
  1416=>"001010000",
  1417=>"110111000",
  1418=>"000000101",
  1419=>"010000000",
  1420=>"010110001",
  1421=>"000111111",
  1422=>"110100100",
  1423=>"010011110",
  1424=>"011011101",
  1425=>"000100010",
  1426=>"001010101",
  1427=>"100000101",
  1428=>"010110010",
  1429=>"111101000",
  1430=>"100100000",
  1431=>"001001110",
  1432=>"111001001",
  1433=>"100001010",
  1434=>"001001110",
  1435=>"001011010",
  1436=>"000101001",
  1437=>"101010101",
  1438=>"111010101",
  1439=>"111111101",
  1440=>"110000010",
  1441=>"111100100",
  1442=>"110000101",
  1443=>"110101110",
  1444=>"011000010",
  1445=>"000010101",
  1446=>"101011110",
  1447=>"001000011",
  1448=>"010001001",
  1449=>"100000010",
  1450=>"100100100",
  1451=>"001101111",
  1452=>"010010010",
  1453=>"010100000",
  1454=>"000000000",
  1455=>"101011100",
  1456=>"000100010",
  1457=>"100100110",
  1458=>"111101111",
  1459=>"011110000",
  1460=>"010100111",
  1461=>"100001111",
  1462=>"100010111",
  1463=>"110100010",
  1464=>"110011010",
  1465=>"110000010",
  1466=>"000011110",
  1467=>"111001000",
  1468=>"110101110",
  1469=>"011000001",
  1470=>"111110111",
  1471=>"010010000",
  1472=>"010001010",
  1473=>"000110001",
  1474=>"010110001",
  1475=>"001111110",
  1476=>"101101100",
  1477=>"110110011",
  1478=>"011000010",
  1479=>"110000100",
  1480=>"001010100",
  1481=>"101111110",
  1482=>"111011010",
  1483=>"010110000",
  1484=>"101100111",
  1485=>"001001001",
  1486=>"011000011",
  1487=>"000111011",
  1488=>"000011001",
  1489=>"110110110",
  1490=>"001111001",
  1491=>"100010111",
  1492=>"001011100",
  1493=>"100101100",
  1494=>"101001100",
  1495=>"110100110",
  1496=>"101011011",
  1497=>"110000110",
  1498=>"000000111",
  1499=>"001111001",
  1500=>"111100110",
  1501=>"000010010",
  1502=>"111110000",
  1503=>"100001100",
  1504=>"111001011",
  1505=>"111101100",
  1506=>"100111010",
  1507=>"100000100",
  1508=>"111101100",
  1509=>"100111110",
  1510=>"011010010",
  1511=>"110101110",
  1512=>"010001101",
  1513=>"000010001",
  1514=>"101010011",
  1515=>"000001111",
  1516=>"001100000",
  1517=>"010001101",
  1518=>"110110111",
  1519=>"110101010",
  1520=>"110101001",
  1521=>"110011000",
  1522=>"100010010",
  1523=>"001011011",
  1524=>"011111001",
  1525=>"110010111",
  1526=>"101111111",
  1527=>"000000001",
  1528=>"100110101",
  1529=>"011000101",
  1530=>"110000001",
  1531=>"001001011",
  1532=>"111111001",
  1533=>"011010110",
  1534=>"001100010",
  1535=>"011110100",
  1536=>"000000111",
  1537=>"010011101",
  1538=>"111010100",
  1539=>"100100101",
  1540=>"000110010",
  1541=>"010010111",
  1542=>"010000001",
  1543=>"111000101",
  1544=>"110111100",
  1545=>"110011100",
  1546=>"110100000",
  1547=>"000011111",
  1548=>"001111011",
  1549=>"011000110",
  1550=>"100100010",
  1551=>"010101110",
  1552=>"000101010",
  1553=>"101110001",
  1554=>"111010110",
  1555=>"000000111",
  1556=>"000010001",
  1557=>"011100111",
  1558=>"110110111",
  1559=>"101101110",
  1560=>"010010111",
  1561=>"100111000",
  1562=>"001000110",
  1563=>"010100001",
  1564=>"100001111",
  1565=>"110000010",
  1566=>"000011001",
  1567=>"110011010",
  1568=>"110100100",
  1569=>"111011011",
  1570=>"101111100",
  1571=>"000101111",
  1572=>"010010011",
  1573=>"001011011",
  1574=>"011110110",
  1575=>"100101110",
  1576=>"100000100",
  1577=>"111100010",
  1578=>"111111011",
  1579=>"100010110",
  1580=>"111001110",
  1581=>"001010111",
  1582=>"110010000",
  1583=>"111010011",
  1584=>"011010101",
  1585=>"011110010",
  1586=>"100100001",
  1587=>"110111101",
  1588=>"100000101",
  1589=>"001000110",
  1590=>"101100000",
  1591=>"110111011",
  1592=>"111100010",
  1593=>"000110111",
  1594=>"110001100",
  1595=>"010000100",
  1596=>"001010011",
  1597=>"100100100",
  1598=>"101000001",
  1599=>"001100110",
  1600=>"001010100",
  1601=>"101011000",
  1602=>"101010001",
  1603=>"010000110",
  1604=>"111010101",
  1605=>"100110100",
  1606=>"100010001",
  1607=>"101011110",
  1608=>"110100100",
  1609=>"010001001",
  1610=>"010110110",
  1611=>"000101100",
  1612=>"010010101",
  1613=>"110111011",
  1614=>"110111011",
  1615=>"111001111",
  1616=>"111001000",
  1617=>"010101100",
  1618=>"000000000",
  1619=>"100011010",
  1620=>"100011001",
  1621=>"001010000",
  1622=>"101011101",
  1623=>"010010111",
  1624=>"001000111",
  1625=>"101111001",
  1626=>"110011000",
  1627=>"110000111",
  1628=>"100111110",
  1629=>"111010100",
  1630=>"111101101",
  1631=>"000101010",
  1632=>"101011111",
  1633=>"001000001",
  1634=>"100000101",
  1635=>"000101100",
  1636=>"100001001",
  1637=>"101111100",
  1638=>"010100100",
  1639=>"011001010",
  1640=>"010011101",
  1641=>"110000010",
  1642=>"111001011",
  1643=>"000010110",
  1644=>"110110110",
  1645=>"001001001",
  1646=>"110001110",
  1647=>"010010111",
  1648=>"111011101",
  1649=>"000101010",
  1650=>"110000001",
  1651=>"101000001",
  1652=>"000110001",
  1653=>"111110011",
  1654=>"010001111",
  1655=>"110110111",
  1656=>"110101000",
  1657=>"000111101",
  1658=>"111111110",
  1659=>"001001010",
  1660=>"001100000",
  1661=>"000010101",
  1662=>"100000100",
  1663=>"110101000",
  1664=>"100000110",
  1665=>"000000000",
  1666=>"101011011",
  1667=>"000001001",
  1668=>"100100000",
  1669=>"011110111",
  1670=>"101001101",
  1671=>"011110001",
  1672=>"101011010",
  1673=>"001001110",
  1674=>"101000001",
  1675=>"101000001",
  1676=>"111010000",
  1677=>"001011100",
  1678=>"100010001",
  1679=>"101100110",
  1680=>"110011010",
  1681=>"000000000",
  1682=>"010001011",
  1683=>"100111011",
  1684=>"101010000",
  1685=>"110111000",
  1686=>"101100001",
  1687=>"000101000",
  1688=>"110001001",
  1689=>"001000100",
  1690=>"000001101",
  1691=>"000001100",
  1692=>"100010011",
  1693=>"011100100",
  1694=>"111000111",
  1695=>"111100111",
  1696=>"111111001",
  1697=>"100110110",
  1698=>"100000101",
  1699=>"001000011",
  1700=>"100100100",
  1701=>"100001000",
  1702=>"101101010",
  1703=>"011010001",
  1704=>"100001101",
  1705=>"110110111",
  1706=>"011000000",
  1707=>"010100010",
  1708=>"000101111",
  1709=>"000000110",
  1710=>"010011110",
  1711=>"001001001",
  1712=>"001111010",
  1713=>"010001111",
  1714=>"111101001",
  1715=>"011011000",
  1716=>"111011101",
  1717=>"000111010",
  1718=>"100101011",
  1719=>"111010100",
  1720=>"000110000",
  1721=>"011011100",
  1722=>"101001000",
  1723=>"000101100",
  1724=>"011101110",
  1725=>"000000001",
  1726=>"100110001",
  1727=>"011110010",
  1728=>"101000000",
  1729=>"001110011",
  1730=>"100001100",
  1731=>"010011010",
  1732=>"000001001",
  1733=>"001011100",
  1734=>"001000010",
  1735=>"011001111",
  1736=>"111000101",
  1737=>"110100000",
  1738=>"111111000",
  1739=>"010001111",
  1740=>"001110000",
  1741=>"001010011",
  1742=>"110010011",
  1743=>"010110110",
  1744=>"011110001",
  1745=>"001000011",
  1746=>"101000001",
  1747=>"000000011",
  1748=>"000110101",
  1749=>"010001101",
  1750=>"110100001",
  1751=>"000010111",
  1752=>"111110111",
  1753=>"000001110",
  1754=>"101110011",
  1755=>"000001010",
  1756=>"011101100",
  1757=>"111110101",
  1758=>"011101010",
  1759=>"110011111",
  1760=>"110111101",
  1761=>"100100010",
  1762=>"011011011",
  1763=>"100100000",
  1764=>"011110111",
  1765=>"110011010",
  1766=>"111010011",
  1767=>"101101111",
  1768=>"110111101",
  1769=>"000000010",
  1770=>"010000000",
  1771=>"110110101",
  1772=>"011010001",
  1773=>"100110110",
  1774=>"110010000",
  1775=>"000010010",
  1776=>"000010010",
  1777=>"110110011",
  1778=>"100010110",
  1779=>"010000100",
  1780=>"110101011",
  1781=>"011001100",
  1782=>"001011000",
  1783=>"110010001",
  1784=>"010110001",
  1785=>"010110101",
  1786=>"001001101",
  1787=>"011000100",
  1788=>"110000001",
  1789=>"110100011",
  1790=>"001110101",
  1791=>"110101011",
  1792=>"000011001",
  1793=>"010000000",
  1794=>"110111110",
  1795=>"110100100",
  1796=>"000000011",
  1797=>"000010011",
  1798=>"001101111",
  1799=>"101111001",
  1800=>"101110001",
  1801=>"001011101",
  1802=>"011111111",
  1803=>"010011111",
  1804=>"000011111",
  1805=>"001001100",
  1806=>"110111001",
  1807=>"100000100",
  1808=>"111101110",
  1809=>"110010010",
  1810=>"010100111",
  1811=>"011011100",
  1812=>"101010110",
  1813=>"011110011",
  1814=>"101011111",
  1815=>"111100001",
  1816=>"000000000",
  1817=>"000010001",
  1818=>"111111000",
  1819=>"001001010",
  1820=>"111000010",
  1821=>"110100011",
  1822=>"110001111",
  1823=>"111110001",
  1824=>"010001110",
  1825=>"101111010",
  1826=>"111101000",
  1827=>"110101101",
  1828=>"101111111",
  1829=>"000010111",
  1830=>"000011001",
  1831=>"010001110",
  1832=>"110010000",
  1833=>"101001001",
  1834=>"001000001",
  1835=>"101000110",
  1836=>"110100110",
  1837=>"101110100",
  1838=>"000000110",
  1839=>"000001101",
  1840=>"111000000",
  1841=>"000111010",
  1842=>"110011101",
  1843=>"001001101",
  1844=>"010010110",
  1845=>"001111111",
  1846=>"110110100",
  1847=>"011000101",
  1848=>"110101110",
  1849=>"110010100",
  1850=>"010000110",
  1851=>"100100010",
  1852=>"101101000",
  1853=>"000000001",
  1854=>"100101101",
  1855=>"100001010",
  1856=>"100101111",
  1857=>"000101011",
  1858=>"110010011",
  1859=>"010001100",
  1860=>"001001000",
  1861=>"100111111",
  1862=>"000101010",
  1863=>"110110100",
  1864=>"001101110",
  1865=>"110000011",
  1866=>"001010110",
  1867=>"000111011",
  1868=>"101001001",
  1869=>"100100010",
  1870=>"110111001",
  1871=>"100001011",
  1872=>"101100111",
  1873=>"110011110",
  1874=>"110111110",
  1875=>"100100010",
  1876=>"001110011",
  1877=>"100101010",
  1878=>"110101010",
  1879=>"001000011",
  1880=>"111001001",
  1881=>"001100111",
  1882=>"100100101",
  1883=>"100110001",
  1884=>"111101001",
  1885=>"101001010",
  1886=>"100110101",
  1887=>"001101001",
  1888=>"110101101",
  1889=>"111101010",
  1890=>"010010001",
  1891=>"101000100",
  1892=>"101110011",
  1893=>"100010010",
  1894=>"100001110",
  1895=>"011011010",
  1896=>"111011110",
  1897=>"100111011",
  1898=>"000011111",
  1899=>"110011110",
  1900=>"101110011",
  1901=>"000001010",
  1902=>"100000001",
  1903=>"110110101",
  1904=>"101011110",
  1905=>"101011011",
  1906=>"001101110",
  1907=>"110111101",
  1908=>"100110100",
  1909=>"000010011",
  1910=>"110000101",
  1911=>"110000100",
  1912=>"010101100",
  1913=>"001100101",
  1914=>"110100111",
  1915=>"010011001",
  1916=>"101010100",
  1917=>"010000001",
  1918=>"110111101",
  1919=>"011110111",
  1920=>"110111000",
  1921=>"000100000",
  1922=>"111110111",
  1923=>"111010010",
  1924=>"010001001",
  1925=>"000101011",
  1926=>"001000100",
  1927=>"110000111",
  1928=>"111100111",
  1929=>"111011000",
  1930=>"000000010",
  1931=>"010001011",
  1932=>"010000010",
  1933=>"010001000",
  1934=>"000000011",
  1935=>"010100000",
  1936=>"110101110",
  1937=>"110000110",
  1938=>"111111111",
  1939=>"001101111",
  1940=>"111110011",
  1941=>"111100110",
  1942=>"010111101",
  1943=>"011000110",
  1944=>"001010101",
  1945=>"001001101",
  1946=>"001000111",
  1947=>"001111011",
  1948=>"101111000",
  1949=>"011101010",
  1950=>"101010000",
  1951=>"000101110",
  1952=>"100000110",
  1953=>"001010010",
  1954=>"000111010",
  1955=>"111001000",
  1956=>"101101111",
  1957=>"000111011",
  1958=>"010011011",
  1959=>"000010011",
  1960=>"100110001",
  1961=>"100001010",
  1962=>"111110111",
  1963=>"011110011",
  1964=>"110001110",
  1965=>"011111100",
  1966=>"110100011",
  1967=>"010000011",
  1968=>"001011010",
  1969=>"101001011",
  1970=>"010010000",
  1971=>"110111001",
  1972=>"011011111",
  1973=>"010100000",
  1974=>"010111101",
  1975=>"110011100",
  1976=>"100111001",
  1977=>"010111100",
  1978=>"100010000",
  1979=>"101111000",
  1980=>"011010010",
  1981=>"100110000",
  1982=>"100110110",
  1983=>"110111100",
  1984=>"001111111",
  1985=>"000000001",
  1986=>"010100010",
  1987=>"010110000",
  1988=>"000111100",
  1989=>"000111000",
  1990=>"011111110",
  1991=>"011001110",
  1992=>"111111111",
  1993=>"100111101",
  1994=>"000010111",
  1995=>"100010101",
  1996=>"110111110",
  1997=>"100000111",
  1998=>"010101110",
  1999=>"100100100",
  2000=>"111101011",
  2001=>"010011110",
  2002=>"011110000",
  2003=>"111100111",
  2004=>"001010011",
  2005=>"000000100",
  2006=>"100000001",
  2007=>"110101001",
  2008=>"110111000",
  2009=>"000011111",
  2010=>"111101000",
  2011=>"111000100",
  2012=>"000001111",
  2013=>"000101101",
  2014=>"000101000",
  2015=>"100001110",
  2016=>"001110110",
  2017=>"000001011",
  2018=>"000010001",
  2019=>"110001000",
  2020=>"000110010",
  2021=>"110001011",
  2022=>"100000011",
  2023=>"111001111",
  2024=>"110000110",
  2025=>"001101010",
  2026=>"111001011",
  2027=>"100010011",
  2028=>"011101011",
  2029=>"110110111",
  2030=>"101001101",
  2031=>"010110010",
  2032=>"110101000",
  2033=>"000010100",
  2034=>"011110010",
  2035=>"111110101",
  2036=>"110101100",
  2037=>"000000000",
  2038=>"111100101",
  2039=>"110101001",
  2040=>"110010000",
  2041=>"101111010",
  2042=>"100000101",
  2043=>"000000000",
  2044=>"000100110",
  2045=>"000010001",
  2046=>"011000100",
  2047=>"110011000",
  2048=>"000110011",
  2049=>"000111101",
  2050=>"100001110",
  2051=>"011001010",
  2052=>"101100100",
  2053=>"110111110",
  2054=>"000111100",
  2055=>"011010000",
  2056=>"100010110",
  2057=>"010101100",
  2058=>"110010111",
  2059=>"110010110",
  2060=>"001011111",
  2061=>"001000010",
  2062=>"001000000",
  2063=>"101100111",
  2064=>"000111010",
  2065=>"010101001",
  2066=>"100100111",
  2067=>"101110001",
  2068=>"111001101",
  2069=>"010011010",
  2070=>"101001101",
  2071=>"001101000",
  2072=>"010001000",
  2073=>"011010010",
  2074=>"110011011",
  2075=>"101101101",
  2076=>"110111110",
  2077=>"100010100",
  2078=>"001011110",
  2079=>"010010001",
  2080=>"001111100",
  2081=>"010000100",
  2082=>"101010111",
  2083=>"110110110",
  2084=>"010100001",
  2085=>"001101000",
  2086=>"100000010",
  2087=>"100110000",
  2088=>"011101010",
  2089=>"001111001",
  2090=>"000111100",
  2091=>"000010010",
  2092=>"100110010",
  2093=>"000101010",
  2094=>"011100100",
  2095=>"010000000",
  2096=>"010110100",
  2097=>"110000010",
  2098=>"011010111",
  2099=>"000001111",
  2100=>"110000110",
  2101=>"011001010",
  2102=>"111011110",
  2103=>"000000011",
  2104=>"111100110",
  2105=>"011100001",
  2106=>"010001000",
  2107=>"101011110",
  2108=>"011000101",
  2109=>"010111001",
  2110=>"011000111",
  2111=>"011010001",
  2112=>"111001010",
  2113=>"000100110",
  2114=>"110111011",
  2115=>"001111101",
  2116=>"101001100",
  2117=>"000110001",
  2118=>"011110111",
  2119=>"101110101",
  2120=>"111100101",
  2121=>"000000000",
  2122=>"011001011",
  2123=>"001111001",
  2124=>"000001010",
  2125=>"010110000",
  2126=>"000101100",
  2127=>"000010101",
  2128=>"000000010",
  2129=>"110001001",
  2130=>"011000011",
  2131=>"100100010",
  2132=>"000110010",
  2133=>"000001111",
  2134=>"111111010",
  2135=>"111001111",
  2136=>"010100111",
  2137=>"001101111",
  2138=>"000110000",
  2139=>"100000000",
  2140=>"100010010",
  2141=>"110010110",
  2142=>"000101110",
  2143=>"110010001",
  2144=>"011110110",
  2145=>"100011111",
  2146=>"000000001",
  2147=>"101110000",
  2148=>"110010010",
  2149=>"000101001",
  2150=>"000111100",
  2151=>"111100111",
  2152=>"011011110",
  2153=>"011011011",
  2154=>"011000111",
  2155=>"101101000",
  2156=>"000101100",
  2157=>"000011100",
  2158=>"111010011",
  2159=>"100010000",
  2160=>"111000000",
  2161=>"100110100",
  2162=>"111001100",
  2163=>"100000110",
  2164=>"001001111",
  2165=>"100101001",
  2166=>"101010111",
  2167=>"011101011",
  2168=>"001001001",
  2169=>"110010010",
  2170=>"000011111",
  2171=>"101001001",
  2172=>"111100011",
  2173=>"110000011",
  2174=>"001011000",
  2175=>"001001000",
  2176=>"111000011",
  2177=>"110000001",
  2178=>"011111100",
  2179=>"000000000",
  2180=>"110000010",
  2181=>"101000110",
  2182=>"111101011",
  2183=>"111100001",
  2184=>"111000101",
  2185=>"101111011",
  2186=>"110101101",
  2187=>"000110010",
  2188=>"010000100",
  2189=>"011111000",
  2190=>"110000100",
  2191=>"110111011",
  2192=>"010001000",
  2193=>"100110000",
  2194=>"100111010",
  2195=>"010101011",
  2196=>"001101011",
  2197=>"001001111",
  2198=>"111111111",
  2199=>"111011011",
  2200=>"011111101",
  2201=>"100000101",
  2202=>"101111001",
  2203=>"001001011",
  2204=>"100011101",
  2205=>"101110101",
  2206=>"011101100",
  2207=>"000100010",
  2208=>"011011100",
  2209=>"011101111",
  2210=>"000010111",
  2211=>"010000001",
  2212=>"100101100",
  2213=>"001100110",
  2214=>"011001111",
  2215=>"110100101",
  2216=>"101100101",
  2217=>"000010010",
  2218=>"111101011",
  2219=>"110010100",
  2220=>"011100001",
  2221=>"001111000",
  2222=>"001110011",
  2223=>"010110100",
  2224=>"110111100",
  2225=>"001000001",
  2226=>"101110101",
  2227=>"100101011",
  2228=>"000110100",
  2229=>"100101010",
  2230=>"011111011",
  2231=>"111010001",
  2232=>"110111011",
  2233=>"111010111",
  2234=>"010000001",
  2235=>"011001001",
  2236=>"100101000",
  2237=>"111100001",
  2238=>"001011111",
  2239=>"100000111",
  2240=>"101001011",
  2241=>"100011011",
  2242=>"100001011",
  2243=>"001001110",
  2244=>"101111010",
  2245=>"100001100",
  2246=>"101111010",
  2247=>"011001010",
  2248=>"110010000",
  2249=>"101011100",
  2250=>"001110011",
  2251=>"011010110",
  2252=>"000101001",
  2253=>"001010001",
  2254=>"101011000",
  2255=>"010100101",
  2256=>"001010001",
  2257=>"110111100",
  2258=>"000010110",
  2259=>"001100110",
  2260=>"111001000",
  2261=>"110010000",
  2262=>"100000100",
  2263=>"010100110",
  2264=>"000000000",
  2265=>"101101000",
  2266=>"000110010",
  2267=>"000110010",
  2268=>"000110010",
  2269=>"011000111",
  2270=>"100010000",
  2271=>"110100100",
  2272=>"101011111",
  2273=>"111110111",
  2274=>"000011010",
  2275=>"110001001",
  2276=>"010010101",
  2277=>"101110110",
  2278=>"111101011",
  2279=>"011110100",
  2280=>"111010111",
  2281=>"100111111",
  2282=>"001100110",
  2283=>"000110101",
  2284=>"100101001",
  2285=>"101111100",
  2286=>"000011111",
  2287=>"101101010",
  2288=>"000100001",
  2289=>"100000101",
  2290=>"010010010",
  2291=>"000000001",
  2292=>"110000011",
  2293=>"001001000",
  2294=>"010110000",
  2295=>"101111110",
  2296=>"011000000",
  2297=>"111011000",
  2298=>"110111011",
  2299=>"101000101",
  2300=>"101001110",
  2301=>"001000010",
  2302=>"011010110",
  2303=>"110111110",
  2304=>"011000001",
  2305=>"101111111",
  2306=>"110000001",
  2307=>"001001011",
  2308=>"010010001",
  2309=>"101001111",
  2310=>"110100101",
  2311=>"100000100",
  2312=>"000111101",
  2313=>"110010110",
  2314=>"000101010",
  2315=>"110111010",
  2316=>"010101111",
  2317=>"100000000",
  2318=>"100001111",
  2319=>"111110010",
  2320=>"001100000",
  2321=>"100101001",
  2322=>"011110110",
  2323=>"001010010",
  2324=>"010101101",
  2325=>"100000101",
  2326=>"101111100",
  2327=>"101011000",
  2328=>"111111010",
  2329=>"111001011",
  2330=>"011110011",
  2331=>"110010010",
  2332=>"101001011",
  2333=>"011000010",
  2334=>"001101000",
  2335=>"100100001",
  2336=>"000000011",
  2337=>"101001101",
  2338=>"111101010",
  2339=>"011100011",
  2340=>"111111000",
  2341=>"010000000",
  2342=>"001000100",
  2343=>"010110100",
  2344=>"000011000",
  2345=>"100010111",
  2346=>"111010011",
  2347=>"101111110",
  2348=>"000001100",
  2349=>"001110000",
  2350=>"110000010",
  2351=>"101010000",
  2352=>"010110000",
  2353=>"111100001",
  2354=>"110111010",
  2355=>"010000000",
  2356=>"111001100",
  2357=>"001110000",
  2358=>"111001111",
  2359=>"010011001",
  2360=>"111111111",
  2361=>"011010101",
  2362=>"011010000",
  2363=>"101101001",
  2364=>"110011101",
  2365=>"011100010",
  2366=>"110111011",
  2367=>"111000000",
  2368=>"100000000",
  2369=>"111101001",
  2370=>"110110011",
  2371=>"111010100",
  2372=>"010101100",
  2373=>"111011110",
  2374=>"111111100",
  2375=>"000110110",
  2376=>"111101011",
  2377=>"101111101",
  2378=>"011000000",
  2379=>"111010011",
  2380=>"110001100",
  2381=>"101000011",
  2382=>"101111111",
  2383=>"111111110",
  2384=>"111000011",
  2385=>"000110110",
  2386=>"110011001",
  2387=>"100000110",
  2388=>"000010000",
  2389=>"100100111",
  2390=>"110111111",
  2391=>"000010101",
  2392=>"110011011",
  2393=>"010010001",
  2394=>"100101111",
  2395=>"111101111",
  2396=>"000010110",
  2397=>"100011100",
  2398=>"101101100",
  2399=>"011011100",
  2400=>"110110001",
  2401=>"010011000",
  2402=>"111100100",
  2403=>"110011010",
  2404=>"001000000",
  2405=>"010010111",
  2406=>"001001011",
  2407=>"011111000",
  2408=>"110101111",
  2409=>"100001010",
  2410=>"011100010",
  2411=>"010101011",
  2412=>"100001110",
  2413=>"010001001",
  2414=>"010110100",
  2415=>"101101011",
  2416=>"000110110",
  2417=>"111110001",
  2418=>"101110000",
  2419=>"011010110",
  2420=>"001101011",
  2421=>"010000101",
  2422=>"110010100",
  2423=>"010010100",
  2424=>"100011010",
  2425=>"010111011",
  2426=>"111111111",
  2427=>"001110100",
  2428=>"010100111",
  2429=>"111101110",
  2430=>"110011100",
  2431=>"001000101",
  2432=>"111011011",
  2433=>"110000100",
  2434=>"000100111",
  2435=>"011001011",
  2436=>"011110110",
  2437=>"101111010",
  2438=>"111111001",
  2439=>"111011110",
  2440=>"101010111",
  2441=>"101110001",
  2442=>"111111100",
  2443=>"111011111",
  2444=>"010001000",
  2445=>"110010000",
  2446=>"000000001",
  2447=>"000000100",
  2448=>"010110011",
  2449=>"010100001",
  2450=>"111011100",
  2451=>"011000101",
  2452=>"101111010",
  2453=>"110001001",
  2454=>"011001100",
  2455=>"010100000",
  2456=>"000111101",
  2457=>"000010000",
  2458=>"011110111",
  2459=>"001110010",
  2460=>"001110100",
  2461=>"010110000",
  2462=>"010010101",
  2463=>"000011110",
  2464=>"101100100",
  2465=>"010010010",
  2466=>"111011010",
  2467=>"011100001",
  2468=>"110100101",
  2469=>"001001001",
  2470=>"110111100",
  2471=>"110101011",
  2472=>"011110100",
  2473=>"101000010",
  2474=>"111111101",
  2475=>"001000100",
  2476=>"001001011",
  2477=>"001100111",
  2478=>"010001100",
  2479=>"000100011",
  2480=>"010100101",
  2481=>"011100010",
  2482=>"011001111",
  2483=>"101000101",
  2484=>"110110001",
  2485=>"111010100",
  2486=>"101100010",
  2487=>"100001111",
  2488=>"001011101",
  2489=>"101110110",
  2490=>"101111010",
  2491=>"111010011",
  2492=>"000100011",
  2493=>"010110011",
  2494=>"011011000",
  2495=>"011011101",
  2496=>"111011010",
  2497=>"110101000",
  2498=>"011110001",
  2499=>"010011111",
  2500=>"000100110",
  2501=>"110011101",
  2502=>"010110010",
  2503=>"110101101",
  2504=>"000101100",
  2505=>"000001001",
  2506=>"001010001",
  2507=>"100101001",
  2508=>"011100010",
  2509=>"100100000",
  2510=>"111110011",
  2511=>"110010011",
  2512=>"010111111",
  2513=>"111110110",
  2514=>"111011111",
  2515=>"000100000",
  2516=>"001001101",
  2517=>"110001100",
  2518=>"011100010",
  2519=>"001110111",
  2520=>"001001001",
  2521=>"010000010",
  2522=>"011100111",
  2523=>"111111011",
  2524=>"101101101",
  2525=>"111010011",
  2526=>"001100011",
  2527=>"111111010",
  2528=>"111000100",
  2529=>"001110010",
  2530=>"101111000",
  2531=>"010101001",
  2532=>"100101100",
  2533=>"010000010",
  2534=>"000111000",
  2535=>"101101011",
  2536=>"110010101",
  2537=>"000011111",
  2538=>"111100010",
  2539=>"010011000",
  2540=>"101100110",
  2541=>"000100101",
  2542=>"110110010",
  2543=>"001101010",
  2544=>"101110111",
  2545=>"110001101",
  2546=>"001001100",
  2547=>"101100100",
  2548=>"110111101",
  2549=>"110100001",
  2550=>"001010011",
  2551=>"001101110",
  2552=>"011011001",
  2553=>"100010010",
  2554=>"010000001",
  2555=>"011111011",
  2556=>"110011111",
  2557=>"001111010",
  2558=>"000000111",
  2559=>"000001011",
  2560=>"110110001",
  2561=>"101011010",
  2562=>"111011111",
  2563=>"000111100",
  2564=>"011100100",
  2565=>"001001100",
  2566=>"110110001",
  2567=>"001100000",
  2568=>"101110110",
  2569=>"100001011",
  2570=>"001010101",
  2571=>"110000001",
  2572=>"011001111",
  2573=>"010001000",
  2574=>"011011001",
  2575=>"101000011",
  2576=>"111000100",
  2577=>"101011110",
  2578=>"000011000",
  2579=>"110100110",
  2580=>"110011110",
  2581=>"000110100",
  2582=>"001100001",
  2583=>"011100010",
  2584=>"111000110",
  2585=>"000111110",
  2586=>"000101010",
  2587=>"100111101",
  2588=>"110111011",
  2589=>"100000111",
  2590=>"101101111",
  2591=>"111001101",
  2592=>"100000110",
  2593=>"001011111",
  2594=>"101011001",
  2595=>"010011110",
  2596=>"011110011",
  2597=>"010111101",
  2598=>"011011100",
  2599=>"011000000",
  2600=>"010011010",
  2601=>"010111101",
  2602=>"011000010",
  2603=>"001110110",
  2604=>"101100000",
  2605=>"011111000",
  2606=>"001110111",
  2607=>"000011111",
  2608=>"000111101",
  2609=>"010001001",
  2610=>"000100100",
  2611=>"000010001",
  2612=>"001110111",
  2613=>"010000110",
  2614=>"001001100",
  2615=>"100000001",
  2616=>"001001001",
  2617=>"111011100",
  2618=>"111110001",
  2619=>"000110111",
  2620=>"001100000",
  2621=>"100111100",
  2622=>"110011010",
  2623=>"100011111",
  2624=>"000010010",
  2625=>"001100000",
  2626=>"110001010",
  2627=>"110111000",
  2628=>"100110101",
  2629=>"000000111",
  2630=>"010111111",
  2631=>"110100001",
  2632=>"110011000",
  2633=>"011101010",
  2634=>"110111000",
  2635=>"101010110",
  2636=>"001101101",
  2637=>"101001110",
  2638=>"001111001",
  2639=>"111011110",
  2640=>"110001011",
  2641=>"111001111",
  2642=>"110000000",
  2643=>"000111000",
  2644=>"100100011",
  2645=>"001101010",
  2646=>"001100111",
  2647=>"000011011",
  2648=>"100010011",
  2649=>"101111001",
  2650=>"111100101",
  2651=>"100101011",
  2652=>"111111010",
  2653=>"100000101",
  2654=>"011010000",
  2655=>"001001011",
  2656=>"010000111",
  2657=>"001010111",
  2658=>"110001101",
  2659=>"110111000",
  2660=>"001010101",
  2661=>"001001111",
  2662=>"001111010",
  2663=>"111001011",
  2664=>"000000111",
  2665=>"000101001",
  2666=>"101000000",
  2667=>"000000110",
  2668=>"011100010",
  2669=>"001101111",
  2670=>"111011101",
  2671=>"010111111",
  2672=>"011111010",
  2673=>"001100111",
  2674=>"000111000",
  2675=>"110100110",
  2676=>"101110010",
  2677=>"100000100",
  2678=>"101101000",
  2679=>"011010100",
  2680=>"110000011",
  2681=>"100100001",
  2682=>"001001010",
  2683=>"000110010",
  2684=>"101011010",
  2685=>"111010001",
  2686=>"100011110",
  2687=>"110100000",
  2688=>"011100110",
  2689=>"111111111",
  2690=>"110001001",
  2691=>"110010011",
  2692=>"100010101",
  2693=>"101011001",
  2694=>"011110010",
  2695=>"011101001",
  2696=>"000010000",
  2697=>"111110101",
  2698=>"111001110",
  2699=>"111100100",
  2700=>"010101000",
  2701=>"011001001",
  2702=>"001001011",
  2703=>"010001110",
  2704=>"010001010",
  2705=>"111110000",
  2706=>"001101011",
  2707=>"000000110",
  2708=>"100110000",
  2709=>"110110111",
  2710=>"001101010",
  2711=>"000010110",
  2712=>"011111111",
  2713=>"100010001",
  2714=>"111011001",
  2715=>"000110001",
  2716=>"111000101",
  2717=>"000000000",
  2718=>"000011100",
  2719=>"000101000",
  2720=>"110011111",
  2721=>"011000110",
  2722=>"110111010",
  2723=>"000110101",
  2724=>"101001011",
  2725=>"100100001",
  2726=>"000000110",
  2727=>"110101110",
  2728=>"000011110",
  2729=>"000010001",
  2730=>"101001100",
  2731=>"111101001",
  2732=>"010011110",
  2733=>"010010111",
  2734=>"101100101",
  2735=>"011001111",
  2736=>"000001010",
  2737=>"010100011",
  2738=>"010111110",
  2739=>"001101000",
  2740=>"001010000",
  2741=>"010111010",
  2742=>"001011110",
  2743=>"111111100",
  2744=>"111000110",
  2745=>"000000000",
  2746=>"010111101",
  2747=>"100000110",
  2748=>"000100010",
  2749=>"110110101",
  2750=>"110101001",
  2751=>"001111100",
  2752=>"101011111",
  2753=>"011100000",
  2754=>"010010101",
  2755=>"010110100",
  2756=>"011110111",
  2757=>"100011010",
  2758=>"101111100",
  2759=>"111010100",
  2760=>"000001000",
  2761=>"011011000",
  2762=>"111111010",
  2763=>"010011101",
  2764=>"001011100",
  2765=>"100010010",
  2766=>"101101010",
  2767=>"101110111",
  2768=>"011111111",
  2769=>"010011001",
  2770=>"111010101",
  2771=>"110110001",
  2772=>"011101010",
  2773=>"111111100",
  2774=>"111110001",
  2775=>"111111110",
  2776=>"011111101",
  2777=>"011011110",
  2778=>"100100110",
  2779=>"001011100",
  2780=>"010100010",
  2781=>"101000001",
  2782=>"010111101",
  2783=>"011101101",
  2784=>"100001010",
  2785=>"000101100",
  2786=>"110000001",
  2787=>"110101011",
  2788=>"111011010",
  2789=>"010100011",
  2790=>"111100100",
  2791=>"101000100",
  2792=>"111110001",
  2793=>"000101110",
  2794=>"010011101",
  2795=>"001010000",
  2796=>"110111111",
  2797=>"111101101",
  2798=>"100100011",
  2799=>"000011011",
  2800=>"100100011",
  2801=>"011001000",
  2802=>"111111111",
  2803=>"111010011",
  2804=>"000010101",
  2805=>"011100011",
  2806=>"100000000",
  2807=>"011100110",
  2808=>"000110000",
  2809=>"100101011",
  2810=>"110111010",
  2811=>"010111110",
  2812=>"000111110",
  2813=>"011101110",
  2814=>"111010110",
  2815=>"000100001",
  2816=>"110000110",
  2817=>"111011111",
  2818=>"001110111",
  2819=>"011011110",
  2820=>"100001000",
  2821=>"100011001",
  2822=>"100001000",
  2823=>"010001010",
  2824=>"011100111",
  2825=>"011001010",
  2826=>"000101100",
  2827=>"111010001",
  2828=>"000100100",
  2829=>"110101111",
  2830=>"100011011",
  2831=>"110100101",
  2832=>"111011101",
  2833=>"100000010",
  2834=>"001111011",
  2835=>"001001110",
  2836=>"001110101",
  2837=>"010010010",
  2838=>"111100110",
  2839=>"000000101",
  2840=>"110001111",
  2841=>"010010001",
  2842=>"000000001",
  2843=>"011011001",
  2844=>"010101011",
  2845=>"101010001",
  2846=>"110000011",
  2847=>"101011101",
  2848=>"100001100",
  2849=>"100111100",
  2850=>"100111111",
  2851=>"011100100",
  2852=>"101111111",
  2853=>"111101101",
  2854=>"000100101",
  2855=>"111000000",
  2856=>"011100110",
  2857=>"110100100",
  2858=>"000110101",
  2859=>"111101001",
  2860=>"011110001",
  2861=>"000100010",
  2862=>"000000010",
  2863=>"000111010",
  2864=>"111100110",
  2865=>"100011001",
  2866=>"001000011",
  2867=>"001000111",
  2868=>"010011011",
  2869=>"000000000",
  2870=>"011001100",
  2871=>"000001011",
  2872=>"100111110",
  2873=>"000100000",
  2874=>"111010000",
  2875=>"000100000",
  2876=>"010100011",
  2877=>"011011000",
  2878=>"000101100",
  2879=>"110100100",
  2880=>"010110100",
  2881=>"110001111",
  2882=>"010100010",
  2883=>"010101100",
  2884=>"011000010",
  2885=>"110101010",
  2886=>"010000110",
  2887=>"011010010",
  2888=>"100001001",
  2889=>"001001001",
  2890=>"010100010",
  2891=>"110110110",
  2892=>"011011101",
  2893=>"000010110",
  2894=>"010000001",
  2895=>"110000100",
  2896=>"101110111",
  2897=>"111110101",
  2898=>"111101001",
  2899=>"000101011",
  2900=>"010000010",
  2901=>"110011100",
  2902=>"011000110",
  2903=>"000111010",
  2904=>"001000000",
  2905=>"101110000",
  2906=>"110100101",
  2907=>"111111110",
  2908=>"011000011",
  2909=>"010001010",
  2910=>"010001100",
  2911=>"110101101",
  2912=>"100110110",
  2913=>"100011000",
  2914=>"110010000",
  2915=>"111000101",
  2916=>"001110111",
  2917=>"000101000",
  2918=>"001101000",
  2919=>"101110010",
  2920=>"111010000",
  2921=>"001111100",
  2922=>"111101011",
  2923=>"101100001",
  2924=>"100000100",
  2925=>"100101110",
  2926=>"010010101",
  2927=>"011011010",
  2928=>"110001001",
  2929=>"000100001",
  2930=>"101000000",
  2931=>"111100010",
  2932=>"110000110",
  2933=>"100110101",
  2934=>"000001011",
  2935=>"000100011",
  2936=>"001001100",
  2937=>"001010010",
  2938=>"110100000",
  2939=>"100010001",
  2940=>"011100100",
  2941=>"111101110",
  2942=>"100011000",
  2943=>"110100110",
  2944=>"101110110",
  2945=>"101110000",
  2946=>"111100010",
  2947=>"110001100",
  2948=>"101111111",
  2949=>"010011101",
  2950=>"011000110",
  2951=>"011110110",
  2952=>"101111111",
  2953=>"001101110",
  2954=>"000010011",
  2955=>"000111000",
  2956=>"010101100",
  2957=>"011111100",
  2958=>"000010000",
  2959=>"000100101",
  2960=>"001000000",
  2961=>"110001000",
  2962=>"011101110",
  2963=>"111011001",
  2964=>"100101010",
  2965=>"001100110",
  2966=>"011000110",
  2967=>"100000101",
  2968=>"110111011",
  2969=>"111110101",
  2970=>"000111110",
  2971=>"010100111",
  2972=>"111000000",
  2973=>"011101111",
  2974=>"100101000",
  2975=>"011001110",
  2976=>"010000010",
  2977=>"011000001",
  2978=>"010011110",
  2979=>"111011101",
  2980=>"101110110",
  2981=>"100101100",
  2982=>"101010111",
  2983=>"001000111",
  2984=>"000001111",
  2985=>"111110111",
  2986=>"111000010",
  2987=>"100010011",
  2988=>"111000011",
  2989=>"000010110",
  2990=>"111000011",
  2991=>"111000111",
  2992=>"000011111",
  2993=>"110011010",
  2994=>"100100111",
  2995=>"001111010",
  2996=>"100101100",
  2997=>"111101011",
  2998=>"000011101",
  2999=>"100001001",
  3000=>"010001111",
  3001=>"011100011",
  3002=>"101011100",
  3003=>"010110110",
  3004=>"111011011",
  3005=>"010110000",
  3006=>"010010101",
  3007=>"111011011",
  3008=>"110100111",
  3009=>"011101111",
  3010=>"000100110",
  3011=>"111111001",
  3012=>"001110100",
  3013=>"011110111",
  3014=>"011110111",
  3015=>"010111110",
  3016=>"100110100",
  3017=>"000011111",
  3018=>"000111011",
  3019=>"100010111",
  3020=>"001001011",
  3021=>"000101100",
  3022=>"101000111",
  3023=>"110111010",
  3024=>"101000101",
  3025=>"001110000",
  3026=>"001001110",
  3027=>"000111100",
  3028=>"010000000",
  3029=>"111100100",
  3030=>"010100100",
  3031=>"100000000",
  3032=>"111001011",
  3033=>"001001000",
  3034=>"000011101",
  3035=>"010001001",
  3036=>"000011000",
  3037=>"000111101",
  3038=>"101101111",
  3039=>"010000110",
  3040=>"010101111",
  3041=>"011000010",
  3042=>"111101001",
  3043=>"010000100",
  3044=>"110011100",
  3045=>"100011101",
  3046=>"110010101",
  3047=>"111000100",
  3048=>"111101010",
  3049=>"111011110",
  3050=>"100000111",
  3051=>"011011011",
  3052=>"000001000",
  3053=>"001010110",
  3054=>"000110111",
  3055=>"001100000",
  3056=>"101000111",
  3057=>"111000111",
  3058=>"111111011",
  3059=>"110010000",
  3060=>"010010100",
  3061=>"000001101",
  3062=>"011001001",
  3063=>"101100000",
  3064=>"001000000",
  3065=>"101000001",
  3066=>"010101000",
  3067=>"101100110",
  3068=>"001111100",
  3069=>"011011011",
  3070=>"010010001",
  3071=>"011101101",
  3072=>"110100100",
  3073=>"111011101",
  3074=>"000010101",
  3075=>"101111011",
  3076=>"000000001",
  3077=>"100010100",
  3078=>"111010000",
  3079=>"001000010",
  3080=>"011111111",
  3081=>"000000110",
  3082=>"011011010",
  3083=>"001111100",
  3084=>"011100000",
  3085=>"100001111",
  3086=>"011000001",
  3087=>"110000010",
  3088=>"001101100",
  3089=>"110110101",
  3090=>"101110101",
  3091=>"000001000",
  3092=>"111111111",
  3093=>"001000000",
  3094=>"110010101",
  3095=>"101001000",
  3096=>"010011011",
  3097=>"000011000",
  3098=>"101011000",
  3099=>"000010010",
  3100=>"101100111",
  3101=>"110010100",
  3102=>"000111011",
  3103=>"101011011",
  3104=>"010000001",
  3105=>"111100111",
  3106=>"111001100",
  3107=>"001100000",
  3108=>"011101001",
  3109=>"001010110",
  3110=>"100101001",
  3111=>"100011001",
  3112=>"110111110",
  3113=>"011100000",
  3114=>"110001010",
  3115=>"101001111",
  3116=>"000010001",
  3117=>"001000011",
  3118=>"101011010",
  3119=>"101000011",
  3120=>"110101111",
  3121=>"100101011",
  3122=>"010011010",
  3123=>"010000000",
  3124=>"011010101",
  3125=>"011010010",
  3126=>"101011010",
  3127=>"010100101",
  3128=>"100110110",
  3129=>"100001111",
  3130=>"110100110",
  3131=>"011101101",
  3132=>"011001101",
  3133=>"010001110",
  3134=>"110000100",
  3135=>"111001011",
  3136=>"111111011",
  3137=>"101000001",
  3138=>"010010000",
  3139=>"001100001",
  3140=>"001000100",
  3141=>"000110000",
  3142=>"101100101",
  3143=>"100100010",
  3144=>"011011100",
  3145=>"101011000",
  3146=>"101000111",
  3147=>"101010001",
  3148=>"110110110",
  3149=>"101010100",
  3150=>"110110000",
  3151=>"001100010",
  3152=>"111100110",
  3153=>"111001010",
  3154=>"110111011",
  3155=>"111100111",
  3156=>"100001000",
  3157=>"111000010",
  3158=>"001111111",
  3159=>"101100101",
  3160=>"011010111",
  3161=>"100111110",
  3162=>"000111010",
  3163=>"011100000",
  3164=>"101011111",
  3165=>"100000010",
  3166=>"000001010",
  3167=>"100000100",
  3168=>"001011110",
  3169=>"110110111",
  3170=>"110111011",
  3171=>"110110100",
  3172=>"110111000",
  3173=>"100000101",
  3174=>"101110110",
  3175=>"100110001",
  3176=>"001110000",
  3177=>"001001110",
  3178=>"011000111",
  3179=>"100100010",
  3180=>"011101010",
  3181=>"101010100",
  3182=>"010000010",
  3183=>"100111010",
  3184=>"010001001",
  3185=>"001100001",
  3186=>"111101001",
  3187=>"000000111",
  3188=>"110001101",
  3189=>"000110000",
  3190=>"011110101",
  3191=>"110111110",
  3192=>"110010110",
  3193=>"111000100",
  3194=>"000010001",
  3195=>"010001000",
  3196=>"111000101",
  3197=>"001101001",
  3198=>"100000010",
  3199=>"001010011",
  3200=>"110001011",
  3201=>"000110011",
  3202=>"010101010",
  3203=>"010110000",
  3204=>"011011001",
  3205=>"110000110",
  3206=>"011001101",
  3207=>"001001001",
  3208=>"110100110",
  3209=>"101001011",
  3210=>"101000011",
  3211=>"000111100",
  3212=>"111011110",
  3213=>"101110101",
  3214=>"111011101",
  3215=>"100100100",
  3216=>"100110110",
  3217=>"001111100",
  3218=>"001111110",
  3219=>"000000000",
  3220=>"000000001",
  3221=>"110000111",
  3222=>"110101110",
  3223=>"010000101",
  3224=>"011001001",
  3225=>"011111001",
  3226=>"010010010",
  3227=>"111000000",
  3228=>"101101111",
  3229=>"110101110",
  3230=>"000101111",
  3231=>"010110000",
  3232=>"001111101",
  3233=>"000000000",
  3234=>"011111100",
  3235=>"011010101",
  3236=>"010010001",
  3237=>"001110110",
  3238=>"000010101",
  3239=>"011001111",
  3240=>"111101001",
  3241=>"010011000",
  3242=>"110110011",
  3243=>"000011100",
  3244=>"100000011",
  3245=>"110011000",
  3246=>"010010000",
  3247=>"000000100",
  3248=>"100110101",
  3249=>"100010000",
  3250=>"111111101",
  3251=>"100000110",
  3252=>"000011001",
  3253=>"101100010",
  3254=>"101001111",
  3255=>"110011011",
  3256=>"101010110",
  3257=>"111110001",
  3258=>"011010111",
  3259=>"001011001",
  3260=>"000000001",
  3261=>"101111011",
  3262=>"000010100",
  3263=>"100100011",
  3264=>"101110001",
  3265=>"000111101",
  3266=>"010110111",
  3267=>"001011000",
  3268=>"011010000",
  3269=>"110110100",
  3270=>"001011110",
  3271=>"110000001",
  3272=>"110101111",
  3273=>"101110011",
  3274=>"010100000",
  3275=>"000111011",
  3276=>"001111010",
  3277=>"100001101",
  3278=>"100101001",
  3279=>"100110110",
  3280=>"000010001",
  3281=>"010110010",
  3282=>"110011010",
  3283=>"101111111",
  3284=>"001001001",
  3285=>"111101011",
  3286=>"000111011",
  3287=>"110011000",
  3288=>"000111010",
  3289=>"001100101",
  3290=>"110000100",
  3291=>"110111001",
  3292=>"010111111",
  3293=>"100001101",
  3294=>"000001110",
  3295=>"001010111",
  3296=>"100011111",
  3297=>"110011111",
  3298=>"001010000",
  3299=>"111001111",
  3300=>"100111110",
  3301=>"100010000",
  3302=>"000010101",
  3303=>"100000110",
  3304=>"110100100",
  3305=>"010111101",
  3306=>"111110000",
  3307=>"101100111",
  3308=>"100111001",
  3309=>"011101111",
  3310=>"111000001",
  3311=>"000010110",
  3312=>"101101100",
  3313=>"101010001",
  3314=>"101010101",
  3315=>"001011010",
  3316=>"101011101",
  3317=>"100111110",
  3318=>"111001001",
  3319=>"110111010",
  3320=>"100001101",
  3321=>"010110110",
  3322=>"011010110",
  3323=>"011111001",
  3324=>"110111110",
  3325=>"110101001",
  3326=>"110010000",
  3327=>"011000010",
  3328=>"001101000",
  3329=>"110001001",
  3330=>"000000011",
  3331=>"001110100",
  3332=>"100111000",
  3333=>"000100011",
  3334=>"011100110",
  3335=>"101100001",
  3336=>"100101101",
  3337=>"011001011",
  3338=>"000010010",
  3339=>"001001011",
  3340=>"011000010",
  3341=>"110011100",
  3342=>"101000100",
  3343=>"100110000",
  3344=>"111010110",
  3345=>"010010000",
  3346=>"000000100",
  3347=>"111011011",
  3348=>"010010110",
  3349=>"110100000",
  3350=>"000010111",
  3351=>"111100100",
  3352=>"011011011",
  3353=>"110011101",
  3354=>"101100110",
  3355=>"111111010",
  3356=>"001001101",
  3357=>"010010101",
  3358=>"110010111",
  3359=>"101111001",
  3360=>"110111011",
  3361=>"110000111",
  3362=>"111000100",
  3363=>"110101101",
  3364=>"101010011",
  3365=>"101010011",
  3366=>"001000001",
  3367=>"110000011",
  3368=>"001011100",
  3369=>"100010000",
  3370=>"111100110",
  3371=>"011000100",
  3372=>"010110000",
  3373=>"000000000",
  3374=>"111100100",
  3375=>"001010110",
  3376=>"011010111",
  3377=>"100010011",
  3378=>"100110011",
  3379=>"110101001",
  3380=>"010110110",
  3381=>"101000110",
  3382=>"111011101",
  3383=>"000100011",
  3384=>"101100100",
  3385=>"010010001",
  3386=>"101111010",
  3387=>"000011110",
  3388=>"000001000",
  3389=>"000101101",
  3390=>"000111100",
  3391=>"110011101",
  3392=>"011110111",
  3393=>"001011001",
  3394=>"000011010",
  3395=>"011110100",
  3396=>"101010111",
  3397=>"110010000",
  3398=>"110011001",
  3399=>"101100101",
  3400=>"001110101",
  3401=>"010001010",
  3402=>"011111011",
  3403=>"110000100",
  3404=>"001100110",
  3405=>"110111111",
  3406=>"110011101",
  3407=>"001001000",
  3408=>"001011110",
  3409=>"011001000",
  3410=>"000010001",
  3411=>"000000000",
  3412=>"111001001",
  3413=>"010111100",
  3414=>"010011001",
  3415=>"000000001",
  3416=>"011111000",
  3417=>"000100111",
  3418=>"111000100",
  3419=>"011100100",
  3420=>"000011110",
  3421=>"111111010",
  3422=>"001110000",
  3423=>"101101011",
  3424=>"100110100",
  3425=>"110000011",
  3426=>"100000001",
  3427=>"111000110",
  3428=>"000000000",
  3429=>"001001000",
  3430=>"000001000",
  3431=>"111100110",
  3432=>"110101110",
  3433=>"101000100",
  3434=>"111000000",
  3435=>"001101100",
  3436=>"001100011",
  3437=>"010101000",
  3438=>"011010001",
  3439=>"111100110",
  3440=>"110001110",
  3441=>"111110011",
  3442=>"111011111",
  3443=>"000010100",
  3444=>"000001100",
  3445=>"010111100",
  3446=>"111001011",
  3447=>"100100001",
  3448=>"000100101",
  3449=>"101011111",
  3450=>"110100001",
  3451=>"100100110",
  3452=>"010011110",
  3453=>"111011000",
  3454=>"111001011",
  3455=>"001011011",
  3456=>"000010001",
  3457=>"111010110",
  3458=>"101101111",
  3459=>"100001010",
  3460=>"011100110",
  3461=>"100011101",
  3462=>"110000101",
  3463=>"010100101",
  3464=>"110010010",
  3465=>"011011000",
  3466=>"010110011",
  3467=>"001011111",
  3468=>"101000000",
  3469=>"100000001",
  3470=>"101111000",
  3471=>"000100001",
  3472=>"110110000",
  3473=>"000000000",
  3474=>"110101111",
  3475=>"010101001",
  3476=>"110110110",
  3477=>"001111101",
  3478=>"000100101",
  3479=>"110101110",
  3480=>"011100101",
  3481=>"010001000",
  3482=>"111110100",
  3483=>"010001111",
  3484=>"101111000",
  3485=>"100110000",
  3486=>"010111111",
  3487=>"010010100",
  3488=>"100111011",
  3489=>"101001000",
  3490=>"110000101",
  3491=>"000000100",
  3492=>"101001101",
  3493=>"110000100",
  3494=>"011010000",
  3495=>"100111111",
  3496=>"111001010",
  3497=>"000000110",
  3498=>"100010111",
  3499=>"000100110",
  3500=>"110100110",
  3501=>"001000001",
  3502=>"110110011",
  3503=>"000111100",
  3504=>"111101110",
  3505=>"000111111",
  3506=>"001010101",
  3507=>"101101110",
  3508=>"011010110",
  3509=>"000111001",
  3510=>"001000100",
  3511=>"110011001",
  3512=>"011011101",
  3513=>"111011011",
  3514=>"011110111",
  3515=>"110011100",
  3516=>"010010011",
  3517=>"110000001",
  3518=>"011010010",
  3519=>"010100111",
  3520=>"011100011",
  3521=>"001101000",
  3522=>"110111010",
  3523=>"101010011",
  3524=>"111011010",
  3525=>"100110100",
  3526=>"110101111",
  3527=>"100110101",
  3528=>"110100001",
  3529=>"101010010",
  3530=>"110000010",
  3531=>"110011000",
  3532=>"100100100",
  3533=>"100000101",
  3534=>"011111111",
  3535=>"110100001",
  3536=>"000101101",
  3537=>"100001101",
  3538=>"101110111",
  3539=>"000000000",
  3540=>"111111111",
  3541=>"100000101",
  3542=>"010000000",
  3543=>"000100001",
  3544=>"010000101",
  3545=>"000000111",
  3546=>"100011001",
  3547=>"001000110",
  3548=>"001010101",
  3549=>"000110100",
  3550=>"101111010",
  3551=>"111000001",
  3552=>"010110000",
  3553=>"100101010",
  3554=>"000101100",
  3555=>"110110001",
  3556=>"010111001",
  3557=>"100010110",
  3558=>"111100101",
  3559=>"101110001",
  3560=>"111110010",
  3561=>"001011001",
  3562=>"110111011",
  3563=>"010011100",
  3564=>"001001110",
  3565=>"011001111",
  3566=>"110001100",
  3567=>"001101100",
  3568=>"101111110",
  3569=>"100011100",
  3570=>"010101100",
  3571=>"010111000",
  3572=>"011110110",
  3573=>"000110010",
  3574=>"101111000",
  3575=>"110110001",
  3576=>"101110000",
  3577=>"011100011",
  3578=>"110011001",
  3579=>"110111101",
  3580=>"100011111",
  3581=>"100101101",
  3582=>"010010101",
  3583=>"100100101",
  3584=>"011111011",
  3585=>"111101100",
  3586=>"011101101",
  3587=>"001001101",
  3588=>"010001011",
  3589=>"111001110",
  3590=>"110000000",
  3591=>"111111111",
  3592=>"101011001",
  3593=>"101000001",
  3594=>"001001110",
  3595=>"010100000",
  3596=>"010110011",
  3597=>"101000000",
  3598=>"100001000",
  3599=>"000010111",
  3600=>"111001011",
  3601=>"000000100",
  3602=>"010111001",
  3603=>"001001101",
  3604=>"011010001",
  3605=>"000111111",
  3606=>"110101111",
  3607=>"000001001",
  3608=>"110110000",
  3609=>"100100110",
  3610=>"000011111",
  3611=>"000010000",
  3612=>"111101001",
  3613=>"000111010",
  3614=>"101111111",
  3615=>"111101011",
  3616=>"101101000",
  3617=>"000000000",
  3618=>"101001111",
  3619=>"000010111",
  3620=>"111111011",
  3621=>"111111100",
  3622=>"010100011",
  3623=>"110100000",
  3624=>"000110000",
  3625=>"000000000",
  3626=>"010011100",
  3627=>"110111010",
  3628=>"010001100",
  3629=>"111001110",
  3630=>"001011110",
  3631=>"001011101",
  3632=>"110101001",
  3633=>"110111111",
  3634=>"111111110",
  3635=>"010101100",
  3636=>"100110111",
  3637=>"110001110",
  3638=>"110000010",
  3639=>"101110111",
  3640=>"110000100",
  3641=>"111110011",
  3642=>"011110010",
  3643=>"011110100",
  3644=>"110000101",
  3645=>"000001000",
  3646=>"001001010",
  3647=>"110010111",
  3648=>"111110101",
  3649=>"010100001",
  3650=>"001000110",
  3651=>"110110010",
  3652=>"011100011",
  3653=>"111100010",
  3654=>"111000010",
  3655=>"010001110",
  3656=>"010011000",
  3657=>"111100000",
  3658=>"010100010",
  3659=>"101011000",
  3660=>"110111100",
  3661=>"111100110",
  3662=>"111011101",
  3663=>"101101000",
  3664=>"100000001",
  3665=>"111011111",
  3666=>"011101110",
  3667=>"010111011",
  3668=>"101101111",
  3669=>"000101010",
  3670=>"001001100",
  3671=>"000101001",
  3672=>"110011001",
  3673=>"000000001",
  3674=>"110001111",
  3675=>"000001001",
  3676=>"110111110",
  3677=>"010001111",
  3678=>"101100000",
  3679=>"111001010",
  3680=>"111101100",
  3681=>"010010011",
  3682=>"011010011",
  3683=>"101000001",
  3684=>"110010001",
  3685=>"001001100",
  3686=>"010111011",
  3687=>"110001011",
  3688=>"011111111",
  3689=>"000111101",
  3690=>"010000111",
  3691=>"000000000",
  3692=>"111100111",
  3693=>"110001110",
  3694=>"111100011",
  3695=>"001011001",
  3696=>"010000000",
  3697=>"000001011",
  3698=>"010101100",
  3699=>"110010101",
  3700=>"100101111",
  3701=>"010110010",
  3702=>"101001101",
  3703=>"101001000",
  3704=>"011110011",
  3705=>"101111110",
  3706=>"000101100",
  3707=>"001101011",
  3708=>"011001101",
  3709=>"010001101",
  3710=>"110100111",
  3711=>"010001100",
  3712=>"010000010",
  3713=>"010000101",
  3714=>"011101001",
  3715=>"001011101",
  3716=>"111001101",
  3717=>"011110110",
  3718=>"011010000",
  3719=>"100000000",
  3720=>"110111001",
  3721=>"011101111",
  3722=>"111110000",
  3723=>"101001100",
  3724=>"011111001",
  3725=>"110111111",
  3726=>"110101110",
  3727=>"110101101",
  3728=>"011101111",
  3729=>"100101010",
  3730=>"010001111",
  3731=>"100001011",
  3732=>"111000010",
  3733=>"010111101",
  3734=>"111100010",
  3735=>"010011100",
  3736=>"011101011",
  3737=>"110110101",
  3738=>"110010110",
  3739=>"000110010",
  3740=>"010011010",
  3741=>"000100010",
  3742=>"000011101",
  3743=>"100110111",
  3744=>"101100001",
  3745=>"101000001",
  3746=>"000100101",
  3747=>"001011100",
  3748=>"010101011",
  3749=>"011110011",
  3750=>"101111111",
  3751=>"010000110",
  3752=>"001100100",
  3753=>"101011001",
  3754=>"100000001",
  3755=>"000001101",
  3756=>"010110100",
  3757=>"101000101",
  3758=>"000110111",
  3759=>"111101100",
  3760=>"010100000",
  3761=>"010011010",
  3762=>"110111000",
  3763=>"000001010",
  3764=>"111000001",
  3765=>"101111110",
  3766=>"100011010",
  3767=>"001101111",
  3768=>"101110011",
  3769=>"010010111",
  3770=>"001001001",
  3771=>"010110100",
  3772=>"110000001",
  3773=>"001111100",
  3774=>"111010111",
  3775=>"100001010",
  3776=>"011000101",
  3777=>"000110100",
  3778=>"111010100",
  3779=>"010101100",
  3780=>"110101100",
  3781=>"111110100",
  3782=>"001100100",
  3783=>"000000111",
  3784=>"011011011",
  3785=>"110010100",
  3786=>"000000110",
  3787=>"011110100",
  3788=>"101011000",
  3789=>"010011100",
  3790=>"111111011",
  3791=>"011001001",
  3792=>"001011111",
  3793=>"111111100",
  3794=>"000101000",
  3795=>"111001011",
  3796=>"001110101",
  3797=>"111001111",
  3798=>"100101100",
  3799=>"110010110",
  3800=>"111101111",
  3801=>"101011010",
  3802=>"001001000",
  3803=>"100000000",
  3804=>"111101101",
  3805=>"000000011",
  3806=>"100011100",
  3807=>"111001011",
  3808=>"100001011",
  3809=>"100101110",
  3810=>"111111000",
  3811=>"001110000",
  3812=>"000101011",
  3813=>"110000100",
  3814=>"111101111",
  3815=>"101011100",
  3816=>"111101000",
  3817=>"101000000",
  3818=>"000110001",
  3819=>"010001011",
  3820=>"001111001",
  3821=>"110111011",
  3822=>"011011011",
  3823=>"111101011",
  3824=>"011000010",
  3825=>"111001011",
  3826=>"111001001",
  3827=>"100100010",
  3828=>"110011100",
  3829=>"111101010",
  3830=>"110010110",
  3831=>"101101001",
  3832=>"011000011",
  3833=>"110100101",
  3834=>"001011011",
  3835=>"011111001",
  3836=>"100010100",
  3837=>"101111101",
  3838=>"011111010",
  3839=>"001111011",
  3840=>"000001000",
  3841=>"000101001",
  3842=>"010100011",
  3843=>"000001111",
  3844=>"110101110",
  3845=>"110010000",
  3846=>"000101001",
  3847=>"101111101",
  3848=>"011100001",
  3849=>"111010110",
  3850=>"011011110",
  3851=>"010010101",
  3852=>"101100000",
  3853=>"000100011",
  3854=>"101010011",
  3855=>"000100100",
  3856=>"011100010",
  3857=>"101101100",
  3858=>"110111010",
  3859=>"000101111",
  3860=>"101010100",
  3861=>"101010110",
  3862=>"001111100",
  3863=>"101101111",
  3864=>"101001101",
  3865=>"111011100",
  3866=>"110100100",
  3867=>"111110001",
  3868=>"010111010",
  3869=>"011110111",
  3870=>"001100011",
  3871=>"100001011",
  3872=>"101011010",
  3873=>"000100000",
  3874=>"111101111",
  3875=>"101010000",
  3876=>"001110111",
  3877=>"001011000",
  3878=>"011101010",
  3879=>"001011001",
  3880=>"000110111",
  3881=>"000100000",
  3882=>"110101111",
  3883=>"010110111",
  3884=>"101110011",
  3885=>"100110111",
  3886=>"100110111",
  3887=>"101100110",
  3888=>"100010110",
  3889=>"011100011",
  3890=>"000001111",
  3891=>"111101111",
  3892=>"010011110",
  3893=>"001110010",
  3894=>"101100001",
  3895=>"010000100",
  3896=>"101100100",
  3897=>"101101101",
  3898=>"011111011",
  3899=>"011001001",
  3900=>"011110111",
  3901=>"001001010",
  3902=>"101111011",
  3903=>"100111101",
  3904=>"000100110",
  3905=>"100110001",
  3906=>"011011010",
  3907=>"001111101",
  3908=>"101001111",
  3909=>"010011110",
  3910=>"110101010",
  3911=>"101101111",
  3912=>"000111011",
  3913=>"110000101",
  3914=>"000101101",
  3915=>"000101100",
  3916=>"111010110",
  3917=>"101010010",
  3918=>"110111000",
  3919=>"011100001",
  3920=>"111111111",
  3921=>"100101011",
  3922=>"001001000",
  3923=>"110000000",
  3924=>"110000001",
  3925=>"111011110",
  3926=>"100110000",
  3927=>"000000100",
  3928=>"001100101",
  3929=>"101011001",
  3930=>"011000100",
  3931=>"100000111",
  3932=>"010010100",
  3933=>"100001110",
  3934=>"101100000",
  3935=>"111110111",
  3936=>"111100001",
  3937=>"010010111",
  3938=>"100001110",
  3939=>"111101101",
  3940=>"110011101",
  3941=>"100101100",
  3942=>"101000010",
  3943=>"000101001",
  3944=>"111010100",
  3945=>"011001001",
  3946=>"011010110",
  3947=>"011011010",
  3948=>"001000001",
  3949=>"011011100",
  3950=>"110010010",
  3951=>"001011101",
  3952=>"001011100",
  3953=>"111101110",
  3954=>"010011100",
  3955=>"000001000",
  3956=>"111001111",
  3957=>"000000101",
  3958=>"011000101",
  3959=>"001111001",
  3960=>"110000111",
  3961=>"011101110",
  3962=>"100111001",
  3963=>"101100010",
  3964=>"011000100",
  3965=>"101001111",
  3966=>"010010001",
  3967=>"110000101",
  3968=>"100100000",
  3969=>"000100110",
  3970=>"001111000",
  3971=>"000001000",
  3972=>"111101111",
  3973=>"101010000",
  3974=>"000000100",
  3975=>"100001111",
  3976=>"001001101",
  3977=>"001011010",
  3978=>"111110100",
  3979=>"101100111",
  3980=>"001100001",
  3981=>"101010001",
  3982=>"011010010",
  3983=>"000101110",
  3984=>"101111111",
  3985=>"111111100",
  3986=>"110110100",
  3987=>"111111111",
  3988=>"001010100",
  3989=>"110111110",
  3990=>"001111010",
  3991=>"000010010",
  3992=>"111111001",
  3993=>"100101111",
  3994=>"110100100",
  3995=>"111101100",
  3996=>"101001101",
  3997=>"011000010",
  3998=>"111100100",
  3999=>"000110001",
  4000=>"011001000",
  4001=>"001011110",
  4002=>"111000100",
  4003=>"011001101",
  4004=>"110100100",
  4005=>"011101000",
  4006=>"101000111",
  4007=>"010001001",
  4008=>"100011000",
  4009=>"001000101",
  4010=>"010111000",
  4011=>"110100111",
  4012=>"100101111",
  4013=>"101111100",
  4014=>"111110100",
  4015=>"110100001",
  4016=>"100101010",
  4017=>"011000111",
  4018=>"111100101",
  4019=>"000110100",
  4020=>"111110010",
  4021=>"010111100",
  4022=>"110111111",
  4023=>"000011011",
  4024=>"110000001",
  4025=>"011001000",
  4026=>"011100100",
  4027=>"111101111",
  4028=>"011010001",
  4029=>"001011001",
  4030=>"000111000",
  4031=>"011101111",
  4032=>"100000000",
  4033=>"111000100",
  4034=>"111010101",
  4035=>"110011000",
  4036=>"111101011",
  4037=>"101101000",
  4038=>"101111100",
  4039=>"100000011",
  4040=>"100101001",
  4041=>"010100000",
  4042=>"111010100",
  4043=>"000100111",
  4044=>"011011001",
  4045=>"101011100",
  4046=>"111010111",
  4047=>"000010011",
  4048=>"101010010",
  4049=>"110101011",
  4050=>"000000011",
  4051=>"011001100",
  4052=>"000000010",
  4053=>"100000000",
  4054=>"110100101",
  4055=>"101101001",
  4056=>"111011011",
  4057=>"010001001",
  4058=>"110011011",
  4059=>"011000101",
  4060=>"001010001",
  4061=>"010111111",
  4062=>"111000010",
  4063=>"001111110",
  4064=>"100101000",
  4065=>"000000110",
  4066=>"100010010",
  4067=>"000001111",
  4068=>"101101001",
  4069=>"010101010",
  4070=>"110101111",
  4071=>"101001000",
  4072=>"010101100",
  4073=>"000111011",
  4074=>"000100110",
  4075=>"101101111",
  4076=>"110000000",
  4077=>"000000001",
  4078=>"101011101",
  4079=>"001001000",
  4080=>"111111010",
  4081=>"000101000",
  4082=>"100101111",
  4083=>"000111011",
  4084=>"110001111",
  4085=>"011011111",
  4086=>"101100111",
  4087=>"110001011",
  4088=>"001100101",
  4089=>"100100111",
  4090=>"111101110",
  4091=>"001010110",
  4092=>"000111001",
  4093=>"110001111",
  4094=>"001110101",
  4095=>"000000001",
  4096=>"001000001",
  4097=>"100111001",
  4098=>"000010011",
  4099=>"000010111",
  4100=>"010010100",
  4101=>"111000000",
  4102=>"100111100",
  4103=>"010100011",
  4104=>"000100110",
  4105=>"001100000",
  4106=>"100000101",
  4107=>"100001110",
  4108=>"010111011",
  4109=>"111111110",
  4110=>"100000110",
  4111=>"111010000",
  4112=>"001010101",
  4113=>"111110000",
  4114=>"001000000",
  4115=>"110111110",
  4116=>"100110110",
  4117=>"111011101",
  4118=>"111101011",
  4119=>"111100000",
  4120=>"010010111",
  4121=>"111100110",
  4122=>"110011000",
  4123=>"010101111",
  4124=>"100111100",
  4125=>"101011100",
  4126=>"001010110",
  4127=>"111011011",
  4128=>"001000000",
  4129=>"010001111",
  4130=>"001111000",
  4131=>"001110100",
  4132=>"111011111",
  4133=>"110101111",
  4134=>"011100110",
  4135=>"000101000",
  4136=>"110010000",
  4137=>"101101111",
  4138=>"100111000",
  4139=>"010100010",
  4140=>"111111101",
  4141=>"011101101",
  4142=>"010001101",
  4143=>"000110010",
  4144=>"111111111",
  4145=>"110100110",
  4146=>"100011101",
  4147=>"101111100",
  4148=>"111011001",
  4149=>"100111100",
  4150=>"110011110",
  4151=>"110000111",
  4152=>"010001101",
  4153=>"000111010",
  4154=>"001000100",
  4155=>"101111000",
  4156=>"110000100",
  4157=>"101110000",
  4158=>"000101000",
  4159=>"010000111",
  4160=>"101110111",
  4161=>"010001011",
  4162=>"110011101",
  4163=>"110100111",
  4164=>"000000110",
  4165=>"011011011",
  4166=>"101001111",
  4167=>"100110001",
  4168=>"101101100",
  4169=>"101011001",
  4170=>"110011111",
  4171=>"001011111",
  4172=>"111100110",
  4173=>"010000100",
  4174=>"111101001",
  4175=>"100001101",
  4176=>"000001010",
  4177=>"110110110",
  4178=>"011001000",
  4179=>"000101000",
  4180=>"010010000",
  4181=>"111100101",
  4182=>"111111011",
  4183=>"010010001",
  4184=>"110001000",
  4185=>"000110001",
  4186=>"001000000",
  4187=>"001010001",
  4188=>"000000100",
  4189=>"110111011",
  4190=>"101010010",
  4191=>"011000110",
  4192=>"100101001",
  4193=>"000101111",
  4194=>"110100010",
  4195=>"001000111",
  4196=>"101001110",
  4197=>"111010100",
  4198=>"111101111",
  4199=>"010010111",
  4200=>"100011110",
  4201=>"001111110",
  4202=>"100011100",
  4203=>"001000101",
  4204=>"111000000",
  4205=>"111111101",
  4206=>"100000100",
  4207=>"000110000",
  4208=>"101101001",
  4209=>"000010000",
  4210=>"011101011",
  4211=>"001100100",
  4212=>"101001001",
  4213=>"011101001",
  4214=>"011111111",
  4215=>"100000101",
  4216=>"010011100",
  4217=>"000100100",
  4218=>"011111100",
  4219=>"010100001",
  4220=>"101000000",
  4221=>"111110010",
  4222=>"000001000",
  4223=>"010111110",
  4224=>"111001100",
  4225=>"001000000",
  4226=>"111010110",
  4227=>"101001110",
  4228=>"000111111",
  4229=>"110011101",
  4230=>"001010000",
  4231=>"110001100",
  4232=>"011111111",
  4233=>"100100010",
  4234=>"110010000",
  4235=>"010010001",
  4236=>"000001010",
  4237=>"100110101",
  4238=>"010111000",
  4239=>"001000010",
  4240=>"111100101",
  4241=>"011110000",
  4242=>"101011010",
  4243=>"110110011",
  4244=>"011011010",
  4245=>"010101111",
  4246=>"110000011",
  4247=>"101010111",
  4248=>"010100001",
  4249=>"100010100",
  4250=>"110100011",
  4251=>"101110111",
  4252=>"110101011",
  4253=>"101100010",
  4254=>"001001110",
  4255=>"011011001",
  4256=>"000011011",
  4257=>"011101110",
  4258=>"000100101",
  4259=>"110011100",
  4260=>"001001000",
  4261=>"011101100",
  4262=>"101100010",
  4263=>"011001010",
  4264=>"000001010",
  4265=>"011011101",
  4266=>"001000101",
  4267=>"101001011",
  4268=>"011010001",
  4269=>"100110100",
  4270=>"001010111",
  4271=>"000000100",
  4272=>"110011100",
  4273=>"100100010",
  4274=>"000100000",
  4275=>"111000001",
  4276=>"010000100",
  4277=>"110100101",
  4278=>"011101001",
  4279=>"111000010",
  4280=>"011001011",
  4281=>"010111101",
  4282=>"000010000",
  4283=>"010000100",
  4284=>"001010000",
  4285=>"100011101",
  4286=>"001100011",
  4287=>"001000001",
  4288=>"110110000",
  4289=>"000111101",
  4290=>"000011011",
  4291=>"000000010",
  4292=>"101100001",
  4293=>"011100000",
  4294=>"100011101",
  4295=>"101001101",
  4296=>"000001000",
  4297=>"000101001",
  4298=>"111110001",
  4299=>"001011001",
  4300=>"000001110",
  4301=>"010010011",
  4302=>"010010110",
  4303=>"100000000",
  4304=>"010000011",
  4305=>"111000000",
  4306=>"100010101",
  4307=>"111011000",
  4308=>"100111100",
  4309=>"011011011",
  4310=>"101011100",
  4311=>"110111100",
  4312=>"100100011",
  4313=>"000111111",
  4314=>"001100110",
  4315=>"101101000",
  4316=>"011001101",
  4317=>"001110111",
  4318=>"110000101",
  4319=>"100110010",
  4320=>"000100001",
  4321=>"011010100",
  4322=>"110100010",
  4323=>"001101010",
  4324=>"101100110",
  4325=>"110100101",
  4326=>"011011110",
  4327=>"111011000",
  4328=>"001010101",
  4329=>"001100001",
  4330=>"101001000",
  4331=>"011011111",
  4332=>"100000001",
  4333=>"000001111",
  4334=>"011011110",
  4335=>"111110101",
  4336=>"000111011",
  4337=>"100111111",
  4338=>"110100111",
  4339=>"011110111",
  4340=>"000001010",
  4341=>"001000010",
  4342=>"111101111",
  4343=>"000011000",
  4344=>"000010000",
  4345=>"110010000",
  4346=>"111110000",
  4347=>"010001101",
  4348=>"111000011",
  4349=>"110100001",
  4350=>"100111011",
  4351=>"011100000",
  4352=>"100111111",
  4353=>"101111011",
  4354=>"000001001",
  4355=>"000101000",
  4356=>"010110010",
  4357=>"010110001",
  4358=>"111110111",
  4359=>"001100111",
  4360=>"000000000",
  4361=>"000111001",
  4362=>"100010100",
  4363=>"000111001",
  4364=>"000100010",
  4365=>"100011111",
  4366=>"010011110",
  4367=>"000001000",
  4368=>"101110000",
  4369=>"010101101",
  4370=>"001111101",
  4371=>"010100100",
  4372=>"101000011",
  4373=>"110100100",
  4374=>"001001000",
  4375=>"110010111",
  4376=>"001110101",
  4377=>"101000001",
  4378=>"001001011",
  4379=>"111011111",
  4380=>"110111111",
  4381=>"101100101",
  4382=>"010011101",
  4383=>"000011000",
  4384=>"100011011",
  4385=>"001110001",
  4386=>"011100110",
  4387=>"111011111",
  4388=>"001100100",
  4389=>"000100011",
  4390=>"010010001",
  4391=>"111111011",
  4392=>"100010000",
  4393=>"000111000",
  4394=>"011000111",
  4395=>"001001000",
  4396=>"111100011",
  4397=>"110101001",
  4398=>"010001010",
  4399=>"001110000",
  4400=>"110000010",
  4401=>"101001000",
  4402=>"011011101",
  4403=>"000111001",
  4404=>"001101110",
  4405=>"000000000",
  4406=>"001100001",
  4407=>"001000001",
  4408=>"011001101",
  4409=>"010010010",
  4410=>"001011111",
  4411=>"011101111",
  4412=>"000000010",
  4413=>"101110011",
  4414=>"010010010",
  4415=>"001010111",
  4416=>"111111111",
  4417=>"111010100",
  4418=>"100000101",
  4419=>"001101001",
  4420=>"111011101",
  4421=>"011110111",
  4422=>"110110000",
  4423=>"110110000",
  4424=>"010111010",
  4425=>"011110010",
  4426=>"101000110",
  4427=>"000001011",
  4428=>"100110110",
  4429=>"011100100",
  4430=>"000001001",
  4431=>"001001000",
  4432=>"010101010",
  4433=>"111011111",
  4434=>"100000000",
  4435=>"010100111",
  4436=>"000101001",
  4437=>"111111110",
  4438=>"111001111",
  4439=>"111000110",
  4440=>"011111000",
  4441=>"010010000",
  4442=>"010111100",
  4443=>"011101101",
  4444=>"011111000",
  4445=>"101000001",
  4446=>"000101010",
  4447=>"000111100",
  4448=>"000101000",
  4449=>"111001111",
  4450=>"011100001",
  4451=>"010100010",
  4452=>"101010101",
  4453=>"011001010",
  4454=>"000001011",
  4455=>"111111110",
  4456=>"000011011",
  4457=>"011001000",
  4458=>"101111010",
  4459=>"100010001",
  4460=>"011011111",
  4461=>"111000100",
  4462=>"000000001",
  4463=>"110011100",
  4464=>"000011110",
  4465=>"011110000",
  4466=>"111011011",
  4467=>"010000000",
  4468=>"001110010",
  4469=>"101001011",
  4470=>"111011101",
  4471=>"010100010",
  4472=>"100100011",
  4473=>"001001001",
  4474=>"011000001",
  4475=>"000001101",
  4476=>"111011000",
  4477=>"111111111",
  4478=>"111110100",
  4479=>"110101011",
  4480=>"011010101",
  4481=>"001101110",
  4482=>"110010001",
  4483=>"011110111",
  4484=>"001010110",
  4485=>"100101001",
  4486=>"011110111",
  4487=>"010010010",
  4488=>"011101011",
  4489=>"000101000",
  4490=>"110001010",
  4491=>"110101001",
  4492=>"100100101",
  4493=>"100001110",
  4494=>"101000011",
  4495=>"111010111",
  4496=>"110100101",
  4497=>"101101110",
  4498=>"011111100",
  4499=>"111110111",
  4500=>"111000000",
  4501=>"110101101",
  4502=>"001000000",
  4503=>"110111100",
  4504=>"100001010",
  4505=>"000101110",
  4506=>"110100100",
  4507=>"110100000",
  4508=>"110010000",
  4509=>"011011110",
  4510=>"010101101",
  4511=>"100001000",
  4512=>"110100001",
  4513=>"001010001",
  4514=>"011010010",
  4515=>"011100111",
  4516=>"001010111",
  4517=>"101001010",
  4518=>"110111101",
  4519=>"101010011",
  4520=>"000001110",
  4521=>"101111011",
  4522=>"011110111",
  4523=>"100001100",
  4524=>"001111010",
  4525=>"101001001",
  4526=>"011111101",
  4527=>"110000000",
  4528=>"110101011",
  4529=>"011111111",
  4530=>"000000011",
  4531=>"000101001",
  4532=>"111011001",
  4533=>"000001000",
  4534=>"001000101",
  4535=>"010001101",
  4536=>"001101000",
  4537=>"100110000",
  4538=>"000011011",
  4539=>"010001101",
  4540=>"111101010",
  4541=>"001100011",
  4542=>"101111011",
  4543=>"110001111",
  4544=>"000101011",
  4545=>"000010011",
  4546=>"111111011",
  4547=>"101011101",
  4548=>"000000000",
  4549=>"011010011",
  4550=>"011011110",
  4551=>"000110001",
  4552=>"110000100",
  4553=>"001110001",
  4554=>"110010000",
  4555=>"101101000",
  4556=>"000101011",
  4557=>"101101101",
  4558=>"000001111",
  4559=>"000010101",
  4560=>"110110101",
  4561=>"011110100",
  4562=>"100000011",
  4563=>"110010100",
  4564=>"110100111",
  4565=>"110100111",
  4566=>"001110001",
  4567=>"010001100",
  4568=>"111111000",
  4569=>"111111001",
  4570=>"001011000",
  4571=>"010000001",
  4572=>"011000111",
  4573=>"111010000",
  4574=>"111100010",
  4575=>"001100111",
  4576=>"000110101",
  4577=>"001000100",
  4578=>"101101101",
  4579=>"011111011",
  4580=>"000000100",
  4581=>"011011010",
  4582=>"000011011",
  4583=>"000100100",
  4584=>"001101011",
  4585=>"011000010",
  4586=>"000110111",
  4587=>"100010111",
  4588=>"000000000",
  4589=>"011110001",
  4590=>"110111100",
  4591=>"010000110",
  4592=>"001000000",
  4593=>"010110000",
  4594=>"111001100",
  4595=>"110000011",
  4596=>"111111010",
  4597=>"111110101",
  4598=>"010111001",
  4599=>"111100000",
  4600=>"111000100",
  4601=>"110100101",
  4602=>"110111010",
  4603=>"010110010",
  4604=>"000000101",
  4605=>"100101010",
  4606=>"001000000",
  4607=>"101010001",
  4608=>"101000000",
  4609=>"101000001",
  4610=>"011010001",
  4611=>"100011101",
  4612=>"011101110",
  4613=>"000000000",
  4614=>"111101101",
  4615=>"101000011",
  4616=>"000001001",
  4617=>"010101110",
  4618=>"111001000",
  4619=>"110111000",
  4620=>"101100000",
  4621=>"001011101",
  4622=>"100111111",
  4623=>"010100101",
  4624=>"000010011",
  4625=>"101101101",
  4626=>"011101010",
  4627=>"111111110",
  4628=>"110011000",
  4629=>"010100001",
  4630=>"001011111",
  4631=>"001100011",
  4632=>"010000110",
  4633=>"001100010",
  4634=>"100001001",
  4635=>"011011001",
  4636=>"111010111",
  4637=>"010100101",
  4638=>"101100000",
  4639=>"111101000",
  4640=>"101000011",
  4641=>"110010101",
  4642=>"000000110",
  4643=>"111000100",
  4644=>"000001011",
  4645=>"110111101",
  4646=>"011110011",
  4647=>"011000100",
  4648=>"100001111",
  4649=>"010110000",
  4650=>"010111101",
  4651=>"101010100",
  4652=>"010100010",
  4653=>"100001011",
  4654=>"110110000",
  4655=>"111101101",
  4656=>"011001111",
  4657=>"110110110",
  4658=>"101101011",
  4659=>"111010001",
  4660=>"000110011",
  4661=>"010111001",
  4662=>"000010111",
  4663=>"010110010",
  4664=>"011001100",
  4665=>"001011111",
  4666=>"110110011",
  4667=>"011000111",
  4668=>"011001011",
  4669=>"000100000",
  4670=>"001001110",
  4671=>"011101011",
  4672=>"010100001",
  4673=>"001001011",
  4674=>"100100100",
  4675=>"000010011",
  4676=>"111000110",
  4677=>"111010110",
  4678=>"110010100",
  4679=>"000010011",
  4680=>"000100111",
  4681=>"111010010",
  4682=>"010010000",
  4683=>"100001101",
  4684=>"100100011",
  4685=>"111100000",
  4686=>"111111111",
  4687=>"111011101",
  4688=>"011000101",
  4689=>"101010100",
  4690=>"001111101",
  4691=>"101101001",
  4692=>"001100101",
  4693=>"100010001",
  4694=>"101111010",
  4695=>"110100110",
  4696=>"111101010",
  4697=>"110100100",
  4698=>"011011101",
  4699=>"001010111",
  4700=>"011001101",
  4701=>"001110000",
  4702=>"111111001",
  4703=>"001100110",
  4704=>"000100110",
  4705=>"010110110",
  4706=>"011101000",
  4707=>"001100000",
  4708=>"001001111",
  4709=>"111000111",
  4710=>"101111011",
  4711=>"011101110",
  4712=>"010011011",
  4713=>"111011100",
  4714=>"110010000",
  4715=>"010000101",
  4716=>"010101001",
  4717=>"011110110",
  4718=>"011010101",
  4719=>"111101011",
  4720=>"101011010",
  4721=>"000010000",
  4722=>"100110010",
  4723=>"100101111",
  4724=>"010101011",
  4725=>"001011101",
  4726=>"110110101",
  4727=>"110000111",
  4728=>"010100000",
  4729=>"011111000",
  4730=>"111000100",
  4731=>"010110110",
  4732=>"001111000",
  4733=>"111000111",
  4734=>"011111000",
  4735=>"101010001",
  4736=>"110111110",
  4737=>"000100001",
  4738=>"110001010",
  4739=>"010110011",
  4740=>"111110111",
  4741=>"101100111",
  4742=>"011010110",
  4743=>"111111010",
  4744=>"011101000",
  4745=>"100011101",
  4746=>"111011101",
  4747=>"101101110",
  4748=>"001101101",
  4749=>"111111010",
  4750=>"110000010",
  4751=>"100011101",
  4752=>"111101110",
  4753=>"110011100",
  4754=>"010101001",
  4755=>"100011001",
  4756=>"101001110",
  4757=>"110111110",
  4758=>"011011011",
  4759=>"101011100",
  4760=>"010111111",
  4761=>"101110111",
  4762=>"010110110",
  4763=>"011001010",
  4764=>"001011110",
  4765=>"000000110",
  4766=>"000100010",
  4767=>"001101111",
  4768=>"111101011",
  4769=>"110010101",
  4770=>"110100011",
  4771=>"000010111",
  4772=>"110011011",
  4773=>"001111001",
  4774=>"110001000",
  4775=>"000011110",
  4776=>"000111111",
  4777=>"011111100",
  4778=>"011101101",
  4779=>"100010010",
  4780=>"000101111",
  4781=>"111110010",
  4782=>"010110011",
  4783=>"101111000",
  4784=>"101010010",
  4785=>"111101011",
  4786=>"011011101",
  4787=>"111100101",
  4788=>"100010110",
  4789=>"100000101",
  4790=>"100011100",
  4791=>"110011111",
  4792=>"111101011",
  4793=>"010100000",
  4794=>"111000110",
  4795=>"100011110",
  4796=>"011010011",
  4797=>"111100001",
  4798=>"010100101",
  4799=>"110100001",
  4800=>"110000111",
  4801=>"101111110",
  4802=>"110110100",
  4803=>"010100010",
  4804=>"111111101",
  4805=>"000000011",
  4806=>"111011010",
  4807=>"101111000",
  4808=>"101110100",
  4809=>"010011000",
  4810=>"000110101",
  4811=>"100000111",
  4812=>"111011010",
  4813=>"001011000",
  4814=>"111010011",
  4815=>"010010111",
  4816=>"000101111",
  4817=>"100011001",
  4818=>"100010011",
  4819=>"001010011",
  4820=>"111101001",
  4821=>"101010111",
  4822=>"001010100",
  4823=>"000101010",
  4824=>"000111110",
  4825=>"100111111",
  4826=>"111111101",
  4827=>"101100001",
  4828=>"011110000",
  4829=>"011110000",
  4830=>"001111000",
  4831=>"110000011",
  4832=>"100100111",
  4833=>"110000011",
  4834=>"101010000",
  4835=>"010000000",
  4836=>"110010110",
  4837=>"111010011",
  4838=>"100111111",
  4839=>"000011000",
  4840=>"001011010",
  4841=>"110001010",
  4842=>"110101110",
  4843=>"101111101",
  4844=>"010100010",
  4845=>"000010110",
  4846=>"010000010",
  4847=>"111110011",
  4848=>"001001111",
  4849=>"000100110",
  4850=>"010011111",
  4851=>"111011100",
  4852=>"000110000",
  4853=>"111110000",
  4854=>"011011110",
  4855=>"111110110",
  4856=>"111000101",
  4857=>"010011010",
  4858=>"011100101",
  4859=>"101011101",
  4860=>"111110101",
  4861=>"001011010",
  4862=>"011000100",
  4863=>"000010000",
  4864=>"111101011",
  4865=>"110100111",
  4866=>"110001101",
  4867=>"110111001",
  4868=>"100001000",
  4869=>"011010100",
  4870=>"110001001",
  4871=>"011110001",
  4872=>"010001101",
  4873=>"010110001",
  4874=>"100101101",
  4875=>"111111111",
  4876=>"010111001",
  4877=>"101100001",
  4878=>"011110001",
  4879=>"101111111",
  4880=>"000011110",
  4881=>"000000011",
  4882=>"111100111",
  4883=>"100110111",
  4884=>"101100011",
  4885=>"001111100",
  4886=>"101100111",
  4887=>"010011001",
  4888=>"001111101",
  4889=>"100101111",
  4890=>"100100000",
  4891=>"110101110",
  4892=>"111100100",
  4893=>"111110011",
  4894=>"111000000",
  4895=>"000111000",
  4896=>"100111001",
  4897=>"111110111",
  4898=>"000000001",
  4899=>"010011000",
  4900=>"011001011",
  4901=>"010111100",
  4902=>"000011010",
  4903=>"000001000",
  4904=>"010000101",
  4905=>"100001101",
  4906=>"101001010",
  4907=>"001001111",
  4908=>"110100101",
  4909=>"000010111",
  4910=>"000111000",
  4911=>"111111101",
  4912=>"110011011",
  4913=>"000111010",
  4914=>"110100000",
  4915=>"111101010",
  4916=>"111110111",
  4917=>"100110111",
  4918=>"111010011",
  4919=>"111100000",
  4920=>"111100000",
  4921=>"000000001",
  4922=>"001000011",
  4923=>"000100000",
  4924=>"100011001",
  4925=>"000011101",
  4926=>"111100101",
  4927=>"101101101",
  4928=>"110000110",
  4929=>"100110000",
  4930=>"010101100",
  4931=>"101000100",
  4932=>"110011100",
  4933=>"110010010",
  4934=>"000011101",
  4935=>"010111000",
  4936=>"101000000",
  4937=>"101110101",
  4938=>"111001000",
  4939=>"101010110",
  4940=>"000001010",
  4941=>"100100101",
  4942=>"110000110",
  4943=>"110011011",
  4944=>"111010110",
  4945=>"000000001",
  4946=>"100101101",
  4947=>"000000111",
  4948=>"111001000",
  4949=>"110011001",
  4950=>"011000110",
  4951=>"101110000",
  4952=>"010001100",
  4953=>"010001101",
  4954=>"100000110",
  4955=>"101111110",
  4956=>"110010011",
  4957=>"001001110",
  4958=>"111001010",
  4959=>"010010101",
  4960=>"101011000",
  4961=>"001000000",
  4962=>"110010111",
  4963=>"100000010",
  4964=>"110101001",
  4965=>"100001111",
  4966=>"101000001",
  4967=>"111101001",
  4968=>"111110011",
  4969=>"101110011",
  4970=>"001011110",
  4971=>"101100101",
  4972=>"100011111",
  4973=>"010100010",
  4974=>"100000101",
  4975=>"010100000",
  4976=>"111111001",
  4977=>"110100110",
  4978=>"010000100",
  4979=>"001100101",
  4980=>"010011000",
  4981=>"000011000",
  4982=>"000011100",
  4983=>"111011000",
  4984=>"011100100",
  4985=>"110111000",
  4986=>"011001101",
  4987=>"011110101",
  4988=>"010000101",
  4989=>"000000010",
  4990=>"011100111",
  4991=>"010010110",
  4992=>"000111100",
  4993=>"101000100",
  4994=>"100111010",
  4995=>"001011101",
  4996=>"100101001",
  4997=>"110110111",
  4998=>"100011001",
  4999=>"111001011",
  5000=>"100111000",
  5001=>"110011101",
  5002=>"010000000",
  5003=>"110111110",
  5004=>"110001001",
  5005=>"010101100",
  5006=>"111000110",
  5007=>"001101001",
  5008=>"011001011",
  5009=>"111101011",
  5010=>"100111101",
  5011=>"010101000",
  5012=>"100011100",
  5013=>"000101100",
  5014=>"011011000",
  5015=>"011010100",
  5016=>"100100000",
  5017=>"000010010",
  5018=>"001011111",
  5019=>"011000100",
  5020=>"010000010",
  5021=>"100110111",
  5022=>"110000111",
  5023=>"111011100",
  5024=>"111000000",
  5025=>"110100000",
  5026=>"000001111",
  5027=>"111011111",
  5028=>"010110111",
  5029=>"011110101",
  5030=>"000110110",
  5031=>"010000000",
  5032=>"010100111",
  5033=>"000110010",
  5034=>"100010010",
  5035=>"100100011",
  5036=>"000011000",
  5037=>"111100110",
  5038=>"111000100",
  5039=>"000011000",
  5040=>"100010111",
  5041=>"010000011",
  5042=>"011000100",
  5043=>"010111011",
  5044=>"000111010",
  5045=>"011111101",
  5046=>"110101010",
  5047=>"111110110",
  5048=>"111101010",
  5049=>"111011011",
  5050=>"010111111",
  5051=>"100000110",
  5052=>"101111111",
  5053=>"010101111",
  5054=>"000101001",
  5055=>"111100100",
  5056=>"111010000",
  5057=>"000100000",
  5058=>"101111110",
  5059=>"100110100",
  5060=>"101001100",
  5061=>"001111011",
  5062=>"010001101",
  5063=>"010001001",
  5064=>"111000001",
  5065=>"001001001",
  5066=>"111001011",
  5067=>"010110110",
  5068=>"001010000",
  5069=>"000100100",
  5070=>"111011111",
  5071=>"000100011",
  5072=>"100101101",
  5073=>"111000010",
  5074=>"001110010",
  5075=>"000010010",
  5076=>"111111111",
  5077=>"101101001",
  5078=>"100010010",
  5079=>"000001110",
  5080=>"011000101",
  5081=>"101000101",
  5082=>"011110111",
  5083=>"001001001",
  5084=>"001010000",
  5085=>"001001110",
  5086=>"101001111",
  5087=>"101001101",
  5088=>"010110010",
  5089=>"110110110",
  5090=>"111100011",
  5091=>"000000010",
  5092=>"001010110",
  5093=>"100001010",
  5094=>"001000011",
  5095=>"111101111",
  5096=>"000101001",
  5097=>"001011000",
  5098=>"101001001",
  5099=>"100110010",
  5100=>"011011111",
  5101=>"011000011",
  5102=>"001110110",
  5103=>"010101001",
  5104=>"010101011",
  5105=>"101111000",
  5106=>"100100000",
  5107=>"000100100",
  5108=>"110011101",
  5109=>"010000100",
  5110=>"100000001",
  5111=>"001111001",
  5112=>"001110111",
  5113=>"101000100",
  5114=>"111001001",
  5115=>"001110001",
  5116=>"000000111",
  5117=>"100001110",
  5118=>"010011011",
  5119=>"011000001",
  5120=>"000000001",
  5121=>"111100000",
  5122=>"111011001",
  5123=>"100011101",
  5124=>"000011100",
  5125=>"000000010",
  5126=>"110110000",
  5127=>"100111011",
  5128=>"010010101",
  5129=>"101111011",
  5130=>"011011100",
  5131=>"010101110",
  5132=>"110011000",
  5133=>"000011101",
  5134=>"111111111",
  5135=>"111101000",
  5136=>"101000011",
  5137=>"001100101",
  5138=>"101110010",
  5139=>"000010001",
  5140=>"000110110",
  5141=>"010100010",
  5142=>"000010001",
  5143=>"111111010",
  5144=>"001010110",
  5145=>"010101111",
  5146=>"100011011",
  5147=>"011010001",
  5148=>"111001011",
  5149=>"001111011",
  5150=>"001000111",
  5151=>"101111011",
  5152=>"110111011",
  5153=>"000010111",
  5154=>"111101000",
  5155=>"000001001",
  5156=>"001110101",
  5157=>"111000100",
  5158=>"000111110",
  5159=>"100001001",
  5160=>"101000111",
  5161=>"111000010",
  5162=>"110101111",
  5163=>"101010011",
  5164=>"010110000",
  5165=>"111000010",
  5166=>"000000011",
  5167=>"111111001",
  5168=>"000000001",
  5169=>"100010000",
  5170=>"100101100",
  5171=>"000111000",
  5172=>"100011010",
  5173=>"100101000",
  5174=>"000000001",
  5175=>"001001111",
  5176=>"111111010",
  5177=>"110110100",
  5178=>"110011010",
  5179=>"001111000",
  5180=>"000100101",
  5181=>"010001111",
  5182=>"111100001",
  5183=>"100001010",
  5184=>"111010101",
  5185=>"100011001",
  5186=>"011010000",
  5187=>"010101010",
  5188=>"111011001",
  5189=>"100000011",
  5190=>"111100111",
  5191=>"011100111",
  5192=>"100010101",
  5193=>"110010010",
  5194=>"000001000",
  5195=>"101111101",
  5196=>"000010101",
  5197=>"001110111",
  5198=>"110100100",
  5199=>"111101111",
  5200=>"101110000",
  5201=>"000011111",
  5202=>"101111000",
  5203=>"011110001",
  5204=>"001111010",
  5205=>"001010111",
  5206=>"111111000",
  5207=>"111100010",
  5208=>"110110110",
  5209=>"011010010",
  5210=>"001111010",
  5211=>"100101101",
  5212=>"010000111",
  5213=>"110111010",
  5214=>"001010100",
  5215=>"010000000",
  5216=>"000011001",
  5217=>"001101111",
  5218=>"110100100",
  5219=>"111001000",
  5220=>"001001010",
  5221=>"110001100",
  5222=>"000001111",
  5223=>"101010001",
  5224=>"101011001",
  5225=>"000101111",
  5226=>"011001010",
  5227=>"010111100",
  5228=>"011111000",
  5229=>"111001101",
  5230=>"001110110",
  5231=>"000101101",
  5232=>"100100010",
  5233=>"100011100",
  5234=>"010010010",
  5235=>"000100000",
  5236=>"011001110",
  5237=>"111011001",
  5238=>"111110010",
  5239=>"010000011",
  5240=>"100101101",
  5241=>"111010010",
  5242=>"000000100",
  5243=>"011110011",
  5244=>"010101011",
  5245=>"111001000",
  5246=>"101000100",
  5247=>"000000101",
  5248=>"111111111",
  5249=>"100111110",
  5250=>"010010101",
  5251=>"101101101",
  5252=>"001111000",
  5253=>"111010110",
  5254=>"101000000",
  5255=>"010100001",
  5256=>"011001100",
  5257=>"000101010",
  5258=>"000101100",
  5259=>"100111010",
  5260=>"011100011",
  5261=>"101111010",
  5262=>"001111000",
  5263=>"011100111",
  5264=>"000011110",
  5265=>"100000110",
  5266=>"001111001",
  5267=>"111011110",
  5268=>"110111001",
  5269=>"101010111",
  5270=>"110111010",
  5271=>"010101000",
  5272=>"111111011",
  5273=>"010110001",
  5274=>"101000001",
  5275=>"001110000",
  5276=>"001011010",
  5277=>"000001010",
  5278=>"000000000",
  5279=>"100111111",
  5280=>"000001100",
  5281=>"110111011",
  5282=>"111100011",
  5283=>"100011110",
  5284=>"111000101",
  5285=>"011110100",
  5286=>"100101110",
  5287=>"110111100",
  5288=>"110101010",
  5289=>"000101111",
  5290=>"111111000",
  5291=>"010010100",
  5292=>"000110001",
  5293=>"100111100",
  5294=>"110110101",
  5295=>"001111000",
  5296=>"001001101",
  5297=>"000000000",
  5298=>"011011100",
  5299=>"010100000",
  5300=>"001111111",
  5301=>"001000000",
  5302=>"101010010",
  5303=>"111011111",
  5304=>"011110101",
  5305=>"010011011",
  5306=>"110010110",
  5307=>"110111110",
  5308=>"101110011",
  5309=>"011001101",
  5310=>"111010010",
  5311=>"011110001",
  5312=>"000011101",
  5313=>"011111110",
  5314=>"100100011",
  5315=>"111100001",
  5316=>"100100101",
  5317=>"111111101",
  5318=>"100100010",
  5319=>"101111100",
  5320=>"100100011",
  5321=>"100111001",
  5322=>"011111001",
  5323=>"010010101",
  5324=>"001000110",
  5325=>"000010001",
  5326=>"101100010",
  5327=>"100101010",
  5328=>"000110111",
  5329=>"001100111",
  5330=>"000100010",
  5331=>"011101111",
  5332=>"110111111",
  5333=>"101101001",
  5334=>"001011001",
  5335=>"110010101",
  5336=>"000011010",
  5337=>"000011100",
  5338=>"001100010",
  5339=>"011001101",
  5340=>"010010111",
  5341=>"000111001",
  5342=>"101100010",
  5343=>"110001111",
  5344=>"111101110",
  5345=>"000011000",
  5346=>"111111111",
  5347=>"110010111",
  5348=>"111101001",
  5349=>"010001110",
  5350=>"011101011",
  5351=>"111100101",
  5352=>"111010011",
  5353=>"110000011",
  5354=>"100111010",
  5355=>"100001000",
  5356=>"110010100",
  5357=>"100000110",
  5358=>"101011001",
  5359=>"110001111",
  5360=>"101001111",
  5361=>"011111010",
  5362=>"000010011",
  5363=>"000011101",
  5364=>"001001101",
  5365=>"100001101",
  5366=>"011010001",
  5367=>"100111010",
  5368=>"010000100",
  5369=>"011010111",
  5370=>"000100111",
  5371=>"000110001",
  5372=>"000011001",
  5373=>"001000010",
  5374=>"110001110",
  5375=>"010000001",
  5376=>"011111100",
  5377=>"111000011",
  5378=>"111011001",
  5379=>"100111100",
  5380=>"101100000",
  5381=>"110110111",
  5382=>"100110111",
  5383=>"000111011",
  5384=>"101001010",
  5385=>"110110101",
  5386=>"010110000",
  5387=>"001001001",
  5388=>"110010000",
  5389=>"111101101",
  5390=>"101110110",
  5391=>"000011010",
  5392=>"101100010",
  5393=>"001111111",
  5394=>"011101010",
  5395=>"111001000",
  5396=>"001101011",
  5397=>"111110000",
  5398=>"100000111",
  5399=>"101111101",
  5400=>"111001000",
  5401=>"000000001",
  5402=>"000111010",
  5403=>"001000001",
  5404=>"001100100",
  5405=>"001011011",
  5406=>"110111001",
  5407=>"000011100",
  5408=>"100111000",
  5409=>"000101011",
  5410=>"111001110",
  5411=>"101110111",
  5412=>"110011011",
  5413=>"111111100",
  5414=>"101010011",
  5415=>"000001001",
  5416=>"101001001",
  5417=>"111110100",
  5418=>"111110111",
  5419=>"100110101",
  5420=>"001101101",
  5421=>"111110110",
  5422=>"000100100",
  5423=>"000000100",
  5424=>"010010110",
  5425=>"011000101",
  5426=>"000000101",
  5427=>"000010001",
  5428=>"110100010",
  5429=>"110110011",
  5430=>"110011010",
  5431=>"000010011",
  5432=>"000000100",
  5433=>"101110101",
  5434=>"101111110",
  5435=>"010101101",
  5436=>"110110011",
  5437=>"001011111",
  5438=>"000110000",
  5439=>"111000110",
  5440=>"100001111",
  5441=>"110111010",
  5442=>"111100010",
  5443=>"100000110",
  5444=>"010111000",
  5445=>"000111100",
  5446=>"101100011",
  5447=>"010111010",
  5448=>"001101111",
  5449=>"001000001",
  5450=>"100100000",
  5451=>"010110011",
  5452=>"110000001",
  5453=>"111110111",
  5454=>"101101110",
  5455=>"111011000",
  5456=>"100110110",
  5457=>"100010100",
  5458=>"000001110",
  5459=>"100100010",
  5460=>"000010000",
  5461=>"001110010",
  5462=>"110001011",
  5463=>"001100011",
  5464=>"001100011",
  5465=>"000111000",
  5466=>"110111001",
  5467=>"001010000",
  5468=>"000000000",
  5469=>"001001010",
  5470=>"101111101",
  5471=>"111011011",
  5472=>"101100010",
  5473=>"000110110",
  5474=>"000010000",
  5475=>"000000011",
  5476=>"011111101",
  5477=>"000000010",
  5478=>"100011011",
  5479=>"010000011",
  5480=>"000010011",
  5481=>"000101011",
  5482=>"100011001",
  5483=>"001000001",
  5484=>"111000100",
  5485=>"000101111",
  5486=>"111100000",
  5487=>"000000000",
  5488=>"010000110",
  5489=>"110101001",
  5490=>"110011101",
  5491=>"110010010",
  5492=>"100110010",
  5493=>"001010010",
  5494=>"111110101",
  5495=>"000001111",
  5496=>"101001001",
  5497=>"001000001",
  5498=>"111011001",
  5499=>"000100011",
  5500=>"111011001",
  5501=>"001001011",
  5502=>"101000110",
  5503=>"101011110",
  5504=>"101010000",
  5505=>"100110100",
  5506=>"110010100",
  5507=>"100110001",
  5508=>"001111101",
  5509=>"101011010",
  5510=>"011000101",
  5511=>"101000010",
  5512=>"100000000",
  5513=>"000010000",
  5514=>"001011001",
  5515=>"000000101",
  5516=>"010010000",
  5517=>"101011011",
  5518=>"000001010",
  5519=>"100111101",
  5520=>"110111100",
  5521=>"111000111",
  5522=>"010011111",
  5523=>"011100010",
  5524=>"100011101",
  5525=>"110110001",
  5526=>"110001111",
  5527=>"001001111",
  5528=>"101001110",
  5529=>"000100110",
  5530=>"110101011",
  5531=>"000010100",
  5532=>"011101010",
  5533=>"010111010",
  5534=>"101010011",
  5535=>"000000001",
  5536=>"001010000",
  5537=>"001011000",
  5538=>"001110100",
  5539=>"010001101",
  5540=>"010111101",
  5541=>"001100101",
  5542=>"100100000",
  5543=>"000100001",
  5544=>"110000110",
  5545=>"101111101",
  5546=>"111101000",
  5547=>"000011011",
  5548=>"001000000",
  5549=>"001100011",
  5550=>"001001000",
  5551=>"010100111",
  5552=>"010010010",
  5553=>"001001100",
  5554=>"101001101",
  5555=>"101110000",
  5556=>"000010010",
  5557=>"010001110",
  5558=>"101000011",
  5559=>"111111010",
  5560=>"000001000",
  5561=>"001100000",
  5562=>"010000000",
  5563=>"000100111",
  5564=>"000011010",
  5565=>"001110011",
  5566=>"001110010",
  5567=>"011010000",
  5568=>"011011100",
  5569=>"001110010",
  5570=>"010101101",
  5571=>"011011100",
  5572=>"100101100",
  5573=>"010101110",
  5574=>"010111101",
  5575=>"100010100",
  5576=>"111110110",
  5577=>"100110001",
  5578=>"011000001",
  5579=>"100001101",
  5580=>"100011110",
  5581=>"101000001",
  5582=>"010000101",
  5583=>"011010101",
  5584=>"011001010",
  5585=>"101111111",
  5586=>"001111101",
  5587=>"111111101",
  5588=>"111010101",
  5589=>"001010010",
  5590=>"100101000",
  5591=>"000001101",
  5592=>"110101000",
  5593=>"110001000",
  5594=>"011110110",
  5595=>"110110101",
  5596=>"011111110",
  5597=>"110100010",
  5598=>"110111100",
  5599=>"111000001",
  5600=>"110000000",
  5601=>"000101110",
  5602=>"000100010",
  5603=>"000001001",
  5604=>"110101111",
  5605=>"100110011",
  5606=>"011001100",
  5607=>"010001001",
  5608=>"101110011",
  5609=>"001110110",
  5610=>"000000111",
  5611=>"110110100",
  5612=>"110010110",
  5613=>"000001011",
  5614=>"110001010",
  5615=>"101000010",
  5616=>"111010001",
  5617=>"010100000",
  5618=>"100010111",
  5619=>"101000110",
  5620=>"110011110",
  5621=>"110010100",
  5622=>"010100111",
  5623=>"011000111",
  5624=>"111110011",
  5625=>"001100101",
  5626=>"000100000",
  5627=>"111100011",
  5628=>"010011000",
  5629=>"000000001",
  5630=>"111101101",
  5631=>"001111001",
  5632=>"001010101",
  5633=>"011000001",
  5634=>"101100011",
  5635=>"001100100",
  5636=>"101111111",
  5637=>"111011001",
  5638=>"011110110",
  5639=>"101001111",
  5640=>"110000001",
  5641=>"100110101",
  5642=>"100100111",
  5643=>"000001100",
  5644=>"101000011",
  5645=>"100001100",
  5646=>"000111001",
  5647=>"110101111",
  5648=>"100111000",
  5649=>"010011111",
  5650=>"101110110",
  5651=>"001001101",
  5652=>"000100111",
  5653=>"000000010",
  5654=>"010101100",
  5655=>"100111110",
  5656=>"111100011",
  5657=>"111111001",
  5658=>"101011111",
  5659=>"011100100",
  5660=>"000101100",
  5661=>"000000000",
  5662=>"011000111",
  5663=>"101000001",
  5664=>"111111111",
  5665=>"000011110",
  5666=>"100101100",
  5667=>"000100110",
  5668=>"101101110",
  5669=>"101100101",
  5670=>"010110111",
  5671=>"000000111",
  5672=>"010001000",
  5673=>"110101101",
  5674=>"000101000",
  5675=>"100001110",
  5676=>"100100011",
  5677=>"101001010",
  5678=>"100001011",
  5679=>"101100000",
  5680=>"100011110",
  5681=>"101100011",
  5682=>"010011011",
  5683=>"101110011",
  5684=>"110001100",
  5685=>"100110101",
  5686=>"011001010",
  5687=>"001001100",
  5688=>"110010010",
  5689=>"011010110",
  5690=>"000110111",
  5691=>"101010011",
  5692=>"101100111",
  5693=>"101110001",
  5694=>"111110111",
  5695=>"111001100",
  5696=>"111111110",
  5697=>"111000011",
  5698=>"000011101",
  5699=>"011011111",
  5700=>"101001101",
  5701=>"111110011",
  5702=>"000001011",
  5703=>"110101100",
  5704=>"010011101",
  5705=>"110111100",
  5706=>"111101101",
  5707=>"111101000",
  5708=>"000110011",
  5709=>"110001011",
  5710=>"111001111",
  5711=>"100100110",
  5712=>"111110111",
  5713=>"011000011",
  5714=>"101111011",
  5715=>"000000000",
  5716=>"100011011",
  5717=>"111010110",
  5718=>"110101011",
  5719=>"100010011",
  5720=>"101011011",
  5721=>"000011111",
  5722=>"101001011",
  5723=>"000000000",
  5724=>"000010011",
  5725=>"001010111",
  5726=>"111101010",
  5727=>"110000010",
  5728=>"011001101",
  5729=>"000110100",
  5730=>"110110011",
  5731=>"000010000",
  5732=>"011101000",
  5733=>"001010000",
  5734=>"110010100",
  5735=>"111110000",
  5736=>"001011100",
  5737=>"110110110",
  5738=>"001010101",
  5739=>"010011001",
  5740=>"000010000",
  5741=>"101001100",
  5742=>"100101111",
  5743=>"000000100",
  5744=>"110011001",
  5745=>"000101100",
  5746=>"111010110",
  5747=>"001000111",
  5748=>"111011000",
  5749=>"010011000",
  5750=>"011010100",
  5751=>"111101000",
  5752=>"110010011",
  5753=>"010001010",
  5754=>"101000100",
  5755=>"001000100",
  5756=>"011011001",
  5757=>"100001100",
  5758=>"000101011",
  5759=>"110111010",
  5760=>"000001101",
  5761=>"101100010",
  5762=>"110000010",
  5763=>"100110010",
  5764=>"110101111",
  5765=>"100010000",
  5766=>"100110111",
  5767=>"000011111",
  5768=>"000001000",
  5769=>"101110010",
  5770=>"000110010",
  5771=>"101100100",
  5772=>"010001000",
  5773=>"100011010",
  5774=>"001010010",
  5775=>"111011110",
  5776=>"111010010",
  5777=>"011101011",
  5778=>"100000100",
  5779=>"001011000",
  5780=>"010000011",
  5781=>"100111001",
  5782=>"000100111",
  5783=>"001101111",
  5784=>"111011101",
  5785=>"001011111",
  5786=>"000000001",
  5787=>"110111001",
  5788=>"001110110",
  5789=>"100110011",
  5790=>"111011000",
  5791=>"001111111",
  5792=>"000000000",
  5793=>"110001100",
  5794=>"111111111",
  5795=>"010100001",
  5796=>"010111111",
  5797=>"110001111",
  5798=>"111111111",
  5799=>"000000101",
  5800=>"011011010",
  5801=>"110000111",
  5802=>"000011100",
  5803=>"010001111",
  5804=>"100100000",
  5805=>"101100110",
  5806=>"100011011",
  5807=>"111111111",
  5808=>"000000100",
  5809=>"101101100",
  5810=>"100111011",
  5811=>"110011100",
  5812=>"011011101",
  5813=>"101110110",
  5814=>"101001001",
  5815=>"001101001",
  5816=>"101111101",
  5817=>"100000001",
  5818=>"101011001",
  5819=>"011011000",
  5820=>"111110000",
  5821=>"101111110",
  5822=>"001000111",
  5823=>"010110101",
  5824=>"101110001",
  5825=>"001110010",
  5826=>"011011010",
  5827=>"000000001",
  5828=>"000011010",
  5829=>"010001001",
  5830=>"101000110",
  5831=>"110000100",
  5832=>"111011101",
  5833=>"011110111",
  5834=>"101001111",
  5835=>"100101111",
  5836=>"000111100",
  5837=>"110100111",
  5838=>"000010110",
  5839=>"100000100",
  5840=>"111110110",
  5841=>"001010001",
  5842=>"111100111",
  5843=>"001001110",
  5844=>"010000001",
  5845=>"001001100",
  5846=>"011101100",
  5847=>"100111010",
  5848=>"100001000",
  5849=>"100000100",
  5850=>"001000001",
  5851=>"000011101",
  5852=>"100000001",
  5853=>"001011100",
  5854=>"100111001",
  5855=>"110111010",
  5856=>"111111111",
  5857=>"001011100",
  5858=>"111100000",
  5859=>"001111100",
  5860=>"110010100",
  5861=>"101010101",
  5862=>"011001001",
  5863=>"001010110",
  5864=>"001101011",
  5865=>"100111000",
  5866=>"011011011",
  5867=>"011000011",
  5868=>"000001001",
  5869=>"100111010",
  5870=>"110101111",
  5871=>"111111000",
  5872=>"011001010",
  5873=>"110011010",
  5874=>"010010000",
  5875=>"010010110",
  5876=>"101010010",
  5877=>"101110001",
  5878=>"100101101",
  5879=>"001011111",
  5880=>"111010101",
  5881=>"101110010",
  5882=>"000011110",
  5883=>"000000011",
  5884=>"000110110",
  5885=>"101000101",
  5886=>"001110101",
  5887=>"000000100",
  5888=>"000010000",
  5889=>"011111001",
  5890=>"100010101",
  5891=>"101101001",
  5892=>"000101101",
  5893=>"011011001",
  5894=>"011110010",
  5895=>"011011111",
  5896=>"101000000",
  5897=>"001000100",
  5898=>"101010101",
  5899=>"100001110",
  5900=>"010100101",
  5901=>"001000001",
  5902=>"110110011",
  5903=>"100011111",
  5904=>"010111101",
  5905=>"100110011",
  5906=>"100011000",
  5907=>"000100000",
  5908=>"100101101",
  5909=>"101010110",
  5910=>"001101010",
  5911=>"101110000",
  5912=>"000000010",
  5913=>"010010110",
  5914=>"000110001",
  5915=>"000111011",
  5916=>"111110000",
  5917=>"011001100",
  5918=>"000100001",
  5919=>"111101000",
  5920=>"111111011",
  5921=>"001101111",
  5922=>"110101000",
  5923=>"011110111",
  5924=>"101111000",
  5925=>"010010110",
  5926=>"000100100",
  5927=>"101001100",
  5928=>"110100110",
  5929=>"001001100",
  5930=>"110111111",
  5931=>"010101100",
  5932=>"011011110",
  5933=>"110110111",
  5934=>"010001010",
  5935=>"000011111",
  5936=>"010001100",
  5937=>"110101101",
  5938=>"111010001",
  5939=>"011101010",
  5940=>"010000100",
  5941=>"111110010",
  5942=>"100010111",
  5943=>"000101001",
  5944=>"000111111",
  5945=>"001010010",
  5946=>"111101010",
  5947=>"111001100",
  5948=>"010010000",
  5949=>"000111110",
  5950=>"000110000",
  5951=>"001100000",
  5952=>"000101001",
  5953=>"011011111",
  5954=>"011000101",
  5955=>"101000000",
  5956=>"001100110",
  5957=>"001110111",
  5958=>"100000111",
  5959=>"001110011",
  5960=>"010101010",
  5961=>"100101100",
  5962=>"101110000",
  5963=>"001000000",
  5964=>"001100010",
  5965=>"100111110",
  5966=>"111011010",
  5967=>"001001000",
  5968=>"000001001",
  5969=>"011111101",
  5970=>"110011110",
  5971=>"100111101",
  5972=>"101101111",
  5973=>"010011011",
  5974=>"001000000",
  5975=>"000111100",
  5976=>"100111110",
  5977=>"000100101",
  5978=>"000000101",
  5979=>"100011010",
  5980=>"100000110",
  5981=>"110100111",
  5982=>"111100100",
  5983=>"100100011",
  5984=>"001100011",
  5985=>"111101011",
  5986=>"111110000",
  5987=>"100010011",
  5988=>"110001010",
  5989=>"110000000",
  5990=>"111100011",
  5991=>"110010010",
  5992=>"010000000",
  5993=>"110001101",
  5994=>"001111010",
  5995=>"100100000",
  5996=>"010010010",
  5997=>"111001000",
  5998=>"111001011",
  5999=>"010100001",
  6000=>"000011110",
  6001=>"101111101",
  6002=>"101010110",
  6003=>"011111000",
  6004=>"101011100",
  6005=>"001010101",
  6006=>"000010010",
  6007=>"010101001",
  6008=>"101100010",
  6009=>"010010100",
  6010=>"011110111",
  6011=>"100011010",
  6012=>"100111100",
  6013=>"111100011",
  6014=>"110101111",
  6015=>"111001001",
  6016=>"011101111",
  6017=>"111111000",
  6018=>"111111010",
  6019=>"100000000",
  6020=>"100100101",
  6021=>"000100110",
  6022=>"110111000",
  6023=>"000100011",
  6024=>"011000010",
  6025=>"111101111",
  6026=>"110111101",
  6027=>"001110111",
  6028=>"100001111",
  6029=>"101101001",
  6030=>"111111010",
  6031=>"000100000",
  6032=>"011111111",
  6033=>"101100000",
  6034=>"000111101",
  6035=>"000110001",
  6036=>"111000100",
  6037=>"011101001",
  6038=>"001000011",
  6039=>"010111110",
  6040=>"111010111",
  6041=>"111001011",
  6042=>"000001100",
  6043=>"000101001",
  6044=>"100010111",
  6045=>"100011000",
  6046=>"110001010",
  6047=>"000010010",
  6048=>"010000110",
  6049=>"010011110",
  6050=>"101100001",
  6051=>"101110000",
  6052=>"010001111",
  6053=>"111100111",
  6054=>"110111011",
  6055=>"110001010",
  6056=>"000111001",
  6057=>"001011100",
  6058=>"111010010",
  6059=>"011010101",
  6060=>"000000010",
  6061=>"100000111",
  6062=>"011101110",
  6063=>"001010110",
  6064=>"011100011",
  6065=>"110100010",
  6066=>"100011100",
  6067=>"100011001",
  6068=>"010100000",
  6069=>"001000000",
  6070=>"001101111",
  6071=>"001010011",
  6072=>"111110101",
  6073=>"110011111",
  6074=>"111111111",
  6075=>"111010000",
  6076=>"111011011",
  6077=>"011001000",
  6078=>"011011100",
  6079=>"000110010",
  6080=>"110001001",
  6081=>"011011000",
  6082=>"010110101",
  6083=>"000001010",
  6084=>"110010000",
  6085=>"000111111",
  6086=>"100001001",
  6087=>"110100011",
  6088=>"100100110",
  6089=>"101111110",
  6090=>"011000100",
  6091=>"111101110",
  6092=>"111110100",
  6093=>"101100110",
  6094=>"111000000",
  6095=>"000110111",
  6096=>"110110011",
  6097=>"001110001",
  6098=>"000110000",
  6099=>"011101111",
  6100=>"011100001",
  6101=>"110100101",
  6102=>"000011011",
  6103=>"111010011",
  6104=>"010011101",
  6105=>"111101101",
  6106=>"100101011",
  6107=>"100110101",
  6108=>"010111110",
  6109=>"010101111",
  6110=>"100110101",
  6111=>"000001001",
  6112=>"000010111",
  6113=>"000000000",
  6114=>"001001000",
  6115=>"111110001",
  6116=>"010101100",
  6117=>"110100000",
  6118=>"001101100",
  6119=>"100110010",
  6120=>"111101001",
  6121=>"111110100",
  6122=>"111001111",
  6123=>"111110011",
  6124=>"111000010",
  6125=>"110001110",
  6126=>"001111000",
  6127=>"100011101",
  6128=>"011010000",
  6129=>"100100100",
  6130=>"111101101",
  6131=>"101101111",
  6132=>"001011111",
  6133=>"111111010",
  6134=>"100000011",
  6135=>"000110100",
  6136=>"101111001",
  6137=>"010001011",
  6138=>"000011001",
  6139=>"000000100",
  6140=>"100101100",
  6141=>"010001100",
  6142=>"001111001",
  6143=>"101100010",
  6144=>"001110111",
  6145=>"101011010",
  6146=>"011110100",
  6147=>"001110000",
  6148=>"101000001",
  6149=>"100010000",
  6150=>"010101100",
  6151=>"001001111",
  6152=>"000101000",
  6153=>"010000010",
  6154=>"001000101",
  6155=>"101101101",
  6156=>"110011001",
  6157=>"011110011",
  6158=>"111100000",
  6159=>"000100010",
  6160=>"000001100",
  6161=>"010001000",
  6162=>"000100000",
  6163=>"110000101",
  6164=>"001101110",
  6165=>"100101000",
  6166=>"111111111",
  6167=>"011111111",
  6168=>"000010111",
  6169=>"101010010",
  6170=>"111110110",
  6171=>"001111101",
  6172=>"001011101",
  6173=>"001000010",
  6174=>"111110001",
  6175=>"101101011",
  6176=>"101101110",
  6177=>"111100100",
  6178=>"100000011",
  6179=>"000110101",
  6180=>"101101101",
  6181=>"111100010",
  6182=>"100001000",
  6183=>"110000101",
  6184=>"011000001",
  6185=>"001111000",
  6186=>"100110001",
  6187=>"101100011",
  6188=>"011000110",
  6189=>"101111110",
  6190=>"001001010",
  6191=>"011000000",
  6192=>"100011000",
  6193=>"010111001",
  6194=>"000001110",
  6195=>"010111110",
  6196=>"000111100",
  6197=>"000010011",
  6198=>"010010100",
  6199=>"001100101",
  6200=>"100101100",
  6201=>"011000000",
  6202=>"101001000",
  6203=>"000000101",
  6204=>"000110101",
  6205=>"111011110",
  6206=>"010001010",
  6207=>"101100000",
  6208=>"110011111",
  6209=>"000110000",
  6210=>"001000001",
  6211=>"100111110",
  6212=>"110000010",
  6213=>"000101110",
  6214=>"010100100",
  6215=>"110101110",
  6216=>"000110110",
  6217=>"110110101",
  6218=>"011101100",
  6219=>"100101001",
  6220=>"000111111",
  6221=>"100111001",
  6222=>"100000001",
  6223=>"000110001",
  6224=>"000101110",
  6225=>"111111101",
  6226=>"111110111",
  6227=>"110110110",
  6228=>"111001111",
  6229=>"101110000",
  6230=>"100010110",
  6231=>"101100100",
  6232=>"011001110",
  6233=>"011001011",
  6234=>"100001101",
  6235=>"101111011",
  6236=>"101000111",
  6237=>"101000000",
  6238=>"011011101",
  6239=>"111111111",
  6240=>"010110001",
  6241=>"110100101",
  6242=>"000010011",
  6243=>"000101000",
  6244=>"110000000",
  6245=>"111001101",
  6246=>"110100001",
  6247=>"100111000",
  6248=>"001111010",
  6249=>"000100010",
  6250=>"111101101",
  6251=>"110111111",
  6252=>"011101110",
  6253=>"011100111",
  6254=>"100111111",
  6255=>"110110100",
  6256=>"000001010",
  6257=>"111100100",
  6258=>"111001101",
  6259=>"100100010",
  6260=>"110001000",
  6261=>"100100010",
  6262=>"001110110",
  6263=>"010011011",
  6264=>"011001000",
  6265=>"101001000",
  6266=>"000000010",
  6267=>"001100101",
  6268=>"011000011",
  6269=>"010111101",
  6270=>"011001101",
  6271=>"100010111",
  6272=>"001000100",
  6273=>"011001100",
  6274=>"101111110",
  6275=>"011100001",
  6276=>"101011101",
  6277=>"000101000",
  6278=>"110010010",
  6279=>"001001001",
  6280=>"111101000",
  6281=>"100010100",
  6282=>"000110010",
  6283=>"010110011",
  6284=>"011000100",
  6285=>"000000000",
  6286=>"100000101",
  6287=>"111110011",
  6288=>"110010001",
  6289=>"100000011",
  6290=>"000001110",
  6291=>"100101001",
  6292=>"001000001",
  6293=>"100111110",
  6294=>"000001101",
  6295=>"001010111",
  6296=>"001000111",
  6297=>"001000111",
  6298=>"001110011",
  6299=>"011001100",
  6300=>"011111000",
  6301=>"101101110",
  6302=>"100010010",
  6303=>"010011111",
  6304=>"110100110",
  6305=>"000000011",
  6306=>"111100000",
  6307=>"101110100",
  6308=>"100000011",
  6309=>"000010010",
  6310=>"010011000",
  6311=>"001001110",
  6312=>"011101011",
  6313=>"010100011",
  6314=>"101011001",
  6315=>"110011110",
  6316=>"110011010",
  6317=>"100000111",
  6318=>"011100110",
  6319=>"100011001",
  6320=>"000111100",
  6321=>"101000011",
  6322=>"011111111",
  6323=>"111100110",
  6324=>"000110001",
  6325=>"101011110",
  6326=>"001011101",
  6327=>"010000100",
  6328=>"010100111",
  6329=>"010100000",
  6330=>"100100101",
  6331=>"001000101",
  6332=>"011000101",
  6333=>"101100010",
  6334=>"110010101",
  6335=>"011011000",
  6336=>"010111110",
  6337=>"111101101",
  6338=>"101111110",
  6339=>"011000101",
  6340=>"111110101",
  6341=>"101011000",
  6342=>"110000100",
  6343=>"001101000",
  6344=>"100010111",
  6345=>"100011101",
  6346=>"010011111",
  6347=>"001111101",
  6348=>"111111011",
  6349=>"111101001",
  6350=>"010000010",
  6351=>"010110110",
  6352=>"111001101",
  6353=>"101000001",
  6354=>"111010110",
  6355=>"111100001",
  6356=>"000101011",
  6357=>"000111101",
  6358=>"111100101",
  6359=>"010101010",
  6360=>"100110110",
  6361=>"000001100",
  6362=>"011111011",
  6363=>"011111100",
  6364=>"011111111",
  6365=>"111001111",
  6366=>"001101000",
  6367=>"110100010",
  6368=>"001101101",
  6369=>"111111111",
  6370=>"011111001",
  6371=>"111110010",
  6372=>"000010100",
  6373=>"011101110",
  6374=>"000011101",
  6375=>"000000111",
  6376=>"000000010",
  6377=>"110111000",
  6378=>"000101110",
  6379=>"011010000",
  6380=>"100111011",
  6381=>"101111010",
  6382=>"111101100",
  6383=>"111011011",
  6384=>"111000000",
  6385=>"001110010",
  6386=>"011111010",
  6387=>"001000111",
  6388=>"000000110",
  6389=>"000001010",
  6390=>"101001100",
  6391=>"000000000",
  6392=>"000101111",
  6393=>"101001000",
  6394=>"100101001",
  6395=>"011111000",
  6396=>"111101101",
  6397=>"110100000",
  6398=>"001111110",
  6399=>"111110100",
  6400=>"001010111",
  6401=>"101010011",
  6402=>"000000010",
  6403=>"000110100",
  6404=>"011100110",
  6405=>"101110011",
  6406=>"000000000",
  6407=>"110010011",
  6408=>"000001000",
  6409=>"010000100",
  6410=>"000000000",
  6411=>"001000110",
  6412=>"001011010",
  6413=>"100101011",
  6414=>"010001000",
  6415=>"111010111",
  6416=>"101001111",
  6417=>"001000010",
  6418=>"111000101",
  6419=>"001100100",
  6420=>"110110011",
  6421=>"000100000",
  6422=>"001100100",
  6423=>"110000010",
  6424=>"111000100",
  6425=>"001111101",
  6426=>"101101001",
  6427=>"000100110",
  6428=>"110111000",
  6429=>"011010100",
  6430=>"110001111",
  6431=>"100011100",
  6432=>"011101100",
  6433=>"101110001",
  6434=>"110111100",
  6435=>"010100010",
  6436=>"110000101",
  6437=>"011101001",
  6438=>"111101010",
  6439=>"000010111",
  6440=>"110101100",
  6441=>"111101010",
  6442=>"011001001",
  6443=>"101101001",
  6444=>"111010000",
  6445=>"101001101",
  6446=>"111001001",
  6447=>"111111011",
  6448=>"101100111",
  6449=>"100010110",
  6450=>"010010101",
  6451=>"111000011",
  6452=>"011000011",
  6453=>"111110010",
  6454=>"010011001",
  6455=>"101101110",
  6456=>"000001101",
  6457=>"011011010",
  6458=>"011101101",
  6459=>"011001001",
  6460=>"101101011",
  6461=>"000101011",
  6462=>"001100110",
  6463=>"111111000",
  6464=>"100011110",
  6465=>"001101101",
  6466=>"001110001",
  6467=>"111000010",
  6468=>"100100010",
  6469=>"110111001",
  6470=>"011011011",
  6471=>"111111101",
  6472=>"001000111",
  6473=>"000001001",
  6474=>"110100010",
  6475=>"101101100",
  6476=>"010010011",
  6477=>"110111100",
  6478=>"111101010",
  6479=>"001010010",
  6480=>"111001100",
  6481=>"111110011",
  6482=>"011010001",
  6483=>"001100111",
  6484=>"010101111",
  6485=>"101101011",
  6486=>"011100000",
  6487=>"111101110",
  6488=>"110100111",
  6489=>"110110011",
  6490=>"110011100",
  6491=>"110111101",
  6492=>"001111010",
  6493=>"010001011",
  6494=>"011101110",
  6495=>"010000100",
  6496=>"101111100",
  6497=>"000010101",
  6498=>"101101101",
  6499=>"011110010",
  6500=>"100001000",
  6501=>"111101010",
  6502=>"011100101",
  6503=>"100001001",
  6504=>"011110100",
  6505=>"110111011",
  6506=>"111001000",
  6507=>"111010110",
  6508=>"101010010",
  6509=>"111111011",
  6510=>"101010100",
  6511=>"000000101",
  6512=>"110100101",
  6513=>"001100000",
  6514=>"001101101",
  6515=>"100111010",
  6516=>"111110100",
  6517=>"100000010",
  6518=>"011000101",
  6519=>"101100110",
  6520=>"101001100",
  6521=>"110001000",
  6522=>"010001101",
  6523=>"011110010",
  6524=>"001001011",
  6525=>"111101001",
  6526=>"111111100",
  6527=>"111010111",
  6528=>"101100110",
  6529=>"001000010",
  6530=>"111100111",
  6531=>"011111011",
  6532=>"001110100",
  6533=>"000001101",
  6534=>"110101001",
  6535=>"101110010",
  6536=>"010111100",
  6537=>"110001110",
  6538=>"110111001",
  6539=>"010000001",
  6540=>"001100111",
  6541=>"001101010",
  6542=>"001101000",
  6543=>"010000111",
  6544=>"101011000",
  6545=>"011010000",
  6546=>"111110110",
  6547=>"011101010",
  6548=>"001100101",
  6549=>"001100011",
  6550=>"111111011",
  6551=>"001111001",
  6552=>"000101101",
  6553=>"011110110",
  6554=>"001101110",
  6555=>"001111100",
  6556=>"011100110",
  6557=>"111111110",
  6558=>"101010101",
  6559=>"011011000",
  6560=>"111110010",
  6561=>"001100110",
  6562=>"101010000",
  6563=>"100000001",
  6564=>"000101110",
  6565=>"111011101",
  6566=>"001110110",
  6567=>"110101011",
  6568=>"001000100",
  6569=>"100100000",
  6570=>"111100000",
  6571=>"100100111",
  6572=>"100100110",
  6573=>"100100011",
  6574=>"101010000",
  6575=>"101010101",
  6576=>"000000001",
  6577=>"011001000",
  6578=>"000111000",
  6579=>"111001001",
  6580=>"111000110",
  6581=>"111111001",
  6582=>"011001100",
  6583=>"111101111",
  6584=>"011010111",
  6585=>"111011011",
  6586=>"010011110",
  6587=>"111010100",
  6588=>"100110010",
  6589=>"000001001",
  6590=>"001000011",
  6591=>"101101111",
  6592=>"111101101",
  6593=>"010000001",
  6594=>"011011001",
  6595=>"101111000",
  6596=>"111101111",
  6597=>"001110010",
  6598=>"011011101",
  6599=>"011011101",
  6600=>"000111100",
  6601=>"100001001",
  6602=>"100001010",
  6603=>"011100011",
  6604=>"100001111",
  6605=>"000000001",
  6606=>"011110110",
  6607=>"111110100",
  6608=>"011000001",
  6609=>"010101011",
  6610=>"111111100",
  6611=>"100001001",
  6612=>"110111111",
  6613=>"011101000",
  6614=>"110100011",
  6615=>"010001010",
  6616=>"100011010",
  6617=>"110100101",
  6618=>"000011000",
  6619=>"011000001",
  6620=>"110100010",
  6621=>"011101100",
  6622=>"101100100",
  6623=>"111100111",
  6624=>"101101011",
  6625=>"111011010",
  6626=>"110001001",
  6627=>"001001100",
  6628=>"010111111",
  6629=>"000011011",
  6630=>"110100110",
  6631=>"001001010",
  6632=>"010111110",
  6633=>"000110110",
  6634=>"101000010",
  6635=>"010111011",
  6636=>"110100100",
  6637=>"100000000",
  6638=>"010011101",
  6639=>"000011111",
  6640=>"010111100",
  6641=>"101111100",
  6642=>"110101111",
  6643=>"101101010",
  6644=>"111111101",
  6645=>"111010101",
  6646=>"110111010",
  6647=>"000011000",
  6648=>"011111010",
  6649=>"100010100",
  6650=>"111101111",
  6651=>"010011111",
  6652=>"010100110",
  6653=>"001111001",
  6654=>"000000100",
  6655=>"101001001",
  6656=>"010101011",
  6657=>"000111010",
  6658=>"000110011",
  6659=>"101001101",
  6660=>"101101100",
  6661=>"101110100",
  6662=>"000100111",
  6663=>"010001110",
  6664=>"111101101",
  6665=>"101100000",
  6666=>"011101010",
  6667=>"001101010",
  6668=>"011100101",
  6669=>"100000001",
  6670=>"100101101",
  6671=>"001000001",
  6672=>"001100101",
  6673=>"001101111",
  6674=>"000000011",
  6675=>"001000001",
  6676=>"000001011",
  6677=>"010001110",
  6678=>"000100110",
  6679=>"001111000",
  6680=>"100111000",
  6681=>"110010011",
  6682=>"111101001",
  6683=>"001110101",
  6684=>"111001001",
  6685=>"111110010",
  6686=>"000101111",
  6687=>"110101101",
  6688=>"010010110",
  6689=>"010110010",
  6690=>"000001001",
  6691=>"010101101",
  6692=>"110100010",
  6693=>"001111000",
  6694=>"110010110",
  6695=>"100100110",
  6696=>"100100100",
  6697=>"001000110",
  6698=>"111010010",
  6699=>"111010100",
  6700=>"001110010",
  6701=>"011100111",
  6702=>"111110110",
  6703=>"111111000",
  6704=>"000111100",
  6705=>"001011111",
  6706=>"010111000",
  6707=>"111011110",
  6708=>"001101101",
  6709=>"101010001",
  6710=>"100101001",
  6711=>"010000011",
  6712=>"101101000",
  6713=>"010001001",
  6714=>"011110001",
  6715=>"110001000",
  6716=>"100000111",
  6717=>"110111111",
  6718=>"010101110",
  6719=>"110110010",
  6720=>"010011111",
  6721=>"010100111",
  6722=>"000101110",
  6723=>"100111110",
  6724=>"101101101",
  6725=>"010001110",
  6726=>"010100101",
  6727=>"110101001",
  6728=>"111111101",
  6729=>"111101100",
  6730=>"100101100",
  6731=>"111000110",
  6732=>"000010011",
  6733=>"101101010",
  6734=>"000011101",
  6735=>"010001101",
  6736=>"010111000",
  6737=>"000000000",
  6738=>"000010101",
  6739=>"001000100",
  6740=>"100110011",
  6741=>"110011011",
  6742=>"111101110",
  6743=>"010001000",
  6744=>"000111000",
  6745=>"010100000",
  6746=>"000011000",
  6747=>"101001101",
  6748=>"111110000",
  6749=>"111101100",
  6750=>"110100010",
  6751=>"001110100",
  6752=>"111001111",
  6753=>"011011010",
  6754=>"101000001",
  6755=>"100010100",
  6756=>"000011101",
  6757=>"000000011",
  6758=>"010010110",
  6759=>"011111110",
  6760=>"010101111",
  6761=>"011101010",
  6762=>"010111001",
  6763=>"111110100",
  6764=>"010010011",
  6765=>"110101011",
  6766=>"111001100",
  6767=>"001111101",
  6768=>"100010110",
  6769=>"110111110",
  6770=>"010110001",
  6771=>"100010100",
  6772=>"010110111",
  6773=>"101000011",
  6774=>"110110100",
  6775=>"000110001",
  6776=>"101110011",
  6777=>"100000011",
  6778=>"010000101",
  6779=>"000010100",
  6780=>"010101101",
  6781=>"111101111",
  6782=>"111100101",
  6783=>"000001111",
  6784=>"010000001",
  6785=>"101011001",
  6786=>"011011001",
  6787=>"110100011",
  6788=>"001100101",
  6789=>"111110010",
  6790=>"100101010",
  6791=>"111000000",
  6792=>"011010100",
  6793=>"000011001",
  6794=>"011010011",
  6795=>"001111010",
  6796=>"110111011",
  6797=>"111101111",
  6798=>"011001110",
  6799=>"001110111",
  6800=>"010110110",
  6801=>"010100100",
  6802=>"010110000",
  6803=>"001101110",
  6804=>"000110110",
  6805=>"001110100",
  6806=>"011011111",
  6807=>"111110110",
  6808=>"000010010",
  6809=>"110111110",
  6810=>"011000001",
  6811=>"101000010",
  6812=>"101111001",
  6813=>"000110101",
  6814=>"010010011",
  6815=>"010010010",
  6816=>"011101001",
  6817=>"010001000",
  6818=>"101011000",
  6819=>"000011100",
  6820=>"100110100",
  6821=>"100100100",
  6822=>"110011000",
  6823=>"000000011",
  6824=>"001100110",
  6825=>"010000110",
  6826=>"110000001",
  6827=>"110001100",
  6828=>"001011101",
  6829=>"110101001",
  6830=>"101011101",
  6831=>"110101100",
  6832=>"000000100",
  6833=>"100011101",
  6834=>"011111001",
  6835=>"111011111",
  6836=>"001100110",
  6837=>"100100000",
  6838=>"001100001",
  6839=>"011000011",
  6840=>"011000100",
  6841=>"111111001",
  6842=>"010001101",
  6843=>"010110111",
  6844=>"101101010",
  6845=>"011001001",
  6846=>"111101001",
  6847=>"000101100",
  6848=>"011101111",
  6849=>"011011001",
  6850=>"000011111",
  6851=>"101101111",
  6852=>"001110110",
  6853=>"101000011",
  6854=>"011101111",
  6855=>"001010111",
  6856=>"001000000",
  6857=>"011010101",
  6858=>"101010001",
  6859=>"000000110",
  6860=>"110101111",
  6861=>"000010100",
  6862=>"000111011",
  6863=>"000100100",
  6864=>"011001011",
  6865=>"001111000",
  6866=>"100010000",
  6867=>"010111010",
  6868=>"001000111",
  6869=>"000011000",
  6870=>"001011000",
  6871=>"010101001",
  6872=>"111111010",
  6873=>"011100100",
  6874=>"010000010",
  6875=>"100010000",
  6876=>"111111011",
  6877=>"100100000",
  6878=>"100100010",
  6879=>"100110100",
  6880=>"011010110",
  6881=>"001011110",
  6882=>"001110100",
  6883=>"011000111",
  6884=>"101101011",
  6885=>"010111010",
  6886=>"011011111",
  6887=>"000001100",
  6888=>"110011101",
  6889=>"111010101",
  6890=>"000001100",
  6891=>"001000000",
  6892=>"111101001",
  6893=>"000100101",
  6894=>"011110000",
  6895=>"101101010",
  6896=>"111111010",
  6897=>"000010010",
  6898=>"010100000",
  6899=>"000001111",
  6900=>"000110011",
  6901=>"011000001",
  6902=>"101010010",
  6903=>"010000111",
  6904=>"110110111",
  6905=>"111100110",
  6906=>"110001001",
  6907=>"000010110",
  6908=>"000101110",
  6909=>"110001110",
  6910=>"010011100",
  6911=>"100110010",
  6912=>"101011011",
  6913=>"010011111",
  6914=>"111101100",
  6915=>"001101111",
  6916=>"111001111",
  6917=>"011000110",
  6918=>"110010100",
  6919=>"101001111",
  6920=>"000010110",
  6921=>"010111001",
  6922=>"111010110",
  6923=>"101010111",
  6924=>"001101111",
  6925=>"101010010",
  6926=>"011001011",
  6927=>"011011001",
  6928=>"001110101",
  6929=>"001010010",
  6930=>"001100000",
  6931=>"010011001",
  6932=>"011111000",
  6933=>"110010101",
  6934=>"001100000",
  6935=>"100110110",
  6936=>"001111010",
  6937=>"010101110",
  6938=>"001000011",
  6939=>"000100010",
  6940=>"000010111",
  6941=>"100111101",
  6942=>"101110001",
  6943=>"110010101",
  6944=>"110001101",
  6945=>"111100011",
  6946=>"010111111",
  6947=>"101100011",
  6948=>"110101010",
  6949=>"111001000",
  6950=>"010101001",
  6951=>"000000011",
  6952=>"100111100",
  6953=>"111000111",
  6954=>"111100110",
  6955=>"010111011",
  6956=>"001001111",
  6957=>"011111110",
  6958=>"101010110",
  6959=>"011111110",
  6960=>"111011001",
  6961=>"110110111",
  6962=>"100011011",
  6963=>"110111000",
  6964=>"100000001",
  6965=>"110101011",
  6966=>"011110100",
  6967=>"111100010",
  6968=>"101110000",
  6969=>"110110110",
  6970=>"111000100",
  6971=>"110110000",
  6972=>"001001001",
  6973=>"000101001",
  6974=>"011111100",
  6975=>"011000011",
  6976=>"111000000",
  6977=>"011101110",
  6978=>"111111100",
  6979=>"101001100",
  6980=>"100001100",
  6981=>"011110100",
  6982=>"100111001",
  6983=>"001011101",
  6984=>"011001000",
  6985=>"100110000",
  6986=>"110110010",
  6987=>"100110101",
  6988=>"010000001",
  6989=>"011011110",
  6990=>"110010000",
  6991=>"101010001",
  6992=>"110110001",
  6993=>"011010011",
  6994=>"100000101",
  6995=>"010110000",
  6996=>"110110101",
  6997=>"111100000",
  6998=>"111111011",
  6999=>"111000110",
  7000=>"100101101",
  7001=>"001001010",
  7002=>"000100010",
  7003=>"111111011",
  7004=>"001010000",
  7005=>"111111111",
  7006=>"001010011",
  7007=>"111101111",
  7008=>"011110011",
  7009=>"000010100",
  7010=>"000000101",
  7011=>"111101110",
  7012=>"010000110",
  7013=>"000111000",
  7014=>"011000101",
  7015=>"010101110",
  7016=>"000010101",
  7017=>"011101000",
  7018=>"110001010",
  7019=>"010010101",
  7020=>"100110100",
  7021=>"111000111",
  7022=>"100100110",
  7023=>"100100000",
  7024=>"011110101",
  7025=>"011111110",
  7026=>"101100010",
  7027=>"011010101",
  7028=>"000001001",
  7029=>"110001101",
  7030=>"101010100",
  7031=>"001011011",
  7032=>"010010010",
  7033=>"101000001",
  7034=>"001000101",
  7035=>"000010011",
  7036=>"010111110",
  7037=>"111111101",
  7038=>"111100000",
  7039=>"010111011",
  7040=>"000011100",
  7041=>"001001101",
  7042=>"100000000",
  7043=>"100110100",
  7044=>"001110011",
  7045=>"010111110",
  7046=>"010011101",
  7047=>"001001101",
  7048=>"000010001",
  7049=>"101111001",
  7050=>"001100111",
  7051=>"101000010",
  7052=>"111111000",
  7053=>"111011001",
  7054=>"010100111",
  7055=>"001111100",
  7056=>"101100101",
  7057=>"000111010",
  7058=>"111001101",
  7059=>"011110110",
  7060=>"100001000",
  7061=>"000111000",
  7062=>"010100101",
  7063=>"110111000",
  7064=>"010011000",
  7065=>"010000011",
  7066=>"000000111",
  7067=>"101000110",
  7068=>"001101101",
  7069=>"011100010",
  7070=>"010010001",
  7071=>"100010011",
  7072=>"110110110",
  7073=>"010111111",
  7074=>"010110011",
  7075=>"011010010",
  7076=>"001101000",
  7077=>"010001001",
  7078=>"100010110",
  7079=>"001000000",
  7080=>"000000110",
  7081=>"101011101",
  7082=>"100001110",
  7083=>"001001100",
  7084=>"111001000",
  7085=>"010110011",
  7086=>"110100011",
  7087=>"000011111",
  7088=>"000110011",
  7089=>"011000101",
  7090=>"011011011",
  7091=>"100111101",
  7092=>"100111000",
  7093=>"011100101",
  7094=>"010110000",
  7095=>"000111010",
  7096=>"100000100",
  7097=>"100000111",
  7098=>"001010111",
  7099=>"110010101",
  7100=>"111111000",
  7101=>"010101100",
  7102=>"110111010",
  7103=>"111111111",
  7104=>"000000001",
  7105=>"111010001",
  7106=>"100010101",
  7107=>"101000000",
  7108=>"101000001",
  7109=>"001000110",
  7110=>"110011011",
  7111=>"001101111",
  7112=>"010001100",
  7113=>"000011110",
  7114=>"101101011",
  7115=>"110101100",
  7116=>"101101111",
  7117=>"111111000",
  7118=>"111001001",
  7119=>"000110100",
  7120=>"100011101",
  7121=>"100101100",
  7122=>"111000100",
  7123=>"110011011",
  7124=>"010101101",
  7125=>"111110100",
  7126=>"010010101",
  7127=>"111011000",
  7128=>"111100111",
  7129=>"010011100",
  7130=>"011111111",
  7131=>"110010100",
  7132=>"001000010",
  7133=>"100000001",
  7134=>"000010011",
  7135=>"100110010",
  7136=>"110111101",
  7137=>"010111000",
  7138=>"010001110",
  7139=>"000110100",
  7140=>"111110110",
  7141=>"111010011",
  7142=>"011010101",
  7143=>"100011100",
  7144=>"000011100",
  7145=>"110110111",
  7146=>"111101111",
  7147=>"100000010",
  7148=>"010111010",
  7149=>"001010001",
  7150=>"000100101",
  7151=>"010011110",
  7152=>"011000000",
  7153=>"100001110",
  7154=>"011010000",
  7155=>"101010101",
  7156=>"001010100",
  7157=>"100110001",
  7158=>"011010110",
  7159=>"111011100",
  7160=>"111011000",
  7161=>"111111100",
  7162=>"101000110",
  7163=>"001101011",
  7164=>"000010000",
  7165=>"110100011",
  7166=>"111111000",
  7167=>"010010001",
  7168=>"001110101",
  7169=>"011001111",
  7170=>"001100100",
  7171=>"100110111",
  7172=>"010111011",
  7173=>"000110111",
  7174=>"010011001",
  7175=>"110111111",
  7176=>"011100000",
  7177=>"111110100",
  7178=>"000000111",
  7179=>"111010011",
  7180=>"010100010",
  7181=>"000100001",
  7182=>"110001111",
  7183=>"010000011",
  7184=>"000111010",
  7185=>"110010011",
  7186=>"001011100",
  7187=>"101010111",
  7188=>"010111010",
  7189=>"011010100",
  7190=>"010100111",
  7191=>"000000011",
  7192=>"111101111",
  7193=>"011001010",
  7194=>"101010111",
  7195=>"100110011",
  7196=>"010011100",
  7197=>"101100101",
  7198=>"001011100",
  7199=>"000110011",
  7200=>"010011001",
  7201=>"010010110",
  7202=>"101010100",
  7203=>"100100111",
  7204=>"011001011",
  7205=>"101110000",
  7206=>"111001110",
  7207=>"111100100",
  7208=>"001010011",
  7209=>"011110001",
  7210=>"011111001",
  7211=>"101101011",
  7212=>"000010100",
  7213=>"010010001",
  7214=>"100010101",
  7215=>"100111011",
  7216=>"011001111",
  7217=>"111110000",
  7218=>"001010000",
  7219=>"011111111",
  7220=>"101001000",
  7221=>"000110100",
  7222=>"111100110",
  7223=>"010011111",
  7224=>"000110010",
  7225=>"100000000",
  7226=>"001011010",
  7227=>"010111110",
  7228=>"011100000",
  7229=>"010000001",
  7230=>"001000010",
  7231=>"111110111",
  7232=>"110011100",
  7233=>"000001011",
  7234=>"001000111",
  7235=>"101100110",
  7236=>"101110001",
  7237=>"011010100",
  7238=>"111110000",
  7239=>"100010111",
  7240=>"100100001",
  7241=>"010011011",
  7242=>"010100100",
  7243=>"101110000",
  7244=>"011000001",
  7245=>"010111011",
  7246=>"001001111",
  7247=>"101000100",
  7248=>"101110011",
  7249=>"110101011",
  7250=>"001101000",
  7251=>"110100101",
  7252=>"100100010",
  7253=>"011110110",
  7254=>"100110111",
  7255=>"101100001",
  7256=>"001101000",
  7257=>"000111000",
  7258=>"000101110",
  7259=>"100001010",
  7260=>"111001010",
  7261=>"100000000",
  7262=>"010110001",
  7263=>"000010010",
  7264=>"000101101",
  7265=>"010110111",
  7266=>"111100111",
  7267=>"000001011",
  7268=>"010010001",
  7269=>"100100111",
  7270=>"010011001",
  7271=>"101111000",
  7272=>"011000100",
  7273=>"000111100",
  7274=>"000001001",
  7275=>"100010001",
  7276=>"101110100",
  7277=>"110110011",
  7278=>"011010000",
  7279=>"001010111",
  7280=>"100110011",
  7281=>"001011011",
  7282=>"011100000",
  7283=>"101110110",
  7284=>"111000001",
  7285=>"000100000",
  7286=>"111100001",
  7287=>"111110111",
  7288=>"010110010",
  7289=>"001011110",
  7290=>"100100101",
  7291=>"000100000",
  7292=>"011000101",
  7293=>"001000111",
  7294=>"000001100",
  7295=>"011110010",
  7296=>"011011001",
  7297=>"101111110",
  7298=>"010011111",
  7299=>"000101001",
  7300=>"010001000",
  7301=>"111100001",
  7302=>"101101111",
  7303=>"000100010",
  7304=>"011111000",
  7305=>"101101010",
  7306=>"101110001",
  7307=>"010000101",
  7308=>"111101110",
  7309=>"100101100",
  7310=>"110011101",
  7311=>"001110010",
  7312=>"000000111",
  7313=>"111010101",
  7314=>"000000101",
  7315=>"111011001",
  7316=>"101001011",
  7317=>"011001110",
  7318=>"110111011",
  7319=>"101110000",
  7320=>"101011111",
  7321=>"000111110",
  7322=>"111001010",
  7323=>"001001000",
  7324=>"110100110",
  7325=>"011000011",
  7326=>"111001011",
  7327=>"010101110",
  7328=>"110111100",
  7329=>"001101111",
  7330=>"000000111",
  7331=>"001111111",
  7332=>"111111111",
  7333=>"101101011",
  7334=>"010011110",
  7335=>"000010101",
  7336=>"000001000",
  7337=>"100111011",
  7338=>"110000100",
  7339=>"010101010",
  7340=>"010001000",
  7341=>"000000110",
  7342=>"010010111",
  7343=>"000100001",
  7344=>"111010101",
  7345=>"100000111",
  7346=>"110010110",
  7347=>"110010011",
  7348=>"110010110",
  7349=>"100101111",
  7350=>"000010001",
  7351=>"001011100",
  7352=>"111000000",
  7353=>"000000111",
  7354=>"100010100",
  7355=>"010100010",
  7356=>"001111110",
  7357=>"101010000",
  7358=>"000010100",
  7359=>"001010011",
  7360=>"000011101",
  7361=>"000000101",
  7362=>"111000010",
  7363=>"011101101",
  7364=>"000000000",
  7365=>"100111000",
  7366=>"001101001",
  7367=>"010000000",
  7368=>"101001011",
  7369=>"101011100",
  7370=>"101100110",
  7371=>"101011101",
  7372=>"010110011",
  7373=>"011100011",
  7374=>"000001111",
  7375=>"101011010",
  7376=>"101110101",
  7377=>"100111000",
  7378=>"100000010",
  7379=>"101111100",
  7380=>"110011000",
  7381=>"011011000",
  7382=>"110000100",
  7383=>"110100010",
  7384=>"100010111",
  7385=>"101010010",
  7386=>"000101000",
  7387=>"001100111",
  7388=>"001101001",
  7389=>"111100101",
  7390=>"001010000",
  7391=>"101000010",
  7392=>"001100001",
  7393=>"101000101",
  7394=>"010100010",
  7395=>"010101011",
  7396=>"101010011",
  7397=>"111011001",
  7398=>"000010010",
  7399=>"010101011",
  7400=>"110010000",
  7401=>"110001001",
  7402=>"000101000",
  7403=>"111010110",
  7404=>"110101000",
  7405=>"100011110",
  7406=>"110111000",
  7407=>"111011000",
  7408=>"011010101",
  7409=>"110111100",
  7410=>"010101100",
  7411=>"010101111",
  7412=>"101001110",
  7413=>"001000001",
  7414=>"010111110",
  7415=>"101000010",
  7416=>"110010111",
  7417=>"001101000",
  7418=>"110100100",
  7419=>"000111011",
  7420=>"010001010",
  7421=>"110111110",
  7422=>"001100101",
  7423=>"101100010",
  7424=>"110100010",
  7425=>"110001111",
  7426=>"000111010",
  7427=>"111111111",
  7428=>"010110110",
  7429=>"010111011",
  7430=>"100100011",
  7431=>"100000110",
  7432=>"000011101",
  7433=>"011101100",
  7434=>"111110001",
  7435=>"111110101",
  7436=>"100001010",
  7437=>"010010000",
  7438=>"010101011",
  7439=>"011001011",
  7440=>"011100010",
  7441=>"011010001",
  7442=>"011100100",
  7443=>"110000110",
  7444=>"011111011",
  7445=>"101001111",
  7446=>"010100100",
  7447=>"100111010",
  7448=>"100011000",
  7449=>"100001110",
  7450=>"100010011",
  7451=>"011001111",
  7452=>"000010011",
  7453=>"111110111",
  7454=>"110111000",
  7455=>"000110110",
  7456=>"000110000",
  7457=>"000001000",
  7458=>"100010000",
  7459=>"101110100",
  7460=>"110101100",
  7461=>"010010100",
  7462=>"001010010",
  7463=>"001010010",
  7464=>"000100110",
  7465=>"111101000",
  7466=>"101110110",
  7467=>"101111101",
  7468=>"101011101",
  7469=>"010000101",
  7470=>"111000001",
  7471=>"111111111",
  7472=>"000110101",
  7473=>"111111000",
  7474=>"011000110",
  7475=>"100000110",
  7476=>"100000011",
  7477=>"100000111",
  7478=>"010000010",
  7479=>"001000110",
  7480=>"101001100",
  7481=>"010101000",
  7482=>"010110001",
  7483=>"111111101",
  7484=>"101011001",
  7485=>"010100001",
  7486=>"000101010",
  7487=>"101010111",
  7488=>"101101011",
  7489=>"111010000",
  7490=>"000011001",
  7491=>"010100110",
  7492=>"000001010",
  7493=>"100101011",
  7494=>"111001000",
  7495=>"111001100",
  7496=>"100110010",
  7497=>"101111001",
  7498=>"101100100",
  7499=>"101100100",
  7500=>"010000000",
  7501=>"000001100",
  7502=>"010101100",
  7503=>"111000001",
  7504=>"011111001",
  7505=>"101001111",
  7506=>"011001110",
  7507=>"110000001",
  7508=>"000000001",
  7509=>"111110111",
  7510=>"110001010",
  7511=>"000000111",
  7512=>"111010111",
  7513=>"001100111",
  7514=>"111001000",
  7515=>"111000010",
  7516=>"010011101",
  7517=>"001101101",
  7518=>"011100011",
  7519=>"010111000",
  7520=>"101001001",
  7521=>"010101111",
  7522=>"010110100",
  7523=>"000111010",
  7524=>"000110000",
  7525=>"010100011",
  7526=>"011101001",
  7527=>"011011110",
  7528=>"111001101",
  7529=>"101010010",
  7530=>"000110111",
  7531=>"101101111",
  7532=>"000101110",
  7533=>"100100000",
  7534=>"010000100",
  7535=>"010010001",
  7536=>"111011011",
  7537=>"111001101",
  7538=>"101000011",
  7539=>"110000001",
  7540=>"110010010",
  7541=>"101101110",
  7542=>"001010001",
  7543=>"000000000",
  7544=>"000011010",
  7545=>"101101101",
  7546=>"011101001",
  7547=>"000110011",
  7548=>"110011111",
  7549=>"100101101",
  7550=>"100110100",
  7551=>"101101100",
  7552=>"101001111",
  7553=>"011000011",
  7554=>"110011011",
  7555=>"111110100",
  7556=>"011010001",
  7557=>"000000010",
  7558=>"011000100",
  7559=>"100011111",
  7560=>"010010001",
  7561=>"000101010",
  7562=>"110111010",
  7563=>"111011010",
  7564=>"100111100",
  7565=>"111110101",
  7566=>"010000001",
  7567=>"101011000",
  7568=>"001010101",
  7569=>"000101001",
  7570=>"101100100",
  7571=>"111101100",
  7572=>"100001100",
  7573=>"000001001",
  7574=>"010100000",
  7575=>"010000000",
  7576=>"111110101",
  7577=>"100010011",
  7578=>"101111000",
  7579=>"100111011",
  7580=>"101110100",
  7581=>"000100101",
  7582=>"101010001",
  7583=>"100101100",
  7584=>"101000000",
  7585=>"110111110",
  7586=>"100010100",
  7587=>"111111011",
  7588=>"110110000",
  7589=>"000010000",
  7590=>"001110111",
  7591=>"101011100",
  7592=>"011011101",
  7593=>"100011000",
  7594=>"100110011",
  7595=>"100000110",
  7596=>"100101100",
  7597=>"011110011",
  7598=>"000011100",
  7599=>"011010010",
  7600=>"001101101",
  7601=>"100001110",
  7602=>"100100101",
  7603=>"011111111",
  7604=>"001001110",
  7605=>"011100000",
  7606=>"101101101",
  7607=>"010111100",
  7608=>"001110111",
  7609=>"001000110",
  7610=>"000000000",
  7611=>"010001011",
  7612=>"111010011",
  7613=>"011001010",
  7614=>"001001010",
  7615=>"110011001",
  7616=>"111110100",
  7617=>"100000010",
  7618=>"100011010",
  7619=>"101001100",
  7620=>"101001010",
  7621=>"110010011",
  7622=>"011111010",
  7623=>"100000001",
  7624=>"101110111",
  7625=>"110101011",
  7626=>"110011110",
  7627=>"011001110",
  7628=>"000011001",
  7629=>"010000010",
  7630=>"100001111",
  7631=>"100010010",
  7632=>"001101000",
  7633=>"100101100",
  7634=>"100000100",
  7635=>"100000001",
  7636=>"111110110",
  7637=>"001011101",
  7638=>"110011110",
  7639=>"101111110",
  7640=>"110000010",
  7641=>"000000111",
  7642=>"011111101",
  7643=>"101000000",
  7644=>"110001110",
  7645=>"101111001",
  7646=>"100111010",
  7647=>"101010100",
  7648=>"000100110",
  7649=>"110010001",
  7650=>"111111011",
  7651=>"001110000",
  7652=>"000010101",
  7653=>"000010001",
  7654=>"000011010",
  7655=>"001001001",
  7656=>"111101010",
  7657=>"111110011",
  7658=>"110101111",
  7659=>"101010010",
  7660=>"011000100",
  7661=>"000101000",
  7662=>"011111101",
  7663=>"010010000",
  7664=>"111011010",
  7665=>"010010011",
  7666=>"110111101",
  7667=>"101000100",
  7668=>"110110100",
  7669=>"000111110",
  7670=>"111010110",
  7671=>"001110010",
  7672=>"001000100",
  7673=>"100011111",
  7674=>"110011010",
  7675=>"101010100",
  7676=>"101011010",
  7677=>"001100100",
  7678=>"010100000",
  7679=>"000110000",
  7680=>"100001100",
  7681=>"001100001",
  7682=>"101110110",
  7683=>"100111011",
  7684=>"011000110",
  7685=>"010101010",
  7686=>"111000000",
  7687=>"000100000",
  7688=>"001101000",
  7689=>"010110010",
  7690=>"100001011",
  7691=>"001001101",
  7692=>"010110110",
  7693=>"001010110",
  7694=>"000000010",
  7695=>"101110100",
  7696=>"001000101",
  7697=>"001011110",
  7698=>"011001100",
  7699=>"111101101",
  7700=>"100100010",
  7701=>"111101100",
  7702=>"100010100",
  7703=>"111001011",
  7704=>"110110110",
  7705=>"110101100",
  7706=>"000001111",
  7707=>"101001101",
  7708=>"010111011",
  7709=>"111101100",
  7710=>"100111001",
  7711=>"101011110",
  7712=>"010010000",
  7713=>"001010001",
  7714=>"011110100",
  7715=>"111101110",
  7716=>"000001111",
  7717=>"100101100",
  7718=>"110100100",
  7719=>"000000110",
  7720=>"100000011",
  7721=>"001001100",
  7722=>"010111100",
  7723=>"001110000",
  7724=>"100111011",
  7725=>"011001101",
  7726=>"001101111",
  7727=>"000110101",
  7728=>"011111100",
  7729=>"010000000",
  7730=>"010010000",
  7731=>"101110101",
  7732=>"011111101",
  7733=>"110110110",
  7734=>"010000111",
  7735=>"101111000",
  7736=>"101111111",
  7737=>"010110011",
  7738=>"011000010",
  7739=>"101010111",
  7740=>"110000111",
  7741=>"011101011",
  7742=>"000000000",
  7743=>"000001110",
  7744=>"011010101",
  7745=>"011001010",
  7746=>"000001000",
  7747=>"111111000",
  7748=>"101110011",
  7749=>"100100000",
  7750=>"000000001",
  7751=>"110001100",
  7752=>"000001110",
  7753=>"011111011",
  7754=>"001000100",
  7755=>"000010110",
  7756=>"011000001",
  7757=>"001110000",
  7758=>"110100000",
  7759=>"110110000",
  7760=>"100001010",
  7761=>"001110110",
  7762=>"111100110",
  7763=>"110001110",
  7764=>"010100010",
  7765=>"001101111",
  7766=>"110100010",
  7767=>"110001010",
  7768=>"000111000",
  7769=>"111111011",
  7770=>"010110110",
  7771=>"111011010",
  7772=>"111011100",
  7773=>"110111110",
  7774=>"010111000",
  7775=>"000000000",
  7776=>"000111101",
  7777=>"100011011",
  7778=>"111110101",
  7779=>"010010010",
  7780=>"011100001",
  7781=>"001111111",
  7782=>"111100100",
  7783=>"110011011",
  7784=>"010011011",
  7785=>"110010100",
  7786=>"011000001",
  7787=>"011010000",
  7788=>"101111110",
  7789=>"000011100",
  7790=>"111110010",
  7791=>"110011000",
  7792=>"000001001",
  7793=>"000000000",
  7794=>"110110011",
  7795=>"110100010",
  7796=>"001111000",
  7797=>"110001011",
  7798=>"100010111",
  7799=>"010100001",
  7800=>"000010110",
  7801=>"000010110",
  7802=>"101001000",
  7803=>"000000110",
  7804=>"110100100",
  7805=>"000110111",
  7806=>"011011100",
  7807=>"110001000",
  7808=>"001000010",
  7809=>"101011001",
  7810=>"011010110",
  7811=>"110101010",
  7812=>"100010000",
  7813=>"111010111",
  7814=>"110000011",
  7815=>"110101111",
  7816=>"010100011",
  7817=>"001100001",
  7818=>"000101000",
  7819=>"101111101",
  7820=>"000110100",
  7821=>"001100100",
  7822=>"111001100",
  7823=>"000100000",
  7824=>"110011100",
  7825=>"001100001",
  7826=>"100100101",
  7827=>"000101100",
  7828=>"001000011",
  7829=>"011111000",
  7830=>"110111100",
  7831=>"100110101",
  7832=>"001111100",
  7833=>"111110001",
  7834=>"001010011",
  7835=>"101110001",
  7836=>"100111000",
  7837=>"111111011",
  7838=>"110100010",
  7839=>"110011010",
  7840=>"001100110",
  7841=>"110001010",
  7842=>"111101011",
  7843=>"000011011",
  7844=>"111110101",
  7845=>"100101100",
  7846=>"100010100",
  7847=>"001010000",
  7848=>"010111011",
  7849=>"001110100",
  7850=>"010000001",
  7851=>"001111010",
  7852=>"111111111",
  7853=>"101101001",
  7854=>"001110100",
  7855=>"011101011",
  7856=>"100001111",
  7857=>"001101111",
  7858=>"111010001",
  7859=>"101110110",
  7860=>"010100110",
  7861=>"010011010",
  7862=>"011011101",
  7863=>"111010000",
  7864=>"000100111",
  7865=>"111000101",
  7866=>"110011111",
  7867=>"001100001",
  7868=>"010011110",
  7869=>"000110010",
  7870=>"011110000",
  7871=>"011001010",
  7872=>"001011101",
  7873=>"111111101",
  7874=>"010101000",
  7875=>"111000110",
  7876=>"100001101",
  7877=>"101000111",
  7878=>"110110010",
  7879=>"110101001",
  7880=>"101010000",
  7881=>"101010110",
  7882=>"010101101",
  7883=>"001001001",
  7884=>"010110010",
  7885=>"110000010",
  7886=>"011101110",
  7887=>"011100011",
  7888=>"010110000",
  7889=>"100001000",
  7890=>"011011011",
  7891=>"111001110",
  7892=>"100101110",
  7893=>"100001111",
  7894=>"101101001",
  7895=>"101010111",
  7896=>"010111110",
  7897=>"001001011",
  7898=>"000100100",
  7899=>"111001010",
  7900=>"111000101",
  7901=>"110111111",
  7902=>"000000011",
  7903=>"100100100",
  7904=>"010101111",
  7905=>"000000010",
  7906=>"010101000",
  7907=>"001001101",
  7908=>"111010001",
  7909=>"111010011",
  7910=>"100110001",
  7911=>"000010110",
  7912=>"000001101",
  7913=>"001110111",
  7914=>"100100111",
  7915=>"000001110",
  7916=>"100111111",
  7917=>"110100111",
  7918=>"100011100",
  7919=>"101101101",
  7920=>"010010110",
  7921=>"001000010",
  7922=>"001001010",
  7923=>"110010110",
  7924=>"110111111",
  7925=>"000011111",
  7926=>"101110000",
  7927=>"011001100",
  7928=>"110111000",
  7929=>"010010110",
  7930=>"011010001",
  7931=>"101010001",
  7932=>"011011011",
  7933=>"110101001",
  7934=>"100000101",
  7935=>"010110101",
  7936=>"111001101",
  7937=>"100110101",
  7938=>"110010110",
  7939=>"110101110",
  7940=>"110001010",
  7941=>"100100010",
  7942=>"011011110",
  7943=>"111111101",
  7944=>"011000100",
  7945=>"100001111",
  7946=>"100110000",
  7947=>"010101100",
  7948=>"100000100",
  7949=>"100010100",
  7950=>"110000000",
  7951=>"110110000",
  7952=>"111101010",
  7953=>"101101001",
  7954=>"111110111",
  7955=>"100011110",
  7956=>"011100000",
  7957=>"100101001",
  7958=>"010000011",
  7959=>"000111100",
  7960=>"001101101",
  7961=>"001010001",
  7962=>"010001010",
  7963=>"011100011",
  7964=>"011101101",
  7965=>"111111101",
  7966=>"110100111",
  7967=>"101001100",
  7968=>"011000000",
  7969=>"100111011",
  7970=>"101111000",
  7971=>"010110001",
  7972=>"100100001",
  7973=>"110110000",
  7974=>"111110011",
  7975=>"000000000",
  7976=>"101011111",
  7977=>"100111011",
  7978=>"011000110",
  7979=>"111001101",
  7980=>"110011011",
  7981=>"010110011",
  7982=>"001111011",
  7983=>"110000101",
  7984=>"011110001",
  7985=>"011111010",
  7986=>"110001110",
  7987=>"100110111",
  7988=>"010100010",
  7989=>"010011000",
  7990=>"110111110",
  7991=>"100101100",
  7992=>"011110100",
  7993=>"110001111",
  7994=>"111101100",
  7995=>"111100000",
  7996=>"010011100",
  7997=>"011000100",
  7998=>"101110111",
  7999=>"001011111",
  8000=>"001101100",
  8001=>"000110110",
  8002=>"000100111",
  8003=>"001110100",
  8004=>"001001111",
  8005=>"011100101",
  8006=>"010001110",
  8007=>"100110011",
  8008=>"011011101",
  8009=>"000101000",
  8010=>"001110111",
  8011=>"001000110",
  8012=>"011011000",
  8013=>"010001000",
  8014=>"010100000",
  8015=>"110111111",
  8016=>"001011100",
  8017=>"100000000",
  8018=>"010110101",
  8019=>"010110100",
  8020=>"000000001",
  8021=>"010110001",
  8022=>"110101011",
  8023=>"000010111",
  8024=>"000011011",
  8025=>"110011100",
  8026=>"000000011",
  8027=>"111010000",
  8028=>"011000010",
  8029=>"001001000",
  8030=>"111010011",
  8031=>"100100000",
  8032=>"010110111",
  8033=>"100111101",
  8034=>"000001000",
  8035=>"111001010",
  8036=>"110000101",
  8037=>"000111010",
  8038=>"100010000",
  8039=>"111000011",
  8040=>"000000001",
  8041=>"010011111",
  8042=>"101110101",
  8043=>"010010001",
  8044=>"010011101",
  8045=>"101001101",
  8046=>"011101001",
  8047=>"001111110",
  8048=>"111111010",
  8049=>"110101011",
  8050=>"010100111",
  8051=>"011011100",
  8052=>"100101011",
  8053=>"101100001",
  8054=>"011011000",
  8055=>"000001001",
  8056=>"001001100",
  8057=>"000000110",
  8058=>"010111100",
  8059=>"110100100",
  8060=>"000110111",
  8061=>"110000010",
  8062=>"111010000",
  8063=>"111101111",
  8064=>"010110011",
  8065=>"000110001",
  8066=>"000001000",
  8067=>"001101000",
  8068=>"100010100",
  8069=>"011101010",
  8070=>"100011010",
  8071=>"100100100",
  8072=>"000010000",
  8073=>"000110111",
  8074=>"100101100",
  8075=>"001010001",
  8076=>"000111010",
  8077=>"111101111",
  8078=>"110110101",
  8079=>"000000110",
  8080=>"000011111",
  8081=>"100101101",
  8082=>"001100001",
  8083=>"010101011",
  8084=>"100001110",
  8085=>"110111111",
  8086=>"110101001",
  8087=>"101000000",
  8088=>"110111100",
  8089=>"010011000",
  8090=>"100111001",
  8091=>"010101010",
  8092=>"111000110",
  8093=>"011011111",
  8094=>"011101000",
  8095=>"001001100",
  8096=>"011000001",
  8097=>"011101001",
  8098=>"100110111",
  8099=>"010111000",
  8100=>"110110000",
  8101=>"010000001",
  8102=>"011110110",
  8103=>"100100001",
  8104=>"000000101",
  8105=>"001011010",
  8106=>"111111111",
  8107=>"101010101",
  8108=>"000010110",
  8109=>"011000001",
  8110=>"111100110",
  8111=>"010101100",
  8112=>"010001010",
  8113=>"111000101",
  8114=>"001001111",
  8115=>"101101111",
  8116=>"110000100",
  8117=>"001010100",
  8118=>"011100101",
  8119=>"001010011",
  8120=>"011000001",
  8121=>"011001000",
  8122=>"111001100",
  8123=>"000110100",
  8124=>"001100101",
  8125=>"111000010",
  8126=>"010100010",
  8127=>"010110011",
  8128=>"101000001",
  8129=>"011101101",
  8130=>"101110010",
  8131=>"111000101",
  8132=>"001101100",
  8133=>"011111001",
  8134=>"111000011",
  8135=>"000000001",
  8136=>"011001100",
  8137=>"111011111",
  8138=>"010100000",
  8139=>"001001011",
  8140=>"010101010",
  8141=>"111010011",
  8142=>"110001110",
  8143=>"110111100",
  8144=>"101110111",
  8145=>"010100010",
  8146=>"111101110",
  8147=>"111001000",
  8148=>"001000101",
  8149=>"111100100",
  8150=>"010000001",
  8151=>"001101100",
  8152=>"001111110",
  8153=>"110110101",
  8154=>"111010110",
  8155=>"001001101",
  8156=>"110000011",
  8157=>"010101110",
  8158=>"100010100",
  8159=>"101000101",
  8160=>"100110111",
  8161=>"000101100",
  8162=>"001111001",
  8163=>"100010110",
  8164=>"001100011",
  8165=>"100001101",
  8166=>"111111101",
  8167=>"010000001",
  8168=>"000010010",
  8169=>"110000011",
  8170=>"001111010",
  8171=>"110000000",
  8172=>"011011101",
  8173=>"101101100",
  8174=>"001111100",
  8175=>"110000111",
  8176=>"101011000",
  8177=>"111100111",
  8178=>"011110010",
  8179=>"011001111",
  8180=>"100010111",
  8181=>"010000001",
  8182=>"100111010",
  8183=>"011001011",
  8184=>"111111110",
  8185=>"010111001",
  8186=>"011010110",
  8187=>"100001111",
  8188=>"110100001",
  8189=>"101000110",
  8190=>"111000011",
  8191=>"010110000",
  8192=>"111100111",
  8193=>"100111111",
  8194=>"111110111",
  8195=>"010101010",
  8196=>"010000001",
  8197=>"101101111",
  8198=>"110111101",
  8199=>"111000000",
  8200=>"100000010",
  8201=>"100001100",
  8202=>"001000000",
  8203=>"111101010",
  8204=>"100011100",
  8205=>"100111111",
  8206=>"001101111",
  8207=>"000010111",
  8208=>"000000101",
  8209=>"101000000",
  8210=>"110000110",
  8211=>"111011110",
  8212=>"101100011",
  8213=>"100111110",
  8214=>"111010111",
  8215=>"001100101",
  8216=>"111101100",
  8217=>"010110011",
  8218=>"100111011",
  8219=>"001001010",
  8220=>"100011111",
  8221=>"100111000",
  8222=>"000000110",
  8223=>"010110101",
  8224=>"011111011",
  8225=>"011001001",
  8226=>"100100011",
  8227=>"101111000",
  8228=>"111001011",
  8229=>"110101000",
  8230=>"000010010",
  8231=>"101010101",
  8232=>"011010000",
  8233=>"000011011",
  8234=>"100100100",
  8235=>"001110011",
  8236=>"010111010",
  8237=>"100110110",
  8238=>"001100000",
  8239=>"110110101",
  8240=>"001001011",
  8241=>"101100011",
  8242=>"101110100",
  8243=>"001001111",
  8244=>"100110011",
  8245=>"010110000",
  8246=>"001000101",
  8247=>"101101011",
  8248=>"011001010",
  8249=>"001101011",
  8250=>"000001000",
  8251=>"111111001",
  8252=>"000011000",
  8253=>"110101000",
  8254=>"110111010",
  8255=>"011010100",
  8256=>"110000101",
  8257=>"100001010",
  8258=>"001100000",
  8259=>"101010111",
  8260=>"101000001",
  8261=>"101011010",
  8262=>"001001000",
  8263=>"000000101",
  8264=>"011000110",
  8265=>"101000110",
  8266=>"010101000",
  8267=>"111000001",
  8268=>"100111101",
  8269=>"011000100",
  8270=>"000010101",
  8271=>"001001001",
  8272=>"001110011",
  8273=>"001110001",
  8274=>"001101001",
  8275=>"010111100",
  8276=>"010100100",
  8277=>"000100000",
  8278=>"011000010",
  8279=>"001011000",
  8280=>"100001000",
  8281=>"010010110",
  8282=>"000101110",
  8283=>"100100001",
  8284=>"001000100",
  8285=>"101110000",
  8286=>"110111111",
  8287=>"111011111",
  8288=>"000000001",
  8289=>"100001000",
  8290=>"111001010",
  8291=>"100111100",
  8292=>"110101101",
  8293=>"100000100",
  8294=>"010110000",
  8295=>"110111000",
  8296=>"100010011",
  8297=>"110001001",
  8298=>"101111011",
  8299=>"010011000",
  8300=>"010111010",
  8301=>"000110000",
  8302=>"010000011",
  8303=>"100001001",
  8304=>"001101110",
  8305=>"001111010",
  8306=>"101101000",
  8307=>"010100010",
  8308=>"110000000",
  8309=>"011000000",
  8310=>"110010010",
  8311=>"000100000",
  8312=>"001000010",
  8313=>"011110010",
  8314=>"011000000",
  8315=>"000111000",
  8316=>"111110011",
  8317=>"010010011",
  8318=>"111101001",
  8319=>"110101111",
  8320=>"110101100",
  8321=>"010000000",
  8322=>"001000011",
  8323=>"100000000",
  8324=>"110111100",
  8325=>"101011001",
  8326=>"101001100",
  8327=>"001000100",
  8328=>"110101010",
  8329=>"001111011",
  8330=>"000010101",
  8331=>"010001000",
  8332=>"101011111",
  8333=>"011010001",
  8334=>"101001111",
  8335=>"010001010",
  8336=>"100011111",
  8337=>"111000010",
  8338=>"001010001",
  8339=>"111110011",
  8340=>"010000100",
  8341=>"110010100",
  8342=>"001001010",
  8343=>"000111010",
  8344=>"000001000",
  8345=>"011100000",
  8346=>"000110111",
  8347=>"100111000",
  8348=>"000101101",
  8349=>"010010000",
  8350=>"011010011",
  8351=>"010110011",
  8352=>"101111001",
  8353=>"101001100",
  8354=>"011100000",
  8355=>"001011111",
  8356=>"111011010",
  8357=>"111110110",
  8358=>"010110010",
  8359=>"010101111",
  8360=>"110101001",
  8361=>"000101010",
  8362=>"100011000",
  8363=>"001000101",
  8364=>"000100110",
  8365=>"100011000",
  8366=>"000000011",
  8367=>"001000000",
  8368=>"010111010",
  8369=>"101000010",
  8370=>"110001101",
  8371=>"010110111",
  8372=>"011101110",
  8373=>"010101000",
  8374=>"100101101",
  8375=>"010101100",
  8376=>"001010011",
  8377=>"011000101",
  8378=>"011011110",
  8379=>"010101101",
  8380=>"110010010",
  8381=>"100000000",
  8382=>"011001011",
  8383=>"000001000",
  8384=>"011101110",
  8385=>"111101100",
  8386=>"101000100",
  8387=>"001100110",
  8388=>"110100100",
  8389=>"000011000",
  8390=>"111000100",
  8391=>"010101100",
  8392=>"110101010",
  8393=>"001100100",
  8394=>"010000111",
  8395=>"011001100",
  8396=>"001110010",
  8397=>"000100010",
  8398=>"000101100",
  8399=>"010001000",
  8400=>"001110111",
  8401=>"000000000",
  8402=>"010000110",
  8403=>"011101111",
  8404=>"011111100",
  8405=>"011010101",
  8406=>"010000001",
  8407=>"001100111",
  8408=>"101010100",
  8409=>"010100001",
  8410=>"111001111",
  8411=>"110000101",
  8412=>"001001101",
  8413=>"000100100",
  8414=>"110101010",
  8415=>"001011110",
  8416=>"011011111",
  8417=>"110101010",
  8418=>"001000011",
  8419=>"001011101",
  8420=>"110111110",
  8421=>"110010101",
  8422=>"000001011",
  8423=>"101001000",
  8424=>"000100101",
  8425=>"101100100",
  8426=>"111011011",
  8427=>"000110000",
  8428=>"101001000",
  8429=>"001010011",
  8430=>"100010011",
  8431=>"110000010",
  8432=>"011000011",
  8433=>"101011001",
  8434=>"001001010",
  8435=>"001100001",
  8436=>"110110000",
  8437=>"001110001",
  8438=>"011001011",
  8439=>"101100110",
  8440=>"010011100",
  8441=>"011100011",
  8442=>"111000110",
  8443=>"011010100",
  8444=>"001000101",
  8445=>"000111010",
  8446=>"010101011",
  8447=>"011110000",
  8448=>"100001100",
  8449=>"010110101",
  8450=>"111110111",
  8451=>"000110101",
  8452=>"001010100",
  8453=>"001100010",
  8454=>"001011011",
  8455=>"100000010",
  8456=>"001000101",
  8457=>"010111001",
  8458=>"010101001",
  8459=>"100101100",
  8460=>"000101011",
  8461=>"101000100",
  8462=>"000000100",
  8463=>"011001010",
  8464=>"110110111",
  8465=>"111101101",
  8466=>"111111111",
  8467=>"111010111",
  8468=>"111111111",
  8469=>"101111000",
  8470=>"111100011",
  8471=>"000101110",
  8472=>"000100011",
  8473=>"000001110",
  8474=>"110101011",
  8475=>"000101101",
  8476=>"001010010",
  8477=>"010001011",
  8478=>"001110101",
  8479=>"100010010",
  8480=>"001100111",
  8481=>"000001001",
  8482=>"100111100",
  8483=>"001110101",
  8484=>"010101110",
  8485=>"100010001",
  8486=>"110100110",
  8487=>"111111101",
  8488=>"100100000",
  8489=>"110100101",
  8490=>"000001110",
  8491=>"001111011",
  8492=>"100111000",
  8493=>"100001010",
  8494=>"101010110",
  8495=>"110100100",
  8496=>"111101011",
  8497=>"010111100",
  8498=>"000111110",
  8499=>"101000101",
  8500=>"101110010",
  8501=>"010110000",
  8502=>"011010011",
  8503=>"110101011",
  8504=>"010011101",
  8505=>"001011001",
  8506=>"101100111",
  8507=>"101010000",
  8508=>"001101100",
  8509=>"100010001",
  8510=>"101011010",
  8511=>"101111011",
  8512=>"110111101",
  8513=>"000000001",
  8514=>"011110001",
  8515=>"000101001",
  8516=>"001111101",
  8517=>"110010001",
  8518=>"101111111",
  8519=>"110100010",
  8520=>"001110101",
  8521=>"101000001",
  8522=>"111110110",
  8523=>"001000101",
  8524=>"111110000",
  8525=>"111110001",
  8526=>"010011001",
  8527=>"101101111",
  8528=>"101001110",
  8529=>"110000010",
  8530=>"000111101",
  8531=>"111000010",
  8532=>"001011111",
  8533=>"000110110",
  8534=>"100101010",
  8535=>"001001011",
  8536=>"010000000",
  8537=>"110010001",
  8538=>"100010101",
  8539=>"101011110",
  8540=>"100000001",
  8541=>"110010110",
  8542=>"010000010",
  8543=>"010111100",
  8544=>"011010000",
  8545=>"111111001",
  8546=>"111100110",
  8547=>"010100001",
  8548=>"101101000",
  8549=>"101110011",
  8550=>"111100010",
  8551=>"101011110",
  8552=>"010110000",
  8553=>"010111011",
  8554=>"110001100",
  8555=>"100111000",
  8556=>"100000001",
  8557=>"110100010",
  8558=>"111011110",
  8559=>"011101000",
  8560=>"000101100",
  8561=>"100001000",
  8562=>"001011001",
  8563=>"010011000",
  8564=>"001101100",
  8565=>"010001010",
  8566=>"111100101",
  8567=>"111110010",
  8568=>"001000000",
  8569=>"100000100",
  8570=>"011100100",
  8571=>"101111000",
  8572=>"110001000",
  8573=>"100101110",
  8574=>"111000101",
  8575=>"111100000",
  8576=>"001011011",
  8577=>"001000001",
  8578=>"001110111",
  8579=>"010111111",
  8580=>"000100011",
  8581=>"101101100",
  8582=>"110111101",
  8583=>"001101100",
  8584=>"000100101",
  8585=>"010101100",
  8586=>"000000101",
  8587=>"110011101",
  8588=>"011100011",
  8589=>"101111100",
  8590=>"000000000",
  8591=>"011111111",
  8592=>"111111001",
  8593=>"111100000",
  8594=>"010110000",
  8595=>"001011111",
  8596=>"110001011",
  8597=>"000001101",
  8598=>"000010010",
  8599=>"101010000",
  8600=>"011101010",
  8601=>"110001101",
  8602=>"010111011",
  8603=>"100100100",
  8604=>"110010100",
  8605=>"011001000",
  8606=>"010110011",
  8607=>"001101001",
  8608=>"001000100",
  8609=>"101011011",
  8610=>"110001011",
  8611=>"011000000",
  8612=>"101000001",
  8613=>"011101111",
  8614=>"001100101",
  8615=>"001100001",
  8616=>"100111000",
  8617=>"100001101",
  8618=>"011101100",
  8619=>"110011100",
  8620=>"101111001",
  8621=>"010010000",
  8622=>"111100111",
  8623=>"001110011",
  8624=>"111101111",
  8625=>"110000100",
  8626=>"001001111",
  8627=>"000010000",
  8628=>"101001001",
  8629=>"000110011",
  8630=>"011101000",
  8631=>"011100000",
  8632=>"101001101",
  8633=>"100111010",
  8634=>"100011000",
  8635=>"000000001",
  8636=>"011110010",
  8637=>"111101000",
  8638=>"000000000",
  8639=>"111010010",
  8640=>"011010000",
  8641=>"111011110",
  8642=>"111000110",
  8643=>"010001000",
  8644=>"010000011",
  8645=>"100100101",
  8646=>"100000010",
  8647=>"001010111",
  8648=>"111001100",
  8649=>"110011100",
  8650=>"110000101",
  8651=>"001000001",
  8652=>"100111001",
  8653=>"101000001",
  8654=>"001011110",
  8655=>"001011001",
  8656=>"010000010",
  8657=>"110010101",
  8658=>"110000111",
  8659=>"110001000",
  8660=>"101101001",
  8661=>"110100011",
  8662=>"000000111",
  8663=>"011110110",
  8664=>"011110011",
  8665=>"110111011",
  8666=>"110000101",
  8667=>"111110011",
  8668=>"010111011",
  8669=>"100011010",
  8670=>"011000001",
  8671=>"010000110",
  8672=>"100110111",
  8673=>"111011111",
  8674=>"000011111",
  8675=>"011011111",
  8676=>"001001000",
  8677=>"010000011",
  8678=>"011111100",
  8679=>"101000100",
  8680=>"101100001",
  8681=>"010011011",
  8682=>"001100010",
  8683=>"110111011",
  8684=>"100011100",
  8685=>"000011101",
  8686=>"000011111",
  8687=>"101110111",
  8688=>"011100101",
  8689=>"001000110",
  8690=>"101101111",
  8691=>"101000010",
  8692=>"010000110",
  8693=>"010010100",
  8694=>"110010100",
  8695=>"100110000",
  8696=>"001000101",
  8697=>"011111110",
  8698=>"111000101",
  8699=>"000100000",
  8700=>"000000011",
  8701=>"101010111",
  8702=>"101110101",
  8703=>"101001101",
  8704=>"101001001",
  8705=>"001000001",
  8706=>"001100101",
  8707=>"011000110",
  8708=>"100111010",
  8709=>"000000010",
  8710=>"100001010",
  8711=>"001001111",
  8712=>"000111101",
  8713=>"001101110",
  8714=>"111010101",
  8715=>"111111001",
  8716=>"101010100",
  8717=>"111010011",
  8718=>"010011100",
  8719=>"101110001",
  8720=>"011111011",
  8721=>"010000001",
  8722=>"110110100",
  8723=>"110110011",
  8724=>"010100010",
  8725=>"100001100",
  8726=>"111111101",
  8727=>"010110110",
  8728=>"100000100",
  8729=>"011111010",
  8730=>"011010000",
  8731=>"101110100",
  8732=>"001111011",
  8733=>"010101000",
  8734=>"111101011",
  8735=>"010110001",
  8736=>"011110101",
  8737=>"101110100",
  8738=>"100010101",
  8739=>"100110000",
  8740=>"100011010",
  8741=>"001001110",
  8742=>"101100001",
  8743=>"010100010",
  8744=>"110000111",
  8745=>"100101011",
  8746=>"100011100",
  8747=>"000110100",
  8748=>"010100001",
  8749=>"111111101",
  8750=>"010001010",
  8751=>"111010111",
  8752=>"010100101",
  8753=>"111010111",
  8754=>"101001001",
  8755=>"110011110",
  8756=>"000000111",
  8757=>"011101011",
  8758=>"110101111",
  8759=>"100111000",
  8760=>"111000111",
  8761=>"010011100",
  8762=>"001010010",
  8763=>"010000100",
  8764=>"110101111",
  8765=>"100110100",
  8766=>"101001001",
  8767=>"100101100",
  8768=>"100111111",
  8769=>"011011110",
  8770=>"001011001",
  8771=>"000100110",
  8772=>"100010111",
  8773=>"111011110",
  8774=>"001101011",
  8775=>"010001000",
  8776=>"010000100",
  8777=>"001000100",
  8778=>"101000101",
  8779=>"111010101",
  8780=>"110000011",
  8781=>"000011000",
  8782=>"100111001",
  8783=>"011101111",
  8784=>"010101000",
  8785=>"111101001",
  8786=>"011111111",
  8787=>"011010011",
  8788=>"110011010",
  8789=>"010111101",
  8790=>"000000101",
  8791=>"011110011",
  8792=>"101000100",
  8793=>"101000101",
  8794=>"101100001",
  8795=>"111111010",
  8796=>"000000001",
  8797=>"010111111",
  8798=>"001110101",
  8799=>"100111010",
  8800=>"100000100",
  8801=>"011011000",
  8802=>"001100101",
  8803=>"100101010",
  8804=>"000011010",
  8805=>"010101111",
  8806=>"011010110",
  8807=>"001111111",
  8808=>"110010010",
  8809=>"100110001",
  8810=>"100010100",
  8811=>"111100010",
  8812=>"001000101",
  8813=>"110101000",
  8814=>"000011110",
  8815=>"011010001",
  8816=>"001010010",
  8817=>"111101011",
  8818=>"000001011",
  8819=>"111011101",
  8820=>"110010111",
  8821=>"110011000",
  8822=>"001010000",
  8823=>"111010100",
  8824=>"001010110",
  8825=>"011011011",
  8826=>"101001100",
  8827=>"011100000",
  8828=>"111110100",
  8829=>"101110101",
  8830=>"001011000",
  8831=>"001000010",
  8832=>"011011001",
  8833=>"010000111",
  8834=>"111101011",
  8835=>"110001110",
  8836=>"110000001",
  8837=>"111111000",
  8838=>"110100100",
  8839=>"011011010",
  8840=>"011001110",
  8841=>"001100110",
  8842=>"111101100",
  8843=>"000001101",
  8844=>"101000100",
  8845=>"001101011",
  8846=>"010000101",
  8847=>"000100111",
  8848=>"001100100",
  8849=>"001000111",
  8850=>"001100111",
  8851=>"101010001",
  8852=>"000001110",
  8853=>"101000000",
  8854=>"110010100",
  8855=>"001101000",
  8856=>"001100111",
  8857=>"111111010",
  8858=>"000010100",
  8859=>"111101111",
  8860=>"011100101",
  8861=>"100011101",
  8862=>"100011100",
  8863=>"100001100",
  8864=>"101111011",
  8865=>"011111110",
  8866=>"110100101",
  8867=>"001101011",
  8868=>"001101000",
  8869=>"000011011",
  8870=>"110000010",
  8871=>"010110111",
  8872=>"110001011",
  8873=>"110101011",
  8874=>"011110000",
  8875=>"101101100",
  8876=>"001100100",
  8877=>"111111110",
  8878=>"101011000",
  8879=>"100011100",
  8880=>"101011010",
  8881=>"100010000",
  8882=>"001001101",
  8883=>"010000110",
  8884=>"011110011",
  8885=>"010010011",
  8886=>"101100111",
  8887=>"101000001",
  8888=>"011011011",
  8889=>"110001100",
  8890=>"111011100",
  8891=>"101110110",
  8892=>"001100011",
  8893=>"011011111",
  8894=>"001101000",
  8895=>"101001100",
  8896=>"011010010",
  8897=>"110001110",
  8898=>"100000101",
  8899=>"100011111",
  8900=>"011010010",
  8901=>"111100010",
  8902=>"111111110",
  8903=>"110111001",
  8904=>"010001000",
  8905=>"010101000",
  8906=>"000110010",
  8907=>"011110100",
  8908=>"101110000",
  8909=>"110000011",
  8910=>"001100010",
  8911=>"011101000",
  8912=>"101111011",
  8913=>"111011001",
  8914=>"111010101",
  8915=>"001000001",
  8916=>"100000111",
  8917=>"011010110",
  8918=>"101110001",
  8919=>"111000110",
  8920=>"001011011",
  8921=>"110111101",
  8922=>"111000111",
  8923=>"110011000",
  8924=>"000000110",
  8925=>"110001101",
  8926=>"000100011",
  8927=>"011110100",
  8928=>"001000000",
  8929=>"101101000",
  8930=>"001110000",
  8931=>"001110111",
  8932=>"101001111",
  8933=>"010000010",
  8934=>"001101010",
  8935=>"110000100",
  8936=>"000000100",
  8937=>"100011111",
  8938=>"101011101",
  8939=>"110010101",
  8940=>"110010110",
  8941=>"010001010",
  8942=>"111010110",
  8943=>"111100111",
  8944=>"001010101",
  8945=>"000010101",
  8946=>"111010110",
  8947=>"110110001",
  8948=>"001110000",
  8949=>"010110110",
  8950=>"101001111",
  8951=>"111100100",
  8952=>"100000101",
  8953=>"101011000",
  8954=>"111011000",
  8955=>"010111101",
  8956=>"110110010",
  8957=>"010000001",
  8958=>"110100011",
  8959=>"001001110",
  8960=>"010001100",
  8961=>"001001000",
  8962=>"000011000",
  8963=>"001001011",
  8964=>"010011001",
  8965=>"101110001",
  8966=>"111110110",
  8967=>"001000010",
  8968=>"000001011",
  8969=>"011111100",
  8970=>"100011000",
  8971=>"111011111",
  8972=>"010000011",
  8973=>"111011011",
  8974=>"111100100",
  8975=>"110100000",
  8976=>"000010001",
  8977=>"110100101",
  8978=>"001001101",
  8979=>"000110000",
  8980=>"000101110",
  8981=>"100000010",
  8982=>"110101111",
  8983=>"010110000",
  8984=>"101101001",
  8985=>"110100101",
  8986=>"010011001",
  8987=>"111001100",
  8988=>"101000101",
  8989=>"111101100",
  8990=>"101100000",
  8991=>"101111010",
  8992=>"100111111",
  8993=>"111011001",
  8994=>"011101000",
  8995=>"010001010",
  8996=>"000101110",
  8997=>"011110000",
  8998=>"110010110",
  8999=>"001101100",
  9000=>"101000000",
  9001=>"001100011",
  9002=>"001110000",
  9003=>"001011100",
  9004=>"011011101",
  9005=>"011011100",
  9006=>"111101011",
  9007=>"100001110",
  9008=>"000000100",
  9009=>"101001011",
  9010=>"010110011",
  9011=>"100111110",
  9012=>"101001010",
  9013=>"111111111",
  9014=>"010100011",
  9015=>"010001111",
  9016=>"100101111",
  9017=>"110011110",
  9018=>"101000010",
  9019=>"011001111",
  9020=>"111000000",
  9021=>"110000101",
  9022=>"010101000",
  9023=>"111001101",
  9024=>"101011011",
  9025=>"000000100",
  9026=>"001011101",
  9027=>"000111100",
  9028=>"001110011",
  9029=>"000101010",
  9030=>"101101001",
  9031=>"011000001",
  9032=>"001110100",
  9033=>"011110000",
  9034=>"110110010",
  9035=>"000001100",
  9036=>"100011000",
  9037=>"001000111",
  9038=>"011011100",
  9039=>"010011010",
  9040=>"001100011",
  9041=>"101001111",
  9042=>"111101111",
  9043=>"110101011",
  9044=>"111001110",
  9045=>"100101110",
  9046=>"011011001",
  9047=>"100100001",
  9048=>"110001101",
  9049=>"011010110",
  9050=>"110001110",
  9051=>"000100110",
  9052=>"110101000",
  9053=>"001000011",
  9054=>"011000000",
  9055=>"100110111",
  9056=>"011110101",
  9057=>"111110001",
  9058=>"000111100",
  9059=>"011000101",
  9060=>"011101010",
  9061=>"110010100",
  9062=>"100011010",
  9063=>"100110000",
  9064=>"000011001",
  9065=>"110111000",
  9066=>"001011000",
  9067=>"101001000",
  9068=>"010110010",
  9069=>"010011000",
  9070=>"111110110",
  9071=>"001111000",
  9072=>"110010001",
  9073=>"111000000",
  9074=>"001010001",
  9075=>"110011111",
  9076=>"101101001",
  9077=>"111100111",
  9078=>"100100101",
  9079=>"101111100",
  9080=>"010011000",
  9081=>"110110100",
  9082=>"001100110",
  9083=>"111110111",
  9084=>"100101111",
  9085=>"011010011",
  9086=>"001010101",
  9087=>"001010010",
  9088=>"010111101",
  9089=>"000111000",
  9090=>"111001001",
  9091=>"111100110",
  9092=>"110101010",
  9093=>"100010101",
  9094=>"111101011",
  9095=>"111100000",
  9096=>"111011110",
  9097=>"111111001",
  9098=>"110110000",
  9099=>"110110111",
  9100=>"111000101",
  9101=>"010101110",
  9102=>"011000011",
  9103=>"110101001",
  9104=>"101000011",
  9105=>"111111111",
  9106=>"100011100",
  9107=>"111001011",
  9108=>"100001010",
  9109=>"011111111",
  9110=>"110001100",
  9111=>"011001011",
  9112=>"000001110",
  9113=>"111000110",
  9114=>"111111000",
  9115=>"001101001",
  9116=>"000100011",
  9117=>"000010000",
  9118=>"100000001",
  9119=>"011001111",
  9120=>"110011011",
  9121=>"010010011",
  9122=>"100101001",
  9123=>"111111001",
  9124=>"101000000",
  9125=>"111011101",
  9126=>"111101001",
  9127=>"101000111",
  9128=>"000010001",
  9129=>"000100011",
  9130=>"011010111",
  9131=>"010100010",
  9132=>"010100111",
  9133=>"000010111",
  9134=>"010100110",
  9135=>"011011111",
  9136=>"010101101",
  9137=>"011111000",
  9138=>"101100111",
  9139=>"011001101",
  9140=>"100000111",
  9141=>"001110010",
  9142=>"001010010",
  9143=>"110100100",
  9144=>"100100100",
  9145=>"111100111",
  9146=>"010111101",
  9147=>"110011110",
  9148=>"001111010",
  9149=>"111001100",
  9150=>"101000101",
  9151=>"000000000",
  9152=>"110110001",
  9153=>"010011101",
  9154=>"100100111",
  9155=>"001111010",
  9156=>"100011110",
  9157=>"000110101",
  9158=>"101110110",
  9159=>"111100010",
  9160=>"100001000",
  9161=>"111110001",
  9162=>"010000001",
  9163=>"010111010",
  9164=>"100011001",
  9165=>"000010110",
  9166=>"001110001",
  9167=>"100110100",
  9168=>"100111101",
  9169=>"000100110",
  9170=>"000000001",
  9171=>"101101011",
  9172=>"110010100",
  9173=>"010101001",
  9174=>"101011000",
  9175=>"011010000",
  9176=>"001010011",
  9177=>"011110010",
  9178=>"001000011",
  9179=>"111111010",
  9180=>"000000111",
  9181=>"101111000",
  9182=>"001001111",
  9183=>"001001101",
  9184=>"001101000",
  9185=>"001001010",
  9186=>"101000010",
  9187=>"110111110",
  9188=>"001110010",
  9189=>"011010101",
  9190=>"111110100",
  9191=>"101001100",
  9192=>"100100101",
  9193=>"000011111",
  9194=>"110000100",
  9195=>"000010011",
  9196=>"001000011",
  9197=>"001100001",
  9198=>"110010111",
  9199=>"111001001",
  9200=>"000000110",
  9201=>"011100001",
  9202=>"010000010",
  9203=>"100001110",
  9204=>"011110010",
  9205=>"111100101",
  9206=>"001001110",
  9207=>"110111001",
  9208=>"101011001",
  9209=>"001000110",
  9210=>"010111101",
  9211=>"101001001",
  9212=>"011101010",
  9213=>"100101010",
  9214=>"110001100",
  9215=>"011111110",
  9216=>"101111101",
  9217=>"111001010",
  9218=>"001111111",
  9219=>"010100001",
  9220=>"110110011",
  9221=>"100011011",
  9222=>"100101110",
  9223=>"000100111",
  9224=>"101000000",
  9225=>"111011010",
  9226=>"110110100",
  9227=>"110100000",
  9228=>"101100111",
  9229=>"101010011",
  9230=>"010110001",
  9231=>"011011111",
  9232=>"010101000",
  9233=>"000010010",
  9234=>"111101000",
  9235=>"010111101",
  9236=>"101101100",
  9237=>"110011001",
  9238=>"010011010",
  9239=>"100100111",
  9240=>"000000001",
  9241=>"010011011",
  9242=>"000000010",
  9243=>"011110000",
  9244=>"110011011",
  9245=>"001101110",
  9246=>"110001011",
  9247=>"001000111",
  9248=>"010011101",
  9249=>"100101101",
  9250=>"111001101",
  9251=>"110110011",
  9252=>"111101001",
  9253=>"110111011",
  9254=>"100110000",
  9255=>"010011011",
  9256=>"111011001",
  9257=>"001100101",
  9258=>"000110111",
  9259=>"000000001",
  9260=>"010111110",
  9261=>"110111000",
  9262=>"001110000",
  9263=>"011010000",
  9264=>"101111100",
  9265=>"011010111",
  9266=>"100101001",
  9267=>"100000110",
  9268=>"111100110",
  9269=>"110100001",
  9270=>"010010111",
  9271=>"010000001",
  9272=>"101100111",
  9273=>"011101110",
  9274=>"000001111",
  9275=>"011001100",
  9276=>"011101111",
  9277=>"010011011",
  9278=>"000011110",
  9279=>"110010010",
  9280=>"000010110",
  9281=>"010000101",
  9282=>"001010000",
  9283=>"010001100",
  9284=>"010100000",
  9285=>"010000000",
  9286=>"111100010",
  9287=>"000011111",
  9288=>"110001111",
  9289=>"010011100",
  9290=>"010001100",
  9291=>"001011000",
  9292=>"001111000",
  9293=>"000000010",
  9294=>"111001001",
  9295=>"100001000",
  9296=>"000100100",
  9297=>"110011011",
  9298=>"001100001",
  9299=>"101100010",
  9300=>"001101000",
  9301=>"100111111",
  9302=>"111000000",
  9303=>"000000111",
  9304=>"011111100",
  9305=>"001000001",
  9306=>"110011100",
  9307=>"110010101",
  9308=>"100011000",
  9309=>"110110111",
  9310=>"001100000",
  9311=>"000010101",
  9312=>"110110101",
  9313=>"111100100",
  9314=>"000011000",
  9315=>"011000000",
  9316=>"111111010",
  9317=>"001110010",
  9318=>"111011101",
  9319=>"011100001",
  9320=>"000010101",
  9321=>"000001111",
  9322=>"100101100",
  9323=>"010111000",
  9324=>"001001110",
  9325=>"101000010",
  9326=>"111010000",
  9327=>"000011000",
  9328=>"011011100",
  9329=>"101000010",
  9330=>"001100011",
  9331=>"001000010",
  9332=>"011000111",
  9333=>"010000110",
  9334=>"100000111",
  9335=>"111010000",
  9336=>"000101100",
  9337=>"000010011",
  9338=>"001100000",
  9339=>"011111011",
  9340=>"110011001",
  9341=>"110110010",
  9342=>"001110000",
  9343=>"010111000",
  9344=>"010000011",
  9345=>"111111110",
  9346=>"010101110",
  9347=>"001110011",
  9348=>"001011100",
  9349=>"001111111",
  9350=>"111101011",
  9351=>"100100100",
  9352=>"101110000",
  9353=>"100111000",
  9354=>"100000100",
  9355=>"111111110",
  9356=>"110000000",
  9357=>"010011010",
  9358=>"100101101",
  9359=>"010101011",
  9360=>"111110011",
  9361=>"101111110",
  9362=>"100011110",
  9363=>"010101000",
  9364=>"010101000",
  9365=>"000011001",
  9366=>"011101101",
  9367=>"010111010",
  9368=>"101000110",
  9369=>"010101010",
  9370=>"000010010",
  9371=>"011001010",
  9372=>"001001001",
  9373=>"110010000",
  9374=>"000101011",
  9375=>"111011111",
  9376=>"010111000",
  9377=>"000110000",
  9378=>"000101000",
  9379=>"100011111",
  9380=>"001100101",
  9381=>"100101010",
  9382=>"011110101",
  9383=>"011011001",
  9384=>"000000011",
  9385=>"010000010",
  9386=>"000110000",
  9387=>"100111111",
  9388=>"100010110",
  9389=>"011000110",
  9390=>"100100011",
  9391=>"101000111",
  9392=>"011011001",
  9393=>"111001101",
  9394=>"111101110",
  9395=>"110100011",
  9396=>"000111110",
  9397=>"100001001",
  9398=>"001000111",
  9399=>"101100101",
  9400=>"100111000",
  9401=>"101101000",
  9402=>"100100111",
  9403=>"010011110",
  9404=>"101100001",
  9405=>"101111101",
  9406=>"011000000",
  9407=>"100101001",
  9408=>"100011110",
  9409=>"111011110",
  9410=>"001001101",
  9411=>"001010000",
  9412=>"100010100",
  9413=>"111111111",
  9414=>"001111111",
  9415=>"100101101",
  9416=>"110000011",
  9417=>"101011101",
  9418=>"110110100",
  9419=>"111111010",
  9420=>"100011101",
  9421=>"101110100",
  9422=>"111001110",
  9423=>"100110110",
  9424=>"010110100",
  9425=>"111110010",
  9426=>"010100101",
  9427=>"010010010",
  9428=>"111001110",
  9429=>"011110101",
  9430=>"111001001",
  9431=>"110110001",
  9432=>"010100101",
  9433=>"111000010",
  9434=>"111101001",
  9435=>"101001101",
  9436=>"010110111",
  9437=>"000100111",
  9438=>"100010000",
  9439=>"011110010",
  9440=>"001100100",
  9441=>"111101111",
  9442=>"001110000",
  9443=>"000101100",
  9444=>"100101010",
  9445=>"010101011",
  9446=>"111110101",
  9447=>"010000011",
  9448=>"000110110",
  9449=>"000011110",
  9450=>"100010100",
  9451=>"000101000",
  9452=>"100010000",
  9453=>"011100111",
  9454=>"111010010",
  9455=>"010111001",
  9456=>"001011100",
  9457=>"110111111",
  9458=>"100000111",
  9459=>"011000011",
  9460=>"110011011",
  9461=>"001101100",
  9462=>"100111110",
  9463=>"001111011",
  9464=>"101100011",
  9465=>"110111101",
  9466=>"000001000",
  9467=>"100100000",
  9468=>"110011100",
  9469=>"011101011",
  9470=>"101011100",
  9471=>"111000010",
  9472=>"011110011",
  9473=>"000100110",
  9474=>"101101010",
  9475=>"100001101",
  9476=>"110011001",
  9477=>"001001100",
  9478=>"111110111",
  9479=>"101101000",
  9480=>"100101111",
  9481=>"001000011",
  9482=>"010011011",
  9483=>"000101011",
  9484=>"100011010",
  9485=>"100111010",
  9486=>"110000100",
  9487=>"000010101",
  9488=>"011000001",
  9489=>"101010101",
  9490=>"101000010",
  9491=>"000010001",
  9492=>"111000110",
  9493=>"001101101",
  9494=>"101110101",
  9495=>"111000010",
  9496=>"010110110",
  9497=>"001101001",
  9498=>"010101100",
  9499=>"110011001",
  9500=>"100011100",
  9501=>"100011010",
  9502=>"000001000",
  9503=>"001100001",
  9504=>"000011010",
  9505=>"001000100",
  9506=>"110011010",
  9507=>"010010000",
  9508=>"110110100",
  9509=>"101100010",
  9510=>"011001001",
  9511=>"011010000",
  9512=>"001111110",
  9513=>"100100110",
  9514=>"101000101",
  9515=>"011110000",
  9516=>"110110111",
  9517=>"110010101",
  9518=>"011101110",
  9519=>"111111110",
  9520=>"001100000",
  9521=>"100000111",
  9522=>"110100001",
  9523=>"110001011",
  9524=>"100110111",
  9525=>"010100110",
  9526=>"001110101",
  9527=>"000110000",
  9528=>"001001101",
  9529=>"101001111",
  9530=>"111111100",
  9531=>"011001000",
  9532=>"000000111",
  9533=>"001100001",
  9534=>"011100110",
  9535=>"100111111",
  9536=>"100111100",
  9537=>"000100011",
  9538=>"111100111",
  9539=>"111010111",
  9540=>"001100000",
  9541=>"000001010",
  9542=>"110101011",
  9543=>"000110101",
  9544=>"101000001",
  9545=>"010001101",
  9546=>"001011111",
  9547=>"101010011",
  9548=>"101011101",
  9549=>"010010101",
  9550=>"011111101",
  9551=>"010101110",
  9552=>"100100000",
  9553=>"010000101",
  9554=>"010001100",
  9555=>"111011111",
  9556=>"100010101",
  9557=>"101111111",
  9558=>"110101000",
  9559=>"011110000",
  9560=>"001100011",
  9561=>"101100101",
  9562=>"000100101",
  9563=>"000101011",
  9564=>"101010011",
  9565=>"101110100",
  9566=>"111110011",
  9567=>"101111101",
  9568=>"100000001",
  9569=>"000011011",
  9570=>"010011110",
  9571=>"001111100",
  9572=>"001000000",
  9573=>"001111011",
  9574=>"101011001",
  9575=>"000000101",
  9576=>"101010010",
  9577=>"111010010",
  9578=>"000000011",
  9579=>"001001110",
  9580=>"011011000",
  9581=>"000111101",
  9582=>"111000011",
  9583=>"000110011",
  9584=>"100011100",
  9585=>"000010010",
  9586=>"011110001",
  9587=>"001001010",
  9588=>"111001010",
  9589=>"110100111",
  9590=>"101101011",
  9591=>"101011001",
  9592=>"110100100",
  9593=>"010100111",
  9594=>"111111111",
  9595=>"011010111",
  9596=>"111011111",
  9597=>"111111110",
  9598=>"101100111",
  9599=>"001110100",
  9600=>"101101111",
  9601=>"011100000",
  9602=>"010010000",
  9603=>"010111000",
  9604=>"011000010",
  9605=>"000110101",
  9606=>"000011110",
  9607=>"101101110",
  9608=>"111000011",
  9609=>"011010001",
  9610=>"101011001",
  9611=>"010000001",
  9612=>"001000010",
  9613=>"010010010",
  9614=>"000000101",
  9615=>"011110001",
  9616=>"001000001",
  9617=>"101000010",
  9618=>"010101111",
  9619=>"111001000",
  9620=>"111111110",
  9621=>"010010000",
  9622=>"100100000",
  9623=>"010000010",
  9624=>"011001000",
  9625=>"001001111",
  9626=>"111011110",
  9627=>"001010010",
  9628=>"010111000",
  9629=>"001111001",
  9630=>"110001001",
  9631=>"110111011",
  9632=>"100100000",
  9633=>"101000101",
  9634=>"011110111",
  9635=>"100001011",
  9636=>"110000101",
  9637=>"111000001",
  9638=>"101011000",
  9639=>"101111100",
  9640=>"010010001",
  9641=>"000000111",
  9642=>"000000000",
  9643=>"001000111",
  9644=>"011100110",
  9645=>"000011010",
  9646=>"111001111",
  9647=>"101100101",
  9648=>"101100100",
  9649=>"111101111",
  9650=>"000010101",
  9651=>"100000001",
  9652=>"001111011",
  9653=>"100000110",
  9654=>"001101101",
  9655=>"010100010",
  9656=>"001101000",
  9657=>"110010111",
  9658=>"110101110",
  9659=>"000000001",
  9660=>"111001011",
  9661=>"111001011",
  9662=>"010101010",
  9663=>"000000011",
  9664=>"010001000",
  9665=>"111001110",
  9666=>"101111001",
  9667=>"010111100",
  9668=>"010100101",
  9669=>"111101101",
  9670=>"001000110",
  9671=>"111100101",
  9672=>"110001011",
  9673=>"011111110",
  9674=>"001101111",
  9675=>"011011001",
  9676=>"101111000",
  9677=>"010001001",
  9678=>"101110100",
  9679=>"011010100",
  9680=>"101001110",
  9681=>"111010001",
  9682=>"011101001",
  9683=>"101001111",
  9684=>"101111010",
  9685=>"010100001",
  9686=>"101010000",
  9687=>"111000001",
  9688=>"110110011",
  9689=>"111010100",
  9690=>"000100001",
  9691=>"101000100",
  9692=>"010101111",
  9693=>"111110001",
  9694=>"010111111",
  9695=>"010001110",
  9696=>"011011001",
  9697=>"001101000",
  9698=>"110100110",
  9699=>"101110111",
  9700=>"011100100",
  9701=>"000110100",
  9702=>"110110111",
  9703=>"111001001",
  9704=>"011001011",
  9705=>"111111111",
  9706=>"000010101",
  9707=>"001111101",
  9708=>"101111101",
  9709=>"010101101",
  9710=>"011001111",
  9711=>"011001100",
  9712=>"110110100",
  9713=>"101010111",
  9714=>"100010111",
  9715=>"001101001",
  9716=>"101010111",
  9717=>"001100001",
  9718=>"001110111",
  9719=>"011111111",
  9720=>"000111110",
  9721=>"000011010",
  9722=>"100010100",
  9723=>"101101110",
  9724=>"100110001",
  9725=>"100111011",
  9726=>"111101111",
  9727=>"011100100",
  9728=>"110110101",
  9729=>"111100111",
  9730=>"011010101",
  9731=>"001001111",
  9732=>"011100101",
  9733=>"010101000",
  9734=>"101110110",
  9735=>"100010011",
  9736=>"011101011",
  9737=>"001000000",
  9738=>"000010111",
  9739=>"011001001",
  9740=>"000001000",
  9741=>"001101110",
  9742=>"100000000",
  9743=>"001111000",
  9744=>"010010100",
  9745=>"100000110",
  9746=>"101001011",
  9747=>"000001011",
  9748=>"010100101",
  9749=>"010111111",
  9750=>"001100011",
  9751=>"110001010",
  9752=>"111000110",
  9753=>"101110111",
  9754=>"100001101",
  9755=>"111001100",
  9756=>"000000111",
  9757=>"010100110",
  9758=>"001001001",
  9759=>"000001000",
  9760=>"101100011",
  9761=>"011100111",
  9762=>"000000010",
  9763=>"100111011",
  9764=>"111100011",
  9765=>"100010011",
  9766=>"010001110",
  9767=>"011111011",
  9768=>"100111010",
  9769=>"011011001",
  9770=>"110010011",
  9771=>"101011111",
  9772=>"111100100",
  9773=>"010000110",
  9774=>"111101111",
  9775=>"110101010",
  9776=>"010011111",
  9777=>"110100110",
  9778=>"111001111",
  9779=>"000010000",
  9780=>"001011110",
  9781=>"000101100",
  9782=>"001110110",
  9783=>"101001101",
  9784=>"111111001",
  9785=>"111101100",
  9786=>"111000100",
  9787=>"001001000",
  9788=>"000010010",
  9789=>"001000001",
  9790=>"000001000",
  9791=>"010000101",
  9792=>"111110101",
  9793=>"110011111",
  9794=>"110100000",
  9795=>"001001101",
  9796=>"000111110",
  9797=>"011011010",
  9798=>"011111000",
  9799=>"000100011",
  9800=>"101010010",
  9801=>"001000100",
  9802=>"101101101",
  9803=>"100101010",
  9804=>"110000001",
  9805=>"101100010",
  9806=>"101000111",
  9807=>"010100011",
  9808=>"001010010",
  9809=>"010110111",
  9810=>"001111000",
  9811=>"111000011",
  9812=>"010010011",
  9813=>"000100110",
  9814=>"001111000",
  9815=>"001000000",
  9816=>"100111000",
  9817=>"100100111",
  9818=>"100101111",
  9819=>"100001010",
  9820=>"101010000",
  9821=>"000010000",
  9822=>"100010111",
  9823=>"001111101",
  9824=>"010101000",
  9825=>"010000001",
  9826=>"001001101",
  9827=>"011011011",
  9828=>"111011101",
  9829=>"110010011",
  9830=>"011101101",
  9831=>"110001111",
  9832=>"001010001",
  9833=>"001000110",
  9834=>"010000100",
  9835=>"100110000",
  9836=>"111101000",
  9837=>"001111011",
  9838=>"000010111",
  9839=>"100110100",
  9840=>"110100110",
  9841=>"010011001",
  9842=>"010001101",
  9843=>"100011001",
  9844=>"100100111",
  9845=>"010001000",
  9846=>"001111101",
  9847=>"111000101",
  9848=>"100011010",
  9849=>"101101001",
  9850=>"001100011",
  9851=>"000100000",
  9852=>"000000011",
  9853=>"110110011",
  9854=>"110100000",
  9855=>"101001010",
  9856=>"111111101",
  9857=>"000110110",
  9858=>"110100001",
  9859=>"001011110",
  9860=>"111011111",
  9861=>"101011000",
  9862=>"110110010",
  9863=>"010100010",
  9864=>"111011010",
  9865=>"001101111",
  9866=>"001011110",
  9867=>"010001111",
  9868=>"111011001",
  9869=>"001100011",
  9870=>"100101001",
  9871=>"101110000",
  9872=>"001001101",
  9873=>"100000111",
  9874=>"110111010",
  9875=>"011000101",
  9876=>"011010000",
  9877=>"011100110",
  9878=>"101111101",
  9879=>"101011001",
  9880=>"011110100",
  9881=>"000010110",
  9882=>"000100110",
  9883=>"000111100",
  9884=>"111011010",
  9885=>"110111011",
  9886=>"101010010",
  9887=>"001100110",
  9888=>"111010000",
  9889=>"101100110",
  9890=>"111000111",
  9891=>"010011011",
  9892=>"010011110",
  9893=>"001111101",
  9894=>"111101110",
  9895=>"111001010",
  9896=>"100010110",
  9897=>"110100110",
  9898=>"000110010",
  9899=>"011000001",
  9900=>"011000010",
  9901=>"110111010",
  9902=>"001111110",
  9903=>"011000001",
  9904=>"001110110",
  9905=>"011001000",
  9906=>"111111101",
  9907=>"001111000",
  9908=>"111100100",
  9909=>"010100101",
  9910=>"101001000",
  9911=>"100000100",
  9912=>"011101100",
  9913=>"110101001",
  9914=>"111010010",
  9915=>"110000110",
  9916=>"011010100",
  9917=>"111111111",
  9918=>"101010110",
  9919=>"111001111",
  9920=>"010101010",
  9921=>"100000100",
  9922=>"110111110",
  9923=>"111011000",
  9924=>"011010010",
  9925=>"010110101",
  9926=>"101100111",
  9927=>"010000000",
  9928=>"010101000",
  9929=>"111000000",
  9930=>"010000111",
  9931=>"000011010",
  9932=>"000010001",
  9933=>"011101011",
  9934=>"001110110",
  9935=>"100000011",
  9936=>"000001001",
  9937=>"100100001",
  9938=>"101010010",
  9939=>"001011001",
  9940=>"000110001",
  9941=>"110010011",
  9942=>"011001111",
  9943=>"001001001",
  9944=>"101111101",
  9945=>"100110001",
  9946=>"010100111",
  9947=>"011101001",
  9948=>"001101111",
  9949=>"101101000",
  9950=>"001000011",
  9951=>"001101111",
  9952=>"110001011",
  9953=>"100100111",
  9954=>"111101111",
  9955=>"101011101",
  9956=>"001011000",
  9957=>"111010110",
  9958=>"000010000",
  9959=>"011001000",
  9960=>"000100110",
  9961=>"101010011",
  9962=>"111011110",
  9963=>"111010101",
  9964=>"010000011",
  9965=>"100010101",
  9966=>"011111011",
  9967=>"111011001",
  9968=>"000100100",
  9969=>"100110000",
  9970=>"000111011",
  9971=>"001001001",
  9972=>"110000100",
  9973=>"100001000",
  9974=>"000110011",
  9975=>"100101000",
  9976=>"110110100",
  9977=>"110111000",
  9978=>"001000000",
  9979=>"100000010",
  9980=>"011101000",
  9981=>"111101100",
  9982=>"011011110",
  9983=>"011001000",
  9984=>"101010110",
  9985=>"001110011",
  9986=>"100100101",
  9987=>"110000000",
  9988=>"101100101",
  9989=>"101100111",
  9990=>"010110011",
  9991=>"100110101",
  9992=>"001001011",
  9993=>"111011100",
  9994=>"111001000",
  9995=>"101011000",
  9996=>"111101110",
  9997=>"001011001",
  9998=>"010001000",
  9999=>"111011101",
  10000=>"100110100",
  10001=>"111111100",
  10002=>"000001000",
  10003=>"100010010",
  10004=>"110001001",
  10005=>"001010110",
  10006=>"111101010",
  10007=>"110101001",
  10008=>"101001001",
  10009=>"011101000",
  10010=>"000110101",
  10011=>"000101110",
  10012=>"111010011",
  10013=>"001111111",
  10014=>"100101101",
  10015=>"101110110",
  10016=>"000110100",
  10017=>"111011011",
  10018=>"110100101",
  10019=>"101011001",
  10020=>"001010111",
  10021=>"101101011",
  10022=>"000001100",
  10023=>"101011100",
  10024=>"100110100",
  10025=>"100100001",
  10026=>"010011001",
  10027=>"110111110",
  10028=>"001110110",
  10029=>"000011010",
  10030=>"110110101",
  10031=>"010110010",
  10032=>"000110001",
  10033=>"101011101",
  10034=>"001000010",
  10035=>"111100101",
  10036=>"011001100",
  10037=>"010100111",
  10038=>"010000001",
  10039=>"001011011",
  10040=>"110101101",
  10041=>"010101010",
  10042=>"001001010",
  10043=>"110001001",
  10044=>"011101101",
  10045=>"100101000",
  10046=>"001101010",
  10047=>"110100000",
  10048=>"001011110",
  10049=>"101100000",
  10050=>"001001010",
  10051=>"100010101",
  10052=>"001011000",
  10053=>"101101111",
  10054=>"101111110",
  10055=>"001011101",
  10056=>"001010000",
  10057=>"111000001",
  10058=>"111101001",
  10059=>"011000100",
  10060=>"111100110",
  10061=>"110111101",
  10062=>"111110101",
  10063=>"100010110",
  10064=>"001100101",
  10065=>"000111010",
  10066=>"101101111",
  10067=>"000101010",
  10068=>"111111000",
  10069=>"000101010",
  10070=>"001111101",
  10071=>"001000000",
  10072=>"111100010",
  10073=>"000010101",
  10074=>"101111000",
  10075=>"000100011",
  10076=>"000001000",
  10077=>"000000011",
  10078=>"111100010",
  10079=>"011110111",
  10080=>"111000001",
  10081=>"110100000",
  10082=>"101111111",
  10083=>"111100111",
  10084=>"001111101",
  10085=>"010100101",
  10086=>"111111100",
  10087=>"001101111",
  10088=>"111000111",
  10089=>"001101100",
  10090=>"101101000",
  10091=>"000000010",
  10092=>"000000100",
  10093=>"001111001",
  10094=>"100101110",
  10095=>"101010110",
  10096=>"110101010",
  10097=>"000011010",
  10098=>"111110111",
  10099=>"101001101",
  10100=>"001001011",
  10101=>"010010011",
  10102=>"001010111",
  10103=>"000001110",
  10104=>"101010110",
  10105=>"111110100",
  10106=>"110001100",
  10107=>"110001110",
  10108=>"111101101",
  10109=>"111110111",
  10110=>"011000010",
  10111=>"111110101",
  10112=>"001001110",
  10113=>"000100111",
  10114=>"110101001",
  10115=>"111010001",
  10116=>"100001100",
  10117=>"111011010",
  10118=>"000110001",
  10119=>"101001001",
  10120=>"100011110",
  10121=>"100000110",
  10122=>"000001010",
  10123=>"111111111",
  10124=>"110000011",
  10125=>"111111010",
  10126=>"101101000",
  10127=>"001111011",
  10128=>"101111011",
  10129=>"111011111",
  10130=>"101110110",
  10131=>"001010100",
  10132=>"011111011",
  10133=>"100110110",
  10134=>"101110101",
  10135=>"100111100",
  10136=>"011100110",
  10137=>"111100110",
  10138=>"111101100",
  10139=>"111100100",
  10140=>"100111101",
  10141=>"010001110",
  10142=>"110100101",
  10143=>"010110010",
  10144=>"111110001",
  10145=>"110000000",
  10146=>"101000010",
  10147=>"111001000",
  10148=>"100100101",
  10149=>"001000010",
  10150=>"101100100",
  10151=>"110000010",
  10152=>"010101110",
  10153=>"111000011",
  10154=>"101101100",
  10155=>"010010110",
  10156=>"111111111",
  10157=>"011111101",
  10158=>"000101111",
  10159=>"100000100",
  10160=>"000000111",
  10161=>"011010100",
  10162=>"100001100",
  10163=>"000111101",
  10164=>"111100110",
  10165=>"001111010",
  10166=>"111001101",
  10167=>"000110001",
  10168=>"110100001",
  10169=>"101101001",
  10170=>"010100110",
  10171=>"000100111",
  10172=>"011110010",
  10173=>"000000000",
  10174=>"010011101",
  10175=>"001101101",
  10176=>"000111011",
  10177=>"110001011",
  10178=>"001011111",
  10179=>"110101101",
  10180=>"000000100",
  10181=>"100011111",
  10182=>"110001111",
  10183=>"011110000",
  10184=>"111001000",
  10185=>"101001000",
  10186=>"101101100",
  10187=>"100000100",
  10188=>"100100100",
  10189=>"000001010",
  10190=>"010001010",
  10191=>"110111111",
  10192=>"000111001",
  10193=>"000001110",
  10194=>"001010110",
  10195=>"100110100",
  10196=>"010101011",
  10197=>"010011000",
  10198=>"111110100",
  10199=>"101110000",
  10200=>"010000110",
  10201=>"010000001",
  10202=>"110111101",
  10203=>"000101110",
  10204=>"011011000",
  10205=>"011101111",
  10206=>"011010111",
  10207=>"000100001",
  10208=>"110100010",
  10209=>"011111111",
  10210=>"001100010",
  10211=>"111010101",
  10212=>"101111111",
  10213=>"111101101",
  10214=>"101010101",
  10215=>"010100000",
  10216=>"000100001",
  10217=>"101101101",
  10218=>"101100111",
  10219=>"110000101",
  10220=>"000100101",
  10221=>"011110000",
  10222=>"110111101",
  10223=>"110001010",
  10224=>"100110011",
  10225=>"101111111",
  10226=>"001011001",
  10227=>"010011101",
  10228=>"110101111",
  10229=>"110010110",
  10230=>"111100011",
  10231=>"001110000",
  10232=>"100001000",
  10233=>"100010111",
  10234=>"110011111",
  10235=>"001000110",
  10236=>"001011100",
  10237=>"011001101",
  10238=>"101001001",
  10239=>"000100010",
  10240=>"011110110",
  10241=>"001111010",
  10242=>"001001101",
  10243=>"000101000",
  10244=>"011110011",
  10245=>"001001010",
  10246=>"101111001",
  10247=>"111010110",
  10248=>"100110011",
  10249=>"010111010",
  10250=>"010111011",
  10251=>"111111101",
  10252=>"011000010",
  10253=>"001001111",
  10254=>"110100011",
  10255=>"111101001",
  10256=>"101111001",
  10257=>"111010000",
  10258=>"110101101",
  10259=>"111001110",
  10260=>"101010110",
  10261=>"100111010",
  10262=>"110101101",
  10263=>"000001001",
  10264=>"011001101",
  10265=>"100111111",
  10266=>"110000011",
  10267=>"110001011",
  10268=>"111011111",
  10269=>"001000000",
  10270=>"110110100",
  10271=>"000001111",
  10272=>"111000010",
  10273=>"111011100",
  10274=>"101001100",
  10275=>"010100111",
  10276=>"100110101",
  10277=>"010110001",
  10278=>"100001100",
  10279=>"110010110",
  10280=>"100110100",
  10281=>"111100111",
  10282=>"011101110",
  10283=>"000000110",
  10284=>"011111001",
  10285=>"101010011",
  10286=>"100011001",
  10287=>"101011111",
  10288=>"001011001",
  10289=>"100001101",
  10290=>"010011011",
  10291=>"101011000",
  10292=>"001111001",
  10293=>"010000001",
  10294=>"010100010",
  10295=>"110011110",
  10296=>"110101001",
  10297=>"011110110",
  10298=>"000000101",
  10299=>"011001011",
  10300=>"011001111",
  10301=>"010110000",
  10302=>"011010101",
  10303=>"000100111",
  10304=>"000111111",
  10305=>"000111100",
  10306=>"110001100",
  10307=>"010010101",
  10308=>"000100110",
  10309=>"000100010",
  10310=>"011011000",
  10311=>"101101001",
  10312=>"001010111",
  10313=>"000010000",
  10314=>"010100001",
  10315=>"000010100",
  10316=>"100001011",
  10317=>"111000111",
  10318=>"000001000",
  10319=>"101100000",
  10320=>"110011011",
  10321=>"000000101",
  10322=>"110100010",
  10323=>"011110100",
  10324=>"111101110",
  10325=>"010000000",
  10326=>"010110011",
  10327=>"100011001",
  10328=>"001101011",
  10329=>"100100011",
  10330=>"000011001",
  10331=>"110111110",
  10332=>"011001100",
  10333=>"000110011",
  10334=>"110111011",
  10335=>"000110110",
  10336=>"001110111",
  10337=>"111110101",
  10338=>"011001011",
  10339=>"000101011",
  10340=>"000101010",
  10341=>"101110010",
  10342=>"011001111",
  10343=>"001101101",
  10344=>"011101011",
  10345=>"010010101",
  10346=>"101001001",
  10347=>"010001111",
  10348=>"111001101",
  10349=>"001110000",
  10350=>"101111111",
  10351=>"000011001",
  10352=>"110010010",
  10353=>"010101010",
  10354=>"101011101",
  10355=>"001111011",
  10356=>"001111100",
  10357=>"101100100",
  10358=>"000001111",
  10359=>"000110101",
  10360=>"110111001",
  10361=>"111101000",
  10362=>"100010111",
  10363=>"001001000",
  10364=>"101011000",
  10365=>"010111000",
  10366=>"010011001",
  10367=>"000100110",
  10368=>"011011100",
  10369=>"010100001",
  10370=>"111010100",
  10371=>"001000110",
  10372=>"001110011",
  10373=>"010001011",
  10374=>"010111111",
  10375=>"011000001",
  10376=>"101011111",
  10377=>"111010101",
  10378=>"001001111",
  10379=>"011111000",
  10380=>"010101011",
  10381=>"100100001",
  10382=>"010110001",
  10383=>"010101110",
  10384=>"101010100",
  10385=>"011011011",
  10386=>"101100100",
  10387=>"110010011",
  10388=>"011110100",
  10389=>"111101010",
  10390=>"110000011",
  10391=>"011000111",
  10392=>"010011000",
  10393=>"011001110",
  10394=>"011101110",
  10395=>"001110000",
  10396=>"000010001",
  10397=>"100100100",
  10398=>"010101010",
  10399=>"110111000",
  10400=>"101111110",
  10401=>"000110101",
  10402=>"010000100",
  10403=>"110010000",
  10404=>"000111111",
  10405=>"000011000",
  10406=>"101001100",
  10407=>"001110101",
  10408=>"100111011",
  10409=>"100010000",
  10410=>"111000001",
  10411=>"000100111",
  10412=>"110010000",
  10413=>"100100100",
  10414=>"001101100",
  10415=>"011001011",
  10416=>"001011111",
  10417=>"000011000",
  10418=>"000010011",
  10419=>"101101111",
  10420=>"110010110",
  10421=>"011010001",
  10422=>"000001110",
  10423=>"000001011",
  10424=>"100100100",
  10425=>"110000101",
  10426=>"001111110",
  10427=>"101110010",
  10428=>"111000101",
  10429=>"001110001",
  10430=>"000100000",
  10431=>"001110000",
  10432=>"111001010",
  10433=>"000011000",
  10434=>"110101101",
  10435=>"100101110",
  10436=>"011001100",
  10437=>"010000100",
  10438=>"010001110",
  10439=>"001001000",
  10440=>"110100010",
  10441=>"011101010",
  10442=>"111101101",
  10443=>"010010101",
  10444=>"111010001",
  10445=>"100100000",
  10446=>"011001010",
  10447=>"001010101",
  10448=>"100010010",
  10449=>"101110100",
  10450=>"111100000",
  10451=>"010011001",
  10452=>"010101101",
  10453=>"001100100",
  10454=>"000110000",
  10455=>"100010111",
  10456=>"100000011",
  10457=>"001010000",
  10458=>"110100010",
  10459=>"011011000",
  10460=>"111111101",
  10461=>"101010111",
  10462=>"001011101",
  10463=>"111100001",
  10464=>"011000110",
  10465=>"001101111",
  10466=>"010101001",
  10467=>"010001011",
  10468=>"111111110",
  10469=>"000001000",
  10470=>"111101110",
  10471=>"110001111",
  10472=>"101011011",
  10473=>"001101011",
  10474=>"010100100",
  10475=>"101011010",
  10476=>"000100100",
  10477=>"010011000",
  10478=>"110010100",
  10479=>"001000000",
  10480=>"010110110",
  10481=>"100101000",
  10482=>"000110101",
  10483=>"110001011",
  10484=>"011000100",
  10485=>"010001000",
  10486=>"101101111",
  10487=>"010010101",
  10488=>"111100001",
  10489=>"110000011",
  10490=>"100010101",
  10491=>"110010100",
  10492=>"111011100",
  10493=>"001110000",
  10494=>"000011011",
  10495=>"010100111",
  10496=>"100110100",
  10497=>"101111010",
  10498=>"000110001",
  10499=>"001001010",
  10500=>"111111001",
  10501=>"011100101",
  10502=>"000011111",
  10503=>"101100001",
  10504=>"010011100",
  10505=>"101111011",
  10506=>"000110111",
  10507=>"110101011",
  10508=>"111011010",
  10509=>"011111011",
  10510=>"100100100",
  10511=>"101000100",
  10512=>"011111011",
  10513=>"000111000",
  10514=>"000111011",
  10515=>"011101110",
  10516=>"110000100",
  10517=>"100011101",
  10518=>"101010010",
  10519=>"101011001",
  10520=>"101010001",
  10521=>"111100010",
  10522=>"001101101",
  10523=>"010100110",
  10524=>"000100110",
  10525=>"010000110",
  10526=>"101101101",
  10527=>"100001001",
  10528=>"000100100",
  10529=>"111101101",
  10530=>"011111010",
  10531=>"000100000",
  10532=>"111101001",
  10533=>"111001001",
  10534=>"001011000",
  10535=>"000110110",
  10536=>"011011111",
  10537=>"100100000",
  10538=>"000111000",
  10539=>"100111111",
  10540=>"000000011",
  10541=>"111110111",
  10542=>"010111111",
  10543=>"100011110",
  10544=>"010100110",
  10545=>"101110110",
  10546=>"010010110",
  10547=>"011010010",
  10548=>"101100111",
  10549=>"111110001",
  10550=>"110100011",
  10551=>"100111110",
  10552=>"101000000",
  10553=>"001100001",
  10554=>"000000110",
  10555=>"110001011",
  10556=>"110000111",
  10557=>"000111001",
  10558=>"110011010",
  10559=>"010011011",
  10560=>"011011011",
  10561=>"100011111",
  10562=>"000100100",
  10563=>"101110010",
  10564=>"000110101",
  10565=>"010001001",
  10566=>"011110001",
  10567=>"101111110",
  10568=>"001100010",
  10569=>"111111000",
  10570=>"100001110",
  10571=>"011111010",
  10572=>"000101110",
  10573=>"010011011",
  10574=>"111001011",
  10575=>"101001011",
  10576=>"000100001",
  10577=>"111100010",
  10578=>"010110011",
  10579=>"101101111",
  10580=>"010111000",
  10581=>"010111111",
  10582=>"000000110",
  10583=>"000010111",
  10584=>"010001100",
  10585=>"010110011",
  10586=>"010001000",
  10587=>"011001010",
  10588=>"100111111",
  10589=>"010100100",
  10590=>"111011101",
  10591=>"100101101",
  10592=>"100111010",
  10593=>"101110100",
  10594=>"010010100",
  10595=>"101100011",
  10596=>"110001000",
  10597=>"111110000",
  10598=>"001111011",
  10599=>"111010111",
  10600=>"011101000",
  10601=>"111110110",
  10602=>"011001011",
  10603=>"101000111",
  10604=>"001110111",
  10605=>"110101100",
  10606=>"111010100",
  10607=>"010101010",
  10608=>"110011010",
  10609=>"000001000",
  10610=>"000001111",
  10611=>"001101100",
  10612=>"010100101",
  10613=>"000000111",
  10614=>"011011001",
  10615=>"000010000",
  10616=>"011100010",
  10617=>"000011100",
  10618=>"111001111",
  10619=>"101001100",
  10620=>"101010010",
  10621=>"001011001",
  10622=>"000101001",
  10623=>"000010100",
  10624=>"111010100",
  10625=>"011001111",
  10626=>"000000000",
  10627=>"010111001",
  10628=>"110101101",
  10629=>"010010011",
  10630=>"011001111",
  10631=>"001110111",
  10632=>"000010000",
  10633=>"101011110",
  10634=>"000000100",
  10635=>"001100010",
  10636=>"110000000",
  10637=>"100000001",
  10638=>"101111001",
  10639=>"101010001",
  10640=>"000011001",
  10641=>"000011110",
  10642=>"001011101",
  10643=>"111011111",
  10644=>"001110100",
  10645=>"001001111",
  10646=>"101000010",
  10647=>"110010010",
  10648=>"111000010",
  10649=>"101000001",
  10650=>"111100110",
  10651=>"011001001",
  10652=>"010001011",
  10653=>"000011110",
  10654=>"001001001",
  10655=>"101100101",
  10656=>"111011110",
  10657=>"110100110",
  10658=>"111111000",
  10659=>"010000111",
  10660=>"111000000",
  10661=>"111011110",
  10662=>"110000101",
  10663=>"111100111",
  10664=>"010010010",
  10665=>"100000000",
  10666=>"000010101",
  10667=>"000100101",
  10668=>"100001000",
  10669=>"111001100",
  10670=>"101001101",
  10671=>"100010111",
  10672=>"000111010",
  10673=>"101001110",
  10674=>"110101111",
  10675=>"011001011",
  10676=>"110000111",
  10677=>"111100111",
  10678=>"111100000",
  10679=>"110011110",
  10680=>"111110010",
  10681=>"111110001",
  10682=>"100100111",
  10683=>"101011101",
  10684=>"001110111",
  10685=>"010101010",
  10686=>"011000001",
  10687=>"001010101",
  10688=>"010011011",
  10689=>"101101100",
  10690=>"010001110",
  10691=>"011111101",
  10692=>"001001010",
  10693=>"100110001",
  10694=>"100010000",
  10695=>"010001010",
  10696=>"011011100",
  10697=>"001100011",
  10698=>"111101000",
  10699=>"010000111",
  10700=>"101110100",
  10701=>"111001001",
  10702=>"010011100",
  10703=>"111000100",
  10704=>"001000011",
  10705=>"000001010",
  10706=>"010000101",
  10707=>"100001011",
  10708=>"110011110",
  10709=>"000001101",
  10710=>"000010101",
  10711=>"111000010",
  10712=>"110100100",
  10713=>"111011001",
  10714=>"110111001",
  10715=>"111010000",
  10716=>"100010110",
  10717=>"000000110",
  10718=>"000011111",
  10719=>"000010001",
  10720=>"111111001",
  10721=>"111001011",
  10722=>"001011011",
  10723=>"111111011",
  10724=>"001010110",
  10725=>"101100010",
  10726=>"010011001",
  10727=>"000010010",
  10728=>"011111110",
  10729=>"011101001",
  10730=>"111011001",
  10731=>"100110010",
  10732=>"011110101",
  10733=>"110001000",
  10734=>"110101111",
  10735=>"110110110",
  10736=>"111111101",
  10737=>"000101010",
  10738=>"100000100",
  10739=>"110010101",
  10740=>"101110100",
  10741=>"010000011",
  10742=>"100001101",
  10743=>"100010101",
  10744=>"100000011",
  10745=>"101101101",
  10746=>"111001011",
  10747=>"010001010",
  10748=>"101100010",
  10749=>"001001100",
  10750=>"110001110",
  10751=>"110110110",
  10752=>"110001111",
  10753=>"100111101",
  10754=>"100010011",
  10755=>"100010100",
  10756=>"010000001",
  10757=>"001010100",
  10758=>"001011101",
  10759=>"110010101",
  10760=>"111010000",
  10761=>"010100010",
  10762=>"100000011",
  10763=>"110011011",
  10764=>"001011101",
  10765=>"111000011",
  10766=>"100110111",
  10767=>"111001111",
  10768=>"011010111",
  10769=>"100011100",
  10770=>"110000010",
  10771=>"001111111",
  10772=>"100000010",
  10773=>"100100011",
  10774=>"111100111",
  10775=>"101001010",
  10776=>"110001101",
  10777=>"000110110",
  10778=>"110011111",
  10779=>"100001110",
  10780=>"000111001",
  10781=>"100011001",
  10782=>"001101110",
  10783=>"111111011",
  10784=>"001101011",
  10785=>"110001100",
  10786=>"110100001",
  10787=>"000100101",
  10788=>"101100111",
  10789=>"111101000",
  10790=>"111011110",
  10791=>"000010100",
  10792=>"000101100",
  10793=>"000100010",
  10794=>"001010010",
  10795=>"000001100",
  10796=>"100010101",
  10797=>"001000011",
  10798=>"000101010",
  10799=>"010011001",
  10800=>"101100001",
  10801=>"110111011",
  10802=>"101011000",
  10803=>"000100000",
  10804=>"111000100",
  10805=>"001100100",
  10806=>"000011100",
  10807=>"010110111",
  10808=>"110010110",
  10809=>"011010111",
  10810=>"010011110",
  10811=>"000110011",
  10812=>"011110110",
  10813=>"110011010",
  10814=>"000000100",
  10815=>"110100111",
  10816=>"011000001",
  10817=>"011110011",
  10818=>"100010110",
  10819=>"100001001",
  10820=>"110011111",
  10821=>"010100011",
  10822=>"001011100",
  10823=>"011100100",
  10824=>"001001000",
  10825=>"001011110",
  10826=>"111110101",
  10827=>"111000001",
  10828=>"101110111",
  10829=>"001100101",
  10830=>"101000111",
  10831=>"011010001",
  10832=>"001010100",
  10833=>"011110011",
  10834=>"110010000",
  10835=>"111100001",
  10836=>"001001101",
  10837=>"010100000",
  10838=>"100100110",
  10839=>"101010010",
  10840=>"010110000",
  10841=>"111100000",
  10842=>"100010001",
  10843=>"111110001",
  10844=>"001010111",
  10845=>"111000111",
  10846=>"010001110",
  10847=>"101010010",
  10848=>"001000011",
  10849=>"001101011",
  10850=>"100000100",
  10851=>"001011110",
  10852=>"011010111",
  10853=>"010011010",
  10854=>"010011101",
  10855=>"000110010",
  10856=>"110101001",
  10857=>"010010110",
  10858=>"110001110",
  10859=>"011101001",
  10860=>"010111011",
  10861=>"011001101",
  10862=>"001000011",
  10863=>"101000101",
  10864=>"101110011",
  10865=>"000100110",
  10866=>"101000111",
  10867=>"100100010",
  10868=>"110111101",
  10869=>"010000110",
  10870=>"010101100",
  10871=>"001000101",
  10872=>"011001001",
  10873=>"101101110",
  10874=>"100111101",
  10875=>"110110010",
  10876=>"000010111",
  10877=>"010101010",
  10878=>"001101001",
  10879=>"011011111",
  10880=>"001010111",
  10881=>"001000101",
  10882=>"001001110",
  10883=>"100111101",
  10884=>"110100100",
  10885=>"101111100",
  10886=>"010101100",
  10887=>"011110000",
  10888=>"111111011",
  10889=>"101100111",
  10890=>"110111000",
  10891=>"000000010",
  10892=>"100110011",
  10893=>"110100101",
  10894=>"110110111",
  10895=>"110110110",
  10896=>"010101100",
  10897=>"101100100",
  10898=>"001100110",
  10899=>"011111111",
  10900=>"100100001",
  10901=>"011010000",
  10902=>"101100000",
  10903=>"110101100",
  10904=>"000101101",
  10905=>"100000101",
  10906=>"110111110",
  10907=>"101100100",
  10908=>"101000001",
  10909=>"101110100",
  10910=>"101010011",
  10911=>"010000100",
  10912=>"011111100",
  10913=>"010010010",
  10914=>"110000101",
  10915=>"101001100",
  10916=>"010010100",
  10917=>"011101111",
  10918=>"000100101",
  10919=>"000001111",
  10920=>"000000010",
  10921=>"011110010",
  10922=>"000010001",
  10923=>"111111101",
  10924=>"101001001",
  10925=>"010011101",
  10926=>"100010101",
  10927=>"001011010",
  10928=>"110001101",
  10929=>"010100011",
  10930=>"111000101",
  10931=>"101101111",
  10932=>"000001010",
  10933=>"000010000",
  10934=>"010011101",
  10935=>"100010001",
  10936=>"001111111",
  10937=>"101101000",
  10938=>"101111101",
  10939=>"010101010",
  10940=>"010000011",
  10941=>"011011101",
  10942=>"101101011",
  10943=>"110111010",
  10944=>"000101111",
  10945=>"011110101",
  10946=>"000100110",
  10947=>"101001000",
  10948=>"011100101",
  10949=>"010101010",
  10950=>"000000001",
  10951=>"001000101",
  10952=>"010010110",
  10953=>"111100100",
  10954=>"100001110",
  10955=>"010000000",
  10956=>"011111001",
  10957=>"100111001",
  10958=>"110100010",
  10959=>"000110100",
  10960=>"010000110",
  10961=>"110010001",
  10962=>"110101010",
  10963=>"000010100",
  10964=>"010010111",
  10965=>"010101000",
  10966=>"101111001",
  10967=>"001111100",
  10968=>"110011110",
  10969=>"000000010",
  10970=>"101101100",
  10971=>"010010111",
  10972=>"000101111",
  10973=>"011001100",
  10974=>"111110001",
  10975=>"001010111",
  10976=>"000000000",
  10977=>"001110011",
  10978=>"001001011",
  10979=>"101010100",
  10980=>"011111101",
  10981=>"000110111",
  10982=>"001111101",
  10983=>"100101110",
  10984=>"010110010",
  10985=>"101100000",
  10986=>"111111111",
  10987=>"001000101",
  10988=>"000011001",
  10989=>"000001111",
  10990=>"110000111",
  10991=>"001111101",
  10992=>"001010000",
  10993=>"000110000",
  10994=>"100001010",
  10995=>"110101110",
  10996=>"111001001",
  10997=>"001111100",
  10998=>"101101010",
  10999=>"111001001",
  11000=>"100100011",
  11001=>"001011010",
  11002=>"010011100",
  11003=>"000100110",
  11004=>"111000000",
  11005=>"111001011",
  11006=>"110100001",
  11007=>"010010000",
  11008=>"000101100",
  11009=>"111100100",
  11010=>"001110101",
  11011=>"001010110",
  11012=>"001000011",
  11013=>"001101100",
  11014=>"000101101",
  11015=>"110011101",
  11016=>"100000011",
  11017=>"111001101",
  11018=>"010011111",
  11019=>"000101011",
  11020=>"001010010",
  11021=>"011000001",
  11022=>"110011011",
  11023=>"011001111",
  11024=>"010110010",
  11025=>"010111001",
  11026=>"001000100",
  11027=>"001101000",
  11028=>"100100001",
  11029=>"000110111",
  11030=>"000110111",
  11031=>"101000010",
  11032=>"011011011",
  11033=>"000011011",
  11034=>"111110100",
  11035=>"111011001",
  11036=>"010100000",
  11037=>"111000001",
  11038=>"011010011",
  11039=>"100001101",
  11040=>"010001111",
  11041=>"010100101",
  11042=>"101110101",
  11043=>"000010000",
  11044=>"011001001",
  11045=>"010000000",
  11046=>"010100110",
  11047=>"100110111",
  11048=>"001000011",
  11049=>"101101001",
  11050=>"001110101",
  11051=>"001110011",
  11052=>"101011010",
  11053=>"110101110",
  11054=>"001001000",
  11055=>"010000110",
  11056=>"011000111",
  11057=>"001010100",
  11058=>"101010111",
  11059=>"010011000",
  11060=>"110010110",
  11061=>"011011110",
  11062=>"000100110",
  11063=>"110101011",
  11064=>"010110001",
  11065=>"011100111",
  11066=>"010000011",
  11067=>"011110010",
  11068=>"110001011",
  11069=>"111011101",
  11070=>"111111000",
  11071=>"010001010",
  11072=>"011011011",
  11073=>"101001111",
  11074=>"110001010",
  11075=>"001001010",
  11076=>"111010110",
  11077=>"111101100",
  11078=>"101111010",
  11079=>"001011100",
  11080=>"101011011",
  11081=>"001010101",
  11082=>"111101101",
  11083=>"100100100",
  11084=>"001111011",
  11085=>"110110000",
  11086=>"111001111",
  11087=>"110111100",
  11088=>"010101000",
  11089=>"011010110",
  11090=>"010001001",
  11091=>"111001101",
  11092=>"001101110",
  11093=>"000001110",
  11094=>"111011011",
  11095=>"100000000",
  11096=>"110001110",
  11097=>"001111010",
  11098=>"100110101",
  11099=>"110010110",
  11100=>"001011000",
  11101=>"100100010",
  11102=>"001000100",
  11103=>"100011110",
  11104=>"111010111",
  11105=>"011101011",
  11106=>"110011011",
  11107=>"111011110",
  11108=>"011100011",
  11109=>"011000001",
  11110=>"010001110",
  11111=>"100111001",
  11112=>"011010111",
  11113=>"000000001",
  11114=>"100111001",
  11115=>"100110101",
  11116=>"111000111",
  11117=>"000011110",
  11118=>"010011101",
  11119=>"011010011",
  11120=>"010111111",
  11121=>"001110010",
  11122=>"001011000",
  11123=>"000001101",
  11124=>"000111000",
  11125=>"100101111",
  11126=>"010101101",
  11127=>"011101011",
  11128=>"011011110",
  11129=>"011100111",
  11130=>"101001000",
  11131=>"111011000",
  11132=>"010001010",
  11133=>"111001000",
  11134=>"001100110",
  11135=>"010010101",
  11136=>"010110000",
  11137=>"101000011",
  11138=>"001100010",
  11139=>"000110000",
  11140=>"000000000",
  11141=>"111000101",
  11142=>"000011110",
  11143=>"010011000",
  11144=>"111101011",
  11145=>"100000111",
  11146=>"001010110",
  11147=>"100010011",
  11148=>"100110101",
  11149=>"110111000",
  11150=>"000001101",
  11151=>"100110110",
  11152=>"000001111",
  11153=>"001100110",
  11154=>"111001010",
  11155=>"100110110",
  11156=>"000100111",
  11157=>"110100001",
  11158=>"100011100",
  11159=>"111001001",
  11160=>"111011011",
  11161=>"100001111",
  11162=>"001011000",
  11163=>"111101100",
  11164=>"000010000",
  11165=>"010000010",
  11166=>"010001100",
  11167=>"111111101",
  11168=>"011111101",
  11169=>"100111000",
  11170=>"000011111",
  11171=>"000111010",
  11172=>"000101101",
  11173=>"001000110",
  11174=>"101110111",
  11175=>"000101101",
  11176=>"110001010",
  11177=>"000010001",
  11178=>"000111001",
  11179=>"101110101",
  11180=>"111101101",
  11181=>"000010111",
  11182=>"010110110",
  11183=>"000111000",
  11184=>"100101100",
  11185=>"111111111",
  11186=>"001010110",
  11187=>"010010101",
  11188=>"110110111",
  11189=>"011110101",
  11190=>"011000110",
  11191=>"011001011",
  11192=>"010000001",
  11193=>"011011111",
  11194=>"010111111",
  11195=>"001100010",
  11196=>"000010000",
  11197=>"100000110",
  11198=>"101111110",
  11199=>"110000101",
  11200=>"100110111",
  11201=>"010101110",
  11202=>"101110000",
  11203=>"111000001",
  11204=>"100000100",
  11205=>"110001101",
  11206=>"011100010",
  11207=>"011011010",
  11208=>"110101010",
  11209=>"000101111",
  11210=>"110000101",
  11211=>"110100010",
  11212=>"111001111",
  11213=>"010000010",
  11214=>"000110000",
  11215=>"010110011",
  11216=>"100101001",
  11217=>"010100010",
  11218=>"101001000",
  11219=>"111111000",
  11220=>"101010010",
  11221=>"100010011",
  11222=>"001010010",
  11223=>"000001111",
  11224=>"101001011",
  11225=>"011001011",
  11226=>"010011100",
  11227=>"110010000",
  11228=>"001110101",
  11229=>"100000011",
  11230=>"101101111",
  11231=>"101101001",
  11232=>"111000110",
  11233=>"010111011",
  11234=>"111001110",
  11235=>"110101110",
  11236=>"010110111",
  11237=>"011000000",
  11238=>"001010001",
  11239=>"011001100",
  11240=>"101000011",
  11241=>"001000001",
  11242=>"001000111",
  11243=>"001011100",
  11244=>"000100110",
  11245=>"110001010",
  11246=>"101110010",
  11247=>"111011111",
  11248=>"100001111",
  11249=>"100101111",
  11250=>"010011101",
  11251=>"111000110",
  11252=>"010010110",
  11253=>"111101000",
  11254=>"110111100",
  11255=>"110000001",
  11256=>"000111110",
  11257=>"111010110",
  11258=>"000110010",
  11259=>"000111001",
  11260=>"111010110",
  11261=>"001011111",
  11262=>"101001101",
  11263=>"000101010",
  11264=>"000111010",
  11265=>"110000101",
  11266=>"011001010",
  11267=>"111011000",
  11268=>"111010111",
  11269=>"000000100",
  11270=>"110100010",
  11271=>"011111011",
  11272=>"111111010",
  11273=>"011110011",
  11274=>"010101000",
  11275=>"111101010",
  11276=>"101010110",
  11277=>"001101101",
  11278=>"100001110",
  11279=>"111011100",
  11280=>"010010111",
  11281=>"000001001",
  11282=>"100010100",
  11283=>"000010010",
  11284=>"111100011",
  11285=>"101110010",
  11286=>"100111001",
  11287=>"011010000",
  11288=>"001100110",
  11289=>"111000000",
  11290=>"010111100",
  11291=>"001011001",
  11292=>"100000101",
  11293=>"000011111",
  11294=>"111000110",
  11295=>"111111011",
  11296=>"111010100",
  11297=>"101010010",
  11298=>"011111010",
  11299=>"100011001",
  11300=>"000110011",
  11301=>"101000011",
  11302=>"100010010",
  11303=>"001101100",
  11304=>"110100011",
  11305=>"011010111",
  11306=>"001101000",
  11307=>"111010111",
  11308=>"000111101",
  11309=>"101101100",
  11310=>"000101111",
  11311=>"100001100",
  11312=>"011111001",
  11313=>"010010111",
  11314=>"010010011",
  11315=>"001011110",
  11316=>"000000111",
  11317=>"100010111",
  11318=>"101001000",
  11319=>"001010101",
  11320=>"000010111",
  11321=>"101101010",
  11322=>"101100111",
  11323=>"100011001",
  11324=>"111101000",
  11325=>"011001110",
  11326=>"011110100",
  11327=>"011001010",
  11328=>"000000000",
  11329=>"100000001",
  11330=>"100011001",
  11331=>"111111101",
  11332=>"100100001",
  11333=>"001000000",
  11334=>"110101001",
  11335=>"111111111",
  11336=>"010101111",
  11337=>"110110000",
  11338=>"110010101",
  11339=>"100100011",
  11340=>"101001101",
  11341=>"110000001",
  11342=>"100000000",
  11343=>"000001011",
  11344=>"110100110",
  11345=>"101110110",
  11346=>"100010011",
  11347=>"100111010",
  11348=>"000100111",
  11349=>"111100011",
  11350=>"101111111",
  11351=>"111101111",
  11352=>"011001100",
  11353=>"101101111",
  11354=>"111101101",
  11355=>"101110110",
  11356=>"000011111",
  11357=>"100100111",
  11358=>"110000011",
  11359=>"000000010",
  11360=>"101110000",
  11361=>"111000101",
  11362=>"101010000",
  11363=>"101100001",
  11364=>"110001011",
  11365=>"001000010",
  11366=>"010101101",
  11367=>"110111111",
  11368=>"011101111",
  11369=>"011000111",
  11370=>"010011001",
  11371=>"110100000",
  11372=>"001001111",
  11373=>"100100100",
  11374=>"110000001",
  11375=>"110110001",
  11376=>"010011110",
  11377=>"100000010",
  11378=>"001000011",
  11379=>"101101011",
  11380=>"100100101",
  11381=>"110001111",
  11382=>"101101111",
  11383=>"010111011",
  11384=>"100011010",
  11385=>"011000110",
  11386=>"001011110",
  11387=>"010000010",
  11388=>"101100101",
  11389=>"101000001",
  11390=>"101000001",
  11391=>"110101100",
  11392=>"000001001",
  11393=>"000001011",
  11394=>"001000101",
  11395=>"000111001",
  11396=>"100100011",
  11397=>"110100011",
  11398=>"111100010",
  11399=>"100000100",
  11400=>"100101001",
  11401=>"010111100",
  11402=>"100010000",
  11403=>"010001000",
  11404=>"110010011",
  11405=>"100100101",
  11406=>"001101011",
  11407=>"111000100",
  11408=>"011101010",
  11409=>"101101111",
  11410=>"011110101",
  11411=>"111101101",
  11412=>"000000000",
  11413=>"101111001",
  11414=>"011101101",
  11415=>"001010101",
  11416=>"111100011",
  11417=>"001100101",
  11418=>"100011010",
  11419=>"011000100",
  11420=>"110000010",
  11421=>"111101001",
  11422=>"000100010",
  11423=>"101100011",
  11424=>"110110000",
  11425=>"001111011",
  11426=>"110111011",
  11427=>"010010101",
  11428=>"001000001",
  11429=>"000100111",
  11430=>"100000101",
  11431=>"100100101",
  11432=>"111010100",
  11433=>"001011110",
  11434=>"010010001",
  11435=>"111010000",
  11436=>"100000111",
  11437=>"101111011",
  11438=>"100010001",
  11439=>"100101001",
  11440=>"000011010",
  11441=>"011010100",
  11442=>"101110010",
  11443=>"011001000",
  11444=>"110001011",
  11445=>"111011101",
  11446=>"100010100",
  11447=>"101001010",
  11448=>"010111110",
  11449=>"111010110",
  11450=>"110000111",
  11451=>"000100001",
  11452=>"111011011",
  11453=>"010110101",
  11454=>"000110011",
  11455=>"110111000",
  11456=>"100011000",
  11457=>"011011111",
  11458=>"000111101",
  11459=>"111000001",
  11460=>"011001100",
  11461=>"011111010",
  11462=>"011110111",
  11463=>"001001011",
  11464=>"111111111",
  11465=>"110111110",
  11466=>"110010010",
  11467=>"100101110",
  11468=>"000111110",
  11469=>"101001000",
  11470=>"000001011",
  11471=>"000010000",
  11472=>"010101111",
  11473=>"010101001",
  11474=>"101010011",
  11475=>"100011010",
  11476=>"001110010",
  11477=>"110111010",
  11478=>"000011010",
  11479=>"001000001",
  11480=>"001000111",
  11481=>"000001010",
  11482=>"101010000",
  11483=>"000010111",
  11484=>"110110011",
  11485=>"001010001",
  11486=>"000011110",
  11487=>"000101110",
  11488=>"111001001",
  11489=>"000000100",
  11490=>"001100111",
  11491=>"010001111",
  11492=>"100110110",
  11493=>"111111111",
  11494=>"011111111",
  11495=>"010110001",
  11496=>"000011110",
  11497=>"111111001",
  11498=>"011011010",
  11499=>"111010110",
  11500=>"011100010",
  11501=>"000001100",
  11502=>"110111101",
  11503=>"100110111",
  11504=>"000010011",
  11505=>"011110101",
  11506=>"111000001",
  11507=>"100101010",
  11508=>"010111010",
  11509=>"110000010",
  11510=>"001111010",
  11511=>"100000010",
  11512=>"001010101",
  11513=>"011111011",
  11514=>"011011111",
  11515=>"000001001",
  11516=>"101000110",
  11517=>"110101101",
  11518=>"010011100",
  11519=>"000111111",
  11520=>"100010110",
  11521=>"100000110",
  11522=>"100111000",
  11523=>"110000010",
  11524=>"001111100",
  11525=>"011010001",
  11526=>"011011110",
  11527=>"010001011",
  11528=>"111001001",
  11529=>"000000010",
  11530=>"100001010",
  11531=>"010111000",
  11532=>"000010001",
  11533=>"001100101",
  11534=>"111001011",
  11535=>"000000111",
  11536=>"001011110",
  11537=>"000000100",
  11538=>"000001110",
  11539=>"110111000",
  11540=>"001100100",
  11541=>"001010011",
  11542=>"010111011",
  11543=>"111101011",
  11544=>"010010100",
  11545=>"110100111",
  11546=>"100010100",
  11547=>"110110111",
  11548=>"000101111",
  11549=>"100100000",
  11550=>"001111000",
  11551=>"011010000",
  11552=>"100100000",
  11553=>"001011001",
  11554=>"100110110",
  11555=>"111010010",
  11556=>"110000000",
  11557=>"100001101",
  11558=>"010000110",
  11559=>"100011100",
  11560=>"000001110",
  11561=>"110010110",
  11562=>"010110110",
  11563=>"101110010",
  11564=>"010001111",
  11565=>"101111101",
  11566=>"011000001",
  11567=>"011111000",
  11568=>"111101110",
  11569=>"110110001",
  11570=>"010011110",
  11571=>"111110001",
  11572=>"111111001",
  11573=>"001000100",
  11574=>"010001100",
  11575=>"001110010",
  11576=>"001110101",
  11577=>"011011101",
  11578=>"001100011",
  11579=>"101001100",
  11580=>"001110001",
  11581=>"111101110",
  11582=>"100100000",
  11583=>"000000011",
  11584=>"010100100",
  11585=>"110101111",
  11586=>"000000110",
  11587=>"101101101",
  11588=>"010011111",
  11589=>"001101110",
  11590=>"100000110",
  11591=>"110110101",
  11592=>"010011110",
  11593=>"110011011",
  11594=>"011100010",
  11595=>"001010100",
  11596=>"110001100",
  11597=>"010011010",
  11598=>"011100001",
  11599=>"100001000",
  11600=>"011011011",
  11601=>"010000000",
  11602=>"110100001",
  11603=>"110011010",
  11604=>"001011000",
  11605=>"000001010",
  11606=>"110010011",
  11607=>"001110011",
  11608=>"000011101",
  11609=>"001000000",
  11610=>"010101010",
  11611=>"100100110",
  11612=>"000010000",
  11613=>"111111101",
  11614=>"001111110",
  11615=>"000001001",
  11616=>"110001010",
  11617=>"011001111",
  11618=>"111001111",
  11619=>"110011011",
  11620=>"111000101",
  11621=>"110100010",
  11622=>"001011111",
  11623=>"000010010",
  11624=>"010010101",
  11625=>"000000000",
  11626=>"000110010",
  11627=>"000010011",
  11628=>"010011000",
  11629=>"011101100",
  11630=>"000000110",
  11631=>"111101110",
  11632=>"010010000",
  11633=>"001011100",
  11634=>"101101100",
  11635=>"011101001",
  11636=>"100011011",
  11637=>"111010100",
  11638=>"100010101",
  11639=>"010001010",
  11640=>"110011110",
  11641=>"010101110",
  11642=>"101011011",
  11643=>"110110111",
  11644=>"010111110",
  11645=>"101110111",
  11646=>"101111111",
  11647=>"100110100",
  11648=>"001001001",
  11649=>"011111111",
  11650=>"010111011",
  11651=>"011011100",
  11652=>"100000001",
  11653=>"100111101",
  11654=>"101100111",
  11655=>"100101010",
  11656=>"111010001",
  11657=>"000100001",
  11658=>"000011101",
  11659=>"010000100",
  11660=>"110101100",
  11661=>"101011100",
  11662=>"000101010",
  11663=>"111000110",
  11664=>"000101011",
  11665=>"000100100",
  11666=>"110101010",
  11667=>"101111000",
  11668=>"011111011",
  11669=>"011111100",
  11670=>"111110111",
  11671=>"110111011",
  11672=>"110000111",
  11673=>"010010010",
  11674=>"001011001",
  11675=>"100000100",
  11676=>"100101100",
  11677=>"110000001",
  11678=>"011100010",
  11679=>"011111000",
  11680=>"111101101",
  11681=>"100001000",
  11682=>"001000011",
  11683=>"000010011",
  11684=>"110100100",
  11685=>"101111101",
  11686=>"011011001",
  11687=>"000010011",
  11688=>"101100001",
  11689=>"110111111",
  11690=>"000011011",
  11691=>"101011011",
  11692=>"000011010",
  11693=>"101011110",
  11694=>"011101111",
  11695=>"111101101",
  11696=>"111101000",
  11697=>"111101110",
  11698=>"010010100",
  11699=>"111001100",
  11700=>"010010011",
  11701=>"101111100",
  11702=>"100010101",
  11703=>"111111000",
  11704=>"101011111",
  11705=>"011011110",
  11706=>"111010010",
  11707=>"110100110",
  11708=>"100011100",
  11709=>"010000101",
  11710=>"101111111",
  11711=>"000111100",
  11712=>"010100111",
  11713=>"001111111",
  11714=>"011010001",
  11715=>"101001000",
  11716=>"101011111",
  11717=>"110111001",
  11718=>"100100011",
  11719=>"001000010",
  11720=>"110111111",
  11721=>"101010101",
  11722=>"110000010",
  11723=>"110011001",
  11724=>"010001110",
  11725=>"011101111",
  11726=>"000010001",
  11727=>"011111010",
  11728=>"110011100",
  11729=>"001101001",
  11730=>"001011100",
  11731=>"100001000",
  11732=>"100000001",
  11733=>"010011011",
  11734=>"011110000",
  11735=>"011100000",
  11736=>"111100100",
  11737=>"100001010",
  11738=>"100000000",
  11739=>"001111000",
  11740=>"100111001",
  11741=>"111001010",
  11742=>"100111100",
  11743=>"110110100",
  11744=>"111000001",
  11745=>"001001000",
  11746=>"111100011",
  11747=>"010111000",
  11748=>"000011110",
  11749=>"100001100",
  11750=>"100111001",
  11751=>"101010101",
  11752=>"101111111",
  11753=>"111110101",
  11754=>"101000000",
  11755=>"001111010",
  11756=>"000011001",
  11757=>"001110100",
  11758=>"001001101",
  11759=>"001111111",
  11760=>"001001001",
  11761=>"010011101",
  11762=>"000001100",
  11763=>"110000100",
  11764=>"111001111",
  11765=>"010010001",
  11766=>"101010011",
  11767=>"010100110",
  11768=>"011011010",
  11769=>"000111100",
  11770=>"000010011",
  11771=>"001110110",
  11772=>"011100101",
  11773=>"000011100",
  11774=>"010100000",
  11775=>"010010100",
  11776=>"100110101",
  11777=>"001100111",
  11778=>"001000100",
  11779=>"001110011",
  11780=>"000010000",
  11781=>"100010100",
  11782=>"110101101",
  11783=>"100110110",
  11784=>"111010001",
  11785=>"000110011",
  11786=>"001100100",
  11787=>"010010000",
  11788=>"000011010",
  11789=>"101000111",
  11790=>"011001010",
  11791=>"101110011",
  11792=>"101011011",
  11793=>"011101101",
  11794=>"111010101",
  11795=>"111100110",
  11796=>"110110010",
  11797=>"110100001",
  11798=>"111010000",
  11799=>"101110000",
  11800=>"000001110",
  11801=>"001110100",
  11802=>"011011011",
  11803=>"010111001",
  11804=>"010010110",
  11805=>"011010111",
  11806=>"011101000",
  11807=>"010110010",
  11808=>"111110011",
  11809=>"011100101",
  11810=>"001100000",
  11811=>"010011010",
  11812=>"111000100",
  11813=>"000011000",
  11814=>"110111000",
  11815=>"000110000",
  11816=>"011001100",
  11817=>"001110100",
  11818=>"010110110",
  11819=>"000100010",
  11820=>"011101101",
  11821=>"001011001",
  11822=>"100000111",
  11823=>"101011101",
  11824=>"100101010",
  11825=>"111100110",
  11826=>"000101100",
  11827=>"000101000",
  11828=>"000000011",
  11829=>"010110010",
  11830=>"101111110",
  11831=>"011010100",
  11832=>"000111100",
  11833=>"000101000",
  11834=>"011010010",
  11835=>"101101111",
  11836=>"011000010",
  11837=>"100010110",
  11838=>"001111010",
  11839=>"010101101",
  11840=>"101001100",
  11841=>"111100011",
  11842=>"010011011",
  11843=>"011010110",
  11844=>"101111001",
  11845=>"010010010",
  11846=>"001101100",
  11847=>"010110110",
  11848=>"001110011",
  11849=>"001001011",
  11850=>"110011000",
  11851=>"010110001",
  11852=>"010010100",
  11853=>"111100100",
  11854=>"100111101",
  11855=>"000011111",
  11856=>"010110101",
  11857=>"110100100",
  11858=>"111110111",
  11859=>"110000101",
  11860=>"110100111",
  11861=>"000111011",
  11862=>"011000110",
  11863=>"000000010",
  11864=>"100011101",
  11865=>"001011111",
  11866=>"011000101",
  11867=>"001000101",
  11868=>"000001110",
  11869=>"110010010",
  11870=>"110011010",
  11871=>"000111010",
  11872=>"011000111",
  11873=>"000010110",
  11874=>"101000101",
  11875=>"001000011",
  11876=>"111011110",
  11877=>"001010001",
  11878=>"101000101",
  11879=>"001110000",
  11880=>"110001110",
  11881=>"001111100",
  11882=>"111001111",
  11883=>"001010000",
  11884=>"100001110",
  11885=>"010100010",
  11886=>"010110100",
  11887=>"010110011",
  11888=>"111100001",
  11889=>"011100100",
  11890=>"011010111",
  11891=>"101010111",
  11892=>"011101011",
  11893=>"011110010",
  11894=>"000000101",
  11895=>"111101111",
  11896=>"111100011",
  11897=>"111000001",
  11898=>"011111001",
  11899=>"011011111",
  11900=>"111101001",
  11901=>"110110100",
  11902=>"101010001",
  11903=>"110111100",
  11904=>"111111100",
  11905=>"110101000",
  11906=>"000000111",
  11907=>"000110111",
  11908=>"110100010",
  11909=>"101010010",
  11910=>"100010110",
  11911=>"010000101",
  11912=>"111011110",
  11913=>"101010000",
  11914=>"011111100",
  11915=>"000000001",
  11916=>"111011111",
  11917=>"011011001",
  11918=>"101101010",
  11919=>"110011111",
  11920=>"110110011",
  11921=>"011101000",
  11922=>"000010001",
  11923=>"001000111",
  11924=>"000000001",
  11925=>"011110000",
  11926=>"011001110",
  11927=>"011010101",
  11928=>"101000000",
  11929=>"111000111",
  11930=>"110110111",
  11931=>"101110000",
  11932=>"111011101",
  11933=>"010111000",
  11934=>"000001110",
  11935=>"010010010",
  11936=>"100100101",
  11937=>"000000011",
  11938=>"010110001",
  11939=>"100111000",
  11940=>"000011011",
  11941=>"101110100",
  11942=>"110101101",
  11943=>"111111011",
  11944=>"000000011",
  11945=>"000001100",
  11946=>"111011111",
  11947=>"110010000",
  11948=>"110100010",
  11949=>"010101001",
  11950=>"101101101",
  11951=>"010011010",
  11952=>"111010101",
  11953=>"110000000",
  11954=>"101001010",
  11955=>"001001011",
  11956=>"000011000",
  11957=>"011001111",
  11958=>"011101110",
  11959=>"111000100",
  11960=>"000111011",
  11961=>"110100001",
  11962=>"000010000",
  11963=>"011001011",
  11964=>"011000111",
  11965=>"101001110",
  11966=>"111010100",
  11967=>"110001101",
  11968=>"001110100",
  11969=>"100011101",
  11970=>"011100100",
  11971=>"001011011",
  11972=>"000110100",
  11973=>"100000100",
  11974=>"011000110",
  11975=>"101110100",
  11976=>"100100000",
  11977=>"001101010",
  11978=>"000100011",
  11979=>"100010110",
  11980=>"100111110",
  11981=>"011110111",
  11982=>"110111111",
  11983=>"000000011",
  11984=>"101001110",
  11985=>"000000010",
  11986=>"100001010",
  11987=>"000100101",
  11988=>"000111111",
  11989=>"110011010",
  11990=>"001000001",
  11991=>"101010111",
  11992=>"010110011",
  11993=>"011011000",
  11994=>"000101100",
  11995=>"100101110",
  11996=>"111110110",
  11997=>"001110011",
  11998=>"010010001",
  11999=>"010010011",
  12000=>"111101110",
  12001=>"100010010",
  12002=>"100000110",
  12003=>"010011001",
  12004=>"001101000",
  12005=>"110100101",
  12006=>"000111100",
  12007=>"001111001",
  12008=>"100010100",
  12009=>"001101011",
  12010=>"101000101",
  12011=>"000001111",
  12012=>"001000001",
  12013=>"100001010",
  12014=>"010000001",
  12015=>"101011000",
  12016=>"000001110",
  12017=>"110101101",
  12018=>"111100000",
  12019=>"101001111",
  12020=>"100110110",
  12021=>"100101101",
  12022=>"000101011",
  12023=>"010101101",
  12024=>"100011000",
  12025=>"011110111",
  12026=>"100000110",
  12027=>"011100011",
  12028=>"100101001",
  12029=>"111001011",
  12030=>"001010101",
  12031=>"101101000",
  12032=>"010100001",
  12033=>"010000100",
  12034=>"011010111",
  12035=>"111111010",
  12036=>"000110010",
  12037=>"100000111",
  12038=>"101010110",
  12039=>"110101010",
  12040=>"010010111",
  12041=>"100101101",
  12042=>"110100000",
  12043=>"100001011",
  12044=>"000001101",
  12045=>"010001000",
  12046=>"100101101",
  12047=>"111110101",
  12048=>"001011011",
  12049=>"100011101",
  12050=>"000011100",
  12051=>"111001100",
  12052=>"000000110",
  12053=>"000001101",
  12054=>"001011011",
  12055=>"101010101",
  12056=>"011000111",
  12057=>"100010010",
  12058=>"010010000",
  12059=>"110100101",
  12060=>"001110111",
  12061=>"100010001",
  12062=>"010010110",
  12063=>"011011110",
  12064=>"111101100",
  12065=>"101111111",
  12066=>"111111101",
  12067=>"010110000",
  12068=>"111010100",
  12069=>"011011011",
  12070=>"101001100",
  12071=>"011111010",
  12072=>"101101110",
  12073=>"101010111",
  12074=>"101000011",
  12075=>"101010010",
  12076=>"101011011",
  12077=>"111101101",
  12078=>"101001001",
  12079=>"101110111",
  12080=>"000000111",
  12081=>"111000111",
  12082=>"101110111",
  12083=>"111111000",
  12084=>"010101001",
  12085=>"001001000",
  12086=>"010011111",
  12087=>"101010001",
  12088=>"110101000",
  12089=>"100010011",
  12090=>"111011011",
  12091=>"100101110",
  12092=>"110111011",
  12093=>"101000001",
  12094=>"101101110",
  12095=>"111101110",
  12096=>"000011101",
  12097=>"100101111",
  12098=>"110111111",
  12099=>"101111111",
  12100=>"101000100",
  12101=>"010000001",
  12102=>"001101000",
  12103=>"000101100",
  12104=>"110000001",
  12105=>"000011000",
  12106=>"000101001",
  12107=>"010111111",
  12108=>"000111000",
  12109=>"011111110",
  12110=>"010100110",
  12111=>"101100100",
  12112=>"000110000",
  12113=>"111110001",
  12114=>"100111110",
  12115=>"110111111",
  12116=>"111110111",
  12117=>"010100110",
  12118=>"000101010",
  12119=>"000101010",
  12120=>"110111100",
  12121=>"010000101",
  12122=>"001101001",
  12123=>"111000011",
  12124=>"011011100",
  12125=>"000111001",
  12126=>"110011111",
  12127=>"000010001",
  12128=>"110010011",
  12129=>"001000011",
  12130=>"010001110",
  12131=>"000100011",
  12132=>"001011010",
  12133=>"000010100",
  12134=>"110011000",
  12135=>"000011011",
  12136=>"010000110",
  12137=>"101000001",
  12138=>"010001100",
  12139=>"100010101",
  12140=>"011111101",
  12141=>"010011011",
  12142=>"110011110",
  12143=>"100001011",
  12144=>"011010110",
  12145=>"111000001",
  12146=>"010001110",
  12147=>"101011000",
  12148=>"111000011",
  12149=>"101110101",
  12150=>"110111110",
  12151=>"010100010",
  12152=>"110100011",
  12153=>"010011000",
  12154=>"010100010",
  12155=>"011010011",
  12156=>"111100101",
  12157=>"010110010",
  12158=>"011001011",
  12159=>"011001110",
  12160=>"000010000",
  12161=>"011110001",
  12162=>"101010010",
  12163=>"111000101",
  12164=>"110101010",
  12165=>"101111110",
  12166=>"100000000",
  12167=>"011100110",
  12168=>"110010000",
  12169=>"001100100",
  12170=>"100011101",
  12171=>"101011000",
  12172=>"110100110",
  12173=>"110111110",
  12174=>"000101001",
  12175=>"111101001",
  12176=>"000100011",
  12177=>"111100010",
  12178=>"000110111",
  12179=>"011100111",
  12180=>"111100001",
  12181=>"011001000",
  12182=>"000001101",
  12183=>"111110110",
  12184=>"111000110",
  12185=>"101011001",
  12186=>"001000100",
  12187=>"111001111",
  12188=>"011001110",
  12189=>"101101111",
  12190=>"110011010",
  12191=>"111010101",
  12192=>"100011100",
  12193=>"110110101",
  12194=>"001010101",
  12195=>"001111001",
  12196=>"100010001",
  12197=>"000010110",
  12198=>"110100100",
  12199=>"111001010",
  12200=>"001010011",
  12201=>"111111011",
  12202=>"110011100",
  12203=>"101010111",
  12204=>"010110100",
  12205=>"111000010",
  12206=>"000001010",
  12207=>"011011111",
  12208=>"110000010",
  12209=>"100011100",
  12210=>"001111111",
  12211=>"111010111",
  12212=>"110111010",
  12213=>"101010001",
  12214=>"111000110",
  12215=>"101010110",
  12216=>"011111011",
  12217=>"011011100",
  12218=>"011011011",
  12219=>"010010001",
  12220=>"011001001",
  12221=>"100010110",
  12222=>"111011110",
  12223=>"101101111",
  12224=>"000011100",
  12225=>"010010011",
  12226=>"110100100",
  12227=>"110000010",
  12228=>"100110101",
  12229=>"011110111",
  12230=>"000110111",
  12231=>"001010110",
  12232=>"111010001",
  12233=>"101101000",
  12234=>"111101101",
  12235=>"111000100",
  12236=>"000110011",
  12237=>"101101101",
  12238=>"111111110",
  12239=>"001001000",
  12240=>"101100000",
  12241=>"010111100",
  12242=>"000101010",
  12243=>"000000010",
  12244=>"001101110",
  12245=>"010101011",
  12246=>"100100010",
  12247=>"110000100",
  12248=>"100111011",
  12249=>"010010011",
  12250=>"111100100",
  12251=>"101111000",
  12252=>"000001111",
  12253=>"000100111",
  12254=>"101011110",
  12255=>"100000000",
  12256=>"001101000",
  12257=>"001101000",
  12258=>"000011110",
  12259=>"001000110",
  12260=>"100111001",
  12261=>"000110110",
  12262=>"010010010",
  12263=>"010101001",
  12264=>"110110100",
  12265=>"010001000",
  12266=>"000101010",
  12267=>"001101110",
  12268=>"011011101",
  12269=>"110111110",
  12270=>"000100110",
  12271=>"010011001",
  12272=>"001010111",
  12273=>"000010111",
  12274=>"101010001",
  12275=>"000110110",
  12276=>"001000010",
  12277=>"101000101",
  12278=>"111110111",
  12279=>"111000011",
  12280=>"000100000",
  12281=>"101001000",
  12282=>"010010000",
  12283=>"001000111",
  12284=>"001010001",
  12285=>"011111101",
  12286=>"001000010",
  12287=>"101011001",
  12288=>"111011001",
  12289=>"001111000",
  12290=>"011110011",
  12291=>"011000011",
  12292=>"010110110",
  12293=>"010001010",
  12294=>"001010111",
  12295=>"100100101",
  12296=>"010000010",
  12297=>"011011110",
  12298=>"100110001",
  12299=>"000011011",
  12300=>"110110111",
  12301=>"110101000",
  12302=>"101000001",
  12303=>"000110011",
  12304=>"111101101",
  12305=>"101010100",
  12306=>"001111101",
  12307=>"100101010",
  12308=>"110100000",
  12309=>"100111100",
  12310=>"100111000",
  12311=>"001000010",
  12312=>"111100001",
  12313=>"100100110",
  12314=>"101100101",
  12315=>"110100111",
  12316=>"100010101",
  12317=>"100000110",
  12318=>"000101001",
  12319=>"001001000",
  12320=>"001000100",
  12321=>"000001100",
  12322=>"110101101",
  12323=>"111011111",
  12324=>"010010011",
  12325=>"010011001",
  12326=>"101111010",
  12327=>"010111100",
  12328=>"010100111",
  12329=>"010010001",
  12330=>"111000010",
  12331=>"110001010",
  12332=>"110000110",
  12333=>"111111011",
  12334=>"111111010",
  12335=>"010000100",
  12336=>"111100011",
  12337=>"101010010",
  12338=>"111010101",
  12339=>"110001001",
  12340=>"001101100",
  12341=>"000010000",
  12342=>"110100110",
  12343=>"010001100",
  12344=>"110111101",
  12345=>"101100110",
  12346=>"000011010",
  12347=>"100000001",
  12348=>"110010010",
  12349=>"101100101",
  12350=>"100101000",
  12351=>"000010101",
  12352=>"100011010",
  12353=>"010011111",
  12354=>"110100001",
  12355=>"001001101",
  12356=>"111111000",
  12357=>"101111000",
  12358=>"010111101",
  12359=>"100101011",
  12360=>"101011001",
  12361=>"110011111",
  12362=>"001000010",
  12363=>"000100111",
  12364=>"110011011",
  12365=>"001110110",
  12366=>"000100000",
  12367=>"111100101",
  12368=>"100101000",
  12369=>"001100110",
  12370=>"010110000",
  12371=>"101000101",
  12372=>"011111010",
  12373=>"110110000",
  12374=>"010000010",
  12375=>"101010100",
  12376=>"100011010",
  12377=>"000010000",
  12378=>"011100101",
  12379=>"001000000",
  12380=>"100010111",
  12381=>"100101100",
  12382=>"010111101",
  12383=>"001010110",
  12384=>"011001000",
  12385=>"000000101",
  12386=>"010001101",
  12387=>"100100100",
  12388=>"110011100",
  12389=>"010000100",
  12390=>"011111010",
  12391=>"000110110",
  12392=>"010000111",
  12393=>"101111010",
  12394=>"100000001",
  12395=>"010111111",
  12396=>"001111011",
  12397=>"010110011",
  12398=>"000010101",
  12399=>"000101001",
  12400=>"011110110",
  12401=>"010001000",
  12402=>"010011100",
  12403=>"000001111",
  12404=>"011110101",
  12405=>"001100010",
  12406=>"000000011",
  12407=>"010010100",
  12408=>"000111011",
  12409=>"111110010",
  12410=>"000101000",
  12411=>"000000111",
  12412=>"010011111",
  12413=>"111001000",
  12414=>"101010000",
  12415=>"111010000",
  12416=>"010101000",
  12417=>"000001101",
  12418=>"011101000",
  12419=>"000100101",
  12420=>"111110010",
  12421=>"001100100",
  12422=>"100110010",
  12423=>"000101101",
  12424=>"100111000",
  12425=>"000111101",
  12426=>"101100100",
  12427=>"100011110",
  12428=>"001110101",
  12429=>"101101111",
  12430=>"110110011",
  12431=>"011111111",
  12432=>"110111011",
  12433=>"000110111",
  12434=>"100101110",
  12435=>"111010011",
  12436=>"000111000",
  12437=>"101001110",
  12438=>"001010110",
  12439=>"100100101",
  12440=>"011110100",
  12441=>"111100000",
  12442=>"000111010",
  12443=>"111011010",
  12444=>"000010010",
  12445=>"011100100",
  12446=>"001010100",
  12447=>"001001111",
  12448=>"001011001",
  12449=>"100111100",
  12450=>"000101001",
  12451=>"001001100",
  12452=>"011100001",
  12453=>"110000111",
  12454=>"111001000",
  12455=>"110010110",
  12456=>"101010010",
  12457=>"110100000",
  12458=>"110000001",
  12459=>"101011001",
  12460=>"111010010",
  12461=>"000010110",
  12462=>"111100111",
  12463=>"110000100",
  12464=>"101111001",
  12465=>"000100111",
  12466=>"111101001",
  12467=>"011000000",
  12468=>"011101011",
  12469=>"011100110",
  12470=>"011001110",
  12471=>"111100010",
  12472=>"000011011",
  12473=>"001111110",
  12474=>"001101011",
  12475=>"111011011",
  12476=>"110101001",
  12477=>"001010000",
  12478=>"100100000",
  12479=>"100000011",
  12480=>"101100011",
  12481=>"111110101",
  12482=>"000000000",
  12483=>"111000000",
  12484=>"011110101",
  12485=>"010100000",
  12486=>"100110100",
  12487=>"101000100",
  12488=>"011011011",
  12489=>"001010011",
  12490=>"011010111",
  12491=>"011011101",
  12492=>"010100100",
  12493=>"110001010",
  12494=>"000001011",
  12495=>"111010100",
  12496=>"011000010",
  12497=>"001110111",
  12498=>"110111100",
  12499=>"011100010",
  12500=>"000000001",
  12501=>"001101010",
  12502=>"010110000",
  12503=>"101000011",
  12504=>"101001101",
  12505=>"011010100",
  12506=>"011011010",
  12507=>"011100110",
  12508=>"111010000",
  12509=>"101001110",
  12510=>"101111000",
  12511=>"101110100",
  12512=>"001101100",
  12513=>"111101000",
  12514=>"011001000",
  12515=>"000001000",
  12516=>"100000100",
  12517=>"001101011",
  12518=>"111000000",
  12519=>"011010010",
  12520=>"111001110",
  12521=>"001001001",
  12522=>"011000110",
  12523=>"101111011",
  12524=>"010101001",
  12525=>"011000101",
  12526=>"000110100",
  12527=>"110000110",
  12528=>"001111111",
  12529=>"010110001",
  12530=>"010100011",
  12531=>"010111111",
  12532=>"000110110",
  12533=>"100100000",
  12534=>"000001001",
  12535=>"011000101",
  12536=>"000011111",
  12537=>"111000001",
  12538=>"011010001",
  12539=>"000000010",
  12540=>"011111110",
  12541=>"011100000",
  12542=>"111111110",
  12543=>"001001000",
  12544=>"111011101",
  12545=>"010111010",
  12546=>"011011101",
  12547=>"000000111",
  12548=>"000111001",
  12549=>"110011101",
  12550=>"011001011",
  12551=>"100111110",
  12552=>"000000110",
  12553=>"110010011",
  12554=>"100001110",
  12555=>"011110100",
  12556=>"011010010",
  12557=>"001110000",
  12558=>"110100001",
  12559=>"000100110",
  12560=>"011000000",
  12561=>"000110101",
  12562=>"101001001",
  12563=>"110110100",
  12564=>"100100011",
  12565=>"011110101",
  12566=>"101011100",
  12567=>"101001010",
  12568=>"100011111",
  12569=>"001111001",
  12570=>"010110010",
  12571=>"011001001",
  12572=>"000100001",
  12573=>"011111110",
  12574=>"110010101",
  12575=>"000010001",
  12576=>"010001001",
  12577=>"110101011",
  12578=>"000011110",
  12579=>"111101100",
  12580=>"110011100",
  12581=>"001010111",
  12582=>"000001010",
  12583=>"111110101",
  12584=>"111111101",
  12585=>"110011101",
  12586=>"101111000",
  12587=>"000100010",
  12588=>"111101111",
  12589=>"000100100",
  12590=>"010111101",
  12591=>"011000000",
  12592=>"001010011",
  12593=>"100101010",
  12594=>"101010010",
  12595=>"000111000",
  12596=>"110111010",
  12597=>"110011101",
  12598=>"001111000",
  12599=>"111101100",
  12600=>"000001101",
  12601=>"101110101",
  12602=>"101001110",
  12603=>"000001111",
  12604=>"010001000",
  12605=>"000010010",
  12606=>"101011001",
  12607=>"011000111",
  12608=>"110101111",
  12609=>"010110101",
  12610=>"000111010",
  12611=>"011101010",
  12612=>"011001100",
  12613=>"100011110",
  12614=>"000001001",
  12615=>"100010000",
  12616=>"100011100",
  12617=>"011101110",
  12618=>"010101010",
  12619=>"101000010",
  12620=>"111101011",
  12621=>"000001101",
  12622=>"010111110",
  12623=>"110000100",
  12624=>"011011001",
  12625=>"011101110",
  12626=>"111011010",
  12627=>"000011001",
  12628=>"100011010",
  12629=>"110001000",
  12630=>"101110100",
  12631=>"100011000",
  12632=>"000110111",
  12633=>"000110011",
  12634=>"101110100",
  12635=>"010101100",
  12636=>"110011001",
  12637=>"000000010",
  12638=>"101111011",
  12639=>"000011110",
  12640=>"101010000",
  12641=>"110001100",
  12642=>"000001010",
  12643=>"001110001",
  12644=>"000101101",
  12645=>"101101110",
  12646=>"111110100",
  12647=>"110110111",
  12648=>"000010100",
  12649=>"101110001",
  12650=>"100111100",
  12651=>"000000101",
  12652=>"000111111",
  12653=>"100100001",
  12654=>"100000011",
  12655=>"011000101",
  12656=>"011010010",
  12657=>"111011100",
  12658=>"000110000",
  12659=>"110100000",
  12660=>"101011111",
  12661=>"001011001",
  12662=>"101111000",
  12663=>"001110001",
  12664=>"001110001",
  12665=>"000010110",
  12666=>"101000110",
  12667=>"100100100",
  12668=>"110110010",
  12669=>"110010110",
  12670=>"000001011",
  12671=>"000001001",
  12672=>"010100001",
  12673=>"000001011",
  12674=>"001100001",
  12675=>"000011000",
  12676=>"110101000",
  12677=>"110110111",
  12678=>"111110111",
  12679=>"000011000",
  12680=>"100000100",
  12681=>"110010000",
  12682=>"111101111",
  12683=>"010111001",
  12684=>"110001010",
  12685=>"101111000",
  12686=>"100011100",
  12687=>"011010010",
  12688=>"001101111",
  12689=>"000000111",
  12690=>"000010111",
  12691=>"101000100",
  12692=>"110101110",
  12693=>"100101101",
  12694=>"110110011",
  12695=>"111111101",
  12696=>"110010100",
  12697=>"001001010",
  12698=>"100101100",
  12699=>"001111000",
  12700=>"110100000",
  12701=>"000101101",
  12702=>"110110011",
  12703=>"110011001",
  12704=>"101000101",
  12705=>"000001111",
  12706=>"110110111",
  12707=>"001101100",
  12708=>"011011001",
  12709=>"000111000",
  12710=>"010010011",
  12711=>"000001101",
  12712=>"111010011",
  12713=>"011011000",
  12714=>"000101011",
  12715=>"100001001",
  12716=>"000001010",
  12717=>"101101010",
  12718=>"111110000",
  12719=>"011101000",
  12720=>"001100011",
  12721=>"101001110",
  12722=>"001100100",
  12723=>"101110100",
  12724=>"110110110",
  12725=>"010111001",
  12726=>"010001110",
  12727=>"011000111",
  12728=>"000001110",
  12729=>"001001001",
  12730=>"000000010",
  12731=>"000000010",
  12732=>"111000100",
  12733=>"111111001",
  12734=>"100011100",
  12735=>"100001000",
  12736=>"001111111",
  12737=>"000000010",
  12738=>"110111011",
  12739=>"111110001",
  12740=>"110001110",
  12741=>"010011010",
  12742=>"011100110",
  12743=>"101100101",
  12744=>"000101010",
  12745=>"110000011",
  12746=>"010110100",
  12747=>"101011000",
  12748=>"001101001",
  12749=>"001110110",
  12750=>"000110010",
  12751=>"001101100",
  12752=>"101000000",
  12753=>"001100000",
  12754=>"100100010",
  12755=>"000111000",
  12756=>"010100100",
  12757=>"100000010",
  12758=>"111111111",
  12759=>"000011010",
  12760=>"100001100",
  12761=>"110000111",
  12762=>"101011001",
  12763=>"010011011",
  12764=>"011001000",
  12765=>"001010101",
  12766=>"110011110",
  12767=>"010011010",
  12768=>"001010010",
  12769=>"110101110",
  12770=>"111111011",
  12771=>"101111110",
  12772=>"101011001",
  12773=>"101111000",
  12774=>"000100001",
  12775=>"010000010",
  12776=>"101111001",
  12777=>"011000000",
  12778=>"010110100",
  12779=>"001100011",
  12780=>"111011110",
  12781=>"110001010",
  12782=>"110100111",
  12783=>"111111000",
  12784=>"001001101",
  12785=>"011101001",
  12786=>"110110001",
  12787=>"111111101",
  12788=>"110001010",
  12789=>"101111110",
  12790=>"100111111",
  12791=>"001010111",
  12792=>"011001010",
  12793=>"111111100",
  12794=>"101010110",
  12795=>"010000010",
  12796=>"011100000",
  12797=>"110000100",
  12798=>"001010000",
  12799=>"100010101",
  12800=>"011011011",
  12801=>"000101010",
  12802=>"101010011",
  12803=>"010100001",
  12804=>"110111011",
  12805=>"110010011",
  12806=>"001101001",
  12807=>"010011011",
  12808=>"010100001",
  12809=>"001010011",
  12810=>"110100101",
  12811=>"011001100",
  12812=>"101100111",
  12813=>"110110110",
  12814=>"111110000",
  12815=>"010010111",
  12816=>"011111011",
  12817=>"000101101",
  12818=>"100001001",
  12819=>"111111000",
  12820=>"011110100",
  12821=>"101011000",
  12822=>"011000010",
  12823=>"101100110",
  12824=>"000100110",
  12825=>"010001011",
  12826=>"100101001",
  12827=>"111100101",
  12828=>"010100100",
  12829=>"110101010",
  12830=>"100111001",
  12831=>"000101001",
  12832=>"000111101",
  12833=>"101101110",
  12834=>"000101100",
  12835=>"000000001",
  12836=>"010011101",
  12837=>"100111110",
  12838=>"001011110",
  12839=>"110100001",
  12840=>"110000001",
  12841=>"010001100",
  12842=>"111111111",
  12843=>"001001000",
  12844=>"000000110",
  12845=>"001011000",
  12846=>"101110110",
  12847=>"011001100",
  12848=>"100001111",
  12849=>"011010111",
  12850=>"000111001",
  12851=>"010010011",
  12852=>"000000010",
  12853=>"010100010",
  12854=>"000100010",
  12855=>"100001110",
  12856=>"000101101",
  12857=>"001111000",
  12858=>"110011010",
  12859=>"010100111",
  12860=>"010010010",
  12861=>"011010101",
  12862=>"110110000",
  12863=>"100000110",
  12864=>"010110101",
  12865=>"000010110",
  12866=>"101011101",
  12867=>"111010100",
  12868=>"101100100",
  12869=>"101101001",
  12870=>"101100011",
  12871=>"110010011",
  12872=>"010010000",
  12873=>"011110000",
  12874=>"010111110",
  12875=>"010001000",
  12876=>"111110100",
  12877=>"100110001",
  12878=>"111000010",
  12879=>"000111110",
  12880=>"001001100",
  12881=>"011110011",
  12882=>"100111110",
  12883=>"000010100",
  12884=>"111100010",
  12885=>"000111100",
  12886=>"011110101",
  12887=>"001101011",
  12888=>"101011001",
  12889=>"100000000",
  12890=>"000111101",
  12891=>"000000010",
  12892=>"001101111",
  12893=>"000000100",
  12894=>"000011110",
  12895=>"010110010",
  12896=>"111000011",
  12897=>"100000000",
  12898=>"001101110",
  12899=>"110010110",
  12900=>"100001100",
  12901=>"011110000",
  12902=>"011011110",
  12903=>"110011001",
  12904=>"010011011",
  12905=>"000111111",
  12906=>"011100111",
  12907=>"000000000",
  12908=>"000110111",
  12909=>"111000111",
  12910=>"010011011",
  12911=>"000000110",
  12912=>"011001011",
  12913=>"010111010",
  12914=>"100100010",
  12915=>"110100111",
  12916=>"011010000",
  12917=>"110000000",
  12918=>"010110000",
  12919=>"011100000",
  12920=>"101000010",
  12921=>"111001110",
  12922=>"111000110",
  12923=>"010101011",
  12924=>"010100110",
  12925=>"011001011",
  12926=>"011010101",
  12927=>"110100111",
  12928=>"001011000",
  12929=>"001111111",
  12930=>"110101111",
  12931=>"000011000",
  12932=>"100011010",
  12933=>"101000001",
  12934=>"000100010",
  12935=>"011110111",
  12936=>"101101110",
  12937=>"110010110",
  12938=>"000101010",
  12939=>"010011111",
  12940=>"110010000",
  12941=>"101000000",
  12942=>"011100001",
  12943=>"011001000",
  12944=>"010100101",
  12945=>"101011101",
  12946=>"110011011",
  12947=>"100111101",
  12948=>"000100110",
  12949=>"000000011",
  12950=>"111101110",
  12951=>"111111110",
  12952=>"111100101",
  12953=>"000100110",
  12954=>"110011001",
  12955=>"100101101",
  12956=>"110100100",
  12957=>"111010011",
  12958=>"010010100",
  12959=>"111010000",
  12960=>"100000100",
  12961=>"010101010",
  12962=>"101100100",
  12963=>"111011111",
  12964=>"110011010",
  12965=>"011011000",
  12966=>"110010101",
  12967=>"010010111",
  12968=>"000000011",
  12969=>"010010100",
  12970=>"110100101",
  12971=>"111000011",
  12972=>"010010000",
  12973=>"001000110",
  12974=>"111111001",
  12975=>"100110010",
  12976=>"010101000",
  12977=>"100011000",
  12978=>"011111001",
  12979=>"000110001",
  12980=>"010100111",
  12981=>"001100011",
  12982=>"001100001",
  12983=>"110010001",
  12984=>"110100111",
  12985=>"001101100",
  12986=>"110100000",
  12987=>"011001011",
  12988=>"111011000",
  12989=>"101100000",
  12990=>"100000111",
  12991=>"000010100",
  12992=>"101010010",
  12993=>"000111010",
  12994=>"100110011",
  12995=>"011110000",
  12996=>"001101011",
  12997=>"000001110",
  12998=>"101110000",
  12999=>"010100100",
  13000=>"111011101",
  13001=>"011101011",
  13002=>"100111100",
  13003=>"110000111",
  13004=>"001011110",
  13005=>"110010010",
  13006=>"001001100",
  13007=>"101001000",
  13008=>"000010001",
  13009=>"110111111",
  13010=>"010100001",
  13011=>"011111000",
  13012=>"001101010",
  13013=>"000000111",
  13014=>"110001001",
  13015=>"101100100",
  13016=>"100001001",
  13017=>"100010001",
  13018=>"001000100",
  13019=>"111011111",
  13020=>"100100110",
  13021=>"001110111",
  13022=>"011111001",
  13023=>"011111000",
  13024=>"111110101",
  13025=>"111100100",
  13026=>"000010111",
  13027=>"110111111",
  13028=>"100101110",
  13029=>"011001111",
  13030=>"110101100",
  13031=>"111010010",
  13032=>"000111010",
  13033=>"010100100",
  13034=>"001111101",
  13035=>"110001010",
  13036=>"010011101",
  13037=>"110000001",
  13038=>"110111011",
  13039=>"101010000",
  13040=>"111111111",
  13041=>"101101110",
  13042=>"101100011",
  13043=>"111101000",
  13044=>"010111111",
  13045=>"010001010",
  13046=>"000011001",
  13047=>"111011110",
  13048=>"001000011",
  13049=>"011101000",
  13050=>"001101011",
  13051=>"011101110",
  13052=>"010001100",
  13053=>"100001000",
  13054=>"000110010",
  13055=>"010100000",
  13056=>"111100110",
  13057=>"110011011",
  13058=>"000000000",
  13059=>"011001010",
  13060=>"011101000",
  13061=>"010110011",
  13062=>"111101110",
  13063=>"111101001",
  13064=>"110010110",
  13065=>"101111111",
  13066=>"000010011",
  13067=>"101101000",
  13068=>"110100001",
  13069=>"010111000",
  13070=>"100100110",
  13071=>"011100001",
  13072=>"000011111",
  13073=>"011111100",
  13074=>"111001110",
  13075=>"010001000",
  13076=>"101000100",
  13077=>"110110100",
  13078=>"010001001",
  13079=>"110000111",
  13080=>"011001111",
  13081=>"101111101",
  13082=>"000101010",
  13083=>"000000101",
  13084=>"111011000",
  13085=>"001100010",
  13086=>"011000000",
  13087=>"101010001",
  13088=>"010101001",
  13089=>"001101111",
  13090=>"100001111",
  13091=>"000000110",
  13092=>"000100000",
  13093=>"101111101",
  13094=>"011111100",
  13095=>"101011110",
  13096=>"000100110",
  13097=>"111000000",
  13098=>"010011011",
  13099=>"000000100",
  13100=>"001011101",
  13101=>"101000011",
  13102=>"010101100",
  13103=>"100000000",
  13104=>"110010011",
  13105=>"001001000",
  13106=>"000100011",
  13107=>"101111000",
  13108=>"100000111",
  13109=>"101011010",
  13110=>"000110110",
  13111=>"110110110",
  13112=>"010100100",
  13113=>"110010010",
  13114=>"111111010",
  13115=>"000000000",
  13116=>"101110110",
  13117=>"101011011",
  13118=>"110000100",
  13119=>"001111010",
  13120=>"001010111",
  13121=>"111111111",
  13122=>"110001111",
  13123=>"110010010",
  13124=>"010111101",
  13125=>"010110010",
  13126=>"110111000",
  13127=>"010110111",
  13128=>"100001100",
  13129=>"100100011",
  13130=>"100001111",
  13131=>"110110111",
  13132=>"010111110",
  13133=>"110100101",
  13134=>"111000011",
  13135=>"101000110",
  13136=>"110110000",
  13137=>"101010101",
  13138=>"011111111",
  13139=>"101010100",
  13140=>"010001011",
  13141=>"000001101",
  13142=>"011101111",
  13143=>"111111001",
  13144=>"001001110",
  13145=>"010011111",
  13146=>"100111011",
  13147=>"111111010",
  13148=>"110111001",
  13149=>"100010100",
  13150=>"110001010",
  13151=>"000000010",
  13152=>"000110110",
  13153=>"111101001",
  13154=>"000101110",
  13155=>"000110101",
  13156=>"001000001",
  13157=>"110000000",
  13158=>"010001011",
  13159=>"001011001",
  13160=>"111110110",
  13161=>"100010110",
  13162=>"111010100",
  13163=>"110001010",
  13164=>"101001111",
  13165=>"110101001",
  13166=>"101111011",
  13167=>"001101011",
  13168=>"001101001",
  13169=>"110010000",
  13170=>"111111001",
  13171=>"100111001",
  13172=>"000010000",
  13173=>"001110100",
  13174=>"000001111",
  13175=>"101100100",
  13176=>"100000010",
  13177=>"110011001",
  13178=>"111001111",
  13179=>"000001111",
  13180=>"000010000",
  13181=>"010000101",
  13182=>"100100101",
  13183=>"000011011",
  13184=>"000110010",
  13185=>"010110111",
  13186=>"000000111",
  13187=>"010101010",
  13188=>"110100011",
  13189=>"110000010",
  13190=>"001010010",
  13191=>"000101111",
  13192=>"001111100",
  13193=>"001000011",
  13194=>"000010000",
  13195=>"001000101",
  13196=>"111100011",
  13197=>"001010011",
  13198=>"000000001",
  13199=>"001010100",
  13200=>"011000111",
  13201=>"011010000",
  13202=>"101001000",
  13203=>"111101111",
  13204=>"111111110",
  13205=>"101011100",
  13206=>"111100111",
  13207=>"010011101",
  13208=>"001111000",
  13209=>"111000100",
  13210=>"010100000",
  13211=>"000110100",
  13212=>"000100111",
  13213=>"101001101",
  13214=>"101001100",
  13215=>"100001001",
  13216=>"111011111",
  13217=>"111100110",
  13218=>"100001000",
  13219=>"000010111",
  13220=>"100111101",
  13221=>"101111100",
  13222=>"100111010",
  13223=>"000101001",
  13224=>"011000100",
  13225=>"100011000",
  13226=>"111011010",
  13227=>"110111110",
  13228=>"110100011",
  13229=>"010110011",
  13230=>"110111101",
  13231=>"111101111",
  13232=>"010010101",
  13233=>"101001010",
  13234=>"011011100",
  13235=>"001000000",
  13236=>"110111011",
  13237=>"001111010",
  13238=>"111101100",
  13239=>"111010100",
  13240=>"011000101",
  13241=>"011001101",
  13242=>"100110011",
  13243=>"110010110",
  13244=>"011111100",
  13245=>"001011010",
  13246=>"101000001",
  13247=>"001001000",
  13248=>"010101001",
  13249=>"010000000",
  13250=>"100111011",
  13251=>"101111001",
  13252=>"000110011",
  13253=>"001110010",
  13254=>"111111011",
  13255=>"110110010",
  13256=>"000100100",
  13257=>"101100111",
  13258=>"100100111",
  13259=>"001100101",
  13260=>"101010110",
  13261=>"110110100",
  13262=>"100110001",
  13263=>"111000011",
  13264=>"011101010",
  13265=>"101001110",
  13266=>"111110110",
  13267=>"100101000",
  13268=>"101011011",
  13269=>"101101110",
  13270=>"110000111",
  13271=>"000100000",
  13272=>"000000011",
  13273=>"110010000",
  13274=>"011011011",
  13275=>"010001010",
  13276=>"111001100",
  13277=>"111000111",
  13278=>"110110000",
  13279=>"011000011",
  13280=>"101001101",
  13281=>"100100011",
  13282=>"000101011",
  13283=>"010111011",
  13284=>"001100000",
  13285=>"110010001",
  13286=>"100110111",
  13287=>"000100101",
  13288=>"001010010",
  13289=>"001101011",
  13290=>"000101010",
  13291=>"100011010",
  13292=>"100111000",
  13293=>"111010101",
  13294=>"010001110",
  13295=>"101110000",
  13296=>"001100100",
  13297=>"011000111",
  13298=>"001111111",
  13299=>"011101101",
  13300=>"110100100",
  13301=>"111000010",
  13302=>"110110000",
  13303=>"010010010",
  13304=>"000100111",
  13305=>"010111111",
  13306=>"111001101",
  13307=>"101010111",
  13308=>"010010100",
  13309=>"101001001",
  13310=>"011110100",
  13311=>"011001000",
  13312=>"000100011",
  13313=>"011111111",
  13314=>"000010000",
  13315=>"101010010",
  13316=>"101001001",
  13317=>"000001000",
  13318=>"111111011",
  13319=>"001011001",
  13320=>"110110000",
  13321=>"111010110",
  13322=>"111111001",
  13323=>"000011011",
  13324=>"001110100",
  13325=>"001111010",
  13326=>"101001001",
  13327=>"000101100",
  13328=>"001111101",
  13329=>"010000001",
  13330=>"110111011",
  13331=>"101111101",
  13332=>"111010101",
  13333=>"001001001",
  13334=>"101011011",
  13335=>"001101111",
  13336=>"010111100",
  13337=>"010100010",
  13338=>"001110110",
  13339=>"100001111",
  13340=>"001011110",
  13341=>"111000101",
  13342=>"000011001",
  13343=>"011100001",
  13344=>"110010110",
  13345=>"011111001",
  13346=>"111111001",
  13347=>"010111111",
  13348=>"011010100",
  13349=>"100100010",
  13350=>"000100101",
  13351=>"101100011",
  13352=>"100101011",
  13353=>"000101010",
  13354=>"010010101",
  13355=>"010001010",
  13356=>"111101000",
  13357=>"000001111",
  13358=>"011111101",
  13359=>"100100001",
  13360=>"011111101",
  13361=>"010110110",
  13362=>"110000111",
  13363=>"001110100",
  13364=>"111010110",
  13365=>"111100000",
  13366=>"111010110",
  13367=>"000101111",
  13368=>"000010110",
  13369=>"111001011",
  13370=>"100111100",
  13371=>"001001111",
  13372=>"001111110",
  13373=>"011100010",
  13374=>"110000001",
  13375=>"010100101",
  13376=>"011111110",
  13377=>"100001011",
  13378=>"110011110",
  13379=>"000010111",
  13380=>"101100101",
  13381=>"001001100",
  13382=>"000001110",
  13383=>"100100000",
  13384=>"111000010",
  13385=>"101111010",
  13386=>"100000011",
  13387=>"101011101",
  13388=>"100111010",
  13389=>"110101110",
  13390=>"010110110",
  13391=>"110100001",
  13392=>"110000110",
  13393=>"010110111",
  13394=>"011000011",
  13395=>"001001011",
  13396=>"101011001",
  13397=>"101000101",
  13398=>"001111110",
  13399=>"000001100",
  13400=>"111011101",
  13401=>"011110100",
  13402=>"001000110",
  13403=>"000101011",
  13404=>"101000000",
  13405=>"110100111",
  13406=>"100011001",
  13407=>"011001110",
  13408=>"101011001",
  13409=>"011110111",
  13410=>"010000011",
  13411=>"100010010",
  13412=>"110100010",
  13413=>"010000110",
  13414=>"111010100",
  13415=>"000110110",
  13416=>"010011110",
  13417=>"100000010",
  13418=>"010001111",
  13419=>"110011000",
  13420=>"000011101",
  13421=>"100110000",
  13422=>"111010010",
  13423=>"010111101",
  13424=>"011001000",
  13425=>"101111100",
  13426=>"010111111",
  13427=>"101111111",
  13428=>"001110000",
  13429=>"110001001",
  13430=>"010110111",
  13431=>"000000001",
  13432=>"010000100",
  13433=>"101001001",
  13434=>"010001100",
  13435=>"100111011",
  13436=>"011100011",
  13437=>"010110010",
  13438=>"011011000",
  13439=>"110011000",
  13440=>"001101010",
  13441=>"000101001",
  13442=>"000101111",
  13443=>"100101010",
  13444=>"000000010",
  13445=>"001110101",
  13446=>"110011000",
  13447=>"101000011",
  13448=>"001011000",
  13449=>"001110000",
  13450=>"101001011",
  13451=>"010100011",
  13452=>"010101011",
  13453=>"101110100",
  13454=>"000011110",
  13455=>"101101101",
  13456=>"001011111",
  13457=>"101000011",
  13458=>"010110101",
  13459=>"001001111",
  13460=>"000000000",
  13461=>"000110001",
  13462=>"111000111",
  13463=>"100011101",
  13464=>"000101001",
  13465=>"010100100",
  13466=>"101100110",
  13467=>"000010100",
  13468=>"001000001",
  13469=>"101100111",
  13470=>"000011010",
  13471=>"111000011",
  13472=>"111000000",
  13473=>"111110001",
  13474=>"000001011",
  13475=>"010101000",
  13476=>"110101001",
  13477=>"101100111",
  13478=>"111111111",
  13479=>"010000100",
  13480=>"110110011",
  13481=>"110010101",
  13482=>"110000111",
  13483=>"010010001",
  13484=>"111000111",
  13485=>"101111101",
  13486=>"101101100",
  13487=>"000101000",
  13488=>"000111001",
  13489=>"011010110",
  13490=>"111110010",
  13491=>"011001000",
  13492=>"110010010",
  13493=>"010000001",
  13494=>"000000111",
  13495=>"011000011",
  13496=>"001110001",
  13497=>"001001000",
  13498=>"001000111",
  13499=>"111000101",
  13500=>"011111010",
  13501=>"001011110",
  13502=>"010000111",
  13503=>"110111000",
  13504=>"000001110",
  13505=>"100111011",
  13506=>"000001010",
  13507=>"100000110",
  13508=>"001100001",
  13509=>"000111010",
  13510=>"111011100",
  13511=>"111100100",
  13512=>"010111010",
  13513=>"010011111",
  13514=>"101111110",
  13515=>"111110010",
  13516=>"111110101",
  13517=>"101111110",
  13518=>"000101010",
  13519=>"111100001",
  13520=>"101001111",
  13521=>"101010000",
  13522=>"101011010",
  13523=>"111011011",
  13524=>"110101100",
  13525=>"110100110",
  13526=>"111011110",
  13527=>"110011100",
  13528=>"100111011",
  13529=>"110000100",
  13530=>"100110101",
  13531=>"000110010",
  13532=>"101010010",
  13533=>"111000101",
  13534=>"101010000",
  13535=>"011111101",
  13536=>"010000111",
  13537=>"011111101",
  13538=>"000011100",
  13539=>"100000111",
  13540=>"111010010",
  13541=>"011111010",
  13542=>"010101011",
  13543=>"101000100",
  13544=>"101000101",
  13545=>"000110000",
  13546=>"110000100",
  13547=>"000011100",
  13548=>"010001101",
  13549=>"001000101",
  13550=>"101001111",
  13551=>"101111000",
  13552=>"010110100",
  13553=>"011110111",
  13554=>"001100100",
  13555=>"000000110",
  13556=>"100000001",
  13557=>"011100110",
  13558=>"000001111",
  13559=>"001111010",
  13560=>"000000100",
  13561=>"110001001",
  13562=>"001110001",
  13563=>"011111000",
  13564=>"010110101",
  13565=>"011011011",
  13566=>"000001001",
  13567=>"100111111",
  13568=>"011000000",
  13569=>"011001011",
  13570=>"011001000",
  13571=>"000101110",
  13572=>"000000100",
  13573=>"011101111",
  13574=>"100110101",
  13575=>"100101011",
  13576=>"000100100",
  13577=>"010001010",
  13578=>"011011110",
  13579=>"001110000",
  13580=>"011010010",
  13581=>"000011011",
  13582=>"010100001",
  13583=>"111111001",
  13584=>"111101111",
  13585=>"101001100",
  13586=>"101110010",
  13587=>"011011101",
  13588=>"101011100",
  13589=>"110011000",
  13590=>"010100001",
  13591=>"101110000",
  13592=>"001000010",
  13593=>"111010001",
  13594=>"010110000",
  13595=>"111011110",
  13596=>"000111001",
  13597=>"100001101",
  13598=>"101110010",
  13599=>"010100110",
  13600=>"000001110",
  13601=>"000110110",
  13602=>"100111001",
  13603=>"000110001",
  13604=>"111001001",
  13605=>"100111000",
  13606=>"001011110",
  13607=>"110110010",
  13608=>"000010111",
  13609=>"000110110",
  13610=>"001001110",
  13611=>"100000000",
  13612=>"101000101",
  13613=>"010000011",
  13614=>"000101011",
  13615=>"100111101",
  13616=>"110000110",
  13617=>"000001101",
  13618=>"010011110",
  13619=>"011011101",
  13620=>"110001010",
  13621=>"000010101",
  13622=>"010010111",
  13623=>"000000000",
  13624=>"100001111",
  13625=>"011101001",
  13626=>"100111111",
  13627=>"100010000",
  13628=>"011111111",
  13629=>"000110100",
  13630=>"111101111",
  13631=>"101001100",
  13632=>"011000001",
  13633=>"010001010",
  13634=>"010000101",
  13635=>"101111111",
  13636=>"111100000",
  13637=>"110001000",
  13638=>"001001000",
  13639=>"100001111",
  13640=>"000000101",
  13641=>"001111011",
  13642=>"000111111",
  13643=>"101100000",
  13644=>"110000000",
  13645=>"000110111",
  13646=>"101110011",
  13647=>"111111001",
  13648=>"101000010",
  13649=>"110011001",
  13650=>"001110110",
  13651=>"100100101",
  13652=>"110100011",
  13653=>"010100000",
  13654=>"111100100",
  13655=>"111101101",
  13656=>"010010011",
  13657=>"001110001",
  13658=>"000100111",
  13659=>"000110011",
  13660=>"101011110",
  13661=>"011101001",
  13662=>"010111010",
  13663=>"000001111",
  13664=>"100001100",
  13665=>"110010101",
  13666=>"011100001",
  13667=>"101010111",
  13668=>"010101111",
  13669=>"000001011",
  13670=>"100001111",
  13671=>"000000000",
  13672=>"000101101",
  13673=>"101110110",
  13674=>"011100011",
  13675=>"010001101",
  13676=>"000010000",
  13677=>"101101001",
  13678=>"000110110",
  13679=>"000010010",
  13680=>"100100101",
  13681=>"011000010",
  13682=>"010111110",
  13683=>"000000101",
  13684=>"111001000",
  13685=>"110101111",
  13686=>"000011101",
  13687=>"101111110",
  13688=>"001011001",
  13689=>"011100111",
  13690=>"110111100",
  13691=>"010000001",
  13692=>"111111001",
  13693=>"001010101",
  13694=>"011011001",
  13695=>"001001010",
  13696=>"100100110",
  13697=>"100000011",
  13698=>"110011011",
  13699=>"111001000",
  13700=>"111010010",
  13701=>"010010101",
  13702=>"000001100",
  13703=>"111010011",
  13704=>"000100110",
  13705=>"100001110",
  13706=>"001101001",
  13707=>"100010100",
  13708=>"001111010",
  13709=>"001011010",
  13710=>"111110011",
  13711=>"010000000",
  13712=>"101100001",
  13713=>"000010111",
  13714=>"011011101",
  13715=>"101100100",
  13716=>"011011111",
  13717=>"111100100",
  13718=>"011110110",
  13719=>"100000010",
  13720=>"111011100",
  13721=>"011010010",
  13722=>"011110011",
  13723=>"011011111",
  13724=>"010100011",
  13725=>"001010000",
  13726=>"001111110",
  13727=>"111001011",
  13728=>"100000011",
  13729=>"011000011",
  13730=>"111001111",
  13731=>"011100110",
  13732=>"010100010",
  13733=>"100001101",
  13734=>"100001000",
  13735=>"101000000",
  13736=>"101111111",
  13737=>"011000011",
  13738=>"011110111",
  13739=>"101010111",
  13740=>"000011000",
  13741=>"001111100",
  13742=>"101000011",
  13743=>"001110010",
  13744=>"010101001",
  13745=>"101110000",
  13746=>"101100001",
  13747=>"111111100",
  13748=>"010100110",
  13749=>"010100011",
  13750=>"011001010",
  13751=>"101000000",
  13752=>"110011101",
  13753=>"101111000",
  13754=>"001110011",
  13755=>"010011100",
  13756=>"101010001",
  13757=>"100101110",
  13758=>"010000110",
  13759=>"110011111",
  13760=>"101111110",
  13761=>"111001101",
  13762=>"001011110",
  13763=>"111001001",
  13764=>"011011011",
  13765=>"111110101",
  13766=>"011000010",
  13767=>"010010101",
  13768=>"001111110",
  13769=>"101110001",
  13770=>"000111111",
  13771=>"100110000",
  13772=>"101010110",
  13773=>"100000011",
  13774=>"000100111",
  13775=>"010000000",
  13776=>"111110111",
  13777=>"010001010",
  13778=>"111101001",
  13779=>"110110111",
  13780=>"111010100",
  13781=>"111010001",
  13782=>"110100001",
  13783=>"010011101",
  13784=>"011000101",
  13785=>"000100001",
  13786=>"001011111",
  13787=>"001001011",
  13788=>"110101010",
  13789=>"000101100",
  13790=>"110010011",
  13791=>"100110110",
  13792=>"010000101",
  13793=>"011111100",
  13794=>"010100010",
  13795=>"011001111",
  13796=>"100000000",
  13797=>"111010000",
  13798=>"110111000",
  13799=>"100001110",
  13800=>"010110010",
  13801=>"011111100",
  13802=>"100101010",
  13803=>"001010001",
  13804=>"111001110",
  13805=>"010111110",
  13806=>"101001110",
  13807=>"111010011",
  13808=>"111101011",
  13809=>"011111011",
  13810=>"110100100",
  13811=>"011101101",
  13812=>"000110001",
  13813=>"100101001",
  13814=>"010011000",
  13815=>"010111010",
  13816=>"010101000",
  13817=>"000101010",
  13818=>"001001101",
  13819=>"001110001",
  13820=>"011111111",
  13821=>"110001010",
  13822=>"111101001",
  13823=>"000011001",
  13824=>"010100100",
  13825=>"100101001",
  13826=>"001100001",
  13827=>"001010101",
  13828=>"101010011",
  13829=>"110100100",
  13830=>"100100111",
  13831=>"111100111",
  13832=>"100010011",
  13833=>"001010111",
  13834=>"111010011",
  13835=>"011011000",
  13836=>"101001011",
  13837=>"001111000",
  13838=>"111011010",
  13839=>"101010000",
  13840=>"100110010",
  13841=>"101000111",
  13842=>"110011111",
  13843=>"101000010",
  13844=>"111010100",
  13845=>"101110011",
  13846=>"111100010",
  13847=>"111110110",
  13848=>"110000100",
  13849=>"101100111",
  13850=>"100110011",
  13851=>"101100100",
  13852=>"010001001",
  13853=>"000011001",
  13854=>"100001111",
  13855=>"010101111",
  13856=>"101110001",
  13857=>"110111000",
  13858=>"101101011",
  13859=>"100001011",
  13860=>"101000111",
  13861=>"010010000",
  13862=>"100101001",
  13863=>"111001101",
  13864=>"110100101",
  13865=>"010101000",
  13866=>"000111100",
  13867=>"000110010",
  13868=>"011110000",
  13869=>"111011011",
  13870=>"010010100",
  13871=>"001011110",
  13872=>"011111001",
  13873=>"011111100",
  13874=>"001000010",
  13875=>"101011101",
  13876=>"011010110",
  13877=>"010111110",
  13878=>"101110110",
  13879=>"010000101",
  13880=>"110100110",
  13881=>"010010111",
  13882=>"100110010",
  13883=>"000101000",
  13884=>"110111100",
  13885=>"001000111",
  13886=>"111000010",
  13887=>"000010001",
  13888=>"000010001",
  13889=>"000100101",
  13890=>"111111001",
  13891=>"000010110",
  13892=>"000001101",
  13893=>"010111001",
  13894=>"101010100",
  13895=>"110000100",
  13896=>"010000011",
  13897=>"100101011",
  13898=>"101101101",
  13899=>"110010110",
  13900=>"010010000",
  13901=>"111011010",
  13902=>"100111110",
  13903=>"100111011",
  13904=>"010110011",
  13905=>"000010001",
  13906=>"011010001",
  13907=>"001011000",
  13908=>"010010000",
  13909=>"011111100",
  13910=>"111100110",
  13911=>"001110010",
  13912=>"101100100",
  13913=>"010000001",
  13914=>"000100001",
  13915=>"100101011",
  13916=>"101000110",
  13917=>"111001010",
  13918=>"000111010",
  13919=>"101100000",
  13920=>"110111111",
  13921=>"001011000",
  13922=>"110010001",
  13923=>"011111111",
  13924=>"001000000",
  13925=>"000000100",
  13926=>"101000100",
  13927=>"010001011",
  13928=>"111110000",
  13929=>"101011010",
  13930=>"100110010",
  13931=>"001111101",
  13932=>"011010010",
  13933=>"001110000",
  13934=>"010110111",
  13935=>"000101010",
  13936=>"110100110",
  13937=>"110010001",
  13938=>"110000111",
  13939=>"000110000",
  13940=>"100101011",
  13941=>"010010000",
  13942=>"101010111",
  13943=>"011000000",
  13944=>"001011010",
  13945=>"000101111",
  13946=>"100101010",
  13947=>"001101101",
  13948=>"011101000",
  13949=>"011111000",
  13950=>"010100000",
  13951=>"001110111",
  13952=>"010010110",
  13953=>"101011001",
  13954=>"000100001",
  13955=>"110000111",
  13956=>"011000111",
  13957=>"001000001",
  13958=>"110111110",
  13959=>"111101100",
  13960=>"101110111",
  13961=>"101010010",
  13962=>"011011011",
  13963=>"100100111",
  13964=>"100010000",
  13965=>"101100110",
  13966=>"101011010",
  13967=>"111110110",
  13968=>"101111110",
  13969=>"000010100",
  13970=>"110101110",
  13971=>"110000100",
  13972=>"011100010",
  13973=>"110101010",
  13974=>"110101010",
  13975=>"100110111",
  13976=>"011000000",
  13977=>"000000001",
  13978=>"000011111",
  13979=>"011100000",
  13980=>"010101001",
  13981=>"000100010",
  13982=>"010010100",
  13983=>"011001111",
  13984=>"001000110",
  13985=>"100001010",
  13986=>"001000011",
  13987=>"111011011",
  13988=>"001000101",
  13989=>"000000111",
  13990=>"010011111",
  13991=>"010000000",
  13992=>"001101111",
  13993=>"000111001",
  13994=>"011001110",
  13995=>"011000010",
  13996=>"110010001",
  13997=>"000001110",
  13998=>"110011010",
  13999=>"100111011",
  14000=>"000011001",
  14001=>"011010100",
  14002=>"001001111",
  14003=>"001000110",
  14004=>"100101010",
  14005=>"000011011",
  14006=>"000110001",
  14007=>"100111101",
  14008=>"001000111",
  14009=>"000001000",
  14010=>"111101011",
  14011=>"101110000",
  14012=>"010000101",
  14013=>"011101001",
  14014=>"011000100",
  14015=>"110000100",
  14016=>"001100111",
  14017=>"000011110",
  14018=>"010011100",
  14019=>"010111011",
  14020=>"011010001",
  14021=>"101101010",
  14022=>"110111001",
  14023=>"001110100",
  14024=>"000000101",
  14025=>"000001100",
  14026=>"001010110",
  14027=>"000000101",
  14028=>"001111011",
  14029=>"011110011",
  14030=>"110101100",
  14031=>"000101101",
  14032=>"011010011",
  14033=>"101111011",
  14034=>"100100001",
  14035=>"000101111",
  14036=>"100111111",
  14037=>"010010010",
  14038=>"101111011",
  14039=>"001101011",
  14040=>"011101101",
  14041=>"011000001",
  14042=>"001000100",
  14043=>"110111001",
  14044=>"110001000",
  14045=>"010011110",
  14046=>"111010000",
  14047=>"011011011",
  14048=>"111101001",
  14049=>"010100010",
  14050=>"001001100",
  14051=>"010110110",
  14052=>"010101010",
  14053=>"110110011",
  14054=>"111111010",
  14055=>"001101001",
  14056=>"101110111",
  14057=>"011110010",
  14058=>"011001010",
  14059=>"100011011",
  14060=>"111000001",
  14061=>"110010100",
  14062=>"101111011",
  14063=>"001000110",
  14064=>"011111010",
  14065=>"000011011",
  14066=>"000010110",
  14067=>"000001000",
  14068=>"111111001",
  14069=>"110001100",
  14070=>"111100101",
  14071=>"100100001",
  14072=>"010010110",
  14073=>"000101111",
  14074=>"110111001",
  14075=>"010001100",
  14076=>"100111101",
  14077=>"011011110",
  14078=>"010000000",
  14079=>"010011000",
  14080=>"111010011",
  14081=>"000000010",
  14082=>"001001000",
  14083=>"111001101",
  14084=>"101110001",
  14085=>"101011010",
  14086=>"101000101",
  14087=>"011010011",
  14088=>"000101010",
  14089=>"110010100",
  14090=>"010000010",
  14091=>"000100000",
  14092=>"000101110",
  14093=>"101100001",
  14094=>"110111101",
  14095=>"111101011",
  14096=>"100101000",
  14097=>"111100001",
  14098=>"000111101",
  14099=>"100101010",
  14100=>"000011010",
  14101=>"010010001",
  14102=>"010110001",
  14103=>"011011101",
  14104=>"001000111",
  14105=>"110101111",
  14106=>"000101111",
  14107=>"101100011",
  14108=>"000100100",
  14109=>"110010011",
  14110=>"000000110",
  14111=>"010111110",
  14112=>"110011011",
  14113=>"111010110",
  14114=>"110011011",
  14115=>"000000110",
  14116=>"110111010",
  14117=>"000100100",
  14118=>"110100011",
  14119=>"100100111",
  14120=>"011100000",
  14121=>"011011000",
  14122=>"101000110",
  14123=>"110101100",
  14124=>"100010001",
  14125=>"110100110",
  14126=>"100000100",
  14127=>"010111101",
  14128=>"101101000",
  14129=>"001100010",
  14130=>"010100100",
  14131=>"101001001",
  14132=>"101111000",
  14133=>"110000111",
  14134=>"000000001",
  14135=>"001011011",
  14136=>"110101001",
  14137=>"100001010",
  14138=>"110001011",
  14139=>"000101100",
  14140=>"111110000",
  14141=>"000000111",
  14142=>"011110111",
  14143=>"100000001",
  14144=>"001010101",
  14145=>"010000000",
  14146=>"001110000",
  14147=>"000100111",
  14148=>"001001010",
  14149=>"110100010",
  14150=>"100100010",
  14151=>"001010010",
  14152=>"000011111",
  14153=>"101101001",
  14154=>"011110100",
  14155=>"100000000",
  14156=>"010010001",
  14157=>"111111111",
  14158=>"001001000",
  14159=>"111011000",
  14160=>"001110111",
  14161=>"000110111",
  14162=>"001100100",
  14163=>"000010010",
  14164=>"100011010",
  14165=>"100110000",
  14166=>"111001111",
  14167=>"001101001",
  14168=>"110000011",
  14169=>"111111001",
  14170=>"001111001",
  14171=>"000101011",
  14172=>"001110110",
  14173=>"110010011",
  14174=>"100101101",
  14175=>"000000100",
  14176=>"001010100",
  14177=>"010010001",
  14178=>"001110101",
  14179=>"100100110",
  14180=>"101000111",
  14181=>"000100100",
  14182=>"011111111",
  14183=>"000001010",
  14184=>"001000101",
  14185=>"000001001",
  14186=>"110010101",
  14187=>"111011000",
  14188=>"000111100",
  14189=>"000011001",
  14190=>"100001100",
  14191=>"001000110",
  14192=>"110101100",
  14193=>"111100010",
  14194=>"111001110",
  14195=>"010001101",
  14196=>"001100111",
  14197=>"110011110",
  14198=>"111111000",
  14199=>"110100111",
  14200=>"100000100",
  14201=>"101110110",
  14202=>"010101101",
  14203=>"011100010",
  14204=>"000010011",
  14205=>"111110100",
  14206=>"111010011",
  14207=>"111001011",
  14208=>"000001111",
  14209=>"100000000",
  14210=>"011001100",
  14211=>"101110010",
  14212=>"010101011",
  14213=>"110000000",
  14214=>"101110111",
  14215=>"001100101",
  14216=>"011001111",
  14217=>"110001001",
  14218=>"000110111",
  14219=>"101010101",
  14220=>"010010101",
  14221=>"010010001",
  14222=>"110110011",
  14223=>"110000111",
  14224=>"100011100",
  14225=>"111001011",
  14226=>"000010010",
  14227=>"010001110",
  14228=>"000011000",
  14229=>"000100000",
  14230=>"011110100",
  14231=>"011111001",
  14232=>"011010101",
  14233=>"000010111",
  14234=>"000011000",
  14235=>"100001010",
  14236=>"100111000",
  14237=>"000010010",
  14238=>"101000111",
  14239=>"001000101",
  14240=>"001001001",
  14241=>"111101101",
  14242=>"000001110",
  14243=>"000001101",
  14244=>"100000101",
  14245=>"011001100",
  14246=>"011100101",
  14247=>"010111111",
  14248=>"011001001",
  14249=>"111101101",
  14250=>"010000011",
  14251=>"111101011",
  14252=>"011011110",
  14253=>"100110100",
  14254=>"000100110",
  14255=>"000101100",
  14256=>"101000010",
  14257=>"110101000",
  14258=>"001001100",
  14259=>"010111111",
  14260=>"000111010",
  14261=>"011011100",
  14262=>"010000100",
  14263=>"111001111",
  14264=>"000000001",
  14265=>"010001110",
  14266=>"110101100",
  14267=>"110010100",
  14268=>"110110110",
  14269=>"100101101",
  14270=>"000101111",
  14271=>"100000011",
  14272=>"011101010",
  14273=>"110101000",
  14274=>"001000000",
  14275=>"000010100",
  14276=>"000111101",
  14277=>"001001001",
  14278=>"111101001",
  14279=>"100111011",
  14280=>"001000011",
  14281=>"100011010",
  14282=>"011100101",
  14283=>"000010011",
  14284=>"011011001",
  14285=>"000000000",
  14286=>"010001000",
  14287=>"000010111",
  14288=>"110010001",
  14289=>"000100010",
  14290=>"010101110",
  14291=>"001010000",
  14292=>"111001010",
  14293=>"100111010",
  14294=>"010011010",
  14295=>"000010100",
  14296=>"001010010",
  14297=>"001000110",
  14298=>"010110010",
  14299=>"011001001",
  14300=>"111111100",
  14301=>"011001010",
  14302=>"100001110",
  14303=>"111111000",
  14304=>"000100000",
  14305=>"011110110",
  14306=>"101101010",
  14307=>"101011011",
  14308=>"000001010",
  14309=>"111100100",
  14310=>"110111010",
  14311=>"010100100",
  14312=>"000100111",
  14313=>"101011110",
  14314=>"001001000",
  14315=>"000010011",
  14316=>"001111101",
  14317=>"000010001",
  14318=>"000110001",
  14319=>"010101001",
  14320=>"011100010",
  14321=>"100100100",
  14322=>"100010100",
  14323=>"010111110",
  14324=>"101101111",
  14325=>"011111110",
  14326=>"001010110",
  14327=>"000011111",
  14328=>"100010001",
  14329=>"001100001",
  14330=>"110000111",
  14331=>"011100111",
  14332=>"110101111",
  14333=>"000110000",
  14334=>"011110111",
  14335=>"100101111",
  14336=>"001111010",
  14337=>"011111011",
  14338=>"100111100",
  14339=>"101100000",
  14340=>"111001010",
  14341=>"100101110",
  14342=>"010100101",
  14343=>"100001101",
  14344=>"111011100",
  14345=>"001110100",
  14346=>"000110010",
  14347=>"110111110",
  14348=>"010011010",
  14349=>"110011011",
  14350=>"101111111",
  14351=>"000011111",
  14352=>"001101000",
  14353=>"010110100",
  14354=>"010100101",
  14355=>"101110000",
  14356=>"000010010",
  14357=>"101010001",
  14358=>"100111000",
  14359=>"001110010",
  14360=>"001000000",
  14361=>"100010010",
  14362=>"111101011",
  14363=>"101110110",
  14364=>"010011011",
  14365=>"100000110",
  14366=>"100011010",
  14367=>"100100001",
  14368=>"011110010",
  14369=>"000101011",
  14370=>"100000001",
  14371=>"000001101",
  14372=>"011010110",
  14373=>"111010111",
  14374=>"111100100",
  14375=>"101110011",
  14376=>"010111001",
  14377=>"001001101",
  14378=>"100010001",
  14379=>"100110111",
  14380=>"010000001",
  14381=>"100010100",
  14382=>"000011010",
  14383=>"000000101",
  14384=>"011000110",
  14385=>"110111001",
  14386=>"110011010",
  14387=>"000100100",
  14388=>"110000000",
  14389=>"000001000",
  14390=>"000111001",
  14391=>"000001100",
  14392=>"111010000",
  14393=>"001000101",
  14394=>"000111010",
  14395=>"000100010",
  14396=>"100010011",
  14397=>"011010110",
  14398=>"011110001",
  14399=>"010111100",
  14400=>"000011010",
  14401=>"001101010",
  14402=>"011101010",
  14403=>"110101100",
  14404=>"101111101",
  14405=>"011110111",
  14406=>"111001101",
  14407=>"010000111",
  14408=>"100010000",
  14409=>"111110010",
  14410=>"001010010",
  14411=>"000001110",
  14412=>"111111110",
  14413=>"000010111",
  14414=>"111001010",
  14415=>"100110111",
  14416=>"000001000",
  14417=>"000001000",
  14418=>"011101101",
  14419=>"111011100",
  14420=>"101001011",
  14421=>"001001111",
  14422=>"000111011",
  14423=>"001001101",
  14424=>"100110111",
  14425=>"000111111",
  14426=>"111000010",
  14427=>"110001000",
  14428=>"101011111",
  14429=>"001111000",
  14430=>"000100001",
  14431=>"111011101",
  14432=>"001000101",
  14433=>"101100010",
  14434=>"111011111",
  14435=>"001001101",
  14436=>"101100010",
  14437=>"100001000",
  14438=>"110101101",
  14439=>"000111111",
  14440=>"001000010",
  14441=>"001111001",
  14442=>"111101001",
  14443=>"101101110",
  14444=>"100010011",
  14445=>"110001000",
  14446=>"010010101",
  14447=>"000100001",
  14448=>"110001010",
  14449=>"001000100",
  14450=>"011111101",
  14451=>"000001000",
  14452=>"011100111",
  14453=>"001011010",
  14454=>"000010010",
  14455=>"001101111",
  14456=>"101000010",
  14457=>"111011111",
  14458=>"100000010",
  14459=>"111100110",
  14460=>"011011111",
  14461=>"111011010",
  14462=>"101010000",
  14463=>"000010001",
  14464=>"011000001",
  14465=>"001011110",
  14466=>"001110100",
  14467=>"000101100",
  14468=>"100100101",
  14469=>"101010000",
  14470=>"100100101",
  14471=>"110010011",
  14472=>"101000111",
  14473=>"101100010",
  14474=>"010010110",
  14475=>"001111101",
  14476=>"110100100",
  14477=>"000110001",
  14478=>"110001011",
  14479=>"111111101",
  14480=>"010001111",
  14481=>"111100000",
  14482=>"000110101",
  14483=>"001000011",
  14484=>"100001100",
  14485=>"010111110",
  14486=>"100111101",
  14487=>"000011001",
  14488=>"110111011",
  14489=>"111101001",
  14490=>"111110000",
  14491=>"000100000",
  14492=>"101111110",
  14493=>"010010101",
  14494=>"101100001",
  14495=>"011010110",
  14496=>"000000011",
  14497=>"000001000",
  14498=>"001100100",
  14499=>"110110011",
  14500=>"100111011",
  14501=>"111000100",
  14502=>"010010011",
  14503=>"111001100",
  14504=>"001001001",
  14505=>"001001001",
  14506=>"101110100",
  14507=>"111111000",
  14508=>"100000000",
  14509=>"001110000",
  14510=>"000110100",
  14511=>"100100000",
  14512=>"110010110",
  14513=>"000011111",
  14514=>"000001011",
  14515=>"101110110",
  14516=>"111110100",
  14517=>"110001001",
  14518=>"011101010",
  14519=>"101100100",
  14520=>"010000110",
  14521=>"000100111",
  14522=>"000000011",
  14523=>"111001010",
  14524=>"101001101",
  14525=>"111111001",
  14526=>"011101101",
  14527=>"111101110",
  14528=>"001001110",
  14529=>"010011100",
  14530=>"000111011",
  14531=>"000011111",
  14532=>"001010010",
  14533=>"001101011",
  14534=>"000010110",
  14535=>"001000100",
  14536=>"001100010",
  14537=>"001100000",
  14538=>"100101000",
  14539=>"011011101",
  14540=>"001111111",
  14541=>"110000011",
  14542=>"010011010",
  14543=>"010101111",
  14544=>"100001000",
  14545=>"000001010",
  14546=>"100000000",
  14547=>"000100100",
  14548=>"111111111",
  14549=>"100000101",
  14550=>"110100110",
  14551=>"011100000",
  14552=>"000110101",
  14553=>"011100101",
  14554=>"000100100",
  14555=>"100111001",
  14556=>"001111011",
  14557=>"010010111",
  14558=>"100001011",
  14559=>"110101110",
  14560=>"111110000",
  14561=>"011010100",
  14562=>"001101010",
  14563=>"110101110",
  14564=>"100110111",
  14565=>"011100110",
  14566=>"000011111",
  14567=>"010000011",
  14568=>"010011001",
  14569=>"011001011",
  14570=>"101101010",
  14571=>"011101000",
  14572=>"101100010",
  14573=>"000100111",
  14574=>"010100001",
  14575=>"010001100",
  14576=>"011011001",
  14577=>"011001110",
  14578=>"101000111",
  14579=>"011000011",
  14580=>"100110101",
  14581=>"010110001",
  14582=>"110111101",
  14583=>"101001101",
  14584=>"011100000",
  14585=>"111011111",
  14586=>"011001100",
  14587=>"000001000",
  14588=>"110000011",
  14589=>"100100111",
  14590=>"001011001",
  14591=>"000100001",
  14592=>"010111001",
  14593=>"010000111",
  14594=>"000010000",
  14595=>"111011110",
  14596=>"000001000",
  14597=>"001000001",
  14598=>"101010001",
  14599=>"111111100",
  14600=>"101011110",
  14601=>"001010000",
  14602=>"101010001",
  14603=>"011100011",
  14604=>"000011111",
  14605=>"001010000",
  14606=>"011110101",
  14607=>"100111000",
  14608=>"101111001",
  14609=>"100101101",
  14610=>"100101010",
  14611=>"001101111",
  14612=>"100011000",
  14613=>"101101100",
  14614=>"001100100",
  14615=>"011001011",
  14616=>"010010101",
  14617=>"001111000",
  14618=>"100101010",
  14619=>"010101001",
  14620=>"000010100",
  14621=>"111010000",
  14622=>"111101101",
  14623=>"100010111",
  14624=>"000000011",
  14625=>"010100100",
  14626=>"110010100",
  14627=>"001000011",
  14628=>"100000001",
  14629=>"011000110",
  14630=>"011001000",
  14631=>"011101000",
  14632=>"010100011",
  14633=>"011110010",
  14634=>"111101001",
  14635=>"000010110",
  14636=>"100101111",
  14637=>"110110100",
  14638=>"001000111",
  14639=>"100001111",
  14640=>"000101000",
  14641=>"001111010",
  14642=>"001011101",
  14643=>"001011000",
  14644=>"001011001",
  14645=>"010000010",
  14646=>"110101110",
  14647=>"010011001",
  14648=>"001000000",
  14649=>"110111010",
  14650=>"101100001",
  14651=>"110010001",
  14652=>"110000011",
  14653=>"100101011",
  14654=>"011110101",
  14655=>"001000101",
  14656=>"110111001",
  14657=>"011101011",
  14658=>"101000110",
  14659=>"101001100",
  14660=>"010010011",
  14661=>"101011010",
  14662=>"011110100",
  14663=>"010001111",
  14664=>"011101010",
  14665=>"111000010",
  14666=>"001010011",
  14667=>"011010000",
  14668=>"110010110",
  14669=>"011110001",
  14670=>"111001000",
  14671=>"011110011",
  14672=>"010000110",
  14673=>"001000100",
  14674=>"100110101",
  14675=>"000110000",
  14676=>"111101111",
  14677=>"101100001",
  14678=>"010111011",
  14679=>"101101001",
  14680=>"001010010",
  14681=>"001110000",
  14682=>"010101000",
  14683=>"001010000",
  14684=>"001010000",
  14685=>"111111101",
  14686=>"110001100",
  14687=>"000001110",
  14688=>"000101011",
  14689=>"110100100",
  14690=>"000101010",
  14691=>"000110010",
  14692=>"111100101",
  14693=>"100011000",
  14694=>"010001101",
  14695=>"101101110",
  14696=>"110000100",
  14697=>"101001010",
  14698=>"100000000",
  14699=>"010011010",
  14700=>"110010011",
  14701=>"101110101",
  14702=>"011111110",
  14703=>"100101110",
  14704=>"000000000",
  14705=>"111001111",
  14706=>"010101111",
  14707=>"110101111",
  14708=>"111111010",
  14709=>"010111100",
  14710=>"111001110",
  14711=>"001101100",
  14712=>"111110101",
  14713=>"111101111",
  14714=>"111101000",
  14715=>"100111010",
  14716=>"111000011",
  14717=>"111101110",
  14718=>"111110110",
  14719=>"100000000",
  14720=>"111111101",
  14721=>"100110011",
  14722=>"111011011",
  14723=>"111110110",
  14724=>"100001100",
  14725=>"101000001",
  14726=>"010010001",
  14727=>"110000111",
  14728=>"101010100",
  14729=>"000010101",
  14730=>"110011001",
  14731=>"110111100",
  14732=>"001111011",
  14733=>"000010010",
  14734=>"001000000",
  14735=>"001111111",
  14736=>"101111110",
  14737=>"000000011",
  14738=>"000100111",
  14739=>"110101000",
  14740=>"010101010",
  14741=>"011100001",
  14742=>"011100101",
  14743=>"011011001",
  14744=>"110000110",
  14745=>"001100001",
  14746=>"001100111",
  14747=>"000110010",
  14748=>"010100001",
  14749=>"000011010",
  14750=>"000000100",
  14751=>"110101000",
  14752=>"000101000",
  14753=>"000111101",
  14754=>"111111111",
  14755=>"110001010",
  14756=>"000111000",
  14757=>"011010010",
  14758=>"010111010",
  14759=>"011101110",
  14760=>"111110011",
  14761=>"110000011",
  14762=>"000000111",
  14763=>"000011101",
  14764=>"000110110",
  14765=>"100000010",
  14766=>"000000010",
  14767=>"010011010",
  14768=>"000100110",
  14769=>"011101100",
  14770=>"111011111",
  14771=>"011100100",
  14772=>"001101110",
  14773=>"000101101",
  14774=>"000000111",
  14775=>"111011000",
  14776=>"101111001",
  14777=>"000101101",
  14778=>"001000000",
  14779=>"001011111",
  14780=>"110110111",
  14781=>"100000000",
  14782=>"111111101",
  14783=>"000010110",
  14784=>"101100110",
  14785=>"011101010",
  14786=>"100011110",
  14787=>"000101011",
  14788=>"111010111",
  14789=>"110000110",
  14790=>"001110100",
  14791=>"000010000",
  14792=>"001100011",
  14793=>"101110100",
  14794=>"100000100",
  14795=>"101010100",
  14796=>"101100101",
  14797=>"011011101",
  14798=>"001111100",
  14799=>"111101100",
  14800=>"100000011",
  14801=>"000100110",
  14802=>"000101010",
  14803=>"010101111",
  14804=>"110001110",
  14805=>"101110000",
  14806=>"100100010",
  14807=>"100010100",
  14808=>"011110111",
  14809=>"111001000",
  14810=>"011110111",
  14811=>"010000100",
  14812=>"111000011",
  14813=>"100111100",
  14814=>"000000000",
  14815=>"101001111",
  14816=>"100000011",
  14817=>"111000000",
  14818=>"111101110",
  14819=>"000100111",
  14820=>"111110100",
  14821=>"001000111",
  14822=>"011001010",
  14823=>"101011101",
  14824=>"010001111",
  14825=>"000000110",
  14826=>"001101001",
  14827=>"000000000",
  14828=>"000101101",
  14829=>"011000000",
  14830=>"000111001",
  14831=>"010110001",
  14832=>"101111010",
  14833=>"000101011",
  14834=>"101110000",
  14835=>"111001010",
  14836=>"100010000",
  14837=>"000101000",
  14838=>"101110101",
  14839=>"000001001",
  14840=>"110111110",
  14841=>"000100010",
  14842=>"100000101",
  14843=>"001011000",
  14844=>"001011111",
  14845=>"101010111",
  14846=>"110110101",
  14847=>"010000000",
  14848=>"011111111",
  14849=>"100111101",
  14850=>"100101010",
  14851=>"111010110",
  14852=>"110011000",
  14853=>"011101100",
  14854=>"111111011",
  14855=>"010000001",
  14856=>"010001100",
  14857=>"000110011",
  14858=>"101100000",
  14859=>"000001000",
  14860=>"000110000",
  14861=>"001100010",
  14862=>"101000111",
  14863=>"111111101",
  14864=>"100110101",
  14865=>"101101100",
  14866=>"101010000",
  14867=>"001001001",
  14868=>"010010100",
  14869=>"101110000",
  14870=>"011111011",
  14871=>"011101101",
  14872=>"001011001",
  14873=>"111101001",
  14874=>"110110011",
  14875=>"011011001",
  14876=>"010000011",
  14877=>"101110101",
  14878=>"111110111",
  14879=>"010001100",
  14880=>"010000011",
  14881=>"010111001",
  14882=>"010001111",
  14883=>"010011011",
  14884=>"011111010",
  14885=>"100110110",
  14886=>"000000101",
  14887=>"110011011",
  14888=>"111111000",
  14889=>"010101011",
  14890=>"010100010",
  14891=>"001011110",
  14892=>"111001101",
  14893=>"001100001",
  14894=>"000110010",
  14895=>"010000000",
  14896=>"111110010",
  14897=>"101100111",
  14898=>"011010001",
  14899=>"100011000",
  14900=>"011110000",
  14901=>"000001011",
  14902=>"101111101",
  14903=>"101111000",
  14904=>"100010000",
  14905=>"011101111",
  14906=>"010111100",
  14907=>"011110011",
  14908=>"100111001",
  14909=>"110000001",
  14910=>"010111001",
  14911=>"111001001",
  14912=>"010101110",
  14913=>"000010001",
  14914=>"010001000",
  14915=>"110011010",
  14916=>"001010101",
  14917=>"110111100",
  14918=>"111000100",
  14919=>"100110111",
  14920=>"110001101",
  14921=>"001010101",
  14922=>"001100110",
  14923=>"101000110",
  14924=>"100000010",
  14925=>"111101010",
  14926=>"001010111",
  14927=>"001000001",
  14928=>"111101111",
  14929=>"010001010",
  14930=>"100001001",
  14931=>"010011101",
  14932=>"010101001",
  14933=>"111000001",
  14934=>"001011010",
  14935=>"011010111",
  14936=>"001010110",
  14937=>"001110100",
  14938=>"110100000",
  14939=>"101011001",
  14940=>"001001011",
  14941=>"110000100",
  14942=>"110111111",
  14943=>"101111001",
  14944=>"001001000",
  14945=>"000100011",
  14946=>"011101110",
  14947=>"011010110",
  14948=>"001110000",
  14949=>"010001010",
  14950=>"001111101",
  14951=>"110101111",
  14952=>"000100010",
  14953=>"111010010",
  14954=>"100110001",
  14955=>"110000001",
  14956=>"101001010",
  14957=>"010010101",
  14958=>"101011000",
  14959=>"011000111",
  14960=>"010100101",
  14961=>"101111011",
  14962=>"001010011",
  14963=>"011001001",
  14964=>"010110001",
  14965=>"010000001",
  14966=>"001010111",
  14967=>"001011011",
  14968=>"100000010",
  14969=>"001000110",
  14970=>"010000100",
  14971=>"111001010",
  14972=>"010100000",
  14973=>"000011100",
  14974=>"000110010",
  14975=>"001011000",
  14976=>"111111101",
  14977=>"101111101",
  14978=>"101101111",
  14979=>"001010110",
  14980=>"111001001",
  14981=>"011010000",
  14982=>"100000010",
  14983=>"010001010",
  14984=>"100000010",
  14985=>"011011101",
  14986=>"101101111",
  14987=>"000000100",
  14988=>"011001001",
  14989=>"001000001",
  14990=>"101011001",
  14991=>"110011100",
  14992=>"000101010",
  14993=>"110111011",
  14994=>"011110000",
  14995=>"100010001",
  14996=>"000000101",
  14997=>"010111010",
  14998=>"000101110",
  14999=>"000100001",
  15000=>"000001101",
  15001=>"010110010",
  15002=>"001010110",
  15003=>"011111111",
  15004=>"111001011",
  15005=>"101100111",
  15006=>"000110101",
  15007=>"101000110",
  15008=>"011101000",
  15009=>"101000010",
  15010=>"111101000",
  15011=>"101111110",
  15012=>"010011001",
  15013=>"111100001",
  15014=>"001000001",
  15015=>"010000101",
  15016=>"000011001",
  15017=>"100010000",
  15018=>"000100010",
  15019=>"011001001",
  15020=>"110111111",
  15021=>"001001101",
  15022=>"110111111",
  15023=>"011000011",
  15024=>"000110101",
  15025=>"000011111",
  15026=>"000111011",
  15027=>"000101101",
  15028=>"010010010",
  15029=>"111000011",
  15030=>"100011101",
  15031=>"110110111",
  15032=>"100100110",
  15033=>"011001010",
  15034=>"011110000",
  15035=>"010110011",
  15036=>"000101010",
  15037=>"100101101",
  15038=>"000100111",
  15039=>"000101101",
  15040=>"000100011",
  15041=>"111001110",
  15042=>"110000000",
  15043=>"111010110",
  15044=>"000100011",
  15045=>"001010111",
  15046=>"101001110",
  15047=>"110111111",
  15048=>"001010100",
  15049=>"111000001",
  15050=>"101100010",
  15051=>"011110011",
  15052=>"100001100",
  15053=>"111001111",
  15054=>"001000000",
  15055=>"110111111",
  15056=>"111110001",
  15057=>"001000110",
  15058=>"001011100",
  15059=>"010101100",
  15060=>"011111110",
  15061=>"001111111",
  15062=>"001001000",
  15063=>"001101000",
  15064=>"101100010",
  15065=>"111010000",
  15066=>"011100110",
  15067=>"110011111",
  15068=>"001101000",
  15069=>"001001011",
  15070=>"001101001",
  15071=>"100110111",
  15072=>"000001100",
  15073=>"111100001",
  15074=>"001100101",
  15075=>"000110111",
  15076=>"101101111",
  15077=>"100100010",
  15078=>"011001000",
  15079=>"111011000",
  15080=>"010111011",
  15081=>"011100010",
  15082=>"100100001",
  15083=>"011010000",
  15084=>"101101110",
  15085=>"111010000",
  15086=>"010110101",
  15087=>"000101111",
  15088=>"111010101",
  15089=>"011011110",
  15090=>"001010010",
  15091=>"010000000",
  15092=>"110110111",
  15093=>"001010000",
  15094=>"000100101",
  15095=>"110111000",
  15096=>"100001000",
  15097=>"110000010",
  15098=>"011001010",
  15099=>"001011011",
  15100=>"100011011",
  15101=>"001010111",
  15102=>"010111000",
  15103=>"110110100",
  15104=>"111000010",
  15105=>"010100001",
  15106=>"110010101",
  15107=>"100100100",
  15108=>"110000110",
  15109=>"101000100",
  15110=>"110111111",
  15111=>"000101010",
  15112=>"000110011",
  15113=>"100101001",
  15114=>"000101000",
  15115=>"001010000",
  15116=>"111000000",
  15117=>"011011011",
  15118=>"000101010",
  15119=>"110101010",
  15120=>"001111010",
  15121=>"000010001",
  15122=>"111000100",
  15123=>"001111100",
  15124=>"111011011",
  15125=>"111110001",
  15126=>"011010011",
  15127=>"000001000",
  15128=>"011011000",
  15129=>"100000000",
  15130=>"001111000",
  15131=>"101101010",
  15132=>"101111011",
  15133=>"101100001",
  15134=>"101111011",
  15135=>"010100101",
  15136=>"101010111",
  15137=>"100000000",
  15138=>"101110111",
  15139=>"000000000",
  15140=>"011011010",
  15141=>"010101000",
  15142=>"110001000",
  15143=>"101101001",
  15144=>"111111000",
  15145=>"111010000",
  15146=>"010101111",
  15147=>"110010010",
  15148=>"011110100",
  15149=>"001110011",
  15150=>"000000001",
  15151=>"011001011",
  15152=>"000111101",
  15153=>"111000111",
  15154=>"110101101",
  15155=>"001110000",
  15156=>"111100111",
  15157=>"010110001",
  15158=>"111101010",
  15159=>"001100001",
  15160=>"000111000",
  15161=>"111101111",
  15162=>"010100101",
  15163=>"110001100",
  15164=>"101101100",
  15165=>"011000100",
  15166=>"101100011",
  15167=>"100100101",
  15168=>"010011000",
  15169=>"110111001",
  15170=>"111100100",
  15171=>"010101101",
  15172=>"111001010",
  15173=>"000000111",
  15174=>"101100101",
  15175=>"101001001",
  15176=>"111111001",
  15177=>"011111010",
  15178=>"100011001",
  15179=>"101001110",
  15180=>"111101000",
  15181=>"011111001",
  15182=>"000010001",
  15183=>"000110011",
  15184=>"101000100",
  15185=>"100110100",
  15186=>"011111100",
  15187=>"110000111",
  15188=>"101111001",
  15189=>"010111010",
  15190=>"001110101",
  15191=>"100111011",
  15192=>"010000010",
  15193=>"111001110",
  15194=>"111000100",
  15195=>"101110111",
  15196=>"111110000",
  15197=>"101010100",
  15198=>"100111110",
  15199=>"001101001",
  15200=>"110100010",
  15201=>"101111111",
  15202=>"000111001",
  15203=>"111111000",
  15204=>"011101011",
  15205=>"110100101",
  15206=>"010100101",
  15207=>"100111101",
  15208=>"011011000",
  15209=>"110000101",
  15210=>"110001101",
  15211=>"110001100",
  15212=>"010010100",
  15213=>"001001111",
  15214=>"001001000",
  15215=>"010110000",
  15216=>"110001000",
  15217=>"110101011",
  15218=>"100011001",
  15219=>"111101111",
  15220=>"101110100",
  15221=>"111000001",
  15222=>"010011110",
  15223=>"001011111",
  15224=>"100001011",
  15225=>"001011000",
  15226=>"101100100",
  15227=>"111110010",
  15228=>"111001100",
  15229=>"101001001",
  15230=>"000011010",
  15231=>"000000010",
  15232=>"100101011",
  15233=>"110100010",
  15234=>"111001001",
  15235=>"000000111",
  15236=>"100110110",
  15237=>"000011001",
  15238=>"000001101",
  15239=>"101011011",
  15240=>"101101111",
  15241=>"110011000",
  15242=>"011011110",
  15243=>"111011110",
  15244=>"101010000",
  15245=>"110111000",
  15246=>"101111110",
  15247=>"011011110",
  15248=>"000001001",
  15249=>"010110111",
  15250=>"000000111",
  15251=>"111010010",
  15252=>"000000011",
  15253=>"001111110",
  15254=>"111011111",
  15255=>"000001001",
  15256=>"001100110",
  15257=>"101101110",
  15258=>"001011000",
  15259=>"000010011",
  15260=>"111110001",
  15261=>"101101100",
  15262=>"110101100",
  15263=>"000011100",
  15264=>"001100000",
  15265=>"101010000",
  15266=>"001011101",
  15267=>"100000101",
  15268=>"000101110",
  15269=>"001001011",
  15270=>"011100111",
  15271=>"011011100",
  15272=>"001000110",
  15273=>"000001000",
  15274=>"011101111",
  15275=>"011011011",
  15276=>"001111100",
  15277=>"000110110",
  15278=>"000111101",
  15279=>"001010001",
  15280=>"110011000",
  15281=>"000110011",
  15282=>"001100011",
  15283=>"010010111",
  15284=>"011100111",
  15285=>"000001010",
  15286=>"001011011",
  15287=>"100001011",
  15288=>"011011111",
  15289=>"011011010",
  15290=>"101110110",
  15291=>"001100000",
  15292=>"111011110",
  15293=>"101010011",
  15294=>"011011010",
  15295=>"100111010",
  15296=>"010110100",
  15297=>"101100010",
  15298=>"100111111",
  15299=>"101010100",
  15300=>"000100111",
  15301=>"000011100",
  15302=>"010100110",
  15303=>"011010000",
  15304=>"011110001",
  15305=>"110011110",
  15306=>"100000000",
  15307=>"010100001",
  15308=>"111101110",
  15309=>"001100000",
  15310=>"010110100",
  15311=>"110101010",
  15312=>"001111110",
  15313=>"110000101",
  15314=>"100101111",
  15315=>"001100001",
  15316=>"000110000",
  15317=>"010000100",
  15318=>"011010111",
  15319=>"011010000",
  15320=>"100111000",
  15321=>"011010011",
  15322=>"000000000",
  15323=>"111110110",
  15324=>"110111001",
  15325=>"111010101",
  15326=>"011110101",
  15327=>"110001101",
  15328=>"000000100",
  15329=>"100001011",
  15330=>"101001100",
  15331=>"010001100",
  15332=>"011000101",
  15333=>"111000001",
  15334=>"100111010",
  15335=>"010000011",
  15336=>"001100101",
  15337=>"111100111",
  15338=>"100101100",
  15339=>"000110111",
  15340=>"101000011",
  15341=>"111100001",
  15342=>"001001010",
  15343=>"000100111",
  15344=>"111000101",
  15345=>"001111101",
  15346=>"011110100",
  15347=>"000100000",
  15348=>"000110111",
  15349=>"100111111",
  15350=>"000100000",
  15351=>"011110011",
  15352=>"000000010",
  15353=>"000111010",
  15354=>"101100010",
  15355=>"011100011",
  15356=>"111110010",
  15357=>"110010000",
  15358=>"110000010",
  15359=>"011010101",
  15360=>"000000000",
  15361=>"111111111",
  15362=>"011000010",
  15363=>"000010110",
  15364=>"001000000",
  15365=>"101010001",
  15366=>"100000010",
  15367=>"110011101",
  15368=>"011000010",
  15369=>"010001010",
  15370=>"111100010",
  15371=>"110011001",
  15372=>"101110111",
  15373=>"000010010",
  15374=>"110101110",
  15375=>"011000001",
  15376=>"011001100",
  15377=>"100001010",
  15378=>"011101110",
  15379=>"110100011",
  15380=>"000011100",
  15381=>"011111111",
  15382=>"001101110",
  15383=>"001101001",
  15384=>"000011001",
  15385=>"110100110",
  15386=>"010010000",
  15387=>"011011101",
  15388=>"111100101",
  15389=>"111000110",
  15390=>"100000100",
  15391=>"100001010",
  15392=>"110101010",
  15393=>"001001110",
  15394=>"011000111",
  15395=>"000101111",
  15396=>"110100111",
  15397=>"111110001",
  15398=>"011111011",
  15399=>"001111010",
  15400=>"111101100",
  15401=>"110011111",
  15402=>"100101001",
  15403=>"100101100",
  15404=>"010001001",
  15405=>"100111100",
  15406=>"000100001",
  15407=>"110000111",
  15408=>"100101010",
  15409=>"101010011",
  15410=>"111111111",
  15411=>"111101111",
  15412=>"010100011",
  15413=>"111010001",
  15414=>"111110010",
  15415=>"101110110",
  15416=>"011001111",
  15417=>"010000101",
  15418=>"000001011",
  15419=>"000101100",
  15420=>"010001000",
  15421=>"110111001",
  15422=>"001110011",
  15423=>"111101101",
  15424=>"011111010",
  15425=>"110011011",
  15426=>"001010000",
  15427=>"101110110",
  15428=>"011111001",
  15429=>"110110001",
  15430=>"000101110",
  15431=>"001110000",
  15432=>"000101101",
  15433=>"000000010",
  15434=>"110001110",
  15435=>"000001110",
  15436=>"010000001",
  15437=>"111111011",
  15438=>"111111001",
  15439=>"011000111",
  15440=>"111001000",
  15441=>"110101001",
  15442=>"100101110",
  15443=>"100010000",
  15444=>"101001011",
  15445=>"111110111",
  15446=>"101101001",
  15447=>"110010110",
  15448=>"010011001",
  15449=>"110100001",
  15450=>"010000001",
  15451=>"110000011",
  15452=>"011101000",
  15453=>"110001000",
  15454=>"110001101",
  15455=>"010110101",
  15456=>"011101011",
  15457=>"001000111",
  15458=>"001100000",
  15459=>"011101100",
  15460=>"110000010",
  15461=>"000000001",
  15462=>"110011010",
  15463=>"111001000",
  15464=>"001010001",
  15465=>"000011001",
  15466=>"000101001",
  15467=>"000011111",
  15468=>"011101111",
  15469=>"001000010",
  15470=>"000001000",
  15471=>"000110111",
  15472=>"000011001",
  15473=>"001011110",
  15474=>"001101110",
  15475=>"000001101",
  15476=>"011100101",
  15477=>"101100111",
  15478=>"011100100",
  15479=>"111110110",
  15480=>"001101000",
  15481=>"110100001",
  15482=>"001100010",
  15483=>"010101101",
  15484=>"101001011",
  15485=>"010100011",
  15486=>"101010111",
  15487=>"010100101",
  15488=>"010000111",
  15489=>"001101001",
  15490=>"010000101",
  15491=>"011001101",
  15492=>"101100010",
  15493=>"001110000",
  15494=>"001101111",
  15495=>"100000000",
  15496=>"011101010",
  15497=>"100010011",
  15498=>"101101101",
  15499=>"011110000",
  15500=>"100100010",
  15501=>"110101010",
  15502=>"110100010",
  15503=>"111010011",
  15504=>"101010000",
  15505=>"000000100",
  15506=>"010000101",
  15507=>"000001001",
  15508=>"001010100",
  15509=>"111010000",
  15510=>"101101110",
  15511=>"010100110",
  15512=>"001100000",
  15513=>"101011101",
  15514=>"100100000",
  15515=>"111010011",
  15516=>"000101000",
  15517=>"101011110",
  15518=>"010010010",
  15519=>"000011010",
  15520=>"000010100",
  15521=>"111111010",
  15522=>"110101001",
  15523=>"010010000",
  15524=>"100110111",
  15525=>"010100110",
  15526=>"010111001",
  15527=>"110100001",
  15528=>"000111000",
  15529=>"001010110",
  15530=>"110111111",
  15531=>"111111111",
  15532=>"111110100",
  15533=>"110000000",
  15534=>"100011001",
  15535=>"100010010",
  15536=>"111110010",
  15537=>"000110111",
  15538=>"000010100",
  15539=>"100011010",
  15540=>"110000010",
  15541=>"001010001",
  15542=>"011110010",
  15543=>"110001000",
  15544=>"111100100",
  15545=>"110100101",
  15546=>"100001011",
  15547=>"000011011",
  15548=>"100000011",
  15549=>"111011111",
  15550=>"010000010",
  15551=>"111100000",
  15552=>"110001110",
  15553=>"101011011",
  15554=>"000101000",
  15555=>"011000111",
  15556=>"010011110",
  15557=>"101011111",
  15558=>"010100011",
  15559=>"101110011",
  15560=>"011001001",
  15561=>"100010101",
  15562=>"011100001",
  15563=>"100100110",
  15564=>"001010100",
  15565=>"101011100",
  15566=>"110110011",
  15567=>"111001101",
  15568=>"001011100",
  15569=>"101000010",
  15570=>"101110110",
  15571=>"011000110",
  15572=>"110010110",
  15573=>"110110110",
  15574=>"000010011",
  15575=>"010000101",
  15576=>"001101000",
  15577=>"010110101",
  15578=>"101010111",
  15579=>"010000110",
  15580=>"010000001",
  15581=>"010010101",
  15582=>"001101101",
  15583=>"010001110",
  15584=>"111110010",
  15585=>"011011011",
  15586=>"100010001",
  15587=>"100111010",
  15588=>"010000010",
  15589=>"111110101",
  15590=>"100000010",
  15591=>"101001110",
  15592=>"111110100",
  15593=>"110100011",
  15594=>"010011010",
  15595=>"101101001",
  15596=>"101111011",
  15597=>"111010101",
  15598=>"001000011",
  15599=>"001101001",
  15600=>"101110000",
  15601=>"111101000",
  15602=>"110000111",
  15603=>"000011111",
  15604=>"101101111",
  15605=>"111110110",
  15606=>"000010011",
  15607=>"011101001",
  15608=>"011000101",
  15609=>"111000001",
  15610=>"011011001",
  15611=>"110100001",
  15612=>"011011101",
  15613=>"010101000",
  15614=>"001000001",
  15615=>"101101111",
  15616=>"001000000",
  15617=>"010010111",
  15618=>"000110111",
  15619=>"110101100",
  15620=>"010110100",
  15621=>"000001001",
  15622=>"100110010",
  15623=>"001001000",
  15624=>"010000101",
  15625=>"010011110",
  15626=>"101110101",
  15627=>"000110010",
  15628=>"111111001",
  15629=>"100000011",
  15630=>"011011001",
  15631=>"011100100",
  15632=>"000011011",
  15633=>"010100011",
  15634=>"001010100",
  15635=>"101101101",
  15636=>"000011111",
  15637=>"000000011",
  15638=>"000100001",
  15639=>"100011110",
  15640=>"100010001",
  15641=>"101110001",
  15642=>"010010010",
  15643=>"011100100",
  15644=>"011001101",
  15645=>"000111000",
  15646=>"000011011",
  15647=>"010111010",
  15648=>"010000100",
  15649=>"000101111",
  15650=>"100110101",
  15651=>"001001100",
  15652=>"010000001",
  15653=>"001111011",
  15654=>"011010000",
  15655=>"000000110",
  15656=>"001101000",
  15657=>"110000010",
  15658=>"011100010",
  15659=>"001101000",
  15660=>"001110100",
  15661=>"000110000",
  15662=>"101111110",
  15663=>"101111001",
  15664=>"001100001",
  15665=>"010010110",
  15666=>"101010101",
  15667=>"010100111",
  15668=>"100110011",
  15669=>"110000000",
  15670=>"001001001",
  15671=>"000011100",
  15672=>"110001010",
  15673=>"111101111",
  15674=>"011110111",
  15675=>"000001100",
  15676=>"111101101",
  15677=>"101001001",
  15678=>"011100110",
  15679=>"111101100",
  15680=>"111101101",
  15681=>"100000100",
  15682=>"110101101",
  15683=>"101011101",
  15684=>"000011100",
  15685=>"011100000",
  15686=>"100011010",
  15687=>"111101001",
  15688=>"000111110",
  15689=>"110001110",
  15690=>"000110110",
  15691=>"110010000",
  15692=>"010011100",
  15693=>"011111001",
  15694=>"010001111",
  15695=>"000000011",
  15696=>"001001000",
  15697=>"001100111",
  15698=>"100010010",
  15699=>"110110111",
  15700=>"000100011",
  15701=>"110011000",
  15702=>"100001010",
  15703=>"011100100",
  15704=>"101011000",
  15705=>"011000110",
  15706=>"000011001",
  15707=>"001010000",
  15708=>"010111000",
  15709=>"011011100",
  15710=>"001011111",
  15711=>"101000011",
  15712=>"101111101",
  15713=>"011100101",
  15714=>"010010000",
  15715=>"000000001",
  15716=>"111111111",
  15717=>"100110100",
  15718=>"100011001",
  15719=>"001110100",
  15720=>"001010110",
  15721=>"010100110",
  15722=>"010100100",
  15723=>"011001001",
  15724=>"100101100",
  15725=>"001011011",
  15726=>"111111011",
  15727=>"100010101",
  15728=>"111110000",
  15729=>"011100101",
  15730=>"001101111",
  15731=>"001111110",
  15732=>"000101010",
  15733=>"100010001",
  15734=>"010111001",
  15735=>"000011110",
  15736=>"111101011",
  15737=>"101100000",
  15738=>"111110010",
  15739=>"110111110",
  15740=>"010110101",
  15741=>"101000111",
  15742=>"011001100",
  15743=>"010111111",
  15744=>"111111010",
  15745=>"111101101",
  15746=>"001101100",
  15747=>"111011100",
  15748=>"110110101",
  15749=>"110001010",
  15750=>"110010100",
  15751=>"110010111",
  15752=>"101000101",
  15753=>"111111010",
  15754=>"010101101",
  15755=>"010111110",
  15756=>"010000001",
  15757=>"100011100",
  15758=>"110110101",
  15759=>"101111011",
  15760=>"000000010",
  15761=>"011001110",
  15762=>"110101100",
  15763=>"000110110",
  15764=>"001100010",
  15765=>"000110000",
  15766=>"100001000",
  15767=>"000111001",
  15768=>"111000001",
  15769=>"000100000",
  15770=>"100011100",
  15771=>"011000101",
  15772=>"011100110",
  15773=>"001010100",
  15774=>"101100101",
  15775=>"100000111",
  15776=>"011110100",
  15777=>"101011110",
  15778=>"100010000",
  15779=>"100100011",
  15780=>"100101010",
  15781=>"000000110",
  15782=>"011101110",
  15783=>"000000001",
  15784=>"100011111",
  15785=>"000000010",
  15786=>"010010011",
  15787=>"101010101",
  15788=>"010011101",
  15789=>"001101110",
  15790=>"000111101",
  15791=>"101001111",
  15792=>"000000001",
  15793=>"111111111",
  15794=>"111000111",
  15795=>"110000001",
  15796=>"110111001",
  15797=>"001111110",
  15798=>"001001001",
  15799=>"010011111",
  15800=>"111011101",
  15801=>"100111111",
  15802=>"010101010",
  15803=>"000100010",
  15804=>"011111011",
  15805=>"100110010",
  15806=>"110110001",
  15807=>"111000001",
  15808=>"100011111",
  15809=>"010101100",
  15810=>"001011111",
  15811=>"101111001",
  15812=>"111100011",
  15813=>"010100001",
  15814=>"101111011",
  15815=>"001011111",
  15816=>"111111001",
  15817=>"110010000",
  15818=>"010110110",
  15819=>"000000100",
  15820=>"000010001",
  15821=>"101100101",
  15822=>"111100001",
  15823=>"011000101",
  15824=>"101100001",
  15825=>"111110011",
  15826=>"101011101",
  15827=>"100101111",
  15828=>"000111001",
  15829=>"111001001",
  15830=>"101101001",
  15831=>"100100111",
  15832=>"110000010",
  15833=>"111010001",
  15834=>"111001101",
  15835=>"110110001",
  15836=>"001100011",
  15837=>"110111011",
  15838=>"011111110",
  15839=>"110111101",
  15840=>"111110101",
  15841=>"001101100",
  15842=>"011111101",
  15843=>"001001111",
  15844=>"001011000",
  15845=>"101110010",
  15846=>"110000000",
  15847=>"110001100",
  15848=>"100001111",
  15849=>"000000000",
  15850=>"111001011",
  15851=>"111000110",
  15852=>"110011111",
  15853=>"100111001",
  15854=>"100001100",
  15855=>"000011000",
  15856=>"011010000",
  15857=>"110000001",
  15858=>"000000110",
  15859=>"010000001",
  15860=>"110101100",
  15861=>"100100100",
  15862=>"000101011",
  15863=>"100000000",
  15864=>"011001000",
  15865=>"001110100",
  15866=>"001001101",
  15867=>"110001110",
  15868=>"000100100",
  15869=>"110001101",
  15870=>"000010001",
  15871=>"100111111",
  15872=>"011001000",
  15873=>"001101101",
  15874=>"101101111",
  15875=>"101000010",
  15876=>"001010110",
  15877=>"000001111",
  15878=>"111010101",
  15879=>"111011110",
  15880=>"101010110",
  15881=>"110000011",
  15882=>"000011110",
  15883=>"110011001",
  15884=>"011000011",
  15885=>"110100100",
  15886=>"010101001",
  15887=>"111101001",
  15888=>"011001011",
  15889=>"010101100",
  15890=>"000000101",
  15891=>"011000101",
  15892=>"001000011",
  15893=>"111110010",
  15894=>"011100100",
  15895=>"011101100",
  15896=>"010101111",
  15897=>"000000100",
  15898=>"000100000",
  15899=>"111101000",
  15900=>"011010000",
  15901=>"100100111",
  15902=>"000010010",
  15903=>"110010111",
  15904=>"101010100",
  15905=>"100000010",
  15906=>"100100101",
  15907=>"100100000",
  15908=>"101111000",
  15909=>"111100010",
  15910=>"000100011",
  15911=>"001000001",
  15912=>"010001000",
  15913=>"001010111",
  15914=>"111010011",
  15915=>"001000011",
  15916=>"011000001",
  15917=>"000000101",
  15918=>"011101100",
  15919=>"000000110",
  15920=>"011011011",
  15921=>"110110111",
  15922=>"000100111",
  15923=>"011011100",
  15924=>"101100100",
  15925=>"001110010",
  15926=>"010011111",
  15927=>"111110001",
  15928=>"011100110",
  15929=>"011000010",
  15930=>"111111001",
  15931=>"101001111",
  15932=>"011010000",
  15933=>"101011000",
  15934=>"100010001",
  15935=>"100000001",
  15936=>"000101000",
  15937=>"000001111",
  15938=>"011111000",
  15939=>"001011111",
  15940=>"001111101",
  15941=>"011010110",
  15942=>"111101011",
  15943=>"100111100",
  15944=>"010001101",
  15945=>"101100011",
  15946=>"010110010",
  15947=>"000010010",
  15948=>"011000110",
  15949=>"101001001",
  15950=>"110111010",
  15951=>"000001001",
  15952=>"011011011",
  15953=>"100000101",
  15954=>"101101110",
  15955=>"100100011",
  15956=>"011010000",
  15957=>"101111010",
  15958=>"000000110",
  15959=>"101100010",
  15960=>"010101001",
  15961=>"011011010",
  15962=>"100100101",
  15963=>"000110110",
  15964=>"000000111",
  15965=>"101100011",
  15966=>"001010010",
  15967=>"111101110",
  15968=>"001001000",
  15969=>"101010000",
  15970=>"000111111",
  15971=>"101110100",
  15972=>"011100111",
  15973=>"110100000",
  15974=>"100110010",
  15975=>"101010111",
  15976=>"101111111",
  15977=>"010000000",
  15978=>"111100000",
  15979=>"000011100",
  15980=>"100011000",
  15981=>"111100101",
  15982=>"100000110",
  15983=>"011100111",
  15984=>"101011001",
  15985=>"100011111",
  15986=>"111001111",
  15987=>"011111110",
  15988=>"011000011",
  15989=>"111101001",
  15990=>"001000101",
  15991=>"101000011",
  15992=>"011010101",
  15993=>"100001010",
  15994=>"011001000",
  15995=>"000000001",
  15996=>"101001010",
  15997=>"000001100",
  15998=>"011100010",
  15999=>"000011111",
  16000=>"010111101",
  16001=>"110001100",
  16002=>"101001100",
  16003=>"100010110",
  16004=>"100101000",
  16005=>"000001011",
  16006=>"011110100",
  16007=>"111111101",
  16008=>"110001101",
  16009=>"100110111",
  16010=>"101101111",
  16011=>"010011111",
  16012=>"000100000",
  16013=>"111100000",
  16014=>"010100000",
  16015=>"001000110",
  16016=>"101110011",
  16017=>"001111011",
  16018=>"011111011",
  16019=>"100011111",
  16020=>"010100001",
  16021=>"100111111",
  16022=>"001110000",
  16023=>"101101110",
  16024=>"110011111",
  16025=>"100000001",
  16026=>"010010100",
  16027=>"111111100",
  16028=>"010001010",
  16029=>"011010001",
  16030=>"000111100",
  16031=>"101010101",
  16032=>"101010000",
  16033=>"011011111",
  16034=>"111001111",
  16035=>"001100010",
  16036=>"011100010",
  16037=>"001000000",
  16038=>"011110011",
  16039=>"000100000",
  16040=>"010011101",
  16041=>"001001000",
  16042=>"000000001",
  16043=>"010110000",
  16044=>"000001010",
  16045=>"100011000",
  16046=>"100110111",
  16047=>"100100011",
  16048=>"111001001",
  16049=>"011010010",
  16050=>"110101110",
  16051=>"110010110",
  16052=>"101001011",
  16053=>"111100011",
  16054=>"100110010",
  16055=>"010100000",
  16056=>"000001100",
  16057=>"001101011",
  16058=>"101110101",
  16059=>"000001111",
  16060=>"001111101",
  16061=>"111001111",
  16062=>"011000001",
  16063=>"000011111",
  16064=>"100011011",
  16065=>"011111110",
  16066=>"111001000",
  16067=>"001010001",
  16068=>"101100111",
  16069=>"000001110",
  16070=>"101111110",
  16071=>"100001000",
  16072=>"010111000",
  16073=>"001011111",
  16074=>"001111000",
  16075=>"000111110",
  16076=>"100000100",
  16077=>"111001011",
  16078=>"100000010",
  16079=>"010110010",
  16080=>"111101010",
  16081=>"001000000",
  16082=>"100100011",
  16083=>"011110101",
  16084=>"111110100",
  16085=>"111111110",
  16086=>"110101001",
  16087=>"011100100",
  16088=>"001111101",
  16089=>"010000000",
  16090=>"010100010",
  16091=>"011101011",
  16092=>"100001100",
  16093=>"111000000",
  16094=>"010011100",
  16095=>"101101110",
  16096=>"101011101",
  16097=>"101111000",
  16098=>"011010011",
  16099=>"000111000",
  16100=>"110011001",
  16101=>"111011001",
  16102=>"000110100",
  16103=>"101110101",
  16104=>"101000000",
  16105=>"100111110",
  16106=>"000110010",
  16107=>"010000100",
  16108=>"011011101",
  16109=>"011100011",
  16110=>"111100101",
  16111=>"001100111",
  16112=>"100110100",
  16113=>"101111111",
  16114=>"010011010",
  16115=>"111000011",
  16116=>"001001011",
  16117=>"101110010",
  16118=>"100011111",
  16119=>"100101011",
  16120=>"000001110",
  16121=>"100010011",
  16122=>"011011001",
  16123=>"010111011",
  16124=>"111011010",
  16125=>"101100000",
  16126=>"111100010",
  16127=>"100001100",
  16128=>"010010101",
  16129=>"011000001",
  16130=>"111101111",
  16131=>"111101101",
  16132=>"010011100",
  16133=>"001010100",
  16134=>"010101110",
  16135=>"110010000",
  16136=>"011110001",
  16137=>"100011010",
  16138=>"000011101",
  16139=>"001010000",
  16140=>"010101100",
  16141=>"101100110",
  16142=>"110011101",
  16143=>"100101100",
  16144=>"100110001",
  16145=>"111000111",
  16146=>"011000000",
  16147=>"100111010",
  16148=>"000001010",
  16149=>"000011011",
  16150=>"010111011",
  16151=>"000001010",
  16152=>"001001000",
  16153=>"000110001",
  16154=>"110000101",
  16155=>"001110101",
  16156=>"011011011",
  16157=>"011011011",
  16158=>"100011000",
  16159=>"100110111",
  16160=>"001111110",
  16161=>"010010100",
  16162=>"101010111",
  16163=>"101111000",
  16164=>"001011000",
  16165=>"110000001",
  16166=>"000111010",
  16167=>"011011101",
  16168=>"101101000",
  16169=>"101001101",
  16170=>"011111011",
  16171=>"011100000",
  16172=>"000011100",
  16173=>"110011000",
  16174=>"110111010",
  16175=>"000100000",
  16176=>"000100010",
  16177=>"111011011",
  16178=>"010000010",
  16179=>"111001101",
  16180=>"100100110",
  16181=>"010110110",
  16182=>"101001010",
  16183=>"001100000",
  16184=>"010011101",
  16185=>"111010000",
  16186=>"101000110",
  16187=>"110000110",
  16188=>"010010110",
  16189=>"000000000",
  16190=>"000100001",
  16191=>"100010111",
  16192=>"001010100",
  16193=>"101011001",
  16194=>"010000111",
  16195=>"101010001",
  16196=>"011010011",
  16197=>"111110110",
  16198=>"001010101",
  16199=>"111001010",
  16200=>"110000000",
  16201=>"010001001",
  16202=>"011111101",
  16203=>"111100011",
  16204=>"111001110",
  16205=>"011101110",
  16206=>"010000100",
  16207=>"000011000",
  16208=>"011011111",
  16209=>"001010111",
  16210=>"111010011",
  16211=>"010011001",
  16212=>"110101110",
  16213=>"001001100",
  16214=>"110110101",
  16215=>"110000010",
  16216=>"010001001",
  16217=>"100111011",
  16218=>"000000001",
  16219=>"010010101",
  16220=>"101011111",
  16221=>"011010101",
  16222=>"001001111",
  16223=>"110010000",
  16224=>"010100111",
  16225=>"101010001",
  16226=>"000001011",
  16227=>"111110111",
  16228=>"110100110",
  16229=>"000000101",
  16230=>"000010100",
  16231=>"000001000",
  16232=>"100000001",
  16233=>"010101000",
  16234=>"100111011",
  16235=>"101001000",
  16236=>"011110110",
  16237=>"101110111",
  16238=>"001011011",
  16239=>"010000101",
  16240=>"001100100",
  16241=>"101000111",
  16242=>"011011100",
  16243=>"110010001",
  16244=>"000000011",
  16245=>"001000010",
  16246=>"110100010",
  16247=>"001001010",
  16248=>"011000101",
  16249=>"000100001",
  16250=>"001111010",
  16251=>"111101101",
  16252=>"000001001",
  16253=>"100100110",
  16254=>"011111011",
  16255=>"110111111",
  16256=>"001000001",
  16257=>"100110100",
  16258=>"101000110",
  16259=>"010001110",
  16260=>"010101101",
  16261=>"011000000",
  16262=>"100101001",
  16263=>"101100101",
  16264=>"101001111",
  16265=>"110000001",
  16266=>"000011001",
  16267=>"101011010",
  16268=>"111001111",
  16269=>"111011011",
  16270=>"100111101",
  16271=>"001010000",
  16272=>"011100111",
  16273=>"101111011",
  16274=>"100110000",
  16275=>"010011110",
  16276=>"111101101",
  16277=>"101101110",
  16278=>"000001000",
  16279=>"101100101",
  16280=>"111001111",
  16281=>"111101111",
  16282=>"100110101",
  16283=>"001110001",
  16284=>"001110011",
  16285=>"001111011",
  16286=>"111011001",
  16287=>"000011011",
  16288=>"000010110",
  16289=>"110100000",
  16290=>"010011000",
  16291=>"010100100",
  16292=>"111100000",
  16293=>"111110100",
  16294=>"101000000",
  16295=>"110101000",
  16296=>"100001011",
  16297=>"111100000",
  16298=>"011111101",
  16299=>"010100010",
  16300=>"000110111",
  16301=>"000100111",
  16302=>"011001001",
  16303=>"101101000",
  16304=>"011110010",
  16305=>"010111110",
  16306=>"000011101",
  16307=>"111011111",
  16308=>"111010011",
  16309=>"011111000",
  16310=>"101110111",
  16311=>"110111001",
  16312=>"000011111",
  16313=>"001000001",
  16314=>"011001011",
  16315=>"011110100",
  16316=>"111000001",
  16317=>"001011001",
  16318=>"000111001",
  16319=>"001000000",
  16320=>"000011001",
  16321=>"111010111",
  16322=>"100000010",
  16323=>"100100010",
  16324=>"000100110",
  16325=>"101111101",
  16326=>"000100001",
  16327=>"010010100",
  16328=>"000010100",
  16329=>"111000101",
  16330=>"100111000",
  16331=>"001101101",
  16332=>"101010110",
  16333=>"001101100",
  16334=>"010100010",
  16335=>"001101010",
  16336=>"000101001",
  16337=>"110000010",
  16338=>"100110001",
  16339=>"110000110",
  16340=>"100010110",
  16341=>"000101111",
  16342=>"010111101",
  16343=>"111001100",
  16344=>"101011011",
  16345=>"111110010",
  16346=>"011001111",
  16347=>"000001000",
  16348=>"010110011",
  16349=>"011101001",
  16350=>"010111010",
  16351=>"001101000",
  16352=>"001101111",
  16353=>"010110011",
  16354=>"000001011",
  16355=>"010111110",
  16356=>"111110110",
  16357=>"101111100",
  16358=>"001011111",
  16359=>"001100010",
  16360=>"010000011",
  16361=>"000010000",
  16362=>"111100010",
  16363=>"100110101",
  16364=>"110110101",
  16365=>"000001010",
  16366=>"101010001",
  16367=>"110010110",
  16368=>"110111101",
  16369=>"101111110",
  16370=>"101110110",
  16371=>"011100010",
  16372=>"010100101",
  16373=>"010110010",
  16374=>"110111110",
  16375=>"000001000",
  16376=>"111000100",
  16377=>"011000100",
  16378=>"000100100",
  16379=>"110000111",
  16380=>"001000010",
  16381=>"100000010",
  16382=>"111100000",
  16383=>"101000110",
  16384=>"101110100",
  16385=>"001111011",
  16386=>"110110111",
  16387=>"110000110",
  16388=>"110110110",
  16389=>"010100001",
  16390=>"000011011",
  16391=>"100000011",
  16392=>"000000001",
  16393=>"001101101",
  16394=>"111010110",
  16395=>"100111010",
  16396=>"001101101",
  16397=>"101011100",
  16398=>"100000111",
  16399=>"101101110",
  16400=>"110100100",
  16401=>"000001011",
  16402=>"101011000",
  16403=>"001010001",
  16404=>"100000000",
  16405=>"011001111",
  16406=>"100001000",
  16407=>"001100101",
  16408=>"011001001",
  16409=>"110011000",
  16410=>"111011011",
  16411=>"110111111",
  16412=>"011111100",
  16413=>"011010010",
  16414=>"100111100",
  16415=>"010011011",
  16416=>"001110001",
  16417=>"111110111",
  16418=>"010100111",
  16419=>"101001011",
  16420=>"101110110",
  16421=>"000110100",
  16422=>"101101010",
  16423=>"010010000",
  16424=>"011100010",
  16425=>"000010000",
  16426=>"010100101",
  16427=>"100101101",
  16428=>"101110101",
  16429=>"110111001",
  16430=>"011010010",
  16431=>"001000111",
  16432=>"001000011",
  16433=>"110101110",
  16434=>"000000110",
  16435=>"010011001",
  16436=>"100000011",
  16437=>"011100001",
  16438=>"101001111",
  16439=>"010011000",
  16440=>"110000001",
  16441=>"011011100",
  16442=>"111100000",
  16443=>"010000110",
  16444=>"010111000",
  16445=>"101100110",
  16446=>"101000000",
  16447=>"011110110",
  16448=>"111101001",
  16449=>"111011011",
  16450=>"010011011",
  16451=>"011101010",
  16452=>"110101100",
  16453=>"000001110",
  16454=>"010001110",
  16455=>"101101010",
  16456=>"111011000",
  16457=>"000000111",
  16458=>"110001011",
  16459=>"111100011",
  16460=>"000011100",
  16461=>"001111100",
  16462=>"001100011",
  16463=>"010011000",
  16464=>"001111111",
  16465=>"011111011",
  16466=>"001100010",
  16467=>"101011100",
  16468=>"101011001",
  16469=>"000000101",
  16470=>"001000001",
  16471=>"100011101",
  16472=>"101010011",
  16473=>"101110001",
  16474=>"001000101",
  16475=>"100000000",
  16476=>"111000001",
  16477=>"111111110",
  16478=>"110100111",
  16479=>"100100001",
  16480=>"001100111",
  16481=>"010101101",
  16482=>"001110000",
  16483=>"111100000",
  16484=>"110001011",
  16485=>"001001111",
  16486=>"010001101",
  16487=>"101000001",
  16488=>"111111010",
  16489=>"011010010",
  16490=>"110111111",
  16491=>"001010110",
  16492=>"011101000",
  16493=>"000001000",
  16494=>"110111010",
  16495=>"111101111",
  16496=>"001001111",
  16497=>"011011101",
  16498=>"010100001",
  16499=>"010111100",
  16500=>"011101011",
  16501=>"111111010",
  16502=>"100100001",
  16503=>"011111111",
  16504=>"010111111",
  16505=>"110100000",
  16506=>"110110100",
  16507=>"011101010",
  16508=>"110000101",
  16509=>"001100010",
  16510=>"111110000",
  16511=>"100001100",
  16512=>"111011110",
  16513=>"111101000",
  16514=>"000111111",
  16515=>"101000100",
  16516=>"100111100",
  16517=>"000111100",
  16518=>"100100101",
  16519=>"101111110",
  16520=>"111111100",
  16521=>"101110100",
  16522=>"011110001",
  16523=>"011101001",
  16524=>"100010011",
  16525=>"110010110",
  16526=>"100101001",
  16527=>"100000011",
  16528=>"011000001",
  16529=>"001101000",
  16530=>"110100111",
  16531=>"110101000",
  16532=>"110100011",
  16533=>"010011100",
  16534=>"111011011",
  16535=>"000101111",
  16536=>"010000001",
  16537=>"011001011",
  16538=>"100111101",
  16539=>"001001011",
  16540=>"001001110",
  16541=>"001011110",
  16542=>"011001100",
  16543=>"001100100",
  16544=>"000010010",
  16545=>"000010111",
  16546=>"111111111",
  16547=>"111001100",
  16548=>"110110011",
  16549=>"010001101",
  16550=>"000100100",
  16551=>"111010011",
  16552=>"001111011",
  16553=>"010000000",
  16554=>"000110010",
  16555=>"110001100",
  16556=>"000010011",
  16557=>"111011101",
  16558=>"000010011",
  16559=>"011111011",
  16560=>"000101100",
  16561=>"000110101",
  16562=>"111010101",
  16563=>"001010010",
  16564=>"100010111",
  16565=>"000110110",
  16566=>"111101101",
  16567=>"110101010",
  16568=>"010010010",
  16569=>"100111110",
  16570=>"111110011",
  16571=>"100010111",
  16572=>"101011011",
  16573=>"000010011",
  16574=>"010011101",
  16575=>"101101111",
  16576=>"000111101",
  16577=>"100110110",
  16578=>"110011011",
  16579=>"010100001",
  16580=>"001100011",
  16581=>"001000111",
  16582=>"110010001",
  16583=>"001011011",
  16584=>"111010110",
  16585=>"001011110",
  16586=>"001100110",
  16587=>"011000100",
  16588=>"101011101",
  16589=>"111100111",
  16590=>"011101110",
  16591=>"000001001",
  16592=>"001111011",
  16593=>"111110010",
  16594=>"000000101",
  16595=>"100011011",
  16596=>"110101111",
  16597=>"100001100",
  16598=>"000011110",
  16599=>"011011101",
  16600=>"111010100",
  16601=>"111110011",
  16602=>"111011110",
  16603=>"001011100",
  16604=>"110011001",
  16605=>"001100100",
  16606=>"011100001",
  16607=>"100101111",
  16608=>"111100100",
  16609=>"110111100",
  16610=>"100001010",
  16611=>"111111101",
  16612=>"111101100",
  16613=>"011100010",
  16614=>"001011010",
  16615=>"000110100",
  16616=>"001110111",
  16617=>"111111110",
  16618=>"100100000",
  16619=>"001000000",
  16620=>"111010111",
  16621=>"001101110",
  16622=>"010010101",
  16623=>"000111000",
  16624=>"111010010",
  16625=>"010011101",
  16626=>"001010000",
  16627=>"010100101",
  16628=>"011010010",
  16629=>"001101100",
  16630=>"011101000",
  16631=>"011011100",
  16632=>"010000010",
  16633=>"110000010",
  16634=>"001000110",
  16635=>"100110100",
  16636=>"010110110",
  16637=>"110010110",
  16638=>"011100010",
  16639=>"110110111",
  16640=>"111001010",
  16641=>"000111101",
  16642=>"000011101",
  16643=>"001110001",
  16644=>"000011110",
  16645=>"001111000",
  16646=>"011111111",
  16647=>"100001011",
  16648=>"000111001",
  16649=>"110010111",
  16650=>"001100000",
  16651=>"011111001",
  16652=>"011001011",
  16653=>"100101111",
  16654=>"100101111",
  16655=>"000000001",
  16656=>"110000101",
  16657=>"011001011",
  16658=>"111001101",
  16659=>"000011110",
  16660=>"100111011",
  16661=>"111001111",
  16662=>"100110110",
  16663=>"101101111",
  16664=>"010100110",
  16665=>"011100011",
  16666=>"101111101",
  16667=>"110000011",
  16668=>"110110011",
  16669=>"101111111",
  16670=>"000110010",
  16671=>"100010010",
  16672=>"110000101",
  16673=>"111111011",
  16674=>"001111111",
  16675=>"010111100",
  16676=>"101100111",
  16677=>"001101010",
  16678=>"010111011",
  16679=>"111001101",
  16680=>"100001001",
  16681=>"111100010",
  16682=>"011010001",
  16683=>"111010101",
  16684=>"000001001",
  16685=>"111111100",
  16686=>"011000001",
  16687=>"001110001",
  16688=>"000000101",
  16689=>"101000110",
  16690=>"111111011",
  16691=>"001101000",
  16692=>"000010010",
  16693=>"000111001",
  16694=>"001111010",
  16695=>"010000111",
  16696=>"111010010",
  16697=>"010001010",
  16698=>"000010111",
  16699=>"100110111",
  16700=>"100000110",
  16701=>"010110011",
  16702=>"011101100",
  16703=>"100010101",
  16704=>"110110011",
  16705=>"011000001",
  16706=>"000010110",
  16707=>"000011011",
  16708=>"110010100",
  16709=>"001101010",
  16710=>"010000001",
  16711=>"011111010",
  16712=>"010100110",
  16713=>"010100100",
  16714=>"110111010",
  16715=>"100010010",
  16716=>"100010110",
  16717=>"111100001",
  16718=>"110111011",
  16719=>"011101100",
  16720=>"010101000",
  16721=>"100010111",
  16722=>"101000001",
  16723=>"000001100",
  16724=>"100101000",
  16725=>"100000111",
  16726=>"111011001",
  16727=>"010001101",
  16728=>"110001011",
  16729=>"111100111",
  16730=>"000011010",
  16731=>"011101010",
  16732=>"011111100",
  16733=>"111110101",
  16734=>"111111110",
  16735=>"011001000",
  16736=>"011000110",
  16737=>"100111010",
  16738=>"010010100",
  16739=>"010000000",
  16740=>"010011100",
  16741=>"110011011",
  16742=>"011010000",
  16743=>"010111011",
  16744=>"101001111",
  16745=>"110000011",
  16746=>"011111101",
  16747=>"110010011",
  16748=>"111001100",
  16749=>"001110101",
  16750=>"110010010",
  16751=>"010110101",
  16752=>"011010010",
  16753=>"111000101",
  16754=>"101011110",
  16755=>"001010000",
  16756=>"001101011",
  16757=>"101011000",
  16758=>"111001000",
  16759=>"001100111",
  16760=>"001110001",
  16761=>"001001001",
  16762=>"001111100",
  16763=>"010110111",
  16764=>"110010000",
  16765=>"110111011",
  16766=>"000000100",
  16767=>"011000010",
  16768=>"111110000",
  16769=>"011001010",
  16770=>"000000111",
  16771=>"010000001",
  16772=>"110100000",
  16773=>"001000111",
  16774=>"011110111",
  16775=>"111100000",
  16776=>"111111000",
  16777=>"100001111",
  16778=>"011011011",
  16779=>"110011110",
  16780=>"010001011",
  16781=>"011010100",
  16782=>"000110010",
  16783=>"111101000",
  16784=>"000011011",
  16785=>"110101000",
  16786=>"111100100",
  16787=>"010011011",
  16788=>"011111001",
  16789=>"000110011",
  16790=>"000101000",
  16791=>"001111010",
  16792=>"010101101",
  16793=>"010000010",
  16794=>"001100011",
  16795=>"001010101",
  16796=>"011100100",
  16797=>"110100111",
  16798=>"101001110",
  16799=>"001001001",
  16800=>"010100000",
  16801=>"110110111",
  16802=>"111011111",
  16803=>"000111000",
  16804=>"011101110",
  16805=>"011100010",
  16806=>"100110111",
  16807=>"110000111",
  16808=>"110010101",
  16809=>"111001000",
  16810=>"000010111",
  16811=>"111010110",
  16812=>"111100111",
  16813=>"000110100",
  16814=>"000001000",
  16815=>"000110001",
  16816=>"100010110",
  16817=>"111110110",
  16818=>"110000010",
  16819=>"101111101",
  16820=>"011111110",
  16821=>"110100111",
  16822=>"000111111",
  16823=>"001000100",
  16824=>"001001101",
  16825=>"111101011",
  16826=>"110110111",
  16827=>"001000001",
  16828=>"111111001",
  16829=>"011110100",
  16830=>"111010000",
  16831=>"111110101",
  16832=>"011011111",
  16833=>"110001011",
  16834=>"011111011",
  16835=>"011001001",
  16836=>"100001111",
  16837=>"111111001",
  16838=>"110111111",
  16839=>"000110011",
  16840=>"100110000",
  16841=>"101000101",
  16842=>"111011011",
  16843=>"111000010",
  16844=>"101001100",
  16845=>"101110001",
  16846=>"000100110",
  16847=>"100001101",
  16848=>"010010100",
  16849=>"110111010",
  16850=>"011110010",
  16851=>"101010110",
  16852=>"100000010",
  16853=>"000011010",
  16854=>"000100000",
  16855=>"110110000",
  16856=>"100100010",
  16857=>"110111101",
  16858=>"100100110",
  16859=>"000111011",
  16860=>"111111000",
  16861=>"000111011",
  16862=>"011110111",
  16863=>"010010110",
  16864=>"110110010",
  16865=>"110101111",
  16866=>"110110011",
  16867=>"011000100",
  16868=>"001101100",
  16869=>"011100011",
  16870=>"111001010",
  16871=>"011110010",
  16872=>"000010010",
  16873=>"010011000",
  16874=>"000011001",
  16875=>"000110100",
  16876=>"101001011",
  16877=>"011101101",
  16878=>"010110001",
  16879=>"101110101",
  16880=>"101011101",
  16881=>"110001110",
  16882=>"111101100",
  16883=>"111001011",
  16884=>"101000011",
  16885=>"101000111",
  16886=>"010100011",
  16887=>"000110101",
  16888=>"000101100",
  16889=>"100101110",
  16890=>"001100001",
  16891=>"101000100",
  16892=>"001011011",
  16893=>"111110111",
  16894=>"100100001",
  16895=>"111000100",
  16896=>"000011001",
  16897=>"001000100",
  16898=>"110100100",
  16899=>"001110111",
  16900=>"101110111",
  16901=>"111100110",
  16902=>"011000111",
  16903=>"111011000",
  16904=>"110001111",
  16905=>"111010000",
  16906=>"000110101",
  16907=>"010101100",
  16908=>"011010000",
  16909=>"101011111",
  16910=>"101000010",
  16911=>"011000011",
  16912=>"100011010",
  16913=>"100001011",
  16914=>"101011100",
  16915=>"110100010",
  16916=>"110011001",
  16917=>"111100111",
  16918=>"000000001",
  16919=>"101110110",
  16920=>"010010000",
  16921=>"000000010",
  16922=>"100111010",
  16923=>"111101011",
  16924=>"100000001",
  16925=>"010000110",
  16926=>"000010011",
  16927=>"011111111",
  16928=>"001110111",
  16929=>"100101111",
  16930=>"011011111",
  16931=>"010010011",
  16932=>"111101010",
  16933=>"100000000",
  16934=>"000101101",
  16935=>"010111011",
  16936=>"001001101",
  16937=>"011111110",
  16938=>"000111111",
  16939=>"010000100",
  16940=>"101011010",
  16941=>"001000000",
  16942=>"111111101",
  16943=>"011111000",
  16944=>"101010111",
  16945=>"100001011",
  16946=>"111011001",
  16947=>"010011010",
  16948=>"011110010",
  16949=>"111110110",
  16950=>"101101111",
  16951=>"000010011",
  16952=>"011101000",
  16953=>"100100110",
  16954=>"001110101",
  16955=>"100111001",
  16956=>"111011011",
  16957=>"111111111",
  16958=>"101001000",
  16959=>"100101101",
  16960=>"000101011",
  16961=>"100011111",
  16962=>"111001111",
  16963=>"101000100",
  16964=>"000000001",
  16965=>"011000100",
  16966=>"000000010",
  16967=>"110001001",
  16968=>"110101000",
  16969=>"101001010",
  16970=>"110111011",
  16971=>"101000110",
  16972=>"101100000",
  16973=>"011000001",
  16974=>"011101110",
  16975=>"110100000",
  16976=>"100011100",
  16977=>"010011111",
  16978=>"000100101",
  16979=>"011010011",
  16980=>"100101010",
  16981=>"111010110",
  16982=>"111101100",
  16983=>"101011100",
  16984=>"111110100",
  16985=>"011110110",
  16986=>"001101010",
  16987=>"010100001",
  16988=>"101111000",
  16989=>"100011111",
  16990=>"000100011",
  16991=>"010100010",
  16992=>"000110111",
  16993=>"000110001",
  16994=>"110010111",
  16995=>"100010100",
  16996=>"110001101",
  16997=>"110011101",
  16998=>"111000111",
  16999=>"001011101",
  17000=>"000111100",
  17001=>"011010101",
  17002=>"101110001",
  17003=>"010000010",
  17004=>"000101001",
  17005=>"101100111",
  17006=>"001001101",
  17007=>"101110001",
  17008=>"100100000",
  17009=>"110010110",
  17010=>"000001000",
  17011=>"000001110",
  17012=>"001111011",
  17013=>"011100001",
  17014=>"111010101",
  17015=>"111001101",
  17016=>"100110000",
  17017=>"001000100",
  17018=>"000110010",
  17019=>"100011100",
  17020=>"111101101",
  17021=>"100100001",
  17022=>"010001101",
  17023=>"010010100",
  17024=>"001001010",
  17025=>"000000010",
  17026=>"000010000",
  17027=>"101011011",
  17028=>"111111010",
  17029=>"001010110",
  17030=>"011011010",
  17031=>"111111111",
  17032=>"010011000",
  17033=>"000100001",
  17034=>"001001110",
  17035=>"000011101",
  17036=>"000000111",
  17037=>"000100111",
  17038=>"001111101",
  17039=>"011000010",
  17040=>"110010000",
  17041=>"110111000",
  17042=>"010101101",
  17043=>"001010100",
  17044=>"011111100",
  17045=>"001000101",
  17046=>"011011000",
  17047=>"101100011",
  17048=>"101000100",
  17049=>"011000010",
  17050=>"101111110",
  17051=>"111110110",
  17052=>"110001100",
  17053=>"101111111",
  17054=>"010011011",
  17055=>"101000101",
  17056=>"100110001",
  17057=>"010100110",
  17058=>"111111101",
  17059=>"110001110",
  17060=>"001110001",
  17061=>"001110001",
  17062=>"001001011",
  17063=>"111010001",
  17064=>"110100100",
  17065=>"011011100",
  17066=>"111000000",
  17067=>"110110100",
  17068=>"001011000",
  17069=>"111101100",
  17070=>"010000111",
  17071=>"100000110",
  17072=>"011110000",
  17073=>"001011101",
  17074=>"111111100",
  17075=>"010000111",
  17076=>"000001001",
  17077=>"110101111",
  17078=>"011110111",
  17079=>"011111001",
  17080=>"100001000",
  17081=>"110001100",
  17082=>"010101000",
  17083=>"100101110",
  17084=>"110100110",
  17085=>"010110110",
  17086=>"010010101",
  17087=>"101111001",
  17088=>"010000101",
  17089=>"001110000",
  17090=>"111101011",
  17091=>"010000101",
  17092=>"001101001",
  17093=>"101011111",
  17094=>"111000101",
  17095=>"000000000",
  17096=>"110111111",
  17097=>"111110010",
  17098=>"111110101",
  17099=>"001101110",
  17100=>"100101110",
  17101=>"000100111",
  17102=>"011101110",
  17103=>"010000001",
  17104=>"001101100",
  17105=>"000101111",
  17106=>"111110101",
  17107=>"011111000",
  17108=>"010001011",
  17109=>"001110000",
  17110=>"100001001",
  17111=>"000001011",
  17112=>"001000001",
  17113=>"111101110",
  17114=>"111111100",
  17115=>"110001011",
  17116=>"001010101",
  17117=>"110100000",
  17118=>"001100110",
  17119=>"010110111",
  17120=>"000101011",
  17121=>"000000011",
  17122=>"001010010",
  17123=>"100101101",
  17124=>"001001111",
  17125=>"111110001",
  17126=>"100011100",
  17127=>"000010001",
  17128=>"111100000",
  17129=>"111011001",
  17130=>"010000100",
  17131=>"000101001",
  17132=>"000001001",
  17133=>"011111100",
  17134=>"010011011",
  17135=>"011000010",
  17136=>"100001010",
  17137=>"011011110",
  17138=>"010111010",
  17139=>"101111010",
  17140=>"101000010",
  17141=>"100001101",
  17142=>"011111011",
  17143=>"110110111",
  17144=>"100110011",
  17145=>"111100001",
  17146=>"110011000",
  17147=>"100011011",
  17148=>"101000001",
  17149=>"111000110",
  17150=>"101111011",
  17151=>"101011001",
  17152=>"110001000",
  17153=>"101111011",
  17154=>"111110000",
  17155=>"000011101",
  17156=>"100010110",
  17157=>"111111000",
  17158=>"010001101",
  17159=>"101111111",
  17160=>"010010101",
  17161=>"010101010",
  17162=>"111101010",
  17163=>"010110001",
  17164=>"100011101",
  17165=>"001101010",
  17166=>"101000000",
  17167=>"011001010",
  17168=>"011010101",
  17169=>"111011000",
  17170=>"110101100",
  17171=>"001110111",
  17172=>"000110100",
  17173=>"110101001",
  17174=>"110011110",
  17175=>"111000001",
  17176=>"110111101",
  17177=>"011010010",
  17178=>"000101011",
  17179=>"110001110",
  17180=>"101010000",
  17181=>"111000011",
  17182=>"000100110",
  17183=>"110101111",
  17184=>"111110011",
  17185=>"110011001",
  17186=>"110001000",
  17187=>"101011100",
  17188=>"000000000",
  17189=>"010100101",
  17190=>"111111110",
  17191=>"000111010",
  17192=>"100001011",
  17193=>"110111000",
  17194=>"100010101",
  17195=>"101100101",
  17196=>"001010000",
  17197=>"000001010",
  17198=>"110101001",
  17199=>"010000000",
  17200=>"101100011",
  17201=>"000010111",
  17202=>"110100110",
  17203=>"010111000",
  17204=>"110000000",
  17205=>"101010110",
  17206=>"111001110",
  17207=>"001011001",
  17208=>"111110111",
  17209=>"110110110",
  17210=>"110010000",
  17211=>"111100101",
  17212=>"110101001",
  17213=>"101101010",
  17214=>"101110011",
  17215=>"111000111",
  17216=>"101010111",
  17217=>"110001111",
  17218=>"000111000",
  17219=>"111000001",
  17220=>"000011000",
  17221=>"011101011",
  17222=>"000000000",
  17223=>"001111001",
  17224=>"001010101",
  17225=>"011110110",
  17226=>"011110010",
  17227=>"010111000",
  17228=>"011100000",
  17229=>"001101111",
  17230=>"111110110",
  17231=>"100100111",
  17232=>"101111101",
  17233=>"110000100",
  17234=>"001011101",
  17235=>"101001010",
  17236=>"010010101",
  17237=>"101000111",
  17238=>"110110000",
  17239=>"110010001",
  17240=>"011011010",
  17241=>"000000111",
  17242=>"100011111",
  17243=>"101111010",
  17244=>"011110101",
  17245=>"110101010",
  17246=>"000100111",
  17247=>"000111111",
  17248=>"000101010",
  17249=>"100001011",
  17250=>"000001011",
  17251=>"010010000",
  17252=>"100000000",
  17253=>"110011100",
  17254=>"101011010",
  17255=>"111111111",
  17256=>"000010000",
  17257=>"001011000",
  17258=>"101011110",
  17259=>"001001011",
  17260=>"100001110",
  17261=>"011010010",
  17262=>"111110111",
  17263=>"101111000",
  17264=>"111000000",
  17265=>"000001000",
  17266=>"101111011",
  17267=>"011010101",
  17268=>"000101100",
  17269=>"111001010",
  17270=>"010001100",
  17271=>"011111100",
  17272=>"100101011",
  17273=>"101001001",
  17274=>"001111000",
  17275=>"011110011",
  17276=>"000010100",
  17277=>"101010001",
  17278=>"100010111",
  17279=>"010101001",
  17280=>"101001110",
  17281=>"111111110",
  17282=>"110001000",
  17283=>"110110110",
  17284=>"101100111",
  17285=>"110001000",
  17286=>"101100011",
  17287=>"001110010",
  17288=>"010000111",
  17289=>"101010100",
  17290=>"100000110",
  17291=>"110001000",
  17292=>"001000111",
  17293=>"000011111",
  17294=>"101100101",
  17295=>"000001001",
  17296=>"010001001",
  17297=>"011010110",
  17298=>"100010000",
  17299=>"010000010",
  17300=>"100100110",
  17301=>"110011101",
  17302=>"110100101",
  17303=>"001011110",
  17304=>"001101100",
  17305=>"000110111",
  17306=>"010100011",
  17307=>"001000010",
  17308=>"111011101",
  17309=>"110001110",
  17310=>"101000011",
  17311=>"001010100",
  17312=>"110110010",
  17313=>"110111100",
  17314=>"000000100",
  17315=>"100101110",
  17316=>"111010000",
  17317=>"010011111",
  17318=>"110011011",
  17319=>"000101001",
  17320=>"110110101",
  17321=>"111111101",
  17322=>"110010010",
  17323=>"011100110",
  17324=>"000000111",
  17325=>"100100100",
  17326=>"010100010",
  17327=>"110000111",
  17328=>"000100000",
  17329=>"101001011",
  17330=>"001110101",
  17331=>"010111010",
  17332=>"001110001",
  17333=>"001111001",
  17334=>"100000100",
  17335=>"001111000",
  17336=>"011011101",
  17337=>"010110011",
  17338=>"111111110",
  17339=>"011101000",
  17340=>"011101111",
  17341=>"001010010",
  17342=>"000010000",
  17343=>"111001001",
  17344=>"101101001",
  17345=>"111101110",
  17346=>"001000101",
  17347=>"011111001",
  17348=>"011100101",
  17349=>"000000000",
  17350=>"111011110",
  17351=>"011010111",
  17352=>"001100000",
  17353=>"101010010",
  17354=>"111110100",
  17355=>"111101100",
  17356=>"000101001",
  17357=>"111010100",
  17358=>"010010111",
  17359=>"100011100",
  17360=>"111010011",
  17361=>"110110010",
  17362=>"111110111",
  17363=>"111101011",
  17364=>"000001111",
  17365=>"100011110",
  17366=>"100111111",
  17367=>"010011111",
  17368=>"000101111",
  17369=>"110000000",
  17370=>"001010001",
  17371=>"111000000",
  17372=>"110001000",
  17373=>"010101000",
  17374=>"111000100",
  17375=>"110001000",
  17376=>"101000011",
  17377=>"110001111",
  17378=>"011110011",
  17379=>"100101101",
  17380=>"110100110",
  17381=>"011101110",
  17382=>"010111010",
  17383=>"100000111",
  17384=>"000001001",
  17385=>"101011010",
  17386=>"111100111",
  17387=>"110100100",
  17388=>"111010011",
  17389=>"100100101",
  17390=>"000110110",
  17391=>"111110110",
  17392=>"101100000",
  17393=>"000001111",
  17394=>"111100101",
  17395=>"111111101",
  17396=>"101010001",
  17397=>"010110110",
  17398=>"111110100",
  17399=>"101001001",
  17400=>"001001000",
  17401=>"001101011",
  17402=>"010010011",
  17403=>"011100011",
  17404=>"000101101",
  17405=>"011110001",
  17406=>"101001001",
  17407=>"011001110",
  17408=>"000000101",
  17409=>"001010101",
  17410=>"000011110",
  17411=>"111100011",
  17412=>"000010000",
  17413=>"010001000",
  17414=>"001110011",
  17415=>"110011000",
  17416=>"100010111",
  17417=>"100000010",
  17418=>"101000001",
  17419=>"110011110",
  17420=>"000100001",
  17421=>"011101000",
  17422=>"101001000",
  17423=>"011110111",
  17424=>"011000101",
  17425=>"000100001",
  17426=>"011011100",
  17427=>"000001010",
  17428=>"110101101",
  17429=>"111111011",
  17430=>"101000011",
  17431=>"000011101",
  17432=>"011111100",
  17433=>"010011110",
  17434=>"000000110",
  17435=>"000010000",
  17436=>"101101100",
  17437=>"100100011",
  17438=>"000111000",
  17439=>"111000000",
  17440=>"011001001",
  17441=>"101011111",
  17442=>"011010001",
  17443=>"111011010",
  17444=>"111100000",
  17445=>"011101111",
  17446=>"100101111",
  17447=>"110101101",
  17448=>"000011110",
  17449=>"111000110",
  17450=>"011011110",
  17451=>"010111100",
  17452=>"110001010",
  17453=>"010001001",
  17454=>"000001001",
  17455=>"100100110",
  17456=>"011111100",
  17457=>"011111010",
  17458=>"000111000",
  17459=>"000000010",
  17460=>"000011100",
  17461=>"110110010",
  17462=>"100010100",
  17463=>"111101010",
  17464=>"001100110",
  17465=>"101010100",
  17466=>"010000000",
  17467=>"101100111",
  17468=>"110100000",
  17469=>"100010110",
  17470=>"111111100",
  17471=>"010101100",
  17472=>"010001010",
  17473=>"000000101",
  17474=>"111110001",
  17475=>"101110101",
  17476=>"001101110",
  17477=>"110010000",
  17478=>"101000011",
  17479=>"001010100",
  17480=>"110011110",
  17481=>"100011101",
  17482=>"000111000",
  17483=>"101100101",
  17484=>"011111010",
  17485=>"110011001",
  17486=>"100000001",
  17487=>"000110110",
  17488=>"010101001",
  17489=>"000010001",
  17490=>"110110010",
  17491=>"111111110",
  17492=>"000000000",
  17493=>"110110110",
  17494=>"000100100",
  17495=>"000010101",
  17496=>"110011100",
  17497=>"101000000",
  17498=>"100000110",
  17499=>"100000000",
  17500=>"001101000",
  17501=>"101001010",
  17502=>"101010100",
  17503=>"110000000",
  17504=>"001010111",
  17505=>"100100100",
  17506=>"100100011",
  17507=>"111100000",
  17508=>"101110110",
  17509=>"101111010",
  17510=>"001001011",
  17511=>"100111100",
  17512=>"111010100",
  17513=>"101111101",
  17514=>"001011000",
  17515=>"111011000",
  17516=>"011001101",
  17517=>"111010101",
  17518=>"010100001",
  17519=>"110110000",
  17520=>"100111101",
  17521=>"110101010",
  17522=>"101010000",
  17523=>"000101110",
  17524=>"100100000",
  17525=>"100110010",
  17526=>"111101111",
  17527=>"001001100",
  17528=>"110100101",
  17529=>"011000101",
  17530=>"000001000",
  17531=>"001111010",
  17532=>"001010101",
  17533=>"001100000",
  17534=>"010100000",
  17535=>"001010110",
  17536=>"011000101",
  17537=>"000010111",
  17538=>"011010001",
  17539=>"101011110",
  17540=>"010011111",
  17541=>"110111001",
  17542=>"110011011",
  17543=>"010001111",
  17544=>"101001011",
  17545=>"000001011",
  17546=>"010100011",
  17547=>"010111110",
  17548=>"000001011",
  17549=>"000110111",
  17550=>"110011111",
  17551=>"001111000",
  17552=>"100011110",
  17553=>"111010011",
  17554=>"110001101",
  17555=>"100111000",
  17556=>"000000000",
  17557=>"101100011",
  17558=>"001101000",
  17559=>"101000010",
  17560=>"000111110",
  17561=>"101010111",
  17562=>"111000100",
  17563=>"110110111",
  17564=>"011010001",
  17565=>"010010100",
  17566=>"100010010",
  17567=>"000100010",
  17568=>"010000101",
  17569=>"001101101",
  17570=>"111011101",
  17571=>"000010101",
  17572=>"100001001",
  17573=>"111011001",
  17574=>"110000100",
  17575=>"001000111",
  17576=>"001011110",
  17577=>"011000011",
  17578=>"110000001",
  17579=>"000010100",
  17580=>"101001101",
  17581=>"000000100",
  17582=>"110111110",
  17583=>"011010010",
  17584=>"001010100",
  17585=>"111111101",
  17586=>"001111110",
  17587=>"110011111",
  17588=>"011001100",
  17589=>"110101000",
  17590=>"110000011",
  17591=>"001100111",
  17592=>"011000001",
  17593=>"111010110",
  17594=>"100101100",
  17595=>"110111011",
  17596=>"111111010",
  17597=>"110000110",
  17598=>"011100010",
  17599=>"001110101",
  17600=>"010011001",
  17601=>"111100101",
  17602=>"000111000",
  17603=>"000110010",
  17604=>"100000000",
  17605=>"110011000",
  17606=>"000001100",
  17607=>"100100101",
  17608=>"110100001",
  17609=>"001101110",
  17610=>"100001111",
  17611=>"010010001",
  17612=>"110010110",
  17613=>"011011111",
  17614=>"111101000",
  17615=>"000000000",
  17616=>"001111001",
  17617=>"111111100",
  17618=>"000011100",
  17619=>"101110001",
  17620=>"111001101",
  17621=>"111100000",
  17622=>"000001011",
  17623=>"111100111",
  17624=>"010101111",
  17625=>"110111000",
  17626=>"011101110",
  17627=>"000110010",
  17628=>"111101000",
  17629=>"011010111",
  17630=>"101100001",
  17631=>"101100111",
  17632=>"001000000",
  17633=>"000011001",
  17634=>"001010100",
  17635=>"010001011",
  17636=>"010000111",
  17637=>"011001000",
  17638=>"101101110",
  17639=>"010000000",
  17640=>"101011111",
  17641=>"100010101",
  17642=>"100101011",
  17643=>"010000000",
  17644=>"100000001",
  17645=>"000010101",
  17646=>"110110101",
  17647=>"110110100",
  17648=>"001000010",
  17649=>"001000110",
  17650=>"101000111",
  17651=>"010000000",
  17652=>"010101101",
  17653=>"110011111",
  17654=>"111111001",
  17655=>"000101011",
  17656=>"100001001",
  17657=>"111111001",
  17658=>"010111000",
  17659=>"110101011",
  17660=>"000111001",
  17661=>"010011011",
  17662=>"010110011",
  17663=>"010011010",
  17664=>"011100000",
  17665=>"110011101",
  17666=>"011111101",
  17667=>"111111101",
  17668=>"010001010",
  17669=>"000010011",
  17670=>"100110111",
  17671=>"101101110",
  17672=>"001011100",
  17673=>"000011000",
  17674=>"100110000",
  17675=>"010011000",
  17676=>"110101000",
  17677=>"011011011",
  17678=>"100000110",
  17679=>"010010100",
  17680=>"010010000",
  17681=>"011101010",
  17682=>"011011000",
  17683=>"000100001",
  17684=>"110110101",
  17685=>"111110111",
  17686=>"111011111",
  17687=>"110001100",
  17688=>"111100001",
  17689=>"111000000",
  17690=>"011101000",
  17691=>"010010001",
  17692=>"110000000",
  17693=>"111110110",
  17694=>"100111011",
  17695=>"100011101",
  17696=>"010101011",
  17697=>"000111111",
  17698=>"101011011",
  17699=>"000101011",
  17700=>"010011100",
  17701=>"010010110",
  17702=>"101101101",
  17703=>"100011110",
  17704=>"100000011",
  17705=>"110111001",
  17706=>"011111010",
  17707=>"101100001",
  17708=>"110111100",
  17709=>"000010000",
  17710=>"000110010",
  17711=>"110001100",
  17712=>"101111010",
  17713=>"110101001",
  17714=>"110000010",
  17715=>"001011000",
  17716=>"111100101",
  17717=>"000010101",
  17718=>"100000111",
  17719=>"101010101",
  17720=>"110000011",
  17721=>"111010111",
  17722=>"010010001",
  17723=>"011011000",
  17724=>"001110011",
  17725=>"011101111",
  17726=>"011001010",
  17727=>"000001110",
  17728=>"011101110",
  17729=>"011000101",
  17730=>"110011000",
  17731=>"001001001",
  17732=>"101011111",
  17733=>"110000100",
  17734=>"110111000",
  17735=>"001001000",
  17736=>"101110011",
  17737=>"011001110",
  17738=>"111111110",
  17739=>"010001000",
  17740=>"000000011",
  17741=>"111010111",
  17742=>"101101010",
  17743=>"111010111",
  17744=>"011110001",
  17745=>"010011000",
  17746=>"111001010",
  17747=>"010111011",
  17748=>"011001011",
  17749=>"111110101",
  17750=>"001100100",
  17751=>"100011011",
  17752=>"000101101",
  17753=>"010001100",
  17754=>"010110100",
  17755=>"101000010",
  17756=>"101100001",
  17757=>"101111000",
  17758=>"110110111",
  17759=>"111010000",
  17760=>"001000101",
  17761=>"001111110",
  17762=>"010011001",
  17763=>"001100100",
  17764=>"101010001",
  17765=>"111100011",
  17766=>"000111100",
  17767=>"111110000",
  17768=>"011000000",
  17769=>"001100001",
  17770=>"010111001",
  17771=>"101111010",
  17772=>"101000001",
  17773=>"111001100",
  17774=>"010001010",
  17775=>"001010010",
  17776=>"001011101",
  17777=>"110001110",
  17778=>"011111101",
  17779=>"101011011",
  17780=>"111100101",
  17781=>"110100110",
  17782=>"100010100",
  17783=>"111001111",
  17784=>"000000111",
  17785=>"100000000",
  17786=>"101110101",
  17787=>"010101101",
  17788=>"001100101",
  17789=>"111000100",
  17790=>"111001110",
  17791=>"011011100",
  17792=>"110011110",
  17793=>"000001011",
  17794=>"001010010",
  17795=>"001000100",
  17796=>"100010011",
  17797=>"001101011",
  17798=>"110011100",
  17799=>"101111111",
  17800=>"001011110",
  17801=>"101011101",
  17802=>"100110010",
  17803=>"001010000",
  17804=>"011011101",
  17805=>"100000000",
  17806=>"111100011",
  17807=>"010010000",
  17808=>"001010000",
  17809=>"001000000",
  17810=>"000000110",
  17811=>"000010111",
  17812=>"110001001",
  17813=>"100011111",
  17814=>"110001001",
  17815=>"000010001",
  17816=>"101110101",
  17817=>"110010110",
  17818=>"000011010",
  17819=>"000001010",
  17820=>"010110001",
  17821=>"111111111",
  17822=>"100010101",
  17823=>"000001101",
  17824=>"001100010",
  17825=>"111111101",
  17826=>"011110001",
  17827=>"111101101",
  17828=>"001111011",
  17829=>"101010010",
  17830=>"010000010",
  17831=>"100001111",
  17832=>"110010100",
  17833=>"011101011",
  17834=>"011110001",
  17835=>"100110111",
  17836=>"110001110",
  17837=>"110000011",
  17838=>"110110101",
  17839=>"111110100",
  17840=>"110010000",
  17841=>"110100111",
  17842=>"111100011",
  17843=>"011111000",
  17844=>"111101110",
  17845=>"001110100",
  17846=>"101110101",
  17847=>"110001011",
  17848=>"111010110",
  17849=>"000101101",
  17850=>"000010000",
  17851=>"110101111",
  17852=>"000110001",
  17853=>"001101011",
  17854=>"011100000",
  17855=>"001010101",
  17856=>"101001000",
  17857=>"100010001",
  17858=>"111111111",
  17859=>"011110000",
  17860=>"000000111",
  17861=>"110101101",
  17862=>"000000111",
  17863=>"011111001",
  17864=>"000000010",
  17865=>"001111111",
  17866=>"111010010",
  17867=>"011101000",
  17868=>"001110101",
  17869=>"011010000",
  17870=>"110111010",
  17871=>"011010001",
  17872=>"001111011",
  17873=>"000111101",
  17874=>"010110001",
  17875=>"000000101",
  17876=>"111011001",
  17877=>"001011110",
  17878=>"101111111",
  17879=>"011000000",
  17880=>"001111101",
  17881=>"010110010",
  17882=>"111110101",
  17883=>"101000000",
  17884=>"000100000",
  17885=>"111110101",
  17886=>"010110110",
  17887=>"010010101",
  17888=>"010001110",
  17889=>"110111000",
  17890=>"110100000",
  17891=>"101101101",
  17892=>"001000001",
  17893=>"111101111",
  17894=>"010001010",
  17895=>"000001110",
  17896=>"010111111",
  17897=>"111001111",
  17898=>"011000111",
  17899=>"111010001",
  17900=>"101001110",
  17901=>"001000111",
  17902=>"010110111",
  17903=>"100100111",
  17904=>"100100101",
  17905=>"010110010",
  17906=>"101000111",
  17907=>"000100100",
  17908=>"011110011",
  17909=>"000011001",
  17910=>"010010010",
  17911=>"100110010",
  17912=>"001000110",
  17913=>"110010010",
  17914=>"001101000",
  17915=>"111101111",
  17916=>"000111101",
  17917=>"001010000",
  17918=>"101110110",
  17919=>"100110110",
  17920=>"101100111",
  17921=>"010100010",
  17922=>"100100010",
  17923=>"111100101",
  17924=>"110100100",
  17925=>"000010010",
  17926=>"111100100",
  17927=>"111001101",
  17928=>"011100100",
  17929=>"010101000",
  17930=>"110111000",
  17931=>"100000010",
  17932=>"111110101",
  17933=>"110100011",
  17934=>"110000010",
  17935=>"000111010",
  17936=>"110111101",
  17937=>"111111111",
  17938=>"101011101",
  17939=>"110001010",
  17940=>"101100001",
  17941=>"111110001",
  17942=>"110000111",
  17943=>"111010011",
  17944=>"011011111",
  17945=>"011011000",
  17946=>"101000010",
  17947=>"000010111",
  17948=>"110110010",
  17949=>"110100101",
  17950=>"100001111",
  17951=>"111001110",
  17952=>"101110011",
  17953=>"101100001",
  17954=>"111000111",
  17955=>"110011011",
  17956=>"110011011",
  17957=>"010110111",
  17958=>"001000000",
  17959=>"000000110",
  17960=>"110101100",
  17961=>"010101101",
  17962=>"001010101",
  17963=>"000000111",
  17964=>"011111111",
  17965=>"001100000",
  17966=>"101101010",
  17967=>"111011101",
  17968=>"010111101",
  17969=>"010010111",
  17970=>"110101100",
  17971=>"100100000",
  17972=>"001000011",
  17973=>"100101100",
  17974=>"001111011",
  17975=>"100100111",
  17976=>"111010011",
  17977=>"010000110",
  17978=>"100010101",
  17979=>"101001001",
  17980=>"110010100",
  17981=>"000010100",
  17982=>"000101100",
  17983=>"010010000",
  17984=>"010011101",
  17985=>"000010000",
  17986=>"101000111",
  17987=>"011011110",
  17988=>"101001000",
  17989=>"011111000",
  17990=>"001000000",
  17991=>"100110000",
  17992=>"001110000",
  17993=>"100100111",
  17994=>"010111111",
  17995=>"110001110",
  17996=>"010011000",
  17997=>"111101110",
  17998=>"011111110",
  17999=>"111111100",
  18000=>"011111001",
  18001=>"001100111",
  18002=>"110100101",
  18003=>"110101010",
  18004=>"100110001",
  18005=>"000010011",
  18006=>"010000101",
  18007=>"000001101",
  18008=>"110010100",
  18009=>"000011111",
  18010=>"101100111",
  18011=>"101000110",
  18012=>"000101111",
  18013=>"000000000",
  18014=>"000001000",
  18015=>"111000100",
  18016=>"110001101",
  18017=>"110000011",
  18018=>"100011100",
  18019=>"010100010",
  18020=>"101100101",
  18021=>"011011011",
  18022=>"011011010",
  18023=>"101100010",
  18024=>"111101001",
  18025=>"010110100",
  18026=>"000000010",
  18027=>"000101001",
  18028=>"100011101",
  18029=>"111000011",
  18030=>"000111100",
  18031=>"110111111",
  18032=>"101001010",
  18033=>"010000100",
  18034=>"000110001",
  18035=>"111010111",
  18036=>"110000001",
  18037=>"101111010",
  18038=>"001101000",
  18039=>"110110110",
  18040=>"011011100",
  18041=>"110010011",
  18042=>"100001010",
  18043=>"001111010",
  18044=>"010111001",
  18045=>"001000100",
  18046=>"111110111",
  18047=>"101000101",
  18048=>"001010010",
  18049=>"010101101",
  18050=>"100111000",
  18051=>"101111001",
  18052=>"001010100",
  18053=>"110010100",
  18054=>"001011010",
  18055=>"001100101",
  18056=>"110000111",
  18057=>"011101111",
  18058=>"110110010",
  18059=>"000100001",
  18060=>"000001000",
  18061=>"011000100",
  18062=>"100001101",
  18063=>"110000111",
  18064=>"110111000",
  18065=>"110010011",
  18066=>"110111010",
  18067=>"010001010",
  18068=>"101101000",
  18069=>"110001100",
  18070=>"000111110",
  18071=>"010100101",
  18072=>"111000111",
  18073=>"001111000",
  18074=>"001011111",
  18075=>"010111001",
  18076=>"000000100",
  18077=>"011111100",
  18078=>"100101111",
  18079=>"001111111",
  18080=>"000010110",
  18081=>"011001011",
  18082=>"101001010",
  18083=>"011110111",
  18084=>"101110111",
  18085=>"010011001",
  18086=>"111000010",
  18087=>"011000101",
  18088=>"111001011",
  18089=>"000100110",
  18090=>"000010110",
  18091=>"011101101",
  18092=>"010011000",
  18093=>"000001000",
  18094=>"111010110",
  18095=>"101111111",
  18096=>"101011000",
  18097=>"001100001",
  18098=>"100001111",
  18099=>"011000011",
  18100=>"010001011",
  18101=>"100110011",
  18102=>"011110101",
  18103=>"000110000",
  18104=>"100100101",
  18105=>"001000101",
  18106=>"000101000",
  18107=>"000111001",
  18108=>"011010111",
  18109=>"110111001",
  18110=>"111010010",
  18111=>"111100100",
  18112=>"001011010",
  18113=>"010011011",
  18114=>"010010110",
  18115=>"011001001",
  18116=>"101110000",
  18117=>"101001101",
  18118=>"101001111",
  18119=>"001010110",
  18120=>"000010010",
  18121=>"000100001",
  18122=>"001101111",
  18123=>"111111101",
  18124=>"011010110",
  18125=>"001000100",
  18126=>"111010010",
  18127=>"111010010",
  18128=>"111110111",
  18129=>"011111010",
  18130=>"110010011",
  18131=>"001101100",
  18132=>"110010111",
  18133=>"010010100",
  18134=>"100110111",
  18135=>"110101101",
  18136=>"000100111",
  18137=>"010111100",
  18138=>"100110000",
  18139=>"101011110",
  18140=>"101011010",
  18141=>"100000101",
  18142=>"111101010",
  18143=>"101001100",
  18144=>"110110111",
  18145=>"101100010",
  18146=>"111010001",
  18147=>"011001010",
  18148=>"111010010",
  18149=>"010010000",
  18150=>"100100011",
  18151=>"010010000",
  18152=>"001101111",
  18153=>"011001110",
  18154=>"111011110",
  18155=>"110001010",
  18156=>"011111101",
  18157=>"010001000",
  18158=>"101101001",
  18159=>"100110100",
  18160=>"001000111",
  18161=>"010110110",
  18162=>"011011111",
  18163=>"010010010",
  18164=>"100000111",
  18165=>"010110001",
  18166=>"110000111",
  18167=>"111101001",
  18168=>"011000010",
  18169=>"110110010",
  18170=>"000000011",
  18171=>"110000100",
  18172=>"111010010",
  18173=>"011010100",
  18174=>"000001001",
  18175=>"000100001",
  18176=>"000101011",
  18177=>"110100100",
  18178=>"101101001",
  18179=>"011000011",
  18180=>"001010011",
  18181=>"111010001",
  18182=>"100110110",
  18183=>"000110000",
  18184=>"010110011",
  18185=>"110111110",
  18186=>"000011000",
  18187=>"111010111",
  18188=>"101111100",
  18189=>"101000011",
  18190=>"110011011",
  18191=>"100100010",
  18192=>"011111110",
  18193=>"011111111",
  18194=>"101100010",
  18195=>"110010101",
  18196=>"100100111",
  18197=>"111111011",
  18198=>"001000100",
  18199=>"100111011",
  18200=>"010010100",
  18201=>"110110100",
  18202=>"101000111",
  18203=>"011101110",
  18204=>"101100011",
  18205=>"001001111",
  18206=>"001001101",
  18207=>"010101001",
  18208=>"111110011",
  18209=>"100100101",
  18210=>"110100011",
  18211=>"010011100",
  18212=>"001101010",
  18213=>"100111111",
  18214=>"111100000",
  18215=>"111110111",
  18216=>"010100011",
  18217=>"000000010",
  18218=>"100010111",
  18219=>"001110011",
  18220=>"010101000",
  18221=>"011010101",
  18222=>"110100010",
  18223=>"101000101",
  18224=>"001011001",
  18225=>"011011101",
  18226=>"011011010",
  18227=>"000010001",
  18228=>"000100101",
  18229=>"000000001",
  18230=>"111011111",
  18231=>"011111111",
  18232=>"000110101",
  18233=>"101101000",
  18234=>"011101101",
  18235=>"000100011",
  18236=>"100000111",
  18237=>"010100100",
  18238=>"110100100",
  18239=>"100111011",
  18240=>"111001101",
  18241=>"111111101",
  18242=>"001001100",
  18243=>"001010111",
  18244=>"010100110",
  18245=>"010000110",
  18246=>"100110110",
  18247=>"000110000",
  18248=>"100001000",
  18249=>"100011110",
  18250=>"000001000",
  18251=>"000001000",
  18252=>"010001000",
  18253=>"100001000",
  18254=>"100011110",
  18255=>"001000101",
  18256=>"010100000",
  18257=>"111111111",
  18258=>"100100001",
  18259=>"010001000",
  18260=>"110101001",
  18261=>"000011111",
  18262=>"000000001",
  18263=>"000001010",
  18264=>"000001011",
  18265=>"110001110",
  18266=>"010001100",
  18267=>"110111110",
  18268=>"101001100",
  18269=>"101110001",
  18270=>"011000100",
  18271=>"100011000",
  18272=>"100111110",
  18273=>"010110001",
  18274=>"001011111",
  18275=>"100110011",
  18276=>"111000110",
  18277=>"111100100",
  18278=>"110010000",
  18279=>"011001111",
  18280=>"011011111",
  18281=>"111011110",
  18282=>"101110110",
  18283=>"111011111",
  18284=>"100001010",
  18285=>"000100001",
  18286=>"011010011",
  18287=>"011110100",
  18288=>"100000000",
  18289=>"100000011",
  18290=>"001011100",
  18291=>"111011011",
  18292=>"000110011",
  18293=>"000001001",
  18294=>"100011100",
  18295=>"001011011",
  18296=>"111001111",
  18297=>"010010000",
  18298=>"010001001",
  18299=>"001110011",
  18300=>"011001000",
  18301=>"110110001",
  18302=>"111011011",
  18303=>"111110111",
  18304=>"011000000",
  18305=>"000101111",
  18306=>"011000101",
  18307=>"010101010",
  18308=>"110000101",
  18309=>"010000001",
  18310=>"001111111",
  18311=>"111111011",
  18312=>"001111001",
  18313=>"001110100",
  18314=>"111110010",
  18315=>"001010010",
  18316=>"110011010",
  18317=>"111100111",
  18318=>"010001010",
  18319=>"010001001",
  18320=>"001000000",
  18321=>"101101101",
  18322=>"011110100",
  18323=>"100000110",
  18324=>"011001011",
  18325=>"110110011",
  18326=>"000011111",
  18327=>"001011000",
  18328=>"100111101",
  18329=>"111101011",
  18330=>"101000001",
  18331=>"001100111",
  18332=>"001000001",
  18333=>"000001010",
  18334=>"000000111",
  18335=>"111101011",
  18336=>"000001111",
  18337=>"010100001",
  18338=>"001111000",
  18339=>"011100000",
  18340=>"101111111",
  18341=>"110110010",
  18342=>"111111111",
  18343=>"100011001",
  18344=>"100011000",
  18345=>"000000101",
  18346=>"101111111",
  18347=>"011110111",
  18348=>"100001100",
  18349=>"101111100",
  18350=>"111110010",
  18351=>"011010100",
  18352=>"010010000",
  18353=>"100110110",
  18354=>"111101110",
  18355=>"001010100",
  18356=>"011101010",
  18357=>"010011010",
  18358=>"100011100",
  18359=>"001010101",
  18360=>"001100101",
  18361=>"000100010",
  18362=>"110000111",
  18363=>"011110000",
  18364=>"101010011",
  18365=>"011010101",
  18366=>"000101100",
  18367=>"010000010",
  18368=>"101100011",
  18369=>"000001101",
  18370=>"100001010",
  18371=>"100110110",
  18372=>"100100111",
  18373=>"010000011",
  18374=>"110111100",
  18375=>"010110001",
  18376=>"110000100",
  18377=>"100010111",
  18378=>"110011011",
  18379=>"011111001",
  18380=>"100011001",
  18381=>"000100011",
  18382=>"110000101",
  18383=>"111001100",
  18384=>"001111110",
  18385=>"001010001",
  18386=>"010110010",
  18387=>"000101000",
  18388=>"000011010",
  18389=>"111010111",
  18390=>"000011010",
  18391=>"000001010",
  18392=>"000101000",
  18393=>"110101001",
  18394=>"111000011",
  18395=>"010101110",
  18396=>"000010110",
  18397=>"111111010",
  18398=>"011101011",
  18399=>"101001001",
  18400=>"110111010",
  18401=>"111101101",
  18402=>"010101101",
  18403=>"110001110",
  18404=>"100101010",
  18405=>"100101110",
  18406=>"100010000",
  18407=>"010110101",
  18408=>"000100111",
  18409=>"110101111",
  18410=>"101000000",
  18411=>"000001010",
  18412=>"010111010",
  18413=>"100010011",
  18414=>"000001101",
  18415=>"111111110",
  18416=>"101100111",
  18417=>"111001100",
  18418=>"010010000",
  18419=>"100011011",
  18420=>"011010000",
  18421=>"011011100",
  18422=>"101111011",
  18423=>"100001101",
  18424=>"100001011",
  18425=>"100100000",
  18426=>"010110010",
  18427=>"010110000",
  18428=>"000011010",
  18429=>"000010000",
  18430=>"100101000",
  18431=>"110110000",
  18432=>"100100000",
  18433=>"110101000",
  18434=>"000110111",
  18435=>"000111110",
  18436=>"000010000",
  18437=>"010011101",
  18438=>"101111101",
  18439=>"010000101",
  18440=>"110011100",
  18441=>"011110011",
  18442=>"111011001",
  18443=>"110111111",
  18444=>"010110001",
  18445=>"010001100",
  18446=>"111001111",
  18447=>"010011010",
  18448=>"001110011",
  18449=>"010100011",
  18450=>"011100100",
  18451=>"001101000",
  18452=>"000111010",
  18453=>"101001111",
  18454=>"100010100",
  18455=>"111011100",
  18456=>"001111000",
  18457=>"111110111",
  18458=>"011100101",
  18459=>"100111111",
  18460=>"111011010",
  18461=>"001110101",
  18462=>"010001110",
  18463=>"001110100",
  18464=>"001000000",
  18465=>"010001111",
  18466=>"011100000",
  18467=>"000111001",
  18468=>"000111000",
  18469=>"011010001",
  18470=>"001011000",
  18471=>"011101101",
  18472=>"101010111",
  18473=>"001000010",
  18474=>"101001100",
  18475=>"110111111",
  18476=>"111011001",
  18477=>"001110101",
  18478=>"000001010",
  18479=>"001100010",
  18480=>"110100000",
  18481=>"100010110",
  18482=>"100100110",
  18483=>"010011000",
  18484=>"110101000",
  18485=>"110011011",
  18486=>"101001010",
  18487=>"000010111",
  18488=>"010111011",
  18489=>"110100001",
  18490=>"111011100",
  18491=>"011001010",
  18492=>"001111101",
  18493=>"010010111",
  18494=>"101001011",
  18495=>"111011111",
  18496=>"000011110",
  18497=>"111101010",
  18498=>"111111011",
  18499=>"010101011",
  18500=>"111000011",
  18501=>"000000011",
  18502=>"011110010",
  18503=>"010011001",
  18504=>"010110001",
  18505=>"000010111",
  18506=>"001100100",
  18507=>"000001101",
  18508=>"000101101",
  18509=>"101101111",
  18510=>"011000111",
  18511=>"101011100",
  18512=>"001001101",
  18513=>"111100101",
  18514=>"000110101",
  18515=>"100100101",
  18516=>"010000000",
  18517=>"101101101",
  18518=>"010000001",
  18519=>"110111110",
  18520=>"111101000",
  18521=>"000001000",
  18522=>"011001011",
  18523=>"011100011",
  18524=>"101111011",
  18525=>"010001100",
  18526=>"011110100",
  18527=>"110001000",
  18528=>"001111111",
  18529=>"001110011",
  18530=>"100000001",
  18531=>"000001010",
  18532=>"110111000",
  18533=>"011001011",
  18534=>"101101010",
  18535=>"001100100",
  18536=>"000010001",
  18537=>"001001100",
  18538=>"000010000",
  18539=>"010001111",
  18540=>"011001100",
  18541=>"011101111",
  18542=>"011110100",
  18543=>"010011100",
  18544=>"110101110",
  18545=>"000001000",
  18546=>"110010010",
  18547=>"000010010",
  18548=>"111111010",
  18549=>"000110111",
  18550=>"110010101",
  18551=>"111010001",
  18552=>"100100011",
  18553=>"001101111",
  18554=>"011101000",
  18555=>"111101010",
  18556=>"110000011",
  18557=>"110011110",
  18558=>"101010110",
  18559=>"100110100",
  18560=>"000111011",
  18561=>"011010110",
  18562=>"111100011",
  18563=>"010100100",
  18564=>"110001010",
  18565=>"100011010",
  18566=>"000001011",
  18567=>"001010001",
  18568=>"010100010",
  18569=>"010000000",
  18570=>"000101111",
  18571=>"001110110",
  18572=>"011111101",
  18573=>"001101101",
  18574=>"101001001",
  18575=>"110101111",
  18576=>"011111001",
  18577=>"000011100",
  18578=>"100000010",
  18579=>"000011001",
  18580=>"111011101",
  18581=>"110111111",
  18582=>"101011010",
  18583=>"101010000",
  18584=>"000110101",
  18585=>"101010011",
  18586=>"001100001",
  18587=>"111011101",
  18588=>"101011011",
  18589=>"011011001",
  18590=>"000001100",
  18591=>"010110101",
  18592=>"101111000",
  18593=>"011010101",
  18594=>"001101001",
  18595=>"000000011",
  18596=>"110000000",
  18597=>"101011011",
  18598=>"001100000",
  18599=>"111001000",
  18600=>"011011010",
  18601=>"100100111",
  18602=>"100011101",
  18603=>"100101101",
  18604=>"000000000",
  18605=>"000001100",
  18606=>"000101110",
  18607=>"111011110",
  18608=>"000111000",
  18609=>"111010010",
  18610=>"000001100",
  18611=>"100100101",
  18612=>"111011111",
  18613=>"000011011",
  18614=>"110110100",
  18615=>"101111110",
  18616=>"011110100",
  18617=>"110000011",
  18618=>"001000101",
  18619=>"111101111",
  18620=>"101011011",
  18621=>"110101100",
  18622=>"111110110",
  18623=>"110111011",
  18624=>"100100110",
  18625=>"101010100",
  18626=>"111011000",
  18627=>"101000000",
  18628=>"101010000",
  18629=>"111110101",
  18630=>"100010100",
  18631=>"110000100",
  18632=>"000010000",
  18633=>"000000000",
  18634=>"001000101",
  18635=>"101000111",
  18636=>"110001001",
  18637=>"110000110",
  18638=>"000000001",
  18639=>"111011001",
  18640=>"111101110",
  18641=>"011110110",
  18642=>"011101000",
  18643=>"100000010",
  18644=>"110101110",
  18645=>"011101001",
  18646=>"101000101",
  18647=>"111011010",
  18648=>"010011001",
  18649=>"011110100",
  18650=>"010111000",
  18651=>"111110000",
  18652=>"111110001",
  18653=>"101001001",
  18654=>"110111101",
  18655=>"010011100",
  18656=>"111000001",
  18657=>"011001001",
  18658=>"011000000",
  18659=>"110011101",
  18660=>"010110100",
  18661=>"101000010",
  18662=>"111111010",
  18663=>"110011011",
  18664=>"101110011",
  18665=>"101110011",
  18666=>"111010100",
  18667=>"101000011",
  18668=>"001111101",
  18669=>"100111000",
  18670=>"000001010",
  18671=>"000000100",
  18672=>"111010011",
  18673=>"010001101",
  18674=>"011000111",
  18675=>"011101111",
  18676=>"111111001",
  18677=>"110100111",
  18678=>"100101101",
  18679=>"010100101",
  18680=>"001001001",
  18681=>"000110011",
  18682=>"111101100",
  18683=>"110111001",
  18684=>"001010010",
  18685=>"110001111",
  18686=>"111111001",
  18687=>"110101101",
  18688=>"010111110",
  18689=>"110011000",
  18690=>"111001001",
  18691=>"000010000",
  18692=>"010000001",
  18693=>"000111100",
  18694=>"101000011",
  18695=>"101011000",
  18696=>"010011111",
  18697=>"001110111",
  18698=>"100011011",
  18699=>"101011101",
  18700=>"000001110",
  18701=>"101001111",
  18702=>"111011011",
  18703=>"111001100",
  18704=>"000110001",
  18705=>"100111010",
  18706=>"010101111",
  18707=>"110010101",
  18708=>"010110100",
  18709=>"111110001",
  18710=>"101100100",
  18711=>"001000000",
  18712=>"110000001",
  18713=>"100100000",
  18714=>"100100000",
  18715=>"110100010",
  18716=>"010011100",
  18717=>"111001010",
  18718=>"101101011",
  18719=>"000010011",
  18720=>"101100011",
  18721=>"100011011",
  18722=>"011100001",
  18723=>"010001000",
  18724=>"111011010",
  18725=>"011000100",
  18726=>"100111000",
  18727=>"000000111",
  18728=>"010110010",
  18729=>"111110111",
  18730=>"011010100",
  18731=>"111100100",
  18732=>"010111000",
  18733=>"001010000",
  18734=>"011011010",
  18735=>"100010001",
  18736=>"011101110",
  18737=>"010110100",
  18738=>"010111000",
  18739=>"001011101",
  18740=>"010101101",
  18741=>"010000011",
  18742=>"101000100",
  18743=>"011111001",
  18744=>"100110000",
  18745=>"000001000",
  18746=>"001000000",
  18747=>"110010111",
  18748=>"000110011",
  18749=>"011001011",
  18750=>"010001100",
  18751=>"101100101",
  18752=>"111010001",
  18753=>"100110111",
  18754=>"011110011",
  18755=>"001000100",
  18756=>"011110001",
  18757=>"011111100",
  18758=>"100010100",
  18759=>"010010111",
  18760=>"011101111",
  18761=>"011101111",
  18762=>"001110000",
  18763=>"001101101",
  18764=>"010100110",
  18765=>"011110000",
  18766=>"100000101",
  18767=>"011001111",
  18768=>"100111100",
  18769=>"011100101",
  18770=>"001111111",
  18771=>"001110011",
  18772=>"011110000",
  18773=>"111001000",
  18774=>"010110110",
  18775=>"100011001",
  18776=>"001101001",
  18777=>"101000000",
  18778=>"100001010",
  18779=>"011110010",
  18780=>"011110101",
  18781=>"010101011",
  18782=>"110011000",
  18783=>"111110010",
  18784=>"111110101",
  18785=>"000001000",
  18786=>"011111101",
  18787=>"000010011",
  18788=>"000111110",
  18789=>"100000010",
  18790=>"011101111",
  18791=>"011010110",
  18792=>"011110101",
  18793=>"011010110",
  18794=>"100011001",
  18795=>"001011000",
  18796=>"000111011",
  18797=>"110000010",
  18798=>"010111101",
  18799=>"010100000",
  18800=>"100101101",
  18801=>"001101101",
  18802=>"111101111",
  18803=>"010111101",
  18804=>"100110101",
  18805=>"000000011",
  18806=>"100110100",
  18807=>"010001101",
  18808=>"000010110",
  18809=>"010111000",
  18810=>"001101010",
  18811=>"011101011",
  18812=>"101001000",
  18813=>"001100010",
  18814=>"011011111",
  18815=>"110001010",
  18816=>"111011000",
  18817=>"010010000",
  18818=>"101111100",
  18819=>"100001110",
  18820=>"001101111",
  18821=>"101101111",
  18822=>"110101010",
  18823=>"000010000",
  18824=>"000001100",
  18825=>"110011000",
  18826=>"011001111",
  18827=>"010101011",
  18828=>"101101111",
  18829=>"101101011",
  18830=>"011110000",
  18831=>"110001011",
  18832=>"011111111",
  18833=>"110011010",
  18834=>"011010111",
  18835=>"001010000",
  18836=>"111011010",
  18837=>"010110001",
  18838=>"001100111",
  18839=>"000101001",
  18840=>"010100010",
  18841=>"001101100",
  18842=>"100000010",
  18843=>"111001101",
  18844=>"001010111",
  18845=>"101011101",
  18846=>"100110011",
  18847=>"001000000",
  18848=>"000011010",
  18849=>"101100110",
  18850=>"011111001",
  18851=>"000000001",
  18852=>"111110001",
  18853=>"100100011",
  18854=>"001010011",
  18855=>"000001011",
  18856=>"111001000",
  18857=>"111001000",
  18858=>"101010000",
  18859=>"011100111",
  18860=>"011011001",
  18861=>"111001010",
  18862=>"011000001",
  18863=>"000110101",
  18864=>"001000011",
  18865=>"100000110",
  18866=>"011000000",
  18867=>"111001001",
  18868=>"111011111",
  18869=>"101011011",
  18870=>"001111111",
  18871=>"110000111",
  18872=>"110001010",
  18873=>"110000000",
  18874=>"110001100",
  18875=>"100011111",
  18876=>"011000000",
  18877=>"001110000",
  18878=>"001110100",
  18879=>"011010101",
  18880=>"111000000",
  18881=>"101111110",
  18882=>"001010000",
  18883=>"000001000",
  18884=>"100110111",
  18885=>"000011010",
  18886=>"010010100",
  18887=>"101100100",
  18888=>"010101000",
  18889=>"010100111",
  18890=>"011010001",
  18891=>"000010100",
  18892=>"101001011",
  18893=>"110110101",
  18894=>"100110011",
  18895=>"010101001",
  18896=>"111100010",
  18897=>"000101100",
  18898=>"000011001",
  18899=>"011110101",
  18900=>"111010000",
  18901=>"100011100",
  18902=>"011011011",
  18903=>"101000000",
  18904=>"011110011",
  18905=>"011100101",
  18906=>"010101111",
  18907=>"000011100",
  18908=>"000101001",
  18909=>"110101010",
  18910=>"010010011",
  18911=>"111010011",
  18912=>"101101011",
  18913=>"111010011",
  18914=>"111010010",
  18915=>"000010010",
  18916=>"010111010",
  18917=>"011101111",
  18918=>"110001000",
  18919=>"111100001",
  18920=>"101001000",
  18921=>"111011111",
  18922=>"000010110",
  18923=>"110110110",
  18924=>"010000001",
  18925=>"111001010",
  18926=>"000001000",
  18927=>"011100000",
  18928=>"100110101",
  18929=>"101001010",
  18930=>"110101101",
  18931=>"011111001",
  18932=>"000010100",
  18933=>"001001100",
  18934=>"010000101",
  18935=>"100111110",
  18936=>"101111001",
  18937=>"111001100",
  18938=>"101111001",
  18939=>"100001110",
  18940=>"111110111",
  18941=>"001001011",
  18942=>"110001111",
  18943=>"010100000",
  18944=>"110000100",
  18945=>"100001110",
  18946=>"010001100",
  18947=>"111010010",
  18948=>"111101011",
  18949=>"111001011",
  18950=>"001101000",
  18951=>"000010010",
  18952=>"010110011",
  18953=>"000100110",
  18954=>"001110011",
  18955=>"011111000",
  18956=>"100000000",
  18957=>"101111010",
  18958=>"010010111",
  18959=>"011011110",
  18960=>"100001110",
  18961=>"001011110",
  18962=>"100111110",
  18963=>"000001101",
  18964=>"000100111",
  18965=>"111110101",
  18966=>"111010100",
  18967=>"011001000",
  18968=>"110001100",
  18969=>"001111001",
  18970=>"011000001",
  18971=>"011001111",
  18972=>"111011101",
  18973=>"011001111",
  18974=>"101001011",
  18975=>"101100111",
  18976=>"100010010",
  18977=>"110100000",
  18978=>"001000111",
  18979=>"000010100",
  18980=>"100100110",
  18981=>"000011011",
  18982=>"111101111",
  18983=>"000101101",
  18984=>"001001000",
  18985=>"010101011",
  18986=>"101011101",
  18987=>"000000000",
  18988=>"111110011",
  18989=>"101111000",
  18990=>"011010010",
  18991=>"011000000",
  18992=>"000100001",
  18993=>"101111010",
  18994=>"100001010",
  18995=>"111100000",
  18996=>"010101110",
  18997=>"101100111",
  18998=>"110010110",
  18999=>"110010010",
  19000=>"000010110",
  19001=>"100001101",
  19002=>"000111000",
  19003=>"011110101",
  19004=>"010111101",
  19005=>"110010000",
  19006=>"000001001",
  19007=>"111011010",
  19008=>"100010101",
  19009=>"100000110",
  19010=>"100010010",
  19011=>"101111101",
  19012=>"010111000",
  19013=>"110111110",
  19014=>"010011100",
  19015=>"101101101",
  19016=>"101111110",
  19017=>"010110111",
  19018=>"001101010",
  19019=>"110000100",
  19020=>"011100010",
  19021=>"010001110",
  19022=>"100011010",
  19023=>"110110111",
  19024=>"001110111",
  19025=>"110110010",
  19026=>"110010001",
  19027=>"011100001",
  19028=>"101001100",
  19029=>"001101101",
  19030=>"000110010",
  19031=>"001001111",
  19032=>"011011010",
  19033=>"000001001",
  19034=>"011111110",
  19035=>"010010010",
  19036=>"101000110",
  19037=>"110001011",
  19038=>"001000100",
  19039=>"111001100",
  19040=>"011001011",
  19041=>"010001000",
  19042=>"000000000",
  19043=>"011010000",
  19044=>"111011101",
  19045=>"101010100",
  19046=>"101110000",
  19047=>"111100111",
  19048=>"000000001",
  19049=>"101010101",
  19050=>"011110001",
  19051=>"010001000",
  19052=>"110010110",
  19053=>"011110111",
  19054=>"000001011",
  19055=>"000010101",
  19056=>"001100000",
  19057=>"011010000",
  19058=>"010001001",
  19059=>"011000111",
  19060=>"111011010",
  19061=>"001001011",
  19062=>"110100100",
  19063=>"100111111",
  19064=>"001100110",
  19065=>"110110100",
  19066=>"101011011",
  19067=>"000111101",
  19068=>"101000000",
  19069=>"000100000",
  19070=>"010111011",
  19071=>"000100101",
  19072=>"000010000",
  19073=>"111110000",
  19074=>"100111001",
  19075=>"000010010",
  19076=>"001110111",
  19077=>"101001001",
  19078=>"001111111",
  19079=>"010000110",
  19080=>"101101000",
  19081=>"111010000",
  19082=>"100001111",
  19083=>"011011011",
  19084=>"011111000",
  19085=>"001111100",
  19086=>"110111001",
  19087=>"100100101",
  19088=>"001000101",
  19089=>"111101100",
  19090=>"101101110",
  19091=>"101110100",
  19092=>"101111110",
  19093=>"010110011",
  19094=>"010111110",
  19095=>"101001110",
  19096=>"000111111",
  19097=>"010100011",
  19098=>"100001111",
  19099=>"001110100",
  19100=>"101000101",
  19101=>"111100100",
  19102=>"101100000",
  19103=>"000011000",
  19104=>"111001011",
  19105=>"010100111",
  19106=>"101111101",
  19107=>"001001111",
  19108=>"011011000",
  19109=>"111010111",
  19110=>"001000000",
  19111=>"101100111",
  19112=>"001101001",
  19113=>"000011001",
  19114=>"110100101",
  19115=>"011101101",
  19116=>"000101010",
  19117=>"110011000",
  19118=>"100010101",
  19119=>"111001010",
  19120=>"101101010",
  19121=>"000010111",
  19122=>"100011101",
  19123=>"011111100",
  19124=>"010000110",
  19125=>"111000010",
  19126=>"011010101",
  19127=>"110000110",
  19128=>"011010001",
  19129=>"000001100",
  19130=>"111111110",
  19131=>"110111101",
  19132=>"111111000",
  19133=>"101000001",
  19134=>"000010010",
  19135=>"011110010",
  19136=>"001011101",
  19137=>"011111010",
  19138=>"000001101",
  19139=>"101101000",
  19140=>"001010101",
  19141=>"001101000",
  19142=>"101101000",
  19143=>"101110011",
  19144=>"011111000",
  19145=>"011110000",
  19146=>"010101010",
  19147=>"101000000",
  19148=>"011000010",
  19149=>"000011110",
  19150=>"000110001",
  19151=>"111110111",
  19152=>"010001001",
  19153=>"010101110",
  19154=>"100101000",
  19155=>"111010100",
  19156=>"111001110",
  19157=>"001000010",
  19158=>"100000100",
  19159=>"000110100",
  19160=>"101110000",
  19161=>"101001111",
  19162=>"110001100",
  19163=>"101010111",
  19164=>"000100011",
  19165=>"000000000",
  19166=>"110010010",
  19167=>"010100111",
  19168=>"000100010",
  19169=>"001101000",
  19170=>"111010010",
  19171=>"110010110",
  19172=>"000011001",
  19173=>"110111011",
  19174=>"010111001",
  19175=>"111101010",
  19176=>"011111000",
  19177=>"101011010",
  19178=>"000010010",
  19179=>"100100001",
  19180=>"000000110",
  19181=>"000010100",
  19182=>"100010111",
  19183=>"111011001",
  19184=>"101101111",
  19185=>"011101101",
  19186=>"100110110",
  19187=>"100010001",
  19188=>"000110000",
  19189=>"010011111",
  19190=>"000110100",
  19191=>"110101000",
  19192=>"010000001",
  19193=>"010101111",
  19194=>"000101110",
  19195=>"100001001",
  19196=>"110111111",
  19197=>"000010000",
  19198=>"010001001",
  19199=>"010000000",
  19200=>"101110000",
  19201=>"001101000",
  19202=>"110100111",
  19203=>"010010111",
  19204=>"111111011",
  19205=>"010100111",
  19206=>"010011001",
  19207=>"110111110",
  19208=>"000001011",
  19209=>"111101100",
  19210=>"111000000",
  19211=>"111011010",
  19212=>"110101110",
  19213=>"000110010",
  19214=>"110111011",
  19215=>"001010011",
  19216=>"000010111",
  19217=>"101011010",
  19218=>"110000100",
  19219=>"010111000",
  19220=>"000000000",
  19221=>"111000100",
  19222=>"101000000",
  19223=>"100011000",
  19224=>"111100000",
  19225=>"111010000",
  19226=>"101101101",
  19227=>"110100000",
  19228=>"101001011",
  19229=>"111101001",
  19230=>"010001001",
  19231=>"110101100",
  19232=>"111000100",
  19233=>"111101100",
  19234=>"101010111",
  19235=>"010100001",
  19236=>"001001111",
  19237=>"011100010",
  19238=>"010111111",
  19239=>"100000000",
  19240=>"100111111",
  19241=>"111001011",
  19242=>"111111101",
  19243=>"001101110",
  19244=>"101011011",
  19245=>"001000011",
  19246=>"011110000",
  19247=>"000100100",
  19248=>"110010110",
  19249=>"001001010",
  19250=>"101110100",
  19251=>"101111111",
  19252=>"000010010",
  19253=>"110000001",
  19254=>"010010110",
  19255=>"111111110",
  19256=>"000001100",
  19257=>"010000101",
  19258=>"000001000",
  19259=>"101101110",
  19260=>"111011000",
  19261=>"111111101",
  19262=>"101011111",
  19263=>"101100100",
  19264=>"000000100",
  19265=>"100101010",
  19266=>"101100100",
  19267=>"110001100",
  19268=>"101000010",
  19269=>"101010100",
  19270=>"110010000",
  19271=>"011010110",
  19272=>"100000101",
  19273=>"000010100",
  19274=>"100001000",
  19275=>"000000000",
  19276=>"111001111",
  19277=>"001001000",
  19278=>"011110000",
  19279=>"010100010",
  19280=>"111010100",
  19281=>"110000010",
  19282=>"010111111",
  19283=>"101010000",
  19284=>"101101100",
  19285=>"000100110",
  19286=>"100101011",
  19287=>"001011110",
  19288=>"000010101",
  19289=>"000101010",
  19290=>"100000100",
  19291=>"101101010",
  19292=>"110110000",
  19293=>"010000111",
  19294=>"110010011",
  19295=>"110010001",
  19296=>"100010011",
  19297=>"110110111",
  19298=>"100010101",
  19299=>"110101011",
  19300=>"000010010",
  19301=>"101000110",
  19302=>"110111001",
  19303=>"100010010",
  19304=>"010010000",
  19305=>"111110111",
  19306=>"011010100",
  19307=>"001000010",
  19308=>"101111000",
  19309=>"110011001",
  19310=>"010111001",
  19311=>"111110000",
  19312=>"100001000",
  19313=>"101010000",
  19314=>"111100001",
  19315=>"100100000",
  19316=>"100101111",
  19317=>"110111010",
  19318=>"100110100",
  19319=>"111000011",
  19320=>"100100111",
  19321=>"010000000",
  19322=>"110001001",
  19323=>"111001011",
  19324=>"000000001",
  19325=>"001001000",
  19326=>"111100101",
  19327=>"000011110",
  19328=>"100000000",
  19329=>"111010111",
  19330=>"001100001",
  19331=>"101010000",
  19332=>"101001011",
  19333=>"000010111",
  19334=>"110111000",
  19335=>"001100100",
  19336=>"001111110",
  19337=>"110111111",
  19338=>"001010000",
  19339=>"101110000",
  19340=>"000011101",
  19341=>"110000000",
  19342=>"010100011",
  19343=>"100100101",
  19344=>"010000010",
  19345=>"011000011",
  19346=>"011010000",
  19347=>"001010011",
  19348=>"110000100",
  19349=>"001011110",
  19350=>"111001101",
  19351=>"010111010",
  19352=>"110110110",
  19353=>"110011110",
  19354=>"110010001",
  19355=>"010101101",
  19356=>"111100111",
  19357=>"111101010",
  19358=>"001100111",
  19359=>"111000010",
  19360=>"101001011",
  19361=>"011011010",
  19362=>"101101011",
  19363=>"100111001",
  19364=>"001011101",
  19365=>"110101010",
  19366=>"000110110",
  19367=>"011010001",
  19368=>"111000110",
  19369=>"000010000",
  19370=>"010001000",
  19371=>"000000101",
  19372=>"011100011",
  19373=>"100001011",
  19374=>"110001101",
  19375=>"000001100",
  19376=>"111100111",
  19377=>"011000110",
  19378=>"010001001",
  19379=>"010011001",
  19380=>"010001111",
  19381=>"000110010",
  19382=>"111111100",
  19383=>"011011101",
  19384=>"001010101",
  19385=>"111000000",
  19386=>"111001111",
  19387=>"000000001",
  19388=>"000111000",
  19389=>"110000100",
  19390=>"101111101",
  19391=>"000000000",
  19392=>"010011001",
  19393=>"110010000",
  19394=>"100010001",
  19395=>"110110101",
  19396=>"111011010",
  19397=>"110111000",
  19398=>"111100000",
  19399=>"100110001",
  19400=>"000100110",
  19401=>"010001011",
  19402=>"101001001",
  19403=>"111111010",
  19404=>"100010010",
  19405=>"001000110",
  19406=>"101000010",
  19407=>"101011001",
  19408=>"010110101",
  19409=>"100010100",
  19410=>"000100110",
  19411=>"011111101",
  19412=>"011110011",
  19413=>"110011110",
  19414=>"001101010",
  19415=>"010110101",
  19416=>"100100100",
  19417=>"010000111",
  19418=>"111111111",
  19419=>"000100110",
  19420=>"111011101",
  19421=>"100110101",
  19422=>"101000111",
  19423=>"100001111",
  19424=>"101101011",
  19425=>"000001111",
  19426=>"001000101",
  19427=>"001001011",
  19428=>"101011010",
  19429=>"111101100",
  19430=>"110101000",
  19431=>"110110011",
  19432=>"001110100",
  19433=>"110111000",
  19434=>"000001010",
  19435=>"101000100",
  19436=>"111111101",
  19437=>"110110010",
  19438=>"001010010",
  19439=>"100110001",
  19440=>"100111110",
  19441=>"111010001",
  19442=>"011111110",
  19443=>"001010111",
  19444=>"011000010",
  19445=>"111011101",
  19446=>"000110010",
  19447=>"101010001",
  19448=>"000100101",
  19449=>"000010001",
  19450=>"011100100",
  19451=>"000011111",
  19452=>"010111000",
  19453=>"100110011",
  19454=>"111111111",
  19455=>"111111101",
  19456=>"011000110",
  19457=>"101110001",
  19458=>"001100011",
  19459=>"010011000",
  19460=>"111110101",
  19461=>"010001110",
  19462=>"101110110",
  19463=>"110000000",
  19464=>"010010110",
  19465=>"110110101",
  19466=>"101001101",
  19467=>"101111010",
  19468=>"100111100",
  19469=>"001010000",
  19470=>"111010011",
  19471=>"110001001",
  19472=>"000010000",
  19473=>"000010001",
  19474=>"010010111",
  19475=>"100111100",
  19476=>"000101011",
  19477=>"000001000",
  19478=>"111101010",
  19479=>"010100011",
  19480=>"011100100",
  19481=>"010000001",
  19482=>"000110110",
  19483=>"000001001",
  19484=>"111111110",
  19485=>"000110000",
  19486=>"100110000",
  19487=>"101111110",
  19488=>"011010011",
  19489=>"100010010",
  19490=>"010101101",
  19491=>"011010000",
  19492=>"011010011",
  19493=>"000010110",
  19494=>"001000100",
  19495=>"011010011",
  19496=>"011101010",
  19497=>"011101000",
  19498=>"101000110",
  19499=>"000101100",
  19500=>"000111000",
  19501=>"000101110",
  19502=>"000001000",
  19503=>"011100101",
  19504=>"111001101",
  19505=>"011000110",
  19506=>"101001100",
  19507=>"110011000",
  19508=>"110101001",
  19509=>"000111011",
  19510=>"001001001",
  19511=>"011001111",
  19512=>"000100110",
  19513=>"000001010",
  19514=>"101100110",
  19515=>"000100011",
  19516=>"010011110",
  19517=>"111111010",
  19518=>"111111010",
  19519=>"010000010",
  19520=>"010000000",
  19521=>"101010010",
  19522=>"001011011",
  19523=>"000110000",
  19524=>"000001001",
  19525=>"011000011",
  19526=>"111100001",
  19527=>"000010100",
  19528=>"111111001",
  19529=>"011010101",
  19530=>"000001010",
  19531=>"000101101",
  19532=>"010111100",
  19533=>"111100100",
  19534=>"110101111",
  19535=>"000111011",
  19536=>"101001011",
  19537=>"010101111",
  19538=>"111000000",
  19539=>"101101000",
  19540=>"100100100",
  19541=>"101111010",
  19542=>"000000011",
  19543=>"011110101",
  19544=>"110000000",
  19545=>"111101011",
  19546=>"101011000",
  19547=>"011000010",
  19548=>"111110111",
  19549=>"000101000",
  19550=>"000000110",
  19551=>"000011111",
  19552=>"101111001",
  19553=>"101000001",
  19554=>"101001111",
  19555=>"000011110",
  19556=>"100111101",
  19557=>"011101000",
  19558=>"000010011",
  19559=>"101001111",
  19560=>"011110000",
  19561=>"101001000",
  19562=>"010011101",
  19563=>"111010110",
  19564=>"000110101",
  19565=>"100010000",
  19566=>"100111010",
  19567=>"110000010",
  19568=>"111100100",
  19569=>"000101110",
  19570=>"000100010",
  19571=>"010101111",
  19572=>"111000110",
  19573=>"000111111",
  19574=>"000100111",
  19575=>"100001010",
  19576=>"000110100",
  19577=>"011000001",
  19578=>"110001010",
  19579=>"011100111",
  19580=>"011000011",
  19581=>"101011100",
  19582=>"111011111",
  19583=>"001100001",
  19584=>"110000110",
  19585=>"001001001",
  19586=>"100100011",
  19587=>"100101010",
  19588=>"101111110",
  19589=>"110111001",
  19590=>"101010010",
  19591=>"011001110",
  19592=>"110110010",
  19593=>"110011011",
  19594=>"001001000",
  19595=>"000000011",
  19596=>"001011000",
  19597=>"101100111",
  19598=>"000000100",
  19599=>"100111000",
  19600=>"100100111",
  19601=>"111011000",
  19602=>"100010001",
  19603=>"011001000",
  19604=>"100101011",
  19605=>"111001011",
  19606=>"001000000",
  19607=>"011000000",
  19608=>"101001010",
  19609=>"111001000",
  19610=>"100100111",
  19611=>"110101101",
  19612=>"000000010",
  19613=>"011001101",
  19614=>"111100101",
  19615=>"010001001",
  19616=>"001110110",
  19617=>"111100001",
  19618=>"111000001",
  19619=>"110101100",
  19620=>"111010011",
  19621=>"111011111",
  19622=>"100011010",
  19623=>"100111000",
  19624=>"000110101",
  19625=>"100011110",
  19626=>"110100101",
  19627=>"101101101",
  19628=>"100110000",
  19629=>"111011000",
  19630=>"001001110",
  19631=>"100100110",
  19632=>"110100111",
  19633=>"100101111",
  19634=>"000101111",
  19635=>"100101000",
  19636=>"101111110",
  19637=>"001000011",
  19638=>"110011001",
  19639=>"000000011",
  19640=>"000010000",
  19641=>"110001110",
  19642=>"101100110",
  19643=>"011000110",
  19644=>"010011010",
  19645=>"011110010",
  19646=>"010110000",
  19647=>"111111000",
  19648=>"001001001",
  19649=>"010111001",
  19650=>"011110000",
  19651=>"110011110",
  19652=>"000111100",
  19653=>"101001010",
  19654=>"101100001",
  19655=>"111101110",
  19656=>"010100111",
  19657=>"011111100",
  19658=>"011100100",
  19659=>"000111010",
  19660=>"001001111",
  19661=>"110011111",
  19662=>"000110001",
  19663=>"010000001",
  19664=>"001110101",
  19665=>"110101101",
  19666=>"100001111",
  19667=>"100000100",
  19668=>"000010100",
  19669=>"110111001",
  19670=>"111101100",
  19671=>"001000111",
  19672=>"101011000",
  19673=>"111111100",
  19674=>"101001110",
  19675=>"100111000",
  19676=>"111100001",
  19677=>"010010110",
  19678=>"001001101",
  19679=>"111100111",
  19680=>"100110111",
  19681=>"100011000",
  19682=>"000010110",
  19683=>"000100110",
  19684=>"110111111",
  19685=>"100000100",
  19686=>"101101100",
  19687=>"001101110",
  19688=>"111000000",
  19689=>"010001011",
  19690=>"010010000",
  19691=>"101100011",
  19692=>"111101010",
  19693=>"011001000",
  19694=>"101111101",
  19695=>"111000101",
  19696=>"110110111",
  19697=>"001111011",
  19698=>"110100000",
  19699=>"101010110",
  19700=>"100000010",
  19701=>"101111111",
  19702=>"001011011",
  19703=>"100000011",
  19704=>"011110011",
  19705=>"110010000",
  19706=>"100001100",
  19707=>"010100010",
  19708=>"101001110",
  19709=>"010111001",
  19710=>"100000000",
  19711=>"100111101",
  19712=>"001011111",
  19713=>"000000111",
  19714=>"110100001",
  19715=>"110100000",
  19716=>"010101100",
  19717=>"101010111",
  19718=>"001011110",
  19719=>"101101111",
  19720=>"010100111",
  19721=>"111101111",
  19722=>"000000101",
  19723=>"010101100",
  19724=>"101100010",
  19725=>"000010100",
  19726=>"011100110",
  19727=>"110110111",
  19728=>"000001111",
  19729=>"011111010",
  19730=>"101001011",
  19731=>"110010101",
  19732=>"101101110",
  19733=>"111110011",
  19734=>"000110001",
  19735=>"100000110",
  19736=>"001110100",
  19737=>"011101011",
  19738=>"011101101",
  19739=>"101110100",
  19740=>"011000011",
  19741=>"011110110",
  19742=>"110110011",
  19743=>"100101010",
  19744=>"001101101",
  19745=>"110111101",
  19746=>"110100101",
  19747=>"110100101",
  19748=>"011111000",
  19749=>"010111110",
  19750=>"000100010",
  19751=>"001010001",
  19752=>"110011001",
  19753=>"000001111",
  19754=>"101011001",
  19755=>"001001000",
  19756=>"001011110",
  19757=>"010000111",
  19758=>"111000000",
  19759=>"100111100",
  19760=>"110111100",
  19761=>"011000010",
  19762=>"011000110",
  19763=>"000111011",
  19764=>"111111110",
  19765=>"010101110",
  19766=>"101110001",
  19767=>"101101011",
  19768=>"111110100",
  19769=>"111111110",
  19770=>"010111001",
  19771=>"011100000",
  19772=>"010100000",
  19773=>"001101100",
  19774=>"111000111",
  19775=>"101110001",
  19776=>"110000001",
  19777=>"101100010",
  19778=>"100101001",
  19779=>"110111000",
  19780=>"100010010",
  19781=>"100001110",
  19782=>"101000000",
  19783=>"000010100",
  19784=>"011000110",
  19785=>"010001111",
  19786=>"000010000",
  19787=>"001111100",
  19788=>"110001000",
  19789=>"000001011",
  19790=>"111011100",
  19791=>"010110110",
  19792=>"001101000",
  19793=>"101011110",
  19794=>"110101011",
  19795=>"000010100",
  19796=>"111000110",
  19797=>"000011010",
  19798=>"001110011",
  19799=>"010100000",
  19800=>"000110101",
  19801=>"111101101",
  19802=>"100110101",
  19803=>"010001001",
  19804=>"011011101",
  19805=>"100000111",
  19806=>"010001000",
  19807=>"001100100",
  19808=>"001001000",
  19809=>"011001011",
  19810=>"011101000",
  19811=>"111100000",
  19812=>"010100101",
  19813=>"010100010",
  19814=>"000010111",
  19815=>"101010001",
  19816=>"110010000",
  19817=>"011010001",
  19818=>"101100101",
  19819=>"011100010",
  19820=>"010000000",
  19821=>"010011101",
  19822=>"110100001",
  19823=>"101110010",
  19824=>"000000101",
  19825=>"001000011",
  19826=>"000001110",
  19827=>"100010101",
  19828=>"110001001",
  19829=>"010101011",
  19830=>"101101101",
  19831=>"001110001",
  19832=>"100110011",
  19833=>"111100011",
  19834=>"010100000",
  19835=>"110101110",
  19836=>"101010000",
  19837=>"010010011",
  19838=>"111110001",
  19839=>"100010100",
  19840=>"101010010",
  19841=>"100010010",
  19842=>"101001101",
  19843=>"011110101",
  19844=>"010111101",
  19845=>"101001101",
  19846=>"100010011",
  19847=>"001111000",
  19848=>"011110110",
  19849=>"011000010",
  19850=>"101000001",
  19851=>"111011010",
  19852=>"001101010",
  19853=>"101100010",
  19854=>"011010000",
  19855=>"101111100",
  19856=>"011000000",
  19857=>"110100101",
  19858=>"110001100",
  19859=>"110000011",
  19860=>"011000101",
  19861=>"110111011",
  19862=>"100101001",
  19863=>"100101110",
  19864=>"000101110",
  19865=>"011010010",
  19866=>"110101101",
  19867=>"110110000",
  19868=>"000001001",
  19869=>"110111000",
  19870=>"000011111",
  19871=>"010110100",
  19872=>"111101100",
  19873=>"111010110",
  19874=>"111001001",
  19875=>"001100101",
  19876=>"100111000",
  19877=>"111100110",
  19878=>"100011011",
  19879=>"110101110",
  19880=>"000110011",
  19881=>"001101001",
  19882=>"100101111",
  19883=>"011101011",
  19884=>"000000001",
  19885=>"000111001",
  19886=>"110101110",
  19887=>"010100001",
  19888=>"101010001",
  19889=>"110000010",
  19890=>"011101100",
  19891=>"100011000",
  19892=>"000001001",
  19893=>"111100111",
  19894=>"010111110",
  19895=>"000011101",
  19896=>"010001110",
  19897=>"000111000",
  19898=>"110001010",
  19899=>"000011011",
  19900=>"010011010",
  19901=>"011010001",
  19902=>"101101001",
  19903=>"100000000",
  19904=>"101001111",
  19905=>"011100110",
  19906=>"001001110",
  19907=>"111011010",
  19908=>"101111010",
  19909=>"111000110",
  19910=>"110100000",
  19911=>"011101010",
  19912=>"111001110",
  19913=>"001011100",
  19914=>"111101110",
  19915=>"111111110",
  19916=>"001011101",
  19917=>"101101000",
  19918=>"100101110",
  19919=>"000001101",
  19920=>"100010110",
  19921=>"000111101",
  19922=>"111011000",
  19923=>"010101101",
  19924=>"001011111",
  19925=>"011101001",
  19926=>"011011100",
  19927=>"100001000",
  19928=>"111010001",
  19929=>"110011101",
  19930=>"101110011",
  19931=>"111011100",
  19932=>"001111011",
  19933=>"111000100",
  19934=>"001110101",
  19935=>"001101111",
  19936=>"000000001",
  19937=>"001100001",
  19938=>"000010001",
  19939=>"001000111",
  19940=>"100101010",
  19941=>"100000100",
  19942=>"111001000",
  19943=>"111001110",
  19944=>"000010001",
  19945=>"100111101",
  19946=>"101010111",
  19947=>"111000110",
  19948=>"111111110",
  19949=>"010011111",
  19950=>"011010010",
  19951=>"100100001",
  19952=>"010000100",
  19953=>"001111010",
  19954=>"111100101",
  19955=>"011110110",
  19956=>"011000011",
  19957=>"001110010",
  19958=>"010111101",
  19959=>"000110110",
  19960=>"110111100",
  19961=>"111111000",
  19962=>"000101000",
  19963=>"011111111",
  19964=>"000111010",
  19965=>"100110001",
  19966=>"101010001",
  19967=>"110001111",
  19968=>"001111110",
  19969=>"010111001",
  19970=>"101001110",
  19971=>"111001100",
  19972=>"100100000",
  19973=>"000000111",
  19974=>"111100100",
  19975=>"101010111",
  19976=>"101110010",
  19977=>"000000100",
  19978=>"011110110",
  19979=>"101000001",
  19980=>"000011110",
  19981=>"010000010",
  19982=>"011100101",
  19983=>"101100011",
  19984=>"001011110",
  19985=>"101110100",
  19986=>"100110101",
  19987=>"100101110",
  19988=>"110100000",
  19989=>"010000000",
  19990=>"110010111",
  19991=>"001001010",
  19992=>"100101010",
  19993=>"001111001",
  19994=>"110001001",
  19995=>"111101010",
  19996=>"011100001",
  19997=>"110110100",
  19998=>"100100000",
  19999=>"000110101",
  20000=>"000101111",
  20001=>"110100000",
  20002=>"001000101",
  20003=>"111010100",
  20004=>"110111110",
  20005=>"010111000",
  20006=>"001110111",
  20007=>"111001011",
  20008=>"000001101",
  20009=>"100110110",
  20010=>"000101101",
  20011=>"110011001",
  20012=>"001110010",
  20013=>"001000101",
  20014=>"001100001",
  20015=>"110110110",
  20016=>"101000001",
  20017=>"111110010",
  20018=>"100000111",
  20019=>"001001010",
  20020=>"110000111",
  20021=>"101110110",
  20022=>"000001010",
  20023=>"001110010",
  20024=>"010001101",
  20025=>"010000011",
  20026=>"101000101",
  20027=>"000100000",
  20028=>"101001010",
  20029=>"101010010",
  20030=>"000010111",
  20031=>"111010010",
  20032=>"101110110",
  20033=>"101011101",
  20034=>"100000001",
  20035=>"010000011",
  20036=>"100001110",
  20037=>"111001001",
  20038=>"000011000",
  20039=>"011111110",
  20040=>"011100010",
  20041=>"011100101",
  20042=>"110111101",
  20043=>"000010100",
  20044=>"001011101",
  20045=>"100111100",
  20046=>"111011000",
  20047=>"111000101",
  20048=>"100001010",
  20049=>"110000010",
  20050=>"000010010",
  20051=>"011001000",
  20052=>"110101010",
  20053=>"010100000",
  20054=>"110011101",
  20055=>"001100101",
  20056=>"110000010",
  20057=>"001110010",
  20058=>"010101100",
  20059=>"010101011",
  20060=>"011101111",
  20061=>"001000101",
  20062=>"101001110",
  20063=>"101111001",
  20064=>"000000101",
  20065=>"010000111",
  20066=>"001111100",
  20067=>"011001001",
  20068=>"000001010",
  20069=>"110010010",
  20070=>"101011111",
  20071=>"101000111",
  20072=>"110001011",
  20073=>"110111010",
  20074=>"010101111",
  20075=>"100001100",
  20076=>"110100011",
  20077=>"001101101",
  20078=>"010011101",
  20079=>"101011010",
  20080=>"111110000",
  20081=>"101001101",
  20082=>"001011111",
  20083=>"100001001",
  20084=>"010101101",
  20085=>"010000101",
  20086=>"100000000",
  20087=>"000111110",
  20088=>"100010010",
  20089=>"011010000",
  20090=>"111110011",
  20091=>"110101001",
  20092=>"001010010",
  20093=>"000101001",
  20094=>"001000110",
  20095=>"011100010",
  20096=>"110110001",
  20097=>"010110001",
  20098=>"111101101",
  20099=>"101101100",
  20100=>"011011010",
  20101=>"110000100",
  20102=>"010111110",
  20103=>"001110001",
  20104=>"101001100",
  20105=>"011100010",
  20106=>"001010000",
  20107=>"010001111",
  20108=>"111011101",
  20109=>"010011100",
  20110=>"001010001",
  20111=>"000110100",
  20112=>"011000100",
  20113=>"101000110",
  20114=>"001101001",
  20115=>"011001111",
  20116=>"010100111",
  20117=>"110011101",
  20118=>"101101111",
  20119=>"011100011",
  20120=>"110101111",
  20121=>"001001101",
  20122=>"010011111",
  20123=>"011111101",
  20124=>"110000100",
  20125=>"101011001",
  20126=>"000100111",
  20127=>"011101011",
  20128=>"000101100",
  20129=>"011011111",
  20130=>"101001001",
  20131=>"101111000",
  20132=>"110110001",
  20133=>"110100100",
  20134=>"000001110",
  20135=>"100100011",
  20136=>"010111010",
  20137=>"001100010",
  20138=>"100100011",
  20139=>"101000000",
  20140=>"100010010",
  20141=>"011000100",
  20142=>"010000011",
  20143=>"110001001",
  20144=>"100111000",
  20145=>"000110011",
  20146=>"101000000",
  20147=>"101000011",
  20148=>"100010111",
  20149=>"100111001",
  20150=>"100001101",
  20151=>"100100100",
  20152=>"101100010",
  20153=>"000101001",
  20154=>"000000001",
  20155=>"100000110",
  20156=>"000001101",
  20157=>"101010010",
  20158=>"000100000",
  20159=>"110010001",
  20160=>"100011001",
  20161=>"111111010",
  20162=>"100010010",
  20163=>"100101010",
  20164=>"100110010",
  20165=>"001011111",
  20166=>"101110010",
  20167=>"110110000",
  20168=>"111010011",
  20169=>"001011101",
  20170=>"010100000",
  20171=>"110101110",
  20172=>"100010010",
  20173=>"100110111",
  20174=>"001010101",
  20175=>"000110000",
  20176=>"010000111",
  20177=>"010010000",
  20178=>"111011111",
  20179=>"000010101",
  20180=>"001100010",
  20181=>"000100011",
  20182=>"100111101",
  20183=>"100000101",
  20184=>"001010110",
  20185=>"001000001",
  20186=>"010100101",
  20187=>"001000011",
  20188=>"010101011",
  20189=>"001001110",
  20190=>"111100111",
  20191=>"110110101",
  20192=>"000000001",
  20193=>"111010101",
  20194=>"010110001",
  20195=>"001001100",
  20196=>"100000001",
  20197=>"100111111",
  20198=>"101100100",
  20199=>"000110000",
  20200=>"001010000",
  20201=>"011110110",
  20202=>"001010111",
  20203=>"000111010",
  20204=>"000100100",
  20205=>"101000110",
  20206=>"011011000",
  20207=>"000110111",
  20208=>"100111000",
  20209=>"101100000",
  20210=>"011110111",
  20211=>"000100010",
  20212=>"111101011",
  20213=>"000000000",
  20214=>"001110000",
  20215=>"010101001",
  20216=>"011110101",
  20217=>"000110110",
  20218=>"011010101",
  20219=>"011000000",
  20220=>"000111111",
  20221=>"110111111",
  20222=>"011110000",
  20223=>"001000101",
  20224=>"100011000",
  20225=>"000100100",
  20226=>"001011000",
  20227=>"001010101",
  20228=>"110101100",
  20229=>"010110001",
  20230=>"001011001",
  20231=>"010000100",
  20232=>"000000000",
  20233=>"000000111",
  20234=>"101111010",
  20235=>"011011111",
  20236=>"011000100",
  20237=>"101101100",
  20238=>"000101100",
  20239=>"001001101",
  20240=>"100010101",
  20241=>"011101011",
  20242=>"110110110",
  20243=>"111011101",
  20244=>"001111100",
  20245=>"011001001",
  20246=>"101011000",
  20247=>"110110111",
  20248=>"001000111",
  20249=>"000110001",
  20250=>"001100110",
  20251=>"101110001",
  20252=>"100000100",
  20253=>"111111100",
  20254=>"011010000",
  20255=>"011111011",
  20256=>"110010100",
  20257=>"000000011",
  20258=>"110101000",
  20259=>"000101000",
  20260=>"011001100",
  20261=>"111101111",
  20262=>"000101100",
  20263=>"101010011",
  20264=>"000001101",
  20265=>"011000110",
  20266=>"010111000",
  20267=>"110011001",
  20268=>"000010001",
  20269=>"011101011",
  20270=>"101010100",
  20271=>"110110001",
  20272=>"101001111",
  20273=>"001101000",
  20274=>"010010110",
  20275=>"110100110",
  20276=>"011001110",
  20277=>"100000111",
  20278=>"111100001",
  20279=>"010000000",
  20280=>"101111001",
  20281=>"011010110",
  20282=>"000110000",
  20283=>"110011101",
  20284=>"011101110",
  20285=>"101101010",
  20286=>"000000110",
  20287=>"100001001",
  20288=>"110111101",
  20289=>"011111101",
  20290=>"111110101",
  20291=>"101001100",
  20292=>"111010000",
  20293=>"000100011",
  20294=>"100010001",
  20295=>"101010000",
  20296=>"101100100",
  20297=>"111100100",
  20298=>"011110110",
  20299=>"010100000",
  20300=>"010110110",
  20301=>"011000010",
  20302=>"111111100",
  20303=>"100010100",
  20304=>"001000000",
  20305=>"010000101",
  20306=>"101010100",
  20307=>"001101010",
  20308=>"000100011",
  20309=>"000000101",
  20310=>"010000010",
  20311=>"010011111",
  20312=>"011000000",
  20313=>"101100111",
  20314=>"100001001",
  20315=>"110101000",
  20316=>"111101011",
  20317=>"101011111",
  20318=>"110110100",
  20319=>"100111010",
  20320=>"101111100",
  20321=>"010010001",
  20322=>"111100000",
  20323=>"000001110",
  20324=>"001111000",
  20325=>"011100111",
  20326=>"100100001",
  20327=>"000111000",
  20328=>"111010110",
  20329=>"000000011",
  20330=>"101000011",
  20331=>"000110000",
  20332=>"011000100",
  20333=>"100000001",
  20334=>"001001111",
  20335=>"111111100",
  20336=>"111010000",
  20337=>"110100000",
  20338=>"100010011",
  20339=>"000000101",
  20340=>"111001001",
  20341=>"000000000",
  20342=>"011010000",
  20343=>"000110100",
  20344=>"111000010",
  20345=>"111110110",
  20346=>"101111101",
  20347=>"001010100",
  20348=>"110000100",
  20349=>"011000101",
  20350=>"111100000",
  20351=>"110011010",
  20352=>"100110111",
  20353=>"110000010",
  20354=>"001000000",
  20355=>"011000111",
  20356=>"101010100",
  20357=>"000111011",
  20358=>"111111011",
  20359=>"110000100",
  20360=>"010111100",
  20361=>"001110101",
  20362=>"010000011",
  20363=>"100011000",
  20364=>"001011011",
  20365=>"110001000",
  20366=>"001010110",
  20367=>"101010100",
  20368=>"101111101",
  20369=>"100111111",
  20370=>"110001010",
  20371=>"111111000",
  20372=>"010011000",
  20373=>"110001100",
  20374=>"011011100",
  20375=>"010110011",
  20376=>"100111100",
  20377=>"110100111",
  20378=>"001011101",
  20379=>"100100110",
  20380=>"011101101",
  20381=>"000101110",
  20382=>"111010100",
  20383=>"100001100",
  20384=>"000000101",
  20385=>"011111110",
  20386=>"101001010",
  20387=>"111111001",
  20388=>"111000000",
  20389=>"111010111",
  20390=>"011110010",
  20391=>"110100001",
  20392=>"000000111",
  20393=>"110010101",
  20394=>"000011101",
  20395=>"010001011",
  20396=>"000101000",
  20397=>"001000011",
  20398=>"001111011",
  20399=>"011101100",
  20400=>"000110001",
  20401=>"101011001",
  20402=>"100100000",
  20403=>"010001111",
  20404=>"001010111",
  20405=>"101000111",
  20406=>"111011111",
  20407=>"000001010",
  20408=>"110001111",
  20409=>"000110111",
  20410=>"000110001",
  20411=>"101010110",
  20412=>"010110111",
  20413=>"001010001",
  20414=>"000000010",
  20415=>"011110100",
  20416=>"010011110",
  20417=>"111111101",
  20418=>"000000001",
  20419=>"001100001",
  20420=>"000110011",
  20421=>"000100010",
  20422=>"011001100",
  20423=>"000000100",
  20424=>"001000001",
  20425=>"010110000",
  20426=>"001000110",
  20427=>"100001100",
  20428=>"001100110",
  20429=>"000000100",
  20430=>"001101000",
  20431=>"000111001",
  20432=>"101100111",
  20433=>"110110001",
  20434=>"101100011",
  20435=>"101110110",
  20436=>"101010111",
  20437=>"110000001",
  20438=>"101111000",
  20439=>"010100111",
  20440=>"100100000",
  20441=>"101001111",
  20442=>"101111010",
  20443=>"011010100",
  20444=>"001000100",
  20445=>"001111110",
  20446=>"011000010",
  20447=>"101100110",
  20448=>"100001101",
  20449=>"101011100",
  20450=>"000001110",
  20451=>"111010111",
  20452=>"110000001",
  20453=>"100100001",
  20454=>"001100001",
  20455=>"111100111",
  20456=>"110110101",
  20457=>"001000110",
  20458=>"100100111",
  20459=>"100100000",
  20460=>"111100110",
  20461=>"001001110",
  20462=>"100001001",
  20463=>"001101100",
  20464=>"100011011",
  20465=>"110011100",
  20466=>"000010011",
  20467=>"111111111",
  20468=>"110010101",
  20469=>"010100100",
  20470=>"000001100",
  20471=>"000000011",
  20472=>"101010011",
  20473=>"100010011",
  20474=>"111100101",
  20475=>"110001110",
  20476=>"000001011",
  20477=>"000001001",
  20478=>"001001101",
  20479=>"101011110",
  20480=>"111100011",
  20481=>"101110110",
  20482=>"001001100",
  20483=>"100100001",
  20484=>"001011010",
  20485=>"000110010",
  20486=>"011101110",
  20487=>"000101010",
  20488=>"100011101",
  20489=>"111110010",
  20490=>"010010111",
  20491=>"011011101",
  20492=>"010101011",
  20493=>"000101011",
  20494=>"000001110",
  20495=>"001010000",
  20496=>"001111000",
  20497=>"011100101",
  20498=>"110010100",
  20499=>"100101100",
  20500=>"001000001",
  20501=>"001111111",
  20502=>"011000100",
  20503=>"010101010",
  20504=>"000110000",
  20505=>"001011100",
  20506=>"100000001",
  20507=>"111111011",
  20508=>"101100001",
  20509=>"000000001",
  20510=>"111101011",
  20511=>"011101110",
  20512=>"101101011",
  20513=>"000001110",
  20514=>"111111010",
  20515=>"101110011",
  20516=>"010111111",
  20517=>"110000001",
  20518=>"100110110",
  20519=>"101101101",
  20520=>"000110010",
  20521=>"011011100",
  20522=>"010010010",
  20523=>"110010110",
  20524=>"001000101",
  20525=>"001101010",
  20526=>"011111001",
  20527=>"000100101",
  20528=>"111101001",
  20529=>"001111010",
  20530=>"111110111",
  20531=>"101101010",
  20532=>"110101001",
  20533=>"110000011",
  20534=>"110111111",
  20535=>"000000000",
  20536=>"001100110",
  20537=>"001001101",
  20538=>"010011011",
  20539=>"001000001",
  20540=>"000101111",
  20541=>"111000000",
  20542=>"101110000",
  20543=>"001001100",
  20544=>"000110100",
  20545=>"011000001",
  20546=>"000100100",
  20547=>"100111110",
  20548=>"011010000",
  20549=>"011011011",
  20550=>"100111010",
  20551=>"110001010",
  20552=>"111101000",
  20553=>"111100011",
  20554=>"100101000",
  20555=>"110010100",
  20556=>"011011110",
  20557=>"111101101",
  20558=>"100010010",
  20559=>"111011100",
  20560=>"111100010",
  20561=>"111011110",
  20562=>"100001000",
  20563=>"110001111",
  20564=>"001110011",
  20565=>"110001010",
  20566=>"100110010",
  20567=>"110111000",
  20568=>"101001000",
  20569=>"111111111",
  20570=>"000100110",
  20571=>"011101001",
  20572=>"011000001",
  20573=>"000001010",
  20574=>"010001110",
  20575=>"100000010",
  20576=>"000000010",
  20577=>"101011101",
  20578=>"010001010",
  20579=>"101110101",
  20580=>"110111100",
  20581=>"010010001",
  20582=>"010101010",
  20583=>"000110010",
  20584=>"110011111",
  20585=>"110111001",
  20586=>"101101001",
  20587=>"000101101",
  20588=>"111000101",
  20589=>"101000101",
  20590=>"111000010",
  20591=>"001000101",
  20592=>"111000101",
  20593=>"011010111",
  20594=>"101010111",
  20595=>"101010110",
  20596=>"010100101",
  20597=>"111111010",
  20598=>"111001111",
  20599=>"010111110",
  20600=>"010110001",
  20601=>"111110001",
  20602=>"010101111",
  20603=>"111111011",
  20604=>"010001001",
  20605=>"000010100",
  20606=>"100001101",
  20607=>"001111111",
  20608=>"010011100",
  20609=>"011110101",
  20610=>"101001100",
  20611=>"100110111",
  20612=>"101101011",
  20613=>"111011100",
  20614=>"111111011",
  20615=>"000110111",
  20616=>"111111111",
  20617=>"011100001",
  20618=>"010111110",
  20619=>"001011110",
  20620=>"000011000",
  20621=>"111110101",
  20622=>"100100110",
  20623=>"010111110",
  20624=>"110000101",
  20625=>"100011110",
  20626=>"111010011",
  20627=>"101000100",
  20628=>"100101010",
  20629=>"011101000",
  20630=>"110111110",
  20631=>"001001110",
  20632=>"011001001",
  20633=>"110001111",
  20634=>"000001011",
  20635=>"011011011",
  20636=>"111110000",
  20637=>"011011100",
  20638=>"000010011",
  20639=>"011111010",
  20640=>"100110100",
  20641=>"101111101",
  20642=>"010100010",
  20643=>"001000100",
  20644=>"111101000",
  20645=>"010110011",
  20646=>"000001010",
  20647=>"000100001",
  20648=>"001000000",
  20649=>"110001110",
  20650=>"010111010",
  20651=>"110000111",
  20652=>"000111011",
  20653=>"100111111",
  20654=>"110000010",
  20655=>"000110100",
  20656=>"001000000",
  20657=>"000111110",
  20658=>"100001000",
  20659=>"001010011",
  20660=>"101001001",
  20661=>"010010110",
  20662=>"000000110",
  20663=>"001111000",
  20664=>"010010100",
  20665=>"010000111",
  20666=>"001011011",
  20667=>"000011000",
  20668=>"001111101",
  20669=>"000111111",
  20670=>"010110111",
  20671=>"111001011",
  20672=>"011111110",
  20673=>"011111110",
  20674=>"000001111",
  20675=>"101000110",
  20676=>"110100011",
  20677=>"111100001",
  20678=>"111101101",
  20679=>"011101011",
  20680=>"011111101",
  20681=>"111101100",
  20682=>"111010000",
  20683=>"110111011",
  20684=>"101000011",
  20685=>"001001010",
  20686=>"101110010",
  20687=>"000101111",
  20688=>"110011000",
  20689=>"101001001",
  20690=>"100011010",
  20691=>"110000101",
  20692=>"110101111",
  20693=>"010010111",
  20694=>"011110101",
  20695=>"011110001",
  20696=>"100110000",
  20697=>"011001100",
  20698=>"000100101",
  20699=>"011111110",
  20700=>"000010000",
  20701=>"101001111",
  20702=>"000001100",
  20703=>"011110000",
  20704=>"000100100",
  20705=>"001101100",
  20706=>"110111000",
  20707=>"111101111",
  20708=>"110010000",
  20709=>"111100001",
  20710=>"100000110",
  20711=>"010011111",
  20712=>"110011110",
  20713=>"110011101",
  20714=>"101000010",
  20715=>"001101011",
  20716=>"101101010",
  20717=>"100100101",
  20718=>"010011010",
  20719=>"011010110",
  20720=>"011110011",
  20721=>"000111000",
  20722=>"010010100",
  20723=>"101011111",
  20724=>"010101001",
  20725=>"111000110",
  20726=>"010010110",
  20727=>"111010111",
  20728=>"010110111",
  20729=>"000000101",
  20730=>"100100110",
  20731=>"000000001",
  20732=>"000010100",
  20733=>"110110001",
  20734=>"100100110",
  20735=>"110111111",
  20736=>"011111100",
  20737=>"011000010",
  20738=>"001101010",
  20739=>"010110111",
  20740=>"010111111",
  20741=>"101010010",
  20742=>"100000101",
  20743=>"101100100",
  20744=>"010010011",
  20745=>"001101110",
  20746=>"101101110",
  20747=>"110001010",
  20748=>"010000010",
  20749=>"111111001",
  20750=>"101101000",
  20751=>"111100111",
  20752=>"000000011",
  20753=>"100101001",
  20754=>"001000011",
  20755=>"111000100",
  20756=>"010110111",
  20757=>"010101011",
  20758=>"001011101",
  20759=>"100001000",
  20760=>"111111111",
  20761=>"010100100",
  20762=>"100110100",
  20763=>"110001000",
  20764=>"001101101",
  20765=>"000010001",
  20766=>"000101001",
  20767=>"101000010",
  20768=>"110110110",
  20769=>"001110100",
  20770=>"000001010",
  20771=>"011001011",
  20772=>"110011110",
  20773=>"010000011",
  20774=>"100110101",
  20775=>"111100010",
  20776=>"101100000",
  20777=>"110111010",
  20778=>"010001100",
  20779=>"001000101",
  20780=>"000100010",
  20781=>"101011111",
  20782=>"000111011",
  20783=>"110111011",
  20784=>"111001010",
  20785=>"101010101",
  20786=>"111010011",
  20787=>"000110111",
  20788=>"010110100",
  20789=>"110100110",
  20790=>"111011111",
  20791=>"001101101",
  20792=>"010010111",
  20793=>"010010001",
  20794=>"001110101",
  20795=>"011000001",
  20796=>"000000000",
  20797=>"011011100",
  20798=>"010100110",
  20799=>"011101000",
  20800=>"000010011",
  20801=>"111111111",
  20802=>"011000000",
  20803=>"111000111",
  20804=>"111011000",
  20805=>"000101010",
  20806=>"110010110",
  20807=>"101110000",
  20808=>"111001100",
  20809=>"011000000",
  20810=>"001100010",
  20811=>"100101110",
  20812=>"000010011",
  20813=>"110101011",
  20814=>"001101110",
  20815=>"101101011",
  20816=>"110011101",
  20817=>"011000110",
  20818=>"100110010",
  20819=>"011101010",
  20820=>"010111101",
  20821=>"110001001",
  20822=>"000011110",
  20823=>"111110110",
  20824=>"000000111",
  20825=>"001000100",
  20826=>"011001010",
  20827=>"110001100",
  20828=>"111110111",
  20829=>"110001101",
  20830=>"011100110",
  20831=>"000000001",
  20832=>"111110111",
  20833=>"110110001",
  20834=>"000011000",
  20835=>"100010100",
  20836=>"000000110",
  20837=>"001000101",
  20838=>"000000100",
  20839=>"011110111",
  20840=>"001000000",
  20841=>"011000111",
  20842=>"000001011",
  20843=>"111101111",
  20844=>"111001110",
  20845=>"111111010",
  20846=>"110000010",
  20847=>"101001100",
  20848=>"001101000",
  20849=>"001001110",
  20850=>"101010000",
  20851=>"011011001",
  20852=>"000111110",
  20853=>"101101101",
  20854=>"111001100",
  20855=>"110000100",
  20856=>"001011010",
  20857=>"000100111",
  20858=>"000100010",
  20859=>"000001110",
  20860=>"110110011",
  20861=>"010101001",
  20862=>"010100001",
  20863=>"100000010",
  20864=>"100011001",
  20865=>"010100010",
  20866=>"101101111",
  20867=>"011000111",
  20868=>"000010010",
  20869=>"111111011",
  20870=>"110111101",
  20871=>"010001000",
  20872=>"010100000",
  20873=>"000101101",
  20874=>"101011101",
  20875=>"001100001",
  20876=>"011110010",
  20877=>"000111101",
  20878=>"111111011",
  20879=>"111110011",
  20880=>"011110110",
  20881=>"110000111",
  20882=>"000100011",
  20883=>"010010000",
  20884=>"001101011",
  20885=>"001001101",
  20886=>"111100000",
  20887=>"111101011",
  20888=>"011101110",
  20889=>"000001011",
  20890=>"100111101",
  20891=>"000000010",
  20892=>"110011011",
  20893=>"100000000",
  20894=>"011000111",
  20895=>"001110100",
  20896=>"000100010",
  20897=>"111100001",
  20898=>"101101011",
  20899=>"111010011",
  20900=>"100011111",
  20901=>"100000111",
  20902=>"000010000",
  20903=>"001010101",
  20904=>"001001011",
  20905=>"100000100",
  20906=>"100101111",
  20907=>"111001010",
  20908=>"001100000",
  20909=>"111000100",
  20910=>"111000011",
  20911=>"100001011",
  20912=>"001001100",
  20913=>"100001100",
  20914=>"100000010",
  20915=>"000111011",
  20916=>"100101001",
  20917=>"010011100",
  20918=>"010110001",
  20919=>"110011111",
  20920=>"110100111",
  20921=>"101010010",
  20922=>"101000100",
  20923=>"110110100",
  20924=>"101100000",
  20925=>"111100111",
  20926=>"011001100",
  20927=>"111100110",
  20928=>"110110111",
  20929=>"000000001",
  20930=>"111011111",
  20931=>"101111110",
  20932=>"101011101",
  20933=>"000110101",
  20934=>"011010110",
  20935=>"000010010",
  20936=>"010011011",
  20937=>"101111010",
  20938=>"110100111",
  20939=>"001101100",
  20940=>"011010011",
  20941=>"111000000",
  20942=>"111110011",
  20943=>"111011111",
  20944=>"010011110",
  20945=>"100000101",
  20946=>"101001000",
  20947=>"000000001",
  20948=>"000010110",
  20949=>"110111001",
  20950=>"111011010",
  20951=>"000101001",
  20952=>"011010100",
  20953=>"000101101",
  20954=>"100100001",
  20955=>"000101010",
  20956=>"111111011",
  20957=>"101011010",
  20958=>"100000001",
  20959=>"111000101",
  20960=>"000110110",
  20961=>"100101010",
  20962=>"110001110",
  20963=>"110110110",
  20964=>"110101110",
  20965=>"000010101",
  20966=>"000110100",
  20967=>"011010110",
  20968=>"101111011",
  20969=>"111101001",
  20970=>"010000000",
  20971=>"101010111",
  20972=>"111010001",
  20973=>"001000000",
  20974=>"010000001",
  20975=>"010110111",
  20976=>"110001101",
  20977=>"000011000",
  20978=>"001010101",
  20979=>"111100010",
  20980=>"010001100",
  20981=>"100111001",
  20982=>"100001001",
  20983=>"010101001",
  20984=>"100010010",
  20985=>"011101011",
  20986=>"011000001",
  20987=>"010010010",
  20988=>"101101101",
  20989=>"100110101",
  20990=>"010000001",
  20991=>"101011111",
  20992=>"010000011",
  20993=>"101001101",
  20994=>"110110110",
  20995=>"000011010",
  20996=>"101110100",
  20997=>"011010000",
  20998=>"101000010",
  20999=>"010111000",
  21000=>"110100101",
  21001=>"000000001",
  21002=>"011101010",
  21003=>"110000010",
  21004=>"100111100",
  21005=>"000000100",
  21006=>"011100001",
  21007=>"111100011",
  21008=>"011011010",
  21009=>"110101111",
  21010=>"101100001",
  21011=>"000100110",
  21012=>"000111001",
  21013=>"101011000",
  21014=>"100111110",
  21015=>"000010010",
  21016=>"111101111",
  21017=>"110101000",
  21018=>"010010100",
  21019=>"100101010",
  21020=>"011101110",
  21021=>"100011011",
  21022=>"100010010",
  21023=>"100100010",
  21024=>"011010010",
  21025=>"000110010",
  21026=>"100010110",
  21027=>"100100101",
  21028=>"101011001",
  21029=>"111101111",
  21030=>"000011110",
  21031=>"110110011",
  21032=>"100011110",
  21033=>"111010110",
  21034=>"001011100",
  21035=>"000000110",
  21036=>"111100011",
  21037=>"001110001",
  21038=>"010001000",
  21039=>"111101000",
  21040=>"111000111",
  21041=>"001011011",
  21042=>"000011010",
  21043=>"110011110",
  21044=>"010111100",
  21045=>"111110101",
  21046=>"000001101",
  21047=>"101100100",
  21048=>"000000010",
  21049=>"000011000",
  21050=>"010101101",
  21051=>"011011101",
  21052=>"100001000",
  21053=>"111111011",
  21054=>"101101010",
  21055=>"110010011",
  21056=>"100101011",
  21057=>"100101100",
  21058=>"000101011",
  21059=>"111111111",
  21060=>"011001000",
  21061=>"010010001",
  21062=>"000010100",
  21063=>"000110011",
  21064=>"001000010",
  21065=>"111000010",
  21066=>"001011100",
  21067=>"110110010",
  21068=>"101111100",
  21069=>"001000111",
  21070=>"000001001",
  21071=>"100111111",
  21072=>"101000111",
  21073=>"001000101",
  21074=>"001010111",
  21075=>"001001000",
  21076=>"001010110",
  21077=>"100110011",
  21078=>"011010111",
  21079=>"111100111",
  21080=>"111101001",
  21081=>"011010110",
  21082=>"011001000",
  21083=>"011000101",
  21084=>"101000001",
  21085=>"001100101",
  21086=>"000101111",
  21087=>"110111000",
  21088=>"001000100",
  21089=>"011001001",
  21090=>"001100111",
  21091=>"000000010",
  21092=>"010100100",
  21093=>"011000101",
  21094=>"011001010",
  21095=>"001001101",
  21096=>"000000101",
  21097=>"001101010",
  21098=>"011000001",
  21099=>"111011000",
  21100=>"000111110",
  21101=>"001100110",
  21102=>"111001110",
  21103=>"100110001",
  21104=>"101001000",
  21105=>"011100011",
  21106=>"100000001",
  21107=>"010001000",
  21108=>"111000100",
  21109=>"011100010",
  21110=>"000011100",
  21111=>"101100001",
  21112=>"111110011",
  21113=>"010110100",
  21114=>"100100000",
  21115=>"001010000",
  21116=>"001000010",
  21117=>"111000001",
  21118=>"111010001",
  21119=>"110110110",
  21120=>"000100100",
  21121=>"111110101",
  21122=>"100111011",
  21123=>"001010110",
  21124=>"101001110",
  21125=>"100100000",
  21126=>"101100010",
  21127=>"011110011",
  21128=>"101100011",
  21129=>"110011000",
  21130=>"110101101",
  21131=>"010101011",
  21132=>"101000100",
  21133=>"111111011",
  21134=>"101101000",
  21135=>"111100000",
  21136=>"100111111",
  21137=>"100010011",
  21138=>"000001010",
  21139=>"011011111",
  21140=>"010100100",
  21141=>"010011101",
  21142=>"010010101",
  21143=>"110010001",
  21144=>"000011101",
  21145=>"001100000",
  21146=>"100111111",
  21147=>"010010000",
  21148=>"110001001",
  21149=>"101101011",
  21150=>"111010011",
  21151=>"100110000",
  21152=>"101000100",
  21153=>"101000001",
  21154=>"010010010",
  21155=>"110101000",
  21156=>"100100100",
  21157=>"001101000",
  21158=>"011100101",
  21159=>"001100000",
  21160=>"101100000",
  21161=>"011000010",
  21162=>"000100100",
  21163=>"111101100",
  21164=>"111000110",
  21165=>"011101000",
  21166=>"111010110",
  21167=>"000100000",
  21168=>"011011011",
  21169=>"101010101",
  21170=>"111011001",
  21171=>"011111011",
  21172=>"010011010",
  21173=>"001000100",
  21174=>"110101101",
  21175=>"000011111",
  21176=>"100011110",
  21177=>"011011100",
  21178=>"010001010",
  21179=>"001110101",
  21180=>"110000101",
  21181=>"010100110",
  21182=>"101100110",
  21183=>"110000110",
  21184=>"000000011",
  21185=>"111111101",
  21186=>"001100111",
  21187=>"001001100",
  21188=>"010001111",
  21189=>"011000110",
  21190=>"100010101",
  21191=>"110101001",
  21192=>"011111111",
  21193=>"000011101",
  21194=>"001000000",
  21195=>"101001010",
  21196=>"100001111",
  21197=>"011110000",
  21198=>"100011111",
  21199=>"010111010",
  21200=>"101001001",
  21201=>"000101000",
  21202=>"101111010",
  21203=>"110111110",
  21204=>"100111111",
  21205=>"001100111",
  21206=>"010110001",
  21207=>"010000000",
  21208=>"010000010",
  21209=>"111101110",
  21210=>"111111101",
  21211=>"000101000",
  21212=>"001101101",
  21213=>"011111001",
  21214=>"110100100",
  21215=>"110110111",
  21216=>"001010010",
  21217=>"110010001",
  21218=>"000111111",
  21219=>"100011000",
  21220=>"110010001",
  21221=>"010011001",
  21222=>"010110100",
  21223=>"100011011",
  21224=>"000000110",
  21225=>"011101110",
  21226=>"010101000",
  21227=>"010011001",
  21228=>"010110111",
  21229=>"100011010",
  21230=>"100001000",
  21231=>"101000011",
  21232=>"100100100",
  21233=>"101101010",
  21234=>"100000010",
  21235=>"000011111",
  21236=>"010111010",
  21237=>"011010000",
  21238=>"010011000",
  21239=>"111100111",
  21240=>"110000011",
  21241=>"111100100",
  21242=>"010110110",
  21243=>"001001001",
  21244=>"110010000",
  21245=>"001001110",
  21246=>"111010111",
  21247=>"110111111",
  21248=>"000100110",
  21249=>"000000111",
  21250=>"101010000",
  21251=>"111111111",
  21252=>"101000000",
  21253=>"011000010",
  21254=>"001111100",
  21255=>"001101100",
  21256=>"000100101",
  21257=>"011011111",
  21258=>"011000010",
  21259=>"000000100",
  21260=>"011011111",
  21261=>"111101111",
  21262=>"111110010",
  21263=>"110010110",
  21264=>"000000010",
  21265=>"001100000",
  21266=>"110100001",
  21267=>"001000000",
  21268=>"110101001",
  21269=>"111010111",
  21270=>"111111000",
  21271=>"000001010",
  21272=>"001110101",
  21273=>"010001011",
  21274=>"000110010",
  21275=>"101000100",
  21276=>"010110000",
  21277=>"110001100",
  21278=>"100100101",
  21279=>"111011011",
  21280=>"010111000",
  21281=>"110111011",
  21282=>"000100111",
  21283=>"011101110",
  21284=>"111111000",
  21285=>"011011110",
  21286=>"001010011",
  21287=>"100000101",
  21288=>"111111111",
  21289=>"111011101",
  21290=>"100111001",
  21291=>"101111011",
  21292=>"000111010",
  21293=>"010000100",
  21294=>"011001000",
  21295=>"111010111",
  21296=>"010100000",
  21297=>"100011111",
  21298=>"001001111",
  21299=>"100000110",
  21300=>"000000110",
  21301=>"110001101",
  21302=>"000001011",
  21303=>"001101111",
  21304=>"010001110",
  21305=>"000010110",
  21306=>"001000111",
  21307=>"101000111",
  21308=>"110110000",
  21309=>"111010001",
  21310=>"111010101",
  21311=>"001010110",
  21312=>"100111101",
  21313=>"100111011",
  21314=>"011000001",
  21315=>"011001111",
  21316=>"011001000",
  21317=>"000001011",
  21318=>"000001111",
  21319=>"001011001",
  21320=>"011101100",
  21321=>"100110110",
  21322=>"110000110",
  21323=>"010111111",
  21324=>"000101110",
  21325=>"010101000",
  21326=>"001010110",
  21327=>"000010001",
  21328=>"111010111",
  21329=>"010001010",
  21330=>"101000011",
  21331=>"110111111",
  21332=>"000111110",
  21333=>"011010011",
  21334=>"010000110",
  21335=>"011010001",
  21336=>"000000011",
  21337=>"011000110",
  21338=>"101111110",
  21339=>"111011100",
  21340=>"001011111",
  21341=>"000000000",
  21342=>"100000101",
  21343=>"000110110",
  21344=>"010011101",
  21345=>"000000011",
  21346=>"000000111",
  21347=>"101001001",
  21348=>"111110001",
  21349=>"100011101",
  21350=>"100100111",
  21351=>"100000000",
  21352=>"110000000",
  21353=>"100100010",
  21354=>"011001000",
  21355=>"110101101",
  21356=>"110101101",
  21357=>"000010110",
  21358=>"101000100",
  21359=>"100110001",
  21360=>"101000111",
  21361=>"110111010",
  21362=>"110000001",
  21363=>"100011010",
  21364=>"101011000",
  21365=>"010010010",
  21366=>"101011100",
  21367=>"010011010",
  21368=>"101011100",
  21369=>"111000100",
  21370=>"010001001",
  21371=>"100101001",
  21372=>"101010000",
  21373=>"011011101",
  21374=>"010100001",
  21375=>"111101111",
  21376=>"101010011",
  21377=>"100011001",
  21378=>"110010011",
  21379=>"100011110",
  21380=>"010001001",
  21381=>"111111101",
  21382=>"000011000",
  21383=>"110001100",
  21384=>"000111110",
  21385=>"001110011",
  21386=>"000100100",
  21387=>"000110010",
  21388=>"101010010",
  21389=>"010000011",
  21390=>"001010101",
  21391=>"110101111",
  21392=>"010100100",
  21393=>"011110100",
  21394=>"000000101",
  21395=>"000110000",
  21396=>"001100011",
  21397=>"101100111",
  21398=>"101010111",
  21399=>"111111100",
  21400=>"111110110",
  21401=>"001100111",
  21402=>"110001011",
  21403=>"010011001",
  21404=>"010100101",
  21405=>"010111001",
  21406=>"111010000",
  21407=>"011101011",
  21408=>"010010001",
  21409=>"010011101",
  21410=>"010001001",
  21411=>"101110110",
  21412=>"100101011",
  21413=>"101110011",
  21414=>"111110011",
  21415=>"011011000",
  21416=>"111001001",
  21417=>"000000000",
  21418=>"111111001",
  21419=>"011010111",
  21420=>"010101010",
  21421=>"100011101",
  21422=>"111011100",
  21423=>"011001100",
  21424=>"011110100",
  21425=>"100010100",
  21426=>"100101111",
  21427=>"010001010",
  21428=>"010001111",
  21429=>"111001000",
  21430=>"110100001",
  21431=>"111100011",
  21432=>"100000000",
  21433=>"011001001",
  21434=>"100010110",
  21435=>"010011001",
  21436=>"010111111",
  21437=>"111010100",
  21438=>"111101111",
  21439=>"010111000",
  21440=>"111101111",
  21441=>"100100010",
  21442=>"000001101",
  21443=>"110101100",
  21444=>"000111001",
  21445=>"101100011",
  21446=>"101110010",
  21447=>"011110111",
  21448=>"010000000",
  21449=>"111010011",
  21450=>"001101101",
  21451=>"111101100",
  21452=>"011000000",
  21453=>"110001010",
  21454=>"110100010",
  21455=>"011011100",
  21456=>"111101111",
  21457=>"001010101",
  21458=>"101100100",
  21459=>"000101010",
  21460=>"011011100",
  21461=>"011101111",
  21462=>"110101001",
  21463=>"011000000",
  21464=>"101100001",
  21465=>"000111010",
  21466=>"100000110",
  21467=>"011001010",
  21468=>"100000100",
  21469=>"111101011",
  21470=>"001110011",
  21471=>"100001110",
  21472=>"001110010",
  21473=>"101110001",
  21474=>"111001101",
  21475=>"110101011",
  21476=>"011111100",
  21477=>"111110011",
  21478=>"111111011",
  21479=>"011101000",
  21480=>"000011100",
  21481=>"000110111",
  21482=>"010010011",
  21483=>"001110111",
  21484=>"001010111",
  21485=>"101011100",
  21486=>"100010001",
  21487=>"010001000",
  21488=>"011000111",
  21489=>"001110101",
  21490=>"101111111",
  21491=>"111011010",
  21492=>"011010100",
  21493=>"010010101",
  21494=>"000111111",
  21495=>"111111111",
  21496=>"110101001",
  21497=>"101111111",
  21498=>"100110111",
  21499=>"101011110",
  21500=>"111011000",
  21501=>"000101110",
  21502=>"111111101",
  21503=>"110010110",
  21504=>"101001010",
  21505=>"111011110",
  21506=>"110100111",
  21507=>"011001101",
  21508=>"011000010",
  21509=>"101100011",
  21510=>"010111001",
  21511=>"111101011",
  21512=>"010100001",
  21513=>"000000000",
  21514=>"100000000",
  21515=>"111100111",
  21516=>"010100001",
  21517=>"110000111",
  21518=>"000101011",
  21519=>"110110110",
  21520=>"000000001",
  21521=>"101011000",
  21522=>"011100010",
  21523=>"011000000",
  21524=>"010001101",
  21525=>"000111010",
  21526=>"100001110",
  21527=>"100000001",
  21528=>"001010100",
  21529=>"110110111",
  21530=>"110101010",
  21531=>"001011010",
  21532=>"101110101",
  21533=>"000011101",
  21534=>"000110001",
  21535=>"101001101",
  21536=>"100100111",
  21537=>"000011110",
  21538=>"001001101",
  21539=>"111000010",
  21540=>"101010010",
  21541=>"111010110",
  21542=>"011000011",
  21543=>"001011001",
  21544=>"011001101",
  21545=>"110001110",
  21546=>"000010100",
  21547=>"001000110",
  21548=>"010000010",
  21549=>"110111110",
  21550=>"000110000",
  21551=>"111100001",
  21552=>"001011011",
  21553=>"100110000",
  21554=>"001111000",
  21555=>"101100001",
  21556=>"000100010",
  21557=>"011111100",
  21558=>"000000000",
  21559=>"110100101",
  21560=>"000001110",
  21561=>"110111001",
  21562=>"110110101",
  21563=>"010001001",
  21564=>"101110111",
  21565=>"010001110",
  21566=>"100100010",
  21567=>"101100010",
  21568=>"011111111",
  21569=>"100000011",
  21570=>"000100011",
  21571=>"111111110",
  21572=>"011100111",
  21573=>"000110001",
  21574=>"101110011",
  21575=>"100100011",
  21576=>"110000111",
  21577=>"000100010",
  21578=>"111111010",
  21579=>"000001111",
  21580=>"001011111",
  21581=>"110000100",
  21582=>"100111111",
  21583=>"111110001",
  21584=>"110110011",
  21585=>"101001001",
  21586=>"101110010",
  21587=>"010011110",
  21588=>"111110111",
  21589=>"001010100",
  21590=>"011000010",
  21591=>"001001010",
  21592=>"101011011",
  21593=>"010010100",
  21594=>"011110000",
  21595=>"101100101",
  21596=>"101001111",
  21597=>"110110101",
  21598=>"000001011",
  21599=>"110010011",
  21600=>"010111001",
  21601=>"111110100",
  21602=>"010001010",
  21603=>"100001010",
  21604=>"001110100",
  21605=>"101000111",
  21606=>"000101111",
  21607=>"101000001",
  21608=>"010010001",
  21609=>"010011110",
  21610=>"111100010",
  21611=>"011001010",
  21612=>"010000001",
  21613=>"001010001",
  21614=>"000110110",
  21615=>"010101011",
  21616=>"000000100",
  21617=>"000110001",
  21618=>"101101001",
  21619=>"100001101",
  21620=>"000001000",
  21621=>"101111010",
  21622=>"010101011",
  21623=>"110011100",
  21624=>"010100001",
  21625=>"010110011",
  21626=>"001010100",
  21627=>"101100111",
  21628=>"101111101",
  21629=>"100110011",
  21630=>"100010001",
  21631=>"011010011",
  21632=>"100001010",
  21633=>"000000000",
  21634=>"001100110",
  21635=>"011010110",
  21636=>"111101000",
  21637=>"010111011",
  21638=>"110100111",
  21639=>"011010011",
  21640=>"011000110",
  21641=>"010011110",
  21642=>"111010110",
  21643=>"101001101",
  21644=>"001101010",
  21645=>"011000001",
  21646=>"101001110",
  21647=>"101001010",
  21648=>"111110001",
  21649=>"111111110",
  21650=>"000100010",
  21651=>"110101000",
  21652=>"111001000",
  21653=>"011001011",
  21654=>"001010110",
  21655=>"100111100",
  21656=>"100100100",
  21657=>"010010110",
  21658=>"000000110",
  21659=>"000101000",
  21660=>"011100000",
  21661=>"100010100",
  21662=>"000000011",
  21663=>"101111010",
  21664=>"011111001",
  21665=>"011010110",
  21666=>"110010010",
  21667=>"011011101",
  21668=>"001110001",
  21669=>"011000110",
  21670=>"001101001",
  21671=>"011100011",
  21672=>"101100011",
  21673=>"111111100",
  21674=>"000110000",
  21675=>"110100000",
  21676=>"100100000",
  21677=>"110011010",
  21678=>"100000010",
  21679=>"101001110",
  21680=>"100101101",
  21681=>"000101101",
  21682=>"100001111",
  21683=>"101111111",
  21684=>"111110001",
  21685=>"101010001",
  21686=>"101110111",
  21687=>"011000000",
  21688=>"101111001",
  21689=>"100000000",
  21690=>"011001000",
  21691=>"010110100",
  21692=>"110101110",
  21693=>"010001001",
  21694=>"010000001",
  21695=>"010101101",
  21696=>"110100110",
  21697=>"101000100",
  21698=>"111100111",
  21699=>"111011001",
  21700=>"100110000",
  21701=>"110010010",
  21702=>"111001100",
  21703=>"010101100",
  21704=>"011010111",
  21705=>"101010010",
  21706=>"101011000",
  21707=>"001100111",
  21708=>"100100001",
  21709=>"111011011",
  21710=>"101100010",
  21711=>"001100000",
  21712=>"001001100",
  21713=>"100000001",
  21714=>"000011011",
  21715=>"011010001",
  21716=>"011100111",
  21717=>"101110111",
  21718=>"011010010",
  21719=>"110010010",
  21720=>"101000111",
  21721=>"011011101",
  21722=>"100011001",
  21723=>"110110110",
  21724=>"010001101",
  21725=>"111010010",
  21726=>"000101000",
  21727=>"110001101",
  21728=>"000011001",
  21729=>"000110110",
  21730=>"001001101",
  21731=>"001010000",
  21732=>"100000110",
  21733=>"000011101",
  21734=>"010111101",
  21735=>"001001010",
  21736=>"100111001",
  21737=>"010001011",
  21738=>"111111010",
  21739=>"001010010",
  21740=>"000100100",
  21741=>"000001111",
  21742=>"101101101",
  21743=>"011011101",
  21744=>"100110011",
  21745=>"110100001",
  21746=>"100011000",
  21747=>"111100101",
  21748=>"011111100",
  21749=>"000101111",
  21750=>"100110101",
  21751=>"100000000",
  21752=>"010010011",
  21753=>"011011000",
  21754=>"001110001",
  21755=>"110111011",
  21756=>"101011110",
  21757=>"011111111",
  21758=>"111000010",
  21759=>"011000111",
  21760=>"100110000",
  21761=>"101000100",
  21762=>"010010011",
  21763=>"010100111",
  21764=>"001110010",
  21765=>"011010110",
  21766=>"110001010",
  21767=>"110010000",
  21768=>"010101001",
  21769=>"010000010",
  21770=>"100111001",
  21771=>"000100101",
  21772=>"111010000",
  21773=>"010001000",
  21774=>"000111010",
  21775=>"100000000",
  21776=>"111111111",
  21777=>"001000001",
  21778=>"110110111",
  21779=>"011000110",
  21780=>"010100111",
  21781=>"110101010",
  21782=>"010111100",
  21783=>"010000000",
  21784=>"010011010",
  21785=>"000101101",
  21786=>"101001001",
  21787=>"001111101",
  21788=>"000110001",
  21789=>"100000001",
  21790=>"000011001",
  21791=>"001010011",
  21792=>"000010111",
  21793=>"011010101",
  21794=>"000000010",
  21795=>"010000001",
  21796=>"001101101",
  21797=>"101100110",
  21798=>"010010101",
  21799=>"110110111",
  21800=>"000010111",
  21801=>"100010000",
  21802=>"100001011",
  21803=>"000010010",
  21804=>"111010110",
  21805=>"110011011",
  21806=>"110111010",
  21807=>"011100011",
  21808=>"110010010",
  21809=>"100001100",
  21810=>"111111110",
  21811=>"101011011",
  21812=>"100000011",
  21813=>"001000001",
  21814=>"010100100",
  21815=>"010101001",
  21816=>"101000111",
  21817=>"111111000",
  21818=>"100100011",
  21819=>"110101111",
  21820=>"101101110",
  21821=>"011011110",
  21822=>"111101001",
  21823=>"100100010",
  21824=>"000000001",
  21825=>"000010011",
  21826=>"111110001",
  21827=>"111011000",
  21828=>"100000010",
  21829=>"100001111",
  21830=>"001110010",
  21831=>"110001101",
  21832=>"011101101",
  21833=>"111001011",
  21834=>"111110111",
  21835=>"011010000",
  21836=>"101100010",
  21837=>"010001011",
  21838=>"101011000",
  21839=>"101111011",
  21840=>"000100001",
  21841=>"100111001",
  21842=>"001111101",
  21843=>"000100011",
  21844=>"010110011",
  21845=>"110000001",
  21846=>"100101100",
  21847=>"000100100",
  21848=>"001111100",
  21849=>"010100101",
  21850=>"011110010",
  21851=>"011111111",
  21852=>"100111000",
  21853=>"100110111",
  21854=>"011000101",
  21855=>"010001000",
  21856=>"011000011",
  21857=>"000000011",
  21858=>"001001111",
  21859=>"000100100",
  21860=>"111101011",
  21861=>"000110100",
  21862=>"111101100",
  21863=>"110110110",
  21864=>"111001100",
  21865=>"010000000",
  21866=>"011001100",
  21867=>"010001110",
  21868=>"010111000",
  21869=>"101100011",
  21870=>"101001000",
  21871=>"100101010",
  21872=>"000001100",
  21873=>"010101001",
  21874=>"010110111",
  21875=>"011111011",
  21876=>"101000001",
  21877=>"011110000",
  21878=>"011100011",
  21879=>"101100100",
  21880=>"001111110",
  21881=>"010010111",
  21882=>"110101001",
  21883=>"111111110",
  21884=>"101000101",
  21885=>"110010101",
  21886=>"011101101",
  21887=>"011011110",
  21888=>"100100001",
  21889=>"011000111",
  21890=>"000101111",
  21891=>"101101011",
  21892=>"010100101",
  21893=>"010101100",
  21894=>"100000100",
  21895=>"001001111",
  21896=>"110110001",
  21897=>"111010010",
  21898=>"000100101",
  21899=>"000110111",
  21900=>"101001100",
  21901=>"010101001",
  21902=>"100111000",
  21903=>"010101101",
  21904=>"001101100",
  21905=>"000000010",
  21906=>"100000100",
  21907=>"011101100",
  21908=>"110111001",
  21909=>"101001111",
  21910=>"100010110",
  21911=>"110100001",
  21912=>"111000010",
  21913=>"101100011",
  21914=>"011101100",
  21915=>"100111111",
  21916=>"110111110",
  21917=>"110011110",
  21918=>"100100010",
  21919=>"000101110",
  21920=>"110011010",
  21921=>"011101101",
  21922=>"000101101",
  21923=>"011010011",
  21924=>"110101100",
  21925=>"000101000",
  21926=>"100010011",
  21927=>"010000100",
  21928=>"101010001",
  21929=>"101101100",
  21930=>"101100010",
  21931=>"101101100",
  21932=>"111000101",
  21933=>"101000110",
  21934=>"011000111",
  21935=>"000001100",
  21936=>"100110000",
  21937=>"110110110",
  21938=>"010101111",
  21939=>"100110010",
  21940=>"110011011",
  21941=>"001110111",
  21942=>"010000010",
  21943=>"111101100",
  21944=>"111010010",
  21945=>"011000000",
  21946=>"111101011",
  21947=>"001110010",
  21948=>"100111111",
  21949=>"100011101",
  21950=>"011001110",
  21951=>"000110011",
  21952=>"100101000",
  21953=>"101101001",
  21954=>"111001011",
  21955=>"111010010",
  21956=>"111000001",
  21957=>"101100000",
  21958=>"000000110",
  21959=>"111010111",
  21960=>"000111111",
  21961=>"110111111",
  21962=>"010000001",
  21963=>"101100101",
  21964=>"101101101",
  21965=>"100011100",
  21966=>"010010111",
  21967=>"001101010",
  21968=>"010100110",
  21969=>"111000001",
  21970=>"010101011",
  21971=>"111000011",
  21972=>"110100000",
  21973=>"101100101",
  21974=>"110000000",
  21975=>"000000001",
  21976=>"101000111",
  21977=>"111001001",
  21978=>"101011001",
  21979=>"100110010",
  21980=>"111011010",
  21981=>"100101101",
  21982=>"101000101",
  21983=>"111100101",
  21984=>"001100011",
  21985=>"110100001",
  21986=>"111111001",
  21987=>"100111101",
  21988=>"001101101",
  21989=>"110000011",
  21990=>"100000101",
  21991=>"010010001",
  21992=>"001110101",
  21993=>"001110111",
  21994=>"000100111",
  21995=>"011011101",
  21996=>"001101001",
  21997=>"100100000",
  21998=>"101111010",
  21999=>"100111101",
  22000=>"111010000",
  22001=>"110000101",
  22002=>"000100011",
  22003=>"100010000",
  22004=>"110111000",
  22005=>"100011001",
  22006=>"101101001",
  22007=>"110000000",
  22008=>"101001100",
  22009=>"011001110",
  22010=>"010001100",
  22011=>"101000010",
  22012=>"100111110",
  22013=>"011111101",
  22014=>"110010101",
  22015=>"100111010",
  22016=>"100110100",
  22017=>"101111100",
  22018=>"011101001",
  22019=>"101000001",
  22020=>"100010001",
  22021=>"110110111",
  22022=>"110111010",
  22023=>"100100000",
  22024=>"111000110",
  22025=>"100100101",
  22026=>"111101000",
  22027=>"100101001",
  22028=>"110011010",
  22029=>"010100111",
  22030=>"011000100",
  22031=>"110110111",
  22032=>"110111011",
  22033=>"111101110",
  22034=>"110011101",
  22035=>"011000000",
  22036=>"001010000",
  22037=>"000100011",
  22038=>"111001110",
  22039=>"101100110",
  22040=>"000000101",
  22041=>"000000111",
  22042=>"000110011",
  22043=>"101101111",
  22044=>"011001100",
  22045=>"011001001",
  22046=>"100111110",
  22047=>"110101110",
  22048=>"010011110",
  22049=>"101101001",
  22050=>"010000111",
  22051=>"101110110",
  22052=>"111110001",
  22053=>"011110000",
  22054=>"010100011",
  22055=>"101110110",
  22056=>"000000011",
  22057=>"100010000",
  22058=>"110010100",
  22059=>"010010100",
  22060=>"100111110",
  22061=>"100000000",
  22062=>"100000010",
  22063=>"100111011",
  22064=>"101101010",
  22065=>"011101010",
  22066=>"111110011",
  22067=>"101101010",
  22068=>"001010111",
  22069=>"000110111",
  22070=>"101101010",
  22071=>"000100010",
  22072=>"101111011",
  22073=>"010111011",
  22074=>"011000010",
  22075=>"101101011",
  22076=>"111010001",
  22077=>"010010110",
  22078=>"110010010",
  22079=>"101111000",
  22080=>"101000111",
  22081=>"101111011",
  22082=>"011110110",
  22083=>"010101110",
  22084=>"111100101",
  22085=>"001010100",
  22086=>"011001110",
  22087=>"000001010",
  22088=>"001001110",
  22089=>"000010011",
  22090=>"000000011",
  22091=>"011011100",
  22092=>"010011110",
  22093=>"011010110",
  22094=>"001010110",
  22095=>"110010011",
  22096=>"010010001",
  22097=>"000111110",
  22098=>"101011110",
  22099=>"110000001",
  22100=>"010101000",
  22101=>"011110001",
  22102=>"111001110",
  22103=>"111000111",
  22104=>"001011000",
  22105=>"001000101",
  22106=>"111010110",
  22107=>"000001000",
  22108=>"100111111",
  22109=>"110011110",
  22110=>"000101011",
  22111=>"011011110",
  22112=>"110000001",
  22113=>"000100100",
  22114=>"101011111",
  22115=>"101010111",
  22116=>"101000111",
  22117=>"101001100",
  22118=>"101110101",
  22119=>"011010000",
  22120=>"010101011",
  22121=>"101100110",
  22122=>"100100100",
  22123=>"110000000",
  22124=>"111000000",
  22125=>"010111001",
  22126=>"010011110",
  22127=>"010000010",
  22128=>"111100110",
  22129=>"001111100",
  22130=>"111101101",
  22131=>"010100011",
  22132=>"011011010",
  22133=>"111100110",
  22134=>"011010100",
  22135=>"010000110",
  22136=>"111000101",
  22137=>"100000110",
  22138=>"001101010",
  22139=>"011000000",
  22140=>"101001100",
  22141=>"011010011",
  22142=>"100101110",
  22143=>"111010110",
  22144=>"111110010",
  22145=>"100000100",
  22146=>"110101111",
  22147=>"111001100",
  22148=>"010100101",
  22149=>"100010000",
  22150=>"010011110",
  22151=>"010001110",
  22152=>"001101100",
  22153=>"111000110",
  22154=>"111000100",
  22155=>"000100010",
  22156=>"000011110",
  22157=>"000011000",
  22158=>"110010011",
  22159=>"010111100",
  22160=>"001000001",
  22161=>"011001111",
  22162=>"100000111",
  22163=>"100110000",
  22164=>"000010010",
  22165=>"001100110",
  22166=>"100111100",
  22167=>"110101100",
  22168=>"111010000",
  22169=>"000111000",
  22170=>"101101110",
  22171=>"101110110",
  22172=>"010000000",
  22173=>"111001001",
  22174=>"100101101",
  22175=>"110000001",
  22176=>"100010101",
  22177=>"010001100",
  22178=>"010010110",
  22179=>"001001101",
  22180=>"110101101",
  22181=>"110001001",
  22182=>"101100100",
  22183=>"111000001",
  22184=>"001111110",
  22185=>"100010011",
  22186=>"011101010",
  22187=>"000100100",
  22188=>"010000000",
  22189=>"110011001",
  22190=>"101011001",
  22191=>"101111000",
  22192=>"100101000",
  22193=>"110010110",
  22194=>"101000111",
  22195=>"100111011",
  22196=>"110010011",
  22197=>"111101101",
  22198=>"101110100",
  22199=>"111100001",
  22200=>"011010111",
  22201=>"101110101",
  22202=>"100001110",
  22203=>"111000101",
  22204=>"010010000",
  22205=>"111011111",
  22206=>"110110100",
  22207=>"101100011",
  22208=>"100010101",
  22209=>"011110101",
  22210=>"111111010",
  22211=>"110111110",
  22212=>"110010101",
  22213=>"100001001",
  22214=>"000000010",
  22215=>"110011101",
  22216=>"010011110",
  22217=>"110000110",
  22218=>"011010000",
  22219=>"000001011",
  22220=>"000010101",
  22221=>"111101111",
  22222=>"111001100",
  22223=>"110010100",
  22224=>"111111111",
  22225=>"110011110",
  22226=>"111000011",
  22227=>"111001010",
  22228=>"101111100",
  22229=>"010010010",
  22230=>"001001001",
  22231=>"101001001",
  22232=>"101111001",
  22233=>"011011011",
  22234=>"100101001",
  22235=>"011001110",
  22236=>"101000001",
  22237=>"111110000",
  22238=>"110111011",
  22239=>"011010001",
  22240=>"011101100",
  22241=>"101100011",
  22242=>"001101100",
  22243=>"111011010",
  22244=>"000100010",
  22245=>"000000000",
  22246=>"111100001",
  22247=>"011011111",
  22248=>"111001111",
  22249=>"011101101",
  22250=>"110111001",
  22251=>"101101001",
  22252=>"000100111",
  22253=>"110011000",
  22254=>"111101011",
  22255=>"100001001",
  22256=>"101010010",
  22257=>"100000110",
  22258=>"111111111",
  22259=>"001011010",
  22260=>"000110110",
  22261=>"011101011",
  22262=>"111101011",
  22263=>"111111110",
  22264=>"111101111",
  22265=>"011000111",
  22266=>"110110011",
  22267=>"011011010",
  22268=>"101100001",
  22269=>"000000111",
  22270=>"000000001",
  22271=>"010010101",
  22272=>"010001101",
  22273=>"001001001",
  22274=>"111000000",
  22275=>"000011011",
  22276=>"110100001",
  22277=>"010100010",
  22278=>"010101011",
  22279=>"011010000",
  22280=>"111011110",
  22281=>"011111011",
  22282=>"011110100",
  22283=>"101000110",
  22284=>"000001000",
  22285=>"111101001",
  22286=>"111001100",
  22287=>"011000101",
  22288=>"000010001",
  22289=>"111010110",
  22290=>"100100101",
  22291=>"101100100",
  22292=>"000010101",
  22293=>"010110111",
  22294=>"000101111",
  22295=>"011010110",
  22296=>"011100010",
  22297=>"011011111",
  22298=>"001010000",
  22299=>"110110010",
  22300=>"010000000",
  22301=>"110101010",
  22302=>"100010110",
  22303=>"100011000",
  22304=>"100000101",
  22305=>"011100001",
  22306=>"111010011",
  22307=>"010111011",
  22308=>"001000001",
  22309=>"000110001",
  22310=>"110111100",
  22311=>"100110011",
  22312=>"111011011",
  22313=>"000010001",
  22314=>"001110011",
  22315=>"101101011",
  22316=>"011001011",
  22317=>"110010001",
  22318=>"001010010",
  22319=>"110011111",
  22320=>"100010010",
  22321=>"101111011",
  22322=>"000101011",
  22323=>"111111001",
  22324=>"000101110",
  22325=>"101111100",
  22326=>"100111010",
  22327=>"000100000",
  22328=>"100110110",
  22329=>"101100000",
  22330=>"001111011",
  22331=>"000000100",
  22332=>"111000101",
  22333=>"001100100",
  22334=>"000010000",
  22335=>"110100101",
  22336=>"100100001",
  22337=>"100111111",
  22338=>"000111111",
  22339=>"000000111",
  22340=>"100110111",
  22341=>"110101010",
  22342=>"100010000",
  22343=>"110101111",
  22344=>"101100001",
  22345=>"100001011",
  22346=>"101101110",
  22347=>"000010101",
  22348=>"000101111",
  22349=>"111101101",
  22350=>"010001000",
  22351=>"110101011",
  22352=>"110101011",
  22353=>"100010100",
  22354=>"111110001",
  22355=>"100101000",
  22356=>"111110101",
  22357=>"000010111",
  22358=>"110011010",
  22359=>"011010010",
  22360=>"011011111",
  22361=>"110101000",
  22362=>"110010001",
  22363=>"101010101",
  22364=>"111111001",
  22365=>"000100000",
  22366=>"010001111",
  22367=>"001100010",
  22368=>"011101000",
  22369=>"001011100",
  22370=>"000110110",
  22371=>"101101101",
  22372=>"100011000",
  22373=>"110100000",
  22374=>"111100110",
  22375=>"011001111",
  22376=>"101001001",
  22377=>"110100110",
  22378=>"110001100",
  22379=>"111000011",
  22380=>"001111010",
  22381=>"001000110",
  22382=>"111101011",
  22383=>"011111010",
  22384=>"111110000",
  22385=>"011100010",
  22386=>"101110000",
  22387=>"011111111",
  22388=>"110110110",
  22389=>"101111011",
  22390=>"101101111",
  22391=>"000011011",
  22392=>"000100000",
  22393=>"001100100",
  22394=>"010000010",
  22395=>"111100100",
  22396=>"000001001",
  22397=>"011101100",
  22398=>"011011110",
  22399=>"110111000",
  22400=>"111101010",
  22401=>"011011010",
  22402=>"100111111",
  22403=>"110111101",
  22404=>"111110000",
  22405=>"100010000",
  22406=>"001011010",
  22407=>"011000011",
  22408=>"011111100",
  22409=>"011010000",
  22410=>"011101111",
  22411=>"010011011",
  22412=>"100010010",
  22413=>"100100100",
  22414=>"001111111",
  22415=>"111010101",
  22416=>"111110111",
  22417=>"001101111",
  22418=>"100000000",
  22419=>"001001000",
  22420=>"101111100",
  22421=>"110011111",
  22422=>"010000111",
  22423=>"010101000",
  22424=>"010000001",
  22425=>"101101110",
  22426=>"110101010",
  22427=>"010010001",
  22428=>"010001011",
  22429=>"111000010",
  22430=>"011001011",
  22431=>"111010100",
  22432=>"001000111",
  22433=>"110110100",
  22434=>"001100110",
  22435=>"110011010",
  22436=>"000110010",
  22437=>"010111010",
  22438=>"101100011",
  22439=>"011001101",
  22440=>"000000000",
  22441=>"101100111",
  22442=>"100101111",
  22443=>"101001110",
  22444=>"110011000",
  22445=>"010010010",
  22446=>"110011101",
  22447=>"101010101",
  22448=>"000000110",
  22449=>"101010000",
  22450=>"001001101",
  22451=>"111101010",
  22452=>"001011011",
  22453=>"111010110",
  22454=>"111100000",
  22455=>"001001111",
  22456=>"100000100",
  22457=>"010001101",
  22458=>"100111110",
  22459=>"111100100",
  22460=>"010000010",
  22461=>"100111110",
  22462=>"100101111",
  22463=>"111011111",
  22464=>"110110000",
  22465=>"100010100",
  22466=>"110010111",
  22467=>"101110001",
  22468=>"010110100",
  22469=>"011100101",
  22470=>"001011110",
  22471=>"010100011",
  22472=>"110001110",
  22473=>"010000110",
  22474=>"000000100",
  22475=>"110100010",
  22476=>"011001001",
  22477=>"000000000",
  22478=>"111110001",
  22479=>"010011010",
  22480=>"011100011",
  22481=>"010000101",
  22482=>"101010111",
  22483=>"000000001",
  22484=>"010010010",
  22485=>"100101000",
  22486=>"010101111",
  22487=>"110111010",
  22488=>"100000110",
  22489=>"010111011",
  22490=>"101100100",
  22491=>"110001001",
  22492=>"100010100",
  22493=>"101010011",
  22494=>"011100100",
  22495=>"111110101",
  22496=>"101100000",
  22497=>"101010111",
  22498=>"101000001",
  22499=>"011001100",
  22500=>"010011010",
  22501=>"000000111",
  22502=>"010100000",
  22503=>"000111110",
  22504=>"100011011",
  22505=>"111010011",
  22506=>"100111000",
  22507=>"000110101",
  22508=>"001110001",
  22509=>"011001000",
  22510=>"001011001",
  22511=>"111100010",
  22512=>"000011100",
  22513=>"110011101",
  22514=>"111001000",
  22515=>"000010110",
  22516=>"110110010",
  22517=>"011101111",
  22518=>"100111110",
  22519=>"011001100",
  22520=>"101111000",
  22521=>"101011110",
  22522=>"010011010",
  22523=>"100101100",
  22524=>"111100101",
  22525=>"011100000",
  22526=>"001000001",
  22527=>"001111010",
  22528=>"010011101",
  22529=>"010011010",
  22530=>"100000011",
  22531=>"111110111",
  22532=>"110111000",
  22533=>"100110000",
  22534=>"111001010",
  22535=>"010011011",
  22536=>"010110110",
  22537=>"010101111",
  22538=>"111011001",
  22539=>"010010011",
  22540=>"110011101",
  22541=>"010010010",
  22542=>"100101101",
  22543=>"110111110",
  22544=>"000010111",
  22545=>"100010001",
  22546=>"000100011",
  22547=>"000111010",
  22548=>"000100000",
  22549=>"101110011",
  22550=>"010111011",
  22551=>"111011011",
  22552=>"101010111",
  22553=>"011110110",
  22554=>"011010110",
  22555=>"101000101",
  22556=>"100100010",
  22557=>"011111000",
  22558=>"101110111",
  22559=>"101111010",
  22560=>"111100000",
  22561=>"100000100",
  22562=>"110111111",
  22563=>"000110011",
  22564=>"101100000",
  22565=>"000000101",
  22566=>"011101010",
  22567=>"100010111",
  22568=>"111011100",
  22569=>"100110111",
  22570=>"110001110",
  22571=>"000001101",
  22572=>"010000111",
  22573=>"110010111",
  22574=>"011100100",
  22575=>"111000001",
  22576=>"011011101",
  22577=>"010110100",
  22578=>"001000111",
  22579=>"010000111",
  22580=>"011000100",
  22581=>"101001100",
  22582=>"011001001",
  22583=>"001010000",
  22584=>"111111011",
  22585=>"111101111",
  22586=>"000000101",
  22587=>"011001010",
  22588=>"010110101",
  22589=>"111101100",
  22590=>"011000000",
  22591=>"010011011",
  22592=>"011001001",
  22593=>"000000010",
  22594=>"110001011",
  22595=>"010000011",
  22596=>"111000000",
  22597=>"010000000",
  22598=>"000101010",
  22599=>"001000001",
  22600=>"011110001",
  22601=>"011110111",
  22602=>"011000000",
  22603=>"000011011",
  22604=>"101010000",
  22605=>"101110011",
  22606=>"100111001",
  22607=>"110101011",
  22608=>"100010111",
  22609=>"001101111",
  22610=>"011100111",
  22611=>"100101000",
  22612=>"010100110",
  22613=>"011110111",
  22614=>"111010110",
  22615=>"011001001",
  22616=>"111000000",
  22617=>"011010000",
  22618=>"010111100",
  22619=>"010100110",
  22620=>"110100010",
  22621=>"110101101",
  22622=>"110110010",
  22623=>"000001110",
  22624=>"001011110",
  22625=>"000010011",
  22626=>"011110010",
  22627=>"111011110",
  22628=>"101000011",
  22629=>"111000000",
  22630=>"101000001",
  22631=>"100011010",
  22632=>"001011100",
  22633=>"010101101",
  22634=>"110000000",
  22635=>"110110110",
  22636=>"001010100",
  22637=>"001011000",
  22638=>"001000011",
  22639=>"101010100",
  22640=>"110100000",
  22641=>"001010100",
  22642=>"010001100",
  22643=>"011010101",
  22644=>"000100010",
  22645=>"010111110",
  22646=>"011000100",
  22647=>"001101100",
  22648=>"001110010",
  22649=>"010001101",
  22650=>"100100101",
  22651=>"101110100",
  22652=>"101000010",
  22653=>"111111010",
  22654=>"000000000",
  22655=>"001000100",
  22656=>"000100000",
  22657=>"001111001",
  22658=>"000000110",
  22659=>"000000101",
  22660=>"111101001",
  22661=>"111011000",
  22662=>"101100011",
  22663=>"100010111",
  22664=>"100011011",
  22665=>"000110100",
  22666=>"100101000",
  22667=>"000000011",
  22668=>"001111111",
  22669=>"001000100",
  22670=>"101010010",
  22671=>"110110010",
  22672=>"010111110",
  22673=>"010101011",
  22674=>"110110000",
  22675=>"101000001",
  22676=>"111110101",
  22677=>"010000101",
  22678=>"100010101",
  22679=>"001100100",
  22680=>"100100001",
  22681=>"111110110",
  22682=>"110110011",
  22683=>"001000000",
  22684=>"000010000",
  22685=>"100110100",
  22686=>"001110111",
  22687=>"110110110",
  22688=>"111001111",
  22689=>"111101110",
  22690=>"100101100",
  22691=>"001101001",
  22692=>"011011101",
  22693=>"010111110",
  22694=>"111111101",
  22695=>"011011001",
  22696=>"111011111",
  22697=>"100110011",
  22698=>"100111111",
  22699=>"101011001",
  22700=>"011100101",
  22701=>"100000000",
  22702=>"100010100",
  22703=>"000111010",
  22704=>"000010100",
  22705=>"000101110",
  22706=>"000001010",
  22707=>"000000110",
  22708=>"011011100",
  22709=>"101001110",
  22710=>"011001100",
  22711=>"000101011",
  22712=>"001000100",
  22713=>"111101011",
  22714=>"010100011",
  22715=>"111100111",
  22716=>"001101010",
  22717=>"001011111",
  22718=>"101100110",
  22719=>"111100110",
  22720=>"010010001",
  22721=>"101101110",
  22722=>"010000101",
  22723=>"011110100",
  22724=>"000001011",
  22725=>"011001001",
  22726=>"101000010",
  22727=>"110010111",
  22728=>"001000110",
  22729=>"010011001",
  22730=>"111100000",
  22731=>"111111010",
  22732=>"010000111",
  22733=>"011101101",
  22734=>"101111100",
  22735=>"110001001",
  22736=>"100100000",
  22737=>"111001001",
  22738=>"100011011",
  22739=>"011101011",
  22740=>"111101010",
  22741=>"001101011",
  22742=>"110110010",
  22743=>"101011100",
  22744=>"010000111",
  22745=>"010010000",
  22746=>"011000001",
  22747=>"010000000",
  22748=>"111001101",
  22749=>"110111101",
  22750=>"101101101",
  22751=>"110100111",
  22752=>"000111011",
  22753=>"111101111",
  22754=>"111101111",
  22755=>"001101101",
  22756=>"101100101",
  22757=>"010101100",
  22758=>"000011101",
  22759=>"111101010",
  22760=>"100110010",
  22761=>"000110110",
  22762=>"011010000",
  22763=>"001000101",
  22764=>"100010001",
  22765=>"111001110",
  22766=>"011000010",
  22767=>"001001001",
  22768=>"111111010",
  22769=>"010111000",
  22770=>"100011110",
  22771=>"100011000",
  22772=>"001110100",
  22773=>"110111111",
  22774=>"111101111",
  22775=>"000011100",
  22776=>"011001100",
  22777=>"111101000",
  22778=>"001010100",
  22779=>"110000001",
  22780=>"001000010",
  22781=>"000010011",
  22782=>"110110110",
  22783=>"011011100",
  22784=>"111011011",
  22785=>"011000010",
  22786=>"110110011",
  22787=>"011010111",
  22788=>"110000110",
  22789=>"000111111",
  22790=>"011001000",
  22791=>"101101010",
  22792=>"001010101",
  22793=>"111000100",
  22794=>"101111111",
  22795=>"010011011",
  22796=>"000010101",
  22797=>"001011011",
  22798=>"100111011",
  22799=>"000111011",
  22800=>"011110001",
  22801=>"000011000",
  22802=>"010111010",
  22803=>"111111110",
  22804=>"110101001",
  22805=>"000001001",
  22806=>"111100111",
  22807=>"000000111",
  22808=>"001000011",
  22809=>"011110001",
  22810=>"000001100",
  22811=>"001000010",
  22812=>"010100111",
  22813=>"000000111",
  22814=>"101101110",
  22815=>"110001101",
  22816=>"011010011",
  22817=>"000001111",
  22818=>"111100001",
  22819=>"110101101",
  22820=>"110001001",
  22821=>"111000001",
  22822=>"010100100",
  22823=>"101111101",
  22824=>"101001010",
  22825=>"101100101",
  22826=>"101000111",
  22827=>"010000100",
  22828=>"111111110",
  22829=>"111100000",
  22830=>"000011100",
  22831=>"111111010",
  22832=>"010011111",
  22833=>"000110100",
  22834=>"100100101",
  22835=>"010010011",
  22836=>"001110001",
  22837=>"001110110",
  22838=>"011111001",
  22839=>"011101110",
  22840=>"000000000",
  22841=>"100000000",
  22842=>"101010000",
  22843=>"000110001",
  22844=>"100100010",
  22845=>"100111110",
  22846=>"101110101",
  22847=>"110111100",
  22848=>"101010101",
  22849=>"000100100",
  22850=>"111111100",
  22851=>"001100000",
  22852=>"010000101",
  22853=>"100100111",
  22854=>"010100010",
  22855=>"101011000",
  22856=>"110101001",
  22857=>"010010010",
  22858=>"100100001",
  22859=>"010001010",
  22860=>"110000100",
  22861=>"111011000",
  22862=>"110111011",
  22863=>"000110100",
  22864=>"111011110",
  22865=>"100100001",
  22866=>"111001111",
  22867=>"001000000",
  22868=>"101011000",
  22869=>"010000110",
  22870=>"111000011",
  22871=>"000100000",
  22872=>"001000101",
  22873=>"111000111",
  22874=>"110000110",
  22875=>"101101101",
  22876=>"001111000",
  22877=>"110010101",
  22878=>"011101000",
  22879=>"010010010",
  22880=>"100000111",
  22881=>"101010101",
  22882=>"011101000",
  22883=>"001000010",
  22884=>"000011010",
  22885=>"110101010",
  22886=>"101000010",
  22887=>"000010000",
  22888=>"110001011",
  22889=>"000110000",
  22890=>"001101100",
  22891=>"001000011",
  22892=>"110000110",
  22893=>"001011001",
  22894=>"100001111",
  22895=>"000100010",
  22896=>"010110001",
  22897=>"100100001",
  22898=>"101111100",
  22899=>"101010010",
  22900=>"101000010",
  22901=>"100111010",
  22902=>"101000100",
  22903=>"000010000",
  22904=>"000100010",
  22905=>"101000010",
  22906=>"100101101",
  22907=>"001110100",
  22908=>"001100110",
  22909=>"111011111",
  22910=>"111111000",
  22911=>"111101111",
  22912=>"010000110",
  22913=>"101011110",
  22914=>"111111001",
  22915=>"001000010",
  22916=>"010010001",
  22917=>"011101000",
  22918=>"111111010",
  22919=>"100001001",
  22920=>"100100101",
  22921=>"000101101",
  22922=>"001101000",
  22923=>"101100011",
  22924=>"111100111",
  22925=>"101000000",
  22926=>"011001111",
  22927=>"001010001",
  22928=>"101010001",
  22929=>"111001110",
  22930=>"101111101",
  22931=>"000010001",
  22932=>"010100100",
  22933=>"001001111",
  22934=>"111111101",
  22935=>"100000100",
  22936=>"111110010",
  22937=>"000100101",
  22938=>"101111100",
  22939=>"100011011",
  22940=>"010101101",
  22941=>"011111111",
  22942=>"010010001",
  22943=>"011010001",
  22944=>"011101110",
  22945=>"001101110",
  22946=>"011000001",
  22947=>"110000010",
  22948=>"000010011",
  22949=>"100011010",
  22950=>"000001110",
  22951=>"101100101",
  22952=>"000101010",
  22953=>"010010110",
  22954=>"001000000",
  22955=>"001000000",
  22956=>"010000111",
  22957=>"101011000",
  22958=>"000111010",
  22959=>"000111100",
  22960=>"011110010",
  22961=>"111111101",
  22962=>"010001111",
  22963=>"011111010",
  22964=>"000100110",
  22965=>"011000100",
  22966=>"100001011",
  22967=>"101011110",
  22968=>"100110011",
  22969=>"000100110",
  22970=>"100100000",
  22971=>"011011001",
  22972=>"111000101",
  22973=>"011111101",
  22974=>"110010101",
  22975=>"110000100",
  22976=>"001011100",
  22977=>"110110110",
  22978=>"010000000",
  22979=>"101111010",
  22980=>"111100110",
  22981=>"110111111",
  22982=>"100000010",
  22983=>"000001000",
  22984=>"010001111",
  22985=>"011010010",
  22986=>"000001111",
  22987=>"100101111",
  22988=>"000010100",
  22989=>"001011000",
  22990=>"001000010",
  22991=>"000001101",
  22992=>"001010010",
  22993=>"000001001",
  22994=>"000000001",
  22995=>"010011100",
  22996=>"010001111",
  22997=>"010000110",
  22998=>"000100010",
  22999=>"111010000",
  23000=>"000010101",
  23001=>"110000111",
  23002=>"000011001",
  23003=>"110000001",
  23004=>"000100010",
  23005=>"101001111",
  23006=>"001111010",
  23007=>"000011110",
  23008=>"011110000",
  23009=>"010010010",
  23010=>"111101000",
  23011=>"010001111",
  23012=>"100001100",
  23013=>"011011010",
  23014=>"110010111",
  23015=>"100001100",
  23016=>"000101010",
  23017=>"011001110",
  23018=>"000110000",
  23019=>"001110111",
  23020=>"010101111",
  23021=>"001101101",
  23022=>"000110000",
  23023=>"101011011",
  23024=>"100110001",
  23025=>"011100100",
  23026=>"000001100",
  23027=>"010000001",
  23028=>"110111110",
  23029=>"101110110",
  23030=>"111001000",
  23031=>"111111110",
  23032=>"001100001",
  23033=>"011100000",
  23034=>"100011100",
  23035=>"011100100",
  23036=>"110101010",
  23037=>"000110000",
  23038=>"111000011",
  23039=>"001101111",
  23040=>"100111100",
  23041=>"011100011",
  23042=>"110010000",
  23043=>"100000110",
  23044=>"011000111",
  23045=>"000110111",
  23046=>"010010101",
  23047=>"000010010",
  23048=>"000000111",
  23049=>"111111000",
  23050=>"110000001",
  23051=>"000000011",
  23052=>"101100000",
  23053=>"100110010",
  23054=>"001110010",
  23055=>"001010010",
  23056=>"101110111",
  23057=>"001000001",
  23058=>"001110000",
  23059=>"101111001",
  23060=>"001001000",
  23061=>"010000010",
  23062=>"010000110",
  23063=>"110100101",
  23064=>"001010001",
  23065=>"101000010",
  23066=>"001001111",
  23067=>"000011111",
  23068=>"101100000",
  23069=>"011000101",
  23070=>"000001000",
  23071=>"101011010",
  23072=>"011101011",
  23073=>"100010101",
  23074=>"010000001",
  23075=>"000001000",
  23076=>"010110000",
  23077=>"110110010",
  23078=>"110001010",
  23079=>"000000101",
  23080=>"001111010",
  23081=>"011001100",
  23082=>"111010110",
  23083=>"110101111",
  23084=>"010110100",
  23085=>"000010110",
  23086=>"100001101",
  23087=>"110101001",
  23088=>"010100010",
  23089=>"000101000",
  23090=>"100010100",
  23091=>"100010000",
  23092=>"000010100",
  23093=>"010100011",
  23094=>"001100010",
  23095=>"001101111",
  23096=>"001110011",
  23097=>"001110101",
  23098=>"010111010",
  23099=>"010101110",
  23100=>"000011001",
  23101=>"110001111",
  23102=>"110100010",
  23103=>"110001000",
  23104=>"000110100",
  23105=>"101111011",
  23106=>"111111111",
  23107=>"001010110",
  23108=>"100011010",
  23109=>"100110011",
  23110=>"100010101",
  23111=>"111011101",
  23112=>"100011010",
  23113=>"000011100",
  23114=>"111010100",
  23115=>"100010100",
  23116=>"000110101",
  23117=>"110000100",
  23118=>"010000000",
  23119=>"100011001",
  23120=>"101111110",
  23121=>"010110101",
  23122=>"000111010",
  23123=>"001010101",
  23124=>"011100010",
  23125=>"010001100",
  23126=>"000110110",
  23127=>"110100010",
  23128=>"110100010",
  23129=>"100011111",
  23130=>"000000010",
  23131=>"100010111",
  23132=>"010110000",
  23133=>"010111011",
  23134=>"000101001",
  23135=>"011000000",
  23136=>"100001000",
  23137=>"110100011",
  23138=>"101111011",
  23139=>"111110101",
  23140=>"111001011",
  23141=>"011111100",
  23142=>"001011111",
  23143=>"010110111",
  23144=>"000000100",
  23145=>"111101101",
  23146=>"101100101",
  23147=>"001101110",
  23148=>"100100001",
  23149=>"011011100",
  23150=>"001101100",
  23151=>"001100001",
  23152=>"100010010",
  23153=>"011011010",
  23154=>"100011010",
  23155=>"100000111",
  23156=>"001101001",
  23157=>"010001011",
  23158=>"111101000",
  23159=>"000000000",
  23160=>"101010010",
  23161=>"010111101",
  23162=>"110110111",
  23163=>"101010001",
  23164=>"011000011",
  23165=>"000000100",
  23166=>"100100110",
  23167=>"110011000",
  23168=>"011100001",
  23169=>"111011011",
  23170=>"001010001",
  23171=>"000000000",
  23172=>"111001000",
  23173=>"000010000",
  23174=>"110101010",
  23175=>"011100010",
  23176=>"111000000",
  23177=>"100110111",
  23178=>"000001000",
  23179=>"000101000",
  23180=>"110000000",
  23181=>"100000101",
  23182=>"101100000",
  23183=>"011000101",
  23184=>"010010110",
  23185=>"011011000",
  23186=>"011100001",
  23187=>"100100111",
  23188=>"111010100",
  23189=>"101001101",
  23190=>"110000010",
  23191=>"000001101",
  23192=>"011000001",
  23193=>"101111111",
  23194=>"110001111",
  23195=>"010010001",
  23196=>"001010000",
  23197=>"111111111",
  23198=>"000011000",
  23199=>"101001001",
  23200=>"110110111",
  23201=>"000010000",
  23202=>"010111001",
  23203=>"000011000",
  23204=>"100101001",
  23205=>"011000010",
  23206=>"000111010",
  23207=>"101010000",
  23208=>"110000000",
  23209=>"010101100",
  23210=>"101100110",
  23211=>"111010000",
  23212=>"011111111",
  23213=>"011010010",
  23214=>"000111001",
  23215=>"101011010",
  23216=>"100111100",
  23217=>"100000010",
  23218=>"000101110",
  23219=>"011000101",
  23220=>"011100110",
  23221=>"000001001",
  23222=>"111000111",
  23223=>"111101000",
  23224=>"111101100",
  23225=>"000000100",
  23226=>"100100110",
  23227=>"000110001",
  23228=>"000110110",
  23229=>"111001111",
  23230=>"011011101",
  23231=>"001100110",
  23232=>"010011101",
  23233=>"011100000",
  23234=>"110110110",
  23235=>"000001010",
  23236=>"100000000",
  23237=>"011100111",
  23238=>"110110111",
  23239=>"010100010",
  23240=>"000000010",
  23241=>"010100001",
  23242=>"000010111",
  23243=>"000110001",
  23244=>"100000000",
  23245=>"001001101",
  23246=>"110001011",
  23247=>"101010101",
  23248=>"000111001",
  23249=>"010111011",
  23250=>"100011001",
  23251=>"001001001",
  23252=>"101101110",
  23253=>"011100001",
  23254=>"010110111",
  23255=>"100010110",
  23256=>"101100101",
  23257=>"110101111",
  23258=>"000011001",
  23259=>"100110000",
  23260=>"110111101",
  23261=>"100001010",
  23262=>"100010011",
  23263=>"100110100",
  23264=>"000010101",
  23265=>"110101101",
  23266=>"110100000",
  23267=>"101111011",
  23268=>"000000110",
  23269=>"101000001",
  23270=>"110010100",
  23271=>"101110110",
  23272=>"100000101",
  23273=>"111011110",
  23274=>"011110001",
  23275=>"110010000",
  23276=>"001000110",
  23277=>"100011001",
  23278=>"010010010",
  23279=>"000010111",
  23280=>"100100001",
  23281=>"100010101",
  23282=>"000111110",
  23283=>"011100000",
  23284=>"000000001",
  23285=>"100000110",
  23286=>"010110111",
  23287=>"111101001",
  23288=>"010001010",
  23289=>"100011111",
  23290=>"111011001",
  23291=>"110101000",
  23292=>"111111111",
  23293=>"111111111",
  23294=>"110011010",
  23295=>"010000001",
  23296=>"101010011",
  23297=>"011101111",
  23298=>"010001000",
  23299=>"011010101",
  23300=>"101100000",
  23301=>"111000011",
  23302=>"011101100",
  23303=>"110110011",
  23304=>"010111000",
  23305=>"111101011",
  23306=>"010001011",
  23307=>"010000010",
  23308=>"110110110",
  23309=>"101100101",
  23310=>"000000110",
  23311=>"101111000",
  23312=>"011001010",
  23313=>"101000100",
  23314=>"001010011",
  23315=>"110100010",
  23316=>"110110001",
  23317=>"001001001",
  23318=>"000010110",
  23319=>"101011000",
  23320=>"011101011",
  23321=>"110101011",
  23322=>"000010010",
  23323=>"000010001",
  23324=>"000101110",
  23325=>"011101101",
  23326=>"011001000",
  23327=>"111010000",
  23328=>"000011001",
  23329=>"000100111",
  23330=>"011110111",
  23331=>"100111100",
  23332=>"101101110",
  23333=>"001111111",
  23334=>"010001100",
  23335=>"000001111",
  23336=>"111101101",
  23337=>"001000100",
  23338=>"011111101",
  23339=>"001110000",
  23340=>"000111111",
  23341=>"100011101",
  23342=>"110110011",
  23343=>"110100000",
  23344=>"110000000",
  23345=>"000011111",
  23346=>"010000100",
  23347=>"110011000",
  23348=>"111101101",
  23349=>"100010101",
  23350=>"010010010",
  23351=>"011111101",
  23352=>"011110000",
  23353=>"000000001",
  23354=>"001110111",
  23355=>"010110111",
  23356=>"110010100",
  23357=>"101111011",
  23358=>"100101101",
  23359=>"001101101",
  23360=>"111011100",
  23361=>"111010001",
  23362=>"000000110",
  23363=>"010110000",
  23364=>"111000111",
  23365=>"011111011",
  23366=>"111101111",
  23367=>"001111011",
  23368=>"110010010",
  23369=>"010001001",
  23370=>"111001011",
  23371=>"101111001",
  23372=>"010010000",
  23373=>"001001111",
  23374=>"111000010",
  23375=>"101100000",
  23376=>"110110000",
  23377=>"011010111",
  23378=>"001011110",
  23379=>"100110000",
  23380=>"010010011",
  23381=>"110010000",
  23382=>"101001000",
  23383=>"101100010",
  23384=>"010111001",
  23385=>"110010110",
  23386=>"110110110",
  23387=>"111010000",
  23388=>"011101100",
  23389=>"111011010",
  23390=>"001100101",
  23391=>"101000001",
  23392=>"000101001",
  23393=>"110110010",
  23394=>"001000101",
  23395=>"010000001",
  23396=>"111000000",
  23397=>"010001001",
  23398=>"110110011",
  23399=>"100111101",
  23400=>"011001110",
  23401=>"111111001",
  23402=>"010010000",
  23403=>"011110101",
  23404=>"001001010",
  23405=>"010000000",
  23406=>"000110000",
  23407=>"010101111",
  23408=>"110010101",
  23409=>"001010000",
  23410=>"011101111",
  23411=>"010001001",
  23412=>"000110000",
  23413=>"010011001",
  23414=>"101010001",
  23415=>"010011100",
  23416=>"010010000",
  23417=>"110111111",
  23418=>"001111000",
  23419=>"101001111",
  23420=>"000000000",
  23421=>"010110010",
  23422=>"000111100",
  23423=>"110011111",
  23424=>"000000100",
  23425=>"000100110",
  23426=>"110110000",
  23427=>"110100011",
  23428=>"100110000",
  23429=>"001000110",
  23430=>"100100110",
  23431=>"100011011",
  23432=>"111100110",
  23433=>"000000111",
  23434=>"100011110",
  23435=>"000101100",
  23436=>"101101010",
  23437=>"001111000",
  23438=>"000100000",
  23439=>"010011111",
  23440=>"110100110",
  23441=>"010100110",
  23442=>"000010111",
  23443=>"111100100",
  23444=>"000111000",
  23445=>"011100111",
  23446=>"000010100",
  23447=>"011000011",
  23448=>"011111000",
  23449=>"111001111",
  23450=>"100000011",
  23451=>"100000000",
  23452=>"100010010",
  23453=>"010110011",
  23454=>"100010111",
  23455=>"001000101",
  23456=>"111000011",
  23457=>"101001111",
  23458=>"010010001",
  23459=>"011010010",
  23460=>"100011000",
  23461=>"010100011",
  23462=>"110001110",
  23463=>"010100010",
  23464=>"001000111",
  23465=>"010001100",
  23466=>"001101001",
  23467=>"111011111",
  23468=>"010000010",
  23469=>"001001100",
  23470=>"000000000",
  23471=>"001010111",
  23472=>"111000101",
  23473=>"100011101",
  23474=>"100001000",
  23475=>"000110010",
  23476=>"111011100",
  23477=>"010010001",
  23478=>"000101101",
  23479=>"000010101",
  23480=>"001101111",
  23481=>"101101010",
  23482=>"011101001",
  23483=>"001100111",
  23484=>"000010111",
  23485=>"101101111",
  23486=>"110100001",
  23487=>"100010110",
  23488=>"011101001",
  23489=>"001110101",
  23490=>"001111111",
  23491=>"000010001",
  23492=>"110010111",
  23493=>"001100101",
  23494=>"011000101",
  23495=>"011000000",
  23496=>"000001000",
  23497=>"110000000",
  23498=>"000000110",
  23499=>"111101110",
  23500=>"010111010",
  23501=>"110101100",
  23502=>"000001100",
  23503=>"111101100",
  23504=>"100111010",
  23505=>"011111111",
  23506=>"111101010",
  23507=>"110100100",
  23508=>"111000001",
  23509=>"110011010",
  23510=>"000011110",
  23511=>"111110110",
  23512=>"010010110",
  23513=>"101100101",
  23514=>"111110001",
  23515=>"010100000",
  23516=>"101111011",
  23517=>"000001100",
  23518=>"001011110",
  23519=>"111110000",
  23520=>"001010110",
  23521=>"011001111",
  23522=>"100110100",
  23523=>"011001110",
  23524=>"100111011",
  23525=>"010110000",
  23526=>"101100001",
  23527=>"110011000",
  23528=>"010000000",
  23529=>"101011100",
  23530=>"000001100",
  23531=>"110010110",
  23532=>"011000101",
  23533=>"001110001",
  23534=>"000101011",
  23535=>"001111111",
  23536=>"100111111",
  23537=>"101001001",
  23538=>"000111010",
  23539=>"001010001",
  23540=>"010111110",
  23541=>"100111100",
  23542=>"011010000",
  23543=>"111010110",
  23544=>"010010100",
  23545=>"110010000",
  23546=>"000000101",
  23547=>"111101111",
  23548=>"001110000",
  23549=>"000100010",
  23550=>"011001111",
  23551=>"100000110",
  23552=>"011001100",
  23553=>"101010011",
  23554=>"010000110",
  23555=>"001111110",
  23556=>"000100000",
  23557=>"111000101",
  23558=>"010001001",
  23559=>"110101111",
  23560=>"001101001",
  23561=>"100001110",
  23562=>"001100111",
  23563=>"111000011",
  23564=>"011111110",
  23565=>"110011011",
  23566=>"001011101",
  23567=>"011110100",
  23568=>"100101101",
  23569=>"110010010",
  23570=>"110010011",
  23571=>"111000010",
  23572=>"010100110",
  23573=>"010101111",
  23574=>"101110010",
  23575=>"100100011",
  23576=>"111011000",
  23577=>"001001101",
  23578=>"011101001",
  23579=>"111100010",
  23580=>"001010101",
  23581=>"101100001",
  23582=>"010101110",
  23583=>"101100001",
  23584=>"110100010",
  23585=>"000010110",
  23586=>"000000001",
  23587=>"010010001",
  23588=>"001110101",
  23589=>"100010001",
  23590=>"100110000",
  23591=>"100010010",
  23592=>"000110000",
  23593=>"000001101",
  23594=>"001010101",
  23595=>"101111001",
  23596=>"101100011",
  23597=>"000010000",
  23598=>"011001110",
  23599=>"010010000",
  23600=>"111010010",
  23601=>"110101001",
  23602=>"111100010",
  23603=>"001111011",
  23604=>"100000110",
  23605=>"000111010",
  23606=>"101011001",
  23607=>"011111001",
  23608=>"111001101",
  23609=>"001000001",
  23610=>"010111111",
  23611=>"001010001",
  23612=>"011010101",
  23613=>"101101101",
  23614=>"110011101",
  23615=>"101000000",
  23616=>"000100111",
  23617=>"000101000",
  23618=>"101111011",
  23619=>"011000100",
  23620=>"011000000",
  23621=>"111001110",
  23622=>"011101111",
  23623=>"101011000",
  23624=>"111011110",
  23625=>"100100101",
  23626=>"000000000",
  23627=>"111000000",
  23628=>"100110011",
  23629=>"000101111",
  23630=>"010101000",
  23631=>"000101100",
  23632=>"001010100",
  23633=>"010000110",
  23634=>"110100010",
  23635=>"111010001",
  23636=>"001111111",
  23637=>"011001110",
  23638=>"000111011",
  23639=>"011100110",
  23640=>"110111000",
  23641=>"111001011",
  23642=>"011100111",
  23643=>"110001101",
  23644=>"000000000",
  23645=>"010100110",
  23646=>"110001110",
  23647=>"001111000",
  23648=>"000010011",
  23649=>"001101000",
  23650=>"011100000",
  23651=>"010011001",
  23652=>"110101000",
  23653=>"101101100",
  23654=>"100101011",
  23655=>"111110000",
  23656=>"000011000",
  23657=>"000010111",
  23658=>"010010001",
  23659=>"001110001",
  23660=>"000001110",
  23661=>"101111010",
  23662=>"101000000",
  23663=>"010010101",
  23664=>"010000000",
  23665=>"001010000",
  23666=>"000000010",
  23667=>"110011100",
  23668=>"111110100",
  23669=>"100111000",
  23670=>"111111010",
  23671=>"101000000",
  23672=>"000101011",
  23673=>"111110000",
  23674=>"110101011",
  23675=>"100001101",
  23676=>"000001111",
  23677=>"110001010",
  23678=>"101111001",
  23679=>"111001100",
  23680=>"011000011",
  23681=>"011010011",
  23682=>"010101011",
  23683=>"001011010",
  23684=>"000000100",
  23685=>"011011101",
  23686=>"100111010",
  23687=>"010000011",
  23688=>"100000110",
  23689=>"000010111",
  23690=>"100010001",
  23691=>"100110111",
  23692=>"010000010",
  23693=>"111110011",
  23694=>"001001111",
  23695=>"101010111",
  23696=>"101111110",
  23697=>"111000010",
  23698=>"001110000",
  23699=>"111101101",
  23700=>"111111110",
  23701=>"111011111",
  23702=>"111010100",
  23703=>"011101110",
  23704=>"011101001",
  23705=>"000100010",
  23706=>"111011100",
  23707=>"001111011",
  23708=>"000100010",
  23709=>"101101100",
  23710=>"011001011",
  23711=>"101001010",
  23712=>"101100100",
  23713=>"010000100",
  23714=>"010000000",
  23715=>"010011010",
  23716=>"000000110",
  23717=>"110001011",
  23718=>"010100011",
  23719=>"110100010",
  23720=>"000001101",
  23721=>"111000100",
  23722=>"000101101",
  23723=>"000000100",
  23724=>"111101011",
  23725=>"010010011",
  23726=>"011110010",
  23727=>"100010101",
  23728=>"000000000",
  23729=>"111010110",
  23730=>"011011011",
  23731=>"100001110",
  23732=>"111010110",
  23733=>"101001100",
  23734=>"111100111",
  23735=>"101011111",
  23736=>"110000101",
  23737=>"101101111",
  23738=>"010111011",
  23739=>"000000001",
  23740=>"100101000",
  23741=>"010000111",
  23742=>"001110011",
  23743=>"000001111",
  23744=>"000101100",
  23745=>"111111000",
  23746=>"011110100",
  23747=>"001111101",
  23748=>"101101110",
  23749=>"001010010",
  23750=>"010010010",
  23751=>"110000111",
  23752=>"001000011",
  23753=>"110100001",
  23754=>"100000110",
  23755=>"101011100",
  23756=>"001101001",
  23757=>"000001111",
  23758=>"001010011",
  23759=>"111010100",
  23760=>"110011110",
  23761=>"111111101",
  23762=>"100000101",
  23763=>"111000100",
  23764=>"011011101",
  23765=>"011101001",
  23766=>"011111010",
  23767=>"100100111",
  23768=>"001010100",
  23769=>"111010110",
  23770=>"000110101",
  23771=>"011111101",
  23772=>"000111011",
  23773=>"010001100",
  23774=>"100000000",
  23775=>"100100100",
  23776=>"110010010",
  23777=>"101001011",
  23778=>"111111101",
  23779=>"010100010",
  23780=>"010110000",
  23781=>"101111100",
  23782=>"110101100",
  23783=>"101101110",
  23784=>"000011101",
  23785=>"000010110",
  23786=>"000110011",
  23787=>"110001111",
  23788=>"110110000",
  23789=>"000110110",
  23790=>"011011101",
  23791=>"101110010",
  23792=>"111001001",
  23793=>"010000001",
  23794=>"010110100",
  23795=>"001001000",
  23796=>"100110101",
  23797=>"110111111",
  23798=>"000010010",
  23799=>"011110100",
  23800=>"001100111",
  23801=>"010011100",
  23802=>"100010100",
  23803=>"000001101",
  23804=>"111101010",
  23805=>"111100101",
  23806=>"100100001",
  23807=>"111111010",
  23808=>"111010111",
  23809=>"001000001",
  23810=>"111001111",
  23811=>"010010001",
  23812=>"111000101",
  23813=>"000010010",
  23814=>"000110000",
  23815=>"110000100",
  23816=>"000111110",
  23817=>"110011010",
  23818=>"101110100",
  23819=>"000011000",
  23820=>"101000000",
  23821=>"100101001",
  23822=>"000101000",
  23823=>"111101101",
  23824=>"000101101",
  23825=>"011001100",
  23826=>"100101000",
  23827=>"111101010",
  23828=>"101001000",
  23829=>"010011101",
  23830=>"000000100",
  23831=>"101000010",
  23832=>"100010001",
  23833=>"101110001",
  23834=>"000000101",
  23835=>"101000000",
  23836=>"010111111",
  23837=>"011111000",
  23838=>"100001000",
  23839=>"111000010",
  23840=>"000100110",
  23841=>"000000110",
  23842=>"111101111",
  23843=>"001111111",
  23844=>"100011000",
  23845=>"101001110",
  23846=>"000000101",
  23847=>"110010110",
  23848=>"000001001",
  23849=>"011000011",
  23850=>"001001101",
  23851=>"111001001",
  23852=>"111111011",
  23853=>"101001101",
  23854=>"000010000",
  23855=>"111110100",
  23856=>"010000101",
  23857=>"100010100",
  23858=>"101010100",
  23859=>"010000000",
  23860=>"010101111",
  23861=>"111010011",
  23862=>"100100110",
  23863=>"011010111",
  23864=>"000010000",
  23865=>"000010001",
  23866=>"000000110",
  23867=>"101010100",
  23868=>"100011111",
  23869=>"011010101",
  23870=>"110100000",
  23871=>"100101000",
  23872=>"000110110",
  23873=>"100000001",
  23874=>"011001100",
  23875=>"111011000",
  23876=>"011101111",
  23877=>"111110101",
  23878=>"100000000",
  23879=>"000010001",
  23880=>"001001110",
  23881=>"100001111",
  23882=>"100101010",
  23883=>"101111111",
  23884=>"010101011",
  23885=>"101101000",
  23886=>"100010010",
  23887=>"000100010",
  23888=>"101100100",
  23889=>"100101101",
  23890=>"010011100",
  23891=>"111010010",
  23892=>"000100000",
  23893=>"011100010",
  23894=>"111100100",
  23895=>"101010111",
  23896=>"011001110",
  23897=>"101001111",
  23898=>"010111100",
  23899=>"010111001",
  23900=>"011010010",
  23901=>"110000111",
  23902=>"110011011",
  23903=>"001000010",
  23904=>"010001110",
  23905=>"110101100",
  23906=>"010110111",
  23907=>"010011000",
  23908=>"001001011",
  23909=>"110001100",
  23910=>"110111111",
  23911=>"100101111",
  23912=>"011110100",
  23913=>"111010001",
  23914=>"001000100",
  23915=>"011000010",
  23916=>"111001111",
  23917=>"010011101",
  23918=>"010001000",
  23919=>"010010011",
  23920=>"110010100",
  23921=>"110110100",
  23922=>"101110000",
  23923=>"000001110",
  23924=>"010111001",
  23925=>"011101000",
  23926=>"010001001",
  23927=>"101010101",
  23928=>"011000000",
  23929=>"111110111",
  23930=>"010010101",
  23931=>"000101100",
  23932=>"000110111",
  23933=>"011101101",
  23934=>"101010111",
  23935=>"000101001",
  23936=>"111110010",
  23937=>"001001010",
  23938=>"110001100",
  23939=>"000010101",
  23940=>"101100000",
  23941=>"000001001",
  23942=>"111100011",
  23943=>"001000110",
  23944=>"001011010",
  23945=>"100110111",
  23946=>"011011011",
  23947=>"001100001",
  23948=>"101001110",
  23949=>"011111010",
  23950=>"010001110",
  23951=>"100101001",
  23952=>"101001011",
  23953=>"101000011",
  23954=>"101001101",
  23955=>"000000111",
  23956=>"010011010",
  23957=>"011110110",
  23958=>"100101011",
  23959=>"000100001",
  23960=>"110010111",
  23961=>"011011010",
  23962=>"011000111",
  23963=>"100000001",
  23964=>"101110010",
  23965=>"101001001",
  23966=>"100111111",
  23967=>"100110001",
  23968=>"101111110",
  23969=>"001111000",
  23970=>"010110000",
  23971=>"000100111",
  23972=>"011101100",
  23973=>"101001000",
  23974=>"000101000",
  23975=>"001111111",
  23976=>"001000101",
  23977=>"000100011",
  23978=>"110101010",
  23979=>"000110110",
  23980=>"011111001",
  23981=>"111001100",
  23982=>"010001001",
  23983=>"111000111",
  23984=>"010001001",
  23985=>"110000100",
  23986=>"100010110",
  23987=>"011001000",
  23988=>"010010011",
  23989=>"111100101",
  23990=>"101110110",
  23991=>"101100011",
  23992=>"110001011",
  23993=>"000100010",
  23994=>"001011111",
  23995=>"000111000",
  23996=>"100100001",
  23997=>"010111001",
  23998=>"101011001",
  23999=>"100000001",
  24000=>"100011111",
  24001=>"000010111",
  24002=>"011110000",
  24003=>"100011000",
  24004=>"111000010",
  24005=>"111001001",
  24006=>"101111001",
  24007=>"111000000",
  24008=>"011000111",
  24009=>"001011110",
  24010=>"100010000",
  24011=>"101111110",
  24012=>"001101110",
  24013=>"000100010",
  24014=>"110010110",
  24015=>"000100000",
  24016=>"011100000",
  24017=>"011101101",
  24018=>"011010001",
  24019=>"101111101",
  24020=>"101010011",
  24021=>"100010001",
  24022=>"001100101",
  24023=>"111011010",
  24024=>"111011100",
  24025=>"101010110",
  24026=>"100000111",
  24027=>"101011101",
  24028=>"111001101",
  24029=>"101000111",
  24030=>"101111110",
  24031=>"010000110",
  24032=>"100000000",
  24033=>"000000110",
  24034=>"000111000",
  24035=>"011100101",
  24036=>"000110011",
  24037=>"010101001",
  24038=>"001011011",
  24039=>"110001111",
  24040=>"101010110",
  24041=>"010011101",
  24042=>"100101001",
  24043=>"001100001",
  24044=>"000000101",
  24045=>"100001001",
  24046=>"001100100",
  24047=>"100001000",
  24048=>"000011011",
  24049=>"100100011",
  24050=>"111100001",
  24051=>"001010111",
  24052=>"011001001",
  24053=>"111001010",
  24054=>"000001010",
  24055=>"001011110",
  24056=>"110101110",
  24057=>"001100011",
  24058=>"100010011",
  24059=>"110110011",
  24060=>"001001010",
  24061=>"011110111",
  24062=>"001001110",
  24063=>"011011100",
  24064=>"001001101",
  24065=>"101111011",
  24066=>"000010010",
  24067=>"100011000",
  24068=>"100001010",
  24069=>"110111011",
  24070=>"100001101",
  24071=>"000000111",
  24072=>"110010101",
  24073=>"101011111",
  24074=>"101010100",
  24075=>"100001000",
  24076=>"011001011",
  24077=>"101010001",
  24078=>"011110000",
  24079=>"001101011",
  24080=>"001101000",
  24081=>"010000000",
  24082=>"000111001",
  24083=>"101111001",
  24084=>"100010111",
  24085=>"011000011",
  24086=>"111110101",
  24087=>"001000100",
  24088=>"001101110",
  24089=>"111111110",
  24090=>"000010110",
  24091=>"010011010",
  24092=>"111001111",
  24093=>"000010011",
  24094=>"000110011",
  24095=>"011011110",
  24096=>"001001000",
  24097=>"010111000",
  24098=>"010011101",
  24099=>"110101101",
  24100=>"000110001",
  24101=>"110111101",
  24102=>"101011111",
  24103=>"000011110",
  24104=>"110101101",
  24105=>"001010101",
  24106=>"101111111",
  24107=>"111010001",
  24108=>"101110100",
  24109=>"000010001",
  24110=>"011101000",
  24111=>"001001111",
  24112=>"101010001",
  24113=>"101101100",
  24114=>"000011000",
  24115=>"101100100",
  24116=>"110000011",
  24117=>"111100110",
  24118=>"110010010",
  24119=>"000011110",
  24120=>"101100111",
  24121=>"011111010",
  24122=>"001111001",
  24123=>"010110001",
  24124=>"110110001",
  24125=>"100111111",
  24126=>"011001110",
  24127=>"100010101",
  24128=>"110100110",
  24129=>"101011000",
  24130=>"001101011",
  24131=>"110010000",
  24132=>"111000001",
  24133=>"101000111",
  24134=>"101110001",
  24135=>"011111111",
  24136=>"110111010",
  24137=>"111011011",
  24138=>"011101000",
  24139=>"110100100",
  24140=>"110101011",
  24141=>"110111000",
  24142=>"000011100",
  24143=>"010000010",
  24144=>"001100111",
  24145=>"100100110",
  24146=>"110011100",
  24147=>"101101101",
  24148=>"110111111",
  24149=>"101111110",
  24150=>"010001001",
  24151=>"110111111",
  24152=>"011011101",
  24153=>"000110001",
  24154=>"101101111",
  24155=>"110010110",
  24156=>"100011101",
  24157=>"101001011",
  24158=>"101010110",
  24159=>"010011010",
  24160=>"010011101",
  24161=>"100001111",
  24162=>"001100110",
  24163=>"010011000",
  24164=>"000001001",
  24165=>"100101010",
  24166=>"110110110",
  24167=>"100001111",
  24168=>"000000011",
  24169=>"100011111",
  24170=>"110100011",
  24171=>"011110101",
  24172=>"001001001",
  24173=>"010010001",
  24174=>"101100101",
  24175=>"001011011",
  24176=>"000110011",
  24177=>"000110001",
  24178=>"101100011",
  24179=>"111010010",
  24180=>"111000100",
  24181=>"010111100",
  24182=>"110100001",
  24183=>"111111111",
  24184=>"111100011",
  24185=>"100000010",
  24186=>"001000100",
  24187=>"010000110",
  24188=>"000001001",
  24189=>"010110001",
  24190=>"100101110",
  24191=>"100000000",
  24192=>"110001101",
  24193=>"111101100",
  24194=>"101111101",
  24195=>"010011101",
  24196=>"111010011",
  24197=>"111001101",
  24198=>"000001110",
  24199=>"100110001",
  24200=>"100100100",
  24201=>"001011010",
  24202=>"010101111",
  24203=>"100110001",
  24204=>"000110011",
  24205=>"101100011",
  24206=>"111011000",
  24207=>"101000111",
  24208=>"111110111",
  24209=>"101010101",
  24210=>"111100110",
  24211=>"110101011",
  24212=>"000000111",
  24213=>"001000101",
  24214=>"011111110",
  24215=>"010100000",
  24216=>"010111111",
  24217=>"111111001",
  24218=>"110000001",
  24219=>"110111111",
  24220=>"000110110",
  24221=>"100010010",
  24222=>"100011000",
  24223=>"001101111",
  24224=>"100100111",
  24225=>"010010110",
  24226=>"001111110",
  24227=>"010001100",
  24228=>"101001100",
  24229=>"011000111",
  24230=>"111111000",
  24231=>"000010100",
  24232=>"101001001",
  24233=>"001110101",
  24234=>"110100000",
  24235=>"101001001",
  24236=>"101111101",
  24237=>"010001000",
  24238=>"101010100",
  24239=>"100001100",
  24240=>"011010000",
  24241=>"011001001",
  24242=>"001100001",
  24243=>"000010100",
  24244=>"110010001",
  24245=>"101000001",
  24246=>"100011110",
  24247=>"010101011",
  24248=>"011110101",
  24249=>"011110000",
  24250=>"000111000",
  24251=>"001111100",
  24252=>"111111010",
  24253=>"111100000",
  24254=>"110010111",
  24255=>"101001101",
  24256=>"110110011",
  24257=>"011010111",
  24258=>"110000001",
  24259=>"001011000",
  24260=>"101001010",
  24261=>"100001011",
  24262=>"100100001",
  24263=>"100111111",
  24264=>"100101011",
  24265=>"111111001",
  24266=>"001011011",
  24267=>"100010010",
  24268=>"001100111",
  24269=>"111100000",
  24270=>"101000010",
  24271=>"001101001",
  24272=>"010100010",
  24273=>"001000011",
  24274=>"010010101",
  24275=>"101010101",
  24276=>"101001101",
  24277=>"010100101",
  24278=>"000111000",
  24279=>"101110101",
  24280=>"100100110",
  24281=>"010000011",
  24282=>"100000010",
  24283=>"011101010",
  24284=>"010001100",
  24285=>"100100000",
  24286=>"000001001",
  24287=>"001011000",
  24288=>"011010000",
  24289=>"100011000",
  24290=>"011011100",
  24291=>"000010100",
  24292=>"111010100",
  24293=>"001110110",
  24294=>"010011011",
  24295=>"111111110",
  24296=>"000001001",
  24297=>"100101011",
  24298=>"010000001",
  24299=>"000001100",
  24300=>"010000011",
  24301=>"001101010",
  24302=>"101101010",
  24303=>"001010111",
  24304=>"100001001",
  24305=>"010001010",
  24306=>"001000111",
  24307=>"011100110",
  24308=>"001100010",
  24309=>"011001100",
  24310=>"111111101",
  24311=>"011001100",
  24312=>"111111011",
  24313=>"110001101",
  24314=>"011001101",
  24315=>"110111000",
  24316=>"010000011",
  24317=>"011101111",
  24318=>"010000010",
  24319=>"111111111",
  24320=>"111000000",
  24321=>"010111011",
  24322=>"001000011",
  24323=>"100110100",
  24324=>"000100111",
  24325=>"011100110",
  24326=>"111001101",
  24327=>"100011100",
  24328=>"101101101",
  24329=>"110000100",
  24330=>"111111110",
  24331=>"001111110",
  24332=>"101001100",
  24333=>"110010000",
  24334=>"110000100",
  24335=>"011100010",
  24336=>"000100111",
  24337=>"110001010",
  24338=>"110110111",
  24339=>"111110000",
  24340=>"001001000",
  24341=>"010111111",
  24342=>"110001001",
  24343=>"010110000",
  24344=>"011001011",
  24345=>"000001010",
  24346=>"001100111",
  24347=>"000111101",
  24348=>"101000111",
  24349=>"110110001",
  24350=>"101001100",
  24351=>"111000100",
  24352=>"101111010",
  24353=>"101110101",
  24354=>"100010110",
  24355=>"010010111",
  24356=>"010110100",
  24357=>"010001000",
  24358=>"100100110",
  24359=>"010000110",
  24360=>"011111111",
  24361=>"111111010",
  24362=>"011011111",
  24363=>"001010100",
  24364=>"010000010",
  24365=>"011001100",
  24366=>"000001010",
  24367=>"111111110",
  24368=>"000001000",
  24369=>"110001110",
  24370=>"010101101",
  24371=>"101101110",
  24372=>"101110001",
  24373=>"001110111",
  24374=>"111101110",
  24375=>"011101101",
  24376=>"011110110",
  24377=>"101100000",
  24378=>"011100011",
  24379=>"010101100",
  24380=>"011000111",
  24381=>"101000110",
  24382=>"000100101",
  24383=>"001100110",
  24384=>"100011000",
  24385=>"011110010",
  24386=>"011101100",
  24387=>"111010101",
  24388=>"000001001",
  24389=>"001100101",
  24390=>"110011101",
  24391=>"011111100",
  24392=>"100111110",
  24393=>"010110111",
  24394=>"101000000",
  24395=>"000100001",
  24396=>"111111010",
  24397=>"000000001",
  24398=>"000110001",
  24399=>"011010000",
  24400=>"110101100",
  24401=>"100011000",
  24402=>"111111010",
  24403=>"111010010",
  24404=>"101001011",
  24405=>"000100110",
  24406=>"000010000",
  24407=>"101000101",
  24408=>"111011101",
  24409=>"010110011",
  24410=>"000100000",
  24411=>"111111100",
  24412=>"000110111",
  24413=>"111111110",
  24414=>"110111111",
  24415=>"001110000",
  24416=>"011011101",
  24417=>"101100110",
  24418=>"101110000",
  24419=>"100110000",
  24420=>"010001101",
  24421=>"010011000",
  24422=>"011100000",
  24423=>"110101000",
  24424=>"000000011",
  24425=>"110001111",
  24426=>"111111001",
  24427=>"101010111",
  24428=>"100101111",
  24429=>"011110011",
  24430=>"010111110",
  24431=>"100010010",
  24432=>"001011111",
  24433=>"100100101",
  24434=>"011111001",
  24435=>"010101101",
  24436=>"000111010",
  24437=>"000000100",
  24438=>"100110111",
  24439=>"100010111",
  24440=>"111001101",
  24441=>"101010101",
  24442=>"000111001",
  24443=>"001000001",
  24444=>"111111101",
  24445=>"010110010",
  24446=>"011011100",
  24447=>"000100110",
  24448=>"111100110",
  24449=>"111001111",
  24450=>"100111001",
  24451=>"111000100",
  24452=>"010010010",
  24453=>"111110111",
  24454=>"010010000",
  24455=>"010011001",
  24456=>"000100111",
  24457=>"100010100",
  24458=>"000010011",
  24459=>"000110000",
  24460=>"111110010",
  24461=>"010110000",
  24462=>"011010011",
  24463=>"100011100",
  24464=>"000011011",
  24465=>"111001011",
  24466=>"010110011",
  24467=>"110010000",
  24468=>"011111111",
  24469=>"010100011",
  24470=>"001010010",
  24471=>"001100001",
  24472=>"111101001",
  24473=>"001011011",
  24474=>"111101110",
  24475=>"110110010",
  24476=>"101011010",
  24477=>"011101101",
  24478=>"111110110",
  24479=>"100010111",
  24480=>"001001000",
  24481=>"101110001",
  24482=>"101101101",
  24483=>"011101010",
  24484=>"001011100",
  24485=>"111111011",
  24486=>"110110010",
  24487=>"100101101",
  24488=>"010111000",
  24489=>"000110010",
  24490=>"000110110",
  24491=>"101010100",
  24492=>"011111111",
  24493=>"100000010",
  24494=>"111100001",
  24495=>"100111000",
  24496=>"111010111",
  24497=>"001011011",
  24498=>"010000011",
  24499=>"010111001",
  24500=>"010011000",
  24501=>"101101101",
  24502=>"011101111",
  24503=>"111111001",
  24504=>"111001010",
  24505=>"111111101",
  24506=>"001111010",
  24507=>"010010001",
  24508=>"001010011",
  24509=>"011001111",
  24510=>"011011001",
  24511=>"111111101",
  24512=>"100000111",
  24513=>"001001011",
  24514=>"110111011",
  24515=>"010111000",
  24516=>"101000011",
  24517=>"000101110",
  24518=>"111101100",
  24519=>"011101110",
  24520=>"110000110",
  24521=>"001101010",
  24522=>"100011100",
  24523=>"011101111",
  24524=>"001100100",
  24525=>"100100100",
  24526=>"110101110",
  24527=>"001011110",
  24528=>"010101111",
  24529=>"010000100",
  24530=>"010000000",
  24531=>"001000110",
  24532=>"010010000",
  24533=>"101011011",
  24534=>"000000010",
  24535=>"000110010",
  24536=>"111110110",
  24537=>"011001011",
  24538=>"001111110",
  24539=>"011101100",
  24540=>"100000100",
  24541=>"110000000",
  24542=>"101011010",
  24543=>"000000010",
  24544=>"111111111",
  24545=>"100000101",
  24546=>"110111100",
  24547=>"010011100",
  24548=>"010010010",
  24549=>"111010101",
  24550=>"101001011",
  24551=>"001100000",
  24552=>"011110000",
  24553=>"000110101",
  24554=>"010011111",
  24555=>"010100011",
  24556=>"101111011",
  24557=>"001110010",
  24558=>"110101110",
  24559=>"101110101",
  24560=>"111010011",
  24561=>"001111110",
  24562=>"001101011",
  24563=>"110111001",
  24564=>"101111101",
  24565=>"010011001",
  24566=>"011010010",
  24567=>"000110001",
  24568=>"011011011",
  24569=>"101111010",
  24570=>"011011110",
  24571=>"101001111",
  24572=>"001111010",
  24573=>"111000100",
  24574=>"010011000",
  24575=>"110100100",
  24576=>"001000000",
  24577=>"110101110",
  24578=>"000100101",
  24579=>"010000111",
  24580=>"100101111",
  24581=>"100011100",
  24582=>"000000000",
  24583=>"001001110",
  24584=>"111110011",
  24585=>"111011100",
  24586=>"111101011",
  24587=>"100110111",
  24588=>"111100111",
  24589=>"000101111",
  24590=>"000111111",
  24591=>"010111001",
  24592=>"110101100",
  24593=>"010000000",
  24594=>"011110001",
  24595=>"010111100",
  24596=>"100010000",
  24597=>"000010011",
  24598=>"110110111",
  24599=>"111001000",
  24600=>"010100010",
  24601=>"001011001",
  24602=>"100010011",
  24603=>"100011101",
  24604=>"100110110",
  24605=>"010001001",
  24606=>"100101000",
  24607=>"110100000",
  24608=>"110111111",
  24609=>"001100000",
  24610=>"100100101",
  24611=>"010000010",
  24612=>"111000101",
  24613=>"101000000",
  24614=>"100101101",
  24615=>"111000011",
  24616=>"011010000",
  24617=>"001111001",
  24618=>"100110111",
  24619=>"100111010",
  24620=>"000000000",
  24621=>"101101011",
  24622=>"000101110",
  24623=>"001111000",
  24624=>"101011001",
  24625=>"101000001",
  24626=>"100111100",
  24627=>"110001111",
  24628=>"011010101",
  24629=>"000100011",
  24630=>"110111111",
  24631=>"011011010",
  24632=>"000011001",
  24633=>"011000001",
  24634=>"111101110",
  24635=>"011001100",
  24636=>"101000001",
  24637=>"111111110",
  24638=>"001000000",
  24639=>"101000110",
  24640=>"001011010",
  24641=>"000101100",
  24642=>"011100001",
  24643=>"001111111",
  24644=>"010010110",
  24645=>"101100000",
  24646=>"011111010",
  24647=>"010100110",
  24648=>"001000111",
  24649=>"001110100",
  24650=>"011111011",
  24651=>"001100000",
  24652=>"110011010",
  24653=>"010111011",
  24654=>"111001010",
  24655=>"100111111",
  24656=>"001000100",
  24657=>"100101000",
  24658=>"110100011",
  24659=>"111001000",
  24660=>"100001111",
  24661=>"010110110",
  24662=>"110111111",
  24663=>"001011111",
  24664=>"110100011",
  24665=>"011010001",
  24666=>"010011010",
  24667=>"111001101",
  24668=>"101100000",
  24669=>"000110100",
  24670=>"110001110",
  24671=>"110001001",
  24672=>"001111101",
  24673=>"000101101",
  24674=>"001110011",
  24675=>"110000111",
  24676=>"100010000",
  24677=>"001111110",
  24678=>"001111100",
  24679=>"000001011",
  24680=>"010110010",
  24681=>"111111111",
  24682=>"111111010",
  24683=>"001110010",
  24684=>"000101111",
  24685=>"010111000",
  24686=>"110001101",
  24687=>"000000001",
  24688=>"110000010",
  24689=>"111010110",
  24690=>"100011110",
  24691=>"011101001",
  24692=>"101101000",
  24693=>"101010101",
  24694=>"111010110",
  24695=>"001001000",
  24696=>"111101001",
  24697=>"011101001",
  24698=>"100111111",
  24699=>"010011100",
  24700=>"000010010",
  24701=>"000110010",
  24702=>"000001100",
  24703=>"000100000",
  24704=>"000000011",
  24705=>"000011011",
  24706=>"000100001",
  24707=>"100010010",
  24708=>"010100010",
  24709=>"001110101",
  24710=>"000000100",
  24711=>"110000100",
  24712=>"110110100",
  24713=>"100010111",
  24714=>"001111100",
  24715=>"010001010",
  24716=>"101010001",
  24717=>"100001001",
  24718=>"000000000",
  24719=>"001010000",
  24720=>"011001110",
  24721=>"000101011",
  24722=>"010111101",
  24723=>"101111011",
  24724=>"101101100",
  24725=>"001011101",
  24726=>"010001101",
  24727=>"000011101",
  24728=>"001010011",
  24729=>"101110111",
  24730=>"011101101",
  24731=>"110000110",
  24732=>"101100010",
  24733=>"100011000",
  24734=>"100110111",
  24735=>"100111101",
  24736=>"010000011",
  24737=>"011111100",
  24738=>"000111010",
  24739=>"110011100",
  24740=>"011101010",
  24741=>"011011001",
  24742=>"001010100",
  24743=>"000000000",
  24744=>"000100111",
  24745=>"011100011",
  24746=>"111101110",
  24747=>"110001000",
  24748=>"010011001",
  24749=>"010100000",
  24750=>"111110001",
  24751=>"111001001",
  24752=>"100101000",
  24753=>"011101101",
  24754=>"001011101",
  24755=>"001001000",
  24756=>"000101000",
  24757=>"100011111",
  24758=>"001111010",
  24759=>"001001100",
  24760=>"001101101",
  24761=>"000101010",
  24762=>"000110001",
  24763=>"010100100",
  24764=>"011001011",
  24765=>"001110101",
  24766=>"101011100",
  24767=>"100011111",
  24768=>"101101010",
  24769=>"100101001",
  24770=>"100001000",
  24771=>"000110101",
  24772=>"000000110",
  24773=>"011000010",
  24774=>"100000001",
  24775=>"110011101",
  24776=>"001100000",
  24777=>"011100010",
  24778=>"110100110",
  24779=>"111111000",
  24780=>"110101100",
  24781=>"101101110",
  24782=>"101001110",
  24783=>"101111000",
  24784=>"100010001",
  24785=>"101101001",
  24786=>"100011110",
  24787=>"011011010",
  24788=>"111010000",
  24789=>"001111111",
  24790=>"111011101",
  24791=>"110000010",
  24792=>"100000001",
  24793=>"011100100",
  24794=>"010101010",
  24795=>"100100001",
  24796=>"101001010",
  24797=>"001010101",
  24798=>"100101001",
  24799=>"111000110",
  24800=>"111111110",
  24801=>"101001101",
  24802=>"001100101",
  24803=>"001011100",
  24804=>"111010010",
  24805=>"111110110",
  24806=>"100110000",
  24807=>"001011100",
  24808=>"010111001",
  24809=>"001000110",
  24810=>"000000000",
  24811=>"001011000",
  24812=>"010001001",
  24813=>"000001101",
  24814=>"000000000",
  24815=>"010101010",
  24816=>"010001011",
  24817=>"000101110",
  24818=>"011000001",
  24819=>"001000100",
  24820=>"110110110",
  24821=>"110110111",
  24822=>"101100000",
  24823=>"100011000",
  24824=>"101011110",
  24825=>"111011000",
  24826=>"011000000",
  24827=>"010000000",
  24828=>"011001110",
  24829=>"111001111",
  24830=>"001010001",
  24831=>"100100101",
  24832=>"011110011",
  24833=>"100101001",
  24834=>"110000000",
  24835=>"010010101",
  24836=>"011111100",
  24837=>"110000011",
  24838=>"000010001",
  24839=>"000010101",
  24840=>"000110110",
  24841=>"010100110",
  24842=>"100100001",
  24843=>"100000111",
  24844=>"100010001",
  24845=>"011001000",
  24846=>"110100111",
  24847=>"111110010",
  24848=>"011000011",
  24849=>"110011000",
  24850=>"010000100",
  24851=>"111110101",
  24852=>"001001000",
  24853=>"010000101",
  24854=>"100010111",
  24855=>"101010010",
  24856=>"011001111",
  24857=>"000101110",
  24858=>"000001010",
  24859=>"011001111",
  24860=>"110111111",
  24861=>"010110110",
  24862=>"010011001",
  24863=>"101010110",
  24864=>"010000011",
  24865=>"001101011",
  24866=>"111100011",
  24867=>"010001001",
  24868=>"100010011",
  24869=>"110000101",
  24870=>"000110000",
  24871=>"110000010",
  24872=>"110111011",
  24873=>"011101011",
  24874=>"000001001",
  24875=>"110000010",
  24876=>"010010000",
  24877=>"101101111",
  24878=>"001000101",
  24879=>"111110010",
  24880=>"101110100",
  24881=>"000110111",
  24882=>"000001111",
  24883=>"001001011",
  24884=>"110101110",
  24885=>"000001011",
  24886=>"111111100",
  24887=>"100110010",
  24888=>"001010101",
  24889=>"000000001",
  24890=>"101110010",
  24891=>"011100011",
  24892=>"100111000",
  24893=>"100011000",
  24894=>"101111001",
  24895=>"010101001",
  24896=>"100110011",
  24897=>"000101111",
  24898=>"111101010",
  24899=>"110110101",
  24900=>"001011010",
  24901=>"111000010",
  24902=>"110000101",
  24903=>"000001110",
  24904=>"101010110",
  24905=>"011110000",
  24906=>"000000001",
  24907=>"100001100",
  24908=>"110110111",
  24909=>"010000001",
  24910=>"100100001",
  24911=>"110011000",
  24912=>"101000000",
  24913=>"111110100",
  24914=>"000101000",
  24915=>"001101001",
  24916=>"010101100",
  24917=>"000101101",
  24918=>"100001011",
  24919=>"100110101",
  24920=>"101110010",
  24921=>"101100101",
  24922=>"101101101",
  24923=>"100010010",
  24924=>"101001110",
  24925=>"010011100",
  24926=>"000010000",
  24927=>"010000010",
  24928=>"000010111",
  24929=>"110100000",
  24930=>"111111110",
  24931=>"101010111",
  24932=>"101100110",
  24933=>"110001101",
  24934=>"010111000",
  24935=>"111010000",
  24936=>"000000101",
  24937=>"101111101",
  24938=>"011001010",
  24939=>"111011101",
  24940=>"110100111",
  24941=>"111001110",
  24942=>"000000110",
  24943=>"100100101",
  24944=>"000101001",
  24945=>"100010111",
  24946=>"011000100",
  24947=>"010101011",
  24948=>"100010101",
  24949=>"010000010",
  24950=>"011011101",
  24951=>"111111101",
  24952=>"111111011",
  24953=>"001100011",
  24954=>"110001010",
  24955=>"101000001",
  24956=>"101101010",
  24957=>"101110100",
  24958=>"010101110",
  24959=>"101000001",
  24960=>"001001001",
  24961=>"000101101",
  24962=>"110000100",
  24963=>"111010010",
  24964=>"010000111",
  24965=>"010110000",
  24966=>"100010101",
  24967=>"111111101",
  24968=>"011010011",
  24969=>"010100001",
  24970=>"010011001",
  24971=>"000000001",
  24972=>"101110101",
  24973=>"001001010",
  24974=>"001010110",
  24975=>"000011111",
  24976=>"001101100",
  24977=>"011100101",
  24978=>"111111011",
  24979=>"000101000",
  24980=>"011101111",
  24981=>"010101000",
  24982=>"111111111",
  24983=>"100111100",
  24984=>"110011110",
  24985=>"001100000",
  24986=>"001011010",
  24987=>"001011110",
  24988=>"000111001",
  24989=>"101101101",
  24990=>"110000100",
  24991=>"110100010",
  24992=>"100101010",
  24993=>"111101111",
  24994=>"110010010",
  24995=>"000001110",
  24996=>"100110111",
  24997=>"110000000",
  24998=>"010110101",
  24999=>"011100010",
  25000=>"010101101",
  25001=>"001001011",
  25002=>"101010010",
  25003=>"000001001",
  25004=>"111100100",
  25005=>"000111001",
  25006=>"010111001",
  25007=>"011001001",
  25008=>"000000000",
  25009=>"000111000",
  25010=>"111110111",
  25011=>"011001111",
  25012=>"101010011",
  25013=>"000110011",
  25014=>"101101001",
  25015=>"101000001",
  25016=>"001101001",
  25017=>"000010000",
  25018=>"101101110",
  25019=>"100100100",
  25020=>"110110001",
  25021=>"010111011",
  25022=>"111111111",
  25023=>"011010000",
  25024=>"011010001",
  25025=>"010000110",
  25026=>"000000001",
  25027=>"111000010",
  25028=>"010000010",
  25029=>"011100100",
  25030=>"111101000",
  25031=>"001001000",
  25032=>"011000010",
  25033=>"000101101",
  25034=>"000100010",
  25035=>"000010000",
  25036=>"000111000",
  25037=>"010011001",
  25038=>"001010101",
  25039=>"001010111",
  25040=>"011010000",
  25041=>"001101111",
  25042=>"011010000",
  25043=>"101011001",
  25044=>"111110111",
  25045=>"000100110",
  25046=>"001010001",
  25047=>"001111101",
  25048=>"110101011",
  25049=>"110111101",
  25050=>"001100100",
  25051=>"010010000",
  25052=>"010000001",
  25053=>"011110110",
  25054=>"010000001",
  25055=>"010011110",
  25056=>"100110100",
  25057=>"111001101",
  25058=>"111111111",
  25059=>"100110001",
  25060=>"000110110",
  25061=>"000100110",
  25062=>"011101101",
  25063=>"100010100",
  25064=>"110111010",
  25065=>"001010001",
  25066=>"000101110",
  25067=>"001100000",
  25068=>"000011011",
  25069=>"100100011",
  25070=>"110000000",
  25071=>"101000010",
  25072=>"001111111",
  25073=>"011100001",
  25074=>"001100011",
  25075=>"101101000",
  25076=>"110001001",
  25077=>"001001110",
  25078=>"111010010",
  25079=>"000010101",
  25080=>"001011010",
  25081=>"110101111",
  25082=>"010111011",
  25083=>"001011110",
  25084=>"110100001",
  25085=>"100001110",
  25086=>"000011010",
  25087=>"011100000",
  25088=>"011110010",
  25089=>"111101000",
  25090=>"100011010",
  25091=>"110011000",
  25092=>"010111010",
  25093=>"010101100",
  25094=>"111000010",
  25095=>"111011110",
  25096=>"000001101",
  25097=>"110110111",
  25098=>"111011000",
  25099=>"010000010",
  25100=>"010010011",
  25101=>"110110100",
  25102=>"101100110",
  25103=>"000011111",
  25104=>"100110110",
  25105=>"000111011",
  25106=>"001110111",
  25107=>"110001110",
  25108=>"111100011",
  25109=>"010001010",
  25110=>"010101010",
  25111=>"101111111",
  25112=>"110111101",
  25113=>"000111101",
  25114=>"100100100",
  25115=>"010010101",
  25116=>"111000001",
  25117=>"000011111",
  25118=>"011101100",
  25119=>"010110111",
  25120=>"101011001",
  25121=>"011000010",
  25122=>"111111111",
  25123=>"100001111",
  25124=>"111011101",
  25125=>"100011011",
  25126=>"110010011",
  25127=>"111101111",
  25128=>"000001101",
  25129=>"110000001",
  25130=>"111000011",
  25131=>"110111011",
  25132=>"011100000",
  25133=>"010111101",
  25134=>"011000100",
  25135=>"101010010",
  25136=>"110011101",
  25137=>"100001000",
  25138=>"011010000",
  25139=>"110011000",
  25140=>"000110001",
  25141=>"010110001",
  25142=>"110100101",
  25143=>"010111110",
  25144=>"001000010",
  25145=>"001000010",
  25146=>"101010100",
  25147=>"000110110",
  25148=>"010101000",
  25149=>"001010001",
  25150=>"101100011",
  25151=>"010000000",
  25152=>"110011101",
  25153=>"100010010",
  25154=>"011001000",
  25155=>"100101101",
  25156=>"101010001",
  25157=>"111100000",
  25158=>"001100100",
  25159=>"101010000",
  25160=>"001000010",
  25161=>"011111011",
  25162=>"011101011",
  25163=>"111011011",
  25164=>"111011000",
  25165=>"001000110",
  25166=>"101010000",
  25167=>"100100001",
  25168=>"010111101",
  25169=>"000110000",
  25170=>"001100000",
  25171=>"011110001",
  25172=>"101110001",
  25173=>"001011101",
  25174=>"000001101",
  25175=>"100100011",
  25176=>"010000011",
  25177=>"111110100",
  25178=>"111110101",
  25179=>"101110101",
  25180=>"011100001",
  25181=>"101111111",
  25182=>"000100010",
  25183=>"110110001",
  25184=>"010000010",
  25185=>"101100100",
  25186=>"010101110",
  25187=>"011100100",
  25188=>"010101010",
  25189=>"010101110",
  25190=>"111111111",
  25191=>"001010100",
  25192=>"010000010",
  25193=>"010000001",
  25194=>"111010001",
  25195=>"111100111",
  25196=>"001010111",
  25197=>"111110000",
  25198=>"010000011",
  25199=>"110001111",
  25200=>"110001101",
  25201=>"101001011",
  25202=>"001111011",
  25203=>"001110011",
  25204=>"101000111",
  25205=>"000011110",
  25206=>"100101101",
  25207=>"100101010",
  25208=>"000101000",
  25209=>"100000000",
  25210=>"111011101",
  25211=>"101001000",
  25212=>"111010011",
  25213=>"101001111",
  25214=>"000111110",
  25215=>"001000111",
  25216=>"001111110",
  25217=>"101000101",
  25218=>"011110010",
  25219=>"011001000",
  25220=>"000010111",
  25221=>"000111100",
  25222=>"100010100",
  25223=>"100000000",
  25224=>"000111000",
  25225=>"101010011",
  25226=>"110000111",
  25227=>"001000001",
  25228=>"000000011",
  25229=>"001000001",
  25230=>"101101110",
  25231=>"001100000",
  25232=>"010001101",
  25233=>"011011010",
  25234=>"110000110",
  25235=>"000101101",
  25236=>"101101100",
  25237=>"100010010",
  25238=>"010100111",
  25239=>"111001010",
  25240=>"111111111",
  25241=>"010000100",
  25242=>"010111000",
  25243=>"011111101",
  25244=>"001100010",
  25245=>"100010000",
  25246=>"010000001",
  25247=>"000010110",
  25248=>"100111111",
  25249=>"000000001",
  25250=>"111000011",
  25251=>"011111001",
  25252=>"100001111",
  25253=>"100010000",
  25254=>"011100100",
  25255=>"101001000",
  25256=>"011011101",
  25257=>"101100100",
  25258=>"001101111",
  25259=>"001011110",
  25260=>"100001110",
  25261=>"000010110",
  25262=>"111001001",
  25263=>"101010100",
  25264=>"110011100",
  25265=>"001111001",
  25266=>"000101010",
  25267=>"111101100",
  25268=>"010101100",
  25269=>"110011110",
  25270=>"001010010",
  25271=>"110011110",
  25272=>"100000110",
  25273=>"110101111",
  25274=>"000011101",
  25275=>"011000010",
  25276=>"000100110",
  25277=>"001101001",
  25278=>"001001101",
  25279=>"000110100",
  25280=>"001010011",
  25281=>"110100110",
  25282=>"000001111",
  25283=>"111110111",
  25284=>"011111101",
  25285=>"000010010",
  25286=>"001110100",
  25287=>"000001111",
  25288=>"010010010",
  25289=>"111111111",
  25290=>"110010001",
  25291=>"011100101",
  25292=>"011110010",
  25293=>"100101101",
  25294=>"001001101",
  25295=>"100101111",
  25296=>"110010010",
  25297=>"100101100",
  25298=>"001001011",
  25299=>"001101110",
  25300=>"101000101",
  25301=>"110101010",
  25302=>"000001111",
  25303=>"001100011",
  25304=>"001011110",
  25305=>"101101101",
  25306=>"000001110",
  25307=>"101011001",
  25308=>"100001110",
  25309=>"110110001",
  25310=>"100011001",
  25311=>"000000110",
  25312=>"110001101",
  25313=>"001101001",
  25314=>"010100011",
  25315=>"011000111",
  25316=>"001100100",
  25317=>"111001000",
  25318=>"100101011",
  25319=>"111011010",
  25320=>"000110000",
  25321=>"110100111",
  25322=>"000010110",
  25323=>"001100100",
  25324=>"000000000",
  25325=>"110000101",
  25326=>"101101110",
  25327=>"010110001",
  25328=>"010001010",
  25329=>"111111110",
  25330=>"100111001",
  25331=>"101000010",
  25332=>"001000010",
  25333=>"101010011",
  25334=>"001000011",
  25335=>"111101111",
  25336=>"011010110",
  25337=>"101111111",
  25338=>"100000110",
  25339=>"110101001",
  25340=>"101111100",
  25341=>"110001011",
  25342=>"001101011",
  25343=>"110101011",
  25344=>"111100001",
  25345=>"000001011",
  25346=>"111010111",
  25347=>"010001101",
  25348=>"010011001",
  25349=>"100100000",
  25350=>"000101100",
  25351=>"110110110",
  25352=>"000001111",
  25353=>"011111100",
  25354=>"101100010",
  25355=>"000000001",
  25356=>"010100101",
  25357=>"010111011",
  25358=>"111110000",
  25359=>"000100001",
  25360=>"010000110",
  25361=>"000011011",
  25362=>"001110111",
  25363=>"010000010",
  25364=>"100011000",
  25365=>"100000011",
  25366=>"011101001",
  25367=>"000011101",
  25368=>"001100010",
  25369=>"010000110",
  25370=>"010000110",
  25371=>"110011111",
  25372=>"011101011",
  25373=>"110100001",
  25374=>"100011110",
  25375=>"010011100",
  25376=>"001110000",
  25377=>"111101010",
  25378=>"100011011",
  25379=>"001010110",
  25380=>"011101101",
  25381=>"000100111",
  25382=>"010101100",
  25383=>"001111000",
  25384=>"101100001",
  25385=>"010011011",
  25386=>"010111011",
  25387=>"011110110",
  25388=>"110001111",
  25389=>"101100100",
  25390=>"101111100",
  25391=>"010011000",
  25392=>"010101011",
  25393=>"011110000",
  25394=>"000101110",
  25395=>"000100110",
  25396=>"001011011",
  25397=>"100101110",
  25398=>"001101001",
  25399=>"011101010",
  25400=>"011111001",
  25401=>"111000111",
  25402=>"110100111",
  25403=>"000100001",
  25404=>"001001001",
  25405=>"000000101",
  25406=>"010000111",
  25407=>"101010010",
  25408=>"011001011",
  25409=>"110001000",
  25410=>"000111110",
  25411=>"010100011",
  25412=>"110101101",
  25413=>"110100010",
  25414=>"000110100",
  25415=>"100001111",
  25416=>"010010010",
  25417=>"010101001",
  25418=>"011010111",
  25419=>"000010001",
  25420=>"010001100",
  25421=>"010000110",
  25422=>"000001100",
  25423=>"110010101",
  25424=>"101110111",
  25425=>"100010101",
  25426=>"011001110",
  25427=>"001111110",
  25428=>"001100001",
  25429=>"110001010",
  25430=>"111010100",
  25431=>"100001001",
  25432=>"110001011",
  25433=>"010011110",
  25434=>"011001110",
  25435=>"111010001",
  25436=>"010010011",
  25437=>"010010100",
  25438=>"111011101",
  25439=>"000001010",
  25440=>"000011111",
  25441=>"111110110",
  25442=>"001000001",
  25443=>"111010010",
  25444=>"010101101",
  25445=>"010101010",
  25446=>"000100011",
  25447=>"111100111",
  25448=>"100001100",
  25449=>"101100001",
  25450=>"101111000",
  25451=>"011011001",
  25452=>"001011100",
  25453=>"010010111",
  25454=>"100111001",
  25455=>"110010001",
  25456=>"110000000",
  25457=>"100110001",
  25458=>"111100111",
  25459=>"111111000",
  25460=>"101001000",
  25461=>"010110100",
  25462=>"101101100",
  25463=>"000000100",
  25464=>"110010001",
  25465=>"010111011",
  25466=>"010001110",
  25467=>"011001010",
  25468=>"110110101",
  25469=>"010010001",
  25470=>"001001011",
  25471=>"100000010",
  25472=>"010010100",
  25473=>"101011100",
  25474=>"100000100",
  25475=>"110101111",
  25476=>"100100011",
  25477=>"011101110",
  25478=>"000101000",
  25479=>"111001101",
  25480=>"110001010",
  25481=>"000011110",
  25482=>"100110011",
  25483=>"111000011",
  25484=>"010101001",
  25485=>"011011101",
  25486=>"001100101",
  25487=>"110100000",
  25488=>"101101000",
  25489=>"000001001",
  25490=>"110011000",
  25491=>"100000011",
  25492=>"000011101",
  25493=>"111000001",
  25494=>"001101010",
  25495=>"110000101",
  25496=>"000100110",
  25497=>"000000110",
  25498=>"100110000",
  25499=>"011000110",
  25500=>"110010011",
  25501=>"010111010",
  25502=>"010100010",
  25503=>"110100010",
  25504=>"010100001",
  25505=>"100011110",
  25506=>"100010011",
  25507=>"111011111",
  25508=>"100111110",
  25509=>"100100000",
  25510=>"001011111",
  25511=>"000001101",
  25512=>"001111101",
  25513=>"010001111",
  25514=>"100101111",
  25515=>"100010100",
  25516=>"011000011",
  25517=>"010011000",
  25518=>"000110101",
  25519=>"011011001",
  25520=>"000011000",
  25521=>"101000111",
  25522=>"110011000",
  25523=>"001010100",
  25524=>"011111111",
  25525=>"101100111",
  25526=>"011010011",
  25527=>"111110000",
  25528=>"101011111",
  25529=>"000110110",
  25530=>"110101100",
  25531=>"001101001",
  25532=>"010110010",
  25533=>"100101000",
  25534=>"110001001",
  25535=>"010100101",
  25536=>"000011000",
  25537=>"010011101",
  25538=>"010010111",
  25539=>"111111000",
  25540=>"111101000",
  25541=>"100001110",
  25542=>"100000001",
  25543=>"101100100",
  25544=>"000000100",
  25545=>"000110001",
  25546=>"001011110",
  25547=>"110010000",
  25548=>"001110101",
  25549=>"010110100",
  25550=>"011001110",
  25551=>"011111101",
  25552=>"110011011",
  25553=>"101101110",
  25554=>"000001110",
  25555=>"100000000",
  25556=>"111111111",
  25557=>"001001001",
  25558=>"101000111",
  25559=>"001111111",
  25560=>"110001101",
  25561=>"000000011",
  25562=>"110100000",
  25563=>"110000101",
  25564=>"101000101",
  25565=>"110010010",
  25566=>"010101101",
  25567=>"000110001",
  25568=>"110011101",
  25569=>"110110111",
  25570=>"100010100",
  25571=>"010001010",
  25572=>"101011110",
  25573=>"010100100",
  25574=>"000010011",
  25575=>"010000101",
  25576=>"010100100",
  25577=>"001000101",
  25578=>"110000101",
  25579=>"101011000",
  25580=>"000110000",
  25581=>"011101010",
  25582=>"001010001",
  25583=>"010000011",
  25584=>"011101101",
  25585=>"101000000",
  25586=>"000101101",
  25587=>"011000001",
  25588=>"100111001",
  25589=>"001000101",
  25590=>"110100100",
  25591=>"000010011",
  25592=>"110001011",
  25593=>"111001111",
  25594=>"110000100",
  25595=>"011100111",
  25596=>"001011001",
  25597=>"011110101",
  25598=>"000001000",
  25599=>"110100001",
  25600=>"111001101",
  25601=>"100000011",
  25602=>"001110110",
  25603=>"101101100",
  25604=>"001011100",
  25605=>"010001111",
  25606=>"101010100",
  25607=>"111000000",
  25608=>"111110101",
  25609=>"010110110",
  25610=>"111011010",
  25611=>"110111001",
  25612=>"101010010",
  25613=>"111111110",
  25614=>"111100100",
  25615=>"101000011",
  25616=>"111000000",
  25617=>"000110001",
  25618=>"101010101",
  25619=>"000111000",
  25620=>"011001000",
  25621=>"101100001",
  25622=>"100100101",
  25623=>"110100001",
  25624=>"111000011",
  25625=>"000010001",
  25626=>"100111110",
  25627=>"010101110",
  25628=>"011111011",
  25629=>"101011101",
  25630=>"001010101",
  25631=>"100000101",
  25632=>"111111000",
  25633=>"010001110",
  25634=>"011100001",
  25635=>"000000101",
  25636=>"001011000",
  25637=>"011010010",
  25638=>"011000010",
  25639=>"101111000",
  25640=>"000000010",
  25641=>"100010111",
  25642=>"100011010",
  25643=>"110011110",
  25644=>"001000101",
  25645=>"110010000",
  25646=>"011000101",
  25647=>"001110100",
  25648=>"110000001",
  25649=>"100101000",
  25650=>"000010011",
  25651=>"000011100",
  25652=>"101100101",
  25653=>"010001011",
  25654=>"011000011",
  25655=>"100001101",
  25656=>"011000011",
  25657=>"000000000",
  25658=>"101111100",
  25659=>"000100100",
  25660=>"011111000",
  25661=>"110000110",
  25662=>"000001001",
  25663=>"110101001",
  25664=>"111011000",
  25665=>"011010001",
  25666=>"001011000",
  25667=>"011101101",
  25668=>"111110110",
  25669=>"101111111",
  25670=>"000101101",
  25671=>"000111100",
  25672=>"000011011",
  25673=>"111101010",
  25674=>"101111011",
  25675=>"100100010",
  25676=>"110000101",
  25677=>"010001100",
  25678=>"101111110",
  25679=>"111100001",
  25680=>"010011000",
  25681=>"000000101",
  25682=>"110110110",
  25683=>"111100000",
  25684=>"111111111",
  25685=>"010000100",
  25686=>"011110000",
  25687=>"110101001",
  25688=>"111101100",
  25689=>"010000111",
  25690=>"000111110",
  25691=>"000000000",
  25692=>"001100110",
  25693=>"010100000",
  25694=>"010110100",
  25695=>"010100000",
  25696=>"001101000",
  25697=>"000110101",
  25698=>"000100010",
  25699=>"101111100",
  25700=>"000000111",
  25701=>"011010110",
  25702=>"100010100",
  25703=>"110100110",
  25704=>"101011001",
  25705=>"010010110",
  25706=>"000010110",
  25707=>"101010111",
  25708=>"011100010",
  25709=>"101101011",
  25710=>"001101000",
  25711=>"100010010",
  25712=>"101010011",
  25713=>"011001110",
  25714=>"000011110",
  25715=>"110000000",
  25716=>"001011110",
  25717=>"001010001",
  25718=>"010111111",
  25719=>"010000010",
  25720=>"101100101",
  25721=>"010110111",
  25722=>"111001011",
  25723=>"101101000",
  25724=>"010111111",
  25725=>"100000011",
  25726=>"111101111",
  25727=>"001011101",
  25728=>"010001000",
  25729=>"001101100",
  25730=>"010011000",
  25731=>"011010111",
  25732=>"011010111",
  25733=>"111111101",
  25734=>"001011001",
  25735=>"111011100",
  25736=>"010100110",
  25737=>"000110000",
  25738=>"100110010",
  25739=>"111110101",
  25740=>"110001111",
  25741=>"011011011",
  25742=>"100001101",
  25743=>"110001111",
  25744=>"111110010",
  25745=>"110000100",
  25746=>"000100110",
  25747=>"100111000",
  25748=>"110000000",
  25749=>"010010110",
  25750=>"110000001",
  25751=>"010100110",
  25752=>"011100111",
  25753=>"010100111",
  25754=>"001011000",
  25755=>"101001111",
  25756=>"111110001",
  25757=>"000001101",
  25758=>"110100101",
  25759=>"010111101",
  25760=>"011110010",
  25761=>"010110000",
  25762=>"100000010",
  25763=>"011010010",
  25764=>"010011111",
  25765=>"101111000",
  25766=>"010100001",
  25767=>"111111010",
  25768=>"110000000",
  25769=>"010100111",
  25770=>"100101000",
  25771=>"101001000",
  25772=>"111010001",
  25773=>"111101100",
  25774=>"000001001",
  25775=>"100001000",
  25776=>"110010001",
  25777=>"001100101",
  25778=>"010011010",
  25779=>"110000110",
  25780=>"011111100",
  25781=>"111111110",
  25782=>"110110001",
  25783=>"010101101",
  25784=>"000100100",
  25785=>"001011100",
  25786=>"110100011",
  25787=>"001111000",
  25788=>"000101111",
  25789=>"011000111",
  25790=>"001111101",
  25791=>"100100011",
  25792=>"100011100",
  25793=>"110000101",
  25794=>"100010000",
  25795=>"110110100",
  25796=>"110000000",
  25797=>"101001010",
  25798=>"100001111",
  25799=>"001000001",
  25800=>"111011101",
  25801=>"111010010",
  25802=>"011110001",
  25803=>"000101001",
  25804=>"001110011",
  25805=>"101100001",
  25806=>"110111001",
  25807=>"000110000",
  25808=>"010010000",
  25809=>"111111101",
  25810=>"010001000",
  25811=>"111101100",
  25812=>"011011001",
  25813=>"011001101",
  25814=>"010101100",
  25815=>"110000011",
  25816=>"110111010",
  25817=>"100110101",
  25818=>"001111001",
  25819=>"001011001",
  25820=>"000010101",
  25821=>"000110110",
  25822=>"000100000",
  25823=>"101111111",
  25824=>"010011000",
  25825=>"010000000",
  25826=>"100001011",
  25827=>"011010010",
  25828=>"011101011",
  25829=>"001010101",
  25830=>"111100000",
  25831=>"011101000",
  25832=>"100100010",
  25833=>"100101011",
  25834=>"100110100",
  25835=>"100000001",
  25836=>"010110001",
  25837=>"110101000",
  25838=>"010001111",
  25839=>"010000010",
  25840=>"101110111",
  25841=>"111101011",
  25842=>"010011010",
  25843=>"110000110",
  25844=>"011101101",
  25845=>"110011011",
  25846=>"000000001",
  25847=>"010100101",
  25848=>"011010110",
  25849=>"011110000",
  25850=>"000110000",
  25851=>"000110001",
  25852=>"011010010",
  25853=>"001010101",
  25854=>"110011111",
  25855=>"001100100",
  25856=>"000110011",
  25857=>"000011001",
  25858=>"010011011",
  25859=>"000111100",
  25860=>"001110010",
  25861=>"000110100",
  25862=>"000001111",
  25863=>"001111101",
  25864=>"111111011",
  25865=>"001010110",
  25866=>"100000101",
  25867=>"001101000",
  25868=>"001111111",
  25869=>"000000001",
  25870=>"110101101",
  25871=>"100010110",
  25872=>"011110110",
  25873=>"100101111",
  25874=>"100100000",
  25875=>"111110001",
  25876=>"111110110",
  25877=>"110100100",
  25878=>"000010011",
  25879=>"100111011",
  25880=>"110101000",
  25881=>"101011101",
  25882=>"110001010",
  25883=>"000111000",
  25884=>"011011010",
  25885=>"100010100",
  25886=>"111101010",
  25887=>"101001110",
  25888=>"011110000",
  25889=>"011110110",
  25890=>"000111111",
  25891=>"000001000",
  25892=>"101111001",
  25893=>"100011100",
  25894=>"011000001",
  25895=>"011100001",
  25896=>"011011111",
  25897=>"011101001",
  25898=>"000110100",
  25899=>"001110100",
  25900=>"110101111",
  25901=>"010000010",
  25902=>"000011101",
  25903=>"001001111",
  25904=>"010000100",
  25905=>"010001101",
  25906=>"110101011",
  25907=>"000111011",
  25908=>"011100000",
  25909=>"100110001",
  25910=>"110111010",
  25911=>"111001101",
  25912=>"000000110",
  25913=>"011010000",
  25914=>"011100001",
  25915=>"011010000",
  25916=>"011011000",
  25917=>"111110111",
  25918=>"111100101",
  25919=>"001111101",
  25920=>"110110110",
  25921=>"000100010",
  25922=>"101110101",
  25923=>"001011010",
  25924=>"011011100",
  25925=>"001100011",
  25926=>"010010000",
  25927=>"111110000",
  25928=>"001001001",
  25929=>"011000100",
  25930=>"000011000",
  25931=>"101000011",
  25932=>"000011111",
  25933=>"110100010",
  25934=>"001101100",
  25935=>"110101100",
  25936=>"100111010",
  25937=>"000101101",
  25938=>"110010110",
  25939=>"001001001",
  25940=>"101111010",
  25941=>"100111111",
  25942=>"111010110",
  25943=>"001001111",
  25944=>"011100101",
  25945=>"011010111",
  25946=>"011001010",
  25947=>"101001010",
  25948=>"111001001",
  25949=>"001111111",
  25950=>"110111101",
  25951=>"111100010",
  25952=>"100110011",
  25953=>"010000111",
  25954=>"011000110",
  25955=>"011010101",
  25956=>"101010101",
  25957=>"111111000",
  25958=>"111011000",
  25959=>"111110000",
  25960=>"100101011",
  25961=>"101001101",
  25962=>"011111000",
  25963=>"111011101",
  25964=>"000000000",
  25965=>"101001101",
  25966=>"011011000",
  25967=>"111000110",
  25968=>"001101110",
  25969=>"101000010",
  25970=>"100010111",
  25971=>"101001001",
  25972=>"000111011",
  25973=>"111111011",
  25974=>"010100011",
  25975=>"100110001",
  25976=>"001000000",
  25977=>"001110101",
  25978=>"001010001",
  25979=>"000000010",
  25980=>"111101111",
  25981=>"011000001",
  25982=>"111010100",
  25983=>"101011110",
  25984=>"101111011",
  25985=>"000000000",
  25986=>"001111101",
  25987=>"000101110",
  25988=>"011000000",
  25989=>"101000100",
  25990=>"010001111",
  25991=>"001011101",
  25992=>"001111110",
  25993=>"110100000",
  25994=>"010011001",
  25995=>"101011111",
  25996=>"101010110",
  25997=>"001111010",
  25998=>"111011111",
  25999=>"111111011",
  26000=>"011111110",
  26001=>"110011110",
  26002=>"011110100",
  26003=>"001000010",
  26004=>"110101011",
  26005=>"010000000",
  26006=>"111100110",
  26007=>"000111101",
  26008=>"000111011",
  26009=>"010111110",
  26010=>"001101111",
  26011=>"001000111",
  26012=>"001011111",
  26013=>"000011000",
  26014=>"111100100",
  26015=>"010001100",
  26016=>"011010011",
  26017=>"110111110",
  26018=>"001111011",
  26019=>"100011010",
  26020=>"100101001",
  26021=>"000101000",
  26022=>"100000110",
  26023=>"010100111",
  26024=>"000010111",
  26025=>"011110101",
  26026=>"001011101",
  26027=>"011100101",
  26028=>"111111000",
  26029=>"010100110",
  26030=>"000000000",
  26031=>"010011101",
  26032=>"011001011",
  26033=>"000010101",
  26034=>"100001111",
  26035=>"100011010",
  26036=>"011000110",
  26037=>"000000001",
  26038=>"000010101",
  26039=>"000010011",
  26040=>"100010001",
  26041=>"110110110",
  26042=>"101100001",
  26043=>"101001000",
  26044=>"110101111",
  26045=>"111111100",
  26046=>"100111100",
  26047=>"000000110",
  26048=>"110000101",
  26049=>"111010110",
  26050=>"100101111",
  26051=>"000000101",
  26052=>"100110001",
  26053=>"000101111",
  26054=>"011010100",
  26055=>"000011000",
  26056=>"111000110",
  26057=>"011101000",
  26058=>"001011101",
  26059=>"011101011",
  26060=>"001111101",
  26061=>"100110110",
  26062=>"000101101",
  26063=>"010001011",
  26064=>"110001000",
  26065=>"111110111",
  26066=>"100011011",
  26067=>"011001011",
  26068=>"100001011",
  26069=>"000011001",
  26070=>"100000011",
  26071=>"111110110",
  26072=>"100111011",
  26073=>"001100111",
  26074=>"000000000",
  26075=>"010010101",
  26076=>"101111101",
  26077=>"000001010",
  26078=>"000110101",
  26079=>"111000001",
  26080=>"101011010",
  26081=>"101110100",
  26082=>"101110101",
  26083=>"011110110",
  26084=>"100111110",
  26085=>"011011001",
  26086=>"000001010",
  26087=>"010110000",
  26088=>"001101010",
  26089=>"011101111",
  26090=>"101111111",
  26091=>"010000001",
  26092=>"111101000",
  26093=>"010110101",
  26094=>"001000111",
  26095=>"101100011",
  26096=>"001111100",
  26097=>"100111010",
  26098=>"101100111",
  26099=>"000011100",
  26100=>"011011000",
  26101=>"110010110",
  26102=>"010101100",
  26103=>"111111111",
  26104=>"110110110",
  26105=>"011010101",
  26106=>"001001101",
  26107=>"010011100",
  26108=>"001000110",
  26109=>"010010111",
  26110=>"111001001",
  26111=>"110010000",
  26112=>"011000101",
  26113=>"001010100",
  26114=>"100100111",
  26115=>"011001000",
  26116=>"111001101",
  26117=>"110011110",
  26118=>"001111000",
  26119=>"000110100",
  26120=>"110110101",
  26121=>"010100101",
  26122=>"010100110",
  26123=>"010000101",
  26124=>"001011010",
  26125=>"110110111",
  26126=>"000000101",
  26127=>"101100100",
  26128=>"111100010",
  26129=>"010011110",
  26130=>"100001001",
  26131=>"000100100",
  26132=>"011100111",
  26133=>"001110001",
  26134=>"101110000",
  26135=>"001101110",
  26136=>"011111000",
  26137=>"111010001",
  26138=>"000110101",
  26139=>"000001011",
  26140=>"100100010",
  26141=>"011000011",
  26142=>"011101010",
  26143=>"110101011",
  26144=>"010000100",
  26145=>"100101001",
  26146=>"110100110",
  26147=>"010110010",
  26148=>"011110100",
  26149=>"110001111",
  26150=>"101011000",
  26151=>"001100000",
  26152=>"110000010",
  26153=>"011000010",
  26154=>"101010011",
  26155=>"101111011",
  26156=>"000111010",
  26157=>"000110100",
  26158=>"101011110",
  26159=>"001100010",
  26160=>"001101101",
  26161=>"010000110",
  26162=>"010110110",
  26163=>"110110101",
  26164=>"111101101",
  26165=>"000111101",
  26166=>"010111011",
  26167=>"111101101",
  26168=>"010101110",
  26169=>"000111000",
  26170=>"100001010",
  26171=>"000100010",
  26172=>"110100001",
  26173=>"000000000",
  26174=>"100101000",
  26175=>"101111111",
  26176=>"000110110",
  26177=>"011010110",
  26178=>"111011111",
  26179=>"101101101",
  26180=>"111011000",
  26181=>"001101100",
  26182=>"101010100",
  26183=>"100010100",
  26184=>"101101111",
  26185=>"010101111",
  26186=>"110000110",
  26187=>"100100011",
  26188=>"111110111",
  26189=>"000101100",
  26190=>"001000101",
  26191=>"100001011",
  26192=>"001011001",
  26193=>"001001000",
  26194=>"110100001",
  26195=>"001111010",
  26196=>"101101010",
  26197=>"111010011",
  26198=>"111000011",
  26199=>"001101110",
  26200=>"110111010",
  26201=>"001001011",
  26202=>"011001000",
  26203=>"101111101",
  26204=>"000011011",
  26205=>"000100111",
  26206=>"010100000",
  26207=>"100100011",
  26208=>"001100000",
  26209=>"101011000",
  26210=>"010011000",
  26211=>"010110011",
  26212=>"101110001",
  26213=>"100100001",
  26214=>"000000100",
  26215=>"111101111",
  26216=>"010001100",
  26217=>"110111101",
  26218=>"110110000",
  26219=>"110001110",
  26220=>"001101010",
  26221=>"100110011",
  26222=>"001100000",
  26223=>"001110110",
  26224=>"001111110",
  26225=>"011110101",
  26226=>"010010010",
  26227=>"001110011",
  26228=>"111001010",
  26229=>"000110111",
  26230=>"000101110",
  26231=>"100000000",
  26232=>"011010100",
  26233=>"110111001",
  26234=>"001000000",
  26235=>"000011010",
  26236=>"000000000",
  26237=>"111111100",
  26238=>"101111011",
  26239=>"010110100",
  26240=>"010100001",
  26241=>"111010101",
  26242=>"110011010",
  26243=>"101101000",
  26244=>"000000011",
  26245=>"101001101",
  26246=>"000101100",
  26247=>"100111001",
  26248=>"001100110",
  26249=>"101111011",
  26250=>"100110100",
  26251=>"000111001",
  26252=>"010000100",
  26253=>"000011010",
  26254=>"101110100",
  26255=>"101000011",
  26256=>"000010000",
  26257=>"111000100",
  26258=>"101110011",
  26259=>"100111111",
  26260=>"101001100",
  26261=>"000001010",
  26262=>"001110100",
  26263=>"101000001",
  26264=>"000011101",
  26265=>"001101011",
  26266=>"110010001",
  26267=>"001000011",
  26268=>"100111110",
  26269=>"000110001",
  26270=>"101110101",
  26271=>"110001000",
  26272=>"110000000",
  26273=>"100111111",
  26274=>"111000011",
  26275=>"010110101",
  26276=>"011000111",
  26277=>"001011111",
  26278=>"001011100",
  26279=>"000000000",
  26280=>"010011011",
  26281=>"111100011",
  26282=>"110010101",
  26283=>"000110000",
  26284=>"000010001",
  26285=>"010011010",
  26286=>"110101101",
  26287=>"111111011",
  26288=>"000110011",
  26289=>"001100011",
  26290=>"100111000",
  26291=>"110110111",
  26292=>"001100111",
  26293=>"010111000",
  26294=>"100000011",
  26295=>"011011011",
  26296=>"101011000",
  26297=>"111011101",
  26298=>"111100010",
  26299=>"010010111",
  26300=>"000100001",
  26301=>"111110101",
  26302=>"000000101",
  26303=>"011001111",
  26304=>"101001000",
  26305=>"110101111",
  26306=>"001001001",
  26307=>"001111101",
  26308=>"111001111",
  26309=>"110001000",
  26310=>"110111110",
  26311=>"111101000",
  26312=>"010011011",
  26313=>"000001111",
  26314=>"011000111",
  26315=>"111111110",
  26316=>"000000100",
  26317=>"110101000",
  26318=>"110101000",
  26319=>"111001000",
  26320=>"011110100",
  26321=>"110110110",
  26322=>"101100101",
  26323=>"111111100",
  26324=>"000101101",
  26325=>"100000100",
  26326=>"011001111",
  26327=>"101100000",
  26328=>"010110001",
  26329=>"100001101",
  26330=>"100010011",
  26331=>"000101001",
  26332=>"101110111",
  26333=>"001000100",
  26334=>"001010000",
  26335=>"000000010",
  26336=>"011110000",
  26337=>"110101100",
  26338=>"111010110",
  26339=>"010010100",
  26340=>"110100000",
  26341=>"110101000",
  26342=>"100001001",
  26343=>"110011110",
  26344=>"110001100",
  26345=>"101001101",
  26346=>"111010001",
  26347=>"001011100",
  26348=>"010000011",
  26349=>"010001010",
  26350=>"101011111",
  26351=>"001011100",
  26352=>"100011110",
  26353=>"001100011",
  26354=>"000110111",
  26355=>"010001010",
  26356=>"000100111",
  26357=>"100101111",
  26358=>"100001010",
  26359=>"100011001",
  26360=>"101011010",
  26361=>"111000000",
  26362=>"001000001",
  26363=>"100110010",
  26364=>"000010101",
  26365=>"000010000",
  26366=>"001000101",
  26367=>"111111111",
  26368=>"011110101",
  26369=>"111100011",
  26370=>"111110001",
  26371=>"011110010",
  26372=>"000010111",
  26373=>"001100110",
  26374=>"110110101",
  26375=>"110001101",
  26376=>"000101101",
  26377=>"110010110",
  26378=>"101101101",
  26379=>"100000101",
  26380=>"111011111",
  26381=>"110100010",
  26382=>"101101101",
  26383=>"001101100",
  26384=>"011010100",
  26385=>"101000010",
  26386=>"111111111",
  26387=>"011101010",
  26388=>"100100101",
  26389=>"111010100",
  26390=>"111000011",
  26391=>"000011011",
  26392=>"010110011",
  26393=>"111111100",
  26394=>"000100110",
  26395=>"000001111",
  26396=>"111100000",
  26397=>"010010011",
  26398=>"100100110",
  26399=>"100101011",
  26400=>"111101111",
  26401=>"110000101",
  26402=>"100110110",
  26403=>"001101000",
  26404=>"111011000",
  26405=>"000000010",
  26406=>"110111101",
  26407=>"100101011",
  26408=>"111011100",
  26409=>"110011010",
  26410=>"110110100",
  26411=>"010111110",
  26412=>"010101101",
  26413=>"101101000",
  26414=>"011100100",
  26415=>"010111011",
  26416=>"101000000",
  26417=>"001010101",
  26418=>"001011000",
  26419=>"000001001",
  26420=>"111010111",
  26421=>"010110101",
  26422=>"011000111",
  26423=>"011000011",
  26424=>"001001000",
  26425=>"011010100",
  26426=>"011101100",
  26427=>"101111110",
  26428=>"010100001",
  26429=>"100110100",
  26430=>"010011100",
  26431=>"110111011",
  26432=>"010010011",
  26433=>"001111110",
  26434=>"000100110",
  26435=>"111111110",
  26436=>"101000111",
  26437=>"000011011",
  26438=>"000010010",
  26439=>"100101111",
  26440=>"111011101",
  26441=>"100111001",
  26442=>"100011111",
  26443=>"001110000",
  26444=>"100011000",
  26445=>"101111110",
  26446=>"001010001",
  26447=>"010110011",
  26448=>"110010000",
  26449=>"100101110",
  26450=>"110110001",
  26451=>"100000010",
  26452=>"101011011",
  26453=>"100001111",
  26454=>"011110001",
  26455=>"110111010",
  26456=>"001100000",
  26457=>"110000010",
  26458=>"000000000",
  26459=>"000100111",
  26460=>"011001101",
  26461=>"011011011",
  26462=>"101110110",
  26463=>"011101111",
  26464=>"110111011",
  26465=>"001101101",
  26466=>"111100100",
  26467=>"010011111",
  26468=>"100001011",
  26469=>"001111101",
  26470=>"101011110",
  26471=>"000110000",
  26472=>"100010010",
  26473=>"101110111",
  26474=>"110001001",
  26475=>"001100011",
  26476=>"110111010",
  26477=>"001110001",
  26478=>"000110010",
  26479=>"111101110",
  26480=>"001010100",
  26481=>"110011011",
  26482=>"100010000",
  26483=>"111111100",
  26484=>"101110100",
  26485=>"001001000",
  26486=>"111001011",
  26487=>"011000010",
  26488=>"110111111",
  26489=>"000101011",
  26490=>"101010110",
  26491=>"010000011",
  26492=>"001011100",
  26493=>"011010000",
  26494=>"011110000",
  26495=>"110011100",
  26496=>"111101111",
  26497=>"110111111",
  26498=>"011001111",
  26499=>"001001011",
  26500=>"000111100",
  26501=>"100001010",
  26502=>"010100010",
  26503=>"010111110",
  26504=>"000111111",
  26505=>"111001111",
  26506=>"111011110",
  26507=>"010010000",
  26508=>"001001001",
  26509=>"101100011",
  26510=>"011001111",
  26511=>"000111010",
  26512=>"001100111",
  26513=>"110110100",
  26514=>"011101100",
  26515=>"110010010",
  26516=>"100001001",
  26517=>"011111011",
  26518=>"100000000",
  26519=>"101010110",
  26520=>"000010001",
  26521=>"000101010",
  26522=>"100011001",
  26523=>"001111001",
  26524=>"101110101",
  26525=>"100110000",
  26526=>"010001111",
  26527=>"101010000",
  26528=>"101010110",
  26529=>"001100100",
  26530=>"100111101",
  26531=>"111101001",
  26532=>"111100001",
  26533=>"000110110",
  26534=>"110001001",
  26535=>"110110011",
  26536=>"111111111",
  26537=>"000010000",
  26538=>"001001010",
  26539=>"100101101",
  26540=>"111001101",
  26541=>"111000101",
  26542=>"011001100",
  26543=>"110110100",
  26544=>"111110111",
  26545=>"011111000",
  26546=>"000100101",
  26547=>"110001100",
  26548=>"010101101",
  26549=>"110110101",
  26550=>"000001001",
  26551=>"001101100",
  26552=>"110000000",
  26553=>"011010000",
  26554=>"000100101",
  26555=>"101111100",
  26556=>"000101100",
  26557=>"111100000",
  26558=>"001000110",
  26559=>"110000011",
  26560=>"110111000",
  26561=>"001010010",
  26562=>"011010100",
  26563=>"000001110",
  26564=>"001010011",
  26565=>"010000101",
  26566=>"000111111",
  26567=>"101011110",
  26568=>"010101101",
  26569=>"110000000",
  26570=>"101100101",
  26571=>"000101101",
  26572=>"100100001",
  26573=>"101100100",
  26574=>"000011101",
  26575=>"100001101",
  26576=>"001000111",
  26577=>"010010111",
  26578=>"010001010",
  26579=>"100001001",
  26580=>"010010110",
  26581=>"111110011",
  26582=>"000010001",
  26583=>"001110010",
  26584=>"111110000",
  26585=>"110110010",
  26586=>"100000000",
  26587=>"101111000",
  26588=>"111110001",
  26589=>"111101000",
  26590=>"110010000",
  26591=>"000011110",
  26592=>"010000010",
  26593=>"111100011",
  26594=>"001110110",
  26595=>"001001011",
  26596=>"011010001",
  26597=>"011011000",
  26598=>"011000000",
  26599=>"010001111",
  26600=>"010001101",
  26601=>"100010000",
  26602=>"111111011",
  26603=>"101110111",
  26604=>"111110111",
  26605=>"101111100",
  26606=>"001010000",
  26607=>"100111111",
  26608=>"101011010",
  26609=>"111101100",
  26610=>"000000010",
  26611=>"001111001",
  26612=>"011100100",
  26613=>"001100100",
  26614=>"001110011",
  26615=>"100011100",
  26616=>"010000010",
  26617=>"001010000",
  26618=>"011000111",
  26619=>"111011001",
  26620=>"100001111",
  26621=>"101011110",
  26622=>"010111001",
  26623=>"011101000",
  26624=>"101000001",
  26625=>"001100110",
  26626=>"001101001",
  26627=>"010010011",
  26628=>"001001000",
  26629=>"011100110",
  26630=>"010011000",
  26631=>"100010010",
  26632=>"111100110",
  26633=>"100001111",
  26634=>"010100110",
  26635=>"111011111",
  26636=>"011100111",
  26637=>"000000101",
  26638=>"000000000",
  26639=>"101110001",
  26640=>"010100101",
  26641=>"110110100",
  26642=>"001010001",
  26643=>"010010001",
  26644=>"001000010",
  26645=>"111111101",
  26646=>"101010110",
  26647=>"111001101",
  26648=>"010101001",
  26649=>"101111001",
  26650=>"110100010",
  26651=>"111001110",
  26652=>"101001010",
  26653=>"011111111",
  26654=>"001010010",
  26655=>"000000111",
  26656=>"010100010",
  26657=>"111111001",
  26658=>"000111001",
  26659=>"101010011",
  26660=>"000000010",
  26661=>"001110110",
  26662=>"010000101",
  26663=>"011101001",
  26664=>"000001101",
  26665=>"010001110",
  26666=>"110110011",
  26667=>"101110011",
  26668=>"111011100",
  26669=>"011010101",
  26670=>"101001010",
  26671=>"000110011",
  26672=>"110100101",
  26673=>"100110001",
  26674=>"101001011",
  26675=>"101100101",
  26676=>"101101101",
  26677=>"001000100",
  26678=>"010000001",
  26679=>"101001010",
  26680=>"010111011",
  26681=>"100000000",
  26682=>"011011101",
  26683=>"001000110",
  26684=>"011100000",
  26685=>"011111101",
  26686=>"001010100",
  26687=>"010001011",
  26688=>"100001011",
  26689=>"001111110",
  26690=>"111010000",
  26691=>"011101111",
  26692=>"110001010",
  26693=>"011000001",
  26694=>"001100000",
  26695=>"101001111",
  26696=>"101000111",
  26697=>"011000000",
  26698=>"001100101",
  26699=>"100010011",
  26700=>"011011101",
  26701=>"010000000",
  26702=>"011101010",
  26703=>"110000010",
  26704=>"101111101",
  26705=>"000110000",
  26706=>"000111000",
  26707=>"011001110",
  26708=>"000011100",
  26709=>"110000011",
  26710=>"010000101",
  26711=>"000011110",
  26712=>"111100111",
  26713=>"010010100",
  26714=>"011000011",
  26715=>"010000000",
  26716=>"110000100",
  26717=>"110000001",
  26718=>"000010001",
  26719=>"011001010",
  26720=>"110100111",
  26721=>"001101111",
  26722=>"011101001",
  26723=>"011000001",
  26724=>"101001100",
  26725=>"000100110",
  26726=>"001000110",
  26727=>"001000111",
  26728=>"101110010",
  26729=>"001101011",
  26730=>"100011001",
  26731=>"011010000",
  26732=>"001101000",
  26733=>"100101001",
  26734=>"101111110",
  26735=>"000011111",
  26736=>"111110110",
  26737=>"100000001",
  26738=>"101001000",
  26739=>"010101101",
  26740=>"010011100",
  26741=>"000000110",
  26742=>"100000010",
  26743=>"010110101",
  26744=>"010011101",
  26745=>"011111111",
  26746=>"111011110",
  26747=>"111100110",
  26748=>"110110001",
  26749=>"110110000",
  26750=>"111011001",
  26751=>"100011100",
  26752=>"110100011",
  26753=>"110101100",
  26754=>"001100011",
  26755=>"000101111",
  26756=>"111100100",
  26757=>"101000100",
  26758=>"101110010",
  26759=>"001101100",
  26760=>"000010001",
  26761=>"000000010",
  26762=>"001100101",
  26763=>"011011001",
  26764=>"101001011",
  26765=>"101010100",
  26766=>"010100000",
  26767=>"000011100",
  26768=>"111110111",
  26769=>"100110001",
  26770=>"011011111",
  26771=>"111111111",
  26772=>"000011110",
  26773=>"110001011",
  26774=>"100010001",
  26775=>"010110111",
  26776=>"111100111",
  26777=>"110000110",
  26778=>"101100111",
  26779=>"001110001",
  26780=>"110000011",
  26781=>"001100000",
  26782=>"110011111",
  26783=>"100000101",
  26784=>"110110001",
  26785=>"001111001",
  26786=>"001000010",
  26787=>"100101111",
  26788=>"101000000",
  26789=>"000011000",
  26790=>"000010111",
  26791=>"010000000",
  26792=>"111000001",
  26793=>"001100110",
  26794=>"000111100",
  26795=>"011111011",
  26796=>"001011010",
  26797=>"110001010",
  26798=>"010010101",
  26799=>"001110000",
  26800=>"001001101",
  26801=>"001001111",
  26802=>"011010110",
  26803=>"010011001",
  26804=>"100000101",
  26805=>"100001100",
  26806=>"001001101",
  26807=>"100110101",
  26808=>"011101000",
  26809=>"000011101",
  26810=>"011100100",
  26811=>"000110110",
  26812=>"111010101",
  26813=>"010010011",
  26814=>"010010100",
  26815=>"111000110",
  26816=>"011100100",
  26817=>"000111101",
  26818=>"110010010",
  26819=>"111110111",
  26820=>"111110011",
  26821=>"100101111",
  26822=>"001000010",
  26823=>"100011011",
  26824=>"010010000",
  26825=>"011010100",
  26826=>"110000010",
  26827=>"101111110",
  26828=>"001111110",
  26829=>"000010101",
  26830=>"101001010",
  26831=>"110000101",
  26832=>"010110000",
  26833=>"010011101",
  26834=>"100110110",
  26835=>"011000010",
  26836=>"101111010",
  26837=>"111001100",
  26838=>"000101000",
  26839=>"010100000",
  26840=>"010011000",
  26841=>"111001011",
  26842=>"000010001",
  26843=>"111111100",
  26844=>"000100000",
  26845=>"110000111",
  26846=>"010000000",
  26847=>"000011100",
  26848=>"001101111",
  26849=>"011011000",
  26850=>"101100011",
  26851=>"001010100",
  26852=>"011100100",
  26853=>"000001011",
  26854=>"010101100",
  26855=>"001111111",
  26856=>"001110000",
  26857=>"101110011",
  26858=>"001110011",
  26859=>"101111011",
  26860=>"010000000",
  26861=>"101000011",
  26862=>"001011100",
  26863=>"101011000",
  26864=>"100000111",
  26865=>"111111001",
  26866=>"111110100",
  26867=>"010111110",
  26868=>"101000011",
  26869=>"010100101",
  26870=>"101001111",
  26871=>"011001001",
  26872=>"011010001",
  26873=>"100000001",
  26874=>"011000110",
  26875=>"101100010",
  26876=>"101111111",
  26877=>"110000110",
  26878=>"011111000",
  26879=>"101000111",
  26880=>"001000111",
  26881=>"111110000",
  26882=>"110011010",
  26883=>"000111001",
  26884=>"111110000",
  26885=>"111111010",
  26886=>"011010000",
  26887=>"111110000",
  26888=>"111101110",
  26889=>"001000000",
  26890=>"111111000",
  26891=>"000111011",
  26892=>"011011000",
  26893=>"101010101",
  26894=>"000111100",
  26895=>"000011001",
  26896=>"101000101",
  26897=>"100111100",
  26898=>"100110111",
  26899=>"011010011",
  26900=>"010000001",
  26901=>"111101101",
  26902=>"010000000",
  26903=>"110011000",
  26904=>"100000011",
  26905=>"000110100",
  26906=>"000001101",
  26907=>"001010100",
  26908=>"000000100",
  26909=>"001100100",
  26910=>"111011001",
  26911=>"000100101",
  26912=>"001010000",
  26913=>"011100010",
  26914=>"110000011",
  26915=>"001110100",
  26916=>"101110001",
  26917=>"000101011",
  26918=>"110101000",
  26919=>"000010000",
  26920=>"111001011",
  26921=>"100100010",
  26922=>"110100110",
  26923=>"011000111",
  26924=>"111011011",
  26925=>"000100111",
  26926=>"100010001",
  26927=>"000010110",
  26928=>"001000100",
  26929=>"000101101",
  26930=>"100111101",
  26931=>"111101111",
  26932=>"100010010",
  26933=>"111011001",
  26934=>"101101111",
  26935=>"000101000",
  26936=>"001101010",
  26937=>"011110000",
  26938=>"110000101",
  26939=>"101110101",
  26940=>"001011100",
  26941=>"010110100",
  26942=>"001101101",
  26943=>"010001110",
  26944=>"111111001",
  26945=>"111110010",
  26946=>"000100101",
  26947=>"000100101",
  26948=>"001101000",
  26949=>"100010111",
  26950=>"000001100",
  26951=>"110011011",
  26952=>"100000000",
  26953=>"100000110",
  26954=>"111010010",
  26955=>"101001101",
  26956=>"010001010",
  26957=>"111111000",
  26958=>"010000000",
  26959=>"111100101",
  26960=>"011100001",
  26961=>"001011100",
  26962=>"000111111",
  26963=>"100001011",
  26964=>"001010101",
  26965=>"001011101",
  26966=>"110000100",
  26967=>"001110111",
  26968=>"111100101",
  26969=>"110001110",
  26970=>"100101100",
  26971=>"100100011",
  26972=>"011000101",
  26973=>"111101001",
  26974=>"010010100",
  26975=>"111111001",
  26976=>"110000101",
  26977=>"101000110",
  26978=>"110101110",
  26979=>"011110100",
  26980=>"010101111",
  26981=>"111110011",
  26982=>"110110001",
  26983=>"001011110",
  26984=>"000000000",
  26985=>"000111100",
  26986=>"001110101",
  26987=>"011101111",
  26988=>"011110111",
  26989=>"000101110",
  26990=>"101110111",
  26991=>"010001011",
  26992=>"110101000",
  26993=>"101001101",
  26994=>"101011110",
  26995=>"000000000",
  26996=>"110101000",
  26997=>"010011011",
  26998=>"101011010",
  26999=>"011111100",
  27000=>"110101000",
  27001=>"101011110",
  27002=>"001011100",
  27003=>"101110010",
  27004=>"111111111",
  27005=>"001000011",
  27006=>"100010100",
  27007=>"111000100",
  27008=>"010001010",
  27009=>"011010011",
  27010=>"000001100",
  27011=>"101111001",
  27012=>"010110111",
  27013=>"101000011",
  27014=>"000110000",
  27015=>"111110100",
  27016=>"010110000",
  27017=>"111000010",
  27018=>"001100010",
  27019=>"111111110",
  27020=>"100011011",
  27021=>"111100010",
  27022=>"100010100",
  27023=>"011000111",
  27024=>"111101001",
  27025=>"111111010",
  27026=>"011110000",
  27027=>"101111100",
  27028=>"110101101",
  27029=>"000110100",
  27030=>"000011010",
  27031=>"011010001",
  27032=>"011000100",
  27033=>"010111001",
  27034=>"100000110",
  27035=>"000100101",
  27036=>"001011001",
  27037=>"011100010",
  27038=>"101101000",
  27039=>"111001001",
  27040=>"110001000",
  27041=>"111001110",
  27042=>"110101110",
  27043=>"111010001",
  27044=>"110011110",
  27045=>"001001000",
  27046=>"111101010",
  27047=>"111011010",
  27048=>"111100110",
  27049=>"000010011",
  27050=>"010100111",
  27051=>"101010001",
  27052=>"000101010",
  27053=>"110001111",
  27054=>"111110000",
  27055=>"001110001",
  27056=>"110001011",
  27057=>"000010000",
  27058=>"110110011",
  27059=>"000111100",
  27060=>"010111111",
  27061=>"101000000",
  27062=>"010010011",
  27063=>"000101010",
  27064=>"110011011",
  27065=>"111101000",
  27066=>"010000011",
  27067=>"010100011",
  27068=>"100110010",
  27069=>"011100100",
  27070=>"000110011",
  27071=>"111001010",
  27072=>"000100010",
  27073=>"110111010",
  27074=>"000110001",
  27075=>"101011000",
  27076=>"010101000",
  27077=>"100000010",
  27078=>"110001111",
  27079=>"111100101",
  27080=>"010100011",
  27081=>"001111000",
  27082=>"001111110",
  27083=>"000011010",
  27084=>"011101001",
  27085=>"100100111",
  27086=>"011011110",
  27087=>"100100001",
  27088=>"011010110",
  27089=>"100111001",
  27090=>"011111000",
  27091=>"110100101",
  27092=>"110011000",
  27093=>"000110001",
  27094=>"010111001",
  27095=>"110010110",
  27096=>"100010011",
  27097=>"100111100",
  27098=>"001011100",
  27099=>"100111010",
  27100=>"001000001",
  27101=>"010101001",
  27102=>"001110011",
  27103=>"101100101",
  27104=>"011110001",
  27105=>"110100010",
  27106=>"010110111",
  27107=>"100011111",
  27108=>"011001011",
  27109=>"111111010",
  27110=>"010011010",
  27111=>"111000100",
  27112=>"110101101",
  27113=>"111111011",
  27114=>"011110011",
  27115=>"010001000",
  27116=>"000001001",
  27117=>"011111000",
  27118=>"110001000",
  27119=>"010001110",
  27120=>"110111111",
  27121=>"001101110",
  27122=>"101100011",
  27123=>"010010101",
  27124=>"000101110",
  27125=>"111111010",
  27126=>"100001011",
  27127=>"100110111",
  27128=>"010101001",
  27129=>"000001000",
  27130=>"011000011",
  27131=>"000110010",
  27132=>"110101001",
  27133=>"000001100",
  27134=>"010101011",
  27135=>"100100010",
  27136=>"111111100",
  27137=>"101000000",
  27138=>"110101111",
  27139=>"100000110",
  27140=>"010010001",
  27141=>"001100000",
  27142=>"010011011",
  27143=>"101011000",
  27144=>"110011000",
  27145=>"110000101",
  27146=>"011101001",
  27147=>"110010100",
  27148=>"001110010",
  27149=>"011110001",
  27150=>"010011001",
  27151=>"111100101",
  27152=>"001111010",
  27153=>"101000010",
  27154=>"011100001",
  27155=>"100100011",
  27156=>"010001110",
  27157=>"101100001",
  27158=>"010000010",
  27159=>"100100001",
  27160=>"000010111",
  27161=>"011000011",
  27162=>"100011000",
  27163=>"010011001",
  27164=>"110000110",
  27165=>"001111011",
  27166=>"100010110",
  27167=>"010000111",
  27168=>"110110111",
  27169=>"101111000",
  27170=>"011101110",
  27171=>"001011111",
  27172=>"110110100",
  27173=>"010110100",
  27174=>"001000000",
  27175=>"010111011",
  27176=>"000101000",
  27177=>"011110101",
  27178=>"011111101",
  27179=>"110010011",
  27180=>"011100000",
  27181=>"010011101",
  27182=>"000110000",
  27183=>"010011101",
  27184=>"000000101",
  27185=>"100000001",
  27186=>"101000010",
  27187=>"011010101",
  27188=>"001111100",
  27189=>"011101100",
  27190=>"001100011",
  27191=>"100000000",
  27192=>"100100001",
  27193=>"110100101",
  27194=>"000100110",
  27195=>"001011110",
  27196=>"110111110",
  27197=>"110111100",
  27198=>"100111000",
  27199=>"001011100",
  27200=>"101111000",
  27201=>"001001010",
  27202=>"101001110",
  27203=>"101111111",
  27204=>"010100000",
  27205=>"010110011",
  27206=>"011000010",
  27207=>"101011111",
  27208=>"000101000",
  27209=>"110101111",
  27210=>"111100010",
  27211=>"011101100",
  27212=>"100010001",
  27213=>"110101001",
  27214=>"101000100",
  27215=>"100011111",
  27216=>"000100011",
  27217=>"100101000",
  27218=>"101000000",
  27219=>"000100110",
  27220=>"000010001",
  27221=>"000011111",
  27222=>"100100000",
  27223=>"000100110",
  27224=>"011110000",
  27225=>"101110111",
  27226=>"011110100",
  27227=>"001000000",
  27228=>"101101110",
  27229=>"110111101",
  27230=>"100100011",
  27231=>"100010101",
  27232=>"111110010",
  27233=>"100110011",
  27234=>"101001000",
  27235=>"101001101",
  27236=>"010011001",
  27237=>"100101011",
  27238=>"000100111",
  27239=>"101000111",
  27240=>"110010100",
  27241=>"110100110",
  27242=>"001010101",
  27243=>"110100100",
  27244=>"011111100",
  27245=>"100001110",
  27246=>"100000101",
  27247=>"100100111",
  27248=>"010110111",
  27249=>"000000010",
  27250=>"001001000",
  27251=>"010011000",
  27252=>"001101100",
  27253=>"000000011",
  27254=>"001111111",
  27255=>"011111111",
  27256=>"100000011",
  27257=>"000001010",
  27258=>"000000010",
  27259=>"011011110",
  27260=>"100110000",
  27261=>"110110101",
  27262=>"101010100",
  27263=>"110110101",
  27264=>"000011111",
  27265=>"111111000",
  27266=>"100011010",
  27267=>"011001001",
  27268=>"111011000",
  27269=>"111111010",
  27270=>"100011011",
  27271=>"011111100",
  27272=>"001111110",
  27273=>"010110101",
  27274=>"101010000",
  27275=>"100100000",
  27276=>"110011011",
  27277=>"100100001",
  27278=>"010100010",
  27279=>"001111011",
  27280=>"000111101",
  27281=>"010011000",
  27282=>"000110110",
  27283=>"010010110",
  27284=>"001110001",
  27285=>"011010011",
  27286=>"110110111",
  27287=>"010000101",
  27288=>"001000010",
  27289=>"101011111",
  27290=>"010010000",
  27291=>"101101010",
  27292=>"101110111",
  27293=>"001010100",
  27294=>"011101001",
  27295=>"100101111",
  27296=>"100111100",
  27297=>"110011110",
  27298=>"000001101",
  27299=>"000011010",
  27300=>"001000110",
  27301=>"001100111",
  27302=>"111001101",
  27303=>"010011101",
  27304=>"101011101",
  27305=>"100011001",
  27306=>"100111011",
  27307=>"101101000",
  27308=>"101000000",
  27309=>"010010001",
  27310=>"001111110",
  27311=>"010111101",
  27312=>"110101000",
  27313=>"011001111",
  27314=>"100111011",
  27315=>"001111011",
  27316=>"110000100",
  27317=>"001010010",
  27318=>"001101111",
  27319=>"001010000",
  27320=>"011100100",
  27321=>"111011110",
  27322=>"110100001",
  27323=>"010100010",
  27324=>"101001001",
  27325=>"010010100",
  27326=>"101111101",
  27327=>"110001001",
  27328=>"111111111",
  27329=>"111001101",
  27330=>"010010101",
  27331=>"001010000",
  27332=>"110000111",
  27333=>"111001001",
  27334=>"011000100",
  27335=>"010000111",
  27336=>"000100100",
  27337=>"110010011",
  27338=>"010011100",
  27339=>"110000100",
  27340=>"101100010",
  27341=>"010001011",
  27342=>"001000110",
  27343=>"101000010",
  27344=>"001001100",
  27345=>"110110001",
  27346=>"110110100",
  27347=>"000110101",
  27348=>"010100100",
  27349=>"000100011",
  27350=>"100110011",
  27351=>"111001110",
  27352=>"111101101",
  27353=>"001010010",
  27354=>"011000101",
  27355=>"110100000",
  27356=>"011001001",
  27357=>"111111000",
  27358=>"100000001",
  27359=>"101001110",
  27360=>"110001111",
  27361=>"100110011",
  27362=>"000000011",
  27363=>"011001111",
  27364=>"101111111",
  27365=>"110101110",
  27366=>"001010000",
  27367=>"010010000",
  27368=>"100000111",
  27369=>"110101111",
  27370=>"011100110",
  27371=>"011011110",
  27372=>"010101000",
  27373=>"111001110",
  27374=>"011001110",
  27375=>"101000000",
  27376=>"011111110",
  27377=>"100101110",
  27378=>"111010110",
  27379=>"101011111",
  27380=>"101100001",
  27381=>"100011100",
  27382=>"011010000",
  27383=>"001011010",
  27384=>"110000000",
  27385=>"011110101",
  27386=>"011101010",
  27387=>"001000001",
  27388=>"111011100",
  27389=>"101101010",
  27390=>"100010100",
  27391=>"001000000",
  27392=>"010111001",
  27393=>"011011011",
  27394=>"101000101",
  27395=>"001001101",
  27396=>"011011110",
  27397=>"111001010",
  27398=>"111011010",
  27399=>"010101101",
  27400=>"010000110",
  27401=>"101110001",
  27402=>"001000101",
  27403=>"111011000",
  27404=>"010010101",
  27405=>"011000110",
  27406=>"000000100",
  27407=>"100100111",
  27408=>"010110110",
  27409=>"011000101",
  27410=>"101111010",
  27411=>"011010110",
  27412=>"111100111",
  27413=>"101011110",
  27414=>"110101110",
  27415=>"001011010",
  27416=>"011101001",
  27417=>"000010110",
  27418=>"001110010",
  27419=>"111101101",
  27420=>"010010100",
  27421=>"101100110",
  27422=>"111111111",
  27423=>"000011001",
  27424=>"100010011",
  27425=>"100110111",
  27426=>"000001000",
  27427=>"010111100",
  27428=>"001111101",
  27429=>"000010010",
  27430=>"000101101",
  27431=>"001101011",
  27432=>"000111010",
  27433=>"111111111",
  27434=>"000100011",
  27435=>"000111000",
  27436=>"111000001",
  27437=>"110111011",
  27438=>"011010000",
  27439=>"000000000",
  27440=>"011001001",
  27441=>"101111110",
  27442=>"110100110",
  27443=>"100001110",
  27444=>"101001110",
  27445=>"100000010",
  27446=>"011001100",
  27447=>"110000100",
  27448=>"100011011",
  27449=>"011001010",
  27450=>"001000000",
  27451=>"101111010",
  27452=>"110000100",
  27453=>"111110100",
  27454=>"001001000",
  27455=>"100010110",
  27456=>"111101100",
  27457=>"100000110",
  27458=>"111110001",
  27459=>"001000011",
  27460=>"010010100",
  27461=>"010000011",
  27462=>"011110100",
  27463=>"010010001",
  27464=>"101001011",
  27465=>"110011011",
  27466=>"110011101",
  27467=>"110101101",
  27468=>"111001011",
  27469=>"011110110",
  27470=>"111100000",
  27471=>"101111100",
  27472=>"001111000",
  27473=>"100101000",
  27474=>"000110110",
  27475=>"110101110",
  27476=>"101111100",
  27477=>"000010110",
  27478=>"011001101",
  27479=>"011011111",
  27480=>"100110001",
  27481=>"111010000",
  27482=>"111110011",
  27483=>"010111100",
  27484=>"010010111",
  27485=>"110011100",
  27486=>"110100011",
  27487=>"010001000",
  27488=>"100100111",
  27489=>"100100010",
  27490=>"000100100",
  27491=>"101011110",
  27492=>"101011110",
  27493=>"111010010",
  27494=>"011100010",
  27495=>"001101011",
  27496=>"001010101",
  27497=>"000010010",
  27498=>"010000111",
  27499=>"111111001",
  27500=>"011000101",
  27501=>"100110111",
  27502=>"010110000",
  27503=>"000000000",
  27504=>"000011111",
  27505=>"011100011",
  27506=>"000010001",
  27507=>"000011110",
  27508=>"111011101",
  27509=>"101111011",
  27510=>"111100000",
  27511=>"000111110",
  27512=>"001111000",
  27513=>"110101100",
  27514=>"101011000",
  27515=>"101000111",
  27516=>"100001010",
  27517=>"000011110",
  27518=>"001101100",
  27519=>"101110110",
  27520=>"001100000",
  27521=>"000110110",
  27522=>"011001010",
  27523=>"001111000",
  27524=>"111111100",
  27525=>"010001011",
  27526=>"111001111",
  27527=>"100110010",
  27528=>"111010001",
  27529=>"101001001",
  27530=>"110001100",
  27531=>"111000000",
  27532=>"100001011",
  27533=>"010110000",
  27534=>"101000101",
  27535=>"010011010",
  27536=>"001101000",
  27537=>"001101101",
  27538=>"111001110",
  27539=>"001010001",
  27540=>"110000000",
  27541=>"110100110",
  27542=>"010001000",
  27543=>"101001110",
  27544=>"000010101",
  27545=>"100000010",
  27546=>"000011001",
  27547=>"110110010",
  27548=>"011101000",
  27549=>"011010001",
  27550=>"110101001",
  27551=>"111100100",
  27552=>"101110100",
  27553=>"111110111",
  27554=>"111000101",
  27555=>"100001011",
  27556=>"101010101",
  27557=>"010101111",
  27558=>"001101111",
  27559=>"010110101",
  27560=>"000101010",
  27561=>"111101100",
  27562=>"011111110",
  27563=>"001010001",
  27564=>"100101100",
  27565=>"111110111",
  27566=>"000101110",
  27567=>"011110101",
  27568=>"110001101",
  27569=>"010101000",
  27570=>"011010111",
  27571=>"111010111",
  27572=>"111011110",
  27573=>"000000010",
  27574=>"101101010",
  27575=>"011000001",
  27576=>"011001000",
  27577=>"011100101",
  27578=>"001110100",
  27579=>"101101101",
  27580=>"110101000",
  27581=>"111111101",
  27582=>"001100000",
  27583=>"110000101",
  27584=>"011111010",
  27585=>"001010101",
  27586=>"111001110",
  27587=>"000000001",
  27588=>"111000001",
  27589=>"100001101",
  27590=>"101111010",
  27591=>"010011101",
  27592=>"000010000",
  27593=>"101010111",
  27594=>"011001110",
  27595=>"010011111",
  27596=>"011110011",
  27597=>"111011101",
  27598=>"011100110",
  27599=>"101011000",
  27600=>"010001111",
  27601=>"000011100",
  27602=>"010001010",
  27603=>"110001100",
  27604=>"010000001",
  27605=>"100000110",
  27606=>"011011111",
  27607=>"101111100",
  27608=>"001000111",
  27609=>"000001111",
  27610=>"101011010",
  27611=>"001011100",
  27612=>"100000101",
  27613=>"000011101",
  27614=>"100100111",
  27615=>"001011101",
  27616=>"111100100",
  27617=>"100010011",
  27618=>"011100110",
  27619=>"000000010",
  27620=>"010011111",
  27621=>"111100100",
  27622=>"111100000",
  27623=>"000111100",
  27624=>"011011001",
  27625=>"011111111",
  27626=>"111100011",
  27627=>"011111010",
  27628=>"101100011",
  27629=>"110101100",
  27630=>"100101110",
  27631=>"110111001",
  27632=>"010011000",
  27633=>"010000100",
  27634=>"011111111",
  27635=>"101011000",
  27636=>"000000011",
  27637=>"101101110",
  27638=>"110001001",
  27639=>"000000110",
  27640=>"101110111",
  27641=>"010100111",
  27642=>"111000101",
  27643=>"110011010",
  27644=>"001110000",
  27645=>"110001000",
  27646=>"111101101",
  27647=>"100101100",
  27648=>"000111110",
  27649=>"001011011",
  27650=>"110000101",
  27651=>"011100101",
  27652=>"111111000",
  27653=>"000001010",
  27654=>"000010000",
  27655=>"001001111",
  27656=>"101100010",
  27657=>"110100110",
  27658=>"010001111",
  27659=>"111000001",
  27660=>"000100110",
  27661=>"011011100",
  27662=>"101011001",
  27663=>"111010110",
  27664=>"110000000",
  27665=>"000110100",
  27666=>"110101111",
  27667=>"101100011",
  27668=>"011010111",
  27669=>"111010101",
  27670=>"110011001",
  27671=>"110010101",
  27672=>"110011111",
  27673=>"111001110",
  27674=>"011000100",
  27675=>"000000110",
  27676=>"100001011",
  27677=>"110011110",
  27678=>"000110011",
  27679=>"110101011",
  27680=>"111111111",
  27681=>"110100011",
  27682=>"101010011",
  27683=>"111010100",
  27684=>"110010100",
  27685=>"010100100",
  27686=>"101100000",
  27687=>"000100111",
  27688=>"110011010",
  27689=>"000110010",
  27690=>"011000011",
  27691=>"110010111",
  27692=>"100111111",
  27693=>"010111101",
  27694=>"000110001",
  27695=>"000011110",
  27696=>"011101101",
  27697=>"111000110",
  27698=>"101101011",
  27699=>"100100100",
  27700=>"010000010",
  27701=>"010110000",
  27702=>"001110010",
  27703=>"001100010",
  27704=>"001111000",
  27705=>"110101101",
  27706=>"100010110",
  27707=>"000000011",
  27708=>"100110010",
  27709=>"100011001",
  27710=>"011101010",
  27711=>"000110010",
  27712=>"011100000",
  27713=>"110000001",
  27714=>"101111011",
  27715=>"010001000",
  27716=>"101001110",
  27717=>"110100000",
  27718=>"010110100",
  27719=>"100110111",
  27720=>"000101001",
  27721=>"110111011",
  27722=>"000110110",
  27723=>"111101010",
  27724=>"000111101",
  27725=>"011010001",
  27726=>"111000000",
  27727=>"000000010",
  27728=>"001011011",
  27729=>"011111101",
  27730=>"111011001",
  27731=>"011100100",
  27732=>"000001100",
  27733=>"011010010",
  27734=>"111100110",
  27735=>"101011010",
  27736=>"111111110",
  27737=>"010110010",
  27738=>"100001110",
  27739=>"010100001",
  27740=>"110000010",
  27741=>"000101000",
  27742=>"101110111",
  27743=>"001111001",
  27744=>"111100110",
  27745=>"101111011",
  27746=>"000011000",
  27747=>"100100010",
  27748=>"110000101",
  27749=>"101010111",
  27750=>"000101011",
  27751=>"111101100",
  27752=>"010011100",
  27753=>"110000100",
  27754=>"000011111",
  27755=>"000001110",
  27756=>"001011001",
  27757=>"000100100",
  27758=>"101000011",
  27759=>"000111110",
  27760=>"001000000",
  27761=>"001111000",
  27762=>"111000111",
  27763=>"000111110",
  27764=>"010101010",
  27765=>"001000001",
  27766=>"100101010",
  27767=>"110101101",
  27768=>"111001011",
  27769=>"110010101",
  27770=>"101010010",
  27771=>"110101001",
  27772=>"010000100",
  27773=>"100111011",
  27774=>"010111111",
  27775=>"010111110",
  27776=>"100100000",
  27777=>"101001110",
  27778=>"001000101",
  27779=>"111110111",
  27780=>"101010001",
  27781=>"101011100",
  27782=>"101110011",
  27783=>"101001000",
  27784=>"001001100",
  27785=>"101111111",
  27786=>"110001111",
  27787=>"010101001",
  27788=>"000100100",
  27789=>"001100001",
  27790=>"101001001",
  27791=>"010101001",
  27792=>"000011001",
  27793=>"010100111",
  27794=>"101001101",
  27795=>"001000000",
  27796=>"000111101",
  27797=>"000101001",
  27798=>"001010000",
  27799=>"111010011",
  27800=>"110111000",
  27801=>"001111111",
  27802=>"101001101",
  27803=>"001000011",
  27804=>"000001100",
  27805=>"111010011",
  27806=>"111101110",
  27807=>"111101010",
  27808=>"100100101",
  27809=>"110010101",
  27810=>"111001111",
  27811=>"111111010",
  27812=>"000110101",
  27813=>"101000001",
  27814=>"101011110",
  27815=>"111110111",
  27816=>"000110101",
  27817=>"001011101",
  27818=>"000110000",
  27819=>"100100110",
  27820=>"000101101",
  27821=>"000000101",
  27822=>"011101111",
  27823=>"111001110",
  27824=>"001001010",
  27825=>"011110000",
  27826=>"001110000",
  27827=>"010001011",
  27828=>"111001111",
  27829=>"010110000",
  27830=>"010100111",
  27831=>"110000110",
  27832=>"110111000",
  27833=>"001011011",
  27834=>"000001110",
  27835=>"101011100",
  27836=>"001010000",
  27837=>"101000110",
  27838=>"001100001",
  27839=>"001010101",
  27840=>"001001111",
  27841=>"000000011",
  27842=>"001100111",
  27843=>"110100110",
  27844=>"001111000",
  27845=>"000001100",
  27846=>"100101110",
  27847=>"000101100",
  27848=>"000110001",
  27849=>"010000000",
  27850=>"001000000",
  27851=>"011100000",
  27852=>"110110101",
  27853=>"111010001",
  27854=>"001111110",
  27855=>"010010101",
  27856=>"110111010",
  27857=>"110011001",
  27858=>"100100011",
  27859=>"001001110",
  27860=>"001010101",
  27861=>"000001101",
  27862=>"101010000",
  27863=>"111111001",
  27864=>"111100000",
  27865=>"101111001",
  27866=>"001000000",
  27867=>"010000110",
  27868=>"011011111",
  27869=>"000001000",
  27870=>"010101010",
  27871=>"010111011",
  27872=>"000010010",
  27873=>"010010111",
  27874=>"110101100",
  27875=>"110100000",
  27876=>"110110000",
  27877=>"010111110",
  27878=>"000101100",
  27879=>"000110101",
  27880=>"110011000",
  27881=>"000111100",
  27882=>"100100000",
  27883=>"010011000",
  27884=>"010100110",
  27885=>"000000100",
  27886=>"010110110",
  27887=>"010110010",
  27888=>"001011111",
  27889=>"010111100",
  27890=>"011011111",
  27891=>"100011011",
  27892=>"111100101",
  27893=>"111101101",
  27894=>"000011101",
  27895=>"001101100",
  27896=>"000110100",
  27897=>"010100010",
  27898=>"101101101",
  27899=>"001100101",
  27900=>"110010111",
  27901=>"010101011",
  27902=>"000010100",
  27903=>"100010000",
  27904=>"011010111",
  27905=>"010011010",
  27906=>"001001101",
  27907=>"011011111",
  27908=>"001010110",
  27909=>"111011110",
  27910=>"100011001",
  27911=>"101111101",
  27912=>"100011001",
  27913=>"100110001",
  27914=>"100011101",
  27915=>"110010100",
  27916=>"101011000",
  27917=>"100101010",
  27918=>"100000110",
  27919=>"100111100",
  27920=>"011001101",
  27921=>"000011110",
  27922=>"001110011",
  27923=>"101000111",
  27924=>"001010100",
  27925=>"001111001",
  27926=>"011001000",
  27927=>"001000010",
  27928=>"011101010",
  27929=>"110100000",
  27930=>"100010101",
  27931=>"001010100",
  27932=>"001001111",
  27933=>"100001000",
  27934=>"110011000",
  27935=>"010101110",
  27936=>"010010010",
  27937=>"100100001",
  27938=>"101010101",
  27939=>"010100101",
  27940=>"000101000",
  27941=>"100001000",
  27942=>"101111101",
  27943=>"100011101",
  27944=>"111111111",
  27945=>"010110101",
  27946=>"000000011",
  27947=>"110101000",
  27948=>"110110111",
  27949=>"010110100",
  27950=>"001100011",
  27951=>"101001111",
  27952=>"110110100",
  27953=>"100101101",
  27954=>"111001001",
  27955=>"001110010",
  27956=>"000011110",
  27957=>"010001111",
  27958=>"000000110",
  27959=>"000001111",
  27960=>"101110011",
  27961=>"000000010",
  27962=>"110110000",
  27963=>"111001100",
  27964=>"001111110",
  27965=>"011100110",
  27966=>"001110101",
  27967=>"101100110",
  27968=>"011001010",
  27969=>"110110101",
  27970=>"101011111",
  27971=>"001001011",
  27972=>"110101100",
  27973=>"100111000",
  27974=>"001110100",
  27975=>"000000011",
  27976=>"010100010",
  27977=>"101101101",
  27978=>"111000100",
  27979=>"110101111",
  27980=>"101111011",
  27981=>"001001111",
  27982=>"000100100",
  27983=>"000010010",
  27984=>"101011011",
  27985=>"111110101",
  27986=>"001011111",
  27987=>"011010001",
  27988=>"110100010",
  27989=>"011011001",
  27990=>"101100010",
  27991=>"000001110",
  27992=>"101001101",
  27993=>"000001010",
  27994=>"000010111",
  27995=>"001000010",
  27996=>"000011011",
  27997=>"001010011",
  27998=>"110011100",
  27999=>"101010011",
  28000=>"101100110",
  28001=>"100011110",
  28002=>"111010110",
  28003=>"000100100",
  28004=>"011000011",
  28005=>"111000100",
  28006=>"000000010",
  28007=>"110110100",
  28008=>"111101011",
  28009=>"110000000",
  28010=>"010101001",
  28011=>"000111010",
  28012=>"110111111",
  28013=>"110001011",
  28014=>"001100001",
  28015=>"101000000",
  28016=>"001001001",
  28017=>"101101101",
  28018=>"110100001",
  28019=>"110110111",
  28020=>"001100111",
  28021=>"111100101",
  28022=>"001000000",
  28023=>"110000000",
  28024=>"010110100",
  28025=>"000111111",
  28026=>"000001110",
  28027=>"100001100",
  28028=>"101000101",
  28029=>"011010011",
  28030=>"000000111",
  28031=>"010111110",
  28032=>"110111000",
  28033=>"010111001",
  28034=>"101100100",
  28035=>"100111111",
  28036=>"011000000",
  28037=>"011001100",
  28038=>"001110100",
  28039=>"111101101",
  28040=>"110000100",
  28041=>"110001000",
  28042=>"000110000",
  28043=>"101101001",
  28044=>"001101000",
  28045=>"110001000",
  28046=>"111101101",
  28047=>"000000100",
  28048=>"101101001",
  28049=>"110110110",
  28050=>"000011010",
  28051=>"000100011",
  28052=>"100010011",
  28053=>"000100110",
  28054=>"011000010",
  28055=>"100010110",
  28056=>"111111011",
  28057=>"101101101",
  28058=>"110111111",
  28059=>"111110101",
  28060=>"101011111",
  28061=>"001100001",
  28062=>"001111110",
  28063=>"111101011",
  28064=>"010000010",
  28065=>"100101111",
  28066=>"000000011",
  28067=>"110101001",
  28068=>"101101011",
  28069=>"011110000",
  28070=>"111101010",
  28071=>"110111010",
  28072=>"100101011",
  28073=>"010101000",
  28074=>"000100111",
  28075=>"100000011",
  28076=>"000000000",
  28077=>"001001001",
  28078=>"011011001",
  28079=>"101011100",
  28080=>"111011100",
  28081=>"111010010",
  28082=>"111111110",
  28083=>"010011111",
  28084=>"110001110",
  28085=>"010111000",
  28086=>"100011010",
  28087=>"010001011",
  28088=>"110000010",
  28089=>"001011101",
  28090=>"111011011",
  28091=>"001011111",
  28092=>"101010111",
  28093=>"100111010",
  28094=>"100000100",
  28095=>"000001000",
  28096=>"011010001",
  28097=>"111000111",
  28098=>"000100100",
  28099=>"111110010",
  28100=>"111110000",
  28101=>"011101110",
  28102=>"011111011",
  28103=>"110000010",
  28104=>"101011100",
  28105=>"100111001",
  28106=>"000111010",
  28107=>"111010111",
  28108=>"001010001",
  28109=>"110010000",
  28110=>"000001100",
  28111=>"101010010",
  28112=>"010000011",
  28113=>"100001001",
  28114=>"010000001",
  28115=>"000111011",
  28116=>"010011010",
  28117=>"110111101",
  28118=>"111000110",
  28119=>"110100001",
  28120=>"111100010",
  28121=>"101010110",
  28122=>"000011011",
  28123=>"100011111",
  28124=>"110011100",
  28125=>"000101101",
  28126=>"101101101",
  28127=>"101101000",
  28128=>"100110001",
  28129=>"101100011",
  28130=>"011001100",
  28131=>"001111001",
  28132=>"110000001",
  28133=>"001111110",
  28134=>"100110001",
  28135=>"010110101",
  28136=>"110001111",
  28137=>"011011001",
  28138=>"110110011",
  28139=>"110101001",
  28140=>"101111010",
  28141=>"010000001",
  28142=>"001010000",
  28143=>"111011000",
  28144=>"110101001",
  28145=>"011010110",
  28146=>"011110001",
  28147=>"110010000",
  28148=>"001010011",
  28149=>"011001110",
  28150=>"111010111",
  28151=>"110001110",
  28152=>"110111000",
  28153=>"111101111",
  28154=>"000100011",
  28155=>"100101111",
  28156=>"111100101",
  28157=>"011000011",
  28158=>"100011001",
  28159=>"000001100",
  28160=>"111001001",
  28161=>"111001010",
  28162=>"111001011",
  28163=>"001011100",
  28164=>"000011100",
  28165=>"011101000",
  28166=>"100101110",
  28167=>"111100100",
  28168=>"110001011",
  28169=>"111110011",
  28170=>"010101010",
  28171=>"010110100",
  28172=>"100010010",
  28173=>"001001011",
  28174=>"011001110",
  28175=>"111011001",
  28176=>"111101101",
  28177=>"011011111",
  28178=>"101001000",
  28179=>"110100010",
  28180=>"100100001",
  28181=>"101100000",
  28182=>"000001011",
  28183=>"011011110",
  28184=>"100001011",
  28185=>"000011101",
  28186=>"001101011",
  28187=>"000010101",
  28188=>"010011000",
  28189=>"101110010",
  28190=>"101000101",
  28191=>"010101101",
  28192=>"101000110",
  28193=>"101001011",
  28194=>"000011101",
  28195=>"100010000",
  28196=>"000001001",
  28197=>"111100101",
  28198=>"111100110",
  28199=>"011101111",
  28200=>"010011001",
  28201=>"100010001",
  28202=>"100100100",
  28203=>"010111011",
  28204=>"101101001",
  28205=>"011101011",
  28206=>"111000111",
  28207=>"100011111",
  28208=>"111001010",
  28209=>"001001001",
  28210=>"011101101",
  28211=>"000100110",
  28212=>"111100110",
  28213=>"011111000",
  28214=>"101010101",
  28215=>"101101111",
  28216=>"000111001",
  28217=>"010010000",
  28218=>"011011101",
  28219=>"101100101",
  28220=>"110110101",
  28221=>"000010111",
  28222=>"100100010",
  28223=>"001000010",
  28224=>"010010011",
  28225=>"000000010",
  28226=>"010001101",
  28227=>"001000001",
  28228=>"000010000",
  28229=>"101001010",
  28230=>"001000110",
  28231=>"001011111",
  28232=>"001000011",
  28233=>"000000101",
  28234=>"101001100",
  28235=>"000001110",
  28236=>"111001000",
  28237=>"100101001",
  28238=>"010111110",
  28239=>"011001001",
  28240=>"010000100",
  28241=>"011011100",
  28242=>"010111011",
  28243=>"001001110",
  28244=>"010101111",
  28245=>"000111100",
  28246=>"000110100",
  28247=>"111111101",
  28248=>"100010101",
  28249=>"011110011",
  28250=>"100101010",
  28251=>"011000010",
  28252=>"000011110",
  28253=>"010000001",
  28254=>"111000001",
  28255=>"100111011",
  28256=>"010111110",
  28257=>"110010000",
  28258=>"001110011",
  28259=>"111011100",
  28260=>"001000110",
  28261=>"010011111",
  28262=>"011110100",
  28263=>"111001011",
  28264=>"100000010",
  28265=>"011011111",
  28266=>"010000010",
  28267=>"001000100",
  28268=>"111101101",
  28269=>"010110001",
  28270=>"010010011",
  28271=>"101110100",
  28272=>"110000110",
  28273=>"001100101",
  28274=>"011101000",
  28275=>"101010100",
  28276=>"100000000",
  28277=>"001001000",
  28278=>"110011111",
  28279=>"011111110",
  28280=>"010000001",
  28281=>"111110010",
  28282=>"110011000",
  28283=>"110011000",
  28284=>"101000000",
  28285=>"011001010",
  28286=>"110011010",
  28287=>"001010101",
  28288=>"001000111",
  28289=>"111111111",
  28290=>"010011011",
  28291=>"010001011",
  28292=>"011000111",
  28293=>"001110010",
  28294=>"110001011",
  28295=>"101110001",
  28296=>"111001101",
  28297=>"000000000",
  28298=>"000110001",
  28299=>"110000110",
  28300=>"001110011",
  28301=>"101001111",
  28302=>"100101100",
  28303=>"101000100",
  28304=>"110101011",
  28305=>"011100100",
  28306=>"101101100",
  28307=>"101000110",
  28308=>"000101110",
  28309=>"110101001",
  28310=>"010010110",
  28311=>"000100000",
  28312=>"100011110",
  28313=>"001100101",
  28314=>"111011010",
  28315=>"111111010",
  28316=>"000000000",
  28317=>"000000110",
  28318=>"111101100",
  28319=>"000011100",
  28320=>"101111011",
  28321=>"110000001",
  28322=>"111101011",
  28323=>"110111000",
  28324=>"010011011",
  28325=>"111010010",
  28326=>"111100001",
  28327=>"100111110",
  28328=>"100010111",
  28329=>"000111010",
  28330=>"010001100",
  28331=>"001110101",
  28332=>"111001101",
  28333=>"000000111",
  28334=>"000111100",
  28335=>"110110001",
  28336=>"011010110",
  28337=>"101110101",
  28338=>"001101011",
  28339=>"101010010",
  28340=>"001101111",
  28341=>"110100111",
  28342=>"000111000",
  28343=>"111000000",
  28344=>"011101111",
  28345=>"001111001",
  28346=>"110010000",
  28347=>"000010000",
  28348=>"001111001",
  28349=>"001001001",
  28350=>"000111000",
  28351=>"011110011",
  28352=>"000101101",
  28353=>"110101111",
  28354=>"011101111",
  28355=>"001101111",
  28356=>"000011101",
  28357=>"101011010",
  28358=>"001111110",
  28359=>"001110100",
  28360=>"101000010",
  28361=>"001001000",
  28362=>"011001001",
  28363=>"000010100",
  28364=>"010110101",
  28365=>"000001100",
  28366=>"101110111",
  28367=>"010011011",
  28368=>"001011001",
  28369=>"010011000",
  28370=>"000010011",
  28371=>"000111011",
  28372=>"101101110",
  28373=>"001010101",
  28374=>"111011101",
  28375=>"001101110",
  28376=>"010001010",
  28377=>"000101000",
  28378=>"010101001",
  28379=>"011010001",
  28380=>"100001101",
  28381=>"100011100",
  28382=>"010010001",
  28383=>"111010110",
  28384=>"010101100",
  28385=>"101011100",
  28386=>"101110010",
  28387=>"000111010",
  28388=>"011110111",
  28389=>"100010000",
  28390=>"111000000",
  28391=>"011100000",
  28392=>"111110110",
  28393=>"111101110",
  28394=>"001010011",
  28395=>"111111100",
  28396=>"110110000",
  28397=>"010010101",
  28398=>"001110010",
  28399=>"001000000",
  28400=>"110111100",
  28401=>"011001011",
  28402=>"001001001",
  28403=>"011101000",
  28404=>"111001101",
  28405=>"111111100",
  28406=>"001010011",
  28407=>"110001110",
  28408=>"111001001",
  28409=>"101111010",
  28410=>"010111110",
  28411=>"110011100",
  28412=>"000011111",
  28413=>"101001100",
  28414=>"100000001",
  28415=>"111101011",
  28416=>"100101010",
  28417=>"000001000",
  28418=>"000010111",
  28419=>"110011100",
  28420=>"111100100",
  28421=>"000011101",
  28422=>"010110001",
  28423=>"000011110",
  28424=>"000101111",
  28425=>"111011101",
  28426=>"110111011",
  28427=>"010010000",
  28428=>"001000001",
  28429=>"000101011",
  28430=>"100000000",
  28431=>"111100100",
  28432=>"011011011",
  28433=>"011101011",
  28434=>"001101001",
  28435=>"011100000",
  28436=>"110111110",
  28437=>"000111111",
  28438=>"011011001",
  28439=>"110101100",
  28440=>"000010010",
  28441=>"100011101",
  28442=>"010011010",
  28443=>"110011111",
  28444=>"010011101",
  28445=>"011000000",
  28446=>"110011000",
  28447=>"011111000",
  28448=>"111101001",
  28449=>"110111111",
  28450=>"011101000",
  28451=>"000000000",
  28452=>"110000101",
  28453=>"100010101",
  28454=>"011000110",
  28455=>"011011101",
  28456=>"010000101",
  28457=>"000100110",
  28458=>"110111000",
  28459=>"100100111",
  28460=>"111111001",
  28461=>"011111101",
  28462=>"100010100",
  28463=>"101100110",
  28464=>"101101000",
  28465=>"011101011",
  28466=>"100001010",
  28467=>"110000010",
  28468=>"101001000",
  28469=>"001010110",
  28470=>"000010000",
  28471=>"000011101",
  28472=>"010110010",
  28473=>"100000110",
  28474=>"100010100",
  28475=>"010001001",
  28476=>"111000010",
  28477=>"001100010",
  28478=>"000010111",
  28479=>"101010001",
  28480=>"001000000",
  28481=>"100101110",
  28482=>"110000110",
  28483=>"010101010",
  28484=>"100111010",
  28485=>"100011010",
  28486=>"010111010",
  28487=>"100011010",
  28488=>"010001010",
  28489=>"110101101",
  28490=>"100101000",
  28491=>"111111010",
  28492=>"101011000",
  28493=>"100111000",
  28494=>"110001101",
  28495=>"101100101",
  28496=>"000000111",
  28497=>"100100100",
  28498=>"111111001",
  28499=>"000100111",
  28500=>"011001111",
  28501=>"111011110",
  28502=>"110101110",
  28503=>"110001101",
  28504=>"110111110",
  28505=>"111111001",
  28506=>"101011011",
  28507=>"111001110",
  28508=>"101111110",
  28509=>"010010100",
  28510=>"111000010",
  28511=>"000101010",
  28512=>"010000000",
  28513=>"000011101",
  28514=>"100010000",
  28515=>"100011010",
  28516=>"100101011",
  28517=>"001010101",
  28518=>"101110000",
  28519=>"111100001",
  28520=>"000010110",
  28521=>"000111111",
  28522=>"000000101",
  28523=>"001110111",
  28524=>"110110000",
  28525=>"100100100",
  28526=>"110011000",
  28527=>"000001100",
  28528=>"101011101",
  28529=>"010010010",
  28530=>"101111011",
  28531=>"101001011",
  28532=>"001001010",
  28533=>"010010111",
  28534=>"111111000",
  28535=>"001100101",
  28536=>"110010000",
  28537=>"110010100",
  28538=>"100110011",
  28539=>"110100101",
  28540=>"000100001",
  28541=>"001010101",
  28542=>"010000000",
  28543=>"101110100",
  28544=>"101011010",
  28545=>"011011010",
  28546=>"000110000",
  28547=>"100001110",
  28548=>"110001101",
  28549=>"100011101",
  28550=>"000001101",
  28551=>"000100100",
  28552=>"111001111",
  28553=>"110000100",
  28554=>"101100010",
  28555=>"010110011",
  28556=>"000100110",
  28557=>"111001110",
  28558=>"100011000",
  28559=>"101000100",
  28560=>"010011011",
  28561=>"111111110",
  28562=>"100101111",
  28563=>"001101101",
  28564=>"000010110",
  28565=>"110111011",
  28566=>"100101100",
  28567=>"110000100",
  28568=>"101011011",
  28569=>"000000111",
  28570=>"011001001",
  28571=>"010000000",
  28572=>"010000110",
  28573=>"110111110",
  28574=>"100111111",
  28575=>"000001100",
  28576=>"001000111",
  28577=>"111101111",
  28578=>"110000001",
  28579=>"000000010",
  28580=>"110001000",
  28581=>"000110000",
  28582=>"101000001",
  28583=>"111100111",
  28584=>"101001101",
  28585=>"101011010",
  28586=>"001100100",
  28587=>"100100111",
  28588=>"001010101",
  28589=>"101111110",
  28590=>"100010001",
  28591=>"111001101",
  28592=>"100110111",
  28593=>"000100010",
  28594=>"011011011",
  28595=>"111100101",
  28596=>"011000010",
  28597=>"111101100",
  28598=>"000101100",
  28599=>"100111010",
  28600=>"011110110",
  28601=>"001100000",
  28602=>"111101000",
  28603=>"010000111",
  28604=>"000111011",
  28605=>"111011110",
  28606=>"110010010",
  28607=>"001010100",
  28608=>"000011001",
  28609=>"100011101",
  28610=>"100111110",
  28611=>"001011010",
  28612=>"000100000",
  28613=>"100010111",
  28614=>"001100011",
  28615=>"111000100",
  28616=>"001101011",
  28617=>"000010011",
  28618=>"010010010",
  28619=>"000110001",
  28620=>"110011000",
  28621=>"101111111",
  28622=>"110100010",
  28623=>"100010101",
  28624=>"011110101",
  28625=>"010010110",
  28626=>"111001011",
  28627=>"000010001",
  28628=>"000101011",
  28629=>"000001000",
  28630=>"011000110",
  28631=>"101110111",
  28632=>"110111100",
  28633=>"101101110",
  28634=>"101100111",
  28635=>"111010000",
  28636=>"000110011",
  28637=>"110101111",
  28638=>"111101010",
  28639=>"101110110",
  28640=>"001010010",
  28641=>"010110100",
  28642=>"010010011",
  28643=>"111111111",
  28644=>"001100001",
  28645=>"010110100",
  28646=>"111100001",
  28647=>"011000101",
  28648=>"111111011",
  28649=>"101000011",
  28650=>"001001000",
  28651=>"000101110",
  28652=>"111000010",
  28653=>"110000001",
  28654=>"010010110",
  28655=>"111011010",
  28656=>"010100110",
  28657=>"011100100",
  28658=>"100000011",
  28659=>"111011011",
  28660=>"011110100",
  28661=>"011101110",
  28662=>"010111110",
  28663=>"001011110",
  28664=>"001100111",
  28665=>"000011110",
  28666=>"100110111",
  28667=>"110110111",
  28668=>"001010010",
  28669=>"101000001",
  28670=>"011000101",
  28671=>"101001101",
  28672=>"011001011",
  28673=>"001011100",
  28674=>"101111001",
  28675=>"000101000",
  28676=>"110110110",
  28677=>"000000001",
  28678=>"110110000",
  28679=>"011100101",
  28680=>"011000101",
  28681=>"000100110",
  28682=>"000100010",
  28683=>"011011100",
  28684=>"100000110",
  28685=>"010000010",
  28686=>"000111111",
  28687=>"000100110",
  28688=>"011000100",
  28689=>"100000100",
  28690=>"001010101",
  28691=>"100001110",
  28692=>"000100011",
  28693=>"100011000",
  28694=>"111011111",
  28695=>"111010100",
  28696=>"111111101",
  28697=>"001001100",
  28698=>"001010010",
  28699=>"011100011",
  28700=>"100001000",
  28701=>"100110110",
  28702=>"010101010",
  28703=>"001111000",
  28704=>"001010111",
  28705=>"110111001",
  28706=>"100111100",
  28707=>"110101000",
  28708=>"100111111",
  28709=>"010110010",
  28710=>"100111011",
  28711=>"101001011",
  28712=>"111011111",
  28713=>"010100000",
  28714=>"001010010",
  28715=>"101010001",
  28716=>"100010101",
  28717=>"111100111",
  28718=>"101101111",
  28719=>"010110001",
  28720=>"000111100",
  28721=>"100110001",
  28722=>"000110110",
  28723=>"111101110",
  28724=>"001101101",
  28725=>"110111011",
  28726=>"010010000",
  28727=>"100011001",
  28728=>"000001011",
  28729=>"001000111",
  28730=>"000011101",
  28731=>"010100100",
  28732=>"110100101",
  28733=>"101101111",
  28734=>"101001000",
  28735=>"000101110",
  28736=>"001011011",
  28737=>"101000101",
  28738=>"011010110",
  28739=>"011100110",
  28740=>"011010101",
  28741=>"111000000",
  28742=>"001011001",
  28743=>"000101111",
  28744=>"110001011",
  28745=>"100000011",
  28746=>"000011001",
  28747=>"001010001",
  28748=>"110100010",
  28749=>"110010111",
  28750=>"100010010",
  28751=>"111010010",
  28752=>"001111000",
  28753=>"010001100",
  28754=>"000110010",
  28755=>"111101101",
  28756=>"101011000",
  28757=>"101101000",
  28758=>"010001000",
  28759=>"001101101",
  28760=>"010010010",
  28761=>"110001010",
  28762=>"011000110",
  28763=>"100110101",
  28764=>"001000011",
  28765=>"000110000",
  28766=>"000101011",
  28767=>"000001110",
  28768=>"000010100",
  28769=>"010110100",
  28770=>"111111110",
  28771=>"010000100",
  28772=>"100000010",
  28773=>"001100101",
  28774=>"111100101",
  28775=>"011011111",
  28776=>"000011101",
  28777=>"110100010",
  28778=>"010000101",
  28779=>"101100011",
  28780=>"110111101",
  28781=>"011000000",
  28782=>"101011000",
  28783=>"111111111",
  28784=>"001000110",
  28785=>"101110001",
  28786=>"010100111",
  28787=>"000000111",
  28788=>"011001000",
  28789=>"011000111",
  28790=>"100110111",
  28791=>"011011101",
  28792=>"010100100",
  28793=>"000100111",
  28794=>"101110000",
  28795=>"001111011",
  28796=>"000111001",
  28797=>"101100111",
  28798=>"111101111",
  28799=>"001010001",
  28800=>"100101001",
  28801=>"111011111",
  28802=>"000111100",
  28803=>"100100001",
  28804=>"111000000",
  28805=>"100011001",
  28806=>"111010111",
  28807=>"110011001",
  28808=>"001111100",
  28809=>"000000000",
  28810=>"100000111",
  28811=>"011010001",
  28812=>"111001010",
  28813=>"101001111",
  28814=>"110001011",
  28815=>"010010110",
  28816=>"000010101",
  28817=>"011100011",
  28818=>"000100001",
  28819=>"111111111",
  28820=>"101101001",
  28821=>"101011110",
  28822=>"111110010",
  28823=>"111000000",
  28824=>"110101011",
  28825=>"100011000",
  28826=>"010001011",
  28827=>"110101011",
  28828=>"110110100",
  28829=>"101111101",
  28830=>"111011110",
  28831=>"010010100",
  28832=>"110010101",
  28833=>"100101011",
  28834=>"000001001",
  28835=>"111110011",
  28836=>"010001011",
  28837=>"110001001",
  28838=>"010100111",
  28839=>"110110000",
  28840=>"111101001",
  28841=>"110100100",
  28842=>"110000111",
  28843=>"000000011",
  28844=>"000010100",
  28845=>"001100011",
  28846=>"011011101",
  28847=>"001111011",
  28848=>"000010010",
  28849=>"110011010",
  28850=>"111111001",
  28851=>"101101111",
  28852=>"011001111",
  28853=>"010110001",
  28854=>"000111000",
  28855=>"111001010",
  28856=>"000110011",
  28857=>"000001010",
  28858=>"011011001",
  28859=>"100001000",
  28860=>"100100110",
  28861=>"010001100",
  28862=>"010011111",
  28863=>"010111000",
  28864=>"010110110",
  28865=>"111101001",
  28866=>"111111110",
  28867=>"110010001",
  28868=>"101010010",
  28869=>"011100001",
  28870=>"100001000",
  28871=>"001001110",
  28872=>"010100011",
  28873=>"000101101",
  28874=>"100010111",
  28875=>"111010101",
  28876=>"110010000",
  28877=>"001101001",
  28878=>"101100001",
  28879=>"000111001",
  28880=>"000010111",
  28881=>"101011101",
  28882=>"100111100",
  28883=>"111000100",
  28884=>"010110110",
  28885=>"011010101",
  28886=>"010101111",
  28887=>"001101010",
  28888=>"000001000",
  28889=>"101010110",
  28890=>"000010000",
  28891=>"100110111",
  28892=>"110011100",
  28893=>"001000001",
  28894=>"101000111",
  28895=>"000000101",
  28896=>"011111110",
  28897=>"000001001",
  28898=>"111001111",
  28899=>"100100011",
  28900=>"001100000",
  28901=>"011001101",
  28902=>"110010100",
  28903=>"000101101",
  28904=>"110001001",
  28905=>"110100001",
  28906=>"110101111",
  28907=>"000111111",
  28908=>"100111101",
  28909=>"101100111",
  28910=>"010010010",
  28911=>"111101100",
  28912=>"111010100",
  28913=>"000101001",
  28914=>"111010101",
  28915=>"011101110",
  28916=>"100011100",
  28917=>"110010101",
  28918=>"011000111",
  28919=>"000100011",
  28920=>"100111101",
  28921=>"101011111",
  28922=>"001111100",
  28923=>"011010000",
  28924=>"100011010",
  28925=>"111011101",
  28926=>"100011010",
  28927=>"110100111",
  28928=>"011000110",
  28929=>"111010011",
  28930=>"011111101",
  28931=>"000110011",
  28932=>"011100011",
  28933=>"110011101",
  28934=>"010011101",
  28935=>"000100110",
  28936=>"100110000",
  28937=>"000010011",
  28938=>"110110011",
  28939=>"000101101",
  28940=>"100100001",
  28941=>"011101100",
  28942=>"000100001",
  28943=>"111111110",
  28944=>"001111110",
  28945=>"010110101",
  28946=>"111111111",
  28947=>"110110100",
  28948=>"001110101",
  28949=>"001111011",
  28950=>"001011011",
  28951=>"101110001",
  28952=>"010001110",
  28953=>"001001010",
  28954=>"000010000",
  28955=>"100010110",
  28956=>"010101110",
  28957=>"001001011",
  28958=>"001010101",
  28959=>"111001001",
  28960=>"000100100",
  28961=>"111011100",
  28962=>"010000100",
  28963=>"011111111",
  28964=>"010010011",
  28965=>"110011010",
  28966=>"011000011",
  28967=>"100110111",
  28968=>"000010011",
  28969=>"101111010",
  28970=>"101111100",
  28971=>"100010000",
  28972=>"011001100",
  28973=>"110111111",
  28974=>"000011000",
  28975=>"010011010",
  28976=>"010000101",
  28977=>"110100000",
  28978=>"001010110",
  28979=>"011111000",
  28980=>"110000100",
  28981=>"000100000",
  28982=>"101011111",
  28983=>"101101010",
  28984=>"000100001",
  28985=>"011011011",
  28986=>"011101111",
  28987=>"111110100",
  28988=>"110110001",
  28989=>"111111111",
  28990=>"100100111",
  28991=>"001101010",
  28992=>"010010101",
  28993=>"011100000",
  28994=>"010000000",
  28995=>"101001111",
  28996=>"111010111",
  28997=>"100110000",
  28998=>"100110110",
  28999=>"111000010",
  29000=>"000110000",
  29001=>"010110010",
  29002=>"100101100",
  29003=>"101010011",
  29004=>"110001000",
  29005=>"100001010",
  29006=>"000100000",
  29007=>"010010011",
  29008=>"011110110",
  29009=>"101100010",
  29010=>"111110111",
  29011=>"000010011",
  29012=>"001011000",
  29013=>"000110011",
  29014=>"011000001",
  29015=>"101000110",
  29016=>"001010011",
  29017=>"011101001",
  29018=>"011101100",
  29019=>"100100100",
  29020=>"100101010",
  29021=>"100010110",
  29022=>"101001001",
  29023=>"010010001",
  29024=>"000000000",
  29025=>"101000101",
  29026=>"111111111",
  29027=>"000011001",
  29028=>"010111000",
  29029=>"011100011",
  29030=>"010000101",
  29031=>"110010101",
  29032=>"101101010",
  29033=>"100000101",
  29034=>"101110111",
  29035=>"010110000",
  29036=>"000000111",
  29037=>"111011110",
  29038=>"101100110",
  29039=>"111001000",
  29040=>"001010101",
  29041=>"100100010",
  29042=>"000000100",
  29043=>"111100110",
  29044=>"010110000",
  29045=>"000100011",
  29046=>"000111100",
  29047=>"100101010",
  29048=>"000010001",
  29049=>"111101110",
  29050=>"100010011",
  29051=>"001011010",
  29052=>"110000010",
  29053=>"110100000",
  29054=>"000010010",
  29055=>"001011100",
  29056=>"110011000",
  29057=>"011000100",
  29058=>"101000000",
  29059=>"101010110",
  29060=>"101101010",
  29061=>"110110110",
  29062=>"111111111",
  29063=>"000000010",
  29064=>"000111110",
  29065=>"100101101",
  29066=>"011110010",
  29067=>"100000000",
  29068=>"101010010",
  29069=>"000001100",
  29070=>"000000001",
  29071=>"101001101",
  29072=>"001011110",
  29073=>"100000000",
  29074=>"001010111",
  29075=>"110010000",
  29076=>"100011110",
  29077=>"111001101",
  29078=>"101011111",
  29079=>"100000011",
  29080=>"101100111",
  29081=>"101100010",
  29082=>"011001011",
  29083=>"010110000",
  29084=>"001110111",
  29085=>"111101000",
  29086=>"001101100",
  29087=>"111001001",
  29088=>"000101111",
  29089=>"000100110",
  29090=>"101101001",
  29091=>"101111110",
  29092=>"001011010",
  29093=>"110100110",
  29094=>"111101010",
  29095=>"001010010",
  29096=>"001010010",
  29097=>"100000000",
  29098=>"100011111",
  29099=>"011011100",
  29100=>"001000000",
  29101=>"111111010",
  29102=>"000011111",
  29103=>"010111111",
  29104=>"000010010",
  29105=>"100000000",
  29106=>"010101011",
  29107=>"111111000",
  29108=>"011101011",
  29109=>"100000000",
  29110=>"010111001",
  29111=>"101010011",
  29112=>"100101100",
  29113=>"101011001",
  29114=>"011010110",
  29115=>"000100010",
  29116=>"001000000",
  29117=>"100111110",
  29118=>"110000101",
  29119=>"000110111",
  29120=>"010111111",
  29121=>"000000000",
  29122=>"100110001",
  29123=>"111010100",
  29124=>"101000101",
  29125=>"000110011",
  29126=>"110101100",
  29127=>"011001101",
  29128=>"111010111",
  29129=>"111100011",
  29130=>"010010100",
  29131=>"111111100",
  29132=>"100100011",
  29133=>"101000110",
  29134=>"110000111",
  29135=>"100101001",
  29136=>"111101010",
  29137=>"101101111",
  29138=>"011000000",
  29139=>"111110000",
  29140=>"011101011",
  29141=>"100110011",
  29142=>"001101011",
  29143=>"010100000",
  29144=>"011001101",
  29145=>"111010100",
  29146=>"000011010",
  29147=>"101011110",
  29148=>"011001001",
  29149=>"000111111",
  29150=>"010010000",
  29151=>"101000010",
  29152=>"011001101",
  29153=>"000110111",
  29154=>"110010100",
  29155=>"010100010",
  29156=>"001110011",
  29157=>"111011110",
  29158=>"111011010",
  29159=>"000000000",
  29160=>"011011100",
  29161=>"110101101",
  29162=>"110100101",
  29163=>"010001000",
  29164=>"101000001",
  29165=>"011000101",
  29166=>"000100010",
  29167=>"010001110",
  29168=>"001110111",
  29169=>"000101000",
  29170=>"000000001",
  29171=>"000011100",
  29172=>"111001000",
  29173=>"000010010",
  29174=>"101001110",
  29175=>"000110001",
  29176=>"001010101",
  29177=>"000101110",
  29178=>"010011110",
  29179=>"000101010",
  29180=>"100011101",
  29181=>"100111111",
  29182=>"111111101",
  29183=>"011000000",
  29184=>"100101110",
  29185=>"110000001",
  29186=>"010110000",
  29187=>"100001101",
  29188=>"101111000",
  29189=>"110001111",
  29190=>"001110011",
  29191=>"111001101",
  29192=>"001010001",
  29193=>"001111101",
  29194=>"100101000",
  29195=>"100010100",
  29196=>"111100011",
  29197=>"100001101",
  29198=>"101001101",
  29199=>"110101011",
  29200=>"111010001",
  29201=>"011000111",
  29202=>"011011000",
  29203=>"111101010",
  29204=>"101100100",
  29205=>"110001101",
  29206=>"110001110",
  29207=>"100000000",
  29208=>"010010000",
  29209=>"101000001",
  29210=>"011011100",
  29211=>"100010100",
  29212=>"111010010",
  29213=>"010100000",
  29214=>"100111011",
  29215=>"011101101",
  29216=>"000000111",
  29217=>"000010101",
  29218=>"001111001",
  29219=>"100100010",
  29220=>"110000101",
  29221=>"100101000",
  29222=>"101001000",
  29223=>"010001011",
  29224=>"110000111",
  29225=>"001010000",
  29226=>"000000000",
  29227=>"010001011",
  29228=>"101011101",
  29229=>"100010100",
  29230=>"100010011",
  29231=>"001010110",
  29232=>"011110011",
  29233=>"011000001",
  29234=>"101001100",
  29235=>"010111110",
  29236=>"011010001",
  29237=>"000010001",
  29238=>"100001010",
  29239=>"100111001",
  29240=>"000111011",
  29241=>"111010111",
  29242=>"110001100",
  29243=>"000001100",
  29244=>"000110101",
  29245=>"010100011",
  29246=>"101011111",
  29247=>"010111010",
  29248=>"110110000",
  29249=>"010001100",
  29250=>"000111101",
  29251=>"101100110",
  29252=>"110001010",
  29253=>"011111110",
  29254=>"011001001",
  29255=>"011000111",
  29256=>"001000110",
  29257=>"111010110",
  29258=>"100000110",
  29259=>"000000011",
  29260=>"111100000",
  29261=>"100010100",
  29262=>"100000011",
  29263=>"001110000",
  29264=>"110010010",
  29265=>"100110100",
  29266=>"001000111",
  29267=>"001101100",
  29268=>"001010110",
  29269=>"000111011",
  29270=>"110011100",
  29271=>"100110111",
  29272=>"000101111",
  29273=>"001010111",
  29274=>"110101110",
  29275=>"110111011",
  29276=>"111111011",
  29277=>"011001101",
  29278=>"001111000",
  29279=>"011100101",
  29280=>"001001110",
  29281=>"000001101",
  29282=>"110101110",
  29283=>"010111101",
  29284=>"010001010",
  29285=>"100111111",
  29286=>"111110000",
  29287=>"100010001",
  29288=>"000001010",
  29289=>"011001000",
  29290=>"111111111",
  29291=>"000011010",
  29292=>"100001011",
  29293=>"110101100",
  29294=>"000010011",
  29295=>"011001010",
  29296=>"111101000",
  29297=>"000110000",
  29298=>"100101010",
  29299=>"011011010",
  29300=>"010010001",
  29301=>"111000010",
  29302=>"000000001",
  29303=>"000001010",
  29304=>"011111011",
  29305=>"011001100",
  29306=>"111111000",
  29307=>"000100101",
  29308=>"010010100",
  29309=>"110111111",
  29310=>"110100011",
  29311=>"100011111",
  29312=>"011101111",
  29313=>"101011110",
  29314=>"111100101",
  29315=>"111001010",
  29316=>"101000011",
  29317=>"011011000",
  29318=>"010001010",
  29319=>"111011000",
  29320=>"001001111",
  29321=>"010000000",
  29322=>"011011010",
  29323=>"100001010",
  29324=>"111111101",
  29325=>"111110000",
  29326=>"110100001",
  29327=>"100001111",
  29328=>"111101010",
  29329=>"100101111",
  29330=>"010110011",
  29331=>"011101101",
  29332=>"000010011",
  29333=>"111110000",
  29334=>"000110111",
  29335=>"011110010",
  29336=>"111110011",
  29337=>"100001011",
  29338=>"100011001",
  29339=>"000000011",
  29340=>"010001110",
  29341=>"111000001",
  29342=>"100111111",
  29343=>"111100101",
  29344=>"111101100",
  29345=>"110101110",
  29346=>"011000001",
  29347=>"100111000",
  29348=>"001010110",
  29349=>"000010111",
  29350=>"000000000",
  29351=>"001101001",
  29352=>"010010111",
  29353=>"011001000",
  29354=>"100010101",
  29355=>"001001100",
  29356=>"100100111",
  29357=>"010100001",
  29358=>"000111100",
  29359=>"001100110",
  29360=>"011110111",
  29361=>"010011101",
  29362=>"001101100",
  29363=>"100001110",
  29364=>"010001000",
  29365=>"111000000",
  29366=>"011011110",
  29367=>"010111111",
  29368=>"000100111",
  29369=>"111011100",
  29370=>"100111100",
  29371=>"111101100",
  29372=>"011110110",
  29373=>"010010111",
  29374=>"000100110",
  29375=>"010000011",
  29376=>"000100010",
  29377=>"101110100",
  29378=>"110000110",
  29379=>"010101000",
  29380=>"000000111",
  29381=>"011100011",
  29382=>"110010100",
  29383=>"111111101",
  29384=>"101000001",
  29385=>"000011100",
  29386=>"010000010",
  29387=>"000000100",
  29388=>"100111111",
  29389=>"111101001",
  29390=>"011011100",
  29391=>"110110010",
  29392=>"100111011",
  29393=>"110101001",
  29394=>"000011001",
  29395=>"101101111",
  29396=>"001000000",
  29397=>"001001001",
  29398=>"010011101",
  29399=>"001000110",
  29400=>"000111011",
  29401=>"000100011",
  29402=>"100110101",
  29403=>"110111000",
  29404=>"100110001",
  29405=>"110111000",
  29406=>"011010000",
  29407=>"000000000",
  29408=>"110010100",
  29409=>"001100010",
  29410=>"111110001",
  29411=>"111001110",
  29412=>"111011000",
  29413=>"110111010",
  29414=>"011100111",
  29415=>"001101100",
  29416=>"000100011",
  29417=>"100010100",
  29418=>"100100000",
  29419=>"010000000",
  29420=>"000001011",
  29421=>"101100011",
  29422=>"101001100",
  29423=>"010100101",
  29424=>"010000011",
  29425=>"000011000",
  29426=>"100111000",
  29427=>"001110010",
  29428=>"110001101",
  29429=>"001010100",
  29430=>"000100001",
  29431=>"101110110",
  29432=>"011111100",
  29433=>"110110101",
  29434=>"101110011",
  29435=>"000001001",
  29436=>"101011000",
  29437=>"010101110",
  29438=>"110001110",
  29439=>"111101001",
  29440=>"111101000",
  29441=>"111111000",
  29442=>"101101110",
  29443=>"011110101",
  29444=>"001011111",
  29445=>"000001001",
  29446=>"010000010",
  29447=>"010111101",
  29448=>"000011100",
  29449=>"010000010",
  29450=>"000001011",
  29451=>"111000000",
  29452=>"001001111",
  29453=>"000111111",
  29454=>"001010101",
  29455=>"010110101",
  29456=>"001101000",
  29457=>"000010010",
  29458=>"111000110",
  29459=>"111011101",
  29460=>"100001110",
  29461=>"111100111",
  29462=>"011001000",
  29463=>"001100101",
  29464=>"101100000",
  29465=>"000001110",
  29466=>"000000001",
  29467=>"100010110",
  29468=>"001111100",
  29469=>"011100111",
  29470=>"111000110",
  29471=>"011110001",
  29472=>"001111000",
  29473=>"111001000",
  29474=>"011101101",
  29475=>"011110101",
  29476=>"010111011",
  29477=>"000000000",
  29478=>"010100101",
  29479=>"111101110",
  29480=>"010010111",
  29481=>"010101000",
  29482=>"001110010",
  29483=>"111111100",
  29484=>"011001011",
  29485=>"011101111",
  29486=>"000011101",
  29487=>"111011011",
  29488=>"000100010",
  29489=>"110010100",
  29490=>"001001000",
  29491=>"110000100",
  29492=>"000000000",
  29493=>"010100010",
  29494=>"011110101",
  29495=>"101111101",
  29496=>"111000011",
  29497=>"101100111",
  29498=>"001000000",
  29499=>"100000000",
  29500=>"010010111",
  29501=>"101100100",
  29502=>"110011100",
  29503=>"011100110",
  29504=>"001000100",
  29505=>"001011000",
  29506=>"000011100",
  29507=>"110001000",
  29508=>"000100110",
  29509=>"101000111",
  29510=>"001000100",
  29511=>"101011111",
  29512=>"011101000",
  29513=>"101010110",
  29514=>"011110110",
  29515=>"010001111",
  29516=>"100100001",
  29517=>"000010011",
  29518=>"101010001",
  29519=>"010011101",
  29520=>"001110001",
  29521=>"010010110",
  29522=>"000100001",
  29523=>"101000001",
  29524=>"010010001",
  29525=>"101011111",
  29526=>"111110010",
  29527=>"100111101",
  29528=>"111011010",
  29529=>"010101010",
  29530=>"000110110",
  29531=>"001011110",
  29532=>"100011011",
  29533=>"010011011",
  29534=>"110101100",
  29535=>"000100101",
  29536=>"011010100",
  29537=>"111110111",
  29538=>"001110000",
  29539=>"001010100",
  29540=>"011010111",
  29541=>"011111111",
  29542=>"110001001",
  29543=>"101001100",
  29544=>"110101010",
  29545=>"001101001",
  29546=>"101011101",
  29547=>"110111110",
  29548=>"101011000",
  29549=>"100011000",
  29550=>"100111111",
  29551=>"100110001",
  29552=>"000000100",
  29553=>"000111000",
  29554=>"111101000",
  29555=>"101010000",
  29556=>"101101011",
  29557=>"101111110",
  29558=>"110001001",
  29559=>"110110101",
  29560=>"011001100",
  29561=>"111111010",
  29562=>"111101000",
  29563=>"000001000",
  29564=>"111000111",
  29565=>"011110001",
  29566=>"110000011",
  29567=>"101101010",
  29568=>"110010001",
  29569=>"011000000",
  29570=>"101010111",
  29571=>"100111110",
  29572=>"000110010",
  29573=>"101001111",
  29574=>"000100110",
  29575=>"011011110",
  29576=>"100000001",
  29577=>"100011110",
  29578=>"001011101",
  29579=>"101001001",
  29580=>"111011000",
  29581=>"001000011",
  29582=>"110110011",
  29583=>"010101101",
  29584=>"000001000",
  29585=>"000001011",
  29586=>"010110110",
  29587=>"111001001",
  29588=>"001010010",
  29589=>"101111000",
  29590=>"000101001",
  29591=>"101100001",
  29592=>"101000011",
  29593=>"100000010",
  29594=>"001100110",
  29595=>"010110110",
  29596=>"110010011",
  29597=>"100001110",
  29598=>"011010110",
  29599=>"001100110",
  29600=>"000111100",
  29601=>"001001010",
  29602=>"011000110",
  29603=>"001001101",
  29604=>"001110011",
  29605=>"110110100",
  29606=>"110101010",
  29607=>"100111111",
  29608=>"000000111",
  29609=>"010101101",
  29610=>"110101101",
  29611=>"110001001",
  29612=>"001010001",
  29613=>"000000110",
  29614=>"110010110",
  29615=>"000000110",
  29616=>"000001001",
  29617=>"001101100",
  29618=>"110100111",
  29619=>"100111000",
  29620=>"111111010",
  29621=>"101001001",
  29622=>"010011111",
  29623=>"110111100",
  29624=>"010000100",
  29625=>"010001101",
  29626=>"010010010",
  29627=>"001100111",
  29628=>"001010001",
  29629=>"010100000",
  29630=>"111101010",
  29631=>"111110000",
  29632=>"101100011",
  29633=>"101011000",
  29634=>"010011001",
  29635=>"111101010",
  29636=>"101110001",
  29637=>"011001010",
  29638=>"011110000",
  29639=>"000000011",
  29640=>"000101100",
  29641=>"111111010",
  29642=>"101010110",
  29643=>"100010001",
  29644=>"000011011",
  29645=>"111101000",
  29646=>"111001110",
  29647=>"010101111",
  29648=>"101100010",
  29649=>"001111111",
  29650=>"101100001",
  29651=>"010111100",
  29652=>"010100110",
  29653=>"101110010",
  29654=>"111110010",
  29655=>"000010000",
  29656=>"000101110",
  29657=>"111000100",
  29658=>"001010011",
  29659=>"111001011",
  29660=>"100100000",
  29661=>"110110110",
  29662=>"111101001",
  29663=>"010001001",
  29664=>"111111101",
  29665=>"000011011",
  29666=>"110001100",
  29667=>"000100111",
  29668=>"111001001",
  29669=>"010010100",
  29670=>"000111010",
  29671=>"011101011",
  29672=>"000110001",
  29673=>"111001101",
  29674=>"100100010",
  29675=>"000000001",
  29676=>"110000000",
  29677=>"100011100",
  29678=>"110000001",
  29679=>"111100011",
  29680=>"100100001",
  29681=>"000010000",
  29682=>"111110000",
  29683=>"011101001",
  29684=>"010010000",
  29685=>"111100000",
  29686=>"001000001",
  29687=>"001010000",
  29688=>"110100000",
  29689=>"001110001",
  29690=>"001000100",
  29691=>"010011001",
  29692=>"111110001",
  29693=>"011110100",
  29694=>"010001011",
  29695=>"011010011",
  29696=>"010001011",
  29697=>"011111111",
  29698=>"101000100",
  29699=>"111111100",
  29700=>"100001001",
  29701=>"110111011",
  29702=>"110111011",
  29703=>"111000000",
  29704=>"011101110",
  29705=>"010000110",
  29706=>"101111111",
  29707=>"101000110",
  29708=>"110101111",
  29709=>"111011001",
  29710=>"111101111",
  29711=>"010111100",
  29712=>"001000010",
  29713=>"110100001",
  29714=>"110101110",
  29715=>"101110101",
  29716=>"111001111",
  29717=>"001111000",
  29718=>"111100000",
  29719=>"110000010",
  29720=>"100111001",
  29721=>"010000011",
  29722=>"000110101",
  29723=>"001100011",
  29724=>"100001010",
  29725=>"000010001",
  29726=>"111010100",
  29727=>"110110001",
  29728=>"010011110",
  29729=>"111110111",
  29730=>"100000111",
  29731=>"000101111",
  29732=>"010100010",
  29733=>"001000000",
  29734=>"111100100",
  29735=>"011010000",
  29736=>"110000000",
  29737=>"000000010",
  29738=>"000111011",
  29739=>"010111011",
  29740=>"010101001",
  29741=>"000101011",
  29742=>"011101011",
  29743=>"001011011",
  29744=>"111111100",
  29745=>"101011110",
  29746=>"010000100",
  29747=>"000000010",
  29748=>"111000000",
  29749=>"111011011",
  29750=>"111101011",
  29751=>"011110010",
  29752=>"110111010",
  29753=>"011111101",
  29754=>"000000101",
  29755=>"111000111",
  29756=>"000010011",
  29757=>"111010001",
  29758=>"011011001",
  29759=>"000101011",
  29760=>"110101011",
  29761=>"001000000",
  29762=>"001011110",
  29763=>"101010011",
  29764=>"100110010",
  29765=>"100001101",
  29766=>"100110100",
  29767=>"000100011",
  29768=>"001100101",
  29769=>"010000000",
  29770=>"110010011",
  29771=>"011001111",
  29772=>"001100000",
  29773=>"010010010",
  29774=>"101100010",
  29775=>"010110010",
  29776=>"111101011",
  29777=>"000011001",
  29778=>"011110101",
  29779=>"001011111",
  29780=>"111011100",
  29781=>"011110010",
  29782=>"110011110",
  29783=>"111000110",
  29784=>"111010110",
  29785=>"110101100",
  29786=>"011010000",
  29787=>"101010011",
  29788=>"000000110",
  29789=>"001100100",
  29790=>"111101100",
  29791=>"001010010",
  29792=>"000111110",
  29793=>"110110110",
  29794=>"011110101",
  29795=>"000111110",
  29796=>"001010010",
  29797=>"100011001",
  29798=>"011110000",
  29799=>"001110010",
  29800=>"110111110",
  29801=>"110011011",
  29802=>"101000011",
  29803=>"000001010",
  29804=>"100111001",
  29805=>"000100101",
  29806=>"001010110",
  29807=>"001100000",
  29808=>"100001101",
  29809=>"010001000",
  29810=>"001001011",
  29811=>"110110110",
  29812=>"001010101",
  29813=>"001001111",
  29814=>"111100111",
  29815=>"011100111",
  29816=>"101100010",
  29817=>"000100001",
  29818=>"001110001",
  29819=>"000011001",
  29820=>"000011100",
  29821=>"000011001",
  29822=>"001001011",
  29823=>"110001100",
  29824=>"101110011",
  29825=>"011100001",
  29826=>"010010000",
  29827=>"100001010",
  29828=>"000001000",
  29829=>"111011101",
  29830=>"010000010",
  29831=>"011011110",
  29832=>"000110100",
  29833=>"010011000",
  29834=>"101001010",
  29835=>"000100010",
  29836=>"111100000",
  29837=>"100100101",
  29838=>"011000100",
  29839=>"110000110",
  29840=>"110110000",
  29841=>"110110101",
  29842=>"100001101",
  29843=>"101010111",
  29844=>"110101001",
  29845=>"001100111",
  29846=>"100001001",
  29847=>"000010011",
  29848=>"110101111",
  29849=>"010001010",
  29850=>"011001001",
  29851=>"100101101",
  29852=>"111010110",
  29853=>"100111010",
  29854=>"101111010",
  29855=>"010011111",
  29856=>"010101100",
  29857=>"101011101",
  29858=>"000101001",
  29859=>"001110101",
  29860=>"010001000",
  29861=>"111001100",
  29862=>"000000111",
  29863=>"010101111",
  29864=>"110000010",
  29865=>"000111110",
  29866=>"111011110",
  29867=>"011100001",
  29868=>"010101111",
  29869=>"001000000",
  29870=>"001000001",
  29871=>"001011111",
  29872=>"001011100",
  29873=>"000011111",
  29874=>"011100101",
  29875=>"000011110",
  29876=>"101110011",
  29877=>"101100101",
  29878=>"110101100",
  29879=>"000010110",
  29880=>"111010001",
  29881=>"101001111",
  29882=>"010000001",
  29883=>"100000111",
  29884=>"010000000",
  29885=>"100001010",
  29886=>"010011111",
  29887=>"110000000",
  29888=>"101101000",
  29889=>"011001111",
  29890=>"101000111",
  29891=>"101110110",
  29892=>"001100011",
  29893=>"110011111",
  29894=>"111111111",
  29895=>"101011101",
  29896=>"110001111",
  29897=>"000000111",
  29898=>"101001101",
  29899=>"000011101",
  29900=>"101101101",
  29901=>"000111100",
  29902=>"000111001",
  29903=>"100100011",
  29904=>"101000101",
  29905=>"100101000",
  29906=>"000011101",
  29907=>"011100100",
  29908=>"101111110",
  29909=>"010101001",
  29910=>"000110101",
  29911=>"111111110",
  29912=>"001011110",
  29913=>"111011110",
  29914=>"101000100",
  29915=>"011100110",
  29916=>"010101011",
  29917=>"011001100",
  29918=>"000010001",
  29919=>"111110101",
  29920=>"101010100",
  29921=>"111101010",
  29922=>"101101100",
  29923=>"000111010",
  29924=>"100101100",
  29925=>"001101110",
  29926=>"011001000",
  29927=>"111100000",
  29928=>"001000001",
  29929=>"010011100",
  29930=>"000001001",
  29931=>"011110111",
  29932=>"111010100",
  29933=>"010111000",
  29934=>"001110111",
  29935=>"001100000",
  29936=>"111100100",
  29937=>"111011111",
  29938=>"011010100",
  29939=>"010100100",
  29940=>"101000000",
  29941=>"110001000",
  29942=>"011101100",
  29943=>"010011101",
  29944=>"010111101",
  29945=>"001111001",
  29946=>"000101000",
  29947=>"000100111",
  29948=>"110110110",
  29949=>"100101111",
  29950=>"000100101",
  29951=>"111110110",
  29952=>"001001101",
  29953=>"001001000",
  29954=>"110010001",
  29955=>"001010100",
  29956=>"011101100",
  29957=>"110011001",
  29958=>"000010110",
  29959=>"110111101",
  29960=>"011010000",
  29961=>"010000001",
  29962=>"001001000",
  29963=>"010011001",
  29964=>"010111011",
  29965=>"000011111",
  29966=>"000011111",
  29967=>"000001001",
  29968=>"001111010",
  29969=>"110111100",
  29970=>"000010001",
  29971=>"101000000",
  29972=>"100000010",
  29973=>"100011010",
  29974=>"000001110",
  29975=>"110111111",
  29976=>"110011010",
  29977=>"111000000",
  29978=>"011010010",
  29979=>"001001000",
  29980=>"110010011",
  29981=>"001001110",
  29982=>"101110011",
  29983=>"000000100",
  29984=>"100101100",
  29985=>"001110101",
  29986=>"111111001",
  29987=>"001101010",
  29988=>"101101100",
  29989=>"011001111",
  29990=>"000000100",
  29991=>"101111010",
  29992=>"010011010",
  29993=>"111010101",
  29994=>"010110010",
  29995=>"000001111",
  29996=>"000110100",
  29997=>"000110101",
  29998=>"010011010",
  29999=>"010010100",
  30000=>"011010011",
  30001=>"001010101",
  30002=>"111111010",
  30003=>"111110101",
  30004=>"000111110",
  30005=>"111101000",
  30006=>"000001011",
  30007=>"011110010",
  30008=>"111000101",
  30009=>"010011000",
  30010=>"111011010",
  30011=>"010000011",
  30012=>"101100110",
  30013=>"111010111",
  30014=>"010001010",
  30015=>"111001000",
  30016=>"000111011",
  30017=>"111001011",
  30018=>"000100011",
  30019=>"000101010",
  30020=>"010101000",
  30021=>"100100001",
  30022=>"000001101",
  30023=>"011111111",
  30024=>"010010000",
  30025=>"010100011",
  30026=>"101111100",
  30027=>"010000110",
  30028=>"001001000",
  30029=>"101000010",
  30030=>"111100111",
  30031=>"001000001",
  30032=>"111110110",
  30033=>"110000101",
  30034=>"000101111",
  30035=>"100100001",
  30036=>"010100111",
  30037=>"110111001",
  30038=>"001011100",
  30039=>"100001000",
  30040=>"111011000",
  30041=>"111101111",
  30042=>"101110101",
  30043=>"000010101",
  30044=>"100001000",
  30045=>"011111101",
  30046=>"110101111",
  30047=>"111111110",
  30048=>"110100111",
  30049=>"000001110",
  30050=>"101100011",
  30051=>"010011111",
  30052=>"000000010",
  30053=>"100001110",
  30054=>"100101011",
  30055=>"001011110",
  30056=>"111011010",
  30057=>"111001010",
  30058=>"001110011",
  30059=>"000000101",
  30060=>"111110111",
  30061=>"110110110",
  30062=>"111000111",
  30063=>"010001100",
  30064=>"110010101",
  30065=>"010010000",
  30066=>"111000001",
  30067=>"111111000",
  30068=>"111001101",
  30069=>"000010001",
  30070=>"011101101",
  30071=>"110000100",
  30072=>"111000101",
  30073=>"110010001",
  30074=>"101010111",
  30075=>"011001010",
  30076=>"000011000",
  30077=>"100011100",
  30078=>"010111110",
  30079=>"011110100",
  30080=>"100010110",
  30081=>"011011011",
  30082=>"001001110",
  30083=>"110011000",
  30084=>"110011001",
  30085=>"100000001",
  30086=>"101001100",
  30087=>"100101011",
  30088=>"011100000",
  30089=>"111001010",
  30090=>"110101011",
  30091=>"101111111",
  30092=>"000101010",
  30093=>"001111111",
  30094=>"010010001",
  30095=>"011001011",
  30096=>"001011001",
  30097=>"000011100",
  30098=>"010111110",
  30099=>"101000100",
  30100=>"111101110",
  30101=>"000001101",
  30102=>"000010010",
  30103=>"111110001",
  30104=>"110010111",
  30105=>"011000011",
  30106=>"101010010",
  30107=>"010110011",
  30108=>"010100100",
  30109=>"110010010",
  30110=>"110110001",
  30111=>"101000101",
  30112=>"101110001",
  30113=>"000010111",
  30114=>"110000010",
  30115=>"000101000",
  30116=>"101110100",
  30117=>"011111000",
  30118=>"000110011",
  30119=>"101001000",
  30120=>"011111010",
  30121=>"010111100",
  30122=>"110001010",
  30123=>"000000011",
  30124=>"001111101",
  30125=>"110110000",
  30126=>"100110011",
  30127=>"010000001",
  30128=>"111011100",
  30129=>"100000000",
  30130=>"100100011",
  30131=>"010011111",
  30132=>"000000100",
  30133=>"001001000",
  30134=>"011100001",
  30135=>"100111100",
  30136=>"110111001",
  30137=>"100010101",
  30138=>"000000110",
  30139=>"110101101",
  30140=>"101100011",
  30141=>"000011000",
  30142=>"010011110",
  30143=>"100111110",
  30144=>"011011001",
  30145=>"001011111",
  30146=>"000100010",
  30147=>"111100000",
  30148=>"001001011",
  30149=>"101010000",
  30150=>"101100110",
  30151=>"000001011",
  30152=>"000000101",
  30153=>"100100010",
  30154=>"110101111",
  30155=>"010101101",
  30156=>"001011011",
  30157=>"001101101",
  30158=>"000010010",
  30159=>"001001011",
  30160=>"011010110",
  30161=>"000001100",
  30162=>"011100001",
  30163=>"000000010",
  30164=>"011101010",
  30165=>"000110100",
  30166=>"000000001",
  30167=>"101000111",
  30168=>"101110110",
  30169=>"101111010",
  30170=>"000000100",
  30171=>"100011000",
  30172=>"110110001",
  30173=>"000111111",
  30174=>"111111111",
  30175=>"110001001",
  30176=>"111101010",
  30177=>"111010000",
  30178=>"111001001",
  30179=>"110011100",
  30180=>"111001010",
  30181=>"110111100",
  30182=>"011011000",
  30183=>"010010011",
  30184=>"110001000",
  30185=>"011100000",
  30186=>"100110001",
  30187=>"001011010",
  30188=>"000100000",
  30189=>"111100000",
  30190=>"110011010",
  30191=>"111101000",
  30192=>"111010111",
  30193=>"011001111",
  30194=>"010100100",
  30195=>"000100000",
  30196=>"001100111",
  30197=>"110001011",
  30198=>"000011000",
  30199=>"111111110",
  30200=>"011101001",
  30201=>"100101110",
  30202=>"110100000",
  30203=>"010111001",
  30204=>"100100001",
  30205=>"011111110",
  30206=>"000111010",
  30207=>"010110011",
  30208=>"111011000",
  30209=>"110100100",
  30210=>"001100001",
  30211=>"000011100",
  30212=>"011100110",
  30213=>"110001110",
  30214=>"000011001",
  30215=>"111111001",
  30216=>"111110011",
  30217=>"011110010",
  30218=>"010101001",
  30219=>"101111110",
  30220=>"001001000",
  30221=>"000001001",
  30222=>"000110000",
  30223=>"101011010",
  30224=>"110010001",
  30225=>"000011000",
  30226=>"011011010",
  30227=>"100100000",
  30228=>"010011100",
  30229=>"011101111",
  30230=>"110110011",
  30231=>"011000110",
  30232=>"001110000",
  30233=>"100010000",
  30234=>"101010001",
  30235=>"000111001",
  30236=>"010010100",
  30237=>"111000011",
  30238=>"110111100",
  30239=>"101101001",
  30240=>"011110011",
  30241=>"010000011",
  30242=>"011001000",
  30243=>"000100110",
  30244=>"011101100",
  30245=>"101011000",
  30246=>"111110010",
  30247=>"111100101",
  30248=>"001010000",
  30249=>"100011101",
  30250=>"100101101",
  30251=>"110000010",
  30252=>"101101100",
  30253=>"101010110",
  30254=>"100000011",
  30255=>"010000000",
  30256=>"111001111",
  30257=>"100111011",
  30258=>"001010001",
  30259=>"101001100",
  30260=>"101110011",
  30261=>"000000001",
  30262=>"110100011",
  30263=>"010000011",
  30264=>"010110110",
  30265=>"101110111",
  30266=>"001100011",
  30267=>"011011000",
  30268=>"110100111",
  30269=>"000001101",
  30270=>"001100101",
  30271=>"010101001",
  30272=>"100111111",
  30273=>"001001000",
  30274=>"011010001",
  30275=>"110000011",
  30276=>"110111000",
  30277=>"001011001",
  30278=>"001001100",
  30279=>"000100011",
  30280=>"010011000",
  30281=>"111001110",
  30282=>"000000110",
  30283=>"101001111",
  30284=>"000101011",
  30285=>"011000010",
  30286=>"100010111",
  30287=>"100000010",
  30288=>"101001000",
  30289=>"011001000",
  30290=>"000110011",
  30291=>"001111101",
  30292=>"100110000",
  30293=>"111001111",
  30294=>"110010110",
  30295=>"101111101",
  30296=>"011110011",
  30297=>"111010001",
  30298=>"100011110",
  30299=>"100001000",
  30300=>"111001100",
  30301=>"010111011",
  30302=>"110101111",
  30303=>"110000001",
  30304=>"000101001",
  30305=>"100001011",
  30306=>"110100100",
  30307=>"010010000",
  30308=>"011110110",
  30309=>"100110011",
  30310=>"001010010",
  30311=>"111010101",
  30312=>"000000111",
  30313=>"010101100",
  30314=>"110001111",
  30315=>"010011001",
  30316=>"011011111",
  30317=>"101010001",
  30318=>"011000011",
  30319=>"011111001",
  30320=>"110000011",
  30321=>"011000101",
  30322=>"110110011",
  30323=>"001110000",
  30324=>"100110001",
  30325=>"111111101",
  30326=>"011011110",
  30327=>"101101011",
  30328=>"111011101",
  30329=>"100001001",
  30330=>"101011011",
  30331=>"110000010",
  30332=>"010101100",
  30333=>"110001101",
  30334=>"000010010",
  30335=>"111110010",
  30336=>"100000001",
  30337=>"001101000",
  30338=>"010111011",
  30339=>"010011011",
  30340=>"001001001",
  30341=>"010110101",
  30342=>"111110110",
  30343=>"111011100",
  30344=>"010011001",
  30345=>"001010100",
  30346=>"111000100",
  30347=>"000000110",
  30348=>"101011110",
  30349=>"000100111",
  30350=>"000100001",
  30351=>"011001100",
  30352=>"010011100",
  30353=>"011101111",
  30354=>"010101010",
  30355=>"011111101",
  30356=>"011111010",
  30357=>"011011000",
  30358=>"011010001",
  30359=>"000101111",
  30360=>"111101000",
  30361=>"001011111",
  30362=>"011111110",
  30363=>"100110000",
  30364=>"000010111",
  30365=>"011011001",
  30366=>"000001000",
  30367=>"010011110",
  30368=>"010000101",
  30369=>"111011110",
  30370=>"000000011",
  30371=>"001010111",
  30372=>"110111010",
  30373=>"010011111",
  30374=>"100001011",
  30375=>"000000010",
  30376=>"100001000",
  30377=>"000110000",
  30378=>"001110000",
  30379=>"100110110",
  30380=>"000100010",
  30381=>"001000010",
  30382=>"100111010",
  30383=>"111001000",
  30384=>"001100000",
  30385=>"000010010",
  30386=>"001010000",
  30387=>"000011000",
  30388=>"000011101",
  30389=>"110111101",
  30390=>"000001010",
  30391=>"110101001",
  30392=>"111000100",
  30393=>"011010101",
  30394=>"111001001",
  30395=>"001101110",
  30396=>"111000100",
  30397=>"011110110",
  30398=>"000100110",
  30399=>"111100010",
  30400=>"101111110",
  30401=>"010000011",
  30402=>"001110111",
  30403=>"001010111",
  30404=>"010100100",
  30405=>"010111110",
  30406=>"111100110",
  30407=>"110101110",
  30408=>"000101100",
  30409=>"000101100",
  30410=>"111010001",
  30411=>"110101101",
  30412=>"100010110",
  30413=>"101000001",
  30414=>"111100011",
  30415=>"011110010",
  30416=>"001000000",
  30417=>"001100010",
  30418=>"100010001",
  30419=>"001110000",
  30420=>"010001000",
  30421=>"010110111",
  30422=>"000111101",
  30423=>"000011100",
  30424=>"111110110",
  30425=>"011110110",
  30426=>"000101100",
  30427=>"111000100",
  30428=>"000000001",
  30429=>"000011110",
  30430=>"111001000",
  30431=>"000101000",
  30432=>"000111010",
  30433=>"011000010",
  30434=>"101111000",
  30435=>"011011111",
  30436=>"011000111",
  30437=>"111011010",
  30438=>"101000111",
  30439=>"100000111",
  30440=>"111011010",
  30441=>"110010111",
  30442=>"000001001",
  30443=>"111010001",
  30444=>"110011111",
  30445=>"110011011",
  30446=>"100101011",
  30447=>"011010001",
  30448=>"011100000",
  30449=>"111110101",
  30450=>"100111111",
  30451=>"101011101",
  30452=>"001001000",
  30453=>"100111000",
  30454=>"100001001",
  30455=>"100001010",
  30456=>"110101001",
  30457=>"101110101",
  30458=>"001000001",
  30459=>"010001101",
  30460=>"001110110",
  30461=>"000110110",
  30462=>"111010101",
  30463=>"010000000",
  30464=>"000101000",
  30465=>"011111101",
  30466=>"011101010",
  30467=>"000010111",
  30468=>"101011000",
  30469=>"111101100",
  30470=>"000000110",
  30471=>"011110110",
  30472=>"110000001",
  30473=>"111111000",
  30474=>"010000001",
  30475=>"110110001",
  30476=>"001011111",
  30477=>"111001001",
  30478=>"001011101",
  30479=>"101001011",
  30480=>"100101000",
  30481=>"001000001",
  30482=>"010100000",
  30483=>"001100011",
  30484=>"101010100",
  30485=>"100100001",
  30486=>"001110011",
  30487=>"101000111",
  30488=>"011110010",
  30489=>"000010001",
  30490=>"000011100",
  30491=>"110101101",
  30492=>"110001101",
  30493=>"110100000",
  30494=>"000100100",
  30495=>"110010111",
  30496=>"010011110",
  30497=>"111000110",
  30498=>"011011000",
  30499=>"100101111",
  30500=>"101011111",
  30501=>"000101000",
  30502=>"101001010",
  30503=>"111011111",
  30504=>"000111000",
  30505=>"010111011",
  30506=>"100110011",
  30507=>"010110001",
  30508=>"000011000",
  30509=>"000001111",
  30510=>"000001111",
  30511=>"101000100",
  30512=>"000111000",
  30513=>"100000110",
  30514=>"101110010",
  30515=>"110111111",
  30516=>"111010000",
  30517=>"011010001",
  30518=>"001011101",
  30519=>"010101000",
  30520=>"011011100",
  30521=>"101101110",
  30522=>"011001110",
  30523=>"101001011",
  30524=>"001111011",
  30525=>"101110100",
  30526=>"110001110",
  30527=>"111010110",
  30528=>"110100011",
  30529=>"011101010",
  30530=>"110011011",
  30531=>"011100110",
  30532=>"001111100",
  30533=>"000101101",
  30534=>"000010110",
  30535=>"111000001",
  30536=>"110111111",
  30537=>"110001001",
  30538=>"000111110",
  30539=>"001110111",
  30540=>"011101010",
  30541=>"011101000",
  30542=>"100000111",
  30543=>"011110110",
  30544=>"000000110",
  30545=>"101111001",
  30546=>"001011110",
  30547=>"100011001",
  30548=>"111100001",
  30549=>"000111111",
  30550=>"010011101",
  30551=>"111001010",
  30552=>"000001000",
  30553=>"101110110",
  30554=>"110011000",
  30555=>"100100011",
  30556=>"111010101",
  30557=>"001010000",
  30558=>"000001011",
  30559=>"000000011",
  30560=>"001011110",
  30561=>"101010000",
  30562=>"010100010",
  30563=>"001110111",
  30564=>"001000100",
  30565=>"110011000",
  30566=>"100000000",
  30567=>"101111111",
  30568=>"101100110",
  30569=>"100100001",
  30570=>"000110111",
  30571=>"011110100",
  30572=>"000110111",
  30573=>"010100110",
  30574=>"101000001",
  30575=>"100000001",
  30576=>"001111001",
  30577=>"000010101",
  30578=>"011101100",
  30579=>"011010111",
  30580=>"110000000",
  30581=>"101100111",
  30582=>"011010000",
  30583=>"011100000",
  30584=>"011011001",
  30585=>"001101011",
  30586=>"111101001",
  30587=>"100100111",
  30588=>"010001010",
  30589=>"001111101",
  30590=>"011010111",
  30591=>"100000110",
  30592=>"100100100",
  30593=>"010000011",
  30594=>"110110011",
  30595=>"000001100",
  30596=>"010000010",
  30597=>"101001001",
  30598=>"000000000",
  30599=>"100100110",
  30600=>"000010011",
  30601=>"000111001",
  30602=>"000000110",
  30603=>"111011100",
  30604=>"000100000",
  30605=>"000100101",
  30606=>"110000100",
  30607=>"110111111",
  30608=>"000000111",
  30609=>"011110010",
  30610=>"101111000",
  30611=>"101111111",
  30612=>"010110111",
  30613=>"001111111",
  30614=>"000111000",
  30615=>"000101001",
  30616=>"110101011",
  30617=>"100110010",
  30618=>"100001111",
  30619=>"000011100",
  30620=>"001000001",
  30621=>"100000010",
  30622=>"001011011",
  30623=>"000010001",
  30624=>"100011100",
  30625=>"011110011",
  30626=>"100101111",
  30627=>"011011011",
  30628=>"011001010",
  30629=>"111111110",
  30630=>"101100101",
  30631=>"100001010",
  30632=>"111101011",
  30633=>"111100001",
  30634=>"010011010",
  30635=>"011010001",
  30636=>"101010011",
  30637=>"011100111",
  30638=>"011011000",
  30639=>"001101111",
  30640=>"110000001",
  30641=>"111101010",
  30642=>"100011111",
  30643=>"000011000",
  30644=>"111101011",
  30645=>"111010111",
  30646=>"100010010",
  30647=>"000110110",
  30648=>"011101100",
  30649=>"001110111",
  30650=>"001011101",
  30651=>"110011111",
  30652=>"110111110",
  30653=>"000000110",
  30654=>"100100100",
  30655=>"000011111",
  30656=>"011110101",
  30657=>"110101110",
  30658=>"000010000",
  30659=>"010000011",
  30660=>"111101110",
  30661=>"110111000",
  30662=>"110010111",
  30663=>"000000000",
  30664=>"000001101",
  30665=>"000100011",
  30666=>"000110100",
  30667=>"111010001",
  30668=>"011000111",
  30669=>"000111100",
  30670=>"001001000",
  30671=>"001010001",
  30672=>"110001001",
  30673=>"100100010",
  30674=>"111000110",
  30675=>"011101111",
  30676=>"000110111",
  30677=>"110010110",
  30678=>"110001101",
  30679=>"101110101",
  30680=>"010111010",
  30681=>"010100100",
  30682=>"010010110",
  30683=>"111010010",
  30684=>"001100101",
  30685=>"110000100",
  30686=>"111000110",
  30687=>"110100101",
  30688=>"001101001",
  30689=>"000001000",
  30690=>"010101101",
  30691=>"000000000",
  30692=>"110101011",
  30693=>"101101010",
  30694=>"111101000",
  30695=>"000101101",
  30696=>"101000000",
  30697=>"111100000",
  30698=>"001000110",
  30699=>"011010101",
  30700=>"101111110",
  30701=>"001101001",
  30702=>"100001011",
  30703=>"101001111",
  30704=>"000101000",
  30705=>"011010011",
  30706=>"100011111",
  30707=>"010001110",
  30708=>"100111110",
  30709=>"110010100",
  30710=>"000011111",
  30711=>"001101011",
  30712=>"100010011",
  30713=>"011100111",
  30714=>"001110110",
  30715=>"000111011",
  30716=>"010000000",
  30717=>"000001101",
  30718=>"010001100",
  30719=>"000111011",
  30720=>"111001001",
  30721=>"101000001",
  30722=>"011100100",
  30723=>"011001100",
  30724=>"000000101",
  30725=>"100010000",
  30726=>"111100101",
  30727=>"101111111",
  30728=>"111000001",
  30729=>"111001111",
  30730=>"001110001",
  30731=>"111000010",
  30732=>"000010110",
  30733=>"000111101",
  30734=>"011111000",
  30735=>"001011100",
  30736=>"111000001",
  30737=>"100000100",
  30738=>"111110000",
  30739=>"000000001",
  30740=>"001000100",
  30741=>"100011100",
  30742=>"100111001",
  30743=>"001110101",
  30744=>"100010110",
  30745=>"111110100",
  30746=>"010111110",
  30747=>"011111011",
  30748=>"001110011",
  30749=>"001100100",
  30750=>"000001001",
  30751=>"100111000",
  30752=>"101010001",
  30753=>"000110111",
  30754=>"001000111",
  30755=>"101100100",
  30756=>"011101101",
  30757=>"011101111",
  30758=>"101000000",
  30759=>"111100110",
  30760=>"111010011",
  30761=>"011111001",
  30762=>"111101111",
  30763=>"111010100",
  30764=>"011101000",
  30765=>"101110110",
  30766=>"100011001",
  30767=>"111110011",
  30768=>"110110010",
  30769=>"001100011",
  30770=>"111001011",
  30771=>"111110000",
  30772=>"000100111",
  30773=>"110111101",
  30774=>"000000101",
  30775=>"000111111",
  30776=>"000000001",
  30777=>"101100001",
  30778=>"010000000",
  30779=>"000001110",
  30780=>"010010000",
  30781=>"110000000",
  30782=>"111111110",
  30783=>"111110111",
  30784=>"010001011",
  30785=>"010100001",
  30786=>"000011100",
  30787=>"101101111",
  30788=>"101011000",
  30789=>"111011001",
  30790=>"011101011",
  30791=>"110100011",
  30792=>"100000100",
  30793=>"110011010",
  30794=>"010011000",
  30795=>"111110110",
  30796=>"111110010",
  30797=>"101001011",
  30798=>"011001010",
  30799=>"010100001",
  30800=>"001101100",
  30801=>"010010101",
  30802=>"000111010",
  30803=>"001100111",
  30804=>"001000100",
  30805=>"000110011",
  30806=>"000011111",
  30807=>"110010000",
  30808=>"010110111",
  30809=>"100111001",
  30810=>"111011101",
  30811=>"000000001",
  30812=>"100000101",
  30813=>"101101011",
  30814=>"011000001",
  30815=>"011110001",
  30816=>"000010011",
  30817=>"010101110",
  30818=>"111011010",
  30819=>"000010010",
  30820=>"000001001",
  30821=>"101010101",
  30822=>"100010110",
  30823=>"001110110",
  30824=>"101101001",
  30825=>"100011110",
  30826=>"010011010",
  30827=>"010100100",
  30828=>"010100100",
  30829=>"010111000",
  30830=>"010101110",
  30831=>"100011100",
  30832=>"001001001",
  30833=>"101011001",
  30834=>"110111110",
  30835=>"100100011",
  30836=>"011111101",
  30837=>"111110000",
  30838=>"110011001",
  30839=>"100110010",
  30840=>"010101101",
  30841=>"011111111",
  30842=>"011010110",
  30843=>"010001001",
  30844=>"110010001",
  30845=>"000100000",
  30846=>"010110001",
  30847=>"101101111",
  30848=>"000000110",
  30849=>"111100000",
  30850=>"101101100",
  30851=>"001011010",
  30852=>"001100101",
  30853=>"010101010",
  30854=>"100111110",
  30855=>"100010111",
  30856=>"001001011",
  30857=>"001010110",
  30858=>"010110110",
  30859=>"010110101",
  30860=>"011001101",
  30861=>"001011110",
  30862=>"110001011",
  30863=>"111110111",
  30864=>"011010001",
  30865=>"100000010",
  30866=>"110011001",
  30867=>"111000000",
  30868=>"100111110",
  30869=>"101011100",
  30870=>"010010110",
  30871=>"000111100",
  30872=>"101101001",
  30873=>"101110010",
  30874=>"011000111",
  30875=>"000110110",
  30876=>"011111100",
  30877=>"000010000",
  30878=>"011000110",
  30879=>"111001110",
  30880=>"101110010",
  30881=>"010000010",
  30882=>"111011011",
  30883=>"111000101",
  30884=>"001001111",
  30885=>"110000001",
  30886=>"101000000",
  30887=>"010101001",
  30888=>"010111010",
  30889=>"001011100",
  30890=>"000110010",
  30891=>"101000000",
  30892=>"000010100",
  30893=>"111101110",
  30894=>"010101001",
  30895=>"110000110",
  30896=>"100010000",
  30897=>"110011100",
  30898=>"101111111",
  30899=>"010000111",
  30900=>"001110111",
  30901=>"100111110",
  30902=>"000001010",
  30903=>"111011011",
  30904=>"000010010",
  30905=>"001110111",
  30906=>"100110111",
  30907=>"100111011",
  30908=>"100011000",
  30909=>"010110010",
  30910=>"010010111",
  30911=>"001110101",
  30912=>"000110100",
  30913=>"011011110",
  30914=>"110111000",
  30915=>"101101110",
  30916=>"110011001",
  30917=>"011110011",
  30918=>"100100011",
  30919=>"111110110",
  30920=>"110000010",
  30921=>"101010000",
  30922=>"011111001",
  30923=>"100110000",
  30924=>"000000011",
  30925=>"010111011",
  30926=>"110000101",
  30927=>"000000110",
  30928=>"001110000",
  30929=>"001101010",
  30930=>"010110001",
  30931=>"101101000",
  30932=>"101000100",
  30933=>"000110100",
  30934=>"111001111",
  30935=>"100000101",
  30936=>"110001010",
  30937=>"101100000",
  30938=>"100101101",
  30939=>"001111101",
  30940=>"011000000",
  30941=>"011111010",
  30942=>"000010110",
  30943=>"010000000",
  30944=>"111000111",
  30945=>"110101111",
  30946=>"001010111",
  30947=>"010101011",
  30948=>"101111111",
  30949=>"111110000",
  30950=>"101011010",
  30951=>"101100010",
  30952=>"111100011",
  30953=>"010010011",
  30954=>"110001100",
  30955=>"101010100",
  30956=>"100110000",
  30957=>"010011110",
  30958=>"111001000",
  30959=>"101101111",
  30960=>"011000111",
  30961=>"001110001",
  30962=>"000111111",
  30963=>"001011010",
  30964=>"101111011",
  30965=>"111001111",
  30966=>"110001010",
  30967=>"100111000",
  30968=>"000010100",
  30969=>"011100111",
  30970=>"101111011",
  30971=>"100001011",
  30972=>"011101110",
  30973=>"000100110",
  30974=>"101001110",
  30975=>"000011100",
  30976=>"101100001",
  30977=>"110101101",
  30978=>"100011110",
  30979=>"011011011",
  30980=>"111101000",
  30981=>"101111011",
  30982=>"000010001",
  30983=>"110000000",
  30984=>"011001111",
  30985=>"100011001",
  30986=>"010001111",
  30987=>"100010110",
  30988=>"110000110",
  30989=>"110000000",
  30990=>"000111100",
  30991=>"001111010",
  30992=>"110100001",
  30993=>"010110010",
  30994=>"100010010",
  30995=>"111101100",
  30996=>"100001011",
  30997=>"101110001",
  30998=>"001110010",
  30999=>"000000111",
  31000=>"110100000",
  31001=>"101100001",
  31002=>"011000011",
  31003=>"110100001",
  31004=>"010001100",
  31005=>"110111110",
  31006=>"101100111",
  31007=>"001101011",
  31008=>"101001000",
  31009=>"011010100",
  31010=>"001100001",
  31011=>"101100100",
  31012=>"001000011",
  31013=>"100100000",
  31014=>"100001000",
  31015=>"010101010",
  31016=>"110001111",
  31017=>"101110101",
  31018=>"001111011",
  31019=>"111100111",
  31020=>"100010011",
  31021=>"100011011",
  31022=>"110101010",
  31023=>"011010001",
  31024=>"100011100",
  31025=>"011111001",
  31026=>"101000010",
  31027=>"001111010",
  31028=>"101110010",
  31029=>"011111100",
  31030=>"101011011",
  31031=>"011110101",
  31032=>"110010010",
  31033=>"000011000",
  31034=>"011111011",
  31035=>"111010000",
  31036=>"101101111",
  31037=>"101101111",
  31038=>"101111100",
  31039=>"000011110",
  31040=>"101011010",
  31041=>"100111010",
  31042=>"111010110",
  31043=>"011000000",
  31044=>"011010100",
  31045=>"010111001",
  31046=>"010000011",
  31047=>"000110001",
  31048=>"110010100",
  31049=>"010110000",
  31050=>"100010001",
  31051=>"110011111",
  31052=>"000011110",
  31053=>"011111011",
  31054=>"000010001",
  31055=>"001111100",
  31056=>"000100000",
  31057=>"000110100",
  31058=>"011010100",
  31059=>"111011010",
  31060=>"001000101",
  31061=>"000101000",
  31062=>"111011010",
  31063=>"100110001",
  31064=>"000010000",
  31065=>"100000110",
  31066=>"110000000",
  31067=>"101010001",
  31068=>"001000110",
  31069=>"010000001",
  31070=>"111100010",
  31071=>"100001010",
  31072=>"011110011",
  31073=>"100010101",
  31074=>"010000001",
  31075=>"000011011",
  31076=>"111001000",
  31077=>"001100111",
  31078=>"101110101",
  31079=>"110101000",
  31080=>"110000100",
  31081=>"100000010",
  31082=>"010110000",
  31083=>"011011001",
  31084=>"001110101",
  31085=>"001000100",
  31086=>"001000001",
  31087=>"100110000",
  31088=>"100001111",
  31089=>"011010100",
  31090=>"100101111",
  31091=>"000000100",
  31092=>"000001001",
  31093=>"001100011",
  31094=>"011110100",
  31095=>"111011101",
  31096=>"100000010",
  31097=>"011000110",
  31098=>"100100010",
  31099=>"100110111",
  31100=>"011001001",
  31101=>"110011010",
  31102=>"111111100",
  31103=>"000101011",
  31104=>"100011111",
  31105=>"001010000",
  31106=>"100001000",
  31107=>"100100110",
  31108=>"100111000",
  31109=>"101110010",
  31110=>"000001111",
  31111=>"010010000",
  31112=>"100000010",
  31113=>"000000110",
  31114=>"110010110",
  31115=>"000101001",
  31116=>"111111000",
  31117=>"000111000",
  31118=>"100011101",
  31119=>"100000011",
  31120=>"100010001",
  31121=>"001011010",
  31122=>"001000000",
  31123=>"110110110",
  31124=>"111110110",
  31125=>"001110110",
  31126=>"011011110",
  31127=>"000001010",
  31128=>"011011110",
  31129=>"100000010",
  31130=>"101010001",
  31131=>"011101111",
  31132=>"111010010",
  31133=>"111111101",
  31134=>"000101010",
  31135=>"000010110",
  31136=>"011011001",
  31137=>"111110110",
  31138=>"011001001",
  31139=>"010010011",
  31140=>"101001010",
  31141=>"000011010",
  31142=>"010000010",
  31143=>"100010010",
  31144=>"001110001",
  31145=>"001001010",
  31146=>"000110000",
  31147=>"010000101",
  31148=>"111101101",
  31149=>"111111111",
  31150=>"011111100",
  31151=>"010000001",
  31152=>"000001101",
  31153=>"010100110",
  31154=>"111111100",
  31155=>"111000001",
  31156=>"011111111",
  31157=>"001010000",
  31158=>"000011111",
  31159=>"001000000",
  31160=>"110111010",
  31161=>"000001100",
  31162=>"010100000",
  31163=>"101000111",
  31164=>"001011101",
  31165=>"101101000",
  31166=>"010101000",
  31167=>"000000000",
  31168=>"010010011",
  31169=>"011010110",
  31170=>"101110101",
  31171=>"101000110",
  31172=>"101000010",
  31173=>"100110010",
  31174=>"100011100",
  31175=>"111110001",
  31176=>"110011011",
  31177=>"010101111",
  31178=>"101011010",
  31179=>"000110000",
  31180=>"100111001",
  31181=>"100000000",
  31182=>"110010110",
  31183=>"110110000",
  31184=>"111000100",
  31185=>"000100101",
  31186=>"101110001",
  31187=>"111000101",
  31188=>"111000000",
  31189=>"011011110",
  31190=>"111111010",
  31191=>"010011100",
  31192=>"000000001",
  31193=>"101011010",
  31194=>"110110101",
  31195=>"111100000",
  31196=>"011001101",
  31197=>"100010010",
  31198=>"110100100",
  31199=>"111110110",
  31200=>"110011111",
  31201=>"101110100",
  31202=>"111011111",
  31203=>"110001110",
  31204=>"100100010",
  31205=>"111110010",
  31206=>"000100001",
  31207=>"100101110",
  31208=>"000110001",
  31209=>"111110001",
  31210=>"110010101",
  31211=>"110010001",
  31212=>"000001101",
  31213=>"010101100",
  31214=>"001100101",
  31215=>"010111000",
  31216=>"110100100",
  31217=>"111000011",
  31218=>"010011111",
  31219=>"011011101",
  31220=>"001111110",
  31221=>"111101110",
  31222=>"011101101",
  31223=>"011000101",
  31224=>"111111111",
  31225=>"001010000",
  31226=>"001101111",
  31227=>"101000001",
  31228=>"011000110",
  31229=>"011101110",
  31230=>"011000010",
  31231=>"000000010",
  31232=>"100000100",
  31233=>"011100000",
  31234=>"100101111",
  31235=>"100001000",
  31236=>"100100101",
  31237=>"010100001",
  31238=>"111011101",
  31239=>"110100001",
  31240=>"000111101",
  31241=>"001010001",
  31242=>"000011110",
  31243=>"101101101",
  31244=>"011001101",
  31245=>"010000000",
  31246=>"000011100",
  31247=>"101000101",
  31248=>"100110111",
  31249=>"010110111",
  31250=>"111111111",
  31251=>"101110001",
  31252=>"000101111",
  31253=>"011100001",
  31254=>"111010011",
  31255=>"010100011",
  31256=>"010110011",
  31257=>"110001000",
  31258=>"110011111",
  31259=>"101101001",
  31260=>"000000001",
  31261=>"010101011",
  31262=>"110110111",
  31263=>"010011000",
  31264=>"111110110",
  31265=>"111011110",
  31266=>"101000000",
  31267=>"001110010",
  31268=>"101111000",
  31269=>"111010011",
  31270=>"000110000",
  31271=>"000111111",
  31272=>"100101100",
  31273=>"010110010",
  31274=>"110111001",
  31275=>"011101001",
  31276=>"110000110",
  31277=>"111110001",
  31278=>"100101010",
  31279=>"110100010",
  31280=>"000010111",
  31281=>"011010001",
  31282=>"010101000",
  31283=>"000100110",
  31284=>"010111101",
  31285=>"000011110",
  31286=>"111011011",
  31287=>"011110101",
  31288=>"100001110",
  31289=>"001100000",
  31290=>"100111110",
  31291=>"111100111",
  31292=>"000101101",
  31293=>"000000000",
  31294=>"011000001",
  31295=>"011010110",
  31296=>"100101110",
  31297=>"111010101",
  31298=>"011011100",
  31299=>"111111000",
  31300=>"100011110",
  31301=>"110101000",
  31302=>"010100101",
  31303=>"101100001",
  31304=>"100100010",
  31305=>"110010101",
  31306=>"111010101",
  31307=>"010000000",
  31308=>"101101110",
  31309=>"101011000",
  31310=>"011100100",
  31311=>"011100111",
  31312=>"000110011",
  31313=>"100101000",
  31314=>"010101110",
  31315=>"001110100",
  31316=>"000000011",
  31317=>"011001101",
  31318=>"000001001",
  31319=>"110111111",
  31320=>"000000010",
  31321=>"100110011",
  31322=>"000111110",
  31323=>"010100010",
  31324=>"011110001",
  31325=>"010110000",
  31326=>"100010000",
  31327=>"000010001",
  31328=>"111110111",
  31329=>"000110011",
  31330=>"010101110",
  31331=>"100111001",
  31332=>"001001000",
  31333=>"100100101",
  31334=>"000111110",
  31335=>"001001000",
  31336=>"000000111",
  31337=>"011111101",
  31338=>"101111010",
  31339=>"000010100",
  31340=>"000101111",
  31341=>"110110011",
  31342=>"000011100",
  31343=>"101001111",
  31344=>"010001001",
  31345=>"011010011",
  31346=>"010100011",
  31347=>"100110111",
  31348=>"101101000",
  31349=>"010001110",
  31350=>"000101000",
  31351=>"101011011",
  31352=>"010110000",
  31353=>"000101101",
  31354=>"101111011",
  31355=>"110000101",
  31356=>"100110001",
  31357=>"101101110",
  31358=>"110011100",
  31359=>"110111010",
  31360=>"000101100",
  31361=>"111101010",
  31362=>"101111110",
  31363=>"011001100",
  31364=>"010101001",
  31365=>"000100100",
  31366=>"100110111",
  31367=>"101110100",
  31368=>"111111111",
  31369=>"010000101",
  31370=>"110001100",
  31371=>"000110001",
  31372=>"100100000",
  31373=>"000010100",
  31374=>"110100000",
  31375=>"111000010",
  31376=>"111001111",
  31377=>"111011001",
  31378=>"110000001",
  31379=>"011111111",
  31380=>"001100101",
  31381=>"010010101",
  31382=>"111111001",
  31383=>"110111011",
  31384=>"011001100",
  31385=>"111110011",
  31386=>"110111001",
  31387=>"111000011",
  31388=>"101101111",
  31389=>"010110001",
  31390=>"000011111",
  31391=>"011110100",
  31392=>"110001010",
  31393=>"000001000",
  31394=>"100110000",
  31395=>"011100111",
  31396=>"000010110",
  31397=>"001110110",
  31398=>"001110001",
  31399=>"010000001",
  31400=>"111001101",
  31401=>"100000111",
  31402=>"001111000",
  31403=>"110000001",
  31404=>"110010000",
  31405=>"000000000",
  31406=>"010011101",
  31407=>"001101011",
  31408=>"000000110",
  31409=>"000001111",
  31410=>"000010011",
  31411=>"110101111",
  31412=>"011001100",
  31413=>"100111110",
  31414=>"110001000",
  31415=>"010000101",
  31416=>"101011000",
  31417=>"110001010",
  31418=>"100101001",
  31419=>"100000100",
  31420=>"100011010",
  31421=>"111110010",
  31422=>"011000000",
  31423=>"100101100",
  31424=>"111101110",
  31425=>"101000101",
  31426=>"010010101",
  31427=>"000101001",
  31428=>"110011111",
  31429=>"010110001",
  31430=>"111001010",
  31431=>"100101000",
  31432=>"010101100",
  31433=>"001010101",
  31434=>"011011001",
  31435=>"010100110",
  31436=>"010101001",
  31437=>"110011100",
  31438=>"101110100",
  31439=>"000010100",
  31440=>"111111101",
  31441=>"001010110",
  31442=>"101011111",
  31443=>"010000001",
  31444=>"011111101",
  31445=>"100111110",
  31446=>"001001001",
  31447=>"010100100",
  31448=>"110111110",
  31449=>"101110111",
  31450=>"110010110",
  31451=>"110110001",
  31452=>"010111101",
  31453=>"010110100",
  31454=>"100001010",
  31455=>"100110001",
  31456=>"101100110",
  31457=>"010000000",
  31458=>"010011110",
  31459=>"101111001",
  31460=>"101100010",
  31461=>"001101001",
  31462=>"111100000",
  31463=>"000001100",
  31464=>"000010000",
  31465=>"111101000",
  31466=>"111110010",
  31467=>"011001111",
  31468=>"010001010",
  31469=>"100010110",
  31470=>"100001110",
  31471=>"111111101",
  31472=>"111111111",
  31473=>"101000011",
  31474=>"101001110",
  31475=>"000110101",
  31476=>"000101100",
  31477=>"001100101",
  31478=>"111110111",
  31479=>"110010000",
  31480=>"001101000",
  31481=>"101110011",
  31482=>"100111011",
  31483=>"100001011",
  31484=>"101100111",
  31485=>"100010001",
  31486=>"010101011",
  31487=>"101010010",
  31488=>"000001101",
  31489=>"111110010",
  31490=>"101110001",
  31491=>"111101110",
  31492=>"000110110",
  31493=>"001001111",
  31494=>"101111011",
  31495=>"010000100",
  31496=>"110110100",
  31497=>"100001010",
  31498=>"100100110",
  31499=>"000000000",
  31500=>"100010001",
  31501=>"100001110",
  31502=>"111100011",
  31503=>"101100101",
  31504=>"000100100",
  31505=>"010100010",
  31506=>"101011000",
  31507=>"000001001",
  31508=>"001011001",
  31509=>"001000001",
  31510=>"010010101",
  31511=>"000110111",
  31512=>"001011001",
  31513=>"011100000",
  31514=>"000001100",
  31515=>"110011010",
  31516=>"010110110",
  31517=>"011001110",
  31518=>"000110101",
  31519=>"000010110",
  31520=>"011011100",
  31521=>"100110101",
  31522=>"000101011",
  31523=>"011110101",
  31524=>"010100101",
  31525=>"011011110",
  31526=>"100011011",
  31527=>"001011100",
  31528=>"101101000",
  31529=>"000011011",
  31530=>"110011110",
  31531=>"001111001",
  31532=>"000010111",
  31533=>"100000001",
  31534=>"011010011",
  31535=>"101000110",
  31536=>"000110001",
  31537=>"110001011",
  31538=>"010011000",
  31539=>"111100100",
  31540=>"000100010",
  31541=>"101010111",
  31542=>"011011110",
  31543=>"000000000",
  31544=>"001101011",
  31545=>"010000011",
  31546=>"000000011",
  31547=>"111000010",
  31548=>"110000011",
  31549=>"000000001",
  31550=>"110000001",
  31551=>"001001110",
  31552=>"010100100",
  31553=>"111111011",
  31554=>"110101001",
  31555=>"010010010",
  31556=>"111000101",
  31557=>"011100011",
  31558=>"100101010",
  31559=>"000111011",
  31560=>"110100000",
  31561=>"100000010",
  31562=>"100011000",
  31563=>"010101000",
  31564=>"010100100",
  31565=>"110010111",
  31566=>"001010011",
  31567=>"000001001",
  31568=>"000100010",
  31569=>"011100110",
  31570=>"000100100",
  31571=>"111100111",
  31572=>"111000001",
  31573=>"110001011",
  31574=>"011010100",
  31575=>"110010001",
  31576=>"001101011",
  31577=>"101111010",
  31578=>"000000010",
  31579=>"110001000",
  31580=>"110000011",
  31581=>"111011111",
  31582=>"111110001",
  31583=>"011111101",
  31584=>"100010011",
  31585=>"100110011",
  31586=>"111001010",
  31587=>"100111000",
  31588=>"100000110",
  31589=>"101011001",
  31590=>"111001111",
  31591=>"000101111",
  31592=>"001011001",
  31593=>"001000101",
  31594=>"111001010",
  31595=>"101110000",
  31596=>"110111011",
  31597=>"111001111",
  31598=>"011010011",
  31599=>"101110110",
  31600=>"011100010",
  31601=>"011101010",
  31602=>"100010000",
  31603=>"101111001",
  31604=>"111010000",
  31605=>"010100110",
  31606=>"010101110",
  31607=>"001111100",
  31608=>"011111100",
  31609=>"101110111",
  31610=>"000101111",
  31611=>"111011100",
  31612=>"111110010",
  31613=>"100010111",
  31614=>"011100001",
  31615=>"000110101",
  31616=>"111100111",
  31617=>"011101110",
  31618=>"111011101",
  31619=>"111110000",
  31620=>"101101111",
  31621=>"001100010",
  31622=>"111011011",
  31623=>"000010010",
  31624=>"100111001",
  31625=>"100000111",
  31626=>"110110000",
  31627=>"010110111",
  31628=>"000011011",
  31629=>"011000000",
  31630=>"101001011",
  31631=>"011011111",
  31632=>"001110000",
  31633=>"110111111",
  31634=>"010001000",
  31635=>"010110010",
  31636=>"111100001",
  31637=>"110001011",
  31638=>"100011101",
  31639=>"011010110",
  31640=>"011101111",
  31641=>"111110101",
  31642=>"110100001",
  31643=>"100010001",
  31644=>"111001001",
  31645=>"001001011",
  31646=>"100001011",
  31647=>"111101001",
  31648=>"110010010",
  31649=>"001010100",
  31650=>"111011101",
  31651=>"100111100",
  31652=>"111010011",
  31653=>"000011010",
  31654=>"110000010",
  31655=>"101000001",
  31656=>"000111010",
  31657=>"100010010",
  31658=>"101000100",
  31659=>"000101010",
  31660=>"010110011",
  31661=>"101101111",
  31662=>"111000000",
  31663=>"011001011",
  31664=>"000001110",
  31665=>"110111010",
  31666=>"101100010",
  31667=>"000000010",
  31668=>"010100011",
  31669=>"010001011",
  31670=>"001111100",
  31671=>"101001011",
  31672=>"001000010",
  31673=>"100101010",
  31674=>"101001100",
  31675=>"010000100",
  31676=>"000100001",
  31677=>"011110011",
  31678=>"011111100",
  31679=>"011100101",
  31680=>"110011111",
  31681=>"000101010",
  31682=>"011101111",
  31683=>"001111100",
  31684=>"100000011",
  31685=>"101110111",
  31686=>"111010011",
  31687=>"110000111",
  31688=>"111011001",
  31689=>"001111111",
  31690=>"100001110",
  31691=>"101001111",
  31692=>"111001111",
  31693=>"101011001",
  31694=>"111101101",
  31695=>"101110100",
  31696=>"110000110",
  31697=>"000001010",
  31698=>"110101000",
  31699=>"110001100",
  31700=>"000110101",
  31701=>"100000111",
  31702=>"111110000",
  31703=>"111000011",
  31704=>"110011101",
  31705=>"000100000",
  31706=>"100001001",
  31707=>"011001010",
  31708=>"001110100",
  31709=>"000001101",
  31710=>"001010111",
  31711=>"000000111",
  31712=>"111010100",
  31713=>"111011110",
  31714=>"011001101",
  31715=>"101000000",
  31716=>"000111011",
  31717=>"011000011",
  31718=>"101100110",
  31719=>"110001001",
  31720=>"010010100",
  31721=>"101000010",
  31722=>"111111111",
  31723=>"101111011",
  31724=>"011101000",
  31725=>"100111110",
  31726=>"011010101",
  31727=>"011011110",
  31728=>"100110101",
  31729=>"111101111",
  31730=>"001010010",
  31731=>"111101001",
  31732=>"101011001",
  31733=>"110001010",
  31734=>"101011011",
  31735=>"010100011",
  31736=>"111010101",
  31737=>"111011010",
  31738=>"101001111",
  31739=>"100111001",
  31740=>"011010111",
  31741=>"011001011",
  31742=>"111101001",
  31743=>"000111010",
  31744=>"101000111",
  31745=>"000101010",
  31746=>"000001011",
  31747=>"101011101",
  31748=>"011111110",
  31749=>"000100010",
  31750=>"010010010",
  31751=>"110001001",
  31752=>"011101100",
  31753=>"001101110",
  31754=>"010000010",
  31755=>"101101111",
  31756=>"011110101",
  31757=>"011110111",
  31758=>"010011111",
  31759=>"100010001",
  31760=>"011010100",
  31761=>"101101011",
  31762=>"000010101",
  31763=>"101010010",
  31764=>"001101010",
  31765=>"011100010",
  31766=>"110011000",
  31767=>"100111001",
  31768=>"011111010",
  31769=>"110101010",
  31770=>"110011000",
  31771=>"110011001",
  31772=>"110000000",
  31773=>"001101101",
  31774=>"000111001",
  31775=>"101101111",
  31776=>"010110101",
  31777=>"001110101",
  31778=>"100001000",
  31779=>"101100110",
  31780=>"101001001",
  31781=>"010011101",
  31782=>"001011100",
  31783=>"001100101",
  31784=>"111011011",
  31785=>"100111011",
  31786=>"110100100",
  31787=>"111110000",
  31788=>"000100011",
  31789=>"101111100",
  31790=>"110010101",
  31791=>"011000001",
  31792=>"010111101",
  31793=>"001001100",
  31794=>"001100111",
  31795=>"000001101",
  31796=>"100010111",
  31797=>"101000111",
  31798=>"111010001",
  31799=>"000010100",
  31800=>"110110011",
  31801=>"110000110",
  31802=>"101000100",
  31803=>"110010101",
  31804=>"011100001",
  31805=>"101000010",
  31806=>"001101100",
  31807=>"101100101",
  31808=>"110110111",
  31809=>"010000001",
  31810=>"000110010",
  31811=>"001000011",
  31812=>"110010000",
  31813=>"100010000",
  31814=>"001001101",
  31815=>"011100011",
  31816=>"101111111",
  31817=>"111010100",
  31818=>"000101010",
  31819=>"001000011",
  31820=>"010111011",
  31821=>"101101000",
  31822=>"011000111",
  31823=>"011100011",
  31824=>"101111100",
  31825=>"001111111",
  31826=>"111011111",
  31827=>"111111000",
  31828=>"011100100",
  31829=>"111101101",
  31830=>"100000111",
  31831=>"000110011",
  31832=>"111111101",
  31833=>"100110100",
  31834=>"100111100",
  31835=>"101001001",
  31836=>"111010001",
  31837=>"000100101",
  31838=>"010101011",
  31839=>"011101100",
  31840=>"000010001",
  31841=>"110001100",
  31842=>"001111100",
  31843=>"100111110",
  31844=>"010000010",
  31845=>"000111110",
  31846=>"001000011",
  31847=>"010100100",
  31848=>"000010101",
  31849=>"111111010",
  31850=>"001001011",
  31851=>"101010000",
  31852=>"010001111",
  31853=>"100110110",
  31854=>"011101100",
  31855=>"000000001",
  31856=>"010110011",
  31857=>"011000000",
  31858=>"010001100",
  31859=>"100110011",
  31860=>"110100110",
  31861=>"100000010",
  31862=>"100100110",
  31863=>"101101101",
  31864=>"100100001",
  31865=>"100000101",
  31866=>"101111110",
  31867=>"100011011",
  31868=>"111110110",
  31869=>"000111111",
  31870=>"111001001",
  31871=>"110011110",
  31872=>"100011101",
  31873=>"010111111",
  31874=>"111001100",
  31875=>"100001010",
  31876=>"111001010",
  31877=>"011101011",
  31878=>"011110111",
  31879=>"000100010",
  31880=>"100100100",
  31881=>"010011010",
  31882=>"101000011",
  31883=>"101001100",
  31884=>"110100000",
  31885=>"111101000",
  31886=>"111000000",
  31887=>"011001101",
  31888=>"101010111",
  31889=>"101111101",
  31890=>"000100111",
  31891=>"111001001",
  31892=>"001001010",
  31893=>"100111001",
  31894=>"110001101",
  31895=>"100101111",
  31896=>"110010001",
  31897=>"111100100",
  31898=>"001000100",
  31899=>"011110111",
  31900=>"000001110",
  31901=>"111110010",
  31902=>"100101000",
  31903=>"111001101",
  31904=>"010101010",
  31905=>"011101010",
  31906=>"100110110",
  31907=>"001111011",
  31908=>"100100101",
  31909=>"100111010",
  31910=>"110011110",
  31911=>"010110011",
  31912=>"101111111",
  31913=>"001010011",
  31914=>"011111110",
  31915=>"111000001",
  31916=>"111111011",
  31917=>"000011101",
  31918=>"110110001",
  31919=>"011000101",
  31920=>"101010111",
  31921=>"100110100",
  31922=>"010100001",
  31923=>"000001100",
  31924=>"100100110",
  31925=>"111110000",
  31926=>"111011111",
  31927=>"010111001",
  31928=>"000101110",
  31929=>"111010000",
  31930=>"011100000",
  31931=>"010110011",
  31932=>"101001011",
  31933=>"011011110",
  31934=>"001001001",
  31935=>"101110001",
  31936=>"000110110",
  31937=>"001100000",
  31938=>"000101110",
  31939=>"111100000",
  31940=>"011001001",
  31941=>"001100001",
  31942=>"111001001",
  31943=>"101101110",
  31944=>"010011011",
  31945=>"111111011",
  31946=>"000110111",
  31947=>"000110000",
  31948=>"101000010",
  31949=>"100100100",
  31950=>"010101101",
  31951=>"001010001",
  31952=>"111110100",
  31953=>"000000010",
  31954=>"111001010",
  31955=>"101010111",
  31956=>"101000010",
  31957=>"100010001",
  31958=>"101011111",
  31959=>"110011110",
  31960=>"111101101",
  31961=>"011010111",
  31962=>"101100110",
  31963=>"100111011",
  31964=>"000111111",
  31965=>"110110001",
  31966=>"100111110",
  31967=>"010000001",
  31968=>"000000111",
  31969=>"101010100",
  31970=>"001001111",
  31971=>"111010100",
  31972=>"111001001",
  31973=>"010110000",
  31974=>"111111000",
  31975=>"000110111",
  31976=>"011000000",
  31977=>"001100100",
  31978=>"001011101",
  31979=>"110010001",
  31980=>"101101000",
  31981=>"001001010",
  31982=>"000101011",
  31983=>"001100001",
  31984=>"010110101",
  31985=>"100100001",
  31986=>"100101101",
  31987=>"111110100",
  31988=>"000111110",
  31989=>"010100101",
  31990=>"100011010",
  31991=>"111111001",
  31992=>"110011010",
  31993=>"101111100",
  31994=>"000001100",
  31995=>"110000001",
  31996=>"111101001",
  31997=>"000111010",
  31998=>"110001110",
  31999=>"001111110",
  32000=>"101110101",
  32001=>"001101100",
  32002=>"101101111",
  32003=>"010100001",
  32004=>"100011001",
  32005=>"101010111",
  32006=>"110011110",
  32007=>"110100111",
  32008=>"010010010",
  32009=>"100001001",
  32010=>"110110010",
  32011=>"100111101",
  32012=>"000010110",
  32013=>"011010011",
  32014=>"010101111",
  32015=>"111010100",
  32016=>"111101001",
  32017=>"110000111",
  32018=>"000010100",
  32019=>"010000001",
  32020=>"010101011",
  32021=>"001010110",
  32022=>"010011000",
  32023=>"001101101",
  32024=>"111111101",
  32025=>"111100100",
  32026=>"101001111",
  32027=>"111110010",
  32028=>"100110111",
  32029=>"100101011",
  32030=>"011011010",
  32031=>"100000001",
  32032=>"110001101",
  32033=>"001000010",
  32034=>"111000101",
  32035=>"011010111",
  32036=>"010000101",
  32037=>"111101111",
  32038=>"101011110",
  32039=>"110010000",
  32040=>"101110101",
  32041=>"001110101",
  32042=>"111011110",
  32043=>"101101101",
  32044=>"011010111",
  32045=>"111101111",
  32046=>"110000100",
  32047=>"011110110",
  32048=>"111110000",
  32049=>"001111100",
  32050=>"110100000",
  32051=>"010010011",
  32052=>"111101011",
  32053=>"001000101",
  32054=>"001001100",
  32055=>"100110111",
  32056=>"000101000",
  32057=>"001101110",
  32058=>"100001101",
  32059=>"000000000",
  32060=>"011011011",
  32061=>"110001110",
  32062=>"101001000",
  32063=>"110000110",
  32064=>"000001100",
  32065=>"101010010",
  32066=>"010100100",
  32067=>"100011001",
  32068=>"100011101",
  32069=>"011011101",
  32070=>"100001001",
  32071=>"001101001",
  32072=>"100011000",
  32073=>"101100000",
  32074=>"111010111",
  32075=>"010001001",
  32076=>"101011011",
  32077=>"000101001",
  32078=>"000110111",
  32079=>"011100010",
  32080=>"000101101",
  32081=>"100000111",
  32082=>"110100111",
  32083=>"000001010",
  32084=>"010101010",
  32085=>"001101001",
  32086=>"001001101",
  32087=>"111111010",
  32088=>"011010010",
  32089=>"101011111",
  32090=>"101000011",
  32091=>"001000100",
  32092=>"101010101",
  32093=>"101010010",
  32094=>"010010100",
  32095=>"100001001",
  32096=>"000010100",
  32097=>"101011011",
  32098=>"111101011",
  32099=>"011111111",
  32100=>"111110111",
  32101=>"001011010",
  32102=>"011100000",
  32103=>"100000001",
  32104=>"001001111",
  32105=>"111110010",
  32106=>"100100000",
  32107=>"011101100",
  32108=>"100010000",
  32109=>"010100100",
  32110=>"101011001",
  32111=>"010011111",
  32112=>"110101011",
  32113=>"001111100",
  32114=>"001001110",
  32115=>"101001000",
  32116=>"101101010",
  32117=>"001111111",
  32118=>"000011001",
  32119=>"100100001",
  32120=>"000011110",
  32121=>"000001101",
  32122=>"001000001",
  32123=>"100010100",
  32124=>"111000100",
  32125=>"101000000",
  32126=>"010001110",
  32127=>"111100111",
  32128=>"110100101",
  32129=>"000110010",
  32130=>"000101000",
  32131=>"011010010",
  32132=>"001110110",
  32133=>"101001110",
  32134=>"001111010",
  32135=>"110000100",
  32136=>"010110001",
  32137=>"011101011",
  32138=>"100010110",
  32139=>"110011110",
  32140=>"110110101",
  32141=>"100000001",
  32142=>"111100111",
  32143=>"101010010",
  32144=>"101000101",
  32145=>"111100001",
  32146=>"000010110",
  32147=>"010101011",
  32148=>"001010001",
  32149=>"110100101",
  32150=>"101011011",
  32151=>"100001010",
  32152=>"101110101",
  32153=>"111110101",
  32154=>"001101001",
  32155=>"101001111",
  32156=>"011101000",
  32157=>"110011101",
  32158=>"110010011",
  32159=>"011110010",
  32160=>"001110101",
  32161=>"011101010",
  32162=>"111010001",
  32163=>"010100110",
  32164=>"100100000",
  32165=>"101110000",
  32166=>"011001011",
  32167=>"100100011",
  32168=>"001111001",
  32169=>"110111011",
  32170=>"101010001",
  32171=>"100010000",
  32172=>"000100000",
  32173=>"010010010",
  32174=>"000000111",
  32175=>"010111011",
  32176=>"110101101",
  32177=>"000000001",
  32178=>"010011001",
  32179=>"111100011",
  32180=>"011001101",
  32181=>"111011101",
  32182=>"100001101",
  32183=>"100000001",
  32184=>"110000011",
  32185=>"011100100",
  32186=>"101001100",
  32187=>"010010101",
  32188=>"111010011",
  32189=>"000110000",
  32190=>"010100001",
  32191=>"110011011",
  32192=>"100001101",
  32193=>"111001000",
  32194=>"000010101",
  32195=>"001001110",
  32196=>"110110101",
  32197=>"001001111",
  32198=>"001110001",
  32199=>"100010101",
  32200=>"010111001",
  32201=>"000110000",
  32202=>"101001100",
  32203=>"101100110",
  32204=>"000101010",
  32205=>"000101000",
  32206=>"011111010",
  32207=>"100110011",
  32208=>"110101001",
  32209=>"110110001",
  32210=>"000001010",
  32211=>"111011111",
  32212=>"010110001",
  32213=>"010011100",
  32214=>"001111010",
  32215=>"101110011",
  32216=>"010011101",
  32217=>"011100010",
  32218=>"001000011",
  32219=>"000011011",
  32220=>"111111001",
  32221=>"010010000",
  32222=>"111111100",
  32223=>"101100010",
  32224=>"001111000",
  32225=>"111000100",
  32226=>"000011011",
  32227=>"000101100",
  32228=>"010111110",
  32229=>"010010100",
  32230=>"101010110",
  32231=>"001111100",
  32232=>"101101010",
  32233=>"000101100",
  32234=>"100010100",
  32235=>"000010011",
  32236=>"010100000",
  32237=>"101101100",
  32238=>"001010111",
  32239=>"001111000",
  32240=>"010011111",
  32241=>"011111110",
  32242=>"110100000",
  32243=>"101101010",
  32244=>"100111001",
  32245=>"000111111",
  32246=>"011010110",
  32247=>"110111100",
  32248=>"111011100",
  32249=>"101000011",
  32250=>"010110111",
  32251=>"010000110",
  32252=>"011111010",
  32253=>"001100000",
  32254=>"100101110",
  32255=>"110100111",
  32256=>"011101111",
  32257=>"000011101",
  32258=>"101110011",
  32259=>"001001101",
  32260=>"111110101",
  32261=>"111011000",
  32262=>"110000011",
  32263=>"100100010",
  32264=>"100111111",
  32265=>"000100111",
  32266=>"111010100",
  32267=>"110100011",
  32268=>"111111010",
  32269=>"001111111",
  32270=>"111101000",
  32271=>"011011100",
  32272=>"101111111",
  32273=>"011110111",
  32274=>"000000011",
  32275=>"100110110",
  32276=>"110001111",
  32277=>"010101010",
  32278=>"111000000",
  32279=>"100011001",
  32280=>"011101001",
  32281=>"000010000",
  32282=>"101001111",
  32283=>"001001001",
  32284=>"100111100",
  32285=>"110001010",
  32286=>"011101101",
  32287=>"001000011",
  32288=>"101101100",
  32289=>"111111001",
  32290=>"011000010",
  32291=>"111011001",
  32292=>"100101110",
  32293=>"000110111",
  32294=>"111100010",
  32295=>"000001101",
  32296=>"011010101",
  32297=>"000010111",
  32298=>"011001110",
  32299=>"110001011",
  32300=>"000010011",
  32301=>"110010011",
  32302=>"001001000",
  32303=>"011100101",
  32304=>"111100010",
  32305=>"100101101",
  32306=>"100000110",
  32307=>"000000001",
  32308=>"011011011",
  32309=>"111110111",
  32310=>"100000111",
  32311=>"001100100",
  32312=>"010010001",
  32313=>"101010100",
  32314=>"110011011",
  32315=>"101111000",
  32316=>"011001101",
  32317=>"011101111",
  32318=>"110001001",
  32319=>"000111111",
  32320=>"110110001",
  32321=>"011101111",
  32322=>"110001110",
  32323=>"010001001",
  32324=>"101001000",
  32325=>"101110100",
  32326=>"111111001",
  32327=>"111101010",
  32328=>"010000110",
  32329=>"110001001",
  32330=>"111100000",
  32331=>"100111000",
  32332=>"000100101",
  32333=>"100000011",
  32334=>"110011011",
  32335=>"010100011",
  32336=>"000100111",
  32337=>"000000000",
  32338=>"011001000",
  32339=>"001101101",
  32340=>"101000110",
  32341=>"101011101",
  32342=>"001111110",
  32343=>"001001000",
  32344=>"000010110",
  32345=>"011100111",
  32346=>"011110010",
  32347=>"001001001",
  32348=>"101001010",
  32349=>"110101010",
  32350=>"100000001",
  32351=>"110110111",
  32352=>"000111101",
  32353=>"011100001",
  32354=>"011011010",
  32355=>"011101001",
  32356=>"010000001",
  32357=>"000100111",
  32358=>"101010111",
  32359=>"111000101",
  32360=>"101101001",
  32361=>"001011110",
  32362=>"011111011",
  32363=>"111001000",
  32364=>"000111011",
  32365=>"011000011",
  32366=>"001110101",
  32367=>"100100001",
  32368=>"111101011",
  32369=>"011001000",
  32370=>"110111110",
  32371=>"011010101",
  32372=>"101010010",
  32373=>"101000000",
  32374=>"011010011",
  32375=>"111001111",
  32376=>"011111010",
  32377=>"100101011",
  32378=>"101110011",
  32379=>"010100011",
  32380=>"101011010",
  32381=>"001011101",
  32382=>"101001001",
  32383=>"100001001",
  32384=>"011001100",
  32385=>"110100001",
  32386=>"111010101",
  32387=>"000001110",
  32388=>"110111100",
  32389=>"011000100",
  32390=>"011100010",
  32391=>"001010000",
  32392=>"001010111",
  32393=>"011110011",
  32394=>"111100101",
  32395=>"000001110",
  32396=>"000111001",
  32397=>"001101001",
  32398=>"101110101",
  32399=>"100111000",
  32400=>"100100100",
  32401=>"011001110",
  32402=>"010011110",
  32403=>"001101000",
  32404=>"011010011",
  32405=>"010100101",
  32406=>"010111001",
  32407=>"001010110",
  32408=>"110011101",
  32409=>"000011000",
  32410=>"101110101",
  32411=>"011011001",
  32412=>"011111110",
  32413=>"110011011",
  32414=>"001000000",
  32415=>"101011000",
  32416=>"000000101",
  32417=>"000010100",
  32418=>"000000101",
  32419=>"100001011",
  32420=>"100011111",
  32421=>"001010100",
  32422=>"001010100",
  32423=>"000000010",
  32424=>"010101111",
  32425=>"011100111",
  32426=>"100011000",
  32427=>"101011110",
  32428=>"100001011",
  32429=>"011100000",
  32430=>"011111011",
  32431=>"101110111",
  32432=>"110110010",
  32433=>"101101010",
  32434=>"000111010",
  32435=>"110010100",
  32436=>"110100101",
  32437=>"001101011",
  32438=>"100010111",
  32439=>"101001000",
  32440=>"010101100",
  32441=>"001100011",
  32442=>"001110100",
  32443=>"010000000",
  32444=>"011011001",
  32445=>"010000000",
  32446=>"011101111",
  32447=>"000110111",
  32448=>"101111011",
  32449=>"101100000",
  32450=>"010000000",
  32451=>"010000101",
  32452=>"001111010",
  32453=>"100000010",
  32454=>"010001000",
  32455=>"000001100",
  32456=>"110110110",
  32457=>"100100010",
  32458=>"010111011",
  32459=>"110001010",
  32460=>"000101000",
  32461=>"010000110",
  32462=>"011010011",
  32463=>"010101000",
  32464=>"100000010",
  32465=>"010101000",
  32466=>"111000011",
  32467=>"011010101",
  32468=>"011010010",
  32469=>"011111011",
  32470=>"100000010",
  32471=>"010110000",
  32472=>"111011000",
  32473=>"101011100",
  32474=>"000000111",
  32475=>"000000100",
  32476=>"000000000",
  32477=>"000001100",
  32478=>"101101001",
  32479=>"000011101",
  32480=>"111010010",
  32481=>"010001010",
  32482=>"110111100",
  32483=>"001011011",
  32484=>"000010101",
  32485=>"100000111",
  32486=>"111001100",
  32487=>"101001010",
  32488=>"000011101",
  32489=>"101010010",
  32490=>"111100101",
  32491=>"010000011",
  32492=>"000110000",
  32493=>"100001110",
  32494=>"010010001",
  32495=>"100101000",
  32496=>"111101111",
  32497=>"011010100",
  32498=>"010100000",
  32499=>"001110001",
  32500=>"100111101",
  32501=>"111010011",
  32502=>"001000011",
  32503=>"101010100",
  32504=>"100001101",
  32505=>"011111100",
  32506=>"000010001",
  32507=>"101101001",
  32508=>"000101001",
  32509=>"101100100",
  32510=>"001011100",
  32511=>"111011100",
  32512=>"011101101",
  32513=>"101001101",
  32514=>"110100010",
  32515=>"111001100",
  32516=>"000001010",
  32517=>"000111001",
  32518=>"111111111",
  32519=>"101100011",
  32520=>"000001101",
  32521=>"000001000",
  32522=>"111101010",
  32523=>"101101010",
  32524=>"111010101",
  32525=>"011010100",
  32526=>"111101110",
  32527=>"110111101",
  32528=>"111000111",
  32529=>"010011111",
  32530=>"101111010",
  32531=>"111010111",
  32532=>"010000001",
  32533=>"110101101",
  32534=>"101000111",
  32535=>"111011111",
  32536=>"111110001",
  32537=>"101010010",
  32538=>"111000011",
  32539=>"110110000",
  32540=>"010110000",
  32541=>"100011100",
  32542=>"010010101",
  32543=>"000101110",
  32544=>"011110110",
  32545=>"100111010",
  32546=>"010010011",
  32547=>"001111001",
  32548=>"110101101",
  32549=>"100001010",
  32550=>"110101010",
  32551=>"100000110",
  32552=>"111011011",
  32553=>"000101110",
  32554=>"000111101",
  32555=>"100010111",
  32556=>"100001011",
  32557=>"000000010",
  32558=>"111110111",
  32559=>"111011110",
  32560=>"001110011",
  32561=>"101000011",
  32562=>"111001110",
  32563=>"110101010",
  32564=>"100000110",
  32565=>"010000000",
  32566=>"101010100",
  32567=>"110111111",
  32568=>"011111001",
  32569=>"001101000",
  32570=>"000110101",
  32571=>"101000111",
  32572=>"111000111",
  32573=>"100100110",
  32574=>"111101011",
  32575=>"001011001",
  32576=>"001100101",
  32577=>"110000100",
  32578=>"101100000",
  32579=>"110001100",
  32580=>"100010111",
  32581=>"001000011",
  32582=>"100100010",
  32583=>"110110011",
  32584=>"011111101",
  32585=>"101000101",
  32586=>"101101000",
  32587=>"000011111",
  32588=>"011000110",
  32589=>"000101111",
  32590=>"100101000",
  32591=>"110011001",
  32592=>"001100101",
  32593=>"110100100",
  32594=>"001100010",
  32595=>"111111001",
  32596=>"101110101",
  32597=>"001100000",
  32598=>"101100011",
  32599=>"110010110",
  32600=>"001010101",
  32601=>"001011010",
  32602=>"001010000",
  32603=>"101101100",
  32604=>"100100010",
  32605=>"000010001",
  32606=>"110110001",
  32607=>"000101101",
  32608=>"011010000",
  32609=>"100011001",
  32610=>"010001101",
  32611=>"001000110",
  32612=>"001111001",
  32613=>"001001111",
  32614=>"110111011",
  32615=>"000100010",
  32616=>"000101110",
  32617=>"100000111",
  32618=>"111001001",
  32619=>"010000110",
  32620=>"111000100",
  32621=>"101110111",
  32622=>"100110000",
  32623=>"101111001",
  32624=>"010111000",
  32625=>"110111001",
  32626=>"001001111",
  32627=>"001111000",
  32628=>"011100100",
  32629=>"100011001",
  32630=>"001101101",
  32631=>"111010000",
  32632=>"000001011",
  32633=>"010010011",
  32634=>"011100000",
  32635=>"010111001",
  32636=>"010010000",
  32637=>"001000111",
  32638=>"101100000",
  32639=>"011100100",
  32640=>"010010001",
  32641=>"101111010",
  32642=>"001101001",
  32643=>"111101111",
  32644=>"000000100",
  32645=>"011111110",
  32646=>"000111101",
  32647=>"001001011",
  32648=>"110100110",
  32649=>"101111111",
  32650=>"000010111",
  32651=>"001000111",
  32652=>"101000101",
  32653=>"100000101",
  32654=>"101110000",
  32655=>"010111101",
  32656=>"111110101",
  32657=>"110100100",
  32658=>"111101100",
  32659=>"111111100",
  32660=>"100011110",
  32661=>"101111111",
  32662=>"111001010",
  32663=>"100101111",
  32664=>"100000100",
  32665=>"000110111",
  32666=>"011001100",
  32667=>"011110110",
  32668=>"001011111",
  32669=>"111110011",
  32670=>"001011000",
  32671=>"010111101",
  32672=>"010111010",
  32673=>"001010110",
  32674=>"100011001",
  32675=>"111101111",
  32676=>"000001010",
  32677=>"100100101",
  32678=>"100000010",
  32679=>"011101010",
  32680=>"101011011",
  32681=>"000000111",
  32682=>"110011100",
  32683=>"010000100",
  32684=>"101110100",
  32685=>"011110001",
  32686=>"100001010",
  32687=>"111110110",
  32688=>"100100111",
  32689=>"111110011",
  32690=>"000110000",
  32691=>"011010001",
  32692=>"010010010",
  32693=>"011100011",
  32694=>"010110001",
  32695=>"010000111",
  32696=>"010000000",
  32697=>"000011001",
  32698=>"010001011",
  32699=>"010010111",
  32700=>"001110110",
  32701=>"101110101",
  32702=>"101010111",
  32703=>"011111001",
  32704=>"100100000",
  32705=>"110001011",
  32706=>"011110101",
  32707=>"111101011",
  32708=>"000110001",
  32709=>"011100000",
  32710=>"001010111",
  32711=>"110101100",
  32712=>"111000101",
  32713=>"000010101",
  32714=>"000010101",
  32715=>"011100101",
  32716=>"000111101",
  32717=>"001001100",
  32718=>"101000101",
  32719=>"100101110",
  32720=>"010100001",
  32721=>"010100001",
  32722=>"000000011",
  32723=>"001001101",
  32724=>"001011100",
  32725=>"010001001",
  32726=>"110011000",
  32727=>"100111000",
  32728=>"001001111",
  32729=>"110011111",
  32730=>"110110000",
  32731=>"110001011",
  32732=>"100100010",
  32733=>"101101100",
  32734=>"001001101",
  32735=>"000001101",
  32736=>"001101110",
  32737=>"010011001",
  32738=>"100101010",
  32739=>"011011001",
  32740=>"111111001",
  32741=>"101100111",
  32742=>"000100000",
  32743=>"010000111",
  32744=>"100011011",
  32745=>"001111110",
  32746=>"001000101",
  32747=>"001111000",
  32748=>"110010111",
  32749=>"000110001",
  32750=>"101000001",
  32751=>"000000000",
  32752=>"101011010",
  32753=>"101011001",
  32754=>"001101010",
  32755=>"111100110",
  32756=>"101011101",
  32757=>"000000101",
  32758=>"100011010",
  32759=>"000000001",
  32760=>"011100100",
  32761=>"001000000",
  32762=>"001100100",
  32763=>"101111101",
  32764=>"001011011",
  32765=>"000011000",
  32766=>"001101000",
  32767=>"110111010",
  32768=>"110101000",
  32769=>"111011010",
  32770=>"110010110",
  32771=>"011000100",
  32772=>"000001011",
  32773=>"010001111",
  32774=>"101000100",
  32775=>"001100110",
  32776=>"101001010",
  32777=>"001101001",
  32778=>"000000101",
  32779=>"101011011",
  32780=>"001101000",
  32781=>"000001101",
  32782=>"010111010",
  32783=>"010100000",
  32784=>"001010110",
  32785=>"010111011",
  32786=>"100000100",
  32787=>"010111100",
  32788=>"100100000",
  32789=>"010110101",
  32790=>"110001101",
  32791=>"000100001",
  32792=>"100111100",
  32793=>"000001111",
  32794=>"001010101",
  32795=>"111100100",
  32796=>"001111010",
  32797=>"000111000",
  32798=>"111011010",
  32799=>"001011100",
  32800=>"101110011",
  32801=>"100000110",
  32802=>"001100011",
  32803=>"000101101",
  32804=>"101000110",
  32805=>"110110011",
  32806=>"100001100",
  32807=>"110001010",
  32808=>"011101001",
  32809=>"000000100",
  32810=>"101010011",
  32811=>"010101000",
  32812=>"000111101",
  32813=>"110010011",
  32814=>"101101001",
  32815=>"110010001",
  32816=>"110111101",
  32817=>"111101110",
  32818=>"010001000",
  32819=>"111111101",
  32820=>"111010110",
  32821=>"000011000",
  32822=>"100001010",
  32823=>"101010010",
  32824=>"100000000",
  32825=>"010011001",
  32826=>"000101010",
  32827=>"000100101",
  32828=>"000011101",
  32829=>"001011001",
  32830=>"110001000",
  32831=>"100000001",
  32832=>"011100001",
  32833=>"001000000",
  32834=>"011100001",
  32835=>"011001101",
  32836=>"101110000",
  32837=>"000100111",
  32838=>"101111110",
  32839=>"000001101",
  32840=>"001110110",
  32841=>"110010001",
  32842=>"000001101",
  32843=>"000101111",
  32844=>"110010001",
  32845=>"110010100",
  32846=>"111000000",
  32847=>"011001100",
  32848=>"110100101",
  32849=>"100001011",
  32850=>"001101011",
  32851=>"110110000",
  32852=>"001010000",
  32853=>"000011001",
  32854=>"101010000",
  32855=>"001111101",
  32856=>"101001101",
  32857=>"001000110",
  32858=>"011000110",
  32859=>"000100001",
  32860=>"000001111",
  32861=>"001010000",
  32862=>"000101101",
  32863=>"111001110",
  32864=>"000101010",
  32865=>"011101001",
  32866=>"100111000",
  32867=>"111000011",
  32868=>"111001001",
  32869=>"001110101",
  32870=>"111111100",
  32871=>"101101110",
  32872=>"010010000",
  32873=>"101011110",
  32874=>"010101001",
  32875=>"001010010",
  32876=>"101100111",
  32877=>"001100111",
  32878=>"101101010",
  32879=>"100011111",
  32880=>"111110100",
  32881=>"101111111",
  32882=>"010110010",
  32883=>"011010110",
  32884=>"100010100",
  32885=>"110001001",
  32886=>"100110111",
  32887=>"110110000",
  32888=>"111011001",
  32889=>"011101011",
  32890=>"010000000",
  32891=>"100000100",
  32892=>"010001110",
  32893=>"101010111",
  32894=>"000101100",
  32895=>"001011111",
  32896=>"111101110",
  32897=>"011010000",
  32898=>"001011001",
  32899=>"010001100",
  32900=>"100001101",
  32901=>"001001011",
  32902=>"001111111",
  32903=>"101101000",
  32904=>"000000010",
  32905=>"000001110",
  32906=>"111001101",
  32907=>"101001010",
  32908=>"010100110",
  32909=>"010001001",
  32910=>"101000101",
  32911=>"110010010",
  32912=>"100011000",
  32913=>"010101101",
  32914=>"000101101",
  32915=>"110011011",
  32916=>"101000001",
  32917=>"000000110",
  32918=>"011001011",
  32919=>"110110111",
  32920=>"100010001",
  32921=>"110010001",
  32922=>"010100100",
  32923=>"110011001",
  32924=>"011111000",
  32925=>"110010100",
  32926=>"110001000",
  32927=>"111010110",
  32928=>"000001101",
  32929=>"101010000",
  32930=>"001111111",
  32931=>"010001011",
  32932=>"010000110",
  32933=>"100001000",
  32934=>"010000000",
  32935=>"011010101",
  32936=>"001001100",
  32937=>"111101001",
  32938=>"001100000",
  32939=>"000100101",
  32940=>"100011111",
  32941=>"100111000",
  32942=>"110100000",
  32943=>"011000010",
  32944=>"011100001",
  32945=>"010001001",
  32946=>"111011010",
  32947=>"000101100",
  32948=>"100101101",
  32949=>"010011010",
  32950=>"100010001",
  32951=>"100111000",
  32952=>"100110111",
  32953=>"000100000",
  32954=>"111011111",
  32955=>"110111010",
  32956=>"001011110",
  32957=>"011111011",
  32958=>"000001111",
  32959=>"011011110",
  32960=>"001011000",
  32961=>"010101001",
  32962=>"001001000",
  32963=>"101101101",
  32964=>"110010010",
  32965=>"001111000",
  32966=>"100010111",
  32967=>"101000100",
  32968=>"011111111",
  32969=>"100100110",
  32970=>"001100110",
  32971=>"011011101",
  32972=>"111111100",
  32973=>"001100100",
  32974=>"101000000",
  32975=>"101001111",
  32976=>"110110001",
  32977=>"011101110",
  32978=>"100100011",
  32979=>"111110000",
  32980=>"111101100",
  32981=>"111100001",
  32982=>"101011110",
  32983=>"010100001",
  32984=>"101111100",
  32985=>"011001001",
  32986=>"100100001",
  32987=>"001001001",
  32988=>"100101111",
  32989=>"110101110",
  32990=>"101101111",
  32991=>"100000010",
  32992=>"001111011",
  32993=>"000101010",
  32994=>"000110110",
  32995=>"101000001",
  32996=>"111101001",
  32997=>"000001010",
  32998=>"110011111",
  32999=>"101100111",
  33000=>"011011110",
  33001=>"110111010",
  33002=>"000001000",
  33003=>"111001100",
  33004=>"111100000",
  33005=>"101000111",
  33006=>"000011000",
  33007=>"101010111",
  33008=>"010011010",
  33009=>"100100110",
  33010=>"101011001",
  33011=>"110100011",
  33012=>"110011000",
  33013=>"101111001",
  33014=>"001111111",
  33015=>"111101100",
  33016=>"010001000",
  33017=>"010011011",
  33018=>"110111000",
  33019=>"101101011",
  33020=>"100111011",
  33021=>"010110111",
  33022=>"111011010",
  33023=>"010001100",
  33024=>"111111011",
  33025=>"010110111",
  33026=>"110000111",
  33027=>"010001011",
  33028=>"010111111",
  33029=>"010010010",
  33030=>"010011011",
  33031=>"001000000",
  33032=>"100101001",
  33033=>"010000101",
  33034=>"111001100",
  33035=>"000000010",
  33036=>"010110000",
  33037=>"011000100",
  33038=>"100001011",
  33039=>"000110010",
  33040=>"100010010",
  33041=>"110000000",
  33042=>"110101000",
  33043=>"110100011",
  33044=>"001010011",
  33045=>"101000011",
  33046=>"001110101",
  33047=>"000100100",
  33048=>"010111111",
  33049=>"111001101",
  33050=>"000000101",
  33051=>"000101001",
  33052=>"100001000",
  33053=>"000111000",
  33054=>"111101111",
  33055=>"011000010",
  33056=>"000000100",
  33057=>"100011111",
  33058=>"011001011",
  33059=>"011010000",
  33060=>"110111011",
  33061=>"011100101",
  33062=>"000010000",
  33063=>"000010111",
  33064=>"110010010",
  33065=>"110011111",
  33066=>"111101001",
  33067=>"001110010",
  33068=>"010011100",
  33069=>"010110010",
  33070=>"001001101",
  33071=>"110011001",
  33072=>"011001111",
  33073=>"101110111",
  33074=>"000000101",
  33075=>"010011100",
  33076=>"011000101",
  33077=>"010101001",
  33078=>"000010011",
  33079=>"111001001",
  33080=>"000001001",
  33081=>"100100001",
  33082=>"010000000",
  33083=>"111001010",
  33084=>"010010011",
  33085=>"110110010",
  33086=>"110110100",
  33087=>"010100101",
  33088=>"010000001",
  33089=>"011001110",
  33090=>"000011111",
  33091=>"100111011",
  33092=>"000111111",
  33093=>"011011001",
  33094=>"010011001",
  33095=>"101001000",
  33096=>"110010111",
  33097=>"110000001",
  33098=>"001110010",
  33099=>"100011001",
  33100=>"000000110",
  33101=>"100100000",
  33102=>"000100000",
  33103=>"001110110",
  33104=>"100100101",
  33105=>"001010011",
  33106=>"110110011",
  33107=>"000111011",
  33108=>"000011101",
  33109=>"011101111",
  33110=>"101110100",
  33111=>"101110010",
  33112=>"010110110",
  33113=>"000000010",
  33114=>"110101101",
  33115=>"001001000",
  33116=>"010110100",
  33117=>"110101000",
  33118=>"010101110",
  33119=>"010100100",
  33120=>"000110111",
  33121=>"111101001",
  33122=>"010000101",
  33123=>"000000100",
  33124=>"011111111",
  33125=>"111001101",
  33126=>"001111100",
  33127=>"010000101",
  33128=>"010000000",
  33129=>"001111111",
  33130=>"100010110",
  33131=>"100101000",
  33132=>"011110011",
  33133=>"110100111",
  33134=>"110000000",
  33135=>"001011001",
  33136=>"010011100",
  33137=>"101001100",
  33138=>"111010001",
  33139=>"110011110",
  33140=>"101011100",
  33141=>"110011001",
  33142=>"000000100",
  33143=>"101111111",
  33144=>"010111110",
  33145=>"101010100",
  33146=>"001011101",
  33147=>"000010101",
  33148=>"001100110",
  33149=>"101111010",
  33150=>"111001101",
  33151=>"011000010",
  33152=>"001001110",
  33153=>"000011101",
  33154=>"111001101",
  33155=>"101100110",
  33156=>"110111100",
  33157=>"000010000",
  33158=>"110111110",
  33159=>"100001011",
  33160=>"011000110",
  33161=>"010110000",
  33162=>"010011011",
  33163=>"001100101",
  33164=>"001000111",
  33165=>"010100101",
  33166=>"001100000",
  33167=>"001001111",
  33168=>"010010010",
  33169=>"001001001",
  33170=>"000100000",
  33171=>"110001101",
  33172=>"110000111",
  33173=>"000010010",
  33174=>"111011011",
  33175=>"101000000",
  33176=>"100011000",
  33177=>"001001100",
  33178=>"000101001",
  33179=>"000111010",
  33180=>"110101101",
  33181=>"010110101",
  33182=>"010000001",
  33183=>"111110110",
  33184=>"101001010",
  33185=>"101100110",
  33186=>"000011111",
  33187=>"010100011",
  33188=>"101100001",
  33189=>"011111011",
  33190=>"010111100",
  33191=>"011111101",
  33192=>"110001100",
  33193=>"101110010",
  33194=>"001011000",
  33195=>"100011100",
  33196=>"010111110",
  33197=>"011010010",
  33198=>"011101100",
  33199=>"100010001",
  33200=>"010001001",
  33201=>"000000100",
  33202=>"110111000",
  33203=>"011011001",
  33204=>"001110001",
  33205=>"001010000",
  33206=>"101111011",
  33207=>"101011000",
  33208=>"111001010",
  33209=>"101000000",
  33210=>"000000111",
  33211=>"100010100",
  33212=>"101000101",
  33213=>"101100101",
  33214=>"001010110",
  33215=>"100101100",
  33216=>"011111110",
  33217=>"110110100",
  33218=>"111011111",
  33219=>"000111101",
  33220=>"100101001",
  33221=>"100101000",
  33222=>"011010000",
  33223=>"000101001",
  33224=>"011001011",
  33225=>"101001000",
  33226=>"000001101",
  33227=>"101110110",
  33228=>"011011000",
  33229=>"100001111",
  33230=>"000001100",
  33231=>"010000000",
  33232=>"010000101",
  33233=>"001011000",
  33234=>"100001011",
  33235=>"100101110",
  33236=>"001001100",
  33237=>"111111110",
  33238=>"100000110",
  33239=>"000110010",
  33240=>"001010101",
  33241=>"101010011",
  33242=>"110001010",
  33243=>"000001000",
  33244=>"101111111",
  33245=>"001010110",
  33246=>"011111110",
  33247=>"011101010",
  33248=>"100000110",
  33249=>"110101111",
  33250=>"110101010",
  33251=>"100000101",
  33252=>"011000010",
  33253=>"010001010",
  33254=>"011000010",
  33255=>"101100011",
  33256=>"100100000",
  33257=>"111100110",
  33258=>"001100011",
  33259=>"101010101",
  33260=>"110100000",
  33261=>"101010110",
  33262=>"000010011",
  33263=>"100011000",
  33264=>"011010011",
  33265=>"110101110",
  33266=>"010100100",
  33267=>"110000111",
  33268=>"101111011",
  33269=>"100000001",
  33270=>"000100100",
  33271=>"101101111",
  33272=>"001000101",
  33273=>"000010110",
  33274=>"111111101",
  33275=>"101101001",
  33276=>"000110100",
  33277=>"011100000",
  33278=>"001101110",
  33279=>"011010010",
  33280=>"100110101",
  33281=>"100011001",
  33282=>"010001001",
  33283=>"110101010",
  33284=>"000101010",
  33285=>"101000011",
  33286=>"100001001",
  33287=>"001101100",
  33288=>"100010101",
  33289=>"011100100",
  33290=>"100000011",
  33291=>"001001101",
  33292=>"111100011",
  33293=>"010000111",
  33294=>"100001001",
  33295=>"011011001",
  33296=>"101011000",
  33297=>"110010000",
  33298=>"110110101",
  33299=>"000011010",
  33300=>"100001001",
  33301=>"001100000",
  33302=>"011001010",
  33303=>"010011111",
  33304=>"100000101",
  33305=>"001001011",
  33306=>"001001000",
  33307=>"000010010",
  33308=>"110101110",
  33309=>"011000100",
  33310=>"001110111",
  33311=>"001001111",
  33312=>"010011001",
  33313=>"000100001",
  33314=>"101000110",
  33315=>"100011000",
  33316=>"101110001",
  33317=>"011001010",
  33318=>"010001001",
  33319=>"000100001",
  33320=>"100010110",
  33321=>"111010000",
  33322=>"011110011",
  33323=>"011011110",
  33324=>"110000010",
  33325=>"000100101",
  33326=>"100000001",
  33327=>"000010111",
  33328=>"101100011",
  33329=>"001000010",
  33330=>"111010101",
  33331=>"011111000",
  33332=>"111000100",
  33333=>"011001001",
  33334=>"000000001",
  33335=>"010000000",
  33336=>"011100111",
  33337=>"000010001",
  33338=>"100101001",
  33339=>"000110000",
  33340=>"011001001",
  33341=>"010001010",
  33342=>"011001010",
  33343=>"000010100",
  33344=>"110000100",
  33345=>"110001001",
  33346=>"101001100",
  33347=>"011011111",
  33348=>"000000000",
  33349=>"000011011",
  33350=>"100011001",
  33351=>"101100011",
  33352=>"001110000",
  33353=>"111001110",
  33354=>"011011100",
  33355=>"001110011",
  33356=>"010001010",
  33357=>"101010100",
  33358=>"111100110",
  33359=>"101100111",
  33360=>"110101000",
  33361=>"100100101",
  33362=>"111110001",
  33363=>"000101010",
  33364=>"101010110",
  33365=>"001101100",
  33366=>"110011011",
  33367=>"011111001",
  33368=>"111001100",
  33369=>"010000100",
  33370=>"011001011",
  33371=>"100010101",
  33372=>"101001010",
  33373=>"101110000",
  33374=>"000100000",
  33375=>"000000001",
  33376=>"110011010",
  33377=>"101001001",
  33378=>"000001100",
  33379=>"111001100",
  33380=>"001011100",
  33381=>"111110000",
  33382=>"010010101",
  33383=>"000100010",
  33384=>"000000000",
  33385=>"000001111",
  33386=>"000110011",
  33387=>"010001100",
  33388=>"000011011",
  33389=>"010001011",
  33390=>"010000000",
  33391=>"001000101",
  33392=>"011011011",
  33393=>"001110011",
  33394=>"100000111",
  33395=>"001110110",
  33396=>"100111000",
  33397=>"110000000",
  33398=>"110011000",
  33399=>"111101000",
  33400=>"010100111",
  33401=>"100001010",
  33402=>"011000100",
  33403=>"111101010",
  33404=>"001000001",
  33405=>"010010001",
  33406=>"000011001",
  33407=>"110101101",
  33408=>"000000110",
  33409=>"011101110",
  33410=>"111100100",
  33411=>"111110111",
  33412=>"001001100",
  33413=>"000110000",
  33414=>"101010110",
  33415=>"111111110",
  33416=>"110100000",
  33417=>"010101010",
  33418=>"100100011",
  33419=>"011000111",
  33420=>"111001111",
  33421=>"001011000",
  33422=>"110011001",
  33423=>"101000010",
  33424=>"100110011",
  33425=>"010001011",
  33426=>"111110001",
  33427=>"000110110",
  33428=>"001001111",
  33429=>"001110011",
  33430=>"011100110",
  33431=>"000000001",
  33432=>"000100000",
  33433=>"110111111",
  33434=>"111100110",
  33435=>"111000111",
  33436=>"101001011",
  33437=>"000000010",
  33438=>"001011001",
  33439=>"101010000",
  33440=>"111010100",
  33441=>"100101110",
  33442=>"101010001",
  33443=>"010001011",
  33444=>"001010011",
  33445=>"100001001",
  33446=>"010101100",
  33447=>"101000110",
  33448=>"011101001",
  33449=>"000100000",
  33450=>"100110111",
  33451=>"111000010",
  33452=>"100001100",
  33453=>"101111010",
  33454=>"110100100",
  33455=>"110000110",
  33456=>"101001101",
  33457=>"001100001",
  33458=>"110110101",
  33459=>"000011110",
  33460=>"100011110",
  33461=>"010100000",
  33462=>"000000010",
  33463=>"111100100",
  33464=>"101101000",
  33465=>"111111111",
  33466=>"100110100",
  33467=>"011100000",
  33468=>"011110001",
  33469=>"101111010",
  33470=>"001001001",
  33471=>"000101001",
  33472=>"100000100",
  33473=>"111001111",
  33474=>"000001000",
  33475=>"011101110",
  33476=>"100100101",
  33477=>"010000101",
  33478=>"110111011",
  33479=>"001000100",
  33480=>"010000100",
  33481=>"001010010",
  33482=>"010010001",
  33483=>"111001000",
  33484=>"001110110",
  33485=>"001101101",
  33486=>"011101101",
  33487=>"000111001",
  33488=>"101011000",
  33489=>"110010011",
  33490=>"100001100",
  33491=>"010011001",
  33492=>"001011101",
  33493=>"100111010",
  33494=>"011101010",
  33495=>"101101010",
  33496=>"001001011",
  33497=>"010111011",
  33498=>"101001111",
  33499=>"011110000",
  33500=>"101111001",
  33501=>"100101000",
  33502=>"011010110",
  33503=>"100000001",
  33504=>"010101011",
  33505=>"001001001",
  33506=>"100111010",
  33507=>"000001001",
  33508=>"111011001",
  33509=>"100000010",
  33510=>"100000101",
  33511=>"011011100",
  33512=>"101100100",
  33513=>"111110111",
  33514=>"110111011",
  33515=>"011011001",
  33516=>"000011001",
  33517=>"010111100",
  33518=>"110111000",
  33519=>"000101010",
  33520=>"001100101",
  33521=>"001001011",
  33522=>"010111010",
  33523=>"000000101",
  33524=>"101100010",
  33525=>"010111011",
  33526=>"111111100",
  33527=>"111111011",
  33528=>"111010011",
  33529=>"010000110",
  33530=>"110001111",
  33531=>"001011100",
  33532=>"001110011",
  33533=>"110111100",
  33534=>"110000110",
  33535=>"000101101",
  33536=>"110000110",
  33537=>"000100100",
  33538=>"001110011",
  33539=>"101010100",
  33540=>"100101000",
  33541=>"001101101",
  33542=>"101000011",
  33543=>"000100000",
  33544=>"100111010",
  33545=>"000100111",
  33546=>"111100001",
  33547=>"101111011",
  33548=>"101100000",
  33549=>"100111111",
  33550=>"010100110",
  33551=>"111010011",
  33552=>"000110010",
  33553=>"101100101",
  33554=>"111011010",
  33555=>"001010010",
  33556=>"110111000",
  33557=>"100000001",
  33558=>"001011001",
  33559=>"100010011",
  33560=>"000010100",
  33561=>"101100110",
  33562=>"010001111",
  33563=>"110010000",
  33564=>"100000110",
  33565=>"011101100",
  33566=>"011001011",
  33567=>"101011011",
  33568=>"001110000",
  33569=>"001011110",
  33570=>"000000111",
  33571=>"101010000",
  33572=>"011001001",
  33573=>"100010010",
  33574=>"110000111",
  33575=>"110110100",
  33576=>"011111111",
  33577=>"100011000",
  33578=>"001000110",
  33579=>"001110011",
  33580=>"101011111",
  33581=>"000110100",
  33582=>"110001010",
  33583=>"110011001",
  33584=>"011001000",
  33585=>"111111011",
  33586=>"000000011",
  33587=>"000111110",
  33588=>"001100001",
  33589=>"100010101",
  33590=>"011001010",
  33591=>"000001001",
  33592=>"001111001",
  33593=>"100000000",
  33594=>"001100011",
  33595=>"111100110",
  33596=>"100001111",
  33597=>"001100101",
  33598=>"101100101",
  33599=>"100110000",
  33600=>"011100101",
  33601=>"110001000",
  33602=>"010100000",
  33603=>"110110111",
  33604=>"101100011",
  33605=>"010101100",
  33606=>"011011011",
  33607=>"100001001",
  33608=>"000010100",
  33609=>"001100001",
  33610=>"110101000",
  33611=>"100101010",
  33612=>"100000111",
  33613=>"001000010",
  33614=>"001111111",
  33615=>"000110001",
  33616=>"011100100",
  33617=>"110000110",
  33618=>"001111011",
  33619=>"111011010",
  33620=>"110110010",
  33621=>"001000100",
  33622=>"111100001",
  33623=>"111100101",
  33624=>"100001101",
  33625=>"010000100",
  33626=>"111101111",
  33627=>"100100001",
  33628=>"000101000",
  33629=>"010110100",
  33630=>"011010010",
  33631=>"010001001",
  33632=>"010010011",
  33633=>"111111010",
  33634=>"010100000",
  33635=>"011110110",
  33636=>"111101110",
  33637=>"000101000",
  33638=>"001100001",
  33639=>"101110111",
  33640=>"001110100",
  33641=>"100101000",
  33642=>"110011011",
  33643=>"010010001",
  33644=>"100111011",
  33645=>"100011111",
  33646=>"010101100",
  33647=>"011111100",
  33648=>"011001000",
  33649=>"101000011",
  33650=>"110010101",
  33651=>"000011010",
  33652=>"101011000",
  33653=>"101100100",
  33654=>"110101111",
  33655=>"111101101",
  33656=>"011010000",
  33657=>"110010101",
  33658=>"101010110",
  33659=>"111011100",
  33660=>"110010010",
  33661=>"111001001",
  33662=>"000100010",
  33663=>"111101000",
  33664=>"010111001",
  33665=>"101011000",
  33666=>"010011110",
  33667=>"010110000",
  33668=>"100000000",
  33669=>"010100101",
  33670=>"010000101",
  33671=>"000001001",
  33672=>"110111101",
  33673=>"101101010",
  33674=>"111110110",
  33675=>"001001101",
  33676=>"110000111",
  33677=>"111000111",
  33678=>"011101010",
  33679=>"000100101",
  33680=>"001100001",
  33681=>"001000110",
  33682=>"001000100",
  33683=>"001000111",
  33684=>"001000111",
  33685=>"100000001",
  33686=>"010100000",
  33687=>"100000011",
  33688=>"001101100",
  33689=>"010010110",
  33690=>"001111001",
  33691=>"000000101",
  33692=>"100101011",
  33693=>"000011110",
  33694=>"010001110",
  33695=>"001010011",
  33696=>"011011011",
  33697=>"111001111",
  33698=>"000111111",
  33699=>"000001100",
  33700=>"011010000",
  33701=>"111100010",
  33702=>"111000100",
  33703=>"011001110",
  33704=>"111010000",
  33705=>"000100111",
  33706=>"100010101",
  33707=>"111011110",
  33708=>"000111000",
  33709=>"000110010",
  33710=>"110100011",
  33711=>"101101001",
  33712=>"000110100",
  33713=>"001111101",
  33714=>"111101000",
  33715=>"010100010",
  33716=>"110101011",
  33717=>"111101111",
  33718=>"000101100",
  33719=>"000011101",
  33720=>"001100100",
  33721=>"000010000",
  33722=>"101101010",
  33723=>"100111001",
  33724=>"011100000",
  33725=>"100000100",
  33726=>"101001111",
  33727=>"001011001",
  33728=>"111000110",
  33729=>"111001111",
  33730=>"101001011",
  33731=>"111000111",
  33732=>"100010111",
  33733=>"110101111",
  33734=>"011110101",
  33735=>"011110011",
  33736=>"011011110",
  33737=>"000011110",
  33738=>"001100110",
  33739=>"110111011",
  33740=>"011111111",
  33741=>"110010110",
  33742=>"000100100",
  33743=>"111011100",
  33744=>"100111011",
  33745=>"101100011",
  33746=>"100110000",
  33747=>"000010010",
  33748=>"011011000",
  33749=>"001000110",
  33750=>"101101011",
  33751=>"100110111",
  33752=>"100001001",
  33753=>"011110011",
  33754=>"001111010",
  33755=>"100000111",
  33756=>"110000001",
  33757=>"011111010",
  33758=>"110001010",
  33759=>"011001000",
  33760=>"000011011",
  33761=>"101011101",
  33762=>"001011001",
  33763=>"010001111",
  33764=>"001011101",
  33765=>"011011001",
  33766=>"000100011",
  33767=>"000100100",
  33768=>"010101001",
  33769=>"011010001",
  33770=>"100101001",
  33771=>"111001000",
  33772=>"010111100",
  33773=>"101011110",
  33774=>"011011111",
  33775=>"101100100",
  33776=>"000111000",
  33777=>"000101011",
  33778=>"100110101",
  33779=>"101101101",
  33780=>"110010011",
  33781=>"001101111",
  33782=>"000101111",
  33783=>"011010010",
  33784=>"011111100",
  33785=>"101000010",
  33786=>"000110001",
  33787=>"010110110",
  33788=>"101111111",
  33789=>"101000000",
  33790=>"110011001",
  33791=>"110011000",
  33792=>"010010111",
  33793=>"111111011",
  33794=>"001111000",
  33795=>"010000101",
  33796=>"011010010",
  33797=>"010010110",
  33798=>"010010100",
  33799=>"110110111",
  33800=>"011001000",
  33801=>"100011111",
  33802=>"110110000",
  33803=>"001011111",
  33804=>"100110101",
  33805=>"001001010",
  33806=>"101100111",
  33807=>"101011101",
  33808=>"001110101",
  33809=>"111111111",
  33810=>"010101100",
  33811=>"001000000",
  33812=>"010000100",
  33813=>"111000110",
  33814=>"001110100",
  33815=>"000110001",
  33816=>"110100110",
  33817=>"001110110",
  33818=>"100000000",
  33819=>"110100100",
  33820=>"110101110",
  33821=>"100001000",
  33822=>"111000001",
  33823=>"011001001",
  33824=>"011010110",
  33825=>"001101010",
  33826=>"110101110",
  33827=>"011110100",
  33828=>"110011111",
  33829=>"101111101",
  33830=>"010111011",
  33831=>"100100000",
  33832=>"110000000",
  33833=>"111000010",
  33834=>"101110111",
  33835=>"111000100",
  33836=>"000110001",
  33837=>"011001011",
  33838=>"101101000",
  33839=>"010000010",
  33840=>"110101010",
  33841=>"010000110",
  33842=>"011001111",
  33843=>"111111101",
  33844=>"100011011",
  33845=>"001110001",
  33846=>"110101000",
  33847=>"101100111",
  33848=>"111111001",
  33849=>"110011001",
  33850=>"001111011",
  33851=>"010100000",
  33852=>"010000001",
  33853=>"000000010",
  33854=>"101100000",
  33855=>"001000011",
  33856=>"000001110",
  33857=>"010010100",
  33858=>"101101101",
  33859=>"000011001",
  33860=>"110110110",
  33861=>"001000001",
  33862=>"011101011",
  33863=>"111010111",
  33864=>"111110000",
  33865=>"111010101",
  33866=>"100000100",
  33867=>"000011101",
  33868=>"110101000",
  33869=>"100001111",
  33870=>"000010010",
  33871=>"001011110",
  33872=>"111001111",
  33873=>"000011110",
  33874=>"001010110",
  33875=>"110111011",
  33876=>"110111100",
  33877=>"110101100",
  33878=>"001001011",
  33879=>"000110000",
  33880=>"000010110",
  33881=>"111111001",
  33882=>"101010100",
  33883=>"011010000",
  33884=>"111001110",
  33885=>"101001011",
  33886=>"101100101",
  33887=>"000011010",
  33888=>"000100110",
  33889=>"101010011",
  33890=>"000010010",
  33891=>"101111101",
  33892=>"100010100",
  33893=>"000100110",
  33894=>"000010001",
  33895=>"001001011",
  33896=>"001101000",
  33897=>"101101011",
  33898=>"110001101",
  33899=>"000001010",
  33900=>"000000011",
  33901=>"110011100",
  33902=>"110011111",
  33903=>"110011111",
  33904=>"001001001",
  33905=>"011001110",
  33906=>"011111111",
  33907=>"000111110",
  33908=>"010100000",
  33909=>"110111110",
  33910=>"101100101",
  33911=>"000110100",
  33912=>"100000000",
  33913=>"101010101",
  33914=>"100000101",
  33915=>"000011100",
  33916=>"010001001",
  33917=>"001110001",
  33918=>"100000110",
  33919=>"000001110",
  33920=>"101111011",
  33921=>"100010101",
  33922=>"100110011",
  33923=>"000001100",
  33924=>"000010001",
  33925=>"110011000",
  33926=>"111111111",
  33927=>"011100100",
  33928=>"011100001",
  33929=>"110110101",
  33930=>"111100011",
  33931=>"111110010",
  33932=>"111100000",
  33933=>"010000110",
  33934=>"011111000",
  33935=>"110011101",
  33936=>"010011100",
  33937=>"111001010",
  33938=>"100000011",
  33939=>"111100100",
  33940=>"100110000",
  33941=>"000011010",
  33942=>"111110100",
  33943=>"001000001",
  33944=>"011000101",
  33945=>"011101001",
  33946=>"101000001",
  33947=>"111111100",
  33948=>"111101110",
  33949=>"000111010",
  33950=>"101000100",
  33951=>"110010100",
  33952=>"110110010",
  33953=>"100100111",
  33954=>"101101000",
  33955=>"001010111",
  33956=>"101101110",
  33957=>"100001001",
  33958=>"110010000",
  33959=>"001000100",
  33960=>"111111000",
  33961=>"000001100",
  33962=>"110101100",
  33963=>"100100011",
  33964=>"110111011",
  33965=>"100011010",
  33966=>"011010010",
  33967=>"011001101",
  33968=>"001001001",
  33969=>"001001011",
  33970=>"010000000",
  33971=>"100001011",
  33972=>"011100111",
  33973=>"110000000",
  33974=>"010100000",
  33975=>"110111100",
  33976=>"011100001",
  33977=>"100011000",
  33978=>"110011000",
  33979=>"010010110",
  33980=>"101010001",
  33981=>"111001000",
  33982=>"000001001",
  33983=>"100011010",
  33984=>"010110110",
  33985=>"000010110",
  33986=>"000010111",
  33987=>"010000011",
  33988=>"000011110",
  33989=>"101010101",
  33990=>"111101011",
  33991=>"000001111",
  33992=>"110111111",
  33993=>"101101110",
  33994=>"001001010",
  33995=>"011101001",
  33996=>"111110110",
  33997=>"000100111",
  33998=>"011010110",
  33999=>"000010000",
  34000=>"011100011",
  34001=>"000000111",
  34002=>"000011010",
  34003=>"011100001",
  34004=>"001111010",
  34005=>"011010000",
  34006=>"010111100",
  34007=>"010110111",
  34008=>"011110101",
  34009=>"010010000",
  34010=>"000100100",
  34011=>"011101110",
  34012=>"101101110",
  34013=>"001011100",
  34014=>"000110000",
  34015=>"110110111",
  34016=>"001100011",
  34017=>"010010001",
  34018=>"100110111",
  34019=>"000100101",
  34020=>"100100001",
  34021=>"110000101",
  34022=>"011001101",
  34023=>"111010101",
  34024=>"100110001",
  34025=>"011011111",
  34026=>"001111100",
  34027=>"100001100",
  34028=>"101000101",
  34029=>"001001001",
  34030=>"010000100",
  34031=>"010100000",
  34032=>"110000111",
  34033=>"111001010",
  34034=>"111010011",
  34035=>"110001010",
  34036=>"111110101",
  34037=>"110101001",
  34038=>"110110111",
  34039=>"101100100",
  34040=>"100011101",
  34041=>"110011100",
  34042=>"010110010",
  34043=>"101101010",
  34044=>"000110100",
  34045=>"000100111",
  34046=>"100000111",
  34047=>"111010100",
  34048=>"000000000",
  34049=>"110011001",
  34050=>"001111111",
  34051=>"010010101",
  34052=>"111001101",
  34053=>"001001111",
  34054=>"010010011",
  34055=>"101001011",
  34056=>"001110010",
  34057=>"011110001",
  34058=>"001000010",
  34059=>"000011100",
  34060=>"011100000",
  34061=>"010001101",
  34062=>"000011011",
  34063=>"101011110",
  34064=>"110110000",
  34065=>"110101001",
  34066=>"110110000",
  34067=>"001101011",
  34068=>"001001101",
  34069=>"100001110",
  34070=>"101001011",
  34071=>"111001110",
  34072=>"110110110",
  34073=>"110110000",
  34074=>"000110111",
  34075=>"110110110",
  34076=>"000101101",
  34077=>"111011111",
  34078=>"010100100",
  34079=>"001000101",
  34080=>"010100011",
  34081=>"001100001",
  34082=>"011010000",
  34083=>"100110011",
  34084=>"000001100",
  34085=>"110000011",
  34086=>"010000000",
  34087=>"010110010",
  34088=>"110000000",
  34089=>"010001110",
  34090=>"011100101",
  34091=>"001000100",
  34092=>"111000000",
  34093=>"000000101",
  34094=>"101101000",
  34095=>"010110010",
  34096=>"101000001",
  34097=>"001101000",
  34098=>"010000111",
  34099=>"111000110",
  34100=>"010000000",
  34101=>"110111001",
  34102=>"010000001",
  34103=>"010110011",
  34104=>"000111111",
  34105=>"101001110",
  34106=>"000001100",
  34107=>"101101001",
  34108=>"001100101",
  34109=>"111000000",
  34110=>"110011100",
  34111=>"100110000",
  34112=>"000010010",
  34113=>"111110001",
  34114=>"010010101",
  34115=>"000110000",
  34116=>"010110000",
  34117=>"110110001",
  34118=>"000001101",
  34119=>"000000000",
  34120=>"110101001",
  34121=>"000010101",
  34122=>"000101010",
  34123=>"000001010",
  34124=>"100111110",
  34125=>"111110111",
  34126=>"010100101",
  34127=>"101101110",
  34128=>"011101001",
  34129=>"110101110",
  34130=>"110010000",
  34131=>"100100000",
  34132=>"001010011",
  34133=>"111100100",
  34134=>"011000101",
  34135=>"111111001",
  34136=>"111101100",
  34137=>"111010010",
  34138=>"001101111",
  34139=>"011100001",
  34140=>"011011111",
  34141=>"100011000",
  34142=>"001001100",
  34143=>"000111101",
  34144=>"010011110",
  34145=>"011011110",
  34146=>"111100010",
  34147=>"011011000",
  34148=>"011010010",
  34149=>"011101100",
  34150=>"101001011",
  34151=>"101100100",
  34152=>"100111100",
  34153=>"010010011",
  34154=>"100100100",
  34155=>"011100110",
  34156=>"101101110",
  34157=>"010111110",
  34158=>"000011000",
  34159=>"111101110",
  34160=>"010011100",
  34161=>"100101110",
  34162=>"100000000",
  34163=>"110010000",
  34164=>"011111000",
  34165=>"000010100",
  34166=>"000101001",
  34167=>"011011110",
  34168=>"011001000",
  34169=>"101001011",
  34170=>"000101111",
  34171=>"100010100",
  34172=>"111010110",
  34173=>"110101101",
  34174=>"111011011",
  34175=>"111101100",
  34176=>"111001011",
  34177=>"100110001",
  34178=>"000100101",
  34179=>"011011010",
  34180=>"100101111",
  34181=>"101010010",
  34182=>"100001010",
  34183=>"100010000",
  34184=>"110101010",
  34185=>"001011011",
  34186=>"010110111",
  34187=>"001000011",
  34188=>"110111010",
  34189=>"000010111",
  34190=>"101000111",
  34191=>"001011111",
  34192=>"111011011",
  34193=>"001000111",
  34194=>"110100100",
  34195=>"110011110",
  34196=>"010101110",
  34197=>"100011011",
  34198=>"100111111",
  34199=>"100110101",
  34200=>"111010011",
  34201=>"101101111",
  34202=>"111000001",
  34203=>"100000001",
  34204=>"101101001",
  34205=>"011011110",
  34206=>"010110010",
  34207=>"001101011",
  34208=>"100100101",
  34209=>"000000100",
  34210=>"001100010",
  34211=>"000011010",
  34212=>"000000111",
  34213=>"101010010",
  34214=>"000101011",
  34215=>"111101000",
  34216=>"100101101",
  34217=>"100010001",
  34218=>"010001010",
  34219=>"001011110",
  34220=>"000100100",
  34221=>"101010000",
  34222=>"011000010",
  34223=>"101100011",
  34224=>"101101000",
  34225=>"011001011",
  34226=>"010011011",
  34227=>"000010110",
  34228=>"100001000",
  34229=>"111101011",
  34230=>"111001000",
  34231=>"101000010",
  34232=>"011011000",
  34233=>"101000111",
  34234=>"000010000",
  34235=>"001100110",
  34236=>"101100110",
  34237=>"001111011",
  34238=>"101110101",
  34239=>"101101111",
  34240=>"100100100",
  34241=>"100000000",
  34242=>"101011011",
  34243=>"101100111",
  34244=>"001100111",
  34245=>"001011101",
  34246=>"110101011",
  34247=>"110001000",
  34248=>"011000110",
  34249=>"100011001",
  34250=>"101011010",
  34251=>"000110100",
  34252=>"101111001",
  34253=>"101111101",
  34254=>"011001110",
  34255=>"000010100",
  34256=>"111001101",
  34257=>"111100010",
  34258=>"100100011",
  34259=>"110001110",
  34260=>"001110101",
  34261=>"100001000",
  34262=>"100100101",
  34263=>"110011110",
  34264=>"100111101",
  34265=>"011110000",
  34266=>"011011010",
  34267=>"000000010",
  34268=>"011110000",
  34269=>"010100101",
  34270=>"011100011",
  34271=>"110110010",
  34272=>"101111110",
  34273=>"001011101",
  34274=>"001111111",
  34275=>"111111100",
  34276=>"100100000",
  34277=>"100101011",
  34278=>"111101011",
  34279=>"100001011",
  34280=>"111111011",
  34281=>"101110000",
  34282=>"010100011",
  34283=>"110100111",
  34284=>"011011101",
  34285=>"010011010",
  34286=>"111001110",
  34287=>"111001000",
  34288=>"001101001",
  34289=>"011000111",
  34290=>"101100101",
  34291=>"011010010",
  34292=>"111111001",
  34293=>"111010110",
  34294=>"001100010",
  34295=>"111110110",
  34296=>"010000100",
  34297=>"001001110",
  34298=>"001001111",
  34299=>"010010110",
  34300=>"001011110",
  34301=>"100101111",
  34302=>"101000101",
  34303=>"111010101",
  34304=>"111000001",
  34305=>"001000111",
  34306=>"000101001",
  34307=>"111111010",
  34308=>"101110010",
  34309=>"111110010",
  34310=>"100010011",
  34311=>"111010001",
  34312=>"000111101",
  34313=>"100110110",
  34314=>"010100110",
  34315=>"110001101",
  34316=>"110000111",
  34317=>"110110011",
  34318=>"110000010",
  34319=>"011100010",
  34320=>"000000000",
  34321=>"110001100",
  34322=>"111001010",
  34323=>"100101011",
  34324=>"000111110",
  34325=>"111100000",
  34326=>"101011010",
  34327=>"101111100",
  34328=>"010000111",
  34329=>"000101001",
  34330=>"100111000",
  34331=>"010010110",
  34332=>"100110110",
  34333=>"010111000",
  34334=>"111110000",
  34335=>"001100111",
  34336=>"100110110",
  34337=>"110011111",
  34338=>"011001011",
  34339=>"001101001",
  34340=>"100100001",
  34341=>"001001101",
  34342=>"000000001",
  34343=>"010110110",
  34344=>"111101001",
  34345=>"100011010",
  34346=>"111110000",
  34347=>"001101001",
  34348=>"100100100",
  34349=>"011010010",
  34350=>"111101011",
  34351=>"001000100",
  34352=>"110000111",
  34353=>"010000100",
  34354=>"001111110",
  34355=>"001110100",
  34356=>"010111110",
  34357=>"110111001",
  34358=>"001001101",
  34359=>"000101001",
  34360=>"001110011",
  34361=>"000000011",
  34362=>"010111001",
  34363=>"110100110",
  34364=>"100010111",
  34365=>"100111011",
  34366=>"110011110",
  34367=>"000110001",
  34368=>"011111010",
  34369=>"011100010",
  34370=>"000011111",
  34371=>"111101011",
  34372=>"100011100",
  34373=>"100011110",
  34374=>"001100100",
  34375=>"101011000",
  34376=>"001110111",
  34377=>"011100100",
  34378=>"011101111",
  34379=>"010100010",
  34380=>"100111111",
  34381=>"000101100",
  34382=>"111101111",
  34383=>"100011001",
  34384=>"010111111",
  34385=>"000011000",
  34386=>"101001001",
  34387=>"111010010",
  34388=>"101101101",
  34389=>"101101101",
  34390=>"100001011",
  34391=>"110111011",
  34392=>"001100100",
  34393=>"101111101",
  34394=>"100110011",
  34395=>"111111010",
  34396=>"010100010",
  34397=>"000011000",
  34398=>"111101001",
  34399=>"111010111",
  34400=>"001000110",
  34401=>"100111110",
  34402=>"010011011",
  34403=>"100011000",
  34404=>"000001001",
  34405=>"000010111",
  34406=>"101111001",
  34407=>"101101000",
  34408=>"111000111",
  34409=>"001101011",
  34410=>"011001010",
  34411=>"000010000",
  34412=>"001000110",
  34413=>"100000111",
  34414=>"101101011",
  34415=>"010000001",
  34416=>"101111000",
  34417=>"010000101",
  34418=>"111101111",
  34419=>"010100000",
  34420=>"010000101",
  34421=>"001110001",
  34422=>"000000010",
  34423=>"100001010",
  34424=>"100101110",
  34425=>"011011011",
  34426=>"101001001",
  34427=>"000010101",
  34428=>"111110011",
  34429=>"001000110",
  34430=>"110001101",
  34431=>"000100000",
  34432=>"011011000",
  34433=>"010000010",
  34434=>"001111111",
  34435=>"001000001",
  34436=>"011111101",
  34437=>"010110010",
  34438=>"111111000",
  34439=>"111111101",
  34440=>"010101001",
  34441=>"000000000",
  34442=>"101010000",
  34443=>"110000001",
  34444=>"001010110",
  34445=>"001000000",
  34446=>"000100100",
  34447=>"011101000",
  34448=>"100100110",
  34449=>"110111011",
  34450=>"000101001",
  34451=>"010000011",
  34452=>"000001101",
  34453=>"000011010",
  34454=>"000001000",
  34455=>"101010100",
  34456=>"010011101",
  34457=>"001001111",
  34458=>"010001010",
  34459=>"011110001",
  34460=>"010110111",
  34461=>"000110111",
  34462=>"111100010",
  34463=>"001000001",
  34464=>"101110001",
  34465=>"001011011",
  34466=>"101111010",
  34467=>"110001010",
  34468=>"001001011",
  34469=>"010101100",
  34470=>"110101111",
  34471=>"010101000",
  34472=>"100010100",
  34473=>"001000010",
  34474=>"000110100",
  34475=>"010100001",
  34476=>"011001010",
  34477=>"010111111",
  34478=>"000111111",
  34479=>"110010001",
  34480=>"001111101",
  34481=>"101000010",
  34482=>"101101001",
  34483=>"010111100",
  34484=>"000011110",
  34485=>"001000100",
  34486=>"101010001",
  34487=>"100000110",
  34488=>"010010001",
  34489=>"001111001",
  34490=>"010010011",
  34491=>"101101111",
  34492=>"011111001",
  34493=>"011111010",
  34494=>"001000101",
  34495=>"100011001",
  34496=>"110111010",
  34497=>"010000001",
  34498=>"010110111",
  34499=>"110011101",
  34500=>"011010100",
  34501=>"010110010",
  34502=>"011001010",
  34503=>"100000101",
  34504=>"011101001",
  34505=>"100110111",
  34506=>"000100011",
  34507=>"011011001",
  34508=>"110100001",
  34509=>"011110101",
  34510=>"001001111",
  34511=>"110101100",
  34512=>"100001011",
  34513=>"010011010",
  34514=>"111000000",
  34515=>"011011111",
  34516=>"111000110",
  34517=>"001010101",
  34518=>"010101101",
  34519=>"000010111",
  34520=>"001001111",
  34521=>"010001000",
  34522=>"011111000",
  34523=>"011000101",
  34524=>"001010111",
  34525=>"011111011",
  34526=>"000010000",
  34527=>"110101011",
  34528=>"100010000",
  34529=>"010101011",
  34530=>"001111111",
  34531=>"111011101",
  34532=>"001110110",
  34533=>"111111001",
  34534=>"101001010",
  34535=>"010100100",
  34536=>"000110001",
  34537=>"101110101",
  34538=>"001100001",
  34539=>"110010111",
  34540=>"010000010",
  34541=>"000011100",
  34542=>"011011010",
  34543=>"000001011",
  34544=>"010001110",
  34545=>"101111110",
  34546=>"000100000",
  34547=>"111111001",
  34548=>"100011010",
  34549=>"100000000",
  34550=>"101110100",
  34551=>"101001001",
  34552=>"100001000",
  34553=>"100010000",
  34554=>"000101000",
  34555=>"100001110",
  34556=>"100101100",
  34557=>"011010010",
  34558=>"011010101",
  34559=>"000111000",
  34560=>"100001101",
  34561=>"110101000",
  34562=>"101011111",
  34563=>"110111011",
  34564=>"110111111",
  34565=>"000010010",
  34566=>"111111110",
  34567=>"011110101",
  34568=>"101111110",
  34569=>"000000111",
  34570=>"000010110",
  34571=>"111101111",
  34572=>"010110110",
  34573=>"110111011",
  34574=>"001001111",
  34575=>"111110100",
  34576=>"010111000",
  34577=>"101010010",
  34578=>"110010000",
  34579=>"110110110",
  34580=>"110001001",
  34581=>"011000010",
  34582=>"111000011",
  34583=>"011000101",
  34584=>"100101000",
  34585=>"010001010",
  34586=>"000001110",
  34587=>"011111001",
  34588=>"011011000",
  34589=>"001001010",
  34590=>"110110111",
  34591=>"010111011",
  34592=>"101000010",
  34593=>"001010110",
  34594=>"000010001",
  34595=>"011111110",
  34596=>"000001001",
  34597=>"000101110",
  34598=>"101000000",
  34599=>"000000111",
  34600=>"011111000",
  34601=>"010101110",
  34602=>"000000100",
  34603=>"110010010",
  34604=>"011110010",
  34605=>"000100000",
  34606=>"101111111",
  34607=>"100000100",
  34608=>"101011010",
  34609=>"101101001",
  34610=>"111111100",
  34611=>"110110000",
  34612=>"010101011",
  34613=>"100000001",
  34614=>"101011011",
  34615=>"111000011",
  34616=>"110011011",
  34617=>"000000001",
  34618=>"111100111",
  34619=>"111000111",
  34620=>"101111110",
  34621=>"010011100",
  34622=>"110010110",
  34623=>"010000110",
  34624=>"101111001",
  34625=>"010010101",
  34626=>"101000110",
  34627=>"010011010",
  34628=>"100110100",
  34629=>"101111000",
  34630=>"011111101",
  34631=>"000001011",
  34632=>"111111001",
  34633=>"110010100",
  34634=>"100000101",
  34635=>"111000000",
  34636=>"000001001",
  34637=>"100111000",
  34638=>"111000001",
  34639=>"111110111",
  34640=>"100010010",
  34641=>"100111001",
  34642=>"000010000",
  34643=>"100111000",
  34644=>"100010111",
  34645=>"100100101",
  34646=>"011111010",
  34647=>"111100100",
  34648=>"011010100",
  34649=>"111111001",
  34650=>"001011111",
  34651=>"000011010",
  34652=>"000000001",
  34653=>"100000010",
  34654=>"100110101",
  34655=>"100000000",
  34656=>"111111001",
  34657=>"111110011",
  34658=>"111001010",
  34659=>"000100000",
  34660=>"001010100",
  34661=>"110100111",
  34662=>"010000101",
  34663=>"011001101",
  34664=>"101000111",
  34665=>"100010110",
  34666=>"011111000",
  34667=>"110011111",
  34668=>"011111100",
  34669=>"110001001",
  34670=>"111011110",
  34671=>"010101010",
  34672=>"111100000",
  34673=>"011100111",
  34674=>"111011010",
  34675=>"101010010",
  34676=>"111010001",
  34677=>"000000000",
  34678=>"000001011",
  34679=>"010111111",
  34680=>"100110110",
  34681=>"001000000",
  34682=>"011111110",
  34683=>"000010011",
  34684=>"110011000",
  34685=>"011010000",
  34686=>"111001001",
  34687=>"110011111",
  34688=>"011010000",
  34689=>"011010110",
  34690=>"101010111",
  34691=>"100011111",
  34692=>"011100001",
  34693=>"100110101",
  34694=>"111101100",
  34695=>"100010000",
  34696=>"000010110",
  34697=>"100110000",
  34698=>"001001111",
  34699=>"111111100",
  34700=>"011110111",
  34701=>"111000110",
  34702=>"110100010",
  34703=>"111011000",
  34704=>"000000111",
  34705=>"000101111",
  34706=>"111011011",
  34707=>"111000100",
  34708=>"111111011",
  34709=>"110110100",
  34710=>"001101001",
  34711=>"101110010",
  34712=>"110011010",
  34713=>"101111111",
  34714=>"110010010",
  34715=>"101000000",
  34716=>"111100101",
  34717=>"100010011",
  34718=>"100111100",
  34719=>"000101110",
  34720=>"100100100",
  34721=>"111111111",
  34722=>"101110010",
  34723=>"101101001",
  34724=>"010111101",
  34725=>"110110111",
  34726=>"010110000",
  34727=>"000110110",
  34728=>"111000010",
  34729=>"101110001",
  34730=>"010111011",
  34731=>"111110110",
  34732=>"110100001",
  34733=>"101110111",
  34734=>"000110111",
  34735=>"000110100",
  34736=>"000101001",
  34737=>"110101110",
  34738=>"001111001",
  34739=>"110110101",
  34740=>"110101111",
  34741=>"011110011",
  34742=>"011100001",
  34743=>"001010001",
  34744=>"111010110",
  34745=>"001001000",
  34746=>"100010110",
  34747=>"001111011",
  34748=>"110111111",
  34749=>"101010011",
  34750=>"010001010",
  34751=>"100001000",
  34752=>"010111011",
  34753=>"101000101",
  34754=>"010101011",
  34755=>"111111111",
  34756=>"101101011",
  34757=>"100011111",
  34758=>"010001000",
  34759=>"000111001",
  34760=>"100111111",
  34761=>"100111001",
  34762=>"000010000",
  34763=>"111001100",
  34764=>"111001001",
  34765=>"001011101",
  34766=>"001101010",
  34767=>"010101110",
  34768=>"100010000",
  34769=>"101010000",
  34770=>"110111101",
  34771=>"010000011",
  34772=>"010000110",
  34773=>"111000011",
  34774=>"101001010",
  34775=>"111000100",
  34776=>"101100001",
  34777=>"100101111",
  34778=>"010000011",
  34779=>"000100000",
  34780=>"110100010",
  34781=>"101000110",
  34782=>"011101100",
  34783=>"111011010",
  34784=>"111011100",
  34785=>"011110001",
  34786=>"001000100",
  34787=>"110010110",
  34788=>"111101110",
  34789=>"001100000",
  34790=>"100110011",
  34791=>"010110010",
  34792=>"100011000",
  34793=>"010110000",
  34794=>"010110001",
  34795=>"011111000",
  34796=>"100010001",
  34797=>"100011100",
  34798=>"111100010",
  34799=>"010011110",
  34800=>"101101100",
  34801=>"000110000",
  34802=>"110111111",
  34803=>"010010101",
  34804=>"100000111",
  34805=>"000011000",
  34806=>"010100011",
  34807=>"000000000",
  34808=>"000001111",
  34809=>"110010100",
  34810=>"101100100",
  34811=>"001100010",
  34812=>"001100000",
  34813=>"011010000",
  34814=>"000111101",
  34815=>"100011111",
  34816=>"111100110",
  34817=>"101000101",
  34818=>"111101001",
  34819=>"100110011",
  34820=>"000101011",
  34821=>"000111110",
  34822=>"101110110",
  34823=>"011100010",
  34824=>"111000110",
  34825=>"110000110",
  34826=>"111101010",
  34827=>"111001011",
  34828=>"011100101",
  34829=>"101011011",
  34830=>"001001000",
  34831=>"000010001",
  34832=>"001001001",
  34833=>"111110010",
  34834=>"011010000",
  34835=>"101011100",
  34836=>"000011010",
  34837=>"010000001",
  34838=>"000100010",
  34839=>"000001000",
  34840=>"011101001",
  34841=>"011011010",
  34842=>"110111011",
  34843=>"100011000",
  34844=>"110111011",
  34845=>"000011100",
  34846=>"000001000",
  34847=>"101000100",
  34848=>"100000111",
  34849=>"000011101",
  34850=>"010110100",
  34851=>"001011001",
  34852=>"111010111",
  34853=>"111010010",
  34854=>"101001101",
  34855=>"010000011",
  34856=>"000110111",
  34857=>"001111000",
  34858=>"110001110",
  34859=>"110010011",
  34860=>"001110100",
  34861=>"010100100",
  34862=>"101011000",
  34863=>"100101001",
  34864=>"011011110",
  34865=>"001101111",
  34866=>"001010001",
  34867=>"111011000",
  34868=>"011001011",
  34869=>"111011010",
  34870=>"011110111",
  34871=>"101000010",
  34872=>"000000000",
  34873=>"110001110",
  34874=>"111100000",
  34875=>"111010101",
  34876=>"100000000",
  34877=>"000111111",
  34878=>"101110111",
  34879=>"000101011",
  34880=>"001110001",
  34881=>"110000000",
  34882=>"110010111",
  34883=>"010110101",
  34884=>"111110001",
  34885=>"010001111",
  34886=>"000101001",
  34887=>"110010011",
  34888=>"110010100",
  34889=>"011000101",
  34890=>"100110101",
  34891=>"000000010",
  34892=>"111101110",
  34893=>"100001100",
  34894=>"101101110",
  34895=>"110001000",
  34896=>"100001000",
  34897=>"110010111",
  34898=>"101101010",
  34899=>"101001011",
  34900=>"010010011",
  34901=>"111011011",
  34902=>"110011110",
  34903=>"101101001",
  34904=>"010110011",
  34905=>"010111000",
  34906=>"100010010",
  34907=>"110011111",
  34908=>"000100100",
  34909=>"001101100",
  34910=>"101111100",
  34911=>"001000011",
  34912=>"111110000",
  34913=>"000001000",
  34914=>"101110110",
  34915=>"000001111",
  34916=>"110001001",
  34917=>"010110011",
  34918=>"010110110",
  34919=>"001001001",
  34920=>"110010101",
  34921=>"011000111",
  34922=>"001111001",
  34923=>"010010000",
  34924=>"101100110",
  34925=>"000110110",
  34926=>"001001001",
  34927=>"001001010",
  34928=>"000111110",
  34929=>"001001000",
  34930=>"111110001",
  34931=>"011001111",
  34932=>"110010000",
  34933=>"001001110",
  34934=>"010110010",
  34935=>"111101101",
  34936=>"001110110",
  34937=>"011100111",
  34938=>"111010100",
  34939=>"100000100",
  34940=>"111011111",
  34941=>"101100100",
  34942=>"011011100",
  34943=>"010011011",
  34944=>"110001000",
  34945=>"001101011",
  34946=>"110111011",
  34947=>"111111110",
  34948=>"100111001",
  34949=>"000001000",
  34950=>"001001100",
  34951=>"110110101",
  34952=>"111010000",
  34953=>"001010010",
  34954=>"110100111",
  34955=>"100011011",
  34956=>"001100001",
  34957=>"011101101",
  34958=>"000010000",
  34959=>"110010011",
  34960=>"110011010",
  34961=>"000010010",
  34962=>"111010110",
  34963=>"111000110",
  34964=>"110000000",
  34965=>"011111110",
  34966=>"100000010",
  34967=>"000001001",
  34968=>"110111100",
  34969=>"010110001",
  34970=>"000111111",
  34971=>"011001000",
  34972=>"011101010",
  34973=>"101101101",
  34974=>"111000011",
  34975=>"101000001",
  34976=>"111011001",
  34977=>"001111001",
  34978=>"111000011",
  34979=>"010010111",
  34980=>"010110010",
  34981=>"000010101",
  34982=>"001110011",
  34983=>"001011101",
  34984=>"111011110",
  34985=>"110110000",
  34986=>"111010000",
  34987=>"100010110",
  34988=>"000111001",
  34989=>"101110001",
  34990=>"000100001",
  34991=>"001010111",
  34992=>"111100011",
  34993=>"110100101",
  34994=>"001000101",
  34995=>"100001001",
  34996=>"010010001",
  34997=>"111001000",
  34998=>"011010011",
  34999=>"011001100",
  35000=>"111111011",
  35001=>"010110110",
  35002=>"101000010",
  35003=>"101110011",
  35004=>"000011000",
  35005=>"010011110",
  35006=>"010000000",
  35007=>"010000001",
  35008=>"010110101",
  35009=>"000000110",
  35010=>"011011011",
  35011=>"101100010",
  35012=>"101011110",
  35013=>"011001100",
  35014=>"011011100",
  35015=>"011000101",
  35016=>"101110011",
  35017=>"010111101",
  35018=>"101100010",
  35019=>"111001110",
  35020=>"000111101",
  35021=>"101011100",
  35022=>"111000111",
  35023=>"100011111",
  35024=>"100000001",
  35025=>"000000000",
  35026=>"101111110",
  35027=>"001100010",
  35028=>"001001011",
  35029=>"000110111",
  35030=>"111101101",
  35031=>"101101011",
  35032=>"001001001",
  35033=>"110010010",
  35034=>"100111110",
  35035=>"001001110",
  35036=>"111001010",
  35037=>"111110010",
  35038=>"101101110",
  35039=>"101011100",
  35040=>"110111111",
  35041=>"111111111",
  35042=>"101100100",
  35043=>"100111010",
  35044=>"100101000",
  35045=>"011000000",
  35046=>"001111111",
  35047=>"110010001",
  35048=>"111011000",
  35049=>"000110000",
  35050=>"001100000",
  35051=>"100000001",
  35052=>"101110001",
  35053=>"110101111",
  35054=>"010010110",
  35055=>"111001011",
  35056=>"010010110",
  35057=>"001001010",
  35058=>"001111000",
  35059=>"000110011",
  35060=>"110001000",
  35061=>"010110000",
  35062=>"011010011",
  35063=>"101000110",
  35064=>"101001010",
  35065=>"101001111",
  35066=>"100111000",
  35067=>"100000001",
  35068=>"011100001",
  35069=>"001001110",
  35070=>"101100101",
  35071=>"011111001",
  35072=>"110000100",
  35073=>"010100000",
  35074=>"101000011",
  35075=>"110001111",
  35076=>"000101101",
  35077=>"001101100",
  35078=>"100100010",
  35079=>"111111100",
  35080=>"100111000",
  35081=>"111010011",
  35082=>"010010111",
  35083=>"010101010",
  35084=>"011000000",
  35085=>"110111001",
  35086=>"010001010",
  35087=>"010000011",
  35088=>"010111000",
  35089=>"011111011",
  35090=>"100111111",
  35091=>"010011100",
  35092=>"001110111",
  35093=>"001000001",
  35094=>"101011000",
  35095=>"110000011",
  35096=>"100001011",
  35097=>"000100110",
  35098=>"010010100",
  35099=>"100111110",
  35100=>"011100001",
  35101=>"000011000",
  35102=>"100001110",
  35103=>"000010010",
  35104=>"010101111",
  35105=>"011100000",
  35106=>"111010001",
  35107=>"001000110",
  35108=>"110000011",
  35109=>"000110000",
  35110=>"100000010",
  35111=>"000011001",
  35112=>"111001111",
  35113=>"111101001",
  35114=>"000110110",
  35115=>"001000100",
  35116=>"000101000",
  35117=>"101101101",
  35118=>"011010010",
  35119=>"100001001",
  35120=>"011101000",
  35121=>"011010101",
  35122=>"111111011",
  35123=>"100110111",
  35124=>"001111011",
  35125=>"110001111",
  35126=>"000010001",
  35127=>"111110110",
  35128=>"010001101",
  35129=>"111001011",
  35130=>"010011101",
  35131=>"010110111",
  35132=>"101101100",
  35133=>"101011010",
  35134=>"011100110",
  35135=>"010100110",
  35136=>"000111000",
  35137=>"101000000",
  35138=>"101001010",
  35139=>"110001110",
  35140=>"001100001",
  35141=>"111001001",
  35142=>"001000001",
  35143=>"010110001",
  35144=>"110001111",
  35145=>"110000010",
  35146=>"000010110",
  35147=>"001110101",
  35148=>"010010000",
  35149=>"100000100",
  35150=>"111111011",
  35151=>"111011100",
  35152=>"110001001",
  35153=>"110111111",
  35154=>"111001111",
  35155=>"110110010",
  35156=>"110010001",
  35157=>"100011110",
  35158=>"111011000",
  35159=>"111101111",
  35160=>"000000010",
  35161=>"000000011",
  35162=>"110110101",
  35163=>"100001100",
  35164=>"010110101",
  35165=>"100000011",
  35166=>"110010101",
  35167=>"001100101",
  35168=>"010111111",
  35169=>"110110100",
  35170=>"101001010",
  35171=>"000110000",
  35172=>"010011101",
  35173=>"001001110",
  35174=>"110001110",
  35175=>"100000010",
  35176=>"010111101",
  35177=>"100110000",
  35178=>"110011110",
  35179=>"010001101",
  35180=>"011101001",
  35181=>"011001111",
  35182=>"100101101",
  35183=>"101101100",
  35184=>"100010010",
  35185=>"010100011",
  35186=>"110111100",
  35187=>"011000110",
  35188=>"111000110",
  35189=>"110110011",
  35190=>"000111010",
  35191=>"010111000",
  35192=>"001111001",
  35193=>"000100110",
  35194=>"100001000",
  35195=>"001000011",
  35196=>"001100101",
  35197=>"111011001",
  35198=>"110010101",
  35199=>"011011001",
  35200=>"100110011",
  35201=>"100101101",
  35202=>"000001010",
  35203=>"001001001",
  35204=>"111101101",
  35205=>"000011001",
  35206=>"101011000",
  35207=>"001000000",
  35208=>"001111110",
  35209=>"010011000",
  35210=>"010001101",
  35211=>"010011010",
  35212=>"101101001",
  35213=>"000001111",
  35214=>"100001100",
  35215=>"001000011",
  35216=>"001010000",
  35217=>"011000011",
  35218=>"101011000",
  35219=>"000010000",
  35220=>"000010010",
  35221=>"001010101",
  35222=>"101100110",
  35223=>"011010101",
  35224=>"101101101",
  35225=>"001100010",
  35226=>"010111101",
  35227=>"110010011",
  35228=>"111111001",
  35229=>"111010010",
  35230=>"111001000",
  35231=>"111100011",
  35232=>"000111101",
  35233=>"011101001",
  35234=>"110011010",
  35235=>"000011100",
  35236=>"001100011",
  35237=>"000010101",
  35238=>"001110011",
  35239=>"110000101",
  35240=>"010110000",
  35241=>"011100101",
  35242=>"000010010",
  35243=>"011000110",
  35244=>"000100001",
  35245=>"011010011",
  35246=>"001111101",
  35247=>"011111001",
  35248=>"101001100",
  35249=>"111101011",
  35250=>"011001110",
  35251=>"111010001",
  35252=>"010110110",
  35253=>"100011010",
  35254=>"000110010",
  35255=>"101100000",
  35256=>"011000011",
  35257=>"010010000",
  35258=>"100011011",
  35259=>"101110101",
  35260=>"111000010",
  35261=>"001010101",
  35262=>"011100100",
  35263=>"010010110",
  35264=>"001010010",
  35265=>"110011110",
  35266=>"010000001",
  35267=>"100101110",
  35268=>"000011011",
  35269=>"011000100",
  35270=>"111011100",
  35271=>"101100001",
  35272=>"011111011",
  35273=>"111001110",
  35274=>"111001100",
  35275=>"001110100",
  35276=>"101101001",
  35277=>"101011110",
  35278=>"010111010",
  35279=>"101100101",
  35280=>"011111111",
  35281=>"011011100",
  35282=>"110000110",
  35283=>"001111111",
  35284=>"100000010",
  35285=>"011110011",
  35286=>"010010000",
  35287=>"001111100",
  35288=>"100100101",
  35289=>"100000000",
  35290=>"111111001",
  35291=>"000011001",
  35292=>"001001100",
  35293=>"010001100",
  35294=>"101110100",
  35295=>"101110010",
  35296=>"000111111",
  35297=>"001100111",
  35298=>"111110101",
  35299=>"101100101",
  35300=>"100011001",
  35301=>"101101110",
  35302=>"010001101",
  35303=>"101011000",
  35304=>"010000011",
  35305=>"110010000",
  35306=>"001101000",
  35307=>"101111111",
  35308=>"010110000",
  35309=>"011111001",
  35310=>"010100001",
  35311=>"111001000",
  35312=>"101000101",
  35313=>"100110100",
  35314=>"000011111",
  35315=>"101101101",
  35316=>"101010101",
  35317=>"101011011",
  35318=>"111001011",
  35319=>"000110001",
  35320=>"010101000",
  35321=>"110101011",
  35322=>"001101011",
  35323=>"010001010",
  35324=>"001010011",
  35325=>"101101000",
  35326=>"001011011",
  35327=>"101110011",
  35328=>"111011010",
  35329=>"011000001",
  35330=>"101110010",
  35331=>"000010000",
  35332=>"011111001",
  35333=>"111011001",
  35334=>"111111100",
  35335=>"000000110",
  35336=>"001010101",
  35337=>"011000000",
  35338=>"101000100",
  35339=>"000010010",
  35340=>"001111111",
  35341=>"101000100",
  35342=>"101001111",
  35343=>"000111110",
  35344=>"000000000",
  35345=>"011101100",
  35346=>"101011000",
  35347=>"100001111",
  35348=>"110011101",
  35349=>"000010010",
  35350=>"000100110",
  35351=>"101110100",
  35352=>"010110100",
  35353=>"011010101",
  35354=>"110010010",
  35355=>"010100111",
  35356=>"000011110",
  35357=>"111010001",
  35358=>"100010100",
  35359=>"000101010",
  35360=>"100001101",
  35361=>"110111010",
  35362=>"000101100",
  35363=>"011111111",
  35364=>"100101101",
  35365=>"000110011",
  35366=>"010111010",
  35367=>"011100110",
  35368=>"111000010",
  35369=>"001110110",
  35370=>"010011111",
  35371=>"100000010",
  35372=>"010010010",
  35373=>"110001001",
  35374=>"100100011",
  35375=>"010001110",
  35376=>"110111100",
  35377=>"101101001",
  35378=>"011101111",
  35379=>"111100000",
  35380=>"100000111",
  35381=>"111100010",
  35382=>"100011110",
  35383=>"111111011",
  35384=>"000110000",
  35385=>"000100011",
  35386=>"100000101",
  35387=>"101000100",
  35388=>"011100110",
  35389=>"011110000",
  35390=>"010000101",
  35391=>"100001100",
  35392=>"101011011",
  35393=>"011001100",
  35394=>"000000001",
  35395=>"000101100",
  35396=>"011111101",
  35397=>"000100000",
  35398=>"100111101",
  35399=>"111110000",
  35400=>"101111101",
  35401=>"110101011",
  35402=>"110001010",
  35403=>"100100011",
  35404=>"000000100",
  35405=>"010100010",
  35406=>"111011010",
  35407=>"001010111",
  35408=>"111001100",
  35409=>"101011100",
  35410=>"100110111",
  35411=>"000100100",
  35412=>"010010000",
  35413=>"000011011",
  35414=>"100000000",
  35415=>"011101011",
  35416=>"011110111",
  35417=>"001100001",
  35418=>"111011000",
  35419=>"101011010",
  35420=>"000000100",
  35421=>"011101000",
  35422=>"000011111",
  35423=>"101011010",
  35424=>"011110000",
  35425=>"011000101",
  35426=>"101010011",
  35427=>"011001010",
  35428=>"001001011",
  35429=>"100100101",
  35430=>"101001001",
  35431=>"111010001",
  35432=>"010110100",
  35433=>"000010101",
  35434=>"000011001",
  35435=>"111001100",
  35436=>"001000111",
  35437=>"011001001",
  35438=>"010101010",
  35439=>"000111100",
  35440=>"101001001",
  35441=>"010011010",
  35442=>"111100001",
  35443=>"110010001",
  35444=>"010011001",
  35445=>"100001110",
  35446=>"100100100",
  35447=>"000110001",
  35448=>"000100101",
  35449=>"110011011",
  35450=>"111110010",
  35451=>"000001001",
  35452=>"001101001",
  35453=>"001100110",
  35454=>"010010110",
  35455=>"011001101",
  35456=>"111010100",
  35457=>"101101110",
  35458=>"000110010",
  35459=>"101000001",
  35460=>"010111111",
  35461=>"000011001",
  35462=>"000111001",
  35463=>"110001111",
  35464=>"000011110",
  35465=>"000010100",
  35466=>"101010100",
  35467=>"011000001",
  35468=>"011001111",
  35469=>"010000111",
  35470=>"100000001",
  35471=>"011011000",
  35472=>"010101000",
  35473=>"100100101",
  35474=>"100010000",
  35475=>"010010010",
  35476=>"101011111",
  35477=>"100011100",
  35478=>"110110010",
  35479=>"010110000",
  35480=>"111101111",
  35481=>"101101010",
  35482=>"111100110",
  35483=>"010011111",
  35484=>"111111111",
  35485=>"010010111",
  35486=>"000001001",
  35487=>"000010011",
  35488=>"011010000",
  35489=>"100000011",
  35490=>"111011010",
  35491=>"100111011",
  35492=>"101101011",
  35493=>"101111010",
  35494=>"111010001",
  35495=>"000101010",
  35496=>"100111100",
  35497=>"110000111",
  35498=>"101010100",
  35499=>"110100000",
  35500=>"010000110",
  35501=>"100001010",
  35502=>"010001100",
  35503=>"110111000",
  35504=>"000111001",
  35505=>"101101010",
  35506=>"000011101",
  35507=>"110110001",
  35508=>"001000111",
  35509=>"000000110",
  35510=>"100010110",
  35511=>"010101101",
  35512=>"101011100",
  35513=>"001010110",
  35514=>"111101100",
  35515=>"001001111",
  35516=>"101001111",
  35517=>"000000001",
  35518=>"110000011",
  35519=>"010010010",
  35520=>"011010001",
  35521=>"101101000",
  35522=>"011000011",
  35523=>"001100101",
  35524=>"010100111",
  35525=>"001001000",
  35526=>"010000001",
  35527=>"001001001",
  35528=>"101000010",
  35529=>"011100111",
  35530=>"011101100",
  35531=>"110000011",
  35532=>"010000111",
  35533=>"000110011",
  35534=>"010001110",
  35535=>"011101001",
  35536=>"110010110",
  35537=>"011101100",
  35538=>"100100100",
  35539=>"011111011",
  35540=>"011011001",
  35541=>"000010011",
  35542=>"101101010",
  35543=>"001100110",
  35544=>"110011000",
  35545=>"100000010",
  35546=>"000000001",
  35547=>"111100001",
  35548=>"001101111",
  35549=>"000001100",
  35550=>"000010100",
  35551=>"110111111",
  35552=>"111100101",
  35553=>"011000010",
  35554=>"001001111",
  35555=>"000001110",
  35556=>"000010101",
  35557=>"100101111",
  35558=>"011111111",
  35559=>"111110101",
  35560=>"011100011",
  35561=>"100101000",
  35562=>"110101101",
  35563=>"111000011",
  35564=>"010011000",
  35565=>"110000101",
  35566=>"010100011",
  35567=>"101001010",
  35568=>"110011110",
  35569=>"110100001",
  35570=>"100111000",
  35571=>"101101000",
  35572=>"100101111",
  35573=>"110000001",
  35574=>"111101011",
  35575=>"110110110",
  35576=>"010111101",
  35577=>"101100010",
  35578=>"100011001",
  35579=>"100010011",
  35580=>"100100110",
  35581=>"100000011",
  35582=>"001101110",
  35583=>"101100100",
  35584=>"001100101",
  35585=>"011011001",
  35586=>"000000001",
  35587=>"110101010",
  35588=>"110011011",
  35589=>"100001110",
  35590=>"010000010",
  35591=>"111100111",
  35592=>"000100001",
  35593=>"110100101",
  35594=>"110001111",
  35595=>"011100001",
  35596=>"001001110",
  35597=>"110111010",
  35598=>"011111111",
  35599=>"100110110",
  35600=>"101110010",
  35601=>"000001011",
  35602=>"111011100",
  35603=>"100110010",
  35604=>"101101111",
  35605=>"111110011",
  35606=>"110000010",
  35607=>"001000000",
  35608=>"100001011",
  35609=>"100111110",
  35610=>"010110101",
  35611=>"010111011",
  35612=>"011011101",
  35613=>"100110001",
  35614=>"111000110",
  35615=>"011100100",
  35616=>"000111010",
  35617=>"011010110",
  35618=>"000110110",
  35619=>"001001111",
  35620=>"110000100",
  35621=>"110011010",
  35622=>"001001110",
  35623=>"011101000",
  35624=>"111111011",
  35625=>"110010111",
  35626=>"110110110",
  35627=>"100111111",
  35628=>"110011110",
  35629=>"001001101",
  35630=>"001110111",
  35631=>"100011000",
  35632=>"110011101",
  35633=>"100100001",
  35634=>"011010011",
  35635=>"111011001",
  35636=>"111100101",
  35637=>"110101101",
  35638=>"101100000",
  35639=>"111010100",
  35640=>"001000000",
  35641=>"000111011",
  35642=>"101111010",
  35643=>"111000101",
  35644=>"000011111",
  35645=>"010010110",
  35646=>"110001001",
  35647=>"100101010",
  35648=>"101010010",
  35649=>"100100111",
  35650=>"100110111",
  35651=>"111101101",
  35652=>"100101110",
  35653=>"110000011",
  35654=>"111000111",
  35655=>"100001101",
  35656=>"010100110",
  35657=>"110100010",
  35658=>"110000000",
  35659=>"011110010",
  35660=>"001011110",
  35661=>"110111001",
  35662=>"011110000",
  35663=>"011111001",
  35664=>"010000010",
  35665=>"010110001",
  35666=>"110011100",
  35667=>"100100011",
  35668=>"100110001",
  35669=>"011010001",
  35670=>"100001110",
  35671=>"111000001",
  35672=>"010111010",
  35673=>"001010001",
  35674=>"110111100",
  35675=>"001001000",
  35676=>"110010000",
  35677=>"100100001",
  35678=>"000100001",
  35679=>"000101111",
  35680=>"011001010",
  35681=>"110110100",
  35682=>"000000010",
  35683=>"110010101",
  35684=>"100101010",
  35685=>"010111111",
  35686=>"101011101",
  35687=>"101010010",
  35688=>"100001101",
  35689=>"010001110",
  35690=>"000011100",
  35691=>"010110111",
  35692=>"111011101",
  35693=>"011101001",
  35694=>"100011100",
  35695=>"000110110",
  35696=>"111011010",
  35697=>"010001011",
  35698=>"100000000",
  35699=>"101011100",
  35700=>"000001000",
  35701=>"001101110",
  35702=>"010011010",
  35703=>"111001011",
  35704=>"101100011",
  35705=>"010011010",
  35706=>"110111010",
  35707=>"000000001",
  35708=>"110100010",
  35709=>"101011111",
  35710=>"011101111",
  35711=>"110001110",
  35712=>"101110101",
  35713=>"111000111",
  35714=>"000001000",
  35715=>"010010000",
  35716=>"010001111",
  35717=>"001111001",
  35718=>"010011000",
  35719=>"100000101",
  35720=>"100101011",
  35721=>"011101001",
  35722=>"010010101",
  35723=>"100111110",
  35724=>"111000111",
  35725=>"101011101",
  35726=>"101101100",
  35727=>"111101101",
  35728=>"001101101",
  35729=>"011010111",
  35730=>"001101110",
  35731=>"111011001",
  35732=>"011101100",
  35733=>"001100100",
  35734=>"110101111",
  35735=>"001101100",
  35736=>"011111110",
  35737=>"000111010",
  35738=>"001011000",
  35739=>"000010011",
  35740=>"100111111",
  35741=>"111111101",
  35742=>"111110001",
  35743=>"010001101",
  35744=>"110001100",
  35745=>"000110110",
  35746=>"011100000",
  35747=>"010000011",
  35748=>"010010110",
  35749=>"010111110",
  35750=>"100000101",
  35751=>"111000111",
  35752=>"011000110",
  35753=>"111101010",
  35754=>"000001111",
  35755=>"100110100",
  35756=>"111100110",
  35757=>"000100110",
  35758=>"110001101",
  35759=>"011100101",
  35760=>"100110101",
  35761=>"001100101",
  35762=>"001111001",
  35763=>"000110001",
  35764=>"101110100",
  35765=>"101000001",
  35766=>"100110010",
  35767=>"101101101",
  35768=>"011101000",
  35769=>"011001001",
  35770=>"011001111",
  35771=>"100011100",
  35772=>"101111011",
  35773=>"011010101",
  35774=>"011001011",
  35775=>"010010111",
  35776=>"000010011",
  35777=>"100110001",
  35778=>"011110011",
  35779=>"011000000",
  35780=>"010101111",
  35781=>"011010111",
  35782=>"111101100",
  35783=>"111010000",
  35784=>"100001011",
  35785=>"001010001",
  35786=>"101110100",
  35787=>"101011001",
  35788=>"000110110",
  35789=>"011111011",
  35790=>"001111011",
  35791=>"011101100",
  35792=>"011011111",
  35793=>"010000000",
  35794=>"110110010",
  35795=>"000001111",
  35796=>"100011101",
  35797=>"100100010",
  35798=>"001001100",
  35799=>"101010001",
  35800=>"110000101",
  35801=>"000000111",
  35802=>"001100100",
  35803=>"110101101",
  35804=>"011110000",
  35805=>"111101000",
  35806=>"101100000",
  35807=>"110100100",
  35808=>"000001111",
  35809=>"101011111",
  35810=>"011111110",
  35811=>"100111110",
  35812=>"111110010",
  35813=>"001100100",
  35814=>"100111011",
  35815=>"100100111",
  35816=>"000001101",
  35817=>"010110000",
  35818=>"101000100",
  35819=>"100100110",
  35820=>"100100111",
  35821=>"111101100",
  35822=>"010111100",
  35823=>"000110110",
  35824=>"011000111",
  35825=>"110111011",
  35826=>"100110110",
  35827=>"101110111",
  35828=>"010100110",
  35829=>"101100100",
  35830=>"111010110",
  35831=>"001101001",
  35832=>"000011011",
  35833=>"100101100",
  35834=>"001011010",
  35835=>"110000111",
  35836=>"110100101",
  35837=>"111010101",
  35838=>"101010100",
  35839=>"000001011",
  35840=>"110010011",
  35841=>"010000000",
  35842=>"111001000",
  35843=>"111101010",
  35844=>"000011011",
  35845=>"100110100",
  35846=>"111100000",
  35847=>"010110111",
  35848=>"110010111",
  35849=>"101110001",
  35850=>"111011000",
  35851=>"111001110",
  35852=>"100010011",
  35853=>"000111110",
  35854=>"000110101",
  35855=>"001101111",
  35856=>"011101111",
  35857=>"111011001",
  35858=>"111010111",
  35859=>"101001001",
  35860=>"000100101",
  35861=>"110001000",
  35862=>"011000111",
  35863=>"111110010",
  35864=>"000110100",
  35865=>"000110111",
  35866=>"110000000",
  35867=>"111100010",
  35868=>"000110001",
  35869=>"111110001",
  35870=>"001010010",
  35871=>"100100001",
  35872=>"000010111",
  35873=>"011110100",
  35874=>"011000001",
  35875=>"100110000",
  35876=>"011111110",
  35877=>"111110101",
  35878=>"100001100",
  35879=>"100000000",
  35880=>"110011110",
  35881=>"010011010",
  35882=>"010001010",
  35883=>"010100110",
  35884=>"011100001",
  35885=>"110101010",
  35886=>"110101010",
  35887=>"110101001",
  35888=>"100010110",
  35889=>"111110100",
  35890=>"100010000",
  35891=>"011011011",
  35892=>"100010010",
  35893=>"011100001",
  35894=>"010010110",
  35895=>"101000001",
  35896=>"010000100",
  35897=>"111100000",
  35898=>"110011111",
  35899=>"000001100",
  35900=>"100011111",
  35901=>"100100001",
  35902=>"100001111",
  35903=>"100110110",
  35904=>"111100100",
  35905=>"100111000",
  35906=>"101111101",
  35907=>"100100111",
  35908=>"111001101",
  35909=>"000110010",
  35910=>"111001101",
  35911=>"111100011",
  35912=>"001111001",
  35913=>"100100011",
  35914=>"110110001",
  35915=>"100000000",
  35916=>"110101011",
  35917=>"001010010",
  35918=>"110101111",
  35919=>"010111111",
  35920=>"011011011",
  35921=>"010111100",
  35922=>"000011001",
  35923=>"110100001",
  35924=>"011110110",
  35925=>"100011010",
  35926=>"001001011",
  35927=>"010010100",
  35928=>"000000100",
  35929=>"011101101",
  35930=>"001110101",
  35931=>"000100100",
  35932=>"101011000",
  35933=>"101100110",
  35934=>"000110111",
  35935=>"000110101",
  35936=>"000000101",
  35937=>"101101001",
  35938=>"100110100",
  35939=>"100101110",
  35940=>"000101001",
  35941=>"011101010",
  35942=>"000001010",
  35943=>"000011010",
  35944=>"110111001",
  35945=>"110011110",
  35946=>"001000111",
  35947=>"111110110",
  35948=>"011010111",
  35949=>"000001010",
  35950=>"101111011",
  35951=>"000011011",
  35952=>"001010000",
  35953=>"001000011",
  35954=>"010000011",
  35955=>"001111111",
  35956=>"001010000",
  35957=>"000110001",
  35958=>"101011000",
  35959=>"101110011",
  35960=>"010110010",
  35961=>"000111100",
  35962=>"001101111",
  35963=>"110001101",
  35964=>"101111011",
  35965=>"110100101",
  35966=>"000110000",
  35967=>"011111010",
  35968=>"111011111",
  35969=>"111011110",
  35970=>"010110110",
  35971=>"101011100",
  35972=>"001000000",
  35973=>"001101000",
  35974=>"100111111",
  35975=>"000100110",
  35976=>"001010011",
  35977=>"100000011",
  35978=>"111000111",
  35979=>"011111010",
  35980=>"101010000",
  35981=>"000010000",
  35982=>"000001110",
  35983=>"100000010",
  35984=>"110011000",
  35985=>"101111101",
  35986=>"001111000",
  35987=>"010101101",
  35988=>"111000111",
  35989=>"000011010",
  35990=>"110001010",
  35991=>"010110100",
  35992=>"000000110",
  35993=>"010111000",
  35994=>"010110011",
  35995=>"000010001",
  35996=>"000000100",
  35997=>"011101011",
  35998=>"000001010",
  35999=>"001001111",
  36000=>"011001000",
  36001=>"000110000",
  36002=>"000101100",
  36003=>"100101110",
  36004=>"100101100",
  36005=>"111011111",
  36006=>"000010010",
  36007=>"010000011",
  36008=>"010011110",
  36009=>"100110110",
  36010=>"000101111",
  36011=>"011010110",
  36012=>"000111100",
  36013=>"010011000",
  36014=>"100101000",
  36015=>"011010010",
  36016=>"011010001",
  36017=>"101101001",
  36018=>"110100100",
  36019=>"111111110",
  36020=>"100011010",
  36021=>"010100000",
  36022=>"110100111",
  36023=>"001101011",
  36024=>"101010111",
  36025=>"100111100",
  36026=>"110110010",
  36027=>"000010111",
  36028=>"101110110",
  36029=>"101000010",
  36030=>"100111110",
  36031=>"101100010",
  36032=>"110101111",
  36033=>"000101110",
  36034=>"001001010",
  36035=>"001111110",
  36036=>"110011111",
  36037=>"000110011",
  36038=>"000000110",
  36039=>"000010111",
  36040=>"010110001",
  36041=>"101000100",
  36042=>"101010000",
  36043=>"000001000",
  36044=>"111111000",
  36045=>"011101000",
  36046=>"110100001",
  36047=>"100011100",
  36048=>"111110001",
  36049=>"110101100",
  36050=>"101000100",
  36051=>"101010101",
  36052=>"011101001",
  36053=>"010010101",
  36054=>"111110110",
  36055=>"101000001",
  36056=>"001000010",
  36057=>"110100001",
  36058=>"110100001",
  36059=>"110000111",
  36060=>"000011100",
  36061=>"010110100",
  36062=>"000011011",
  36063=>"111000110",
  36064=>"000000100",
  36065=>"110111001",
  36066=>"100110000",
  36067=>"010111111",
  36068=>"000011100",
  36069=>"011111101",
  36070=>"011001110",
  36071=>"111011011",
  36072=>"100100000",
  36073=>"111010100",
  36074=>"000001010",
  36075=>"110001000",
  36076=>"010110000",
  36077=>"011101110",
  36078=>"011111000",
  36079=>"010110101",
  36080=>"011001010",
  36081=>"101011111",
  36082=>"001101010",
  36083=>"001011001",
  36084=>"100111111",
  36085=>"010001001",
  36086=>"111010011",
  36087=>"111110111",
  36088=>"101001000",
  36089=>"111100001",
  36090=>"101101110",
  36091=>"111110011",
  36092=>"110111101",
  36093=>"110101000",
  36094=>"101101100",
  36095=>"010110011",
  36096=>"101101011",
  36097=>"011000001",
  36098=>"100001001",
  36099=>"100011011",
  36100=>"110010000",
  36101=>"001001000",
  36102=>"111001111",
  36103=>"100000100",
  36104=>"000000000",
  36105=>"001100011",
  36106=>"111010100",
  36107=>"101100010",
  36108=>"101110001",
  36109=>"100111100",
  36110=>"110000101",
  36111=>"001101100",
  36112=>"110001001",
  36113=>"101101001",
  36114=>"000011111",
  36115=>"111111000",
  36116=>"001111100",
  36117=>"001010100",
  36118=>"100111101",
  36119=>"011011010",
  36120=>"001010010",
  36121=>"000100111",
  36122=>"100011101",
  36123=>"000101110",
  36124=>"001111110",
  36125=>"001000001",
  36126=>"011001110",
  36127=>"001011011",
  36128=>"000001111",
  36129=>"010110101",
  36130=>"100100000",
  36131=>"011110011",
  36132=>"110110001",
  36133=>"100010001",
  36134=>"100001000",
  36135=>"000101010",
  36136=>"000000000",
  36137=>"110110100",
  36138=>"100010011",
  36139=>"110100001",
  36140=>"110110000",
  36141=>"000011101",
  36142=>"011111101",
  36143=>"001001101",
  36144=>"001100011",
  36145=>"000101111",
  36146=>"010010000",
  36147=>"111001001",
  36148=>"010011001",
  36149=>"100000100",
  36150=>"010110000",
  36151=>"101111110",
  36152=>"110011101",
  36153=>"110111000",
  36154=>"001101000",
  36155=>"110001101",
  36156=>"001101010",
  36157=>"001100110",
  36158=>"001100100",
  36159=>"111000110",
  36160=>"010110011",
  36161=>"010111001",
  36162=>"010110110",
  36163=>"111111001",
  36164=>"010010000",
  36165=>"001100111",
  36166=>"001010010",
  36167=>"111100100",
  36168=>"110010111",
  36169=>"011011111",
  36170=>"111110101",
  36171=>"110010001",
  36172=>"111100001",
  36173=>"001111001",
  36174=>"111011111",
  36175=>"111011101",
  36176=>"001110111",
  36177=>"110001011",
  36178=>"000110001",
  36179=>"110010010",
  36180=>"111000010",
  36181=>"011111111",
  36182=>"011111000",
  36183=>"110000111",
  36184=>"100110000",
  36185=>"101101101",
  36186=>"101001100",
  36187=>"101010101",
  36188=>"111000110",
  36189=>"100111011",
  36190=>"010010000",
  36191=>"011110111",
  36192=>"110111000",
  36193=>"010111000",
  36194=>"000110111",
  36195=>"011011010",
  36196=>"011100100",
  36197=>"000101010",
  36198=>"010010001",
  36199=>"111001111",
  36200=>"001001000",
  36201=>"000011011",
  36202=>"111111011",
  36203=>"110110001",
  36204=>"011010000",
  36205=>"111100011",
  36206=>"101000010",
  36207=>"111110000",
  36208=>"110001110",
  36209=>"110100000",
  36210=>"111011111",
  36211=>"101111000",
  36212=>"111110111",
  36213=>"001101000",
  36214=>"010111111",
  36215=>"011011001",
  36216=>"001101111",
  36217=>"000100101",
  36218=>"011001110",
  36219=>"111111110",
  36220=>"001010011",
  36221=>"000001000",
  36222=>"001111001",
  36223=>"000011001",
  36224=>"000010000",
  36225=>"000010000",
  36226=>"111001101",
  36227=>"111010110",
  36228=>"110011101",
  36229=>"000000010",
  36230=>"001100011",
  36231=>"001011111",
  36232=>"001101001",
  36233=>"000100101",
  36234=>"110110110",
  36235=>"000101100",
  36236=>"010101011",
  36237=>"001110000",
  36238=>"111110101",
  36239=>"100110010",
  36240=>"100010010",
  36241=>"110001000",
  36242=>"001010011",
  36243=>"100111110",
  36244=>"000010000",
  36245=>"001111010",
  36246=>"101111111",
  36247=>"101001001",
  36248=>"111010111",
  36249=>"101011111",
  36250=>"111111110",
  36251=>"000111111",
  36252=>"100110010",
  36253=>"101001011",
  36254=>"010010111",
  36255=>"111111110",
  36256=>"101110100",
  36257=>"000101011",
  36258=>"001010001",
  36259=>"100000000",
  36260=>"010010011",
  36261=>"011000101",
  36262=>"010111010",
  36263=>"010100111",
  36264=>"101011101",
  36265=>"010100011",
  36266=>"101010000",
  36267=>"011000001",
  36268=>"111101001",
  36269=>"001011110",
  36270=>"000010000",
  36271=>"110000001",
  36272=>"010000001",
  36273=>"110000100",
  36274=>"100001010",
  36275=>"001011111",
  36276=>"110010000",
  36277=>"110110000",
  36278=>"010010011",
  36279=>"001110000",
  36280=>"010001101",
  36281=>"101010100",
  36282=>"110010010",
  36283=>"110111100",
  36284=>"110111111",
  36285=>"101001000",
  36286=>"100010110",
  36287=>"010001100",
  36288=>"000001000",
  36289=>"100011000",
  36290=>"000111110",
  36291=>"101000101",
  36292=>"000100000",
  36293=>"110001001",
  36294=>"110111011",
  36295=>"000110111",
  36296=>"010011000",
  36297=>"010100111",
  36298=>"100110100",
  36299=>"101111111",
  36300=>"111010101",
  36301=>"111001001",
  36302=>"100010001",
  36303=>"111010010",
  36304=>"101010000",
  36305=>"111111110",
  36306=>"100101111",
  36307=>"110110100",
  36308=>"001101010",
  36309=>"100110010",
  36310=>"001101000",
  36311=>"110000010",
  36312=>"101001101",
  36313=>"111011110",
  36314=>"110111001",
  36315=>"111111110",
  36316=>"100011110",
  36317=>"110100100",
  36318=>"000110111",
  36319=>"001110101",
  36320=>"011111000",
  36321=>"001111011",
  36322=>"100111100",
  36323=>"010000011",
  36324=>"010001110",
  36325=>"111010101",
  36326=>"001011101",
  36327=>"100100010",
  36328=>"110010101",
  36329=>"011011001",
  36330=>"111110011",
  36331=>"111110010",
  36332=>"010111001",
  36333=>"011101000",
  36334=>"010000101",
  36335=>"000000010",
  36336=>"101101100",
  36337=>"011100101",
  36338=>"111101000",
  36339=>"101100010",
  36340=>"100001110",
  36341=>"010110110",
  36342=>"001011001",
  36343=>"000001100",
  36344=>"110001110",
  36345=>"000000100",
  36346=>"011111110",
  36347=>"010000010",
  36348=>"111111110",
  36349=>"111010111",
  36350=>"000101111",
  36351=>"111010111",
  36352=>"100001101",
  36353=>"100010001",
  36354=>"010011111",
  36355=>"010111000",
  36356=>"000111000",
  36357=>"100111000",
  36358=>"000001111",
  36359=>"000001101",
  36360=>"011000101",
  36361=>"010010100",
  36362=>"000111010",
  36363=>"110011101",
  36364=>"100101110",
  36365=>"001110111",
  36366=>"011111010",
  36367=>"110100101",
  36368=>"010011100",
  36369=>"101111101",
  36370=>"010000101",
  36371=>"010000110",
  36372=>"001101101",
  36373=>"010101010",
  36374=>"111011111",
  36375=>"001111001",
  36376=>"111101000",
  36377=>"100000111",
  36378=>"000001001",
  36379=>"001111110",
  36380=>"110110010",
  36381=>"110010000",
  36382=>"110110110",
  36383=>"111111111",
  36384=>"001110100",
  36385=>"100101111",
  36386=>"000010001",
  36387=>"100100000",
  36388=>"101111100",
  36389=>"101000100",
  36390=>"111001110",
  36391=>"101011110",
  36392=>"011001010",
  36393=>"101100101",
  36394=>"111011111",
  36395=>"111010101",
  36396=>"101000100",
  36397=>"010100100",
  36398=>"100011000",
  36399=>"101110000",
  36400=>"110110110",
  36401=>"000100110",
  36402=>"110010000",
  36403=>"010111101",
  36404=>"001100100",
  36405=>"111011010",
  36406=>"101101110",
  36407=>"110110011",
  36408=>"101101001",
  36409=>"100011101",
  36410=>"101110101",
  36411=>"010001111",
  36412=>"101000100",
  36413=>"001011101",
  36414=>"101010010",
  36415=>"010100110",
  36416=>"101111010",
  36417=>"001111000",
  36418=>"110011000",
  36419=>"011000100",
  36420=>"000100010",
  36421=>"101010011",
  36422=>"000001111",
  36423=>"010001011",
  36424=>"111010110",
  36425=>"100000000",
  36426=>"000001110",
  36427=>"001011000",
  36428=>"011001010",
  36429=>"000111010",
  36430=>"101001000",
  36431=>"011010000",
  36432=>"111011111",
  36433=>"011010111",
  36434=>"110011111",
  36435=>"011110110",
  36436=>"101111010",
  36437=>"010101010",
  36438=>"010111111",
  36439=>"111111000",
  36440=>"001010000",
  36441=>"110011010",
  36442=>"010100110",
  36443=>"001100111",
  36444=>"010100010",
  36445=>"110011110",
  36446=>"000000110",
  36447=>"100110101",
  36448=>"110101110",
  36449=>"110110010",
  36450=>"111010101",
  36451=>"110111110",
  36452=>"011111101",
  36453=>"000000001",
  36454=>"011011001",
  36455=>"000110001",
  36456=>"010110010",
  36457=>"101100001",
  36458=>"010111100",
  36459=>"111110111",
  36460=>"011101000",
  36461=>"010010101",
  36462=>"000000010",
  36463=>"011111100",
  36464=>"111110000",
  36465=>"000001000",
  36466=>"110111111",
  36467=>"000111011",
  36468=>"101111110",
  36469=>"001110010",
  36470=>"011100110",
  36471=>"010100000",
  36472=>"110111011",
  36473=>"010001001",
  36474=>"001011000",
  36475=>"000110010",
  36476=>"111000111",
  36477=>"010000110",
  36478=>"001010110",
  36479=>"101010101",
  36480=>"000000000",
  36481=>"000001011",
  36482=>"011011111",
  36483=>"000100000",
  36484=>"000110101",
  36485=>"101101000",
  36486=>"110010111",
  36487=>"110011111",
  36488=>"100000101",
  36489=>"111000001",
  36490=>"101100011",
  36491=>"001100110",
  36492=>"011011111",
  36493=>"000000111",
  36494=>"100101000",
  36495=>"011100001",
  36496=>"011011010",
  36497=>"110000100",
  36498=>"100100101",
  36499=>"010100101",
  36500=>"111110101",
  36501=>"000001010",
  36502=>"111011110",
  36503=>"101110011",
  36504=>"000100100",
  36505=>"000111101",
  36506=>"010100010",
  36507=>"100011100",
  36508=>"100011100",
  36509=>"110011000",
  36510=>"010100111",
  36511=>"000000010",
  36512=>"100010010",
  36513=>"101001010",
  36514=>"011010000",
  36515=>"010111010",
  36516=>"001101000",
  36517=>"001011111",
  36518=>"011101000",
  36519=>"100000100",
  36520=>"011110111",
  36521=>"011100011",
  36522=>"001100011",
  36523=>"100111101",
  36524=>"011111000",
  36525=>"011111111",
  36526=>"110110111",
  36527=>"111011010",
  36528=>"100000000",
  36529=>"100111111",
  36530=>"010000011",
  36531=>"111101111",
  36532=>"111001001",
  36533=>"001101010",
  36534=>"001011111",
  36535=>"101000111",
  36536=>"110000110",
  36537=>"111010110",
  36538=>"111000111",
  36539=>"000011001",
  36540=>"000111011",
  36541=>"011000011",
  36542=>"011110011",
  36543=>"110100101",
  36544=>"011111010",
  36545=>"011101100",
  36546=>"100100100",
  36547=>"011100010",
  36548=>"011000001",
  36549=>"111001111",
  36550=>"101101111",
  36551=>"000000111",
  36552=>"001011100",
  36553=>"110101001",
  36554=>"110010111",
  36555=>"110001001",
  36556=>"101011001",
  36557=>"000110000",
  36558=>"010011100",
  36559=>"111100101",
  36560=>"100110010",
  36561=>"011100111",
  36562=>"000111010",
  36563=>"010010000",
  36564=>"110011100",
  36565=>"000001010",
  36566=>"111001101",
  36567=>"110101100",
  36568=>"111100010",
  36569=>"000101000",
  36570=>"010000000",
  36571=>"011100111",
  36572=>"110001011",
  36573=>"001010110",
  36574=>"101010011",
  36575=>"010010100",
  36576=>"000011101",
  36577=>"000100000",
  36578=>"111101100",
  36579=>"101111101",
  36580=>"110000111",
  36581=>"111100010",
  36582=>"101010111",
  36583=>"011001010",
  36584=>"000000101",
  36585=>"000101100",
  36586=>"100001000",
  36587=>"001010000",
  36588=>"000011101",
  36589=>"010110111",
  36590=>"101011111",
  36591=>"100101000",
  36592=>"010011001",
  36593=>"101111011",
  36594=>"011111001",
  36595=>"100000001",
  36596=>"010100100",
  36597=>"001110000",
  36598=>"010100011",
  36599=>"000010011",
  36600=>"101110111",
  36601=>"011001010",
  36602=>"100100001",
  36603=>"000101100",
  36604=>"111111011",
  36605=>"101001011",
  36606=>"101100000",
  36607=>"101000110",
  36608=>"011111100",
  36609=>"011101110",
  36610=>"010101000",
  36611=>"101101100",
  36612=>"110101101",
  36613=>"010100110",
  36614=>"101100111",
  36615=>"011101001",
  36616=>"011101011",
  36617=>"111110100",
  36618=>"100001000",
  36619=>"110111111",
  36620=>"011000101",
  36621=>"110010001",
  36622=>"001000011",
  36623=>"010011100",
  36624=>"000110000",
  36625=>"000001011",
  36626=>"101000000",
  36627=>"000100100",
  36628=>"011001000",
  36629=>"110100011",
  36630=>"100111000",
  36631=>"101000110",
  36632=>"011110011",
  36633=>"011111111",
  36634=>"000100110",
  36635=>"000100011",
  36636=>"110011110",
  36637=>"001111010",
  36638=>"000111110",
  36639=>"101111110",
  36640=>"100000010",
  36641=>"001100001",
  36642=>"100100111",
  36643=>"011011000",
  36644=>"101111100",
  36645=>"101001000",
  36646=>"101111000",
  36647=>"010010001",
  36648=>"001110011",
  36649=>"001001100",
  36650=>"110000111",
  36651=>"110010001",
  36652=>"101010111",
  36653=>"111001101",
  36654=>"110001010",
  36655=>"001110011",
  36656=>"111010001",
  36657=>"110110001",
  36658=>"110000100",
  36659=>"010100001",
  36660=>"101001000",
  36661=>"101000101",
  36662=>"111111111",
  36663=>"101110111",
  36664=>"011110010",
  36665=>"101100101",
  36666=>"110010100",
  36667=>"111000010",
  36668=>"001010101",
  36669=>"010110111",
  36670=>"001101111",
  36671=>"011011001",
  36672=>"110110111",
  36673=>"111100001",
  36674=>"111110100",
  36675=>"110100010",
  36676=>"011011001",
  36677=>"010001100",
  36678=>"100010000",
  36679=>"110101000",
  36680=>"011101101",
  36681=>"111111010",
  36682=>"100111010",
  36683=>"010000000",
  36684=>"100110111",
  36685=>"011101100",
  36686=>"111111011",
  36687=>"100000111",
  36688=>"110101010",
  36689=>"110001100",
  36690=>"100111111",
  36691=>"100110110",
  36692=>"111101010",
  36693=>"001101011",
  36694=>"111111111",
  36695=>"110101100",
  36696=>"011110111",
  36697=>"010101001",
  36698=>"011010000",
  36699=>"010011011",
  36700=>"000101100",
  36701=>"111101000",
  36702=>"010111101",
  36703=>"000000101",
  36704=>"101111001",
  36705=>"100001011",
  36706=>"011001010",
  36707=>"111000001",
  36708=>"011010010",
  36709=>"110000000",
  36710=>"000001000",
  36711=>"010010001",
  36712=>"000100000",
  36713=>"001100101",
  36714=>"101001110",
  36715=>"110111011",
  36716=>"110111000",
  36717=>"100100000",
  36718=>"101000110",
  36719=>"001000000",
  36720=>"011110101",
  36721=>"000000010",
  36722=>"010100000",
  36723=>"111011000",
  36724=>"100011000",
  36725=>"100101101",
  36726=>"000001001",
  36727=>"101100111",
  36728=>"011101010",
  36729=>"111111110",
  36730=>"110111111",
  36731=>"000001101",
  36732=>"101001000",
  36733=>"000010101",
  36734=>"111101110",
  36735=>"000001000",
  36736=>"110100010",
  36737=>"011000111",
  36738=>"000001100",
  36739=>"101110101",
  36740=>"110011100",
  36741=>"011100000",
  36742=>"110110111",
  36743=>"000101011",
  36744=>"001001011",
  36745=>"000001110",
  36746=>"110110001",
  36747=>"111111111",
  36748=>"110111111",
  36749=>"001100011",
  36750=>"110011100",
  36751=>"110010100",
  36752=>"001110100",
  36753=>"110100010",
  36754=>"011111000",
  36755=>"100011010",
  36756=>"001100001",
  36757=>"101110101",
  36758=>"010111111",
  36759=>"000101001",
  36760=>"111100011",
  36761=>"001011001",
  36762=>"001111000",
  36763=>"110100100",
  36764=>"111111010",
  36765=>"011011111",
  36766=>"001111110",
  36767=>"000010000",
  36768=>"010111011",
  36769=>"011101111",
  36770=>"010010110",
  36771=>"111010100",
  36772=>"000001101",
  36773=>"101000011",
  36774=>"101101000",
  36775=>"000000011",
  36776=>"100110001",
  36777=>"111101011",
  36778=>"110010001",
  36779=>"101000001",
  36780=>"110001111",
  36781=>"001010110",
  36782=>"000001101",
  36783=>"110101101",
  36784=>"010000000",
  36785=>"100101011",
  36786=>"100101111",
  36787=>"011001101",
  36788=>"111001101",
  36789=>"011001001",
  36790=>"011100100",
  36791=>"010110000",
  36792=>"111100011",
  36793=>"111101100",
  36794=>"101011100",
  36795=>"101000111",
  36796=>"010010000",
  36797=>"101001110",
  36798=>"000101101",
  36799=>"001111010",
  36800=>"011101011",
  36801=>"100001111",
  36802=>"010011110",
  36803=>"001111000",
  36804=>"001001111",
  36805=>"010001101",
  36806=>"011101010",
  36807=>"100110010",
  36808=>"111101010",
  36809=>"101100000",
  36810=>"000000100",
  36811=>"111000000",
  36812=>"101110111",
  36813=>"011010101",
  36814=>"001000001",
  36815=>"101001001",
  36816=>"010111100",
  36817=>"101011001",
  36818=>"110101110",
  36819=>"101010100",
  36820=>"011001001",
  36821=>"101100100",
  36822=>"001001110",
  36823=>"111010100",
  36824=>"110111001",
  36825=>"010100011",
  36826=>"000101001",
  36827=>"010011100",
  36828=>"001111101",
  36829=>"000100010",
  36830=>"101011000",
  36831=>"011101111",
  36832=>"110101110",
  36833=>"010010101",
  36834=>"110000110",
  36835=>"000110000",
  36836=>"000100101",
  36837=>"000001011",
  36838=>"011011110",
  36839=>"101000001",
  36840=>"111011111",
  36841=>"101001111",
  36842=>"000101100",
  36843=>"010110000",
  36844=>"010100100",
  36845=>"100010000",
  36846=>"001000101",
  36847=>"000010101",
  36848=>"100111110",
  36849=>"001111000",
  36850=>"110011101",
  36851=>"111111111",
  36852=>"010111010",
  36853=>"101100010",
  36854=>"000100001",
  36855=>"011000000",
  36856=>"011101000",
  36857=>"100001100",
  36858=>"110011110",
  36859=>"000001000",
  36860=>"100100101",
  36861=>"111100111",
  36862=>"100100001",
  36863=>"001000001",
  36864=>"110101110",
  36865=>"111100001",
  36866=>"111110110",
  36867=>"011111101",
  36868=>"111110111",
  36869=>"001000001",
  36870=>"110110010",
  36871=>"100100100",
  36872=>"000100110",
  36873=>"111100010",
  36874=>"010010111",
  36875=>"010110101",
  36876=>"110111010",
  36877=>"111001010",
  36878=>"110101111",
  36879=>"101001011",
  36880=>"000010110",
  36881=>"110010100",
  36882=>"101000010",
  36883=>"010100001",
  36884=>"000110010",
  36885=>"110111101",
  36886=>"101000000",
  36887=>"001111010",
  36888=>"101111011",
  36889=>"101100000",
  36890=>"101001101",
  36891=>"000001011",
  36892=>"100011010",
  36893=>"101010101",
  36894=>"110111011",
  36895=>"100011101",
  36896=>"110011111",
  36897=>"101111100",
  36898=>"001010101",
  36899=>"000111010",
  36900=>"011111000",
  36901=>"001001011",
  36902=>"000000100",
  36903=>"110111011",
  36904=>"001100111",
  36905=>"101010001",
  36906=>"110100000",
  36907=>"111111101",
  36908=>"100011000",
  36909=>"000000001",
  36910=>"000001010",
  36911=>"110100101",
  36912=>"000111011",
  36913=>"110100101",
  36914=>"000001111",
  36915=>"101110111",
  36916=>"010010000",
  36917=>"111000100",
  36918=>"100011010",
  36919=>"101011100",
  36920=>"011001111",
  36921=>"000010100",
  36922=>"001000001",
  36923=>"101000011",
  36924=>"110111101",
  36925=>"001010111",
  36926=>"100100101",
  36927=>"100100011",
  36928=>"111110001",
  36929=>"100000111",
  36930=>"000001111",
  36931=>"101010100",
  36932=>"010110100",
  36933=>"010100001",
  36934=>"011001111",
  36935=>"000011011",
  36936=>"001101100",
  36937=>"110010001",
  36938=>"100101101",
  36939=>"000010011",
  36940=>"010001001",
  36941=>"111001000",
  36942=>"111101101",
  36943=>"000101001",
  36944=>"110011010",
  36945=>"010011100",
  36946=>"010011010",
  36947=>"011011010",
  36948=>"001001110",
  36949=>"101110110",
  36950=>"100100101",
  36951=>"001101010",
  36952=>"000110000",
  36953=>"100000011",
  36954=>"110000011",
  36955=>"100000000",
  36956=>"101000000",
  36957=>"110001111",
  36958=>"000011110",
  36959=>"100101101",
  36960=>"000101000",
  36961=>"101101010",
  36962=>"010000101",
  36963=>"011000010",
  36964=>"010010001",
  36965=>"111000000",
  36966=>"101100000",
  36967=>"110010000",
  36968=>"000100001",
  36969=>"010111001",
  36970=>"110110000",
  36971=>"110111110",
  36972=>"101000111",
  36973=>"100110011",
  36974=>"001010110",
  36975=>"101111010",
  36976=>"111001101",
  36977=>"100001010",
  36978=>"110000110",
  36979=>"111100001",
  36980=>"001010101",
  36981=>"001100000",
  36982=>"001101011",
  36983=>"100110110",
  36984=>"100111010",
  36985=>"111101111",
  36986=>"000011111",
  36987=>"000010111",
  36988=>"001010110",
  36989=>"010001110",
  36990=>"011111011",
  36991=>"011011101",
  36992=>"011101101",
  36993=>"110001110",
  36994=>"101110111",
  36995=>"011011001",
  36996=>"111000100",
  36997=>"100001100",
  36998=>"100110101",
  36999=>"010101110",
  37000=>"010000011",
  37001=>"000000000",
  37002=>"100110110",
  37003=>"010100001",
  37004=>"110101000",
  37005=>"010001101",
  37006=>"101010100",
  37007=>"111010110",
  37008=>"110101001",
  37009=>"001110001",
  37010=>"110111001",
  37011=>"000100100",
  37012=>"101001001",
  37013=>"011001011",
  37014=>"110100111",
  37015=>"011101110",
  37016=>"011000001",
  37017=>"000100110",
  37018=>"011111000",
  37019=>"101011111",
  37020=>"101100110",
  37021=>"100000000",
  37022=>"101110101",
  37023=>"010111101",
  37024=>"001001100",
  37025=>"011101101",
  37026=>"011010111",
  37027=>"000011100",
  37028=>"111010101",
  37029=>"001110110",
  37030=>"110111010",
  37031=>"010001101",
  37032=>"110010011",
  37033=>"111100110",
  37034=>"110111101",
  37035=>"111001010",
  37036=>"010001000",
  37037=>"110001011",
  37038=>"011001100",
  37039=>"001111001",
  37040=>"000100100",
  37041=>"100111011",
  37042=>"010001001",
  37043=>"101110000",
  37044=>"001100010",
  37045=>"101111011",
  37046=>"101000000",
  37047=>"001101110",
  37048=>"011010111",
  37049=>"010001010",
  37050=>"010100000",
  37051=>"000100000",
  37052=>"001111011",
  37053=>"000000000",
  37054=>"101000010",
  37055=>"010111010",
  37056=>"000100111",
  37057=>"001110111",
  37058=>"100110000",
  37059=>"111011010",
  37060=>"101001001",
  37061=>"011000000",
  37062=>"000000000",
  37063=>"111001110",
  37064=>"100111100",
  37065=>"110100011",
  37066=>"100001000",
  37067=>"100110011",
  37068=>"100011000",
  37069=>"110001111",
  37070=>"010100100",
  37071=>"111010011",
  37072=>"010110000",
  37073=>"110111100",
  37074=>"011111010",
  37075=>"001011100",
  37076=>"101010010",
  37077=>"001111100",
  37078=>"110110101",
  37079=>"011110010",
  37080=>"001011000",
  37081=>"100111101",
  37082=>"110101011",
  37083=>"101101011",
  37084=>"010110101",
  37085=>"111111101",
  37086=>"111001001",
  37087=>"001101110",
  37088=>"111110100",
  37089=>"001101000",
  37090=>"110110101",
  37091=>"000100001",
  37092=>"110111011",
  37093=>"000011101",
  37094=>"001110011",
  37095=>"111110110",
  37096=>"000101111",
  37097=>"100000011",
  37098=>"001110000",
  37099=>"101101010",
  37100=>"011100100",
  37101=>"011111011",
  37102=>"110100000",
  37103=>"010010110",
  37104=>"011110011",
  37105=>"011110101",
  37106=>"111001001",
  37107=>"000100000",
  37108=>"111111100",
  37109=>"001101101",
  37110=>"010111110",
  37111=>"000110101",
  37112=>"100111011",
  37113=>"001010000",
  37114=>"111111011",
  37115=>"011010011",
  37116=>"000101100",
  37117=>"011010000",
  37118=>"011100101",
  37119=>"010111010",
  37120=>"111001110",
  37121=>"011001111",
  37122=>"110111011",
  37123=>"000011010",
  37124=>"011111101",
  37125=>"011110110",
  37126=>"101001101",
  37127=>"011011000",
  37128=>"001001101",
  37129=>"001010000",
  37130=>"100001000",
  37131=>"101111010",
  37132=>"100010000",
  37133=>"011001110",
  37134=>"000101000",
  37135=>"010001011",
  37136=>"110011100",
  37137=>"010110000",
  37138=>"111001101",
  37139=>"111011010",
  37140=>"010001001",
  37141=>"100100000",
  37142=>"101110000",
  37143=>"000000010",
  37144=>"100111101",
  37145=>"110110000",
  37146=>"100000001",
  37147=>"101000101",
  37148=>"010000001",
  37149=>"110100111",
  37150=>"001001000",
  37151=>"010101000",
  37152=>"101011100",
  37153=>"000110100",
  37154=>"001000001",
  37155=>"001010100",
  37156=>"111000010",
  37157=>"110000000",
  37158=>"110001010",
  37159=>"000100000",
  37160=>"110000010",
  37161=>"010110111",
  37162=>"000101000",
  37163=>"010111011",
  37164=>"010000111",
  37165=>"011011100",
  37166=>"000010011",
  37167=>"010010110",
  37168=>"110110101",
  37169=>"010101010",
  37170=>"010011101",
  37171=>"001010010",
  37172=>"100111101",
  37173=>"001001001",
  37174=>"001001101",
  37175=>"111101011",
  37176=>"110101001",
  37177=>"001100110",
  37178=>"101100000",
  37179=>"101000000",
  37180=>"110010011",
  37181=>"110111000",
  37182=>"110001101",
  37183=>"100001011",
  37184=>"010100001",
  37185=>"111100000",
  37186=>"011000010",
  37187=>"110000000",
  37188=>"101001100",
  37189=>"001111110",
  37190=>"111001001",
  37191=>"001110110",
  37192=>"010111010",
  37193=>"101100100",
  37194=>"011001001",
  37195=>"010001101",
  37196=>"100101111",
  37197=>"110010010",
  37198=>"000100011",
  37199=>"011000110",
  37200=>"001000000",
  37201=>"010100011",
  37202=>"101000010",
  37203=>"000001011",
  37204=>"000010100",
  37205=>"100101000",
  37206=>"011001010",
  37207=>"000100011",
  37208=>"100100011",
  37209=>"110111000",
  37210=>"011110111",
  37211=>"010000001",
  37212=>"001111100",
  37213=>"111110100",
  37214=>"111110101",
  37215=>"001001001",
  37216=>"011000100",
  37217=>"011010101",
  37218=>"011100011",
  37219=>"011001110",
  37220=>"010011110",
  37221=>"111111110",
  37222=>"101111010",
  37223=>"010010000",
  37224=>"001111110",
  37225=>"001000001",
  37226=>"101010110",
  37227=>"001011001",
  37228=>"110011011",
  37229=>"011111000",
  37230=>"111000101",
  37231=>"011101010",
  37232=>"110100110",
  37233=>"011011011",
  37234=>"110001000",
  37235=>"101101111",
  37236=>"010100110",
  37237=>"010011011",
  37238=>"111010100",
  37239=>"010011111",
  37240=>"001111110",
  37241=>"011011111",
  37242=>"110001000",
  37243=>"001000110",
  37244=>"001011011",
  37245=>"110101101",
  37246=>"010110011",
  37247=>"100111110",
  37248=>"111010001",
  37249=>"000001010",
  37250=>"100011110",
  37251=>"010101101",
  37252=>"010100001",
  37253=>"111010011",
  37254=>"111000001",
  37255=>"000101000",
  37256=>"000000101",
  37257=>"111111111",
  37258=>"110100111",
  37259=>"100101111",
  37260=>"000001110",
  37261=>"010001011",
  37262=>"101001010",
  37263=>"010110111",
  37264=>"111000011",
  37265=>"010000100",
  37266=>"111011101",
  37267=>"001100100",
  37268=>"111111011",
  37269=>"001000010",
  37270=>"001100000",
  37271=>"001000001",
  37272=>"010111000",
  37273=>"100001100",
  37274=>"000111001",
  37275=>"101100001",
  37276=>"011100101",
  37277=>"001001111",
  37278=>"001010101",
  37279=>"111111100",
  37280=>"111101000",
  37281=>"011000101",
  37282=>"000111011",
  37283=>"001001011",
  37284=>"001001001",
  37285=>"000010100",
  37286=>"101001010",
  37287=>"000100111",
  37288=>"100111000",
  37289=>"101111000",
  37290=>"010111110",
  37291=>"011000000",
  37292=>"000010110",
  37293=>"100110001",
  37294=>"111111100",
  37295=>"110011011",
  37296=>"100100010",
  37297=>"000010101",
  37298=>"101101100",
  37299=>"110000001",
  37300=>"111111010",
  37301=>"010000011",
  37302=>"100101110",
  37303=>"011100000",
  37304=>"000101101",
  37305=>"000111111",
  37306=>"001110011",
  37307=>"101101110",
  37308=>"101101001",
  37309=>"100111111",
  37310=>"100010010",
  37311=>"010001100",
  37312=>"101101000",
  37313=>"110000010",
  37314=>"100011010",
  37315=>"110011101",
  37316=>"011100110",
  37317=>"101001000",
  37318=>"010100100",
  37319=>"011101110",
  37320=>"111000100",
  37321=>"000111010",
  37322=>"001110111",
  37323=>"101100101",
  37324=>"011000100",
  37325=>"101010100",
  37326=>"000111011",
  37327=>"111011000",
  37328=>"100110100",
  37329=>"010000100",
  37330=>"001101101",
  37331=>"001110110",
  37332=>"010010000",
  37333=>"110101101",
  37334=>"010100110",
  37335=>"111010010",
  37336=>"001010111",
  37337=>"101011011",
  37338=>"101100100",
  37339=>"010011100",
  37340=>"100010110",
  37341=>"101100000",
  37342=>"111010000",
  37343=>"100011010",
  37344=>"100001111",
  37345=>"101000000",
  37346=>"111111010",
  37347=>"101000001",
  37348=>"110111001",
  37349=>"100111000",
  37350=>"101000000",
  37351=>"110010100",
  37352=>"010011000",
  37353=>"001000000",
  37354=>"001110100",
  37355=>"010000101",
  37356=>"011010000",
  37357=>"011111001",
  37358=>"100100010",
  37359=>"001100110",
  37360=>"111010110",
  37361=>"011001000",
  37362=>"111111110",
  37363=>"011111001",
  37364=>"100100011",
  37365=>"000111011",
  37366=>"100101100",
  37367=>"011001010",
  37368=>"000111110",
  37369=>"100110011",
  37370=>"010101001",
  37371=>"001101000",
  37372=>"101010010",
  37373=>"110101111",
  37374=>"011100001",
  37375=>"001010111",
  37376=>"000100110",
  37377=>"001111100",
  37378=>"110010000",
  37379=>"000000010",
  37380=>"110110111",
  37381=>"110101110",
  37382=>"001000101",
  37383=>"011000101",
  37384=>"010100000",
  37385=>"110000100",
  37386=>"001101010",
  37387=>"000100111",
  37388=>"001101001",
  37389=>"100101011",
  37390=>"011001000",
  37391=>"111010110",
  37392=>"110011111",
  37393=>"000100000",
  37394=>"011001011",
  37395=>"011001100",
  37396=>"011110011",
  37397=>"111000101",
  37398=>"110011111",
  37399=>"000110000",
  37400=>"111101101",
  37401=>"000011011",
  37402=>"010101010",
  37403=>"011010011",
  37404=>"011011010",
  37405=>"000101010",
  37406=>"011101011",
  37407=>"110111010",
  37408=>"000100100",
  37409=>"110010110",
  37410=>"001110011",
  37411=>"111001010",
  37412=>"110011010",
  37413=>"110001111",
  37414=>"010011110",
  37415=>"000010111",
  37416=>"101000101",
  37417=>"011011000",
  37418=>"011000011",
  37419=>"011010000",
  37420=>"110000100",
  37421=>"010011000",
  37422=>"000011010",
  37423=>"011001111",
  37424=>"100001111",
  37425=>"101110101",
  37426=>"101011110",
  37427=>"011000011",
  37428=>"001011011",
  37429=>"001000101",
  37430=>"101100110",
  37431=>"100010000",
  37432=>"101000000",
  37433=>"101101100",
  37434=>"010110100",
  37435=>"100000111",
  37436=>"000101001",
  37437=>"011011001",
  37438=>"000110111",
  37439=>"011100110",
  37440=>"010010100",
  37441=>"101101111",
  37442=>"011011001",
  37443=>"000100000",
  37444=>"100100110",
  37445=>"011001110",
  37446=>"001110011",
  37447=>"110111001",
  37448=>"001000011",
  37449=>"100011110",
  37450=>"010000101",
  37451=>"110110001",
  37452=>"110011010",
  37453=>"111010001",
  37454=>"000001010",
  37455=>"010000011",
  37456=>"110101111",
  37457=>"001100100",
  37458=>"010100001",
  37459=>"110010100",
  37460=>"100100101",
  37461=>"100010000",
  37462=>"111111100",
  37463=>"111011010",
  37464=>"100010100",
  37465=>"110000110",
  37466=>"000101111",
  37467=>"101111101",
  37468=>"011010101",
  37469=>"000010010",
  37470=>"010000110",
  37471=>"010110111",
  37472=>"010011101",
  37473=>"100011011",
  37474=>"101100101",
  37475=>"001100010",
  37476=>"100000101",
  37477=>"110101000",
  37478=>"100000011",
  37479=>"000110111",
  37480=>"011001100",
  37481=>"010100111",
  37482=>"000110000",
  37483=>"100011010",
  37484=>"100010010",
  37485=>"111110010",
  37486=>"001011010",
  37487=>"010110010",
  37488=>"011101000",
  37489=>"000010101",
  37490=>"111000010",
  37491=>"101101110",
  37492=>"000001011",
  37493=>"110111010",
  37494=>"001011010",
  37495=>"010000100",
  37496=>"111001000",
  37497=>"010011011",
  37498=>"100001001",
  37499=>"100110101",
  37500=>"111010000",
  37501=>"101001100",
  37502=>"110111101",
  37503=>"000001001",
  37504=>"101100100",
  37505=>"011010110",
  37506=>"111100000",
  37507=>"011101111",
  37508=>"100110100",
  37509=>"001010100",
  37510=>"011000100",
  37511=>"110111010",
  37512=>"010001001",
  37513=>"100000111",
  37514=>"100011000",
  37515=>"101101011",
  37516=>"010100000",
  37517=>"000100101",
  37518=>"110011011",
  37519=>"100001000",
  37520=>"101010001",
  37521=>"101111000",
  37522=>"101101110",
  37523=>"000011000",
  37524=>"000000010",
  37525=>"101010110",
  37526=>"101001111",
  37527=>"001110011",
  37528=>"111001011",
  37529=>"001010000",
  37530=>"000110100",
  37531=>"011001110",
  37532=>"101101011",
  37533=>"000101010",
  37534=>"111111011",
  37535=>"111111000",
  37536=>"011001000",
  37537=>"001011000",
  37538=>"010000101",
  37539=>"110100110",
  37540=>"000001011",
  37541=>"110001100",
  37542=>"001001111",
  37543=>"000010111",
  37544=>"110011000",
  37545=>"010101011",
  37546=>"111110001",
  37547=>"000100000",
  37548=>"100100000",
  37549=>"010001001",
  37550=>"001000100",
  37551=>"011111110",
  37552=>"000001110",
  37553=>"110111101",
  37554=>"110111000",
  37555=>"001000111",
  37556=>"110001001",
  37557=>"111101010",
  37558=>"011111001",
  37559=>"111111110",
  37560=>"100101000",
  37561=>"000011100",
  37562=>"010000000",
  37563=>"111010010",
  37564=>"101100101",
  37565=>"000011110",
  37566=>"000000000",
  37567=>"111101110",
  37568=>"111100111",
  37569=>"001011001",
  37570=>"000111011",
  37571=>"001110000",
  37572=>"001010110",
  37573=>"100101110",
  37574=>"001011101",
  37575=>"100010011",
  37576=>"111000010",
  37577=>"100000101",
  37578=>"001100000",
  37579=>"001001001",
  37580=>"000101100",
  37581=>"101111111",
  37582=>"000010001",
  37583=>"101010001",
  37584=>"111011110",
  37585=>"100100111",
  37586=>"010100011",
  37587=>"110110110",
  37588=>"001101010",
  37589=>"001000011",
  37590=>"101101110",
  37591=>"010001101",
  37592=>"101111111",
  37593=>"101010100",
  37594=>"000101101",
  37595=>"101110011",
  37596=>"110110101",
  37597=>"110000100",
  37598=>"001111110",
  37599=>"111011010",
  37600=>"100000110",
  37601=>"011001111",
  37602=>"010111001",
  37603=>"100001011",
  37604=>"000010101",
  37605=>"111000000",
  37606=>"000100000",
  37607=>"000000001",
  37608=>"100010010",
  37609=>"100101101",
  37610=>"100011001",
  37611=>"100110111",
  37612=>"101001110",
  37613=>"010000101",
  37614=>"000010100",
  37615=>"000111111",
  37616=>"111100111",
  37617=>"001100010",
  37618=>"011111000",
  37619=>"100010000",
  37620=>"101101100",
  37621=>"100111110",
  37622=>"011101011",
  37623=>"110100101",
  37624=>"011110111",
  37625=>"101110011",
  37626=>"101010011",
  37627=>"100010000",
  37628=>"101110001",
  37629=>"010101001",
  37630=>"111100001",
  37631=>"000001010",
  37632=>"011011101",
  37633=>"010011100",
  37634=>"010111001",
  37635=>"001101000",
  37636=>"110100101",
  37637=>"000001101",
  37638=>"011100010",
  37639=>"001000111",
  37640=>"100111000",
  37641=>"001001101",
  37642=>"110011101",
  37643=>"010011100",
  37644=>"111001100",
  37645=>"001010001",
  37646=>"101001110",
  37647=>"001101101",
  37648=>"001111001",
  37649=>"001001000",
  37650=>"000000001",
  37651=>"101111001",
  37652=>"000110100",
  37653=>"111011000",
  37654=>"101000010",
  37655=>"001100100",
  37656=>"000100001",
  37657=>"001100100",
  37658=>"100001001",
  37659=>"001101011",
  37660=>"000001101",
  37661=>"001010101",
  37662=>"001011000",
  37663=>"010011000",
  37664=>"001101111",
  37665=>"001100100",
  37666=>"111000010",
  37667=>"100000101",
  37668=>"011000001",
  37669=>"110110010",
  37670=>"100100100",
  37671=>"010100111",
  37672=>"101011011",
  37673=>"111001001",
  37674=>"010100111",
  37675=>"100011101",
  37676=>"010010111",
  37677=>"010010001",
  37678=>"100010110",
  37679=>"001011100",
  37680=>"101010100",
  37681=>"011101111",
  37682=>"000001001",
  37683=>"111100010",
  37684=>"011011011",
  37685=>"001110000",
  37686=>"001010011",
  37687=>"000000111",
  37688=>"010111100",
  37689=>"010100000",
  37690=>"101101001",
  37691=>"111010111",
  37692=>"100010000",
  37693=>"110001101",
  37694=>"101001100",
  37695=>"100100100",
  37696=>"011010111",
  37697=>"111100110",
  37698=>"000000101",
  37699=>"001100100",
  37700=>"001110001",
  37701=>"110011000",
  37702=>"110000010",
  37703=>"111111011",
  37704=>"111010111",
  37705=>"010000010",
  37706=>"000101001",
  37707=>"000110001",
  37708=>"111100101",
  37709=>"111010000",
  37710=>"111001101",
  37711=>"111101000",
  37712=>"111110001",
  37713=>"010100001",
  37714=>"001000000",
  37715=>"100100010",
  37716=>"101100010",
  37717=>"100111010",
  37718=>"010011011",
  37719=>"111101000",
  37720=>"000000110",
  37721=>"000100100",
  37722=>"111010111",
  37723=>"101101111",
  37724=>"001011010",
  37725=>"100110100",
  37726=>"000110101",
  37727=>"000001111",
  37728=>"101110010",
  37729=>"101101010",
  37730=>"011100000",
  37731=>"000100110",
  37732=>"101010110",
  37733=>"010101001",
  37734=>"100000001",
  37735=>"110111111",
  37736=>"110011111",
  37737=>"011010111",
  37738=>"111001100",
  37739=>"000001001",
  37740=>"110101000",
  37741=>"011110001",
  37742=>"000110000",
  37743=>"111110100",
  37744=>"101110110",
  37745=>"011011011",
  37746=>"001000101",
  37747=>"010111101",
  37748=>"000001101",
  37749=>"110000101",
  37750=>"011001010",
  37751=>"101001010",
  37752=>"010001011",
  37753=>"111011010",
  37754=>"110001000",
  37755=>"111111011",
  37756=>"000110101",
  37757=>"101100111",
  37758=>"010011001",
  37759=>"111110010",
  37760=>"010001101",
  37761=>"010100111",
  37762=>"010010101",
  37763=>"101010001",
  37764=>"111110111",
  37765=>"000101000",
  37766=>"000001101",
  37767=>"101000110",
  37768=>"010110010",
  37769=>"111000100",
  37770=>"111011000",
  37771=>"100111101",
  37772=>"011011011",
  37773=>"001011101",
  37774=>"110000010",
  37775=>"011000001",
  37776=>"110011001",
  37777=>"000001001",
  37778=>"110100001",
  37779=>"100000101",
  37780=>"110000000",
  37781=>"111111101",
  37782=>"010011111",
  37783=>"110100110",
  37784=>"101000011",
  37785=>"100010101",
  37786=>"011111001",
  37787=>"000101001",
  37788=>"110100100",
  37789=>"001101000",
  37790=>"101110000",
  37791=>"111000000",
  37792=>"001001010",
  37793=>"100101000",
  37794=>"000100001",
  37795=>"110010100",
  37796=>"110011000",
  37797=>"110101001",
  37798=>"111001001",
  37799=>"000101001",
  37800=>"111110000",
  37801=>"000000011",
  37802=>"100110111",
  37803=>"110101001",
  37804=>"100001000",
  37805=>"100000011",
  37806=>"010011000",
  37807=>"000101110",
  37808=>"111001000",
  37809=>"000010101",
  37810=>"101110000",
  37811=>"000011110",
  37812=>"110001011",
  37813=>"010000110",
  37814=>"000111100",
  37815=>"000010110",
  37816=>"100011011",
  37817=>"101010001",
  37818=>"110010001",
  37819=>"011100101",
  37820=>"100101000",
  37821=>"110011011",
  37822=>"110101111",
  37823=>"010010100",
  37824=>"010101011",
  37825=>"110100111",
  37826=>"100010101",
  37827=>"110001010",
  37828=>"011011000",
  37829=>"000100000",
  37830=>"000000100",
  37831=>"111101000",
  37832=>"001000110",
  37833=>"111101011",
  37834=>"010000010",
  37835=>"001111101",
  37836=>"111000101",
  37837=>"000010000",
  37838=>"110011000",
  37839=>"011010110",
  37840=>"011100001",
  37841=>"010111111",
  37842=>"101001111",
  37843=>"100000100",
  37844=>"000101010",
  37845=>"110000001",
  37846=>"100010101",
  37847=>"111011110",
  37848=>"010011100",
  37849=>"101101110",
  37850=>"011111000",
  37851=>"110010100",
  37852=>"010011010",
  37853=>"100000100",
  37854=>"000101011",
  37855=>"100101001",
  37856=>"100011000",
  37857=>"000011110",
  37858=>"011101110",
  37859=>"100101001",
  37860=>"010100101",
  37861=>"100110100",
  37862=>"000100000",
  37863=>"001110100",
  37864=>"000101011",
  37865=>"000010111",
  37866=>"001100000",
  37867=>"010010010",
  37868=>"100101110",
  37869=>"110010111",
  37870=>"011001111",
  37871=>"110000001",
  37872=>"101010010",
  37873=>"100111011",
  37874=>"100001100",
  37875=>"010100111",
  37876=>"101000111",
  37877=>"010011010",
  37878=>"011110001",
  37879=>"101010100",
  37880=>"011101000",
  37881=>"010101010",
  37882=>"111101101",
  37883=>"110110100",
  37884=>"000111101",
  37885=>"011110110",
  37886=>"001010011",
  37887=>"110110011",
  37888=>"010010010",
  37889=>"001011001",
  37890=>"110101011",
  37891=>"010111011",
  37892=>"010010001",
  37893=>"111100111",
  37894=>"110010110",
  37895=>"100111000",
  37896=>"001010100",
  37897=>"010110101",
  37898=>"001011011",
  37899=>"111010011",
  37900=>"010000110",
  37901=>"111111011",
  37902=>"101000111",
  37903=>"010110000",
  37904=>"111011001",
  37905=>"010100001",
  37906=>"101010001",
  37907=>"010111011",
  37908=>"010110010",
  37909=>"101000101",
  37910=>"101110011",
  37911=>"101100110",
  37912=>"110011001",
  37913=>"011110111",
  37914=>"111101010",
  37915=>"100000111",
  37916=>"011111100",
  37917=>"110011000",
  37918=>"011010100",
  37919=>"110001000",
  37920=>"111010010",
  37921=>"100100110",
  37922=>"001101111",
  37923=>"011001100",
  37924=>"000000101",
  37925=>"010101111",
  37926=>"100001010",
  37927=>"011000110",
  37928=>"111111101",
  37929=>"000000011",
  37930=>"001011011",
  37931=>"000000111",
  37932=>"011110001",
  37933=>"001011000",
  37934=>"100101010",
  37935=>"010001001",
  37936=>"101010101",
  37937=>"101100011",
  37938=>"000010011",
  37939=>"010111111",
  37940=>"100010000",
  37941=>"000001000",
  37942=>"110000111",
  37943=>"110000110",
  37944=>"100110010",
  37945=>"101001101",
  37946=>"100000011",
  37947=>"110101110",
  37948=>"010010101",
  37949=>"110011111",
  37950=>"111010000",
  37951=>"110000011",
  37952=>"110101100",
  37953=>"001001110",
  37954=>"111010000",
  37955=>"010001010",
  37956=>"110000001",
  37957=>"110010110",
  37958=>"010001100",
  37959=>"000101100",
  37960=>"100100011",
  37961=>"111110000",
  37962=>"111001011",
  37963=>"000000001",
  37964=>"101111101",
  37965=>"100001111",
  37966=>"100001011",
  37967=>"100100011",
  37968=>"100000111",
  37969=>"111101011",
  37970=>"101101111",
  37971=>"101100111",
  37972=>"001000111",
  37973=>"111111000",
  37974=>"100100111",
  37975=>"100011100",
  37976=>"001011110",
  37977=>"111111101",
  37978=>"011110000",
  37979=>"100101100",
  37980=>"000111011",
  37981=>"101001001",
  37982=>"001001110",
  37983=>"011111111",
  37984=>"110000111",
  37985=>"101000010",
  37986=>"000001111",
  37987=>"100001101",
  37988=>"101001010",
  37989=>"111111111",
  37990=>"111010010",
  37991=>"010101101",
  37992=>"110101010",
  37993=>"010000111",
  37994=>"111010110",
  37995=>"011100101",
  37996=>"110001000",
  37997=>"110010010",
  37998=>"001001101",
  37999=>"000010110",
  38000=>"101100000",
  38001=>"001001010",
  38002=>"111111011",
  38003=>"100101010",
  38004=>"010101110",
  38005=>"100110110",
  38006=>"011101001",
  38007=>"011001001",
  38008=>"011101101",
  38009=>"111001101",
  38010=>"111110001",
  38011=>"101100111",
  38012=>"011011111",
  38013=>"000101110",
  38014=>"001000100",
  38015=>"010010001",
  38016=>"111010011",
  38017=>"111001101",
  38018=>"101000100",
  38019=>"100100100",
  38020=>"010101100",
  38021=>"000000001",
  38022=>"000110010",
  38023=>"000000111",
  38024=>"010011110",
  38025=>"011001101",
  38026=>"101000010",
  38027=>"000000101",
  38028=>"101111111",
  38029=>"011000000",
  38030=>"100110011",
  38031=>"110000001",
  38032=>"111100111",
  38033=>"111001000",
  38034=>"100111100",
  38035=>"100100010",
  38036=>"110100111",
  38037=>"100110000",
  38038=>"110011001",
  38039=>"010100100",
  38040=>"000000111",
  38041=>"010111011",
  38042=>"100010011",
  38043=>"011110000",
  38044=>"100010000",
  38045=>"100000110",
  38046=>"011111100",
  38047=>"011001111",
  38048=>"001010010",
  38049=>"110100100",
  38050=>"000101010",
  38051=>"001000001",
  38052=>"110000000",
  38053=>"000101001",
  38054=>"100101100",
  38055=>"111000000",
  38056=>"011010001",
  38057=>"111000101",
  38058=>"011000110",
  38059=>"011001010",
  38060=>"110111010",
  38061=>"110110101",
  38062=>"100000010",
  38063=>"000110101",
  38064=>"100100110",
  38065=>"000011100",
  38066=>"001011100",
  38067=>"100100100",
  38068=>"000001111",
  38069=>"000000011",
  38070=>"110111010",
  38071=>"010111100",
  38072=>"010111100",
  38073=>"101101111",
  38074=>"111001011",
  38075=>"011000100",
  38076=>"011000111",
  38077=>"110110110",
  38078=>"000001101",
  38079=>"001101101",
  38080=>"111011110",
  38081=>"100010011",
  38082=>"110100101",
  38083=>"011001110",
  38084=>"101000101",
  38085=>"100000111",
  38086=>"111110111",
  38087=>"010000011",
  38088=>"001100111",
  38089=>"010110101",
  38090=>"111110101",
  38091=>"101001101",
  38092=>"001000111",
  38093=>"011111100",
  38094=>"100100000",
  38095=>"110110100",
  38096=>"100100101",
  38097=>"001000011",
  38098=>"100111111",
  38099=>"011110110",
  38100=>"100001011",
  38101=>"001110000",
  38102=>"001111111",
  38103=>"100010001",
  38104=>"000010100",
  38105=>"111111101",
  38106=>"110111010",
  38107=>"111001101",
  38108=>"001111110",
  38109=>"101111110",
  38110=>"011101001",
  38111=>"000000000",
  38112=>"111110101",
  38113=>"011000011",
  38114=>"101011010",
  38115=>"111110110",
  38116=>"100001111",
  38117=>"011110111",
  38118=>"111101010",
  38119=>"111111100",
  38120=>"011011100",
  38121=>"111101011",
  38122=>"011000100",
  38123=>"010000000",
  38124=>"110110000",
  38125=>"110110111",
  38126=>"111100011",
  38127=>"101101011",
  38128=>"001011111",
  38129=>"101000000",
  38130=>"000000000",
  38131=>"100010001",
  38132=>"101001111",
  38133=>"011010001",
  38134=>"110110110",
  38135=>"100111000",
  38136=>"001001110",
  38137=>"010010001",
  38138=>"101101101",
  38139=>"010010011",
  38140=>"110010111",
  38141=>"100100101",
  38142=>"111110100",
  38143=>"101000100",
  38144=>"001101101",
  38145=>"001011000",
  38146=>"101100110",
  38147=>"011111010",
  38148=>"100000000",
  38149=>"100011111",
  38150=>"100010100",
  38151=>"101100010",
  38152=>"000001101",
  38153=>"100111011",
  38154=>"010011001",
  38155=>"111111100",
  38156=>"001011000",
  38157=>"100011101",
  38158=>"101011000",
  38159=>"111001101",
  38160=>"011100111",
  38161=>"101010001",
  38162=>"110111001",
  38163=>"000101110",
  38164=>"011000101",
  38165=>"010100101",
  38166=>"100110110",
  38167=>"110010010",
  38168=>"011010011",
  38169=>"111000100",
  38170=>"000110011",
  38171=>"011101001",
  38172=>"110111000",
  38173=>"100100010",
  38174=>"000000000",
  38175=>"010101101",
  38176=>"100111011",
  38177=>"100101010",
  38178=>"000101011",
  38179=>"010101100",
  38180=>"001001110",
  38181=>"001001100",
  38182=>"101111001",
  38183=>"110011101",
  38184=>"001111100",
  38185=>"100111010",
  38186=>"111110100",
  38187=>"100011101",
  38188=>"110110000",
  38189=>"001001010",
  38190=>"011011011",
  38191=>"011111101",
  38192=>"011110000",
  38193=>"000100111",
  38194=>"101000001",
  38195=>"000100011",
  38196=>"001110001",
  38197=>"000000111",
  38198=>"011001110",
  38199=>"101111111",
  38200=>"000010010",
  38201=>"011111000",
  38202=>"111100110",
  38203=>"001010110",
  38204=>"001000100",
  38205=>"010000010",
  38206=>"110010100",
  38207=>"111100110",
  38208=>"111000111",
  38209=>"101011011",
  38210=>"111111101",
  38211=>"110011100",
  38212=>"011010111",
  38213=>"111001001",
  38214=>"111000000",
  38215=>"100100001",
  38216=>"101011100",
  38217=>"100101100",
  38218=>"001010100",
  38219=>"100100001",
  38220=>"000010001",
  38221=>"000010011",
  38222=>"011100100",
  38223=>"101101111",
  38224=>"011110101",
  38225=>"101100010",
  38226=>"000101100",
  38227=>"001001010",
  38228=>"111011111",
  38229=>"001101010",
  38230=>"110011001",
  38231=>"101010101",
  38232=>"001101011",
  38233=>"111110010",
  38234=>"101111101",
  38235=>"111111011",
  38236=>"011010011",
  38237=>"000000000",
  38238=>"111010010",
  38239=>"111100001",
  38240=>"000111101",
  38241=>"001101110",
  38242=>"100110000",
  38243=>"000010001",
  38244=>"100000001",
  38245=>"111011001",
  38246=>"110101110",
  38247=>"010000000",
  38248=>"110101011",
  38249=>"000100011",
  38250=>"111000000",
  38251=>"000001010",
  38252=>"001100100",
  38253=>"000100010",
  38254=>"110000000",
  38255=>"011001010",
  38256=>"011110010",
  38257=>"001011010",
  38258=>"001001111",
  38259=>"111001101",
  38260=>"101001010",
  38261=>"100100011",
  38262=>"000000101",
  38263=>"101000100",
  38264=>"000000111",
  38265=>"000101010",
  38266=>"100001001",
  38267=>"000001111",
  38268=>"001000101",
  38269=>"000101001",
  38270=>"101101010",
  38271=>"011000111",
  38272=>"101111111",
  38273=>"000100101",
  38274=>"101100101",
  38275=>"000100111",
  38276=>"000101100",
  38277=>"010001100",
  38278=>"101001100",
  38279=>"101111111",
  38280=>"001111010",
  38281=>"010001010",
  38282=>"001001110",
  38283=>"000000000",
  38284=>"011010101",
  38285=>"101001101",
  38286=>"001110011",
  38287=>"000001111",
  38288=>"001111000",
  38289=>"000011110",
  38290=>"010111100",
  38291=>"001000100",
  38292=>"111000100",
  38293=>"101100110",
  38294=>"011001000",
  38295=>"001101001",
  38296=>"010000100",
  38297=>"011010011",
  38298=>"100011111",
  38299=>"010000011",
  38300=>"001011000",
  38301=>"110100011",
  38302=>"100111111",
  38303=>"001000000",
  38304=>"110011100",
  38305=>"011100001",
  38306=>"001000110",
  38307=>"000001000",
  38308=>"001000011",
  38309=>"010010000",
  38310=>"000110100",
  38311=>"100001111",
  38312=>"011101100",
  38313=>"011000011",
  38314=>"000000001",
  38315=>"000000101",
  38316=>"101100111",
  38317=>"111110111",
  38318=>"000000111",
  38319=>"000100101",
  38320=>"010111001",
  38321=>"001111110",
  38322=>"000010000",
  38323=>"110110011",
  38324=>"010100000",
  38325=>"011000101",
  38326=>"100010100",
  38327=>"101101111",
  38328=>"111101001",
  38329=>"100110100",
  38330=>"011001000",
  38331=>"101001111",
  38332=>"101011001",
  38333=>"101001110",
  38334=>"100001001",
  38335=>"111011100",
  38336=>"101100000",
  38337=>"101101111",
  38338=>"001000100",
  38339=>"101111011",
  38340=>"101010100",
  38341=>"000111011",
  38342=>"111001011",
  38343=>"011100100",
  38344=>"100001100",
  38345=>"010100100",
  38346=>"110111001",
  38347=>"110110001",
  38348=>"111001011",
  38349=>"110111100",
  38350=>"000010110",
  38351=>"011111111",
  38352=>"101010111",
  38353=>"011000110",
  38354=>"011110001",
  38355=>"001110000",
  38356=>"111110100",
  38357=>"111100111",
  38358=>"100100000",
  38359=>"111110000",
  38360=>"000100010",
  38361=>"100000001",
  38362=>"101111010",
  38363=>"111101111",
  38364=>"101010010",
  38365=>"101010011",
  38366=>"000110000",
  38367=>"000001011",
  38368=>"010110110",
  38369=>"100111000",
  38370=>"111100001",
  38371=>"010101110",
  38372=>"011011110",
  38373=>"111000000",
  38374=>"011111101",
  38375=>"111000101",
  38376=>"010000110",
  38377=>"110011010",
  38378=>"101001011",
  38379=>"001101110",
  38380=>"100001010",
  38381=>"010110100",
  38382=>"001010101",
  38383=>"111010010",
  38384=>"100001101",
  38385=>"101001001",
  38386=>"001100100",
  38387=>"101001010",
  38388=>"001101001",
  38389=>"010110111",
  38390=>"101000101",
  38391=>"101110011",
  38392=>"010001001",
  38393=>"000101001",
  38394=>"100101111",
  38395=>"010010010",
  38396=>"001001111",
  38397=>"001110110",
  38398=>"110001010",
  38399=>"010110001",
  38400=>"011111101",
  38401=>"101011101",
  38402=>"000111111",
  38403=>"011111010",
  38404=>"001001111",
  38405=>"001000000",
  38406=>"010001101",
  38407=>"110110011",
  38408=>"000110000",
  38409=>"010010110",
  38410=>"010001011",
  38411=>"110011011",
  38412=>"111110000",
  38413=>"001000100",
  38414=>"100000110",
  38415=>"011011010",
  38416=>"111110101",
  38417=>"001000111",
  38418=>"100100110",
  38419=>"011100000",
  38420=>"011110100",
  38421=>"101000101",
  38422=>"010000111",
  38423=>"001011110",
  38424=>"001100000",
  38425=>"000100000",
  38426=>"010000000",
  38427=>"100000010",
  38428=>"001111010",
  38429=>"000100110",
  38430=>"001100010",
  38431=>"110001011",
  38432=>"001001111",
  38433=>"110001101",
  38434=>"100010110",
  38435=>"010000101",
  38436=>"011011110",
  38437=>"010110001",
  38438=>"111101001",
  38439=>"101001000",
  38440=>"010101101",
  38441=>"001110011",
  38442=>"001110100",
  38443=>"001011101",
  38444=>"101000100",
  38445=>"000100100",
  38446=>"010100111",
  38447=>"000011001",
  38448=>"111011010",
  38449=>"100111111",
  38450=>"001001001",
  38451=>"101111101",
  38452=>"011011000",
  38453=>"110001101",
  38454=>"110000000",
  38455=>"000100010",
  38456=>"101011010",
  38457=>"110100110",
  38458=>"001000000",
  38459=>"010110011",
  38460=>"111000110",
  38461=>"110010100",
  38462=>"001000001",
  38463=>"101111011",
  38464=>"011010111",
  38465=>"011100011",
  38466=>"101000011",
  38467=>"010010101",
  38468=>"111001000",
  38469=>"111000111",
  38470=>"110010011",
  38471=>"110000000",
  38472=>"000010010",
  38473=>"111111011",
  38474=>"011000110",
  38475=>"101001111",
  38476=>"111101111",
  38477=>"100001110",
  38478=>"001011010",
  38479=>"000110010",
  38480=>"110010101",
  38481=>"000000000",
  38482=>"110110110",
  38483=>"000110100",
  38484=>"010100000",
  38485=>"011111110",
  38486=>"000110100",
  38487=>"001001011",
  38488=>"110110101",
  38489=>"010000011",
  38490=>"000110010",
  38491=>"100000100",
  38492=>"101011011",
  38493=>"101011001",
  38494=>"100010101",
  38495=>"111011101",
  38496=>"111011100",
  38497=>"000010100",
  38498=>"010000110",
  38499=>"100000001",
  38500=>"010001110",
  38501=>"000001101",
  38502=>"011000110",
  38503=>"101100111",
  38504=>"000110001",
  38505=>"101101110",
  38506=>"110100001",
  38507=>"111000101",
  38508=>"110100100",
  38509=>"010011101",
  38510=>"111101010",
  38511=>"011000011",
  38512=>"001101010",
  38513=>"111010111",
  38514=>"101101000",
  38515=>"011100101",
  38516=>"101001110",
  38517=>"110000101",
  38518=>"110111111",
  38519=>"101001100",
  38520=>"110111001",
  38521=>"010011000",
  38522=>"111100000",
  38523=>"001111111",
  38524=>"111001000",
  38525=>"110100101",
  38526=>"111001101",
  38527=>"000100011",
  38528=>"100101000",
  38529=>"010000111",
  38530=>"101011100",
  38531=>"000001001",
  38532=>"111000001",
  38533=>"110100010",
  38534=>"011011110",
  38535=>"010111010",
  38536=>"100110111",
  38537=>"101110000",
  38538=>"011101111",
  38539=>"001101011",
  38540=>"011000011",
  38541=>"011011001",
  38542=>"110011100",
  38543=>"101101011",
  38544=>"011100100",
  38545=>"110110001",
  38546=>"000010000",
  38547=>"111110110",
  38548=>"101100010",
  38549=>"100000111",
  38550=>"100001111",
  38551=>"000000000",
  38552=>"111101001",
  38553=>"001001101",
  38554=>"111010101",
  38555=>"111110010",
  38556=>"111101001",
  38557=>"011001011",
  38558=>"001110110",
  38559=>"001111101",
  38560=>"111001100",
  38561=>"001111000",
  38562=>"100010000",
  38563=>"101110101",
  38564=>"100101000",
  38565=>"101000111",
  38566=>"010010100",
  38567=>"000011000",
  38568=>"100001000",
  38569=>"000000001",
  38570=>"001001110",
  38571=>"101101101",
  38572=>"110010010",
  38573=>"010001110",
  38574=>"001111100",
  38575=>"000001000",
  38576=>"101001111",
  38577=>"001011111",
  38578=>"001010110",
  38579=>"001100100",
  38580=>"011000110",
  38581=>"111000011",
  38582=>"001010000",
  38583=>"101000000",
  38584=>"001111000",
  38585=>"000111101",
  38586=>"101000100",
  38587=>"001000000",
  38588=>"010000011",
  38589=>"100001001",
  38590=>"101100100",
  38591=>"010010110",
  38592=>"100001111",
  38593=>"000110110",
  38594=>"101111010",
  38595=>"000111101",
  38596=>"111011100",
  38597=>"011110110",
  38598=>"010010111",
  38599=>"001101110",
  38600=>"011010000",
  38601=>"001100100",
  38602=>"101000101",
  38603=>"011000010",
  38604=>"011101010",
  38605=>"101001010",
  38606=>"101000010",
  38607=>"010001000",
  38608=>"011000100",
  38609=>"111100111",
  38610=>"100110101",
  38611=>"101110001",
  38612=>"000111100",
  38613=>"111011000",
  38614=>"011101000",
  38615=>"110000010",
  38616=>"000000000",
  38617=>"000010110",
  38618=>"101100000",
  38619=>"100001100",
  38620=>"001010101",
  38621=>"001010100",
  38622=>"010011101",
  38623=>"001101001",
  38624=>"101111001",
  38625=>"101000001",
  38626=>"100101100",
  38627=>"100111000",
  38628=>"010100000",
  38629=>"101100110",
  38630=>"110101011",
  38631=>"101100000",
  38632=>"010101111",
  38633=>"111110100",
  38634=>"100001010",
  38635=>"100011100",
  38636=>"101000110",
  38637=>"011111110",
  38638=>"100110011",
  38639=>"110000000",
  38640=>"000101111",
  38641=>"010001100",
  38642=>"000001100",
  38643=>"000111110",
  38644=>"001011100",
  38645=>"010101011",
  38646=>"000011101",
  38647=>"010000001",
  38648=>"011001100",
  38649=>"000011010",
  38650=>"100000110",
  38651=>"101101111",
  38652=>"011000001",
  38653=>"000001111",
  38654=>"001100010",
  38655=>"111111100",
  38656=>"010111010",
  38657=>"111110111",
  38658=>"110010011",
  38659=>"100001000",
  38660=>"010000010",
  38661=>"001101010",
  38662=>"010011111",
  38663=>"100101010",
  38664=>"111110011",
  38665=>"101011111",
  38666=>"011101101",
  38667=>"010000000",
  38668=>"000001000",
  38669=>"111011100",
  38670=>"101000011",
  38671=>"001000010",
  38672=>"110110101",
  38673=>"000110001",
  38674=>"001001100",
  38675=>"110100101",
  38676=>"111100111",
  38677=>"011000100",
  38678=>"100001001",
  38679=>"000001011",
  38680=>"011100101",
  38681=>"010111111",
  38682=>"100001000",
  38683=>"011011111",
  38684=>"011011010",
  38685=>"110100111",
  38686=>"110101100",
  38687=>"001100100",
  38688=>"011110100",
  38689=>"001001101",
  38690=>"000100001",
  38691=>"110100011",
  38692=>"101100100",
  38693=>"011000000",
  38694=>"011101011",
  38695=>"000011101",
  38696=>"011101011",
  38697=>"011111011",
  38698=>"101111110",
  38699=>"111001001",
  38700=>"101000010",
  38701=>"000000111",
  38702=>"010111001",
  38703=>"101111010",
  38704=>"000100111",
  38705=>"000010000",
  38706=>"010111110",
  38707=>"010100101",
  38708=>"001100000",
  38709=>"111101001",
  38710=>"010100111",
  38711=>"000110110",
  38712=>"001001000",
  38713=>"100110111",
  38714=>"011110100",
  38715=>"000100010",
  38716=>"000001010",
  38717=>"110011110",
  38718=>"101101100",
  38719=>"001100010",
  38720=>"100011010",
  38721=>"101101101",
  38722=>"001100001",
  38723=>"101001001",
  38724=>"110011011",
  38725=>"111101110",
  38726=>"100100101",
  38727=>"100101001",
  38728=>"100000010",
  38729=>"111111111",
  38730=>"000110101",
  38731=>"010001011",
  38732=>"010110000",
  38733=>"101100111",
  38734=>"010000001",
  38735=>"111111101",
  38736=>"010000011",
  38737=>"010000100",
  38738=>"111110000",
  38739=>"000000010",
  38740=>"001110001",
  38741=>"011110101",
  38742=>"100110101",
  38743=>"111011100",
  38744=>"010000000",
  38745=>"110110110",
  38746=>"100001001",
  38747=>"100001100",
  38748=>"011000111",
  38749=>"101011101",
  38750=>"110001010",
  38751=>"000101011",
  38752=>"001001101",
  38753=>"111100000",
  38754=>"101000011",
  38755=>"111101011",
  38756=>"001101101",
  38757=>"000001000",
  38758=>"001001000",
  38759=>"111010000",
  38760=>"000101011",
  38761=>"010000001",
  38762=>"101100111",
  38763=>"110000111",
  38764=>"101000001",
  38765=>"010111100",
  38766=>"100100101",
  38767=>"111011001",
  38768=>"011110011",
  38769=>"100101100",
  38770=>"001101000",
  38771=>"011000011",
  38772=>"110000000",
  38773=>"000101101",
  38774=>"010010110",
  38775=>"001101111",
  38776=>"011000000",
  38777=>"111010000",
  38778=>"010011001",
  38779=>"001111111",
  38780=>"110000100",
  38781=>"010101011",
  38782=>"101110101",
  38783=>"011010011",
  38784=>"010100101",
  38785=>"000011010",
  38786=>"011111110",
  38787=>"011100001",
  38788=>"011101001",
  38789=>"101011000",
  38790=>"101100100",
  38791=>"000000101",
  38792=>"101000000",
  38793=>"111011000",
  38794=>"000111011",
  38795=>"000110101",
  38796=>"000001010",
  38797=>"101001100",
  38798=>"001100001",
  38799=>"010111110",
  38800=>"001101000",
  38801=>"000111110",
  38802=>"000100110",
  38803=>"100111000",
  38804=>"011101011",
  38805=>"101011111",
  38806=>"011010001",
  38807=>"000110000",
  38808=>"110000100",
  38809=>"001000000",
  38810=>"011001110",
  38811=>"101010011",
  38812=>"110110110",
  38813=>"011001001",
  38814=>"001101000",
  38815=>"110001001",
  38816=>"000001101",
  38817=>"100001100",
  38818=>"000000001",
  38819=>"011101000",
  38820=>"001011000",
  38821=>"010011111",
  38822=>"111101011",
  38823=>"000000100",
  38824=>"010010000",
  38825=>"101000000",
  38826=>"011111011",
  38827=>"110011101",
  38828=>"010010100",
  38829=>"010110110",
  38830=>"001010010",
  38831=>"001111111",
  38832=>"101011111",
  38833=>"011001010",
  38834=>"000100101",
  38835=>"011010001",
  38836=>"111010101",
  38837=>"100110010",
  38838=>"010000010",
  38839=>"000110000",
  38840=>"001111100",
  38841=>"011101011",
  38842=>"111001111",
  38843=>"011011100",
  38844=>"101111001",
  38845=>"110011100",
  38846=>"001100111",
  38847=>"000111101",
  38848=>"100110111",
  38849=>"100110111",
  38850=>"101110001",
  38851=>"110011100",
  38852=>"111101101",
  38853=>"010000001",
  38854=>"100000000",
  38855=>"000011110",
  38856=>"010100001",
  38857=>"111001010",
  38858=>"101001011",
  38859=>"101010100",
  38860=>"100111001",
  38861=>"010111010",
  38862=>"111111110",
  38863=>"000001010",
  38864=>"011101010",
  38865=>"111110101",
  38866=>"100101001",
  38867=>"100100000",
  38868=>"101010111",
  38869=>"011101010",
  38870=>"010001000",
  38871=>"000000010",
  38872=>"000111100",
  38873=>"111101101",
  38874=>"111101101",
  38875=>"101011010",
  38876=>"001010000",
  38877=>"010010000",
  38878=>"110100000",
  38879=>"110101101",
  38880=>"111011100",
  38881=>"110001010",
  38882=>"101001101",
  38883=>"010010111",
  38884=>"010011110",
  38885=>"000111011",
  38886=>"011000000",
  38887=>"011010000",
  38888=>"010110110",
  38889=>"000101110",
  38890=>"010000001",
  38891=>"110100111",
  38892=>"110110011",
  38893=>"110111010",
  38894=>"011011000",
  38895=>"001010010",
  38896=>"010010001",
  38897=>"001011010",
  38898=>"100100110",
  38899=>"010100111",
  38900=>"010001110",
  38901=>"111110111",
  38902=>"000011110",
  38903=>"101111110",
  38904=>"111101110",
  38905=>"111010001",
  38906=>"011001100",
  38907=>"010001010",
  38908=>"101010111",
  38909=>"100101010",
  38910=>"000010100",
  38911=>"111100000",
  38912=>"110100110",
  38913=>"000100010",
  38914=>"001110100",
  38915=>"111100110",
  38916=>"001110000",
  38917=>"100110000",
  38918=>"110111110",
  38919=>"111111000",
  38920=>"111001011",
  38921=>"111001101",
  38922=>"000000010",
  38923=>"011011111",
  38924=>"110010000",
  38925=>"111101111",
  38926=>"011010000",
  38927=>"101101001",
  38928=>"001001011",
  38929=>"110110100",
  38930=>"000001001",
  38931=>"000100111",
  38932=>"000001100",
  38933=>"100011100",
  38934=>"010010011",
  38935=>"111001001",
  38936=>"101001101",
  38937=>"110101000",
  38938=>"110111111",
  38939=>"101011001",
  38940=>"111100100",
  38941=>"001011000",
  38942=>"010010100",
  38943=>"110011111",
  38944=>"010100101",
  38945=>"000111111",
  38946=>"000000011",
  38947=>"111100111",
  38948=>"101110001",
  38949=>"101100000",
  38950=>"111101010",
  38951=>"110110000",
  38952=>"000001001",
  38953=>"000111001",
  38954=>"111010000",
  38955=>"100111001",
  38956=>"100100000",
  38957=>"111010111",
  38958=>"001010011",
  38959=>"000010011",
  38960=>"110110011",
  38961=>"111100010",
  38962=>"001000110",
  38963=>"011001110",
  38964=>"110001111",
  38965=>"100010001",
  38966=>"000000011",
  38967=>"101101110",
  38968=>"111110011",
  38969=>"101100000",
  38970=>"000000100",
  38971=>"000011000",
  38972=>"000000010",
  38973=>"011100010",
  38974=>"011011111",
  38975=>"100001110",
  38976=>"000110111",
  38977=>"000111000",
  38978=>"000111100",
  38979=>"100100001",
  38980=>"010001111",
  38981=>"000101111",
  38982=>"011111111",
  38983=>"001101111",
  38984=>"100011001",
  38985=>"100000101",
  38986=>"000001010",
  38987=>"110100011",
  38988=>"100000100",
  38989=>"001001011",
  38990=>"001011010",
  38991=>"110100010",
  38992=>"011011100",
  38993=>"100100100",
  38994=>"011000011",
  38995=>"101010110",
  38996=>"110011000",
  38997=>"111110010",
  38998=>"100010001",
  38999=>"101110101",
  39000=>"001010101",
  39001=>"001000100",
  39002=>"100100010",
  39003=>"100011100",
  39004=>"101101110",
  39005=>"100000001",
  39006=>"011000100",
  39007=>"001011110",
  39008=>"001010001",
  39009=>"101000101",
  39010=>"010000110",
  39011=>"101101100",
  39012=>"101011101",
  39013=>"010100000",
  39014=>"000010000",
  39015=>"010001111",
  39016=>"010011010",
  39017=>"110001000",
  39018=>"111101001",
  39019=>"100101111",
  39020=>"101101011",
  39021=>"100010111",
  39022=>"111111000",
  39023=>"100100000",
  39024=>"000100000",
  39025=>"011110011",
  39026=>"000001100",
  39027=>"110000011",
  39028=>"000010100",
  39029=>"011000110",
  39030=>"101010101",
  39031=>"100011110",
  39032=>"010100100",
  39033=>"111110000",
  39034=>"110000001",
  39035=>"101100000",
  39036=>"011111110",
  39037=>"110100101",
  39038=>"011011110",
  39039=>"010101111",
  39040=>"111111001",
  39041=>"111010111",
  39042=>"110111010",
  39043=>"001001000",
  39044=>"101100001",
  39045=>"001110000",
  39046=>"010010110",
  39047=>"001000010",
  39048=>"011001111",
  39049=>"011100100",
  39050=>"110000110",
  39051=>"010101111",
  39052=>"011000000",
  39053=>"101011011",
  39054=>"011101110",
  39055=>"011010100",
  39056=>"110010010",
  39057=>"000101111",
  39058=>"001010010",
  39059=>"010000110",
  39060=>"000000001",
  39061=>"011000011",
  39062=>"111101010",
  39063=>"110000000",
  39064=>"111100011",
  39065=>"010010001",
  39066=>"110000000",
  39067=>"101001001",
  39068=>"111110011",
  39069=>"110111000",
  39070=>"011110000",
  39071=>"001011110",
  39072=>"011011011",
  39073=>"000111000",
  39074=>"010001001",
  39075=>"000001000",
  39076=>"110110100",
  39077=>"001111011",
  39078=>"110000001",
  39079=>"000001111",
  39080=>"001010100",
  39081=>"011101001",
  39082=>"010010101",
  39083=>"100001010",
  39084=>"101100100",
  39085=>"100001101",
  39086=>"000100100",
  39087=>"111101010",
  39088=>"110101010",
  39089=>"100011100",
  39090=>"101010010",
  39091=>"010011110",
  39092=>"000000100",
  39093=>"000010000",
  39094=>"100010000",
  39095=>"001000000",
  39096=>"000110000",
  39097=>"111110111",
  39098=>"010101011",
  39099=>"110000010",
  39100=>"011111110",
  39101=>"100100110",
  39102=>"011001101",
  39103=>"000111000",
  39104=>"001000010",
  39105=>"110100101",
  39106=>"111001111",
  39107=>"000000110",
  39108=>"100010000",
  39109=>"101010010",
  39110=>"000110111",
  39111=>"010011101",
  39112=>"110000010",
  39113=>"110001110",
  39114=>"011001011",
  39115=>"101100111",
  39116=>"010000010",
  39117=>"001000001",
  39118=>"101000110",
  39119=>"000000101",
  39120=>"000011010",
  39121=>"111110000",
  39122=>"000101010",
  39123=>"000011100",
  39124=>"110000110",
  39125=>"100010011",
  39126=>"111001111",
  39127=>"111000011",
  39128=>"100101111",
  39129=>"010110001",
  39130=>"010111110",
  39131=>"101110000",
  39132=>"100010101",
  39133=>"110110111",
  39134=>"101100111",
  39135=>"110011100",
  39136=>"101111100",
  39137=>"111101100",
  39138=>"101111100",
  39139=>"111110111",
  39140=>"001011010",
  39141=>"101011101",
  39142=>"000110011",
  39143=>"110010100",
  39144=>"001100100",
  39145=>"100011101",
  39146=>"010100011",
  39147=>"000000000",
  39148=>"111001110",
  39149=>"111011111",
  39150=>"000000011",
  39151=>"111000111",
  39152=>"111000110",
  39153=>"101111101",
  39154=>"111111010",
  39155=>"110001000",
  39156=>"001111001",
  39157=>"011011110",
  39158=>"011000011",
  39159=>"111100011",
  39160=>"000100111",
  39161=>"011010111",
  39162=>"001100101",
  39163=>"011011000",
  39164=>"010010010",
  39165=>"010100001",
  39166=>"001101001",
  39167=>"001010010",
  39168=>"101111101",
  39169=>"111010110",
  39170=>"110011100",
  39171=>"000001010",
  39172=>"100110100",
  39173=>"111001000",
  39174=>"000111110",
  39175=>"110110100",
  39176=>"000000101",
  39177=>"111111100",
  39178=>"100011001",
  39179=>"100101010",
  39180=>"100011101",
  39181=>"101000001",
  39182=>"000110001",
  39183=>"011001011",
  39184=>"010010111",
  39185=>"011000001",
  39186=>"101110010",
  39187=>"000101100",
  39188=>"001100011",
  39189=>"111010101",
  39190=>"100000000",
  39191=>"111110001",
  39192=>"110000011",
  39193=>"000010111",
  39194=>"101011011",
  39195=>"001111001",
  39196=>"100111110",
  39197=>"010000111",
  39198=>"111011011",
  39199=>"111100111",
  39200=>"001110111",
  39201=>"110101100",
  39202=>"001101111",
  39203=>"111100011",
  39204=>"111000000",
  39205=>"111010100",
  39206=>"011011001",
  39207=>"110011100",
  39208=>"001001000",
  39209=>"001001011",
  39210=>"001110000",
  39211=>"000101011",
  39212=>"101000000",
  39213=>"101101111",
  39214=>"100001011",
  39215=>"000100100",
  39216=>"111000100",
  39217=>"010010010",
  39218=>"001100000",
  39219=>"101111111",
  39220=>"001111110",
  39221=>"100011000",
  39222=>"000010100",
  39223=>"011101101",
  39224=>"010111010",
  39225=>"101000100",
  39226=>"001111011",
  39227=>"001101000",
  39228=>"100010101",
  39229=>"000101010",
  39230=>"100100111",
  39231=>"111111111",
  39232=>"110100111",
  39233=>"111111000",
  39234=>"001001000",
  39235=>"010110100",
  39236=>"001111000",
  39237=>"011001000",
  39238=>"111011111",
  39239=>"110100000",
  39240=>"000010001",
  39241=>"001101101",
  39242=>"111001011",
  39243=>"101110000",
  39244=>"110111010",
  39245=>"001110011",
  39246=>"101101000",
  39247=>"111010000",
  39248=>"111010111",
  39249=>"011011111",
  39250=>"100000111",
  39251=>"000001011",
  39252=>"010100110",
  39253=>"011011011",
  39254=>"110001110",
  39255=>"101011111",
  39256=>"000011000",
  39257=>"100010001",
  39258=>"011010001",
  39259=>"110101100",
  39260=>"111001011",
  39261=>"000010000",
  39262=>"000100010",
  39263=>"101001101",
  39264=>"111000110",
  39265=>"110101100",
  39266=>"100011011",
  39267=>"101101001",
  39268=>"000110011",
  39269=>"001000001",
  39270=>"100100010",
  39271=>"101111001",
  39272=>"110011001",
  39273=>"110111101",
  39274=>"011110001",
  39275=>"010100010",
  39276=>"111100111",
  39277=>"010011111",
  39278=>"010110111",
  39279=>"111101001",
  39280=>"010000111",
  39281=>"010000011",
  39282=>"111100101",
  39283=>"101011101",
  39284=>"100110001",
  39285=>"011000110",
  39286=>"010100000",
  39287=>"001000100",
  39288=>"000101110",
  39289=>"100110000",
  39290=>"110101100",
  39291=>"100100000",
  39292=>"011001100",
  39293=>"100000010",
  39294=>"111110000",
  39295=>"110111101",
  39296=>"011000111",
  39297=>"000110111",
  39298=>"100111010",
  39299=>"010100011",
  39300=>"110111000",
  39301=>"100011011",
  39302=>"111111001",
  39303=>"000100011",
  39304=>"010100001",
  39305=>"100010011",
  39306=>"011010100",
  39307=>"111101111",
  39308=>"110100000",
  39309=>"001111110",
  39310=>"111010101",
  39311=>"100110111",
  39312=>"111101100",
  39313=>"010000010",
  39314=>"111101111",
  39315=>"000100101",
  39316=>"100000011",
  39317=>"101100010",
  39318=>"010111110",
  39319=>"011101001",
  39320=>"001010110",
  39321=>"100000100",
  39322=>"101100000",
  39323=>"100110001",
  39324=>"011110101",
  39325=>"011101110",
  39326=>"010111101",
  39327=>"101111000",
  39328=>"100101001",
  39329=>"011011001",
  39330=>"000000110",
  39331=>"000001010",
  39332=>"001000100",
  39333=>"011000011",
  39334=>"110101000",
  39335=>"010100000",
  39336=>"001111111",
  39337=>"101000110",
  39338=>"100011000",
  39339=>"000111000",
  39340=>"111111001",
  39341=>"101011101",
  39342=>"101111000",
  39343=>"000100010",
  39344=>"100111010",
  39345=>"010111001",
  39346=>"001010100",
  39347=>"100100110",
  39348=>"100000101",
  39349=>"111011100",
  39350=>"110001001",
  39351=>"111001110",
  39352=>"001100110",
  39353=>"010011110",
  39354=>"101010110",
  39355=>"101111110",
  39356=>"101110101",
  39357=>"111101101",
  39358=>"001000001",
  39359=>"010001001",
  39360=>"101101000",
  39361=>"001011101",
  39362=>"011101001",
  39363=>"100010001",
  39364=>"000100010",
  39365=>"011011011",
  39366=>"101100010",
  39367=>"000000000",
  39368=>"001111000",
  39369=>"101011001",
  39370=>"010001010",
  39371=>"000001001",
  39372=>"101000011",
  39373=>"000010111",
  39374=>"001111100",
  39375=>"110011010",
  39376=>"111100110",
  39377=>"000111001",
  39378=>"000010001",
  39379=>"010000011",
  39380=>"111111111",
  39381=>"100010100",
  39382=>"001100011",
  39383=>"110001001",
  39384=>"001111000",
  39385=>"000011100",
  39386=>"010001100",
  39387=>"101101000",
  39388=>"100010100",
  39389=>"101000001",
  39390=>"001010111",
  39391=>"011110000",
  39392=>"111111011",
  39393=>"111011011",
  39394=>"110010011",
  39395=>"111001000",
  39396=>"010100111",
  39397=>"111110110",
  39398=>"111101010",
  39399=>"101100100",
  39400=>"000000011",
  39401=>"100100100",
  39402=>"001000011",
  39403=>"000111101",
  39404=>"010111010",
  39405=>"000011010",
  39406=>"111000101",
  39407=>"000000111",
  39408=>"011111001",
  39409=>"000010100",
  39410=>"111101001",
  39411=>"111100001",
  39412=>"001100010",
  39413=>"011100000",
  39414=>"111100011",
  39415=>"001100100",
  39416=>"100010100",
  39417=>"001100011",
  39418=>"101001000",
  39419=>"010111011",
  39420=>"110011111",
  39421=>"010101010",
  39422=>"010000111",
  39423=>"110000110",
  39424=>"001011100",
  39425=>"000101011",
  39426=>"011101110",
  39427=>"100001101",
  39428=>"011101100",
  39429=>"100111100",
  39430=>"011101101",
  39431=>"101111100",
  39432=>"100011011",
  39433=>"000101111",
  39434=>"010100110",
  39435=>"111111011",
  39436=>"001010001",
  39437=>"000001001",
  39438=>"101011110",
  39439=>"010000001",
  39440=>"110011000",
  39441=>"000101101",
  39442=>"000111111",
  39443=>"100110010",
  39444=>"000001100",
  39445=>"101101111",
  39446=>"111101100",
  39447=>"011010110",
  39448=>"111111100",
  39449=>"100011000",
  39450=>"101110110",
  39451=>"010100001",
  39452=>"000110011",
  39453=>"101010011",
  39454=>"111111111",
  39455=>"101000100",
  39456=>"000000000",
  39457=>"000001001",
  39458=>"000001010",
  39459=>"110101111",
  39460=>"000011011",
  39461=>"001011001",
  39462=>"111101001",
  39463=>"110101010",
  39464=>"000110110",
  39465=>"000001010",
  39466=>"100100111",
  39467=>"010110011",
  39468=>"000111101",
  39469=>"100010001",
  39470=>"100010000",
  39471=>"000010100",
  39472=>"101001101",
  39473=>"010101010",
  39474=>"101111010",
  39475=>"101001100",
  39476=>"100101001",
  39477=>"100110110",
  39478=>"011110100",
  39479=>"101111011",
  39480=>"111000101",
  39481=>"011001000",
  39482=>"010001001",
  39483=>"100101110",
  39484=>"111111001",
  39485=>"101001110",
  39486=>"010111001",
  39487=>"111100011",
  39488=>"101100010",
  39489=>"100010011",
  39490=>"000001101",
  39491=>"111111100",
  39492=>"111001101",
  39493=>"110110111",
  39494=>"010000001",
  39495=>"111101111",
  39496=>"101001010",
  39497=>"011000011",
  39498=>"000010001",
  39499=>"000010000",
  39500=>"111001101",
  39501=>"001110011",
  39502=>"111001011",
  39503=>"001101011",
  39504=>"000100101",
  39505=>"111001000",
  39506=>"011100111",
  39507=>"010011110",
  39508=>"111110111",
  39509=>"001000000",
  39510=>"111001101",
  39511=>"011010001",
  39512=>"100111111",
  39513=>"101010001",
  39514=>"101101011",
  39515=>"000001101",
  39516=>"010100110",
  39517=>"010100100",
  39518=>"101010000",
  39519=>"110011110",
  39520=>"001111100",
  39521=>"000111111",
  39522=>"111100000",
  39523=>"101000001",
  39524=>"100100000",
  39525=>"100101011",
  39526=>"010010001",
  39527=>"000001000",
  39528=>"100000010",
  39529=>"000100010",
  39530=>"101011011",
  39531=>"111110111",
  39532=>"000101001",
  39533=>"101111010",
  39534=>"011011011",
  39535=>"010010110",
  39536=>"000010110",
  39537=>"101001011",
  39538=>"010101111",
  39539=>"100000000",
  39540=>"101010100",
  39541=>"101001011",
  39542=>"010111111",
  39543=>"101011001",
  39544=>"011110111",
  39545=>"011000111",
  39546=>"000100000",
  39547=>"000100101",
  39548=>"010110000",
  39549=>"110100111",
  39550=>"011000101",
  39551=>"101100100",
  39552=>"000000110",
  39553=>"001111110",
  39554=>"110010101",
  39555=>"001110011",
  39556=>"000110101",
  39557=>"011000100",
  39558=>"000110011",
  39559=>"110101011",
  39560=>"000010001",
  39561=>"100100010",
  39562=>"000001110",
  39563=>"001000000",
  39564=>"101010110",
  39565=>"010001101",
  39566=>"011001011",
  39567=>"111001011",
  39568=>"000100110",
  39569=>"100010010",
  39570=>"001111000",
  39571=>"000000111",
  39572=>"011101010",
  39573=>"010100111",
  39574=>"000100111",
  39575=>"001110111",
  39576=>"101101101",
  39577=>"010010001",
  39578=>"011111011",
  39579=>"101111110",
  39580=>"011110000",
  39581=>"100100000",
  39582=>"000000000",
  39583=>"110010110",
  39584=>"010010111",
  39585=>"000111110",
  39586=>"011110001",
  39587=>"000100110",
  39588=>"001000111",
  39589=>"101101001",
  39590=>"001000010",
  39591=>"110000001",
  39592=>"011001000",
  39593=>"010100100",
  39594=>"101010101",
  39595=>"001111011",
  39596=>"011111011",
  39597=>"100100100",
  39598=>"010111110",
  39599=>"111011000",
  39600=>"111110000",
  39601=>"110000100",
  39602=>"001011101",
  39603=>"100101100",
  39604=>"000000101",
  39605=>"001001011",
  39606=>"000011010",
  39607=>"011011100",
  39608=>"001101001",
  39609=>"011101111",
  39610=>"111110000",
  39611=>"110010101",
  39612=>"110111110",
  39613=>"110100100",
  39614=>"100000100",
  39615=>"101011101",
  39616=>"101101011",
  39617=>"101000100",
  39618=>"001101110",
  39619=>"101100010",
  39620=>"111100100",
  39621=>"000101001",
  39622=>"001100110",
  39623=>"111101111",
  39624=>"101011010",
  39625=>"001100100",
  39626=>"101011111",
  39627=>"001001101",
  39628=>"000101001",
  39629=>"110100101",
  39630=>"000011101",
  39631=>"100000101",
  39632=>"001011011",
  39633=>"011011101",
  39634=>"010010111",
  39635=>"111111011",
  39636=>"101000110",
  39637=>"100001010",
  39638=>"101100110",
  39639=>"010000111",
  39640=>"010000011",
  39641=>"000110000",
  39642=>"110111011",
  39643=>"001000110",
  39644=>"101001100",
  39645=>"010001000",
  39646=>"110001000",
  39647=>"010110101",
  39648=>"000111100",
  39649=>"111000010",
  39650=>"111011000",
  39651=>"111101100",
  39652=>"111110110",
  39653=>"100011001",
  39654=>"100000110",
  39655=>"100000001",
  39656=>"011111111",
  39657=>"111010111",
  39658=>"101100001",
  39659=>"011000110",
  39660=>"111001010",
  39661=>"100111111",
  39662=>"011000100",
  39663=>"010010010",
  39664=>"000000000",
  39665=>"001101111",
  39666=>"011101100",
  39667=>"100000011",
  39668=>"100111100",
  39669=>"010111000",
  39670=>"000001100",
  39671=>"010101110",
  39672=>"101100101",
  39673=>"111100110",
  39674=>"101000000",
  39675=>"001010011",
  39676=>"001001111",
  39677=>"010010110",
  39678=>"101001110",
  39679=>"010100001",
  39680=>"001101110",
  39681=>"000100100",
  39682=>"000111100",
  39683=>"000011011",
  39684=>"100011010",
  39685=>"000110111",
  39686=>"100101011",
  39687=>"110111110",
  39688=>"111100011",
  39689=>"100111111",
  39690=>"110101111",
  39691=>"010001001",
  39692=>"001101011",
  39693=>"111100111",
  39694=>"111010111",
  39695=>"000000101",
  39696=>"111111000",
  39697=>"100010100",
  39698=>"000000011",
  39699=>"110101000",
  39700=>"100010000",
  39701=>"101101110",
  39702=>"010011000",
  39703=>"010100010",
  39704=>"011101100",
  39705=>"001100100",
  39706=>"000000111",
  39707=>"010000000",
  39708=>"011101000",
  39709=>"101010101",
  39710=>"000000111",
  39711=>"101000011",
  39712=>"001001000",
  39713=>"101001111",
  39714=>"101000110",
  39715=>"000111111",
  39716=>"011101110",
  39717=>"010111101",
  39718=>"111001101",
  39719=>"010000001",
  39720=>"100011111",
  39721=>"001011101",
  39722=>"110001100",
  39723=>"100001000",
  39724=>"011001101",
  39725=>"001000000",
  39726=>"100111101",
  39727=>"110111110",
  39728=>"111000111",
  39729=>"000010110",
  39730=>"111001011",
  39731=>"100110110",
  39732=>"101010000",
  39733=>"110001010",
  39734=>"011100101",
  39735=>"110111011",
  39736=>"101000111",
  39737=>"011010011",
  39738=>"001000011",
  39739=>"001010100",
  39740=>"001110000",
  39741=>"100010110",
  39742=>"101111011",
  39743=>"011110110",
  39744=>"010111010",
  39745=>"100101010",
  39746=>"110001000",
  39747=>"111101110",
  39748=>"100011011",
  39749=>"100000000",
  39750=>"010100100",
  39751=>"000110110",
  39752=>"100001111",
  39753=>"110001111",
  39754=>"101011010",
  39755=>"010100100",
  39756=>"011110111",
  39757=>"111101001",
  39758=>"111011011",
  39759=>"100110001",
  39760=>"111110111",
  39761=>"100101001",
  39762=>"000111010",
  39763=>"010100111",
  39764=>"111001111",
  39765=>"001100100",
  39766=>"101100101",
  39767=>"011000010",
  39768=>"000000000",
  39769=>"101011100",
  39770=>"100000101",
  39771=>"111010111",
  39772=>"101011110",
  39773=>"110000111",
  39774=>"111111011",
  39775=>"000100110",
  39776=>"010011001",
  39777=>"110010011",
  39778=>"010100010",
  39779=>"100010100",
  39780=>"010100110",
  39781=>"111010111",
  39782=>"000101101",
  39783=>"011001001",
  39784=>"100100100",
  39785=>"000110000",
  39786=>"001011011",
  39787=>"001010100",
  39788=>"101000001",
  39789=>"111001111",
  39790=>"000000111",
  39791=>"001001000",
  39792=>"011001101",
  39793=>"000101011",
  39794=>"010011101",
  39795=>"000111010",
  39796=>"110110011",
  39797=>"110101001",
  39798=>"101100000",
  39799=>"010001001",
  39800=>"101000010",
  39801=>"011111010",
  39802=>"110010001",
  39803=>"001110000",
  39804=>"111111101",
  39805=>"010010011",
  39806=>"101100100",
  39807=>"100111111",
  39808=>"101001111",
  39809=>"100101111",
  39810=>"101001101",
  39811=>"010110110",
  39812=>"110100000",
  39813=>"111010011",
  39814=>"001110110",
  39815=>"000110110",
  39816=>"100111100",
  39817=>"011011000",
  39818=>"000111111",
  39819=>"000101101",
  39820=>"110011100",
  39821=>"101010110",
  39822=>"111011100",
  39823=>"110111101",
  39824=>"001100110",
  39825=>"010000000",
  39826=>"011011001",
  39827=>"000111101",
  39828=>"000100110",
  39829=>"010111000",
  39830=>"000000001",
  39831=>"110000111",
  39832=>"110010000",
  39833=>"000110110",
  39834=>"100100000",
  39835=>"010011110",
  39836=>"001001110",
  39837=>"001001000",
  39838=>"000010000",
  39839=>"011110000",
  39840=>"110011111",
  39841=>"100110010",
  39842=>"100000011",
  39843=>"011010010",
  39844=>"101100001",
  39845=>"010111010",
  39846=>"010110101",
  39847=>"001000001",
  39848=>"000111110",
  39849=>"111011011",
  39850=>"011010101",
  39851=>"001100000",
  39852=>"010111011",
  39853=>"111100100",
  39854=>"100000011",
  39855=>"111111110",
  39856=>"001001000",
  39857=>"111101110",
  39858=>"011101010",
  39859=>"101110101",
  39860=>"101010101",
  39861=>"100001010",
  39862=>"111100100",
  39863=>"101101111",
  39864=>"100100110",
  39865=>"110111111",
  39866=>"000010111",
  39867=>"101010010",
  39868=>"101100101",
  39869=>"111011000",
  39870=>"110100010",
  39871=>"010100001",
  39872=>"101101101",
  39873=>"011011110",
  39874=>"001111100",
  39875=>"011011010",
  39876=>"101110100",
  39877=>"011001010",
  39878=>"010111111",
  39879=>"010011111",
  39880=>"001001011",
  39881=>"001111100",
  39882=>"110001111",
  39883=>"100010111",
  39884=>"100101110",
  39885=>"111000010",
  39886=>"111111100",
  39887=>"010110001",
  39888=>"111110111",
  39889=>"000000010",
  39890=>"111111010",
  39891=>"111001011",
  39892=>"000101011",
  39893=>"100011101",
  39894=>"000011001",
  39895=>"000010001",
  39896=>"000101000",
  39897=>"110010101",
  39898=>"100000101",
  39899=>"110101100",
  39900=>"100100110",
  39901=>"101101101",
  39902=>"100010000",
  39903=>"101101001",
  39904=>"111100000",
  39905=>"001001111",
  39906=>"100011111",
  39907=>"011001100",
  39908=>"000011010",
  39909=>"011101101",
  39910=>"001100110",
  39911=>"011011101",
  39912=>"001110000",
  39913=>"011111110",
  39914=>"001110000",
  39915=>"000111100",
  39916=>"101010111",
  39917=>"011000001",
  39918=>"000110010",
  39919=>"001001000",
  39920=>"010111000",
  39921=>"000010010",
  39922=>"001010101",
  39923=>"101011001",
  39924=>"000010110",
  39925=>"100011011",
  39926=>"010000011",
  39927=>"010110101",
  39928=>"011110110",
  39929=>"110001010",
  39930=>"111111111",
  39931=>"011010000",
  39932=>"000000101",
  39933=>"110110101",
  39934=>"001000100",
  39935=>"011101010",
  39936=>"001111111",
  39937=>"110100101",
  39938=>"110001101",
  39939=>"101101001",
  39940=>"001010111",
  39941=>"101001101",
  39942=>"010000010",
  39943=>"101111111",
  39944=>"100001101",
  39945=>"100111100",
  39946=>"100000101",
  39947=>"001001000",
  39948=>"001011000",
  39949=>"011011110",
  39950=>"110101001",
  39951=>"110000101",
  39952=>"110111111",
  39953=>"000001111",
  39954=>"010011011",
  39955=>"100011110",
  39956=>"100010001",
  39957=>"100100101",
  39958=>"111100110",
  39959=>"000111110",
  39960=>"000110011",
  39961=>"110101011",
  39962=>"011101111",
  39963=>"000100000",
  39964=>"111000111",
  39965=>"001010100",
  39966=>"111000000",
  39967=>"101010010",
  39968=>"100010100",
  39969=>"000010010",
  39970=>"011110111",
  39971=>"111000110",
  39972=>"000000010",
  39973=>"111010100",
  39974=>"101110000",
  39975=>"111110110",
  39976=>"001010000",
  39977=>"001100110",
  39978=>"000111101",
  39979=>"101010010",
  39980=>"100010000",
  39981=>"001000001",
  39982=>"010111100",
  39983=>"100100101",
  39984=>"000100101",
  39985=>"111011111",
  39986=>"110100010",
  39987=>"000011000",
  39988=>"101100000",
  39989=>"100011011",
  39990=>"111010101",
  39991=>"110111001",
  39992=>"100010001",
  39993=>"100100001",
  39994=>"001011000",
  39995=>"011101100",
  39996=>"010110001",
  39997=>"110010001",
  39998=>"110111111",
  39999=>"110110011",
  40000=>"111111111",
  40001=>"100100000",
  40002=>"110101000",
  40003=>"111101110",
  40004=>"000100101",
  40005=>"010101100",
  40006=>"001110100",
  40007=>"000111100",
  40008=>"001110001",
  40009=>"111001111",
  40010=>"010111111",
  40011=>"101110000",
  40012=>"001100001",
  40013=>"011110000",
  40014=>"101010111",
  40015=>"010101000",
  40016=>"101110011",
  40017=>"011011011",
  40018=>"010010111",
  40019=>"010010101",
  40020=>"111101010",
  40021=>"010111001",
  40022=>"010110010",
  40023=>"111010101",
  40024=>"011111111",
  40025=>"101010101",
  40026=>"011101000",
  40027=>"111100011",
  40028=>"010101110",
  40029=>"101000010",
  40030=>"011010001",
  40031=>"101000100",
  40032=>"010111001",
  40033=>"000001010",
  40034=>"000001010",
  40035=>"001111111",
  40036=>"100100010",
  40037=>"010110011",
  40038=>"001100100",
  40039=>"111001011",
  40040=>"011001010",
  40041=>"100110001",
  40042=>"011000000",
  40043=>"111011011",
  40044=>"101111100",
  40045=>"001100110",
  40046=>"100010001",
  40047=>"110000001",
  40048=>"001100111",
  40049=>"010111110",
  40050=>"111011101",
  40051=>"100100111",
  40052=>"100001100",
  40053=>"010001010",
  40054=>"101001100",
  40055=>"110011010",
  40056=>"010101100",
  40057=>"100000111",
  40058=>"101101111",
  40059=>"100100001",
  40060=>"110011010",
  40061=>"010010001",
  40062=>"100000101",
  40063=>"101001000",
  40064=>"110001001",
  40065=>"101000010",
  40066=>"110001101",
  40067=>"111100100",
  40068=>"111000000",
  40069=>"010110110",
  40070=>"001111011",
  40071=>"000101001",
  40072=>"011111011",
  40073=>"000011100",
  40074=>"000000000",
  40075=>"100111100",
  40076=>"000001010",
  40077=>"100000010",
  40078=>"110011100",
  40079=>"010011010",
  40080=>"010100001",
  40081=>"111011010",
  40082=>"001000110",
  40083=>"101000010",
  40084=>"101101000",
  40085=>"001110101",
  40086=>"110111111",
  40087=>"001011001",
  40088=>"101110110",
  40089=>"100001101",
  40090=>"101101011",
  40091=>"010001010",
  40092=>"111001000",
  40093=>"100110001",
  40094=>"011100101",
  40095=>"110001111",
  40096=>"110100110",
  40097=>"011110000",
  40098=>"000010000",
  40099=>"110101111",
  40100=>"000111010",
  40101=>"011010110",
  40102=>"010011111",
  40103=>"000000010",
  40104=>"011101000",
  40105=>"001001101",
  40106=>"111001101",
  40107=>"000010011",
  40108=>"110011000",
  40109=>"000110010",
  40110=>"100001111",
  40111=>"110010111",
  40112=>"001100101",
  40113=>"110101010",
  40114=>"010110101",
  40115=>"101001000",
  40116=>"010111011",
  40117=>"111110010",
  40118=>"000010000",
  40119=>"000010111",
  40120=>"111100010",
  40121=>"101000000",
  40122=>"110011001",
  40123=>"010100010",
  40124=>"110010101",
  40125=>"010011110",
  40126=>"101000000",
  40127=>"010101101",
  40128=>"001111111",
  40129=>"000010010",
  40130=>"101000011",
  40131=>"111111111",
  40132=>"010101101",
  40133=>"011111010",
  40134=>"110110000",
  40135=>"011110000",
  40136=>"001111100",
  40137=>"111010001",
  40138=>"111111000",
  40139=>"010011010",
  40140=>"111100000",
  40141=>"110110001",
  40142=>"110100110",
  40143=>"011000001",
  40144=>"110110000",
  40145=>"010001100",
  40146=>"100100100",
  40147=>"110101111",
  40148=>"111000100",
  40149=>"000011111",
  40150=>"011101110",
  40151=>"110011010",
  40152=>"001111000",
  40153=>"000101100",
  40154=>"001010100",
  40155=>"111110001",
  40156=>"101001110",
  40157=>"000010000",
  40158=>"101011011",
  40159=>"001100100",
  40160=>"110101011",
  40161=>"100100000",
  40162=>"000110100",
  40163=>"101010000",
  40164=>"011100110",
  40165=>"000010111",
  40166=>"110100001",
  40167=>"101010011",
  40168=>"000011000",
  40169=>"100100100",
  40170=>"010001110",
  40171=>"011101000",
  40172=>"010111111",
  40173=>"110011110",
  40174=>"010111110",
  40175=>"010000010",
  40176=>"001000011",
  40177=>"001110110",
  40178=>"101101000",
  40179=>"110001110",
  40180=>"011001101",
  40181=>"110111110",
  40182=>"000100000",
  40183=>"001001010",
  40184=>"100110111",
  40185=>"000100010",
  40186=>"010101100",
  40187=>"101101111",
  40188=>"111001100",
  40189=>"011111111",
  40190=>"100111000",
  40191=>"100111100",
  40192=>"110111101",
  40193=>"100111100",
  40194=>"100100100",
  40195=>"100010000",
  40196=>"001111011",
  40197=>"111101001",
  40198=>"100001110",
  40199=>"011110010",
  40200=>"111110101",
  40201=>"011001011",
  40202=>"100011001",
  40203=>"111100101",
  40204=>"111110001",
  40205=>"000101110",
  40206=>"111111000",
  40207=>"110011100",
  40208=>"011011010",
  40209=>"011011000",
  40210=>"001000010",
  40211=>"111011111",
  40212=>"000100111",
  40213=>"001001001",
  40214=>"000100110",
  40215=>"100010011",
  40216=>"001011101",
  40217=>"101000101",
  40218=>"101111100",
  40219=>"010000101",
  40220=>"010010001",
  40221=>"010111111",
  40222=>"111010000",
  40223=>"111110110",
  40224=>"110100100",
  40225=>"101010100",
  40226=>"011100000",
  40227=>"110010010",
  40228=>"101011100",
  40229=>"111100101",
  40230=>"101001000",
  40231=>"000101001",
  40232=>"101011011",
  40233=>"101010011",
  40234=>"000000010",
  40235=>"000101010",
  40236=>"010010110",
  40237=>"000110011",
  40238=>"001111001",
  40239=>"100010011",
  40240=>"111110111",
  40241=>"011101010",
  40242=>"100001101",
  40243=>"110001011",
  40244=>"011011101",
  40245=>"111101010",
  40246=>"010100001",
  40247=>"000100100",
  40248=>"000011011",
  40249=>"011000110",
  40250=>"100001010",
  40251=>"010011100",
  40252=>"100100010",
  40253=>"100100010",
  40254=>"010111001",
  40255=>"100010111",
  40256=>"010100100",
  40257=>"000011110",
  40258=>"101110101",
  40259=>"010110000",
  40260=>"111110101",
  40261=>"011011101",
  40262=>"110110011",
  40263=>"010101100",
  40264=>"100000000",
  40265=>"010010001",
  40266=>"010010110",
  40267=>"000110001",
  40268=>"101110111",
  40269=>"100001011",
  40270=>"000011101",
  40271=>"101110000",
  40272=>"101001111",
  40273=>"010000001",
  40274=>"011110111",
  40275=>"110111100",
  40276=>"011101101",
  40277=>"000110111",
  40278=>"110100010",
  40279=>"011011001",
  40280=>"001000001",
  40281=>"010011010",
  40282=>"100011010",
  40283=>"111011111",
  40284=>"100110111",
  40285=>"101111000",
  40286=>"000111001",
  40287=>"011011011",
  40288=>"111111001",
  40289=>"001000101",
  40290=>"111001101",
  40291=>"110101010",
  40292=>"101100010",
  40293=>"011011001",
  40294=>"001110001",
  40295=>"000111111",
  40296=>"100111011",
  40297=>"000000100",
  40298=>"111111010",
  40299=>"011010101",
  40300=>"111111101",
  40301=>"110111000",
  40302=>"011111001",
  40303=>"010100010",
  40304=>"010010010",
  40305=>"101100110",
  40306=>"110111010",
  40307=>"000000111",
  40308=>"010000101",
  40309=>"111110010",
  40310=>"010000111",
  40311=>"111000010",
  40312=>"111011010",
  40313=>"110011000",
  40314=>"110000010",
  40315=>"001100111",
  40316=>"000111101",
  40317=>"101011010",
  40318=>"101110111",
  40319=>"001011101",
  40320=>"001011111",
  40321=>"000010000",
  40322=>"101001101",
  40323=>"111101111",
  40324=>"001001010",
  40325=>"011110011",
  40326=>"001111011",
  40327=>"000110111",
  40328=>"110000001",
  40329=>"000110100",
  40330=>"011010011",
  40331=>"111011001",
  40332=>"000011110",
  40333=>"110101111",
  40334=>"100111111",
  40335=>"110101101",
  40336=>"000010100",
  40337=>"110110001",
  40338=>"010000001",
  40339=>"100000011",
  40340=>"000000001",
  40341=>"000011010",
  40342=>"101111101",
  40343=>"110100011",
  40344=>"011100100",
  40345=>"111011110",
  40346=>"111010111",
  40347=>"110010000",
  40348=>"110101000",
  40349=>"101001100",
  40350=>"101001100",
  40351=>"110110110",
  40352=>"101100100",
  40353=>"001111111",
  40354=>"100110110",
  40355=>"100100110",
  40356=>"111100111",
  40357=>"000000100",
  40358=>"011100100",
  40359=>"010011010",
  40360=>"000010001",
  40361=>"111100010",
  40362=>"011000100",
  40363=>"100100100",
  40364=>"110100100",
  40365=>"100010100",
  40366=>"001010100",
  40367=>"100011010",
  40368=>"101001011",
  40369=>"011111001",
  40370=>"100001001",
  40371=>"111001100",
  40372=>"010001011",
  40373=>"001110010",
  40374=>"100011101",
  40375=>"111101010",
  40376=>"101000001",
  40377=>"101101011",
  40378=>"001001100",
  40379=>"000010000",
  40380=>"011000100",
  40381=>"110011011",
  40382=>"101010000",
  40383=>"000011010",
  40384=>"111100111",
  40385=>"111010000",
  40386=>"000011101",
  40387=>"111110011",
  40388=>"111000000",
  40389=>"101111011",
  40390=>"101110110",
  40391=>"000011101",
  40392=>"010101000",
  40393=>"000101100",
  40394=>"100010000",
  40395=>"000000001",
  40396=>"010000000",
  40397=>"011011101",
  40398=>"011011110",
  40399=>"100100111",
  40400=>"011111101",
  40401=>"011110010",
  40402=>"110110001",
  40403=>"101100111",
  40404=>"001000110",
  40405=>"011011011",
  40406=>"010011000",
  40407=>"111000001",
  40408=>"101001010",
  40409=>"011101000",
  40410=>"100110100",
  40411=>"101101000",
  40412=>"111010101",
  40413=>"010000110",
  40414=>"000101011",
  40415=>"010011111",
  40416=>"110111101",
  40417=>"111111000",
  40418=>"011111000",
  40419=>"000110010",
  40420=>"110100101",
  40421=>"000010011",
  40422=>"111010100",
  40423=>"000011111",
  40424=>"111110111",
  40425=>"000101110",
  40426=>"111000001",
  40427=>"011100111",
  40428=>"000111001",
  40429=>"100010000",
  40430=>"101110100",
  40431=>"001101011",
  40432=>"000001101",
  40433=>"001110101",
  40434=>"110010010",
  40435=>"000000110",
  40436=>"001101101",
  40437=>"111111111",
  40438=>"110010011",
  40439=>"100011110",
  40440=>"110101010",
  40441=>"011101001",
  40442=>"111110100",
  40443=>"011110111",
  40444=>"101101100",
  40445=>"111011000",
  40446=>"000010110",
  40447=>"100010111",
  40448=>"110001010",
  40449=>"110001110",
  40450=>"001110100",
  40451=>"101110101",
  40452=>"001111001",
  40453=>"011001011",
  40454=>"001001011",
  40455=>"101111111",
  40456=>"011001011",
  40457=>"110001001",
  40458=>"101010011",
  40459=>"000010100",
  40460=>"110001110",
  40461=>"010010000",
  40462=>"001010110",
  40463=>"011100110",
  40464=>"110001001",
  40465=>"011011011",
  40466=>"111011110",
  40467=>"001001101",
  40468=>"010111111",
  40469=>"100000001",
  40470=>"101111011",
  40471=>"101010010",
  40472=>"010000110",
  40473=>"111101010",
  40474=>"110000011",
  40475=>"000100111",
  40476=>"100001101",
  40477=>"110100110",
  40478=>"011011101",
  40479=>"111011100",
  40480=>"010101111",
  40481=>"100100011",
  40482=>"111011100",
  40483=>"011000111",
  40484=>"110100001",
  40485=>"010010110",
  40486=>"000110000",
  40487=>"111001101",
  40488=>"110110000",
  40489=>"110101000",
  40490=>"001010000",
  40491=>"110111111",
  40492=>"011000101",
  40493=>"001110100",
  40494=>"011100110",
  40495=>"011100101",
  40496=>"001100111",
  40497=>"010010011",
  40498=>"111111110",
  40499=>"001010010",
  40500=>"000010000",
  40501=>"101100011",
  40502=>"111000101",
  40503=>"000011100",
  40504=>"101010101",
  40505=>"010100100",
  40506=>"001100011",
  40507=>"010111100",
  40508=>"001100001",
  40509=>"000100111",
  40510=>"101010001",
  40511=>"000101101",
  40512=>"000100000",
  40513=>"110000100",
  40514=>"011101101",
  40515=>"110111111",
  40516=>"110011110",
  40517=>"010010100",
  40518=>"001000111",
  40519=>"011010011",
  40520=>"001011110",
  40521=>"111111000",
  40522=>"011010111",
  40523=>"011100101",
  40524=>"011110010",
  40525=>"010001011",
  40526=>"111111001",
  40527=>"011000000",
  40528=>"111101011",
  40529=>"010101010",
  40530=>"101011001",
  40531=>"100000111",
  40532=>"000000001",
  40533=>"011110001",
  40534=>"000100010",
  40535=>"100011111",
  40536=>"000001101",
  40537=>"101100100",
  40538=>"111100111",
  40539=>"001011010",
  40540=>"000101110",
  40541=>"011010101",
  40542=>"111100001",
  40543=>"010101110",
  40544=>"110111010",
  40545=>"001101111",
  40546=>"100100010",
  40547=>"000010010",
  40548=>"101010110",
  40549=>"001000100",
  40550=>"101101111",
  40551=>"011010111",
  40552=>"110011001",
  40553=>"010010111",
  40554=>"100101110",
  40555=>"111011111",
  40556=>"110011001",
  40557=>"101011110",
  40558=>"001000010",
  40559=>"111001111",
  40560=>"011001111",
  40561=>"000100100",
  40562=>"000001010",
  40563=>"100011010",
  40564=>"011010101",
  40565=>"001100111",
  40566=>"110010001",
  40567=>"001000010",
  40568=>"000011010",
  40569=>"001101000",
  40570=>"011110101",
  40571=>"000011111",
  40572=>"010001001",
  40573=>"101000000",
  40574=>"100000101",
  40575=>"101011110",
  40576=>"000001100",
  40577=>"101011010",
  40578=>"111101111",
  40579=>"001001111",
  40580=>"001101111",
  40581=>"110110110",
  40582=>"100011111",
  40583=>"001010110",
  40584=>"100000001",
  40585=>"010100001",
  40586=>"011011001",
  40587=>"000111110",
  40588=>"100111111",
  40589=>"011000110",
  40590=>"010000010",
  40591=>"010000000",
  40592=>"001111110",
  40593=>"011101000",
  40594=>"011001100",
  40595=>"110110111",
  40596=>"111110000",
  40597=>"011011001",
  40598=>"101001000",
  40599=>"101010001",
  40600=>"000110111",
  40601=>"011010011",
  40602=>"101010000",
  40603=>"000111100",
  40604=>"110110001",
  40605=>"111011011",
  40606=>"001110001",
  40607=>"001100010",
  40608=>"000111100",
  40609=>"111011110",
  40610=>"001110100",
  40611=>"000110010",
  40612=>"100011110",
  40613=>"010110111",
  40614=>"110101100",
  40615=>"000000000",
  40616=>"001001000",
  40617=>"101011000",
  40618=>"000010110",
  40619=>"001001011",
  40620=>"000100101",
  40621=>"000001100",
  40622=>"010000111",
  40623=>"011111101",
  40624=>"000110001",
  40625=>"011111101",
  40626=>"000110110",
  40627=>"011011111",
  40628=>"010111010",
  40629=>"001010110",
  40630=>"101000110",
  40631=>"111111101",
  40632=>"110101000",
  40633=>"001111100",
  40634=>"010011001",
  40635=>"111011111",
  40636=>"100110010",
  40637=>"100101000",
  40638=>"111001000",
  40639=>"111001110",
  40640=>"110110111",
  40641=>"111001011",
  40642=>"111101110",
  40643=>"001111110",
  40644=>"011100101",
  40645=>"110011100",
  40646=>"100100100",
  40647=>"111100101",
  40648=>"001100000",
  40649=>"001001100",
  40650=>"101110101",
  40651=>"001001010",
  40652=>"101100011",
  40653=>"001010011",
  40654=>"110010101",
  40655=>"000010000",
  40656=>"010100110",
  40657=>"011100000",
  40658=>"100001110",
  40659=>"111111101",
  40660=>"100101100",
  40661=>"000011001",
  40662=>"111111011",
  40663=>"110000001",
  40664=>"101111010",
  40665=>"110011110",
  40666=>"010001000",
  40667=>"110000001",
  40668=>"001000111",
  40669=>"001111001",
  40670=>"000000101",
  40671=>"010110101",
  40672=>"011100101",
  40673=>"001100101",
  40674=>"011011011",
  40675=>"001001000",
  40676=>"000111010",
  40677=>"100111011",
  40678=>"110101010",
  40679=>"010001100",
  40680=>"111000000",
  40681=>"000101110",
  40682=>"001101011",
  40683=>"110111101",
  40684=>"100010011",
  40685=>"001010001",
  40686=>"110101111",
  40687=>"011000001",
  40688=>"111111111",
  40689=>"110011111",
  40690=>"101110011",
  40691=>"111111001",
  40692=>"010100111",
  40693=>"010111100",
  40694=>"011100111",
  40695=>"110011110",
  40696=>"000001001",
  40697=>"111011101",
  40698=>"010000110",
  40699=>"011000000",
  40700=>"010011111",
  40701=>"011100000",
  40702=>"011011000",
  40703=>"110100101",
  40704=>"111111111",
  40705=>"011000010",
  40706=>"101110001",
  40707=>"000011100",
  40708=>"010010010",
  40709=>"110110010",
  40710=>"000000000",
  40711=>"101110110",
  40712=>"101011111",
  40713=>"100110001",
  40714=>"100001111",
  40715=>"001011001",
  40716=>"101101101",
  40717=>"011000101",
  40718=>"100101000",
  40719=>"001001110",
  40720=>"111000000",
  40721=>"111011110",
  40722=>"000101110",
  40723=>"000110010",
  40724=>"101011101",
  40725=>"100010111",
  40726=>"100110111",
  40727=>"111001001",
  40728=>"000001000",
  40729=>"010100010",
  40730=>"010010001",
  40731=>"000010001",
  40732=>"111011001",
  40733=>"111101111",
  40734=>"111011011",
  40735=>"101100110",
  40736=>"001010111",
  40737=>"000110001",
  40738=>"001101000",
  40739=>"111101101",
  40740=>"010101000",
  40741=>"010111001",
  40742=>"110100001",
  40743=>"011111001",
  40744=>"100011101",
  40745=>"001111111",
  40746=>"011110110",
  40747=>"010001000",
  40748=>"011101010",
  40749=>"101000110",
  40750=>"101110110",
  40751=>"011010011",
  40752=>"100000011",
  40753=>"000100011",
  40754=>"000101001",
  40755=>"100001011",
  40756=>"010101011",
  40757=>"110000010",
  40758=>"011010101",
  40759=>"100100100",
  40760=>"000110010",
  40761=>"000101101",
  40762=>"011111001",
  40763=>"001100101",
  40764=>"101110101",
  40765=>"100000110",
  40766=>"100001010",
  40767=>"100110111",
  40768=>"110010010",
  40769=>"110110010",
  40770=>"100101010",
  40771=>"100011000",
  40772=>"111011001",
  40773=>"111010110",
  40774=>"111011101",
  40775=>"101100001",
  40776=>"100101000",
  40777=>"111010001",
  40778=>"110110011",
  40779=>"101010100",
  40780=>"111111010",
  40781=>"111010000",
  40782=>"111000111",
  40783=>"110010111",
  40784=>"011100000",
  40785=>"001010001",
  40786=>"001000001",
  40787=>"010000111",
  40788=>"010111100",
  40789=>"011011101",
  40790=>"111101011",
  40791=>"111010110",
  40792=>"111000100",
  40793=>"010010000",
  40794=>"011100101",
  40795=>"111001010",
  40796=>"010000100",
  40797=>"100000010",
  40798=>"001010001",
  40799=>"011010000",
  40800=>"001000100",
  40801=>"100110010",
  40802=>"110010000",
  40803=>"110110110",
  40804=>"000101110",
  40805=>"100001011",
  40806=>"110001001",
  40807=>"110010110",
  40808=>"010111111",
  40809=>"010000011",
  40810=>"001110110",
  40811=>"001010101",
  40812=>"010100111",
  40813=>"110000010",
  40814=>"001100011",
  40815=>"001001001",
  40816=>"110110000",
  40817=>"100110111",
  40818=>"110001000",
  40819=>"010100001",
  40820=>"100110011",
  40821=>"001010101",
  40822=>"011110011",
  40823=>"110001000",
  40824=>"101110111",
  40825=>"000101100",
  40826=>"101011101",
  40827=>"010100110",
  40828=>"110101100",
  40829=>"010111011",
  40830=>"110111100",
  40831=>"010000000",
  40832=>"110010101",
  40833=>"001010001",
  40834=>"000110001",
  40835=>"011101111",
  40836=>"100110000",
  40837=>"100001100",
  40838=>"001100011",
  40839=>"111110100",
  40840=>"010011100",
  40841=>"001100110",
  40842=>"001010000",
  40843=>"001001011",
  40844=>"001011110",
  40845=>"001110010",
  40846=>"101101010",
  40847=>"000001000",
  40848=>"011010001",
  40849=>"001001111",
  40850=>"101101011",
  40851=>"010111000",
  40852=>"000011110",
  40853=>"110110011",
  40854=>"100100010",
  40855=>"100011100",
  40856=>"110110101",
  40857=>"000000111",
  40858=>"111110110",
  40859=>"000010101",
  40860=>"111001111",
  40861=>"011110101",
  40862=>"111011000",
  40863=>"010001010",
  40864=>"011110010",
  40865=>"010001101",
  40866=>"010000101",
  40867=>"101100110",
  40868=>"001000101",
  40869=>"110001111",
  40870=>"110001110",
  40871=>"001001110",
  40872=>"000100111",
  40873=>"101011101",
  40874=>"011110011",
  40875=>"010000110",
  40876=>"111001010",
  40877=>"000010100",
  40878=>"100011011",
  40879=>"001011111",
  40880=>"111111011",
  40881=>"001100111",
  40882=>"111111001",
  40883=>"110101000",
  40884=>"001110111",
  40885=>"101011000",
  40886=>"101101011",
  40887=>"001001011",
  40888=>"100111011",
  40889=>"100000110",
  40890=>"010111101",
  40891=>"111001110",
  40892=>"000000010",
  40893=>"101111111",
  40894=>"101010001",
  40895=>"100101001",
  40896=>"000010000",
  40897=>"011110110",
  40898=>"011101101",
  40899=>"010110011",
  40900=>"011101101",
  40901=>"101100101",
  40902=>"010001000",
  40903=>"001011101",
  40904=>"111111110",
  40905=>"001000000",
  40906=>"111111100",
  40907=>"000010010",
  40908=>"111011111",
  40909=>"010111000",
  40910=>"101111111",
  40911=>"100101010",
  40912=>"100110100",
  40913=>"001101010",
  40914=>"101100111",
  40915=>"000100110",
  40916=>"100011001",
  40917=>"011010000",
  40918=>"010111110",
  40919=>"011000100",
  40920=>"111111100",
  40921=>"100010101",
  40922=>"010011000",
  40923=>"100000000",
  40924=>"111101011",
  40925=>"001010110",
  40926=>"010110000",
  40927=>"101110001",
  40928=>"010111111",
  40929=>"000000110",
  40930=>"010110100",
  40931=>"111000101",
  40932=>"111010000",
  40933=>"001101000",
  40934=>"111111000",
  40935=>"001010010",
  40936=>"111100101",
  40937=>"001110000",
  40938=>"111101000",
  40939=>"110011111",
  40940=>"100000000",
  40941=>"111010100",
  40942=>"111100000",
  40943=>"001111000",
  40944=>"101111010",
  40945=>"010101000",
  40946=>"100000100",
  40947=>"100010000",
  40948=>"100111001",
  40949=>"111100010",
  40950=>"011110100",
  40951=>"100011010",
  40952=>"100110111",
  40953=>"110000011",
  40954=>"100110010",
  40955=>"111110100",
  40956=>"111100011",
  40957=>"010000001",
  40958=>"100111110",
  40959=>"000011100",
  40960=>"001111000",
  40961=>"110000000",
  40962=>"011100101",
  40963=>"110001110",
  40964=>"001110110",
  40965=>"001111111",
  40966=>"010010010",
  40967=>"010100011",
  40968=>"011001110",
  40969=>"100000111",
  40970=>"001001111",
  40971=>"111101101",
  40972=>"101111100",
  40973=>"110100111",
  40974=>"010010011",
  40975=>"001011101",
  40976=>"010010000",
  40977=>"101111000",
  40978=>"100000001",
  40979=>"000000111",
  40980=>"100101111",
  40981=>"000001000",
  40982=>"110100101",
  40983=>"001110001",
  40984=>"001101011",
  40985=>"010000100",
  40986=>"011010011",
  40987=>"001011110",
  40988=>"110111000",
  40989=>"010101111",
  40990=>"111000111",
  40991=>"100100000",
  40992=>"100010000",
  40993=>"000011110",
  40994=>"101100001",
  40995=>"001001011",
  40996=>"011111111",
  40997=>"110111101",
  40998=>"100011111",
  40999=>"100000101",
  41000=>"111010000",
  41001=>"010101110",
  41002=>"110010111",
  41003=>"101101111",
  41004=>"011001100",
  41005=>"101001010",
  41006=>"011010000",
  41007=>"001101010",
  41008=>"000010111",
  41009=>"101110101",
  41010=>"100000011",
  41011=>"010001011",
  41012=>"001100011",
  41013=>"101000100",
  41014=>"000110010",
  41015=>"001010101",
  41016=>"010110100",
  41017=>"111010010",
  41018=>"100010111",
  41019=>"110011111",
  41020=>"101101100",
  41021=>"010110110",
  41022=>"001101100",
  41023=>"111101101",
  41024=>"100001010",
  41025=>"101100100",
  41026=>"001010010",
  41027=>"000100100",
  41028=>"111100101",
  41029=>"100000010",
  41030=>"001101111",
  41031=>"111001001",
  41032=>"110010001",
  41033=>"101111101",
  41034=>"001101101",
  41035=>"100011111",
  41036=>"100100000",
  41037=>"110011011",
  41038=>"111100011",
  41039=>"011110101",
  41040=>"011001101",
  41041=>"111100110",
  41042=>"101011000",
  41043=>"001010011",
  41044=>"110000000",
  41045=>"011100001",
  41046=>"100110101",
  41047=>"001011001",
  41048=>"111110001",
  41049=>"100011010",
  41050=>"000010010",
  41051=>"000010011",
  41052=>"101111111",
  41053=>"110101011",
  41054=>"100001101",
  41055=>"111001000",
  41056=>"000110010",
  41057=>"111011111",
  41058=>"101000111",
  41059=>"010010010",
  41060=>"101011011",
  41061=>"110000101",
  41062=>"100111101",
  41063=>"000101000",
  41064=>"010101111",
  41065=>"100001000",
  41066=>"000010100",
  41067=>"011100111",
  41068=>"010001111",
  41069=>"001101101",
  41070=>"110000110",
  41071=>"110111000",
  41072=>"001001011",
  41073=>"010110001",
  41074=>"000101000",
  41075=>"101100101",
  41076=>"011000110",
  41077=>"100010111",
  41078=>"111000000",
  41079=>"010100000",
  41080=>"000010100",
  41081=>"101000111",
  41082=>"110111010",
  41083=>"111111101",
  41084=>"000011100",
  41085=>"010111111",
  41086=>"100101111",
  41087=>"000100110",
  41088=>"100100001",
  41089=>"111110000",
  41090=>"011010000",
  41091=>"100111110",
  41092=>"111111110",
  41093=>"111010000",
  41094=>"001111011",
  41095=>"111011111",
  41096=>"010000110",
  41097=>"010000110",
  41098=>"100011010",
  41099=>"111010001",
  41100=>"010010000",
  41101=>"100010001",
  41102=>"111101100",
  41103=>"110100010",
  41104=>"000001011",
  41105=>"001010101",
  41106=>"000100111",
  41107=>"110011101",
  41108=>"001110111",
  41109=>"110100010",
  41110=>"011110110",
  41111=>"000001000",
  41112=>"010100000",
  41113=>"100001011",
  41114=>"010100001",
  41115=>"100011110",
  41116=>"010100100",
  41117=>"101010000",
  41118=>"011100011",
  41119=>"100110011",
  41120=>"000001000",
  41121=>"110011010",
  41122=>"010010010",
  41123=>"011100000",
  41124=>"011110100",
  41125=>"110100110",
  41126=>"011101100",
  41127=>"111010110",
  41128=>"011100100",
  41129=>"000010001",
  41130=>"110011111",
  41131=>"010111101",
  41132=>"001100100",
  41133=>"010010011",
  41134=>"011110110",
  41135=>"001000000",
  41136=>"011101101",
  41137=>"111110000",
  41138=>"100001100",
  41139=>"110111000",
  41140=>"101100000",
  41141=>"110111111",
  41142=>"000000110",
  41143=>"010100001",
  41144=>"001000111",
  41145=>"000000111",
  41146=>"100100011",
  41147=>"100111101",
  41148=>"001011011",
  41149=>"101000010",
  41150=>"000010011",
  41151=>"001011110",
  41152=>"000011011",
  41153=>"010100100",
  41154=>"111100001",
  41155=>"001111111",
  41156=>"010101000",
  41157=>"101010011",
  41158=>"101011010",
  41159=>"101011111",
  41160=>"100101000",
  41161=>"110000011",
  41162=>"010101010",
  41163=>"101011111",
  41164=>"010011010",
  41165=>"100001100",
  41166=>"001010100",
  41167=>"111011001",
  41168=>"111001111",
  41169=>"011000000",
  41170=>"110100100",
  41171=>"100010001",
  41172=>"010111100",
  41173=>"010000000",
  41174=>"001111001",
  41175=>"110011101",
  41176=>"110111000",
  41177=>"101011111",
  41178=>"111111110",
  41179=>"111100101",
  41180=>"011101001",
  41181=>"000110111",
  41182=>"111100010",
  41183=>"011010100",
  41184=>"111010010",
  41185=>"001010001",
  41186=>"111000000",
  41187=>"011111101",
  41188=>"100101101",
  41189=>"010111111",
  41190=>"010000101",
  41191=>"101101001",
  41192=>"011110111",
  41193=>"101100111",
  41194=>"010110100",
  41195=>"000110000",
  41196=>"110101010",
  41197=>"110111110",
  41198=>"001100001",
  41199=>"110001111",
  41200=>"011010010",
  41201=>"010011110",
  41202=>"010101001",
  41203=>"111111000",
  41204=>"110011101",
  41205=>"000000110",
  41206=>"111110000",
  41207=>"101001010",
  41208=>"100001111",
  41209=>"111101010",
  41210=>"110101111",
  41211=>"011011100",
  41212=>"111011011",
  41213=>"111011010",
  41214=>"001001000",
  41215=>"010000010",
  41216=>"111111000",
  41217=>"111100000",
  41218=>"110011010",
  41219=>"111111100",
  41220=>"001101011",
  41221=>"101111111",
  41222=>"110110001",
  41223=>"001110001",
  41224=>"110001001",
  41225=>"100111011",
  41226=>"000100110",
  41227=>"111000110",
  41228=>"001001001",
  41229=>"000110100",
  41230=>"010111100",
  41231=>"011011011",
  41232=>"001101111",
  41233=>"110000010",
  41234=>"010011001",
  41235=>"011111001",
  41236=>"011011101",
  41237=>"110110011",
  41238=>"010111010",
  41239=>"110101001",
  41240=>"111011110",
  41241=>"011111111",
  41242=>"010111100",
  41243=>"101001111",
  41244=>"100100100",
  41245=>"001111000",
  41246=>"000011111",
  41247=>"111111010",
  41248=>"000011110",
  41249=>"010110000",
  41250=>"011111000",
  41251=>"110011110",
  41252=>"110001111",
  41253=>"101101000",
  41254=>"111110111",
  41255=>"111110111",
  41256=>"000000011",
  41257=>"111000110",
  41258=>"111100101",
  41259=>"001110000",
  41260=>"100011101",
  41261=>"111011010",
  41262=>"111110011",
  41263=>"011010011",
  41264=>"011011101",
  41265=>"100111100",
  41266=>"001011011",
  41267=>"001001010",
  41268=>"101000111",
  41269=>"010100101",
  41270=>"100001101",
  41271=>"011000010",
  41272=>"000000000",
  41273=>"001011100",
  41274=>"011000101",
  41275=>"111111011",
  41276=>"011001100",
  41277=>"100100100",
  41278=>"000001000",
  41279=>"101110011",
  41280=>"100000101",
  41281=>"010100111",
  41282=>"111011010",
  41283=>"011000010",
  41284=>"110010011",
  41285=>"110001001",
  41286=>"110000101",
  41287=>"011000100",
  41288=>"111111101",
  41289=>"100000001",
  41290=>"111000110",
  41291=>"101101111",
  41292=>"010001000",
  41293=>"111101110",
  41294=>"110000001",
  41295=>"001100100",
  41296=>"111101001",
  41297=>"011000001",
  41298=>"100110011",
  41299=>"101001110",
  41300=>"110011000",
  41301=>"010011001",
  41302=>"010001010",
  41303=>"111111000",
  41304=>"101010100",
  41305=>"001011011",
  41306=>"010011011",
  41307=>"110011011",
  41308=>"100011100",
  41309=>"010010101",
  41310=>"011001000",
  41311=>"110001000",
  41312=>"000100100",
  41313=>"000111010",
  41314=>"101011101",
  41315=>"111011110",
  41316=>"111111000",
  41317=>"000001001",
  41318=>"011010000",
  41319=>"111011011",
  41320=>"110110001",
  41321=>"000000001",
  41322=>"001001001",
  41323=>"100101101",
  41324=>"111111101",
  41325=>"000001101",
  41326=>"010001101",
  41327=>"010111111",
  41328=>"001111001",
  41329=>"011001010",
  41330=>"000111011",
  41331=>"100101001",
  41332=>"111001100",
  41333=>"010111011",
  41334=>"000001011",
  41335=>"100111010",
  41336=>"011101101",
  41337=>"101101011",
  41338=>"111110100",
  41339=>"111110000",
  41340=>"010011001",
  41341=>"000000001",
  41342=>"101111100",
  41343=>"110000101",
  41344=>"111001100",
  41345=>"111110101",
  41346=>"110011100",
  41347=>"110100100",
  41348=>"110101011",
  41349=>"001011101",
  41350=>"011000100",
  41351=>"111110000",
  41352=>"111110001",
  41353=>"010011100",
  41354=>"011110001",
  41355=>"010010010",
  41356=>"000111111",
  41357=>"101001010",
  41358=>"010001011",
  41359=>"100010101",
  41360=>"010011110",
  41361=>"111011000",
  41362=>"001101000",
  41363=>"100001101",
  41364=>"100101101",
  41365=>"101000001",
  41366=>"000010101",
  41367=>"001000110",
  41368=>"100001010",
  41369=>"100001010",
  41370=>"101010010",
  41371=>"011100011",
  41372=>"111011100",
  41373=>"011101111",
  41374=>"111010111",
  41375=>"010010111",
  41376=>"111101001",
  41377=>"011111010",
  41378=>"111101100",
  41379=>"111101001",
  41380=>"001001111",
  41381=>"101110101",
  41382=>"001001010",
  41383=>"100000001",
  41384=>"001110011",
  41385=>"111000010",
  41386=>"011010100",
  41387=>"111110010",
  41388=>"001101110",
  41389=>"111011100",
  41390=>"110000001",
  41391=>"011110000",
  41392=>"001010100",
  41393=>"010110000",
  41394=>"000001010",
  41395=>"001101001",
  41396=>"001111111",
  41397=>"011000100",
  41398=>"010110000",
  41399=>"011001011",
  41400=>"110101001",
  41401=>"100001101",
  41402=>"110011001",
  41403=>"100101110",
  41404=>"100101111",
  41405=>"111111101",
  41406=>"101001111",
  41407=>"011011101",
  41408=>"100110000",
  41409=>"000110010",
  41410=>"000011100",
  41411=>"101110100",
  41412=>"111011011",
  41413=>"000101000",
  41414=>"000010000",
  41415=>"110110100",
  41416=>"001011010",
  41417=>"110001011",
  41418=>"111101111",
  41419=>"101100101",
  41420=>"111110011",
  41421=>"111111011",
  41422=>"000011011",
  41423=>"011000111",
  41424=>"100100010",
  41425=>"101011011",
  41426=>"011100100",
  41427=>"000010010",
  41428=>"111101100",
  41429=>"110001000",
  41430=>"011101101",
  41431=>"110111100",
  41432=>"001111101",
  41433=>"101011001",
  41434=>"010111000",
  41435=>"001010011",
  41436=>"100100100",
  41437=>"010001010",
  41438=>"111001100",
  41439=>"001101010",
  41440=>"000010100",
  41441=>"010100100",
  41442=>"000101001",
  41443=>"001010101",
  41444=>"111101011",
  41445=>"001011001",
  41446=>"010110101",
  41447=>"101011011",
  41448=>"111110000",
  41449=>"101111010",
  41450=>"000010000",
  41451=>"110110110",
  41452=>"000100101",
  41453=>"100001111",
  41454=>"111011100",
  41455=>"111111000",
  41456=>"000001000",
  41457=>"111010001",
  41458=>"101000111",
  41459=>"101001000",
  41460=>"110110101",
  41461=>"100000111",
  41462=>"111111000",
  41463=>"010010110",
  41464=>"101100110",
  41465=>"010011100",
  41466=>"111110010",
  41467=>"100101101",
  41468=>"000010011",
  41469=>"101000111",
  41470=>"001111110",
  41471=>"011111011",
  41472=>"000001000",
  41473=>"010000111",
  41474=>"101101001",
  41475=>"101101010",
  41476=>"110110110",
  41477=>"001101010",
  41478=>"100110011",
  41479=>"010011101",
  41480=>"100000000",
  41481=>"011011101",
  41482=>"100111110",
  41483=>"000001110",
  41484=>"100110111",
  41485=>"101000011",
  41486=>"111000101",
  41487=>"100110111",
  41488=>"101100001",
  41489=>"001110010",
  41490=>"101011101",
  41491=>"111110100",
  41492=>"011110010",
  41493=>"001110000",
  41494=>"010010110",
  41495=>"001000010",
  41496=>"110100110",
  41497=>"101110011",
  41498=>"110110100",
  41499=>"101001011",
  41500=>"101001100",
  41501=>"101000011",
  41502=>"000101111",
  41503=>"000011101",
  41504=>"011100010",
  41505=>"101010111",
  41506=>"000011011",
  41507=>"111001011",
  41508=>"010011001",
  41509=>"010010100",
  41510=>"010001101",
  41511=>"010010011",
  41512=>"101000110",
  41513=>"111100101",
  41514=>"100010111",
  41515=>"101001000",
  41516=>"010110111",
  41517=>"010101010",
  41518=>"000110000",
  41519=>"001111000",
  41520=>"100101100",
  41521=>"011111101",
  41522=>"110011101",
  41523=>"001111001",
  41524=>"110100110",
  41525=>"111101100",
  41526=>"101010110",
  41527=>"010010010",
  41528=>"101010011",
  41529=>"101100100",
  41530=>"101101111",
  41531=>"010011001",
  41532=>"001100100",
  41533=>"111001110",
  41534=>"111001101",
  41535=>"101100100",
  41536=>"000001000",
  41537=>"100011000",
  41538=>"110011010",
  41539=>"001000010",
  41540=>"001001000",
  41541=>"001001110",
  41542=>"011000001",
  41543=>"101101001",
  41544=>"101010010",
  41545=>"110110011",
  41546=>"100010110",
  41547=>"001100111",
  41548=>"011100011",
  41549=>"000111010",
  41550=>"011110010",
  41551=>"011101111",
  41552=>"010000100",
  41553=>"001000010",
  41554=>"010111011",
  41555=>"101001000",
  41556=>"100101110",
  41557=>"010000010",
  41558=>"111010010",
  41559=>"101100011",
  41560=>"010010101",
  41561=>"110000111",
  41562=>"101011010",
  41563=>"000111010",
  41564=>"101011000",
  41565=>"100111000",
  41566=>"001000001",
  41567=>"100001000",
  41568=>"010110100",
  41569=>"100100111",
  41570=>"011110100",
  41571=>"000000011",
  41572=>"101110011",
  41573=>"110011000",
  41574=>"101111000",
  41575=>"111101101",
  41576=>"101010000",
  41577=>"111001111",
  41578=>"001011001",
  41579=>"000111000",
  41580=>"110101011",
  41581=>"100010000",
  41582=>"101001100",
  41583=>"111101111",
  41584=>"000100011",
  41585=>"001111000",
  41586=>"000111111",
  41587=>"101000000",
  41588=>"011001101",
  41589=>"111000011",
  41590=>"110101100",
  41591=>"101111100",
  41592=>"110110010",
  41593=>"010010110",
  41594=>"100001101",
  41595=>"001110010",
  41596=>"111100010",
  41597=>"010011011",
  41598=>"110000010",
  41599=>"111111010",
  41600=>"111001000",
  41601=>"001000011",
  41602=>"011101110",
  41603=>"010000001",
  41604=>"110000001",
  41605=>"110110111",
  41606=>"111111011",
  41607=>"100111101",
  41608=>"001011101",
  41609=>"110001100",
  41610=>"100110010",
  41611=>"110011110",
  41612=>"110110101",
  41613=>"111010110",
  41614=>"111110111",
  41615=>"000000001",
  41616=>"001001101",
  41617=>"001000110",
  41618=>"110001101",
  41619=>"110101101",
  41620=>"100000001",
  41621=>"000110100",
  41622=>"111111011",
  41623=>"010101110",
  41624=>"100010100",
  41625=>"000010010",
  41626=>"111011011",
  41627=>"111101110",
  41628=>"100101000",
  41629=>"110101111",
  41630=>"010111101",
  41631=>"010000111",
  41632=>"000111110",
  41633=>"101001001",
  41634=>"011000001",
  41635=>"101001101",
  41636=>"100110111",
  41637=>"101001001",
  41638=>"110011100",
  41639=>"110011000",
  41640=>"010010110",
  41641=>"111111110",
  41642=>"000100100",
  41643=>"001101101",
  41644=>"011111000",
  41645=>"011000111",
  41646=>"110010011",
  41647=>"111111000",
  41648=>"100000010",
  41649=>"101001011",
  41650=>"110001000",
  41651=>"001000100",
  41652=>"101010101",
  41653=>"010101100",
  41654=>"101100111",
  41655=>"101000000",
  41656=>"001110001",
  41657=>"100001100",
  41658=>"110000011",
  41659=>"111101101",
  41660=>"101001100",
  41661=>"101001001",
  41662=>"111010100",
  41663=>"111011111",
  41664=>"110010010",
  41665=>"110011110",
  41666=>"101011110",
  41667=>"110001010",
  41668=>"100000101",
  41669=>"101100101",
  41670=>"111000001",
  41671=>"010110101",
  41672=>"110101111",
  41673=>"000000101",
  41674=>"000010101",
  41675=>"101010000",
  41676=>"010100101",
  41677=>"100111101",
  41678=>"011110110",
  41679=>"101010010",
  41680=>"101001011",
  41681=>"011110110",
  41682=>"100100000",
  41683=>"010000011",
  41684=>"010110110",
  41685=>"001010010",
  41686=>"111111101",
  41687=>"000001101",
  41688=>"011011011",
  41689=>"000110001",
  41690=>"000100001",
  41691=>"001100010",
  41692=>"011001101",
  41693=>"101001100",
  41694=>"101100101",
  41695=>"111010101",
  41696=>"111101111",
  41697=>"000000010",
  41698=>"100000101",
  41699=>"001110001",
  41700=>"000010011",
  41701=>"000110001",
  41702=>"011011111",
  41703=>"111010011",
  41704=>"101001011",
  41705=>"101000100",
  41706=>"001011111",
  41707=>"101101011",
  41708=>"011010100",
  41709=>"000111110",
  41710=>"001000100",
  41711=>"011011011",
  41712=>"011001110",
  41713=>"000011110",
  41714=>"010111001",
  41715=>"000110100",
  41716=>"110110110",
  41717=>"011000110",
  41718=>"010001100",
  41719=>"100010101",
  41720=>"111111101",
  41721=>"000000001",
  41722=>"001001100",
  41723=>"111110110",
  41724=>"001011110",
  41725=>"100111011",
  41726=>"110110001",
  41727=>"010001000",
  41728=>"101110001",
  41729=>"110001100",
  41730=>"000100001",
  41731=>"101100110",
  41732=>"011110000",
  41733=>"100000001",
  41734=>"000100110",
  41735=>"010110001",
  41736=>"010000000",
  41737=>"000101101",
  41738=>"101000000",
  41739=>"110011110",
  41740=>"101011100",
  41741=>"000010011",
  41742=>"101011001",
  41743=>"100100100",
  41744=>"101110001",
  41745=>"100011011",
  41746=>"011110011",
  41747=>"101010011",
  41748=>"001010101",
  41749=>"100000000",
  41750=>"111000000",
  41751=>"110000110",
  41752=>"001111001",
  41753=>"101000001",
  41754=>"001101101",
  41755=>"010000001",
  41756=>"001000000",
  41757=>"001111111",
  41758=>"000011001",
  41759=>"111010001",
  41760=>"100010000",
  41761=>"101000001",
  41762=>"010001111",
  41763=>"000101001",
  41764=>"110100111",
  41765=>"100000101",
  41766=>"101111110",
  41767=>"111000111",
  41768=>"001101010",
  41769=>"001110001",
  41770=>"111010011",
  41771=>"111110010",
  41772=>"101010110",
  41773=>"000110111",
  41774=>"101001010",
  41775=>"110011111",
  41776=>"000010010",
  41777=>"110111101",
  41778=>"000001100",
  41779=>"000100000",
  41780=>"011111000",
  41781=>"110110101",
  41782=>"111110010",
  41783=>"101011100",
  41784=>"111110000",
  41785=>"000000011",
  41786=>"001110011",
  41787=>"110001100",
  41788=>"001001000",
  41789=>"001111011",
  41790=>"101000011",
  41791=>"001001000",
  41792=>"010101010",
  41793=>"110000110",
  41794=>"111111101",
  41795=>"010001101",
  41796=>"010000000",
  41797=>"101010110",
  41798=>"000010000",
  41799=>"010000111",
  41800=>"100010110",
  41801=>"111100111",
  41802=>"000011110",
  41803=>"101101101",
  41804=>"001010001",
  41805=>"000001001",
  41806=>"001001111",
  41807=>"100010010",
  41808=>"110001100",
  41809=>"111001011",
  41810=>"011000111",
  41811=>"010000100",
  41812=>"111100001",
  41813=>"110101000",
  41814=>"001101011",
  41815=>"111000111",
  41816=>"110001100",
  41817=>"101001001",
  41818=>"100100100",
  41819=>"011011100",
  41820=>"100100001",
  41821=>"101000010",
  41822=>"001011000",
  41823=>"101101100",
  41824=>"011000110",
  41825=>"010011101",
  41826=>"000010010",
  41827=>"010011111",
  41828=>"011000100",
  41829=>"000100000",
  41830=>"001111001",
  41831=>"100100101",
  41832=>"100001001",
  41833=>"111100001",
  41834=>"101001111",
  41835=>"110010111",
  41836=>"111101110",
  41837=>"100000010",
  41838=>"110101100",
  41839=>"011110110",
  41840=>"010010001",
  41841=>"001100010",
  41842=>"111011110",
  41843=>"101011000",
  41844=>"100001101",
  41845=>"001000000",
  41846=>"010110110",
  41847=>"000111000",
  41848=>"000000111",
  41849=>"001100111",
  41850=>"001011111",
  41851=>"001001100",
  41852=>"001010000",
  41853=>"111101001",
  41854=>"111101010",
  41855=>"001011000",
  41856=>"001001111",
  41857=>"100000101",
  41858=>"000111000",
  41859=>"000110010",
  41860=>"100100001",
  41861=>"001100010",
  41862=>"100100110",
  41863=>"000001111",
  41864=>"010001111",
  41865=>"001010010",
  41866=>"001110000",
  41867=>"101111111",
  41868=>"110001000",
  41869=>"111100100",
  41870=>"111000111",
  41871=>"111101001",
  41872=>"101110101",
  41873=>"000011001",
  41874=>"111011000",
  41875=>"000010111",
  41876=>"110010000",
  41877=>"000100100",
  41878=>"010111011",
  41879=>"110001101",
  41880=>"010011111",
  41881=>"010001111",
  41882=>"010001111",
  41883=>"000000010",
  41884=>"110111100",
  41885=>"111011101",
  41886=>"000000101",
  41887=>"010110100",
  41888=>"100100100",
  41889=>"101111100",
  41890=>"001011100",
  41891=>"000001110",
  41892=>"011001010",
  41893=>"011000001",
  41894=>"111111101",
  41895=>"111100011",
  41896=>"110100000",
  41897=>"011000001",
  41898=>"101111101",
  41899=>"000000000",
  41900=>"101100101",
  41901=>"100000000",
  41902=>"100100011",
  41903=>"001000100",
  41904=>"010001110",
  41905=>"100100011",
  41906=>"010111001",
  41907=>"001110011",
  41908=>"111101010",
  41909=>"011001111",
  41910=>"001010101",
  41911=>"011001101",
  41912=>"101101001",
  41913=>"001100101",
  41914=>"000011111",
  41915=>"101101001",
  41916=>"110111011",
  41917=>"010000000",
  41918=>"101010110",
  41919=>"100000010",
  41920=>"101111111",
  41921=>"111110111",
  41922=>"101000011",
  41923=>"101101110",
  41924=>"000011000",
  41925=>"001101101",
  41926=>"001011001",
  41927=>"010000101",
  41928=>"010010010",
  41929=>"111100101",
  41930=>"111011000",
  41931=>"001010000",
  41932=>"111011011",
  41933=>"001000101",
  41934=>"101100000",
  41935=>"011000011",
  41936=>"111110111",
  41937=>"001101110",
  41938=>"111001111",
  41939=>"001110000",
  41940=>"001000100",
  41941=>"100000100",
  41942=>"000000000",
  41943=>"001110011",
  41944=>"110111011",
  41945=>"010101111",
  41946=>"010101111",
  41947=>"110100000",
  41948=>"111011011",
  41949=>"110110011",
  41950=>"100100010",
  41951=>"110111101",
  41952=>"000100100",
  41953=>"101001011",
  41954=>"010110110",
  41955=>"100000101",
  41956=>"111101011",
  41957=>"100100000",
  41958=>"001111100",
  41959=>"010110101",
  41960=>"001001100",
  41961=>"001111011",
  41962=>"110000111",
  41963=>"100011010",
  41964=>"010011100",
  41965=>"101001101",
  41966=>"011000101",
  41967=>"000001111",
  41968=>"001101101",
  41969=>"000001010",
  41970=>"010101001",
  41971=>"100000100",
  41972=>"110100111",
  41973=>"110010110",
  41974=>"000000110",
  41975=>"111100001",
  41976=>"111010010",
  41977=>"101111011",
  41978=>"111010111",
  41979=>"011010110",
  41980=>"000000010",
  41981=>"100111100",
  41982=>"011011000",
  41983=>"110011001",
  41984=>"111001011",
  41985=>"001001011",
  41986=>"111010010",
  41987=>"001010110",
  41988=>"100001001",
  41989=>"110100010",
  41990=>"111001101",
  41991=>"101011010",
  41992=>"001100010",
  41993=>"100100100",
  41994=>"111011110",
  41995=>"101110010",
  41996=>"000111111",
  41997=>"101011111",
  41998=>"000001110",
  41999=>"010100101",
  42000=>"010010000",
  42001=>"111110111",
  42002=>"111111111",
  42003=>"001011110",
  42004=>"010111000",
  42005=>"101001111",
  42006=>"111100011",
  42007=>"111011111",
  42008=>"011001111",
  42009=>"000100011",
  42010=>"101100000",
  42011=>"000000001",
  42012=>"000101011",
  42013=>"101100010",
  42014=>"000101010",
  42015=>"010010011",
  42016=>"001000010",
  42017=>"001011101",
  42018=>"001011000",
  42019=>"110111001",
  42020=>"111011011",
  42021=>"101111011",
  42022=>"111011101",
  42023=>"111100001",
  42024=>"011110001",
  42025=>"010110101",
  42026=>"110001010",
  42027=>"001001111",
  42028=>"111011110",
  42029=>"000100010",
  42030=>"011101000",
  42031=>"001101011",
  42032=>"101000000",
  42033=>"110110100",
  42034=>"011111101",
  42035=>"110001010",
  42036=>"010001101",
  42037=>"110001101",
  42038=>"011001010",
  42039=>"010010111",
  42040=>"001111010",
  42041=>"100010100",
  42042=>"110000001",
  42043=>"010000100",
  42044=>"000111000",
  42045=>"101100011",
  42046=>"010000000",
  42047=>"000111111",
  42048=>"110000100",
  42049=>"000000010",
  42050=>"101011110",
  42051=>"111011000",
  42052=>"100101100",
  42053=>"010100000",
  42054=>"101011010",
  42055=>"101111011",
  42056=>"100000101",
  42057=>"101000001",
  42058=>"011101001",
  42059=>"111111011",
  42060=>"001100111",
  42061=>"111110011",
  42062=>"011010001",
  42063=>"111011101",
  42064=>"111000000",
  42065=>"000011111",
  42066=>"011100001",
  42067=>"101101110",
  42068=>"111000010",
  42069=>"010101111",
  42070=>"100010111",
  42071=>"100001100",
  42072=>"010001100",
  42073=>"011010010",
  42074=>"111000100",
  42075=>"000000110",
  42076=>"000100110",
  42077=>"000011101",
  42078=>"000110111",
  42079=>"110001100",
  42080=>"011001100",
  42081=>"001000000",
  42082=>"111101010",
  42083=>"100101000",
  42084=>"111111111",
  42085=>"110000101",
  42086=>"110100100",
  42087=>"100100111",
  42088=>"011101000",
  42089=>"110011111",
  42090=>"001000000",
  42091=>"111000001",
  42092=>"110111011",
  42093=>"110111111",
  42094=>"001111001",
  42095=>"100001100",
  42096=>"110101100",
  42097=>"011001101",
  42098=>"111000111",
  42099=>"011000001",
  42100=>"101111101",
  42101=>"001110100",
  42102=>"111101011",
  42103=>"100000011",
  42104=>"100000000",
  42105=>"101101111",
  42106=>"111011011",
  42107=>"101011000",
  42108=>"100101011",
  42109=>"010110010",
  42110=>"100110101",
  42111=>"011000100",
  42112=>"011000100",
  42113=>"001000110",
  42114=>"000000000",
  42115=>"101011101",
  42116=>"011000001",
  42117=>"101111110",
  42118=>"001110101",
  42119=>"001001010",
  42120=>"101011100",
  42121=>"100000100",
  42122=>"111101110",
  42123=>"111011111",
  42124=>"110011000",
  42125=>"110100010",
  42126=>"101100011",
  42127=>"011010010",
  42128=>"101000110",
  42129=>"110000101",
  42130=>"001011110",
  42131=>"010011001",
  42132=>"000100101",
  42133=>"011100101",
  42134=>"101101010",
  42135=>"110100011",
  42136=>"001101000",
  42137=>"100110001",
  42138=>"110110010",
  42139=>"111011010",
  42140=>"110100011",
  42141=>"010010001",
  42142=>"100111010",
  42143=>"010110111",
  42144=>"011000001",
  42145=>"011010001",
  42146=>"110000110",
  42147=>"011111010",
  42148=>"100110010",
  42149=>"100011111",
  42150=>"011010010",
  42151=>"000001100",
  42152=>"010110001",
  42153=>"101111100",
  42154=>"110011101",
  42155=>"011000010",
  42156=>"110110101",
  42157=>"011010101",
  42158=>"011111100",
  42159=>"011001101",
  42160=>"100011001",
  42161=>"011000010",
  42162=>"011111111",
  42163=>"111000000",
  42164=>"000110100",
  42165=>"110101110",
  42166=>"011100111",
  42167=>"010011111",
  42168=>"010101001",
  42169=>"110010111",
  42170=>"100000100",
  42171=>"101111101",
  42172=>"001001000",
  42173=>"100110111",
  42174=>"010010010",
  42175=>"111111111",
  42176=>"001101111",
  42177=>"011110111",
  42178=>"011010101",
  42179=>"001110000",
  42180=>"010101011",
  42181=>"110001010",
  42182=>"110011110",
  42183=>"110100010",
  42184=>"100011000",
  42185=>"100111111",
  42186=>"010110101",
  42187=>"100001011",
  42188=>"011100111",
  42189=>"111000010",
  42190=>"000101101",
  42191=>"110101100",
  42192=>"110111111",
  42193=>"100111001",
  42194=>"000111011",
  42195=>"011101101",
  42196=>"011001101",
  42197=>"011010001",
  42198=>"011100010",
  42199=>"001111011",
  42200=>"001110010",
  42201=>"111111010",
  42202=>"011110011",
  42203=>"010101111",
  42204=>"111101100",
  42205=>"111111011",
  42206=>"110000100",
  42207=>"010111100",
  42208=>"010011001",
  42209=>"010101000",
  42210=>"101001001",
  42211=>"001000010",
  42212=>"001101011",
  42213=>"000111011",
  42214=>"101000001",
  42215=>"111011110",
  42216=>"100110101",
  42217=>"001110101",
  42218=>"011001111",
  42219=>"101111100",
  42220=>"010011110",
  42221=>"010111110",
  42222=>"000100101",
  42223=>"110100100",
  42224=>"000001100",
  42225=>"110010001",
  42226=>"001101000",
  42227=>"010000111",
  42228=>"001000000",
  42229=>"111111110",
  42230=>"111110101",
  42231=>"010100101",
  42232=>"000000100",
  42233=>"111001100",
  42234=>"010001000",
  42235=>"011110000",
  42236=>"000010010",
  42237=>"110000001",
  42238=>"011011111",
  42239=>"100000010",
  42240=>"100011111",
  42241=>"011011011",
  42242=>"110000101",
  42243=>"011001100",
  42244=>"000011110",
  42245=>"101001100",
  42246=>"010110001",
  42247=>"110100001",
  42248=>"001011101",
  42249=>"110110011",
  42250=>"010100100",
  42251=>"001001111",
  42252=>"111101001",
  42253=>"000011011",
  42254=>"001100010",
  42255=>"000000000",
  42256=>"100100100",
  42257=>"110101110",
  42258=>"101110111",
  42259=>"101001110",
  42260=>"010000010",
  42261=>"001000010",
  42262=>"101000101",
  42263=>"111110101",
  42264=>"111011000",
  42265=>"001111011",
  42266=>"100000000",
  42267=>"010001101",
  42268=>"111111101",
  42269=>"110111001",
  42270=>"101100101",
  42271=>"101011111",
  42272=>"101011100",
  42273=>"110000010",
  42274=>"101101101",
  42275=>"101000011",
  42276=>"110100101",
  42277=>"000101111",
  42278=>"110110101",
  42279=>"100101101",
  42280=>"000101001",
  42281=>"001111011",
  42282=>"100111011",
  42283=>"101001100",
  42284=>"111111011",
  42285=>"100011111",
  42286=>"111000000",
  42287=>"011100011",
  42288=>"010111011",
  42289=>"000000010",
  42290=>"001110000",
  42291=>"010000001",
  42292=>"111100110",
  42293=>"110111110",
  42294=>"001111011",
  42295=>"011010101",
  42296=>"011011011",
  42297=>"010100101",
  42298=>"000100000",
  42299=>"000000011",
  42300=>"111001101",
  42301=>"011111100",
  42302=>"111001000",
  42303=>"011101011",
  42304=>"010101100",
  42305=>"011010011",
  42306=>"000100001",
  42307=>"010011011",
  42308=>"111011001",
  42309=>"100000011",
  42310=>"000101001",
  42311=>"000101101",
  42312=>"101010101",
  42313=>"011011011",
  42314=>"000011111",
  42315=>"110100011",
  42316=>"111000110",
  42317=>"100011101",
  42318=>"000011000",
  42319=>"110001010",
  42320=>"111000011",
  42321=>"111011011",
  42322=>"000111100",
  42323=>"100001100",
  42324=>"101100000",
  42325=>"001001001",
  42326=>"000110100",
  42327=>"011111110",
  42328=>"101011110",
  42329=>"110101011",
  42330=>"011101101",
  42331=>"010010011",
  42332=>"010010010",
  42333=>"110011001",
  42334=>"100111111",
  42335=>"111010100",
  42336=>"101101101",
  42337=>"010010001",
  42338=>"000010100",
  42339=>"011000010",
  42340=>"101011000",
  42341=>"011101111",
  42342=>"000111010",
  42343=>"011110101",
  42344=>"110011110",
  42345=>"111110111",
  42346=>"100010111",
  42347=>"010001001",
  42348=>"001010001",
  42349=>"010111101",
  42350=>"000100110",
  42351=>"011000011",
  42352=>"010010011",
  42353=>"010111000",
  42354=>"110000110",
  42355=>"111110010",
  42356=>"100001000",
  42357=>"011110110",
  42358=>"101100010",
  42359=>"101000011",
  42360=>"110111100",
  42361=>"110101101",
  42362=>"011011010",
  42363=>"011110000",
  42364=>"100010111",
  42365=>"011111111",
  42366=>"111100001",
  42367=>"100001000",
  42368=>"110010010",
  42369=>"100111000",
  42370=>"010010111",
  42371=>"101010000",
  42372=>"110101101",
  42373=>"100110001",
  42374=>"011011101",
  42375=>"000011010",
  42376=>"011011111",
  42377=>"110110001",
  42378=>"001000110",
  42379=>"000001010",
  42380=>"001011001",
  42381=>"000000000",
  42382=>"111110010",
  42383=>"111000001",
  42384=>"100111001",
  42385=>"110000001",
  42386=>"110000110",
  42387=>"010100001",
  42388=>"101110101",
  42389=>"010111011",
  42390=>"110110110",
  42391=>"110110110",
  42392=>"100110100",
  42393=>"010111011",
  42394=>"010110000",
  42395=>"111100001",
  42396=>"110011001",
  42397=>"111100010",
  42398=>"001010010",
  42399=>"000001000",
  42400=>"011011111",
  42401=>"010000010",
  42402=>"001000000",
  42403=>"111000001",
  42404=>"110000011",
  42405=>"111101000",
  42406=>"101001011",
  42407=>"010000100",
  42408=>"011100100",
  42409=>"111111100",
  42410=>"000100111",
  42411=>"110011110",
  42412=>"000100010",
  42413=>"011000111",
  42414=>"010000001",
  42415=>"001110000",
  42416=>"110011100",
  42417=>"101110111",
  42418=>"110101110",
  42419=>"110101001",
  42420=>"000000001",
  42421=>"010001001",
  42422=>"100110011",
  42423=>"110101101",
  42424=>"011101100",
  42425=>"001100011",
  42426=>"011001001",
  42427=>"100111101",
  42428=>"011000010",
  42429=>"001011011",
  42430=>"101100110",
  42431=>"001110000",
  42432=>"110101110",
  42433=>"110011001",
  42434=>"010001110",
  42435=>"001010101",
  42436=>"000110010",
  42437=>"110110001",
  42438=>"100001110",
  42439=>"010000010",
  42440=>"010101001",
  42441=>"000101010",
  42442=>"101011111",
  42443=>"100010011",
  42444=>"110101010",
  42445=>"101111101",
  42446=>"010110010",
  42447=>"010110011",
  42448=>"010000101",
  42449=>"101010110",
  42450=>"001111100",
  42451=>"101000011",
  42452=>"111110100",
  42453=>"110110111",
  42454=>"000000001",
  42455=>"101101010",
  42456=>"010001011",
  42457=>"101001110",
  42458=>"011111001",
  42459=>"101100000",
  42460=>"110110011",
  42461=>"010011110",
  42462=>"101001010",
  42463=>"100010111",
  42464=>"011101110",
  42465=>"101111101",
  42466=>"111001101",
  42467=>"001000111",
  42468=>"010000010",
  42469=>"010011111",
  42470=>"100111011",
  42471=>"011110111",
  42472=>"000000001",
  42473=>"100101110",
  42474=>"001000111",
  42475=>"101111000",
  42476=>"111001101",
  42477=>"011101110",
  42478=>"110011011",
  42479=>"011000100",
  42480=>"000000001",
  42481=>"100010000",
  42482=>"100110000",
  42483=>"101011101",
  42484=>"111101101",
  42485=>"101110100",
  42486=>"110000100",
  42487=>"010010101",
  42488=>"001000001",
  42489=>"010111011",
  42490=>"001101100",
  42491=>"110001101",
  42492=>"000010011",
  42493=>"110001011",
  42494=>"100111010",
  42495=>"111101001",
  42496=>"100000000",
  42497=>"010000000",
  42498=>"000111110",
  42499=>"100111101",
  42500=>"111000000",
  42501=>"100010000",
  42502=>"001001111",
  42503=>"001000000",
  42504=>"101101100",
  42505=>"000010000",
  42506=>"001011101",
  42507=>"000011111",
  42508=>"000111111",
  42509=>"100000001",
  42510=>"001010011",
  42511=>"010000011",
  42512=>"011001000",
  42513=>"111010001",
  42514=>"011000001",
  42515=>"100011111",
  42516=>"101011101",
  42517=>"101100101",
  42518=>"011100010",
  42519=>"110110100",
  42520=>"000110110",
  42521=>"100001000",
  42522=>"101100111",
  42523=>"010110110",
  42524=>"101100000",
  42525=>"010001001",
  42526=>"010000001",
  42527=>"010110011",
  42528=>"110111000",
  42529=>"000110010",
  42530=>"001000001",
  42531=>"110011111",
  42532=>"110101111",
  42533=>"000011000",
  42534=>"110101110",
  42535=>"101111101",
  42536=>"001100110",
  42537=>"000001011",
  42538=>"100000111",
  42539=>"110000001",
  42540=>"011110110",
  42541=>"001110111",
  42542=>"100000000",
  42543=>"010101110",
  42544=>"110000010",
  42545=>"110111110",
  42546=>"001001100",
  42547=>"100011001",
  42548=>"101111100",
  42549=>"011101110",
  42550=>"000000010",
  42551=>"000110110",
  42552=>"010000001",
  42553=>"010101110",
  42554=>"000100000",
  42555=>"111011100",
  42556=>"010010000",
  42557=>"001111100",
  42558=>"010110100",
  42559=>"010000100",
  42560=>"111000011",
  42561=>"010000001",
  42562=>"100100000",
  42563=>"101110110",
  42564=>"110101100",
  42565=>"011011000",
  42566=>"010101001",
  42567=>"110110100",
  42568=>"101100101",
  42569=>"110011000",
  42570=>"111110011",
  42571=>"001001100",
  42572=>"000110101",
  42573=>"101111010",
  42574=>"011011101",
  42575=>"110001110",
  42576=>"111011000",
  42577=>"111110000",
  42578=>"010110010",
  42579=>"010101110",
  42580=>"000101011",
  42581=>"001111101",
  42582=>"101110100",
  42583=>"100011001",
  42584=>"011110111",
  42585=>"011110001",
  42586=>"000100010",
  42587=>"100101010",
  42588=>"000001110",
  42589=>"100101001",
  42590=>"001011110",
  42591=>"101010010",
  42592=>"000100101",
  42593=>"000011011",
  42594=>"000001000",
  42595=>"010111111",
  42596=>"001110000",
  42597=>"011010110",
  42598=>"011101111",
  42599=>"110111111",
  42600=>"000101110",
  42601=>"000110000",
  42602=>"001010011",
  42603=>"010110001",
  42604=>"100001110",
  42605=>"100010111",
  42606=>"011100110",
  42607=>"010110000",
  42608=>"010010011",
  42609=>"011010010",
  42610=>"010011110",
  42611=>"101010110",
  42612=>"110101001",
  42613=>"110011101",
  42614=>"000100001",
  42615=>"111100100",
  42616=>"111000010",
  42617=>"011011111",
  42618=>"110111100",
  42619=>"010011011",
  42620=>"000000111",
  42621=>"100110100",
  42622=>"000000111",
  42623=>"011001111",
  42624=>"100101010",
  42625=>"001110000",
  42626=>"110101000",
  42627=>"001110000",
  42628=>"000011000",
  42629=>"110100010",
  42630=>"101001101",
  42631=>"010111000",
  42632=>"111011111",
  42633=>"011110110",
  42634=>"011000010",
  42635=>"000101101",
  42636=>"000010100",
  42637=>"110000100",
  42638=>"110110100",
  42639=>"001000111",
  42640=>"000101010",
  42641=>"000111000",
  42642=>"100010111",
  42643=>"010100111",
  42644=>"110100010",
  42645=>"010111111",
  42646=>"011110111",
  42647=>"000000000",
  42648=>"110110011",
  42649=>"000010001",
  42650=>"100011110",
  42651=>"000110111",
  42652=>"000001101",
  42653=>"110111011",
  42654=>"000011101",
  42655=>"101100010",
  42656=>"000100011",
  42657=>"101000111",
  42658=>"010010111",
  42659=>"111110000",
  42660=>"100100001",
  42661=>"100111111",
  42662=>"111000001",
  42663=>"010000001",
  42664=>"100000011",
  42665=>"111001110",
  42666=>"011011100",
  42667=>"010001001",
  42668=>"001110100",
  42669=>"001000110",
  42670=>"010001000",
  42671=>"001000000",
  42672=>"000100111",
  42673=>"000011101",
  42674=>"010101100",
  42675=>"100100001",
  42676=>"010011101",
  42677=>"111110000",
  42678=>"111000101",
  42679=>"001001100",
  42680=>"111010100",
  42681=>"000000011",
  42682=>"000111101",
  42683=>"010100011",
  42684=>"111000010",
  42685=>"111010110",
  42686=>"000001110",
  42687=>"001010100",
  42688=>"000010000",
  42689=>"111100110",
  42690=>"001011010",
  42691=>"011011001",
  42692=>"111100111",
  42693=>"000001100",
  42694=>"100000100",
  42695=>"001000111",
  42696=>"011010010",
  42697=>"010110110",
  42698=>"100000101",
  42699=>"000101111",
  42700=>"100001100",
  42701=>"111100110",
  42702=>"001101000",
  42703=>"011101110",
  42704=>"101110111",
  42705=>"010010011",
  42706=>"101101101",
  42707=>"000110011",
  42708=>"110011111",
  42709=>"111101101",
  42710=>"000001000",
  42711=>"000111001",
  42712=>"000011101",
  42713=>"101110110",
  42714=>"000101011",
  42715=>"000101010",
  42716=>"010110101",
  42717=>"111010110",
  42718=>"010011110",
  42719=>"111101110",
  42720=>"010000001",
  42721=>"110111000",
  42722=>"110111111",
  42723=>"011100100",
  42724=>"101011010",
  42725=>"010111011",
  42726=>"001011001",
  42727=>"011101011",
  42728=>"100000011",
  42729=>"100101011",
  42730=>"111001111",
  42731=>"101001101",
  42732=>"100101110",
  42733=>"111001011",
  42734=>"011100110",
  42735=>"000001100",
  42736=>"111111010",
  42737=>"001100101",
  42738=>"100110000",
  42739=>"010011000",
  42740=>"110111110",
  42741=>"000110010",
  42742=>"010101111",
  42743=>"101000100",
  42744=>"011000111",
  42745=>"001011001",
  42746=>"011010011",
  42747=>"101100001",
  42748=>"011011101",
  42749=>"001101110",
  42750=>"010100101",
  42751=>"000000010",
  42752=>"000100100",
  42753=>"010000101",
  42754=>"111101111",
  42755=>"100010001",
  42756=>"010100000",
  42757=>"100010011",
  42758=>"100110111",
  42759=>"011000001",
  42760=>"000011100",
  42761=>"010001100",
  42762=>"011100101",
  42763=>"101100010",
  42764=>"111010001",
  42765=>"101001101",
  42766=>"011010000",
  42767=>"000101000",
  42768=>"000000101",
  42769=>"101000111",
  42770=>"110101111",
  42771=>"001010110",
  42772=>"010101110",
  42773=>"000001010",
  42774=>"100010010",
  42775=>"011011110",
  42776=>"001110111",
  42777=>"100011000",
  42778=>"110110100",
  42779=>"001111011",
  42780=>"110010110",
  42781=>"101011111",
  42782=>"101100101",
  42783=>"001000110",
  42784=>"011110111",
  42785=>"010000011",
  42786=>"110101101",
  42787=>"010111110",
  42788=>"001000110",
  42789=>"010101110",
  42790=>"110010100",
  42791=>"111101101",
  42792=>"101001001",
  42793=>"000010110",
  42794=>"010000110",
  42795=>"111110110",
  42796=>"110100010",
  42797=>"110010011",
  42798=>"011100100",
  42799=>"110010110",
  42800=>"110101111",
  42801=>"000000100",
  42802=>"010110111",
  42803=>"100000010",
  42804=>"111100001",
  42805=>"001011001",
  42806=>"001011011",
  42807=>"001100001",
  42808=>"010011111",
  42809=>"100010011",
  42810=>"000111001",
  42811=>"110101001",
  42812=>"101111011",
  42813=>"101110001",
  42814=>"110111101",
  42815=>"101011001",
  42816=>"000111110",
  42817=>"111111100",
  42818=>"001000010",
  42819=>"000100000",
  42820=>"111011100",
  42821=>"011100010",
  42822=>"110000110",
  42823=>"101001001",
  42824=>"101001010",
  42825=>"001001000",
  42826=>"001100010",
  42827=>"010010001",
  42828=>"100101100",
  42829=>"110101100",
  42830=>"110000111",
  42831=>"011010110",
  42832=>"101101110",
  42833=>"111011111",
  42834=>"000100110",
  42835=>"101110111",
  42836=>"000000101",
  42837=>"010001100",
  42838=>"011000001",
  42839=>"101010111",
  42840=>"010100010",
  42841=>"000110101",
  42842=>"100100001",
  42843=>"101001100",
  42844=>"011110111",
  42845=>"100001111",
  42846=>"001111110",
  42847=>"000011011",
  42848=>"010010010",
  42849=>"110010111",
  42850=>"100101010",
  42851=>"001101000",
  42852=>"010100000",
  42853=>"000000101",
  42854=>"101011010",
  42855=>"011000100",
  42856=>"001010110",
  42857=>"111110101",
  42858=>"000010001",
  42859=>"001100001",
  42860=>"100010111",
  42861=>"001110000",
  42862=>"001111100",
  42863=>"100110010",
  42864=>"010111010",
  42865=>"111000001",
  42866=>"011010100",
  42867=>"000010001",
  42868=>"101011001",
  42869=>"000010001",
  42870=>"000101100",
  42871=>"100100000",
  42872=>"011010010",
  42873=>"000000101",
  42874=>"110010100",
  42875=>"101001111",
  42876=>"111101010",
  42877=>"000000011",
  42878=>"000000101",
  42879=>"111111100",
  42880=>"001110101",
  42881=>"100000111",
  42882=>"110010001",
  42883=>"010001011",
  42884=>"110001100",
  42885=>"110011100",
  42886=>"111111100",
  42887=>"001100101",
  42888=>"000001011",
  42889=>"000111111",
  42890=>"111100000",
  42891=>"000000100",
  42892=>"101000000",
  42893=>"011100010",
  42894=>"101100010",
  42895=>"011001000",
  42896=>"111101010",
  42897=>"101000110",
  42898=>"000000011",
  42899=>"000101011",
  42900=>"101110100",
  42901=>"101101111",
  42902=>"010101110",
  42903=>"101100101",
  42904=>"001100110",
  42905=>"111001101",
  42906=>"101111110",
  42907=>"110110111",
  42908=>"111101111",
  42909=>"011001101",
  42910=>"000001110",
  42911=>"010010110",
  42912=>"001000101",
  42913=>"000000111",
  42914=>"010110011",
  42915=>"011001000",
  42916=>"111000111",
  42917=>"001111011",
  42918=>"110010110",
  42919=>"000010011",
  42920=>"000111111",
  42921=>"000111000",
  42922=>"010000001",
  42923=>"111011100",
  42924=>"110000001",
  42925=>"011111011",
  42926=>"000011000",
  42927=>"010110110",
  42928=>"101100010",
  42929=>"000111100",
  42930=>"100000001",
  42931=>"101110100",
  42932=>"000100101",
  42933=>"011110011",
  42934=>"001111011",
  42935=>"100011001",
  42936=>"101011110",
  42937=>"110001010",
  42938=>"010001111",
  42939=>"010101100",
  42940=>"011111001",
  42941=>"111010010",
  42942=>"001101011",
  42943=>"101010110",
  42944=>"111111100",
  42945=>"010111110",
  42946=>"001111111",
  42947=>"011100011",
  42948=>"110111111",
  42949=>"001111001",
  42950=>"010100111",
  42951=>"100111111",
  42952=>"000011000",
  42953=>"111000100",
  42954=>"110011000",
  42955=>"001010000",
  42956=>"001000101",
  42957=>"000011111",
  42958=>"000000011",
  42959=>"101000110",
  42960=>"001101100",
  42961=>"100111100",
  42962=>"000000000",
  42963=>"101100111",
  42964=>"001000001",
  42965=>"011000000",
  42966=>"011101100",
  42967=>"110011101",
  42968=>"111101010",
  42969=>"101011010",
  42970=>"000001010",
  42971=>"001100111",
  42972=>"001101011",
  42973=>"110111100",
  42974=>"111000110",
  42975=>"100010000",
  42976=>"111100010",
  42977=>"110001010",
  42978=>"001100100",
  42979=>"000011101",
  42980=>"011000111",
  42981=>"010100001",
  42982=>"111101001",
  42983=>"100111011",
  42984=>"000010100",
  42985=>"010110010",
  42986=>"011100001",
  42987=>"101001111",
  42988=>"110010100",
  42989=>"011111100",
  42990=>"100000110",
  42991=>"100101010",
  42992=>"111111000",
  42993=>"111101100",
  42994=>"100011110",
  42995=>"011100100",
  42996=>"000000101",
  42997=>"101001011",
  42998=>"000010011",
  42999=>"101100101",
  43000=>"001011110",
  43001=>"101101001",
  43002=>"000000010",
  43003=>"111011001",
  43004=>"011011001",
  43005=>"110001011",
  43006=>"101000010",
  43007=>"010100000",
  43008=>"111100101",
  43009=>"110111011",
  43010=>"100000000",
  43011=>"011110111",
  43012=>"000111011",
  43013=>"010110001",
  43014=>"110111110",
  43015=>"011001001",
  43016=>"010110110",
  43017=>"011100100",
  43018=>"011101001",
  43019=>"010111000",
  43020=>"011110001",
  43021=>"111001010",
  43022=>"100101100",
  43023=>"111110101",
  43024=>"010011000",
  43025=>"011000011",
  43026=>"010000100",
  43027=>"011000001",
  43028=>"110011111",
  43029=>"000100010",
  43030=>"000110010",
  43031=>"101000101",
  43032=>"000000101",
  43033=>"100010011",
  43034=>"111101010",
  43035=>"100010111",
  43036=>"000111011",
  43037=>"000010110",
  43038=>"100111010",
  43039=>"111011101",
  43040=>"111110111",
  43041=>"101001000",
  43042=>"110111000",
  43043=>"110001111",
  43044=>"100101000",
  43045=>"010011111",
  43046=>"001010110",
  43047=>"110001101",
  43048=>"010110111",
  43049=>"100111000",
  43050=>"100010011",
  43051=>"110001111",
  43052=>"110000100",
  43053=>"000000010",
  43054=>"111001010",
  43055=>"000000011",
  43056=>"111000101",
  43057=>"011100111",
  43058=>"001100110",
  43059=>"111111011",
  43060=>"111111000",
  43061=>"011000100",
  43062=>"101000110",
  43063=>"000011110",
  43064=>"111011100",
  43065=>"010010110",
  43066=>"010100101",
  43067=>"000000001",
  43068=>"101101010",
  43069=>"000110101",
  43070=>"111100000",
  43071=>"011011001",
  43072=>"110001100",
  43073=>"010111111",
  43074=>"110010101",
  43075=>"000101011",
  43076=>"111011000",
  43077=>"100101001",
  43078=>"010100111",
  43079=>"111010110",
  43080=>"101011111",
  43081=>"110101111",
  43082=>"011101000",
  43083=>"101111001",
  43084=>"010100100",
  43085=>"110111110",
  43086=>"100011110",
  43087=>"111011110",
  43088=>"000100000",
  43089=>"111000010",
  43090=>"101011010",
  43091=>"101010111",
  43092=>"111111110",
  43093=>"101011100",
  43094=>"000100110",
  43095=>"001011000",
  43096=>"110010100",
  43097=>"011100101",
  43098=>"110000101",
  43099=>"001101101",
  43100=>"101001010",
  43101=>"000001000",
  43102=>"000010000",
  43103=>"100101101",
  43104=>"010011010",
  43105=>"000000001",
  43106=>"100011101",
  43107=>"111100000",
  43108=>"011001110",
  43109=>"101001110",
  43110=>"010000100",
  43111=>"100010110",
  43112=>"100011001",
  43113=>"111111001",
  43114=>"011010111",
  43115=>"011110111",
  43116=>"000011001",
  43117=>"011011110",
  43118=>"100011000",
  43119=>"000010011",
  43120=>"101000011",
  43121=>"000111100",
  43122=>"010011000",
  43123=>"111001110",
  43124=>"101100010",
  43125=>"010100010",
  43126=>"000100111",
  43127=>"110010100",
  43128=>"010001100",
  43129=>"101010000",
  43130=>"100111111",
  43131=>"011101101",
  43132=>"101001000",
  43133=>"011110100",
  43134=>"101001101",
  43135=>"000000000",
  43136=>"101010001",
  43137=>"001011010",
  43138=>"011000010",
  43139=>"000111000",
  43140=>"011010001",
  43141=>"011101000",
  43142=>"011110100",
  43143=>"010101111",
  43144=>"110110100",
  43145=>"001110101",
  43146=>"111111001",
  43147=>"010011010",
  43148=>"000010100",
  43149=>"000101110",
  43150=>"000100100",
  43151=>"011111101",
  43152=>"000011001",
  43153=>"010011100",
  43154=>"001110000",
  43155=>"011011011",
  43156=>"101000010",
  43157=>"011110010",
  43158=>"110101101",
  43159=>"000001101",
  43160=>"011100110",
  43161=>"010000011",
  43162=>"001111111",
  43163=>"011011011",
  43164=>"101101000",
  43165=>"110110010",
  43166=>"100001101",
  43167=>"110100010",
  43168=>"011000011",
  43169=>"100010011",
  43170=>"011110101",
  43171=>"001111101",
  43172=>"101111011",
  43173=>"001001000",
  43174=>"100100001",
  43175=>"110100010",
  43176=>"000111110",
  43177=>"100110000",
  43178=>"011000110",
  43179=>"001011100",
  43180=>"110111111",
  43181=>"110001010",
  43182=>"101000111",
  43183=>"110100011",
  43184=>"101001011",
  43185=>"010001110",
  43186=>"001111111",
  43187=>"000111101",
  43188=>"001000001",
  43189=>"001000000",
  43190=>"111000111",
  43191=>"111110011",
  43192=>"000100111",
  43193=>"101011001",
  43194=>"001110100",
  43195=>"000110011",
  43196=>"111001011",
  43197=>"111111111",
  43198=>"001000001",
  43199=>"100111101",
  43200=>"101000000",
  43201=>"010111100",
  43202=>"111100000",
  43203=>"010101111",
  43204=>"111001101",
  43205=>"111101101",
  43206=>"100111100",
  43207=>"011011010",
  43208=>"100011010",
  43209=>"101111100",
  43210=>"101110110",
  43211=>"110111001",
  43212=>"100000001",
  43213=>"000010010",
  43214=>"111001001",
  43215=>"100000001",
  43216=>"111010110",
  43217=>"011011010",
  43218=>"011111000",
  43219=>"000111001",
  43220=>"110010001",
  43221=>"011100010",
  43222=>"110100010",
  43223=>"000000000",
  43224=>"110011101",
  43225=>"101101101",
  43226=>"111110010",
  43227=>"100111111",
  43228=>"000000101",
  43229=>"010001011",
  43230=>"100101110",
  43231=>"110011101",
  43232=>"011101000",
  43233=>"000000001",
  43234=>"101000011",
  43235=>"001101101",
  43236=>"100000001",
  43237=>"100101001",
  43238=>"110011110",
  43239=>"010001000",
  43240=>"011001011",
  43241=>"111010110",
  43242=>"111110101",
  43243=>"000011110",
  43244=>"001010100",
  43245=>"000111001",
  43246=>"111010010",
  43247=>"000010110",
  43248=>"000101110",
  43249=>"110110111",
  43250=>"001010111",
  43251=>"000010110",
  43252=>"111111101",
  43253=>"010011100",
  43254=>"011110010",
  43255=>"111100101",
  43256=>"010101100",
  43257=>"101100011",
  43258=>"000010001",
  43259=>"111101111",
  43260=>"010100000",
  43261=>"100010101",
  43262=>"111000011",
  43263=>"100110111",
  43264=>"100111100",
  43265=>"000011110",
  43266=>"101110010",
  43267=>"101000110",
  43268=>"010001100",
  43269=>"110110100",
  43270=>"001110100",
  43271=>"010010100",
  43272=>"000111111",
  43273=>"001110111",
  43274=>"100001011",
  43275=>"100110101",
  43276=>"001011000",
  43277=>"011100011",
  43278=>"111100111",
  43279=>"100110000",
  43280=>"101000100",
  43281=>"001001111",
  43282=>"100001110",
  43283=>"000000101",
  43284=>"000001001",
  43285=>"111111000",
  43286=>"100000010",
  43287=>"011111101",
  43288=>"110100001",
  43289=>"000000110",
  43290=>"000101001",
  43291=>"110001010",
  43292=>"110101110",
  43293=>"101001011",
  43294=>"111100111",
  43295=>"100110000",
  43296=>"010010111",
  43297=>"110011000",
  43298=>"111110100",
  43299=>"001111010",
  43300=>"011101000",
  43301=>"110000010",
  43302=>"011110001",
  43303=>"111000100",
  43304=>"001000001",
  43305=>"111001111",
  43306=>"001100001",
  43307=>"101000011",
  43308=>"101110010",
  43309=>"111111111",
  43310=>"001111100",
  43311=>"100100110",
  43312=>"011111000",
  43313=>"111001001",
  43314=>"111111111",
  43315=>"100101101",
  43316=>"100010000",
  43317=>"001100111",
  43318=>"000100101",
  43319=>"001000101",
  43320=>"111000100",
  43321=>"000101000",
  43322=>"111010110",
  43323=>"100111010",
  43324=>"100001100",
  43325=>"110000101",
  43326=>"000001011",
  43327=>"111000110",
  43328=>"000110000",
  43329=>"111101111",
  43330=>"110111010",
  43331=>"111100101",
  43332=>"101111001",
  43333=>"100010111",
  43334=>"011010000",
  43335=>"011001000",
  43336=>"001011111",
  43337=>"100110000",
  43338=>"010000101",
  43339=>"011111111",
  43340=>"000001011",
  43341=>"011101001",
  43342=>"000111101",
  43343=>"000101001",
  43344=>"011101010",
  43345=>"001101001",
  43346=>"100000100",
  43347=>"111010001",
  43348=>"111111010",
  43349=>"111011000",
  43350=>"001110101",
  43351=>"100110010",
  43352=>"101011010",
  43353=>"001001100",
  43354=>"111100101",
  43355=>"101001101",
  43356=>"111111100",
  43357=>"111000111",
  43358=>"111110011",
  43359=>"000001001",
  43360=>"011000001",
  43361=>"000000000",
  43362=>"111000010",
  43363=>"011110111",
  43364=>"010111011",
  43365=>"000000010",
  43366=>"110000111",
  43367=>"010111011",
  43368=>"010100100",
  43369=>"111101111",
  43370=>"001010010",
  43371=>"110100110",
  43372=>"101101010",
  43373=>"011100110",
  43374=>"001110101",
  43375=>"100111100",
  43376=>"101001000",
  43377=>"001100101",
  43378=>"001100011",
  43379=>"011010111",
  43380=>"011001000",
  43381=>"011010010",
  43382=>"000101100",
  43383=>"100011010",
  43384=>"000010011",
  43385=>"001101101",
  43386=>"110110101",
  43387=>"100001110",
  43388=>"110000111",
  43389=>"011001001",
  43390=>"000011101",
  43391=>"011100111",
  43392=>"000110010",
  43393=>"001111011",
  43394=>"011110110",
  43395=>"111011000",
  43396=>"010110110",
  43397=>"001100000",
  43398=>"110011100",
  43399=>"111110110",
  43400=>"001001000",
  43401=>"100001000",
  43402=>"101000111",
  43403=>"100011101",
  43404=>"111111011",
  43405=>"100111001",
  43406=>"011111111",
  43407=>"111111100",
  43408=>"011100011",
  43409=>"000001111",
  43410=>"110110111",
  43411=>"000001000",
  43412=>"111110011",
  43413=>"001100001",
  43414=>"110000000",
  43415=>"010101100",
  43416=>"011101110",
  43417=>"010100000",
  43418=>"011001111",
  43419=>"010100000",
  43420=>"110110010",
  43421=>"011101101",
  43422=>"111100110",
  43423=>"000111111",
  43424=>"010100110",
  43425=>"011100000",
  43426=>"001010000",
  43427=>"001001011",
  43428=>"101000000",
  43429=>"000001011",
  43430=>"100110111",
  43431=>"111001110",
  43432=>"000100101",
  43433=>"000001000",
  43434=>"111101100",
  43435=>"100100010",
  43436=>"001010000",
  43437=>"011100111",
  43438=>"010100001",
  43439=>"111001101",
  43440=>"010000110",
  43441=>"010100101",
  43442=>"000011001",
  43443=>"010101000",
  43444=>"000101011",
  43445=>"010010000",
  43446=>"000100101",
  43447=>"100010000",
  43448=>"100100110",
  43449=>"010101010",
  43450=>"110101110",
  43451=>"011010111",
  43452=>"111101011",
  43453=>"101000111",
  43454=>"111110100",
  43455=>"001000100",
  43456=>"000110011",
  43457=>"001010100",
  43458=>"111000100",
  43459=>"000000100",
  43460=>"000011010",
  43461=>"111001111",
  43462=>"100001010",
  43463=>"110100110",
  43464=>"011010111",
  43465=>"010010111",
  43466=>"011000111",
  43467=>"100010101",
  43468=>"011110001",
  43469=>"111000001",
  43470=>"110111111",
  43471=>"011101101",
  43472=>"101011101",
  43473=>"001111001",
  43474=>"001001001",
  43475=>"111001011",
  43476=>"111000000",
  43477=>"001111000",
  43478=>"101010001",
  43479=>"001111101",
  43480=>"111010100",
  43481=>"010110001",
  43482=>"100000000",
  43483=>"110011001",
  43484=>"010011101",
  43485=>"101100100",
  43486=>"010000110",
  43487=>"010111100",
  43488=>"101111011",
  43489=>"000111010",
  43490=>"101111111",
  43491=>"111110111",
  43492=>"101100111",
  43493=>"101100011",
  43494=>"001100100",
  43495=>"100110000",
  43496=>"100011011",
  43497=>"111111000",
  43498=>"000110100",
  43499=>"110001111",
  43500=>"110011110",
  43501=>"111110000",
  43502=>"101101111",
  43503=>"011011000",
  43504=>"011100100",
  43505=>"001000110",
  43506=>"101010101",
  43507=>"111001000",
  43508=>"101000010",
  43509=>"001010011",
  43510=>"011101111",
  43511=>"001100011",
  43512=>"110110001",
  43513=>"101000001",
  43514=>"010000000",
  43515=>"001100110",
  43516=>"000011000",
  43517=>"100000011",
  43518=>"111000110",
  43519=>"010000100",
  43520=>"010000111",
  43521=>"000111011",
  43522=>"111011011",
  43523=>"111001000",
  43524=>"000100110",
  43525=>"110101110",
  43526=>"100010010",
  43527=>"111011000",
  43528=>"100100001",
  43529=>"111011111",
  43530=>"110111111",
  43531=>"001110111",
  43532=>"010011100",
  43533=>"011101000",
  43534=>"000101000",
  43535=>"110110111",
  43536=>"011001010",
  43537=>"101001000",
  43538=>"110001011",
  43539=>"011000000",
  43540=>"100101101",
  43541=>"011101000",
  43542=>"000110101",
  43543=>"101000110",
  43544=>"001100111",
  43545=>"100100110",
  43546=>"000100010",
  43547=>"000001000",
  43548=>"100010110",
  43549=>"011010001",
  43550=>"010101000",
  43551=>"000000000",
  43552=>"001000000",
  43553=>"001110011",
  43554=>"010111111",
  43555=>"000000000",
  43556=>"110011111",
  43557=>"000000011",
  43558=>"111011001",
  43559=>"010101101",
  43560=>"000101001",
  43561=>"011000110",
  43562=>"000000011",
  43563=>"010101100",
  43564=>"001110110",
  43565=>"100110011",
  43566=>"000110110",
  43567=>"000101001",
  43568=>"011100111",
  43569=>"011101011",
  43570=>"100010110",
  43571=>"110010111",
  43572=>"001100100",
  43573=>"001001111",
  43574=>"100011111",
  43575=>"010100111",
  43576=>"111111101",
  43577=>"010000000",
  43578=>"001101101",
  43579=>"001010111",
  43580=>"000001011",
  43581=>"010001011",
  43582=>"010111111",
  43583=>"110100111",
  43584=>"111111001",
  43585=>"111110011",
  43586=>"100010011",
  43587=>"001100100",
  43588=>"101111000",
  43589=>"110000100",
  43590=>"111110111",
  43591=>"011101111",
  43592=>"000001001",
  43593=>"100111011",
  43594=>"100000010",
  43595=>"000100010",
  43596=>"101111111",
  43597=>"010100011",
  43598=>"010011110",
  43599=>"010100100",
  43600=>"011001011",
  43601=>"100100010",
  43602=>"111011010",
  43603=>"000000010",
  43604=>"100100010",
  43605=>"110111111",
  43606=>"010000111",
  43607=>"100010010",
  43608=>"100010111",
  43609=>"100110101",
  43610=>"000010100",
  43611=>"001000011",
  43612=>"000001111",
  43613=>"111011101",
  43614=>"111000101",
  43615=>"100111011",
  43616=>"000101111",
  43617=>"101111101",
  43618=>"010111011",
  43619=>"100100000",
  43620=>"100100000",
  43621=>"110100100",
  43622=>"101000100",
  43623=>"101000010",
  43624=>"101100010",
  43625=>"010001101",
  43626=>"100010000",
  43627=>"000010110",
  43628=>"100010101",
  43629=>"000000010",
  43630=>"100101110",
  43631=>"000001110",
  43632=>"101010000",
  43633=>"101110110",
  43634=>"010101010",
  43635=>"101000001",
  43636=>"011000010",
  43637=>"000010000",
  43638=>"011110000",
  43639=>"101100111",
  43640=>"110011111",
  43641=>"100000000",
  43642=>"010000011",
  43643=>"101110000",
  43644=>"011100001",
  43645=>"111111101",
  43646=>"010111010",
  43647=>"111000110",
  43648=>"001111100",
  43649=>"001110011",
  43650=>"110010110",
  43651=>"001011010",
  43652=>"000110111",
  43653=>"100110011",
  43654=>"111001101",
  43655=>"000101010",
  43656=>"000100010",
  43657=>"111111011",
  43658=>"100111101",
  43659=>"011100000",
  43660=>"001011000",
  43661=>"001100011",
  43662=>"000110000",
  43663=>"110110101",
  43664=>"010111111",
  43665=>"101100001",
  43666=>"011000000",
  43667=>"101100110",
  43668=>"000000111",
  43669=>"011010101",
  43670=>"100000111",
  43671=>"000010110",
  43672=>"010111011",
  43673=>"100000100",
  43674=>"100001010",
  43675=>"000100101",
  43676=>"111111101",
  43677=>"011111010",
  43678=>"111000101",
  43679=>"100111011",
  43680=>"101111010",
  43681=>"011001110",
  43682=>"110101111",
  43683=>"100001011",
  43684=>"100000011",
  43685=>"000001100",
  43686=>"000000111",
  43687=>"000001010",
  43688=>"110011000",
  43689=>"010001101",
  43690=>"000101000",
  43691=>"011000110",
  43692=>"011010001",
  43693=>"010100011",
  43694=>"001110001",
  43695=>"110001100",
  43696=>"001111010",
  43697=>"110100111",
  43698=>"011111001",
  43699=>"110111010",
  43700=>"001011001",
  43701=>"010010010",
  43702=>"000100100",
  43703=>"011111000",
  43704=>"001001111",
  43705=>"110100001",
  43706=>"010101001",
  43707=>"010100000",
  43708=>"010100000",
  43709=>"110010001",
  43710=>"011110110",
  43711=>"001000001",
  43712=>"111101000",
  43713=>"011111111",
  43714=>"000010010",
  43715=>"001010010",
  43716=>"111111011",
  43717=>"101000111",
  43718=>"001110010",
  43719=>"000110010",
  43720=>"011110100",
  43721=>"110000011",
  43722=>"111101001",
  43723=>"100111101",
  43724=>"111000001",
  43725=>"110000001",
  43726=>"001100011",
  43727=>"000101001",
  43728=>"111111101",
  43729=>"000110000",
  43730=>"111000010",
  43731=>"000000001",
  43732=>"111110110",
  43733=>"101000011",
  43734=>"001100000",
  43735=>"001001100",
  43736=>"001010101",
  43737=>"110101010",
  43738=>"110100101",
  43739=>"111001001",
  43740=>"000101011",
  43741=>"010000010",
  43742=>"000000000",
  43743=>"011110110",
  43744=>"101001110",
  43745=>"101010000",
  43746=>"001110100",
  43747=>"101000101",
  43748=>"100000000",
  43749=>"110011010",
  43750=>"001101011",
  43751=>"000111000",
  43752=>"100101001",
  43753=>"111110111",
  43754=>"111101111",
  43755=>"100100101",
  43756=>"001001100",
  43757=>"011101011",
  43758=>"011001000",
  43759=>"111000000",
  43760=>"101000010",
  43761=>"111000001",
  43762=>"000100110",
  43763=>"000011101",
  43764=>"101110110",
  43765=>"011011000",
  43766=>"010000010",
  43767=>"100111111",
  43768=>"110111010",
  43769=>"001010001",
  43770=>"110101000",
  43771=>"111010001",
  43772=>"000000111",
  43773=>"010111000",
  43774=>"101100111",
  43775=>"110010101",
  43776=>"100100001",
  43777=>"110100000",
  43778=>"011000010",
  43779=>"011111101",
  43780=>"100000010",
  43781=>"100010001",
  43782=>"111010011",
  43783=>"100010101",
  43784=>"010111000",
  43785=>"001010111",
  43786=>"110010100",
  43787=>"011111000",
  43788=>"011101010",
  43789=>"110000101",
  43790=>"010011001",
  43791=>"111010001",
  43792=>"110011001",
  43793=>"001010000",
  43794=>"000000111",
  43795=>"110110111",
  43796=>"111001100",
  43797=>"011011111",
  43798=>"100101111",
  43799=>"000000000",
  43800=>"101001001",
  43801=>"000010001",
  43802=>"000111111",
  43803=>"010010111",
  43804=>"001111000",
  43805=>"101000101",
  43806=>"001101100",
  43807=>"010010110",
  43808=>"011101110",
  43809=>"000001111",
  43810=>"010101101",
  43811=>"010100001",
  43812=>"010001101",
  43813=>"010000110",
  43814=>"011011000",
  43815=>"000000010",
  43816=>"111100011",
  43817=>"101010011",
  43818=>"100100011",
  43819=>"111110111",
  43820=>"000110011",
  43821=>"101011010",
  43822=>"001001000",
  43823=>"010110110",
  43824=>"100100001",
  43825=>"111011010",
  43826=>"111111001",
  43827=>"010010001",
  43828=>"011111111",
  43829=>"111011110",
  43830=>"110011111",
  43831=>"110001011",
  43832=>"101111101",
  43833=>"101010010",
  43834=>"101000000",
  43835=>"011001101",
  43836=>"110000111",
  43837=>"000001010",
  43838=>"001000001",
  43839=>"100110111",
  43840=>"010100110",
  43841=>"001100111",
  43842=>"010110011",
  43843=>"100110111",
  43844=>"000101000",
  43845=>"101001000",
  43846=>"101010101",
  43847=>"000110101",
  43848=>"111000111",
  43849=>"111111111",
  43850=>"110000100",
  43851=>"100111111",
  43852=>"111001100",
  43853=>"110001100",
  43854=>"011011000",
  43855=>"010100111",
  43856=>"010101010",
  43857=>"010000001",
  43858=>"100001110",
  43859=>"010111110",
  43860=>"110110000",
  43861=>"101101100",
  43862=>"110001111",
  43863=>"010110111",
  43864=>"010001000",
  43865=>"011011111",
  43866=>"001111000",
  43867=>"001001001",
  43868=>"001111010",
  43869=>"001001001",
  43870=>"011011000",
  43871=>"000100100",
  43872=>"010101010",
  43873=>"000101000",
  43874=>"010011110",
  43875=>"111000011",
  43876=>"111101101",
  43877=>"000110100",
  43878=>"101011011",
  43879=>"000000011",
  43880=>"111001101",
  43881=>"101111101",
  43882=>"110011000",
  43883=>"010101100",
  43884=>"111011011",
  43885=>"001000000",
  43886=>"001100100",
  43887=>"111000110",
  43888=>"001100111",
  43889=>"111101110",
  43890=>"100000101",
  43891=>"010001010",
  43892=>"111000001",
  43893=>"110100010",
  43894=>"001101011",
  43895=>"101101011",
  43896=>"111100000",
  43897=>"001010000",
  43898=>"111110111",
  43899=>"110011000",
  43900=>"111110000",
  43901=>"010101101",
  43902=>"010110111",
  43903=>"111110101",
  43904=>"000011000",
  43905=>"010110011",
  43906=>"001001110",
  43907=>"110111100",
  43908=>"001010100",
  43909=>"011010010",
  43910=>"100001111",
  43911=>"001001001",
  43912=>"000101110",
  43913=>"010101011",
  43914=>"111111000",
  43915=>"000010000",
  43916=>"110011010",
  43917=>"110101011",
  43918=>"100011011",
  43919=>"110110011",
  43920=>"100000010",
  43921=>"000110010",
  43922=>"101110100",
  43923=>"011101001",
  43924=>"111111111",
  43925=>"011011110",
  43926=>"000101000",
  43927=>"111100011",
  43928=>"110011000",
  43929=>"011111111",
  43930=>"000011111",
  43931=>"001010000",
  43932=>"000011001",
  43933=>"100100011",
  43934=>"111111001",
  43935=>"110101111",
  43936=>"100000001",
  43937=>"101001111",
  43938=>"101011011",
  43939=>"000110111",
  43940=>"001110100",
  43941=>"000110110",
  43942=>"001000100",
  43943=>"000100000",
  43944=>"100101100",
  43945=>"010011001",
  43946=>"000000101",
  43947=>"111100001",
  43948=>"100001001",
  43949=>"111111100",
  43950=>"010001000",
  43951=>"110110110",
  43952=>"010010000",
  43953=>"111010001",
  43954=>"011111100",
  43955=>"010100101",
  43956=>"011101001",
  43957=>"111010011",
  43958=>"101011011",
  43959=>"010001100",
  43960=>"011000100",
  43961=>"011110101",
  43962=>"101010010",
  43963=>"111100001",
  43964=>"101001000",
  43965=>"010011011",
  43966=>"100101110",
  43967=>"110110011",
  43968=>"111101010",
  43969=>"111000100",
  43970=>"110111100",
  43971=>"011111010",
  43972=>"011011001",
  43973=>"011000001",
  43974=>"000010000",
  43975=>"011010010",
  43976=>"100101010",
  43977=>"101111110",
  43978=>"101000110",
  43979=>"110110101",
  43980=>"100001110",
  43981=>"110010110",
  43982=>"000011010",
  43983=>"000000110",
  43984=>"110011010",
  43985=>"101000000",
  43986=>"111000111",
  43987=>"100000001",
  43988=>"001001000",
  43989=>"111111110",
  43990=>"111101010",
  43991=>"100001010",
  43992=>"000010101",
  43993=>"011011110",
  43994=>"101111000",
  43995=>"001001110",
  43996=>"101101111",
  43997=>"000001000",
  43998=>"111111111",
  43999=>"000101100",
  44000=>"001011111",
  44001=>"110011110",
  44002=>"100011110",
  44003=>"001111010",
  44004=>"010111000",
  44005=>"110100110",
  44006=>"000100001",
  44007=>"101110011",
  44008=>"010111100",
  44009=>"001011100",
  44010=>"100101101",
  44011=>"000000110",
  44012=>"010111100",
  44013=>"110010100",
  44014=>"000111011",
  44015=>"000000111",
  44016=>"011001111",
  44017=>"000011010",
  44018=>"001110101",
  44019=>"111110101",
  44020=>"110011100",
  44021=>"000001001",
  44022=>"001001011",
  44023=>"101011110",
  44024=>"001000010",
  44025=>"000011011",
  44026=>"100000010",
  44027=>"100010101",
  44028=>"111011000",
  44029=>"000011100",
  44030=>"101100001",
  44031=>"001000100",
  44032=>"010101000",
  44033=>"110010110",
  44034=>"011100100",
  44035=>"001011111",
  44036=>"001001001",
  44037=>"001011001",
  44038=>"100000111",
  44039=>"000000110",
  44040=>"100101010",
  44041=>"001001010",
  44042=>"111000001",
  44043=>"101101011",
  44044=>"011001011",
  44045=>"100011111",
  44046=>"100101011",
  44047=>"000001110",
  44048=>"000110101",
  44049=>"111110100",
  44050=>"011100101",
  44051=>"111001011",
  44052=>"011000010",
  44053=>"011011011",
  44054=>"011011111",
  44055=>"000101001",
  44056=>"111011101",
  44057=>"000011101",
  44058=>"111011010",
  44059=>"001000100",
  44060=>"001110010",
  44061=>"010101001",
  44062=>"011111010",
  44063=>"011001001",
  44064=>"101000111",
  44065=>"001000110",
  44066=>"100000100",
  44067=>"101011000",
  44068=>"000010110",
  44069=>"011110111",
  44070=>"000101000",
  44071=>"101011010",
  44072=>"110100111",
  44073=>"111111101",
  44074=>"100001100",
  44075=>"111010010",
  44076=>"100011100",
  44077=>"101100100",
  44078=>"101011110",
  44079=>"100011000",
  44080=>"001010000",
  44081=>"001000101",
  44082=>"001110001",
  44083=>"101000111",
  44084=>"000110011",
  44085=>"111101011",
  44086=>"011010010",
  44087=>"010111000",
  44088=>"100000011",
  44089=>"001111110",
  44090=>"110111011",
  44091=>"101011101",
  44092=>"011111000",
  44093=>"111011011",
  44094=>"011101100",
  44095=>"001000111",
  44096=>"000000000",
  44097=>"110001011",
  44098=>"110011011",
  44099=>"001000110",
  44100=>"111011011",
  44101=>"110101001",
  44102=>"101001011",
  44103=>"000111000",
  44104=>"011111011",
  44105=>"010111001",
  44106=>"010001010",
  44107=>"101000000",
  44108=>"101111101",
  44109=>"011100100",
  44110=>"010011011",
  44111=>"010001010",
  44112=>"000110000",
  44113=>"000001111",
  44114=>"110000111",
  44115=>"000001100",
  44116=>"111010001",
  44117=>"010110011",
  44118=>"010100010",
  44119=>"011101101",
  44120=>"111101000",
  44121=>"110111111",
  44122=>"010100111",
  44123=>"001001110",
  44124=>"010101011",
  44125=>"000100100",
  44126=>"100111101",
  44127=>"101111010",
  44128=>"111001011",
  44129=>"001111011",
  44130=>"110110000",
  44131=>"011001011",
  44132=>"001000100",
  44133=>"100101110",
  44134=>"001010011",
  44135=>"000110101",
  44136=>"001011000",
  44137=>"001100011",
  44138=>"111110010",
  44139=>"111111111",
  44140=>"101101100",
  44141=>"011001100",
  44142=>"101010001",
  44143=>"001110111",
  44144=>"111110111",
  44145=>"001101011",
  44146=>"000011011",
  44147=>"100011010",
  44148=>"101010100",
  44149=>"110111001",
  44150=>"111001111",
  44151=>"010101010",
  44152=>"001101000",
  44153=>"011000101",
  44154=>"010001010",
  44155=>"001010011",
  44156=>"010001101",
  44157=>"010101000",
  44158=>"010010000",
  44159=>"111111001",
  44160=>"101001001",
  44161=>"001001110",
  44162=>"001001010",
  44163=>"110111111",
  44164=>"000101111",
  44165=>"101111111",
  44166=>"011011100",
  44167=>"010000001",
  44168=>"100111001",
  44169=>"111000011",
  44170=>"000110100",
  44171=>"111011010",
  44172=>"100100010",
  44173=>"001000010",
  44174=>"000001111",
  44175=>"011011000",
  44176=>"110100111",
  44177=>"111110010",
  44178=>"101011010",
  44179=>"101011011",
  44180=>"100100011",
  44181=>"010111000",
  44182=>"001111001",
  44183=>"000101011",
  44184=>"000011101",
  44185=>"111111111",
  44186=>"001000000",
  44187=>"000111110",
  44188=>"011110011",
  44189=>"000101001",
  44190=>"000011001",
  44191=>"001100000",
  44192=>"001011001",
  44193=>"010010011",
  44194=>"100110000",
  44195=>"101100101",
  44196=>"100000001",
  44197=>"101101001",
  44198=>"011000001",
  44199=>"010100001",
  44200=>"111001010",
  44201=>"010101100",
  44202=>"100101000",
  44203=>"000101110",
  44204=>"111111010",
  44205=>"001001011",
  44206=>"111100000",
  44207=>"011011010",
  44208=>"111111011",
  44209=>"000110011",
  44210=>"101001000",
  44211=>"101001100",
  44212=>"111111011",
  44213=>"111010110",
  44214=>"111000110",
  44215=>"000000001",
  44216=>"000011100",
  44217=>"001110011",
  44218=>"011010100",
  44219=>"101011111",
  44220=>"011111001",
  44221=>"101100011",
  44222=>"000101010",
  44223=>"100010000",
  44224=>"110001101",
  44225=>"111111110",
  44226=>"111011000",
  44227=>"100100011",
  44228=>"111100000",
  44229=>"000010111",
  44230=>"100100001",
  44231=>"000100110",
  44232=>"111011001",
  44233=>"110110110",
  44234=>"000101001",
  44235=>"001110100",
  44236=>"010100011",
  44237=>"000010101",
  44238=>"111001111",
  44239=>"001010001",
  44240=>"001011001",
  44241=>"110111001",
  44242=>"100001000",
  44243=>"101010111",
  44244=>"101001001",
  44245=>"001101001",
  44246=>"011010000",
  44247=>"000010001",
  44248=>"001001101",
  44249=>"110010000",
  44250=>"110110000",
  44251=>"000001110",
  44252=>"111111010",
  44253=>"011100110",
  44254=>"001011100",
  44255=>"110111100",
  44256=>"001101000",
  44257=>"011000000",
  44258=>"010000001",
  44259=>"011001110",
  44260=>"100110100",
  44261=>"101101011",
  44262=>"010111000",
  44263=>"001111000",
  44264=>"010100000",
  44265=>"110111111",
  44266=>"101111101",
  44267=>"001011000",
  44268=>"000001010",
  44269=>"100111110",
  44270=>"101001001",
  44271=>"111011111",
  44272=>"001010110",
  44273=>"001101000",
  44274=>"010011011",
  44275=>"100010001",
  44276=>"010101011",
  44277=>"000011111",
  44278=>"011101011",
  44279=>"111001111",
  44280=>"001000110",
  44281=>"101001100",
  44282=>"110011000",
  44283=>"100110111",
  44284=>"010000001",
  44285=>"011000010",
  44286=>"010010111",
  44287=>"101010000",
  44288=>"101011010",
  44289=>"101111000",
  44290=>"010001010",
  44291=>"101011000",
  44292=>"010001000",
  44293=>"101010001",
  44294=>"011001100",
  44295=>"101001011",
  44296=>"010111001",
  44297=>"111111001",
  44298=>"000111101",
  44299=>"011110000",
  44300=>"111000001",
  44301=>"100000000",
  44302=>"110111110",
  44303=>"011000011",
  44304=>"111010001",
  44305=>"000001001",
  44306=>"000010011",
  44307=>"110000011",
  44308=>"101000000",
  44309=>"011111111",
  44310=>"111001110",
  44311=>"111100001",
  44312=>"111010111",
  44313=>"000011001",
  44314=>"011011000",
  44315=>"110011011",
  44316=>"100011100",
  44317=>"110110001",
  44318=>"110010110",
  44319=>"100011110",
  44320=>"101001111",
  44321=>"011011000",
  44322=>"001101101",
  44323=>"100011011",
  44324=>"101000010",
  44325=>"110011010",
  44326=>"011101011",
  44327=>"000001100",
  44328=>"001101111",
  44329=>"100111110",
  44330=>"011100000",
  44331=>"000001011",
  44332=>"110001000",
  44333=>"011001101",
  44334=>"100011101",
  44335=>"001011100",
  44336=>"101011011",
  44337=>"010010010",
  44338=>"110101111",
  44339=>"011001010",
  44340=>"100110111",
  44341=>"011110101",
  44342=>"110111000",
  44343=>"000111000",
  44344=>"001001111",
  44345=>"011100100",
  44346=>"000010010",
  44347=>"001001000",
  44348=>"000100010",
  44349=>"110101011",
  44350=>"101111010",
  44351=>"001011101",
  44352=>"111111001",
  44353=>"011001111",
  44354=>"101100001",
  44355=>"111101000",
  44356=>"101110111",
  44357=>"010000111",
  44358=>"001101000",
  44359=>"100001000",
  44360=>"111010110",
  44361=>"111011000",
  44362=>"010010111",
  44363=>"001100010",
  44364=>"100001111",
  44365=>"000111111",
  44366=>"000001011",
  44367=>"101101010",
  44368=>"101111100",
  44369=>"100101101",
  44370=>"000011010",
  44371=>"110111000",
  44372=>"110100111",
  44373=>"111010110",
  44374=>"111101001",
  44375=>"010101101",
  44376=>"100000010",
  44377=>"000000011",
  44378=>"111001110",
  44379=>"000001000",
  44380=>"010011101",
  44381=>"101111011",
  44382=>"010001111",
  44383=>"011100110",
  44384=>"000001111",
  44385=>"011110000",
  44386=>"111111000",
  44387=>"000111110",
  44388=>"001011010",
  44389=>"111110111",
  44390=>"100111000",
  44391=>"001010100",
  44392=>"001101101",
  44393=>"011011100",
  44394=>"011011011",
  44395=>"111010000",
  44396=>"110101010",
  44397=>"000100011",
  44398=>"001000100",
  44399=>"100000110",
  44400=>"011011101",
  44401=>"110011001",
  44402=>"110110011",
  44403=>"010110010",
  44404=>"000100010",
  44405=>"110101111",
  44406=>"111100101",
  44407=>"111001011",
  44408=>"000100100",
  44409=>"110010101",
  44410=>"110001101",
  44411=>"101010100",
  44412=>"010110001",
  44413=>"000001010",
  44414=>"011000111",
  44415=>"011011001",
  44416=>"001011011",
  44417=>"011101100",
  44418=>"101001010",
  44419=>"101011001",
  44420=>"100110100",
  44421=>"111101110",
  44422=>"011111100",
  44423=>"000001011",
  44424=>"111001101",
  44425=>"100100010",
  44426=>"001110010",
  44427=>"000101000",
  44428=>"001001011",
  44429=>"110001111",
  44430=>"111011000",
  44431=>"001110110",
  44432=>"001011111",
  44433=>"111001000",
  44434=>"111000111",
  44435=>"100100110",
  44436=>"010011110",
  44437=>"011011001",
  44438=>"011010011",
  44439=>"101110111",
  44440=>"001001001",
  44441=>"001101001",
  44442=>"000000111",
  44443=>"001010101",
  44444=>"101111011",
  44445=>"011101111",
  44446=>"000110000",
  44447=>"110000010",
  44448=>"111001010",
  44449=>"111100000",
  44450=>"110100010",
  44451=>"110100100",
  44452=>"111100011",
  44453=>"000110100",
  44454=>"001100101",
  44455=>"010000010",
  44456=>"000010001",
  44457=>"010111111",
  44458=>"010101010",
  44459=>"010000111",
  44460=>"010000010",
  44461=>"011011010",
  44462=>"010110110",
  44463=>"101001001",
  44464=>"101001010",
  44465=>"101001011",
  44466=>"101100100",
  44467=>"011011101",
  44468=>"001001011",
  44469=>"101110010",
  44470=>"001010010",
  44471=>"110101011",
  44472=>"111101101",
  44473=>"101110000",
  44474=>"010001110",
  44475=>"101100011",
  44476=>"011100110",
  44477=>"101110000",
  44478=>"100010100",
  44479=>"000000101",
  44480=>"011001000",
  44481=>"110011010",
  44482=>"111110011",
  44483=>"110101000",
  44484=>"000101000",
  44485=>"111000110",
  44486=>"110111101",
  44487=>"111111001",
  44488=>"101101101",
  44489=>"101001010",
  44490=>"000011011",
  44491=>"111110001",
  44492=>"111011100",
  44493=>"001011111",
  44494=>"100000011",
  44495=>"001101100",
  44496=>"100111000",
  44497=>"010100001",
  44498=>"010111111",
  44499=>"010100010",
  44500=>"100011001",
  44501=>"110001010",
  44502=>"000111101",
  44503=>"001000001",
  44504=>"010100000",
  44505=>"110101011",
  44506=>"111001011",
  44507=>"010011111",
  44508=>"111111110",
  44509=>"000101011",
  44510=>"010000000",
  44511=>"111001010",
  44512=>"011000000",
  44513=>"000001000",
  44514=>"010001010",
  44515=>"010101100",
  44516=>"010010011",
  44517=>"000011111",
  44518=>"000010001",
  44519=>"110111111",
  44520=>"111011011",
  44521=>"000011110",
  44522=>"001111101",
  44523=>"111110000",
  44524=>"011111000",
  44525=>"110111011",
  44526=>"010111101",
  44527=>"001101001",
  44528=>"100000010",
  44529=>"110110111",
  44530=>"111010111",
  44531=>"010111010",
  44532=>"100111001",
  44533=>"001101110",
  44534=>"001100110",
  44535=>"111101001",
  44536=>"101101101",
  44537=>"100000100",
  44538=>"000010001",
  44539=>"010011101",
  44540=>"010000110",
  44541=>"010101110",
  44542=>"001100010",
  44543=>"101110011",
  44544=>"101000010",
  44545=>"111001100",
  44546=>"101011101",
  44547=>"010001000",
  44548=>"010011001",
  44549=>"011100011",
  44550=>"010111000",
  44551=>"101111101",
  44552=>"111111101",
  44553=>"010100101",
  44554=>"100011010",
  44555=>"110111001",
  44556=>"000010100",
  44557=>"000000100",
  44558=>"101100111",
  44559=>"011010111",
  44560=>"010100010",
  44561=>"111101010",
  44562=>"001100100",
  44563=>"010001000",
  44564=>"101000101",
  44565=>"110111101",
  44566=>"010000110",
  44567=>"111111110",
  44568=>"000101010",
  44569=>"011111000",
  44570=>"001110111",
  44571=>"000010100",
  44572=>"001111101",
  44573=>"110110010",
  44574=>"000101010",
  44575=>"000101000",
  44576=>"011110111",
  44577=>"010011001",
  44578=>"111000100",
  44579=>"010110001",
  44580=>"111111101",
  44581=>"110000111",
  44582=>"001011100",
  44583=>"000101010",
  44584=>"000001010",
  44585=>"101010001",
  44586=>"111010110",
  44587=>"001010110",
  44588=>"111110101",
  44589=>"100001001",
  44590=>"001001111",
  44591=>"100011111",
  44592=>"011010010",
  44593=>"001001100",
  44594=>"101000000",
  44595=>"001100101",
  44596=>"111111011",
  44597=>"000000101",
  44598=>"001000101",
  44599=>"010001110",
  44600=>"100101011",
  44601=>"000011010",
  44602=>"010010010",
  44603=>"110000001",
  44604=>"100111110",
  44605=>"010000000",
  44606=>"000000100",
  44607=>"011011001",
  44608=>"011000000",
  44609=>"011100111",
  44610=>"010011001",
  44611=>"010100000",
  44612=>"110011000",
  44613=>"001101111",
  44614=>"110000100",
  44615=>"100100101",
  44616=>"111010010",
  44617=>"111001100",
  44618=>"100101111",
  44619=>"010011010",
  44620=>"010101010",
  44621=>"001010110",
  44622=>"010010001",
  44623=>"101010000",
  44624=>"011011101",
  44625=>"001010110",
  44626=>"010001110",
  44627=>"101100010",
  44628=>"011011100",
  44629=>"101101000",
  44630=>"101011000",
  44631=>"010110011",
  44632=>"010111001",
  44633=>"110110100",
  44634=>"101010001",
  44635=>"011011000",
  44636=>"111101101",
  44637=>"101010011",
  44638=>"000001001",
  44639=>"111010001",
  44640=>"100000000",
  44641=>"010000111",
  44642=>"010011101",
  44643=>"100010000",
  44644=>"110101111",
  44645=>"100010010",
  44646=>"010000000",
  44647=>"011000111",
  44648=>"110010101",
  44649=>"011001101",
  44650=>"100011100",
  44651=>"000001001",
  44652=>"111110000",
  44653=>"111100110",
  44654=>"100100110",
  44655=>"110111011",
  44656=>"111010010",
  44657=>"111101000",
  44658=>"000000001",
  44659=>"011000010",
  44660=>"100011110",
  44661=>"110100111",
  44662=>"100101010",
  44663=>"100100100",
  44664=>"001110001",
  44665=>"111111100",
  44666=>"110110101",
  44667=>"011001011",
  44668=>"100011001",
  44669=>"000010011",
  44670=>"110011000",
  44671=>"000010011",
  44672=>"100101110",
  44673=>"110111101",
  44674=>"011111011",
  44675=>"010001100",
  44676=>"011010000",
  44677=>"010001110",
  44678=>"100010101",
  44679=>"111101100",
  44680=>"011011000",
  44681=>"110011111",
  44682=>"110010001",
  44683=>"011100100",
  44684=>"111110100",
  44685=>"000101111",
  44686=>"011101111",
  44687=>"010000001",
  44688=>"101110011",
  44689=>"111011011",
  44690=>"111101110",
  44691=>"001011111",
  44692=>"000101111",
  44693=>"011111101",
  44694=>"000011110",
  44695=>"111011110",
  44696=>"001011011",
  44697=>"100000110",
  44698=>"001100101",
  44699=>"011011011",
  44700=>"011111101",
  44701=>"010001110",
  44702=>"011101010",
  44703=>"110011100",
  44704=>"001001011",
  44705=>"001110111",
  44706=>"000110111",
  44707=>"110001000",
  44708=>"001010111",
  44709=>"010100001",
  44710=>"011010101",
  44711=>"001010000",
  44712=>"011100111",
  44713=>"111001100",
  44714=>"011101111",
  44715=>"011001011",
  44716=>"110000000",
  44717=>"100000001",
  44718=>"001100101",
  44719=>"011100010",
  44720=>"110111001",
  44721=>"100110010",
  44722=>"101000100",
  44723=>"010000000",
  44724=>"100000101",
  44725=>"110000011",
  44726=>"101000010",
  44727=>"001100111",
  44728=>"000101011",
  44729=>"111001100",
  44730=>"000001001",
  44731=>"000000001",
  44732=>"110110101",
  44733=>"011111011",
  44734=>"110001000",
  44735=>"111110010",
  44736=>"000011011",
  44737=>"110000100",
  44738=>"001011101",
  44739=>"111111110",
  44740=>"101110101",
  44741=>"110011111",
  44742=>"111000100",
  44743=>"111010001",
  44744=>"111011110",
  44745=>"010101100",
  44746=>"100110101",
  44747=>"101111100",
  44748=>"010001011",
  44749=>"010011001",
  44750=>"001000111",
  44751=>"111111001",
  44752=>"101110001",
  44753=>"000011001",
  44754=>"011110100",
  44755=>"010001111",
  44756=>"000100101",
  44757=>"000010111",
  44758=>"000001011",
  44759=>"111010101",
  44760=>"100101110",
  44761=>"111111110",
  44762=>"011010001",
  44763=>"000010010",
  44764=>"111010001",
  44765=>"000010101",
  44766=>"001111011",
  44767=>"101101111",
  44768=>"110110001",
  44769=>"001000000",
  44770=>"001010011",
  44771=>"101001010",
  44772=>"011001011",
  44773=>"011010000",
  44774=>"101010100",
  44775=>"110001110",
  44776=>"011000010",
  44777=>"000110010",
  44778=>"111110111",
  44779=>"101010101",
  44780=>"010001111",
  44781=>"010110001",
  44782=>"100111111",
  44783=>"010011001",
  44784=>"010100011",
  44785=>"000000100",
  44786=>"100111111",
  44787=>"001011001",
  44788=>"111101101",
  44789=>"000011111",
  44790=>"101011110",
  44791=>"101011111",
  44792=>"100001111",
  44793=>"100010101",
  44794=>"001011111",
  44795=>"011011000",
  44796=>"110001010",
  44797=>"101010011",
  44798=>"111110010",
  44799=>"100100110",
  44800=>"011100101",
  44801=>"101100010",
  44802=>"100100000",
  44803=>"010101110",
  44804=>"110111001",
  44805=>"111001001",
  44806=>"101100111",
  44807=>"000001100",
  44808=>"011001101",
  44809=>"110110001",
  44810=>"111000101",
  44811=>"111001100",
  44812=>"011110111",
  44813=>"101110101",
  44814=>"100111100",
  44815=>"000010111",
  44816=>"011111101",
  44817=>"010010001",
  44818=>"110100111",
  44819=>"001100101",
  44820=>"100011100",
  44821=>"111001011",
  44822=>"100011110",
  44823=>"000110100",
  44824=>"111011111",
  44825=>"111111010",
  44826=>"111110011",
  44827=>"111100100",
  44828=>"101010110",
  44829=>"111010010",
  44830=>"011000000",
  44831=>"100111101",
  44832=>"000011011",
  44833=>"100101000",
  44834=>"110100000",
  44835=>"101110111",
  44836=>"101011100",
  44837=>"110001100",
  44838=>"000100111",
  44839=>"011111111",
  44840=>"100111110",
  44841=>"100011010",
  44842=>"000001011",
  44843=>"000110110",
  44844=>"101010001",
  44845=>"000011001",
  44846=>"001101011",
  44847=>"010001011",
  44848=>"011011101",
  44849=>"101010000",
  44850=>"011110001",
  44851=>"101100001",
  44852=>"001010001",
  44853=>"010111011",
  44854=>"010101001",
  44855=>"010100101",
  44856=>"100111100",
  44857=>"011100011",
  44858=>"101001101",
  44859=>"110101110",
  44860=>"001110010",
  44861=>"110100101",
  44862=>"010001000",
  44863=>"000011011",
  44864=>"110011111",
  44865=>"111101110",
  44866=>"111011000",
  44867=>"001110110",
  44868=>"100000011",
  44869=>"010100111",
  44870=>"001100010",
  44871=>"111010000",
  44872=>"100011110",
  44873=>"001011010",
  44874=>"001010010",
  44875=>"000100110",
  44876=>"110111111",
  44877=>"110100000",
  44878=>"111101101",
  44879=>"010001101",
  44880=>"101001011",
  44881=>"001000111",
  44882=>"111001010",
  44883=>"011101110",
  44884=>"010011011",
  44885=>"101001101",
  44886=>"001111010",
  44887=>"000010010",
  44888=>"110101111",
  44889=>"000011100",
  44890=>"000110110",
  44891=>"000100011",
  44892=>"100111111",
  44893=>"010101111",
  44894=>"011011111",
  44895=>"101100010",
  44896=>"010101000",
  44897=>"011101010",
  44898=>"010010110",
  44899=>"110101100",
  44900=>"100010100",
  44901=>"011011010",
  44902=>"111101000",
  44903=>"001011010",
  44904=>"111111001",
  44905=>"010000010",
  44906=>"111111011",
  44907=>"000110111",
  44908=>"101111000",
  44909=>"011011001",
  44910=>"001100000",
  44911=>"100001111",
  44912=>"111001010",
  44913=>"111110011",
  44914=>"111111010",
  44915=>"110001010",
  44916=>"010101010",
  44917=>"010000101",
  44918=>"101110110",
  44919=>"111110100",
  44920=>"111101011",
  44921=>"000001101",
  44922=>"110101001",
  44923=>"100110101",
  44924=>"000011000",
  44925=>"110101100",
  44926=>"101001001",
  44927=>"011010000",
  44928=>"000001101",
  44929=>"101011110",
  44930=>"111101101",
  44931=>"111000001",
  44932=>"000110101",
  44933=>"111111011",
  44934=>"000000000",
  44935=>"111011011",
  44936=>"101111000",
  44937=>"110100110",
  44938=>"111011100",
  44939=>"011000011",
  44940=>"110100100",
  44941=>"010010111",
  44942=>"001101101",
  44943=>"101100011",
  44944=>"011101101",
  44945=>"100011000",
  44946=>"111001000",
  44947=>"101011000",
  44948=>"111001111",
  44949=>"101101010",
  44950=>"000011010",
  44951=>"101011100",
  44952=>"011111101",
  44953=>"011011110",
  44954=>"110010001",
  44955=>"110000011",
  44956=>"110111011",
  44957=>"101101101",
  44958=>"110100110",
  44959=>"011111111",
  44960=>"111111001",
  44961=>"011011111",
  44962=>"111011100",
  44963=>"101000101",
  44964=>"110001101",
  44965=>"001000111",
  44966=>"010101000",
  44967=>"100101110",
  44968=>"100111011",
  44969=>"000111100",
  44970=>"000101100",
  44971=>"001110001",
  44972=>"001010100",
  44973=>"000001000",
  44974=>"110000100",
  44975=>"000011110",
  44976=>"001011000",
  44977=>"000000101",
  44978=>"101100001",
  44979=>"001111100",
  44980=>"011110110",
  44981=>"100010011",
  44982=>"010000110",
  44983=>"000011010",
  44984=>"000011111",
  44985=>"010000100",
  44986=>"000011011",
  44987=>"110000000",
  44988=>"101111100",
  44989=>"010110000",
  44990=>"100000100",
  44991=>"111100000",
  44992=>"100110010",
  44993=>"100001011",
  44994=>"010100001",
  44995=>"000100011",
  44996=>"000011100",
  44997=>"000011101",
  44998=>"110001101",
  44999=>"100111001",
  45000=>"000001100",
  45001=>"010001111",
  45002=>"011100001",
  45003=>"100001000",
  45004=>"110100111",
  45005=>"101000000",
  45006=>"111110001",
  45007=>"101101011",
  45008=>"010101010",
  45009=>"010010100",
  45010=>"000111111",
  45011=>"011010110",
  45012=>"000011110",
  45013=>"111111011",
  45014=>"100111111",
  45015=>"101011010",
  45016=>"011100000",
  45017=>"001110000",
  45018=>"101110111",
  45019=>"111010011",
  45020=>"110011110",
  45021=>"111010101",
  45022=>"111111001",
  45023=>"100101001",
  45024=>"010000000",
  45025=>"101101011",
  45026=>"101111100",
  45027=>"110100011",
  45028=>"001011001",
  45029=>"011111011",
  45030=>"000000110",
  45031=>"100010000",
  45032=>"011000101",
  45033=>"111100101",
  45034=>"001111001",
  45035=>"111010101",
  45036=>"111110000",
  45037=>"100000100",
  45038=>"000110111",
  45039=>"010111100",
  45040=>"001111111",
  45041=>"101110011",
  45042=>"001000011",
  45043=>"000000100",
  45044=>"010010010",
  45045=>"011001001",
  45046=>"010011011",
  45047=>"111011000",
  45048=>"001011010",
  45049=>"111000110",
  45050=>"101000000",
  45051=>"100011000",
  45052=>"101111000",
  45053=>"101100010",
  45054=>"111101100",
  45055=>"010111111",
  45056=>"101100111",
  45057=>"110001110",
  45058=>"111100000",
  45059=>"011111101",
  45060=>"110011100",
  45061=>"111101100",
  45062=>"111101011",
  45063=>"100000010",
  45064=>"000010011",
  45065=>"010100010",
  45066=>"010011101",
  45067=>"111111011",
  45068=>"000100000",
  45069=>"010101110",
  45070=>"001000101",
  45071=>"100000100",
  45072=>"110011001",
  45073=>"100111010",
  45074=>"010111011",
  45075=>"111000100",
  45076=>"011010101",
  45077=>"111010111",
  45078=>"101011000",
  45079=>"111000111",
  45080=>"010110010",
  45081=>"101101101",
  45082=>"000011010",
  45083=>"110101110",
  45084=>"000101100",
  45085=>"100010001",
  45086=>"001101111",
  45087=>"101110100",
  45088=>"011101100",
  45089=>"110101100",
  45090=>"011001110",
  45091=>"111000110",
  45092=>"011101000",
  45093=>"010111010",
  45094=>"000101101",
  45095=>"001011010",
  45096=>"110100011",
  45097=>"111010001",
  45098=>"100100111",
  45099=>"110110111",
  45100=>"111111111",
  45101=>"010010011",
  45102=>"110100011",
  45103=>"011000101",
  45104=>"111001011",
  45105=>"010000010",
  45106=>"111000001",
  45107=>"001111011",
  45108=>"110000100",
  45109=>"110100110",
  45110=>"111000010",
  45111=>"101111111",
  45112=>"110001001",
  45113=>"111001011",
  45114=>"010100001",
  45115=>"110111110",
  45116=>"000001000",
  45117=>"000101000",
  45118=>"010010110",
  45119=>"111010101",
  45120=>"111110000",
  45121=>"101111101",
  45122=>"010011001",
  45123=>"101001000",
  45124=>"101000011",
  45125=>"111111100",
  45126=>"001101100",
  45127=>"011101000",
  45128=>"101000010",
  45129=>"000100100",
  45130=>"011011011",
  45131=>"100111101",
  45132=>"010101100",
  45133=>"110111111",
  45134=>"000001101",
  45135=>"000001101",
  45136=>"111101100",
  45137=>"101010101",
  45138=>"110000011",
  45139=>"010001010",
  45140=>"101101111",
  45141=>"001101110",
  45142=>"001110110",
  45143=>"000100001",
  45144=>"110010011",
  45145=>"110011011",
  45146=>"001101010",
  45147=>"001000101",
  45148=>"001000001",
  45149=>"110110010",
  45150=>"010111010",
  45151=>"100101000",
  45152=>"000110110",
  45153=>"001101010",
  45154=>"111010100",
  45155=>"000111001",
  45156=>"001001000",
  45157=>"111101100",
  45158=>"110101010",
  45159=>"001110111",
  45160=>"010010011",
  45161=>"100000101",
  45162=>"000111010",
  45163=>"100000011",
  45164=>"101100101",
  45165=>"001110111",
  45166=>"000010111",
  45167=>"111100010",
  45168=>"011100001",
  45169=>"110010101",
  45170=>"111100111",
  45171=>"111001101",
  45172=>"001100001",
  45173=>"000001111",
  45174=>"111101001",
  45175=>"101100001",
  45176=>"100110100",
  45177=>"011011001",
  45178=>"100101110",
  45179=>"000111111",
  45180=>"101111100",
  45181=>"000001011",
  45182=>"011011101",
  45183=>"000111110",
  45184=>"110111111",
  45185=>"111000101",
  45186=>"110100110",
  45187=>"111101000",
  45188=>"110100101",
  45189=>"100011000",
  45190=>"101001110",
  45191=>"100100010",
  45192=>"100111100",
  45193=>"011000000",
  45194=>"010001100",
  45195=>"100100010",
  45196=>"100010001",
  45197=>"101000110",
  45198=>"100111111",
  45199=>"000001100",
  45200=>"010000110",
  45201=>"111001001",
  45202=>"011110000",
  45203=>"101010111",
  45204=>"001100101",
  45205=>"110101011",
  45206=>"000101010",
  45207=>"110101000",
  45208=>"111111101",
  45209=>"100111101",
  45210=>"100110001",
  45211=>"111101110",
  45212=>"100101110",
  45213=>"110001100",
  45214=>"011000100",
  45215=>"110111001",
  45216=>"101010000",
  45217=>"101010111",
  45218=>"010000000",
  45219=>"100111000",
  45220=>"111000001",
  45221=>"100101010",
  45222=>"010010100",
  45223=>"010110010",
  45224=>"100000111",
  45225=>"010100111",
  45226=>"000100011",
  45227=>"001010100",
  45228=>"011101000",
  45229=>"011000110",
  45230=>"100101111",
  45231=>"011100101",
  45232=>"001001000",
  45233=>"010010000",
  45234=>"101011101",
  45235=>"011000000",
  45236=>"001001101",
  45237=>"000000000",
  45238=>"000010000",
  45239=>"001010000",
  45240=>"000101011",
  45241=>"100101001",
  45242=>"101000110",
  45243=>"000001101",
  45244=>"001001011",
  45245=>"000010101",
  45246=>"011000110",
  45247=>"001000010",
  45248=>"100011110",
  45249=>"100110011",
  45250=>"010101110",
  45251=>"111001111",
  45252=>"000101011",
  45253=>"101010001",
  45254=>"000000001",
  45255=>"101111100",
  45256=>"110010011",
  45257=>"101011101",
  45258=>"000101010",
  45259=>"011011100",
  45260=>"100110000",
  45261=>"110111111",
  45262=>"011100011",
  45263=>"101011011",
  45264=>"001100010",
  45265=>"101011101",
  45266=>"010111110",
  45267=>"110000000",
  45268=>"101000111",
  45269=>"110111110",
  45270=>"001111101",
  45271=>"100000001",
  45272=>"100011100",
  45273=>"000111001",
  45274=>"011011011",
  45275=>"101011001",
  45276=>"000100010",
  45277=>"110001010",
  45278=>"111001000",
  45279=>"110110110",
  45280=>"001011000",
  45281=>"011100110",
  45282=>"110111001",
  45283=>"100101101",
  45284=>"110111000",
  45285=>"100010101",
  45286=>"010000100",
  45287=>"101010001",
  45288=>"010000000",
  45289=>"111010011",
  45290=>"111000101",
  45291=>"100101111",
  45292=>"000001110",
  45293=>"100011011",
  45294=>"100001110",
  45295=>"110010001",
  45296=>"111111100",
  45297=>"101110100",
  45298=>"100111001",
  45299=>"010001111",
  45300=>"010001001",
  45301=>"010100000",
  45302=>"100110100",
  45303=>"001001110",
  45304=>"100110011",
  45305=>"111110101",
  45306=>"101111100",
  45307=>"000000100",
  45308=>"101000010",
  45309=>"010001001",
  45310=>"001010101",
  45311=>"110010100",
  45312=>"010111100",
  45313=>"111010001",
  45314=>"111011111",
  45315=>"001100110",
  45316=>"111000101",
  45317=>"111100001",
  45318=>"011100110",
  45319=>"001101001",
  45320=>"000011011",
  45321=>"110101011",
  45322=>"001010000",
  45323=>"100110110",
  45324=>"001011001",
  45325=>"011010001",
  45326=>"011001011",
  45327=>"100110101",
  45328=>"011001110",
  45329=>"111110001",
  45330=>"110111111",
  45331=>"100101100",
  45332=>"001101110",
  45333=>"110111001",
  45334=>"010100100",
  45335=>"101011111",
  45336=>"000101010",
  45337=>"001101010",
  45338=>"011011111",
  45339=>"110100101",
  45340=>"100000001",
  45341=>"100100010",
  45342=>"011100110",
  45343=>"011110000",
  45344=>"100011110",
  45345=>"011000010",
  45346=>"110000001",
  45347=>"000000100",
  45348=>"001011011",
  45349=>"111101111",
  45350=>"111110100",
  45351=>"011000011",
  45352=>"011001111",
  45353=>"010010011",
  45354=>"100000010",
  45355=>"100000001",
  45356=>"101010100",
  45357=>"011000101",
  45358=>"000110001",
  45359=>"000110000",
  45360=>"100101100",
  45361=>"110101111",
  45362=>"011001111",
  45363=>"101110011",
  45364=>"001000111",
  45365=>"010100010",
  45366=>"000010000",
  45367=>"001110111",
  45368=>"000110011",
  45369=>"000110110",
  45370=>"011010111",
  45371=>"111011101",
  45372=>"010110101",
  45373=>"100101001",
  45374=>"100110000",
  45375=>"001100101",
  45376=>"110111111",
  45377=>"100010110",
  45378=>"110101010",
  45379=>"011011100",
  45380=>"011001011",
  45381=>"000000010",
  45382=>"100001000",
  45383=>"100101000",
  45384=>"011101010",
  45385=>"100000011",
  45386=>"111011001",
  45387=>"000110110",
  45388=>"111111010",
  45389=>"110011110",
  45390=>"001010001",
  45391=>"110100111",
  45392=>"001111100",
  45393=>"110100000",
  45394=>"000001111",
  45395=>"111111101",
  45396=>"001111111",
  45397=>"011000000",
  45398=>"010111111",
  45399=>"000100110",
  45400=>"011010101",
  45401=>"011111011",
  45402=>"000011111",
  45403=>"101101000",
  45404=>"101010010",
  45405=>"001100001",
  45406=>"111111101",
  45407=>"010101000",
  45408=>"111111100",
  45409=>"111110011",
  45410=>"110011001",
  45411=>"111111100",
  45412=>"111000101",
  45413=>"100111100",
  45414=>"010001100",
  45415=>"101111010",
  45416=>"000001110",
  45417=>"111100011",
  45418=>"100010010",
  45419=>"100011101",
  45420=>"011000100",
  45421=>"001000000",
  45422=>"011111111",
  45423=>"001010011",
  45424=>"010101101",
  45425=>"000011100",
  45426=>"101000111",
  45427=>"010101001",
  45428=>"110111000",
  45429=>"101011000",
  45430=>"011001011",
  45431=>"011011011",
  45432=>"111011111",
  45433=>"001011011",
  45434=>"100000000",
  45435=>"001011000",
  45436=>"110111000",
  45437=>"000100011",
  45438=>"101001011",
  45439=>"111010000",
  45440=>"010011011",
  45441=>"101001000",
  45442=>"011101100",
  45443=>"011110000",
  45444=>"010001111",
  45445=>"000001000",
  45446=>"011000010",
  45447=>"100000000",
  45448=>"010100011",
  45449=>"100100011",
  45450=>"111011111",
  45451=>"011001111",
  45452=>"110010100",
  45453=>"110011100",
  45454=>"011111101",
  45455=>"011111010",
  45456=>"101001011",
  45457=>"011000011",
  45458=>"011111010",
  45459=>"101111111",
  45460=>"001100110",
  45461=>"010110110",
  45462=>"001100101",
  45463=>"001011111",
  45464=>"011110100",
  45465=>"100100110",
  45466=>"000111011",
  45467=>"011010000",
  45468=>"111001001",
  45469=>"000001001",
  45470=>"010010110",
  45471=>"110000110",
  45472=>"001000101",
  45473=>"110100101",
  45474=>"111110000",
  45475=>"110100111",
  45476=>"100000100",
  45477=>"101111111",
  45478=>"001010011",
  45479=>"100000000",
  45480=>"101000000",
  45481=>"111000000",
  45482=>"010000100",
  45483=>"011010011",
  45484=>"011011001",
  45485=>"001010000",
  45486=>"000101110",
  45487=>"110001101",
  45488=>"000011000",
  45489=>"000001100",
  45490=>"011100101",
  45491=>"001000101",
  45492=>"111111000",
  45493=>"011010100",
  45494=>"111101111",
  45495=>"000011011",
  45496=>"000001110",
  45497=>"010000000",
  45498=>"101100101",
  45499=>"101011000",
  45500=>"100001100",
  45501=>"110001011",
  45502=>"000011100",
  45503=>"010010110",
  45504=>"111100001",
  45505=>"110111010",
  45506=>"101011100",
  45507=>"010011010",
  45508=>"010011011",
  45509=>"110011110",
  45510=>"011111000",
  45511=>"101111110",
  45512=>"101011100",
  45513=>"000101001",
  45514=>"001001001",
  45515=>"011001001",
  45516=>"011001110",
  45517=>"100000111",
  45518=>"101101010",
  45519=>"000100110",
  45520=>"010100000",
  45521=>"000111100",
  45522=>"010010011",
  45523=>"001110100",
  45524=>"100011101",
  45525=>"010010000",
  45526=>"100011000",
  45527=>"001001110",
  45528=>"000100001",
  45529=>"111110111",
  45530=>"001100110",
  45531=>"101110000",
  45532=>"111101110",
  45533=>"110000011",
  45534=>"110101111",
  45535=>"100011011",
  45536=>"001000101",
  45537=>"010101000",
  45538=>"101100110",
  45539=>"011010100",
  45540=>"001101100",
  45541=>"101111100",
  45542=>"011010000",
  45543=>"011111110",
  45544=>"010110000",
  45545=>"011010100",
  45546=>"000111101",
  45547=>"010100110",
  45548=>"100111010",
  45549=>"011001001",
  45550=>"011001001",
  45551=>"000110001",
  45552=>"011111001",
  45553=>"011101000",
  45554=>"011000000",
  45555=>"011010001",
  45556=>"101100001",
  45557=>"111000001",
  45558=>"010101011",
  45559=>"111010100",
  45560=>"110010101",
  45561=>"011011000",
  45562=>"011111110",
  45563=>"011000100",
  45564=>"000011011",
  45565=>"000001001",
  45566=>"000111000",
  45567=>"110011000",
  45568=>"010101001",
  45569=>"110011100",
  45570=>"010100010",
  45571=>"100000000",
  45572=>"101100111",
  45573=>"001110001",
  45574=>"011011111",
  45575=>"000010010",
  45576=>"010000010",
  45577=>"111100001",
  45578=>"110111101",
  45579=>"011111110",
  45580=>"110111001",
  45581=>"100110011",
  45582=>"100000110",
  45583=>"100000011",
  45584=>"101100011",
  45585=>"010111000",
  45586=>"100000001",
  45587=>"101101011",
  45588=>"000000101",
  45589=>"100011101",
  45590=>"011101010",
  45591=>"010100010",
  45592=>"110010110",
  45593=>"100100000",
  45594=>"011011011",
  45595=>"111100000",
  45596=>"010100101",
  45597=>"100101111",
  45598=>"110001111",
  45599=>"110001100",
  45600=>"110111000",
  45601=>"100111011",
  45602=>"000100011",
  45603=>"100000001",
  45604=>"010010011",
  45605=>"110011111",
  45606=>"011111010",
  45607=>"000101000",
  45608=>"010110101",
  45609=>"001011010",
  45610=>"110110011",
  45611=>"010100110",
  45612=>"111101000",
  45613=>"000001000",
  45614=>"110010000",
  45615=>"100101111",
  45616=>"000001010",
  45617=>"101010100",
  45618=>"010100011",
  45619=>"100100010",
  45620=>"010100000",
  45621=>"111110101",
  45622=>"110110011",
  45623=>"010000010",
  45624=>"111101100",
  45625=>"101110101",
  45626=>"010010110",
  45627=>"101011100",
  45628=>"110111111",
  45629=>"000010001",
  45630=>"111000011",
  45631=>"101001111",
  45632=>"110111011",
  45633=>"001010111",
  45634=>"110111011",
  45635=>"001100101",
  45636=>"000011100",
  45637=>"000100011",
  45638=>"001100111",
  45639=>"100111101",
  45640=>"000011111",
  45641=>"010100110",
  45642=>"010011011",
  45643=>"101000110",
  45644=>"001011011",
  45645=>"100010111",
  45646=>"010100010",
  45647=>"110100001",
  45648=>"010111110",
  45649=>"111111100",
  45650=>"011110011",
  45651=>"000100001",
  45652=>"101110101",
  45653=>"111011000",
  45654=>"111100101",
  45655=>"000000101",
  45656=>"010101110",
  45657=>"110100110",
  45658=>"101011011",
  45659=>"011001111",
  45660=>"010000101",
  45661=>"110010110",
  45662=>"101001010",
  45663=>"111101101",
  45664=>"001111100",
  45665=>"010010010",
  45666=>"010011100",
  45667=>"100101011",
  45668=>"011011110",
  45669=>"111011010",
  45670=>"011110001",
  45671=>"100010001",
  45672=>"111010010",
  45673=>"010110111",
  45674=>"000000101",
  45675=>"001000110",
  45676=>"101000001",
  45677=>"001101101",
  45678=>"110001011",
  45679=>"001001000",
  45680=>"100011011",
  45681=>"101101011",
  45682=>"111110010",
  45683=>"110001011",
  45684=>"111110000",
  45685=>"110001001",
  45686=>"000001100",
  45687=>"101000110",
  45688=>"101000111",
  45689=>"011000111",
  45690=>"001001000",
  45691=>"110111000",
  45692=>"111000011",
  45693=>"011100111",
  45694=>"010101011",
  45695=>"100100011",
  45696=>"011100100",
  45697=>"101011001",
  45698=>"101101000",
  45699=>"111111111",
  45700=>"101110000",
  45701=>"011010100",
  45702=>"101110111",
  45703=>"010010000",
  45704=>"111110111",
  45705=>"100101000",
  45706=>"011100001",
  45707=>"011101000",
  45708=>"010010001",
  45709=>"001110000",
  45710=>"101000000",
  45711=>"100110100",
  45712=>"101011000",
  45713=>"001001111",
  45714=>"010111101",
  45715=>"001010111",
  45716=>"111010010",
  45717=>"100001000",
  45718=>"001001010",
  45719=>"010110011",
  45720=>"011000000",
  45721=>"111001110",
  45722=>"110011010",
  45723=>"111101111",
  45724=>"000010111",
  45725=>"010101001",
  45726=>"010000100",
  45727=>"011100011",
  45728=>"001010011",
  45729=>"010101000",
  45730=>"000000010",
  45731=>"000011111",
  45732=>"000110000",
  45733=>"000010111",
  45734=>"001001001",
  45735=>"100001000",
  45736=>"011010111",
  45737=>"101010100",
  45738=>"100001100",
  45739=>"010101111",
  45740=>"100101101",
  45741=>"101010110",
  45742=>"001010110",
  45743=>"100001101",
  45744=>"001011111",
  45745=>"110001111",
  45746=>"001101110",
  45747=>"000110100",
  45748=>"100101101",
  45749=>"100101100",
  45750=>"111100001",
  45751=>"100110111",
  45752=>"101101010",
  45753=>"100101100",
  45754=>"100110100",
  45755=>"011100110",
  45756=>"111110110",
  45757=>"000110000",
  45758=>"101010110",
  45759=>"010010001",
  45760=>"000010000",
  45761=>"011110011",
  45762=>"100001010",
  45763=>"111011000",
  45764=>"111001100",
  45765=>"110000101",
  45766=>"010100011",
  45767=>"110010010",
  45768=>"111110101",
  45769=>"110000000",
  45770=>"011001110",
  45771=>"110011111",
  45772=>"001011111",
  45773=>"100001111",
  45774=>"001100001",
  45775=>"000100100",
  45776=>"001110011",
  45777=>"110001000",
  45778=>"010010011",
  45779=>"010100100",
  45780=>"101111101",
  45781=>"100101000",
  45782=>"111001001",
  45783=>"111100111",
  45784=>"011011000",
  45785=>"101010001",
  45786=>"101101110",
  45787=>"100001000",
  45788=>"111001101",
  45789=>"001100100",
  45790=>"010010011",
  45791=>"001100000",
  45792=>"000101100",
  45793=>"100000011",
  45794=>"111100010",
  45795=>"000000001",
  45796=>"001000100",
  45797=>"011001000",
  45798=>"010011111",
  45799=>"110010000",
  45800=>"001100111",
  45801=>"111111100",
  45802=>"111101011",
  45803=>"001110100",
  45804=>"110101111",
  45805=>"000001000",
  45806=>"100000001",
  45807=>"110111001",
  45808=>"001101010",
  45809=>"110010001",
  45810=>"011001000",
  45811=>"000001101",
  45812=>"000010100",
  45813=>"101000011",
  45814=>"111110100",
  45815=>"010001111",
  45816=>"011001110",
  45817=>"001110110",
  45818=>"100100000",
  45819=>"000101110",
  45820=>"011011111",
  45821=>"001111110",
  45822=>"000000111",
  45823=>"000000100",
  45824=>"101101010",
  45825=>"010110100",
  45826=>"010100101",
  45827=>"100110111",
  45828=>"011111101",
  45829=>"111011011",
  45830=>"110010000",
  45831=>"101011100",
  45832=>"101000000",
  45833=>"111100110",
  45834=>"010101010",
  45835=>"101010010",
  45836=>"101110010",
  45837=>"010011100",
  45838=>"001100111",
  45839=>"101111111",
  45840=>"111000011",
  45841=>"011000111",
  45842=>"110100100",
  45843=>"111011111",
  45844=>"101110111",
  45845=>"110110100",
  45846=>"000010111",
  45847=>"011100010",
  45848=>"000001101",
  45849=>"101001100",
  45850=>"110111011",
  45851=>"101001110",
  45852=>"001101111",
  45853=>"100000010",
  45854=>"101100100",
  45855=>"011001000",
  45856=>"111110010",
  45857=>"010001000",
  45858=>"010000011",
  45859=>"011011010",
  45860=>"010111000",
  45861=>"101011000",
  45862=>"101101111",
  45863=>"010100011",
  45864=>"010111011",
  45865=>"000001011",
  45866=>"000110010",
  45867=>"010111011",
  45868=>"011001000",
  45869=>"001110101",
  45870=>"001001000",
  45871=>"110011111",
  45872=>"000010001",
  45873=>"000000011",
  45874=>"101011011",
  45875=>"000101010",
  45876=>"101011010",
  45877=>"111010111",
  45878=>"111110011",
  45879=>"110001110",
  45880=>"110000001",
  45881=>"010000001",
  45882=>"001101010",
  45883=>"000101100",
  45884=>"001101011",
  45885=>"000011010",
  45886=>"001100100",
  45887=>"011010110",
  45888=>"010000000",
  45889=>"101101110",
  45890=>"110010100",
  45891=>"101000011",
  45892=>"111110000",
  45893=>"100101001",
  45894=>"000000000",
  45895=>"111011011",
  45896=>"100011011",
  45897=>"100110100",
  45898=>"001011001",
  45899=>"000101100",
  45900=>"000001011",
  45901=>"011110100",
  45902=>"100001100",
  45903=>"100011010",
  45904=>"000111001",
  45905=>"100101000",
  45906=>"000001100",
  45907=>"001110000",
  45908=>"110101011",
  45909=>"100101001",
  45910=>"100111100",
  45911=>"111001101",
  45912=>"001111011",
  45913=>"100110111",
  45914=>"110011111",
  45915=>"010100100",
  45916=>"000000001",
  45917=>"101110111",
  45918=>"011010011",
  45919=>"100001001",
  45920=>"010010110",
  45921=>"000111001",
  45922=>"000100110",
  45923=>"001101110",
  45924=>"011010000",
  45925=>"110110011",
  45926=>"010101101",
  45927=>"011110010",
  45928=>"111110000",
  45929=>"010000000",
  45930=>"011000100",
  45931=>"000010011",
  45932=>"110000000",
  45933=>"001010110",
  45934=>"010010100",
  45935=>"101111010",
  45936=>"000110110",
  45937=>"010111101",
  45938=>"111010010",
  45939=>"010000111",
  45940=>"101010001",
  45941=>"110010001",
  45942=>"000000110",
  45943=>"101100000",
  45944=>"101100110",
  45945=>"100100011",
  45946=>"010000000",
  45947=>"001000100",
  45948=>"010010111",
  45949=>"111100101",
  45950=>"001010000",
  45951=>"010100100",
  45952=>"111111001",
  45953=>"100001111",
  45954=>"111011101",
  45955=>"111011101",
  45956=>"111100100",
  45957=>"011110010",
  45958=>"100011011",
  45959=>"011100011",
  45960=>"000110001",
  45961=>"111111001",
  45962=>"000110001",
  45963=>"101110111",
  45964=>"100111110",
  45965=>"000101010",
  45966=>"000011101",
  45967=>"010010000",
  45968=>"010000001",
  45969=>"111101101",
  45970=>"100000100",
  45971=>"000000101",
  45972=>"110111000",
  45973=>"100101110",
  45974=>"001101000",
  45975=>"000100011",
  45976=>"010001100",
  45977=>"000001110",
  45978=>"100101001",
  45979=>"001010111",
  45980=>"010110100",
  45981=>"101111000",
  45982=>"010111111",
  45983=>"001110000",
  45984=>"010010000",
  45985=>"000010111",
  45986=>"111011100",
  45987=>"110100011",
  45988=>"000100011",
  45989=>"011010001",
  45990=>"110100000",
  45991=>"000110000",
  45992=>"010000000",
  45993=>"011010110",
  45994=>"110011010",
  45995=>"011101101",
  45996=>"000111010",
  45997=>"011100010",
  45998=>"101101101",
  45999=>"010100011",
  46000=>"101000100",
  46001=>"101011010",
  46002=>"100100110",
  46003=>"110110101",
  46004=>"011010111",
  46005=>"110111001",
  46006=>"011111110",
  46007=>"001100101",
  46008=>"111101000",
  46009=>"111010110",
  46010=>"101001101",
  46011=>"101011000",
  46012=>"111100000",
  46013=>"111000011",
  46014=>"101001011",
  46015=>"110001101",
  46016=>"100011000",
  46017=>"100000011",
  46018=>"001101010",
  46019=>"100110110",
  46020=>"111001010",
  46021=>"100101011",
  46022=>"100110010",
  46023=>"010101010",
  46024=>"010110100",
  46025=>"010010010",
  46026=>"111101011",
  46027=>"101000110",
  46028=>"100000101",
  46029=>"110010011",
  46030=>"100100011",
  46031=>"100100010",
  46032=>"101100001",
  46033=>"000100001",
  46034=>"101010111",
  46035=>"111000110",
  46036=>"111100101",
  46037=>"001011011",
  46038=>"010100001",
  46039=>"111101110",
  46040=>"110100011",
  46041=>"011011110",
  46042=>"111111010",
  46043=>"010011000",
  46044=>"101010010",
  46045=>"101101110",
  46046=>"001101111",
  46047=>"011100101",
  46048=>"000101101",
  46049=>"000100111",
  46050=>"100000010",
  46051=>"001010001",
  46052=>"011100110",
  46053=>"000000101",
  46054=>"111111111",
  46055=>"001100101",
  46056=>"110000010",
  46057=>"101010110",
  46058=>"001000101",
  46059=>"111001110",
  46060=>"001111101",
  46061=>"011011010",
  46062=>"111001001",
  46063=>"101011111",
  46064=>"101111010",
  46065=>"000011001",
  46066=>"100000000",
  46067=>"001100111",
  46068=>"111011011",
  46069=>"111000100",
  46070=>"011010010",
  46071=>"000000100",
  46072=>"001000100",
  46073=>"001111010",
  46074=>"100111001",
  46075=>"100111011",
  46076=>"110010101",
  46077=>"011101100",
  46078=>"111001111",
  46079=>"000000100",
  46080=>"111100001",
  46081=>"111000110",
  46082=>"000101011",
  46083=>"010010100",
  46084=>"000100101",
  46085=>"101011000",
  46086=>"000101011",
  46087=>"011110101",
  46088=>"011011110",
  46089=>"111111011",
  46090=>"010101000",
  46091=>"111001001",
  46092=>"010101100",
  46093=>"100001110",
  46094=>"100100110",
  46095=>"000110110",
  46096=>"100010001",
  46097=>"111000010",
  46098=>"110000011",
  46099=>"000100100",
  46100=>"000001111",
  46101=>"001000000",
  46102=>"100011011",
  46103=>"100000001",
  46104=>"001001011",
  46105=>"011101011",
  46106=>"011001001",
  46107=>"111100100",
  46108=>"101011010",
  46109=>"110010001",
  46110=>"100011000",
  46111=>"000001101",
  46112=>"111100100",
  46113=>"000110100",
  46114=>"100110000",
  46115=>"000110010",
  46116=>"000101100",
  46117=>"011011101",
  46118=>"110011001",
  46119=>"100111000",
  46120=>"000100011",
  46121=>"010011110",
  46122=>"101010110",
  46123=>"000000110",
  46124=>"001111111",
  46125=>"101011100",
  46126=>"001000110",
  46127=>"000100010",
  46128=>"011100000",
  46129=>"000100111",
  46130=>"101100010",
  46131=>"100001101",
  46132=>"110100010",
  46133=>"100010010",
  46134=>"000011001",
  46135=>"010010010",
  46136=>"111000001",
  46137=>"001101011",
  46138=>"011001100",
  46139=>"110000101",
  46140=>"011000100",
  46141=>"101011001",
  46142=>"000101000",
  46143=>"001001001",
  46144=>"001010110",
  46145=>"000000001",
  46146=>"101111110",
  46147=>"010010010",
  46148=>"011000100",
  46149=>"101110111",
  46150=>"010110100",
  46151=>"001111101",
  46152=>"110000000",
  46153=>"111110010",
  46154=>"010001000",
  46155=>"010100101",
  46156=>"001001010",
  46157=>"010110000",
  46158=>"110110001",
  46159=>"101010010",
  46160=>"011000110",
  46161=>"011110001",
  46162=>"010101110",
  46163=>"101101111",
  46164=>"100010111",
  46165=>"111001100",
  46166=>"110111101",
  46167=>"011010001",
  46168=>"001100111",
  46169=>"010100101",
  46170=>"010001110",
  46171=>"100100000",
  46172=>"110001111",
  46173=>"010101100",
  46174=>"100101111",
  46175=>"001111111",
  46176=>"111110000",
  46177=>"100010011",
  46178=>"011101011",
  46179=>"011010001",
  46180=>"000111111",
  46181=>"001111001",
  46182=>"111001100",
  46183=>"001011110",
  46184=>"000001010",
  46185=>"101111001",
  46186=>"000101001",
  46187=>"000110101",
  46188=>"000110000",
  46189=>"001101010",
  46190=>"001001010",
  46191=>"010001111",
  46192=>"000000000",
  46193=>"100010111",
  46194=>"000010011",
  46195=>"000100111",
  46196=>"011111111",
  46197=>"111001100",
  46198=>"111110100",
  46199=>"100011001",
  46200=>"101011111",
  46201=>"000011001",
  46202=>"000011100",
  46203=>"101001001",
  46204=>"011011000",
  46205=>"001100010",
  46206=>"110101001",
  46207=>"111001000",
  46208=>"110111000",
  46209=>"100101001",
  46210=>"110001110",
  46211=>"000101001",
  46212=>"110001000",
  46213=>"110110000",
  46214=>"001000001",
  46215=>"100000111",
  46216=>"010010100",
  46217=>"001011010",
  46218=>"000011100",
  46219=>"101010001",
  46220=>"110011100",
  46221=>"111100101",
  46222=>"111111000",
  46223=>"111110110",
  46224=>"011000010",
  46225=>"010001101",
  46226=>"011110000",
  46227=>"111101000",
  46228=>"010001100",
  46229=>"111001010",
  46230=>"100110010",
  46231=>"001110101",
  46232=>"110010110",
  46233=>"101100001",
  46234=>"000110001",
  46235=>"011001000",
  46236=>"100110111",
  46237=>"111000000",
  46238=>"000000001",
  46239=>"100111111",
  46240=>"010100111",
  46241=>"011000111",
  46242=>"001010100",
  46243=>"011000001",
  46244=>"110000010",
  46245=>"110010111",
  46246=>"011011111",
  46247=>"001101001",
  46248=>"010001001",
  46249=>"100000000",
  46250=>"100100100",
  46251=>"101000101",
  46252=>"111001111",
  46253=>"110110100",
  46254=>"110111101",
  46255=>"110100011",
  46256=>"101111100",
  46257=>"010001111",
  46258=>"001001010",
  46259=>"101100000",
  46260=>"110001011",
  46261=>"001110101",
  46262=>"011001011",
  46263=>"101001001",
  46264=>"111111011",
  46265=>"111000110",
  46266=>"000000000",
  46267=>"101100000",
  46268=>"011100001",
  46269=>"011001001",
  46270=>"101010000",
  46271=>"010111001",
  46272=>"111001001",
  46273=>"110011000",
  46274=>"000111111",
  46275=>"101100001",
  46276=>"000000001",
  46277=>"001010000",
  46278=>"100001111",
  46279=>"000000001",
  46280=>"010011011",
  46281=>"101000100",
  46282=>"001011110",
  46283=>"001010000",
  46284=>"101010010",
  46285=>"001101111",
  46286=>"001000101",
  46287=>"111010100",
  46288=>"101010110",
  46289=>"100000011",
  46290=>"010111111",
  46291=>"001000111",
  46292=>"001111100",
  46293=>"000100001",
  46294=>"011101010",
  46295=>"001000101",
  46296=>"110010110",
  46297=>"110010101",
  46298=>"110011000",
  46299=>"001000010",
  46300=>"101011000",
  46301=>"101010000",
  46302=>"101001111",
  46303=>"000111101",
  46304=>"011111001",
  46305=>"001001100",
  46306=>"100101111",
  46307=>"111110101",
  46308=>"111001101",
  46309=>"100010101",
  46310=>"011110001",
  46311=>"000111010",
  46312=>"011111110",
  46313=>"100100011",
  46314=>"000000101",
  46315=>"111100001",
  46316=>"001011110",
  46317=>"110100111",
  46318=>"101100001",
  46319=>"110110110",
  46320=>"101111001",
  46321=>"010011000",
  46322=>"010010111",
  46323=>"101010111",
  46324=>"101111110",
  46325=>"111011110",
  46326=>"001100000",
  46327=>"001011100",
  46328=>"000010011",
  46329=>"111110110",
  46330=>"111100111",
  46331=>"001001011",
  46332=>"100100001",
  46333=>"010110111",
  46334=>"001010011",
  46335=>"001101010",
  46336=>"101011000",
  46337=>"010101111",
  46338=>"101110100",
  46339=>"010100011",
  46340=>"110100111",
  46341=>"010001100",
  46342=>"111100110",
  46343=>"010111101",
  46344=>"101110111",
  46345=>"101100000",
  46346=>"100100101",
  46347=>"010010000",
  46348=>"000101101",
  46349=>"011011100",
  46350=>"110000011",
  46351=>"010001101",
  46352=>"011111100",
  46353=>"100010101",
  46354=>"100100000",
  46355=>"011111110",
  46356=>"101111011",
  46357=>"001100010",
  46358=>"001001101",
  46359=>"000111101",
  46360=>"111011011",
  46361=>"001101001",
  46362=>"001101001",
  46363=>"010101011",
  46364=>"011101010",
  46365=>"010010011",
  46366=>"011111110",
  46367=>"001000101",
  46368=>"110111001",
  46369=>"000000111",
  46370=>"101100100",
  46371=>"000010110",
  46372=>"010000000",
  46373=>"000011011",
  46374=>"010000100",
  46375=>"101011011",
  46376=>"000000110",
  46377=>"010010011",
  46378=>"000100001",
  46379=>"111011000",
  46380=>"101000110",
  46381=>"111001010",
  46382=>"111010011",
  46383=>"100100101",
  46384=>"110000110",
  46385=>"110000110",
  46386=>"111110110",
  46387=>"000100000",
  46388=>"000000001",
  46389=>"101100110",
  46390=>"111010111",
  46391=>"101010111",
  46392=>"000000110",
  46393=>"110111111",
  46394=>"110110111",
  46395=>"100011001",
  46396=>"000110001",
  46397=>"110110001",
  46398=>"000010100",
  46399=>"110000100",
  46400=>"000100111",
  46401=>"010100010",
  46402=>"111101000",
  46403=>"000001111",
  46404=>"011100111",
  46405=>"100111001",
  46406=>"010010101",
  46407=>"001001001",
  46408=>"010010010",
  46409=>"001000110",
  46410=>"001101110",
  46411=>"010100011",
  46412=>"001011000",
  46413=>"111110010",
  46414=>"000101100",
  46415=>"111111101",
  46416=>"001100110",
  46417=>"101010001",
  46418=>"001001000",
  46419=>"010101001",
  46420=>"000100011",
  46421=>"100000011",
  46422=>"011011100",
  46423=>"110011010",
  46424=>"001100011",
  46425=>"100000010",
  46426=>"101001000",
  46427=>"111110110",
  46428=>"010110011",
  46429=>"000111001",
  46430=>"001100111",
  46431=>"111100110",
  46432=>"001111101",
  46433=>"111000110",
  46434=>"110010010",
  46435=>"110111110",
  46436=>"101101101",
  46437=>"101100011",
  46438=>"001001100",
  46439=>"011110001",
  46440=>"110111011",
  46441=>"011100010",
  46442=>"100010000",
  46443=>"000101110",
  46444=>"000010000",
  46445=>"001000000",
  46446=>"001010010",
  46447=>"110011000",
  46448=>"001000100",
  46449=>"011100010",
  46450=>"011010110",
  46451=>"011100011",
  46452=>"000010101",
  46453=>"000111111",
  46454=>"100011110",
  46455=>"111100000",
  46456=>"101010001",
  46457=>"011110000",
  46458=>"001001010",
  46459=>"111010010",
  46460=>"101010000",
  46461=>"010100100",
  46462=>"110001110",
  46463=>"010000101",
  46464=>"100001101",
  46465=>"000111100",
  46466=>"110101101",
  46467=>"010011001",
  46468=>"011011001",
  46469=>"001111101",
  46470=>"111111111",
  46471=>"001000111",
  46472=>"100110011",
  46473=>"100111001",
  46474=>"001111011",
  46475=>"000001000",
  46476=>"000101011",
  46477=>"001100011",
  46478=>"110000000",
  46479=>"001100100",
  46480=>"011111110",
  46481=>"010110000",
  46482=>"011010110",
  46483=>"111000110",
  46484=>"111101111",
  46485=>"100011011",
  46486=>"011010110",
  46487=>"010100000",
  46488=>"110001110",
  46489=>"011001100",
  46490=>"000110101",
  46491=>"011000000",
  46492=>"111100101",
  46493=>"001001000",
  46494=>"011010101",
  46495=>"110001100",
  46496=>"000110010",
  46497=>"000110010",
  46498=>"010111110",
  46499=>"100111000",
  46500=>"000100010",
  46501=>"011001000",
  46502=>"110111001",
  46503=>"000000101",
  46504=>"101011001",
  46505=>"101111011",
  46506=>"100100001",
  46507=>"010010010",
  46508=>"110111100",
  46509=>"101000101",
  46510=>"101100110",
  46511=>"010111011",
  46512=>"101010101",
  46513=>"010110111",
  46514=>"000010110",
  46515=>"110001101",
  46516=>"101011001",
  46517=>"001100010",
  46518=>"101011111",
  46519=>"110101110",
  46520=>"001101110",
  46521=>"001001011",
  46522=>"010010100",
  46523=>"010000110",
  46524=>"110110100",
  46525=>"111001110",
  46526=>"001101001",
  46527=>"001111110",
  46528=>"011100000",
  46529=>"011011111",
  46530=>"111011101",
  46531=>"001100011",
  46532=>"000101110",
  46533=>"011101000",
  46534=>"001111001",
  46535=>"111111010",
  46536=>"111110110",
  46537=>"001100001",
  46538=>"111101001",
  46539=>"100111011",
  46540=>"100010001",
  46541=>"010111100",
  46542=>"010101010",
  46543=>"100011101",
  46544=>"000001001",
  46545=>"101111000",
  46546=>"101001101",
  46547=>"100001101",
  46548=>"000101110",
  46549=>"100011001",
  46550=>"011001011",
  46551=>"100100101",
  46552=>"010100100",
  46553=>"100010111",
  46554=>"011001101",
  46555=>"100110100",
  46556=>"010010010",
  46557=>"010000001",
  46558=>"011110011",
  46559=>"011110000",
  46560=>"001111001",
  46561=>"000000010",
  46562=>"011001001",
  46563=>"111110100",
  46564=>"010000001",
  46565=>"101100010",
  46566=>"011110100",
  46567=>"110000000",
  46568=>"111101110",
  46569=>"001001011",
  46570=>"001111111",
  46571=>"010101000",
  46572=>"100100110",
  46573=>"110001111",
  46574=>"110010000",
  46575=>"000001000",
  46576=>"111011011",
  46577=>"110101011",
  46578=>"001101111",
  46579=>"010001000",
  46580=>"110110001",
  46581=>"111010010",
  46582=>"100111111",
  46583=>"111011100",
  46584=>"111010011",
  46585=>"011111011",
  46586=>"100000010",
  46587=>"000000001",
  46588=>"010110010",
  46589=>"111110100",
  46590=>"001111001",
  46591=>"000110010",
  46592=>"101111010",
  46593=>"010011000",
  46594=>"000001011",
  46595=>"010000000",
  46596=>"001011000",
  46597=>"000000001",
  46598=>"110000110",
  46599=>"111000010",
  46600=>"000001000",
  46601=>"111101111",
  46602=>"011010101",
  46603=>"001001001",
  46604=>"000111000",
  46605=>"101101001",
  46606=>"101000000",
  46607=>"101111001",
  46608=>"100000101",
  46609=>"010011100",
  46610=>"101000011",
  46611=>"011010010",
  46612=>"110000101",
  46613=>"010011001",
  46614=>"011101001",
  46615=>"101100111",
  46616=>"111111000",
  46617=>"101101111",
  46618=>"111010010",
  46619=>"000101101",
  46620=>"000001001",
  46621=>"111000010",
  46622=>"011100101",
  46623=>"111011100",
  46624=>"010111000",
  46625=>"101111101",
  46626=>"000110110",
  46627=>"011001110",
  46628=>"110101100",
  46629=>"011011110",
  46630=>"100101001",
  46631=>"010100000",
  46632=>"001001110",
  46633=>"110110011",
  46634=>"101110011",
  46635=>"111011000",
  46636=>"101011011",
  46637=>"010111000",
  46638=>"101011001",
  46639=>"000000000",
  46640=>"101001000",
  46641=>"110000011",
  46642=>"110010100",
  46643=>"111001000",
  46644=>"100000000",
  46645=>"000001001",
  46646=>"111010110",
  46647=>"110011111",
  46648=>"100100111",
  46649=>"111010001",
  46650=>"010111110",
  46651=>"000000110",
  46652=>"111101000",
  46653=>"001011100",
  46654=>"001010101",
  46655=>"101000010",
  46656=>"111011010",
  46657=>"100111100",
  46658=>"010011111",
  46659=>"000111111",
  46660=>"000010111",
  46661=>"001111010",
  46662=>"111010001",
  46663=>"011101000",
  46664=>"001000010",
  46665=>"101010100",
  46666=>"111101101",
  46667=>"000111101",
  46668=>"001011010",
  46669=>"000010100",
  46670=>"010101101",
  46671=>"101010111",
  46672=>"000100010",
  46673=>"010100101",
  46674=>"010111100",
  46675=>"000110001",
  46676=>"011101111",
  46677=>"101111110",
  46678=>"000100100",
  46679=>"001010100",
  46680=>"111010001",
  46681=>"011101010",
  46682=>"110011110",
  46683=>"000000011",
  46684=>"100000110",
  46685=>"101101100",
  46686=>"111000111",
  46687=>"111111011",
  46688=>"011101111",
  46689=>"010000010",
  46690=>"110110001",
  46691=>"001111101",
  46692=>"000001100",
  46693=>"101100010",
  46694=>"000001100",
  46695=>"001111001",
  46696=>"011000001",
  46697=>"011110011",
  46698=>"111001101",
  46699=>"001001000",
  46700=>"011001101",
  46701=>"001101011",
  46702=>"011111110",
  46703=>"111100101",
  46704=>"001000111",
  46705=>"001011101",
  46706=>"100110010",
  46707=>"101110001",
  46708=>"111101001",
  46709=>"011100000",
  46710=>"010010000",
  46711=>"000100001",
  46712=>"001001000",
  46713=>"101000011",
  46714=>"000101000",
  46715=>"100001110",
  46716=>"100110001",
  46717=>"001011011",
  46718=>"010000110",
  46719=>"100111101",
  46720=>"001111111",
  46721=>"001001010",
  46722=>"001000111",
  46723=>"001101101",
  46724=>"010000011",
  46725=>"011000010",
  46726=>"111010111",
  46727=>"111111000",
  46728=>"001010101",
  46729=>"011000001",
  46730=>"001111110",
  46731=>"000111001",
  46732=>"111101001",
  46733=>"110011010",
  46734=>"101010000",
  46735=>"000100110",
  46736=>"101011100",
  46737=>"100001100",
  46738=>"000001001",
  46739=>"011101000",
  46740=>"111111011",
  46741=>"111110011",
  46742=>"000001100",
  46743=>"001110011",
  46744=>"111111100",
  46745=>"111111111",
  46746=>"110101011",
  46747=>"100100111",
  46748=>"100001100",
  46749=>"111010011",
  46750=>"000111011",
  46751=>"101101100",
  46752=>"100010001",
  46753=>"110011111",
  46754=>"010010111",
  46755=>"111101101",
  46756=>"111110110",
  46757=>"011011010",
  46758=>"110011001",
  46759=>"100000001",
  46760=>"111100000",
  46761=>"010000100",
  46762=>"000000001",
  46763=>"010110101",
  46764=>"110101010",
  46765=>"101010011",
  46766=>"100101001",
  46767=>"000010010",
  46768=>"111110111",
  46769=>"100001100",
  46770=>"111001100",
  46771=>"100100011",
  46772=>"000001101",
  46773=>"111111001",
  46774=>"111001001",
  46775=>"111100011",
  46776=>"111100110",
  46777=>"100000100",
  46778=>"111110001",
  46779=>"101000101",
  46780=>"000001111",
  46781=>"110110001",
  46782=>"110100000",
  46783=>"101010101",
  46784=>"011011000",
  46785=>"010001010",
  46786=>"101010001",
  46787=>"001011111",
  46788=>"001000101",
  46789=>"001100001",
  46790=>"111111101",
  46791=>"000001001",
  46792=>"111111000",
  46793=>"000011011",
  46794=>"011101000",
  46795=>"100100010",
  46796=>"000011111",
  46797=>"101100011",
  46798=>"101010001",
  46799=>"011000100",
  46800=>"001011000",
  46801=>"101101001",
  46802=>"110100000",
  46803=>"111001101",
  46804=>"101100110",
  46805=>"011010101",
  46806=>"111001001",
  46807=>"000010011",
  46808=>"000111010",
  46809=>"101000111",
  46810=>"110110110",
  46811=>"011101110",
  46812=>"110000100",
  46813=>"100111111",
  46814=>"101011111",
  46815=>"111000001",
  46816=>"100000010",
  46817=>"001010110",
  46818=>"011011011",
  46819=>"000010001",
  46820=>"110110100",
  46821=>"110011110",
  46822=>"010000100",
  46823=>"000110010",
  46824=>"000100101",
  46825=>"001110101",
  46826=>"110011111",
  46827=>"110101110",
  46828=>"100011000",
  46829=>"110000110",
  46830=>"001011101",
  46831=>"000011110",
  46832=>"000101010",
  46833=>"010010010",
  46834=>"100010000",
  46835=>"110101111",
  46836=>"000000011",
  46837=>"011110000",
  46838=>"110111100",
  46839=>"010000111",
  46840=>"110100111",
  46841=>"011110100",
  46842=>"100110101",
  46843=>"000101001",
  46844=>"010010101",
  46845=>"110011101",
  46846=>"101101100",
  46847=>"000010001",
  46848=>"110110100",
  46849=>"111111001",
  46850=>"111110111",
  46851=>"111101111",
  46852=>"011001100",
  46853=>"000010111",
  46854=>"101110111",
  46855=>"101001011",
  46856=>"100110010",
  46857=>"101101101",
  46858=>"010101010",
  46859=>"110101100",
  46860=>"000001100",
  46861=>"110010011",
  46862=>"010011100",
  46863=>"111001001",
  46864=>"111101011",
  46865=>"000001001",
  46866=>"001011111",
  46867=>"101101010",
  46868=>"001101111",
  46869=>"110000110",
  46870=>"000010000",
  46871=>"100010001",
  46872=>"111101011",
  46873=>"001010011",
  46874=>"110010111",
  46875=>"000110111",
  46876=>"000011010",
  46877=>"110010111",
  46878=>"101001101",
  46879=>"101001100",
  46880=>"010101100",
  46881=>"000101110",
  46882=>"111111101",
  46883=>"010111110",
  46884=>"111011110",
  46885=>"011011100",
  46886=>"010100000",
  46887=>"100000000",
  46888=>"110110111",
  46889=>"010001101",
  46890=>"000101000",
  46891=>"111000011",
  46892=>"101000000",
  46893=>"001001111",
  46894=>"110111011",
  46895=>"001011000",
  46896=>"011101000",
  46897=>"001111111",
  46898=>"110100000",
  46899=>"001001110",
  46900=>"101101101",
  46901=>"100000011",
  46902=>"101001110",
  46903=>"100100001",
  46904=>"000010110",
  46905=>"000110000",
  46906=>"010101000",
  46907=>"110000010",
  46908=>"001000011",
  46909=>"001111111",
  46910=>"010100000",
  46911=>"101110101",
  46912=>"100111111",
  46913=>"110000001",
  46914=>"010110100",
  46915=>"100100010",
  46916=>"100001100",
  46917=>"100001110",
  46918=>"101111110",
  46919=>"010111101",
  46920=>"001010100",
  46921=>"110100000",
  46922=>"011001001",
  46923=>"101111101",
  46924=>"111001001",
  46925=>"011101000",
  46926=>"010110100",
  46927=>"010000011",
  46928=>"110100010",
  46929=>"000000000",
  46930=>"001011000",
  46931=>"001010101",
  46932=>"111010100",
  46933=>"011010101",
  46934=>"100010100",
  46935=>"001100100",
  46936=>"110110111",
  46937=>"101110101",
  46938=>"000000100",
  46939=>"010110101",
  46940=>"001010111",
  46941=>"100100111",
  46942=>"101011100",
  46943=>"101010011",
  46944=>"111011100",
  46945=>"101000001",
  46946=>"000100000",
  46947=>"111101010",
  46948=>"000010001",
  46949=>"001001010",
  46950=>"100111111",
  46951=>"010011111",
  46952=>"011100110",
  46953=>"010110100",
  46954=>"010000000",
  46955=>"111100001",
  46956=>"101011010",
  46957=>"110110011",
  46958=>"101011110",
  46959=>"100110011",
  46960=>"011000100",
  46961=>"001010110",
  46962=>"100000011",
  46963=>"101000011",
  46964=>"111100101",
  46965=>"101000000",
  46966=>"110000111",
  46967=>"001010111",
  46968=>"010000110",
  46969=>"100011000",
  46970=>"111000001",
  46971=>"101100111",
  46972=>"100001000",
  46973=>"010000011",
  46974=>"110010001",
  46975=>"001111000",
  46976=>"011111001",
  46977=>"100010000",
  46978=>"100110000",
  46979=>"111000011",
  46980=>"001010100",
  46981=>"000000111",
  46982=>"100101100",
  46983=>"101001001",
  46984=>"101010101",
  46985=>"001101101",
  46986=>"100110101",
  46987=>"101100010",
  46988=>"110110000",
  46989=>"001111111",
  46990=>"001100111",
  46991=>"000111100",
  46992=>"000011000",
  46993=>"000110001",
  46994=>"000100010",
  46995=>"100001110",
  46996=>"111101110",
  46997=>"011010010",
  46998=>"100100111",
  46999=>"111101001",
  47000=>"001110111",
  47001=>"110110101",
  47002=>"110101100",
  47003=>"010000101",
  47004=>"001111111",
  47005=>"101001100",
  47006=>"110110011",
  47007=>"011001110",
  47008=>"001001101",
  47009=>"101111100",
  47010=>"000110000",
  47011=>"001000100",
  47012=>"100010000",
  47013=>"000101111",
  47014=>"001000011",
  47015=>"001001111",
  47016=>"011011111",
  47017=>"110111001",
  47018=>"101110111",
  47019=>"111010100",
  47020=>"001010001",
  47021=>"111100001",
  47022=>"111000100",
  47023=>"101011101",
  47024=>"100111100",
  47025=>"010101100",
  47026=>"001001000",
  47027=>"100111111",
  47028=>"110111010",
  47029=>"001110110",
  47030=>"011111001",
  47031=>"111010010",
  47032=>"011100111",
  47033=>"111011100",
  47034=>"111001110",
  47035=>"101101101",
  47036=>"111101111",
  47037=>"100001000",
  47038=>"001101000",
  47039=>"010111000",
  47040=>"011111110",
  47041=>"111110100",
  47042=>"010110111",
  47043=>"100001110",
  47044=>"010101111",
  47045=>"101011100",
  47046=>"100011011",
  47047=>"011100111",
  47048=>"101000001",
  47049=>"001010101",
  47050=>"011110101",
  47051=>"110110001",
  47052=>"000010001",
  47053=>"010011100",
  47054=>"100000010",
  47055=>"001111111",
  47056=>"011000001",
  47057=>"001111111",
  47058=>"100101110",
  47059=>"011011000",
  47060=>"110000101",
  47061=>"001001011",
  47062=>"101000010",
  47063=>"011011010",
  47064=>"010001100",
  47065=>"000101001",
  47066=>"111011110",
  47067=>"111101001",
  47068=>"110101010",
  47069=>"011100011",
  47070=>"111100100",
  47071=>"111001000",
  47072=>"010010000",
  47073=>"000000101",
  47074=>"000111000",
  47075=>"001000111",
  47076=>"110001100",
  47077=>"101100101",
  47078=>"111101100",
  47079=>"101111101",
  47080=>"000001110",
  47081=>"010000010",
  47082=>"001001011",
  47083=>"010000100",
  47084=>"001000000",
  47085=>"111110000",
  47086=>"010011011",
  47087=>"001011000",
  47088=>"010011101",
  47089=>"000001011",
  47090=>"111001111",
  47091=>"101101010",
  47092=>"110111110",
  47093=>"000000110",
  47094=>"001100110",
  47095=>"011110111",
  47096=>"101110010",
  47097=>"101011000",
  47098=>"001111100",
  47099=>"010101100",
  47100=>"110000000",
  47101=>"111101110",
  47102=>"000110001",
  47103=>"101011001",
  47104=>"110100011",
  47105=>"000000101",
  47106=>"011111111",
  47107=>"001011111",
  47108=>"101001010",
  47109=>"001011010",
  47110=>"101110111",
  47111=>"000000001",
  47112=>"000100101",
  47113=>"100101111",
  47114=>"101111010",
  47115=>"111111111",
  47116=>"000110100",
  47117=>"001100011",
  47118=>"011010111",
  47119=>"110110111",
  47120=>"000111111",
  47121=>"111011000",
  47122=>"110001011",
  47123=>"101100001",
  47124=>"111110101",
  47125=>"000110110",
  47126=>"100111011",
  47127=>"100101100",
  47128=>"101111010",
  47129=>"000100110",
  47130=>"001010001",
  47131=>"001100010",
  47132=>"111000011",
  47133=>"111011001",
  47134=>"110010000",
  47135=>"110110010",
  47136=>"000001000",
  47137=>"111010101",
  47138=>"010110101",
  47139=>"001111011",
  47140=>"100111000",
  47141=>"010011001",
  47142=>"101001110",
  47143=>"100110100",
  47144=>"000011001",
  47145=>"111000111",
  47146=>"111100111",
  47147=>"011010101",
  47148=>"010000000",
  47149=>"110101101",
  47150=>"001100100",
  47151=>"010100000",
  47152=>"011111110",
  47153=>"001001001",
  47154=>"100101011",
  47155=>"000101010",
  47156=>"110001100",
  47157=>"000111011",
  47158=>"011101010",
  47159=>"000101101",
  47160=>"000110110",
  47161=>"110010010",
  47162=>"110010110",
  47163=>"101110111",
  47164=>"010101000",
  47165=>"000100100",
  47166=>"110010001",
  47167=>"111000101",
  47168=>"110001110",
  47169=>"111101000",
  47170=>"101111100",
  47171=>"111110111",
  47172=>"110111110",
  47173=>"011100100",
  47174=>"110110001",
  47175=>"101011001",
  47176=>"010001100",
  47177=>"011000000",
  47178=>"101101000",
  47179=>"111110010",
  47180=>"011110011",
  47181=>"101111101",
  47182=>"010000100",
  47183=>"001101010",
  47184=>"100010111",
  47185=>"111111110",
  47186=>"110110001",
  47187=>"011000011",
  47188=>"000001011",
  47189=>"011000111",
  47190=>"101111101",
  47191=>"100001100",
  47192=>"100100000",
  47193=>"111001100",
  47194=>"110001111",
  47195=>"110111101",
  47196=>"111111101",
  47197=>"111011110",
  47198=>"111011110",
  47199=>"110011111",
  47200=>"000000101",
  47201=>"111100110",
  47202=>"011001000",
  47203=>"100110010",
  47204=>"110101111",
  47205=>"110101010",
  47206=>"000011101",
  47207=>"110111110",
  47208=>"111000000",
  47209=>"100100111",
  47210=>"011111111",
  47211=>"111101100",
  47212=>"001101101",
  47213=>"010100110",
  47214=>"111111101",
  47215=>"111101010",
  47216=>"011100010",
  47217=>"110101101",
  47218=>"111101111",
  47219=>"101101001",
  47220=>"111000101",
  47221=>"101111101",
  47222=>"011010111",
  47223=>"101100001",
  47224=>"110000000",
  47225=>"100111110",
  47226=>"111101011",
  47227=>"100110101",
  47228=>"001000101",
  47229=>"010011000",
  47230=>"101100101",
  47231=>"110101010",
  47232=>"010000110",
  47233=>"000001001",
  47234=>"011001000",
  47235=>"100010100",
  47236=>"011000011",
  47237=>"110111100",
  47238=>"110100101",
  47239=>"000011010",
  47240=>"000001001",
  47241=>"111110100",
  47242=>"000000011",
  47243=>"011011011",
  47244=>"000011010",
  47245=>"111110100",
  47246=>"000011111",
  47247=>"000001100",
  47248=>"000101101",
  47249=>"111010001",
  47250=>"011100100",
  47251=>"011101101",
  47252=>"100100111",
  47253=>"101001000",
  47254=>"010111000",
  47255=>"010010000",
  47256=>"000001011",
  47257=>"101000000",
  47258=>"010011011",
  47259=>"000101011",
  47260=>"111111100",
  47261=>"111111000",
  47262=>"000011111",
  47263=>"001100011",
  47264=>"100100010",
  47265=>"110101000",
  47266=>"010010111",
  47267=>"100111011",
  47268=>"010010010",
  47269=>"100001001",
  47270=>"010111101",
  47271=>"000010010",
  47272=>"000100001",
  47273=>"001101010",
  47274=>"010101000",
  47275=>"000100000",
  47276=>"011011101",
  47277=>"101000001",
  47278=>"100000011",
  47279=>"110001001",
  47280=>"100101001",
  47281=>"110000011",
  47282=>"101001100",
  47283=>"000001001",
  47284=>"010011101",
  47285=>"000101011",
  47286=>"001000000",
  47287=>"001111100",
  47288=>"110010100",
  47289=>"100100111",
  47290=>"101000100",
  47291=>"000101000",
  47292=>"011000010",
  47293=>"110010011",
  47294=>"001010110",
  47295=>"010000111",
  47296=>"111100111",
  47297=>"000110100",
  47298=>"111010101",
  47299=>"010000100",
  47300=>"101110000",
  47301=>"111110110",
  47302=>"110000111",
  47303=>"101000011",
  47304=>"110001100",
  47305=>"000100110",
  47306=>"101001000",
  47307=>"101011111",
  47308=>"000000111",
  47309=>"100001101",
  47310=>"110000100",
  47311=>"010000110",
  47312=>"000001101",
  47313=>"000001000",
  47314=>"110111110",
  47315=>"001110100",
  47316=>"011111001",
  47317=>"111001101",
  47318=>"011011001",
  47319=>"111110010",
  47320=>"011100111",
  47321=>"101010111",
  47322=>"101110101",
  47323=>"100011101",
  47324=>"101010001",
  47325=>"001000111",
  47326=>"101100001",
  47327=>"111001111",
  47328=>"010100100",
  47329=>"000100110",
  47330=>"001110011",
  47331=>"101100101",
  47332=>"000001011",
  47333=>"101101111",
  47334=>"110110111",
  47335=>"011010000",
  47336=>"010000101",
  47337=>"001001001",
  47338=>"110011011",
  47339=>"101100101",
  47340=>"001111111",
  47341=>"101100011",
  47342=>"001101100",
  47343=>"001101111",
  47344=>"011101010",
  47345=>"101101000",
  47346=>"110111001",
  47347=>"001000110",
  47348=>"000001000",
  47349=>"010001110",
  47350=>"111011010",
  47351=>"001010101",
  47352=>"101100100",
  47353=>"110111101",
  47354=>"100101101",
  47355=>"000111000",
  47356=>"100100001",
  47357=>"110000101",
  47358=>"111000011",
  47359=>"100000101",
  47360=>"111101100",
  47361=>"001111101",
  47362=>"100100010",
  47363=>"101011111",
  47364=>"101111001",
  47365=>"100001101",
  47366=>"101101101",
  47367=>"100101001",
  47368=>"111001010",
  47369=>"110101010",
  47370=>"101000100",
  47371=>"111110011",
  47372=>"000011010",
  47373=>"111111101",
  47374=>"001110010",
  47375=>"000100000",
  47376=>"101010011",
  47377=>"011110101",
  47378=>"101011100",
  47379=>"110101011",
  47380=>"111111111",
  47381=>"111110000",
  47382=>"010110111",
  47383=>"110011011",
  47384=>"000000110",
  47385=>"001010001",
  47386=>"110110010",
  47387=>"001110010",
  47388=>"110001111",
  47389=>"111100110",
  47390=>"000000101",
  47391=>"011000100",
  47392=>"110011011",
  47393=>"101101110",
  47394=>"011011100",
  47395=>"010010111",
  47396=>"000011011",
  47397=>"000001100",
  47398=>"010010110",
  47399=>"101001110",
  47400=>"011010100",
  47401=>"010100000",
  47402=>"101101110",
  47403=>"110010011",
  47404=>"000011101",
  47405=>"110110010",
  47406=>"000011101",
  47407=>"101101101",
  47408=>"110110111",
  47409=>"100011001",
  47410=>"001000110",
  47411=>"111001100",
  47412=>"111000111",
  47413=>"110100000",
  47414=>"010011110",
  47415=>"000110000",
  47416=>"011111011",
  47417=>"011011000",
  47418=>"100110111",
  47419=>"100000100",
  47420=>"001110100",
  47421=>"010000010",
  47422=>"100000111",
  47423=>"010010000",
  47424=>"110010100",
  47425=>"111011110",
  47426=>"100000100",
  47427=>"011010010",
  47428=>"101100101",
  47429=>"011010000",
  47430=>"101100010",
  47431=>"101000010",
  47432=>"110110100",
  47433=>"101100000",
  47434=>"101100010",
  47435=>"110010000",
  47436=>"001001011",
  47437=>"001000001",
  47438=>"100001000",
  47439=>"111010001",
  47440=>"011101010",
  47441=>"101100000",
  47442=>"110010011",
  47443=>"111010111",
  47444=>"100111101",
  47445=>"010011111",
  47446=>"000101111",
  47447=>"001101101",
  47448=>"110110101",
  47449=>"111010011",
  47450=>"001000110",
  47451=>"110110000",
  47452=>"111111100",
  47453=>"111010100",
  47454=>"010011010",
  47455=>"110100000",
  47456=>"111001010",
  47457=>"001011010",
  47458=>"100111111",
  47459=>"111110110",
  47460=>"101111101",
  47461=>"011111111",
  47462=>"111010100",
  47463=>"110010000",
  47464=>"000001001",
  47465=>"000001111",
  47466=>"000001011",
  47467=>"111101100",
  47468=>"101010010",
  47469=>"100010000",
  47470=>"110110101",
  47471=>"000111100",
  47472=>"000000011",
  47473=>"111111001",
  47474=>"000010010",
  47475=>"101111110",
  47476=>"111001000",
  47477=>"100011011",
  47478=>"100011110",
  47479=>"111011010",
  47480=>"010001110",
  47481=>"000101000",
  47482=>"100010000",
  47483=>"100000001",
  47484=>"011101111",
  47485=>"000100100",
  47486=>"110000101",
  47487=>"101101011",
  47488=>"110001111",
  47489=>"110111100",
  47490=>"100010101",
  47491=>"111100111",
  47492=>"000111100",
  47493=>"111001011",
  47494=>"110001101",
  47495=>"000111110",
  47496=>"001010101",
  47497=>"101010101",
  47498=>"000111100",
  47499=>"000001110",
  47500=>"010001111",
  47501=>"000000010",
  47502=>"000110001",
  47503=>"101010011",
  47504=>"111101110",
  47505=>"100101111",
  47506=>"011011101",
  47507=>"001100010",
  47508=>"010100110",
  47509=>"110111011",
  47510=>"100111111",
  47511=>"111000001",
  47512=>"111111101",
  47513=>"100000110",
  47514=>"001001111",
  47515=>"111101110",
  47516=>"000010110",
  47517=>"011100101",
  47518=>"000011110",
  47519=>"111100100",
  47520=>"110101101",
  47521=>"111110111",
  47522=>"001010000",
  47523=>"101110111",
  47524=>"001011000",
  47525=>"010111101",
  47526=>"011101001",
  47527=>"010101000",
  47528=>"000100001",
  47529=>"010101000",
  47530=>"100101110",
  47531=>"000111111",
  47532=>"111101111",
  47533=>"001001100",
  47534=>"111110111",
  47535=>"001110011",
  47536=>"101101001",
  47537=>"010100110",
  47538=>"000101101",
  47539=>"101101011",
  47540=>"100100010",
  47541=>"000001100",
  47542=>"111011111",
  47543=>"010010111",
  47544=>"111011010",
  47545=>"011101001",
  47546=>"101101011",
  47547=>"110000010",
  47548=>"100001111",
  47549=>"100010011",
  47550=>"111110001",
  47551=>"001100001",
  47552=>"001011010",
  47553=>"110011011",
  47554=>"011001011",
  47555=>"000100000",
  47556=>"100000010",
  47557=>"011100011",
  47558=>"011110101",
  47559=>"001000100",
  47560=>"101010010",
  47561=>"011110010",
  47562=>"011010101",
  47563=>"010001000",
  47564=>"110111011",
  47565=>"110101011",
  47566=>"101011001",
  47567=>"100110100",
  47568=>"011000101",
  47569=>"000110110",
  47570=>"110110001",
  47571=>"001000011",
  47572=>"111011111",
  47573=>"110000011",
  47574=>"000000001",
  47575=>"101100110",
  47576=>"011011001",
  47577=>"101011100",
  47578=>"100100011",
  47579=>"100000010",
  47580=>"000000111",
  47581=>"101100110",
  47582=>"010101000",
  47583=>"010011101",
  47584=>"011101001",
  47585=>"111100001",
  47586=>"000110110",
  47587=>"010110000",
  47588=>"011001100",
  47589=>"000001111",
  47590=>"110100001",
  47591=>"110011011",
  47592=>"011000100",
  47593=>"100001100",
  47594=>"111000100",
  47595=>"010010010",
  47596=>"011101001",
  47597=>"110001101",
  47598=>"000101100",
  47599=>"011000110",
  47600=>"001011000",
  47601=>"000011001",
  47602=>"010101010",
  47603=>"001111011",
  47604=>"100100100",
  47605=>"010011000",
  47606=>"110110100",
  47607=>"011000100",
  47608=>"011111110",
  47609=>"111000011",
  47610=>"100101110",
  47611=>"100001010",
  47612=>"111111101",
  47613=>"101000100",
  47614=>"011110111",
  47615=>"111011000",
  47616=>"011001010",
  47617=>"000110101",
  47618=>"011000001",
  47619=>"110001110",
  47620=>"101111000",
  47621=>"000000111",
  47622=>"110100110",
  47623=>"101101001",
  47624=>"011100110",
  47625=>"011000110",
  47626=>"011001011",
  47627=>"001000000",
  47628=>"010001111",
  47629=>"011100010",
  47630=>"000100111",
  47631=>"110001011",
  47632=>"010011101",
  47633=>"110010010",
  47634=>"101001010",
  47635=>"001100000",
  47636=>"000101001",
  47637=>"101100100",
  47638=>"010001000",
  47639=>"000001101",
  47640=>"111110000",
  47641=>"000111101",
  47642=>"101110001",
  47643=>"110111000",
  47644=>"001001100",
  47645=>"100010110",
  47646=>"100100111",
  47647=>"100111000",
  47648=>"110010000",
  47649=>"111000011",
  47650=>"111101000",
  47651=>"111011110",
  47652=>"000001110",
  47653=>"100101101",
  47654=>"001010100",
  47655=>"000101000",
  47656=>"100001010",
  47657=>"010100000",
  47658=>"100011001",
  47659=>"101100100",
  47660=>"110111111",
  47661=>"000100001",
  47662=>"111000000",
  47663=>"010101100",
  47664=>"000001010",
  47665=>"000011110",
  47666=>"110000011",
  47667=>"111111110",
  47668=>"110110101",
  47669=>"010110111",
  47670=>"010111101",
  47671=>"111101111",
  47672=>"001101010",
  47673=>"110011110",
  47674=>"011101001",
  47675=>"001101101",
  47676=>"101100000",
  47677=>"010111010",
  47678=>"100000111",
  47679=>"001000100",
  47680=>"001010110",
  47681=>"111101000",
  47682=>"110010110",
  47683=>"010010110",
  47684=>"100100100",
  47685=>"101110101",
  47686=>"010001111",
  47687=>"100111111",
  47688=>"000110010",
  47689=>"000000110",
  47690=>"000000000",
  47691=>"111101111",
  47692=>"110111010",
  47693=>"101000100",
  47694=>"111010010",
  47695=>"110110000",
  47696=>"010100110",
  47697=>"011011111",
  47698=>"000110100",
  47699=>"001011010",
  47700=>"110100011",
  47701=>"111110110",
  47702=>"001011111",
  47703=>"100011010",
  47704=>"001111010",
  47705=>"111110001",
  47706=>"001101010",
  47707=>"110100110",
  47708=>"000010000",
  47709=>"110100000",
  47710=>"111101111",
  47711=>"011100101",
  47712=>"010001110",
  47713=>"000001011",
  47714=>"111100111",
  47715=>"111110111",
  47716=>"001001001",
  47717=>"001100001",
  47718=>"110000011",
  47719=>"100100011",
  47720=>"111001001",
  47721=>"110001000",
  47722=>"001001110",
  47723=>"010000011",
  47724=>"111110010",
  47725=>"100011111",
  47726=>"111011010",
  47727=>"001101100",
  47728=>"000011110",
  47729=>"011010011",
  47730=>"101100100",
  47731=>"110010000",
  47732=>"110100001",
  47733=>"000001010",
  47734=>"110110100",
  47735=>"010100100",
  47736=>"011100110",
  47737=>"000010101",
  47738=>"101110000",
  47739=>"001001001",
  47740=>"110101001",
  47741=>"100001100",
  47742=>"101001110",
  47743=>"101010111",
  47744=>"000110100",
  47745=>"111100010",
  47746=>"000011101",
  47747=>"010111000",
  47748=>"111010011",
  47749=>"000100011",
  47750=>"111101011",
  47751=>"100010101",
  47752=>"111011111",
  47753=>"011111111",
  47754=>"111101010",
  47755=>"001010001",
  47756=>"111100100",
  47757=>"010000101",
  47758=>"100010100",
  47759=>"110110001",
  47760=>"111101001",
  47761=>"001100101",
  47762=>"001001110",
  47763=>"001011101",
  47764=>"110010000",
  47765=>"111001001",
  47766=>"011011110",
  47767=>"010000001",
  47768=>"111101011",
  47769=>"100111110",
  47770=>"100011011",
  47771=>"110100000",
  47772=>"000000011",
  47773=>"100101100",
  47774=>"010100011",
  47775=>"011110110",
  47776=>"000000101",
  47777=>"011110011",
  47778=>"101000001",
  47779=>"011000100",
  47780=>"100111000",
  47781=>"101111101",
  47782=>"111111000",
  47783=>"110011000",
  47784=>"011101001",
  47785=>"001110101",
  47786=>"010000111",
  47787=>"000001100",
  47788=>"001101111",
  47789=>"101100110",
  47790=>"001110110",
  47791=>"000100000",
  47792=>"100110001",
  47793=>"111100111",
  47794=>"101011111",
  47795=>"010010100",
  47796=>"101001001",
  47797=>"010111000",
  47798=>"011011011",
  47799=>"001010001",
  47800=>"101101001",
  47801=>"100110110",
  47802=>"101101010",
  47803=>"101101111",
  47804=>"001110111",
  47805=>"000001010",
  47806=>"110100000",
  47807=>"110110001",
  47808=>"000011100",
  47809=>"111111111",
  47810=>"001010100",
  47811=>"110101001",
  47812=>"001010000",
  47813=>"111110101",
  47814=>"110110010",
  47815=>"101101111",
  47816=>"010001010",
  47817=>"001011111",
  47818=>"100011000",
  47819=>"100000001",
  47820=>"011101110",
  47821=>"001000110",
  47822=>"010010010",
  47823=>"101000111",
  47824=>"001111000",
  47825=>"001100011",
  47826=>"011011000",
  47827=>"011000001",
  47828=>"110000111",
  47829=>"111111111",
  47830=>"110111100",
  47831=>"100101100",
  47832=>"011111010",
  47833=>"011000000",
  47834=>"110010101",
  47835=>"010110110",
  47836=>"000101110",
  47837=>"000111000",
  47838=>"011101001",
  47839=>"111011111",
  47840=>"011011111",
  47841=>"001001110",
  47842=>"101011101",
  47843=>"010011001",
  47844=>"110000000",
  47845=>"100000110",
  47846=>"111000010",
  47847=>"000100111",
  47848=>"101100101",
  47849=>"100011110",
  47850=>"001000011",
  47851=>"110011000",
  47852=>"001000010",
  47853=>"010100100",
  47854=>"010010011",
  47855=>"100111110",
  47856=>"100010000",
  47857=>"111001100",
  47858=>"111111110",
  47859=>"111110111",
  47860=>"010101000",
  47861=>"111010001",
  47862=>"010010001",
  47863=>"010010110",
  47864=>"111110100",
  47865=>"011010101",
  47866=>"001010000",
  47867=>"011100000",
  47868=>"111000111",
  47869=>"100100010",
  47870=>"111110001",
  47871=>"101000111",
  47872=>"101101101",
  47873=>"001011111",
  47874=>"110001000",
  47875=>"011011000",
  47876=>"010001100",
  47877=>"101000111",
  47878=>"111111010",
  47879=>"001010000",
  47880=>"101011101",
  47881=>"110001001",
  47882=>"111000101",
  47883=>"001001011",
  47884=>"010111011",
  47885=>"100011000",
  47886=>"110000010",
  47887=>"010111110",
  47888=>"111011001",
  47889=>"110101000",
  47890=>"101011000",
  47891=>"100101000",
  47892=>"011001011",
  47893=>"000010110",
  47894=>"010111111",
  47895=>"101110011",
  47896=>"010010000",
  47897=>"011001000",
  47898=>"011101010",
  47899=>"111100010",
  47900=>"001001001",
  47901=>"111011110",
  47902=>"100111110",
  47903=>"001010110",
  47904=>"100010111",
  47905=>"111111100",
  47906=>"100101110",
  47907=>"111000100",
  47908=>"100110111",
  47909=>"000000101",
  47910=>"001101100",
  47911=>"001101110",
  47912=>"100001010",
  47913=>"000111001",
  47914=>"000010100",
  47915=>"111001010",
  47916=>"001010111",
  47917=>"100111010",
  47918=>"111100001",
  47919=>"100100100",
  47920=>"100010101",
  47921=>"011111111",
  47922=>"001100000",
  47923=>"100010111",
  47924=>"101101010",
  47925=>"111010011",
  47926=>"110110010",
  47927=>"011101111",
  47928=>"001100110",
  47929=>"100101100",
  47930=>"000011000",
  47931=>"001100101",
  47932=>"111011111",
  47933=>"101010111",
  47934=>"001010011",
  47935=>"101100000",
  47936=>"011000010",
  47937=>"011101000",
  47938=>"101100110",
  47939=>"100000111",
  47940=>"011000000",
  47941=>"111010010",
  47942=>"010110011",
  47943=>"110000000",
  47944=>"010010010",
  47945=>"110100010",
  47946=>"010001000",
  47947=>"001010000",
  47948=>"111101011",
  47949=>"100110111",
  47950=>"100111111",
  47951=>"100110110",
  47952=>"110001101",
  47953=>"001111111",
  47954=>"000111111",
  47955=>"100111110",
  47956=>"000100000",
  47957=>"001001101",
  47958=>"111000111",
  47959=>"011010111",
  47960=>"110110111",
  47961=>"000110011",
  47962=>"011010101",
  47963=>"101100101",
  47964=>"000110000",
  47965=>"010101001",
  47966=>"000100111",
  47967=>"011100011",
  47968=>"110110110",
  47969=>"100011011",
  47970=>"111011111",
  47971=>"001111001",
  47972=>"000000111",
  47973=>"111001011",
  47974=>"100100000",
  47975=>"111010010",
  47976=>"111001110",
  47977=>"111000010",
  47978=>"001000001",
  47979=>"010010111",
  47980=>"000001000",
  47981=>"001101111",
  47982=>"010111100",
  47983=>"011011001",
  47984=>"110111110",
  47985=>"110010010",
  47986=>"001110010",
  47987=>"001100010",
  47988=>"000101001",
  47989=>"010011110",
  47990=>"011100001",
  47991=>"110000010",
  47992=>"001001011",
  47993=>"010010011",
  47994=>"000110000",
  47995=>"100110111",
  47996=>"100101111",
  47997=>"011111011",
  47998=>"010001100",
  47999=>"000110100",
  48000=>"101100010",
  48001=>"111011100",
  48002=>"111001010",
  48003=>"110111101",
  48004=>"100110100",
  48005=>"001001100",
  48006=>"010000101",
  48007=>"101010110",
  48008=>"110000000",
  48009=>"001111000",
  48010=>"100111100",
  48011=>"111110010",
  48012=>"111000001",
  48013=>"000110010",
  48014=>"100000001",
  48015=>"101111101",
  48016=>"101100100",
  48017=>"010011110",
  48018=>"000101111",
  48019=>"100011000",
  48020=>"000100011",
  48021=>"011000000",
  48022=>"000111101",
  48023=>"101011000",
  48024=>"111110001",
  48025=>"010110110",
  48026=>"101010100",
  48027=>"101100010",
  48028=>"100000000",
  48029=>"001111001",
  48030=>"110111111",
  48031=>"000110011",
  48032=>"000000010",
  48033=>"010000000",
  48034=>"010100110",
  48035=>"011010101",
  48036=>"100110000",
  48037=>"000001011",
  48038=>"110110000",
  48039=>"100100000",
  48040=>"000110111",
  48041=>"101011001",
  48042=>"111000101",
  48043=>"101000111",
  48044=>"111101001",
  48045=>"101010101",
  48046=>"001111010",
  48047=>"100001001",
  48048=>"001000110",
  48049=>"111011001",
  48050=>"001010100",
  48051=>"000000001",
  48052=>"111000110",
  48053=>"001010100",
  48054=>"100011100",
  48055=>"000001110",
  48056=>"010000110",
  48057=>"101011110",
  48058=>"010101011",
  48059=>"111011000",
  48060=>"101001000",
  48061=>"000000011",
  48062=>"110110000",
  48063=>"100001101",
  48064=>"000001000",
  48065=>"111011001",
  48066=>"001000100",
  48067=>"100100100",
  48068=>"111100110",
  48069=>"110101000",
  48070=>"111011000",
  48071=>"000110110",
  48072=>"011100100",
  48073=>"111011000",
  48074=>"111001101",
  48075=>"110110101",
  48076=>"011001011",
  48077=>"111110011",
  48078=>"001101010",
  48079=>"011000000",
  48080=>"101000111",
  48081=>"000101011",
  48082=>"001010000",
  48083=>"101110100",
  48084=>"110100110",
  48085=>"000000100",
  48086=>"010100000",
  48087=>"111100101",
  48088=>"111101111",
  48089=>"101011000",
  48090=>"101011101",
  48091=>"000101001",
  48092=>"010101100",
  48093=>"001001100",
  48094=>"001100110",
  48095=>"001000101",
  48096=>"111100011",
  48097=>"101010010",
  48098=>"000111001",
  48099=>"000000110",
  48100=>"110111000",
  48101=>"000110101",
  48102=>"111100101",
  48103=>"100010011",
  48104=>"101000111",
  48105=>"000111101",
  48106=>"000100010",
  48107=>"010110110",
  48108=>"111110101",
  48109=>"001000100",
  48110=>"101111101",
  48111=>"110010001",
  48112=>"101111110",
  48113=>"100010001",
  48114=>"101001101",
  48115=>"100110101",
  48116=>"000101100",
  48117=>"001101101",
  48118=>"100000011",
  48119=>"000000101",
  48120=>"011111001",
  48121=>"001011011",
  48122=>"111101110",
  48123=>"010001010",
  48124=>"100010111",
  48125=>"101101011",
  48126=>"111010010",
  48127=>"000101101",
  48128=>"010110111",
  48129=>"010001111",
  48130=>"110000010",
  48131=>"011011111",
  48132=>"000101100",
  48133=>"101001101",
  48134=>"001101100",
  48135=>"100100011",
  48136=>"110100011",
  48137=>"010011011",
  48138=>"100000000",
  48139=>"101101011",
  48140=>"111100100",
  48141=>"101000001",
  48142=>"010011001",
  48143=>"111100010",
  48144=>"011000100",
  48145=>"011110010",
  48146=>"101100100",
  48147=>"111011011",
  48148=>"001000101",
  48149=>"011011100",
  48150=>"110011000",
  48151=>"110011000",
  48152=>"001110000",
  48153=>"010010110",
  48154=>"001110010",
  48155=>"110001110",
  48156=>"000000110",
  48157=>"000000000",
  48158=>"000010110",
  48159=>"111010100",
  48160=>"110110001",
  48161=>"100111100",
  48162=>"100111101",
  48163=>"101011000",
  48164=>"111000111",
  48165=>"101110010",
  48166=>"100111001",
  48167=>"100011011",
  48168=>"100000010",
  48169=>"101111111",
  48170=>"111010001",
  48171=>"001110001",
  48172=>"110101010",
  48173=>"011101100",
  48174=>"110111111",
  48175=>"111000010",
  48176=>"101000110",
  48177=>"101100010",
  48178=>"101011111",
  48179=>"110111001",
  48180=>"000001011",
  48181=>"010100000",
  48182=>"100010000",
  48183=>"110001111",
  48184=>"100010101",
  48185=>"110011000",
  48186=>"001011101",
  48187=>"010101100",
  48188=>"110110010",
  48189=>"010101011",
  48190=>"000011100",
  48191=>"101010001",
  48192=>"111000001",
  48193=>"010101000",
  48194=>"101011011",
  48195=>"100010001",
  48196=>"101001101",
  48197=>"100000001",
  48198=>"111111001",
  48199=>"000110101",
  48200=>"000011010",
  48201=>"110010011",
  48202=>"011000001",
  48203=>"110110011",
  48204=>"101111001",
  48205=>"110000001",
  48206=>"111000000",
  48207=>"100100000",
  48208=>"011101010",
  48209=>"010101110",
  48210=>"100011001",
  48211=>"110111111",
  48212=>"100100000",
  48213=>"110111011",
  48214=>"101110110",
  48215=>"010100100",
  48216=>"101101100",
  48217=>"111110011",
  48218=>"001110010",
  48219=>"011010001",
  48220=>"111101000",
  48221=>"111000010",
  48222=>"111001000",
  48223=>"100000010",
  48224=>"001111010",
  48225=>"111110011",
  48226=>"110011110",
  48227=>"111010000",
  48228=>"000000010",
  48229=>"001000001",
  48230=>"011010101",
  48231=>"000101011",
  48232=>"010001001",
  48233=>"111111011",
  48234=>"111100100",
  48235=>"011010101",
  48236=>"010001001",
  48237=>"011100110",
  48238=>"101100010",
  48239=>"000010111",
  48240=>"011010111",
  48241=>"100001010",
  48242=>"101110111",
  48243=>"000010000",
  48244=>"100001001",
  48245=>"101101110",
  48246=>"100111101",
  48247=>"000111111",
  48248=>"101010011",
  48249=>"000101001",
  48250=>"000010100",
  48251=>"000110100",
  48252=>"111100010",
  48253=>"001101010",
  48254=>"110110110",
  48255=>"001000010",
  48256=>"110110111",
  48257=>"011000001",
  48258=>"101110010",
  48259=>"000111101",
  48260=>"111001000",
  48261=>"001010101",
  48262=>"101111000",
  48263=>"110110101",
  48264=>"101001011",
  48265=>"001000100",
  48266=>"000100001",
  48267=>"111000110",
  48268=>"110000000",
  48269=>"111111011",
  48270=>"000100100",
  48271=>"001101101",
  48272=>"110010100",
  48273=>"000100001",
  48274=>"101100111",
  48275=>"011011000",
  48276=>"000111100",
  48277=>"110001010",
  48278=>"100111110",
  48279=>"010110010",
  48280=>"101010101",
  48281=>"000010000",
  48282=>"011000010",
  48283=>"010010110",
  48284=>"001101010",
  48285=>"101101011",
  48286=>"010000101",
  48287=>"000111000",
  48288=>"011011010",
  48289=>"100110010",
  48290=>"111111100",
  48291=>"011011010",
  48292=>"011110101",
  48293=>"111000111",
  48294=>"000010101",
  48295=>"011110001",
  48296=>"100101110",
  48297=>"101011111",
  48298=>"011010000",
  48299=>"110000100",
  48300=>"011101001",
  48301=>"011010110",
  48302=>"101100100",
  48303=>"000110101",
  48304=>"111101001",
  48305=>"000100000",
  48306=>"111101000",
  48307=>"011011101",
  48308=>"111000101",
  48309=>"100000111",
  48310=>"010100001",
  48311=>"000111110",
  48312=>"111010010",
  48313=>"100100101",
  48314=>"001101100",
  48315=>"100000111",
  48316=>"110001010",
  48317=>"111000110",
  48318=>"111101101",
  48319=>"100100110",
  48320=>"110010010",
  48321=>"010010000",
  48322=>"111111000",
  48323=>"010100111",
  48324=>"111110010",
  48325=>"110110001",
  48326=>"000000011",
  48327=>"110100100",
  48328=>"101000011",
  48329=>"101101010",
  48330=>"000000101",
  48331=>"110010111",
  48332=>"001111000",
  48333=>"011100110",
  48334=>"110010011",
  48335=>"110110000",
  48336=>"000110011",
  48337=>"001110001",
  48338=>"010101000",
  48339=>"000011101",
  48340=>"100111011",
  48341=>"101011110",
  48342=>"110111000",
  48343=>"001101011",
  48344=>"000111100",
  48345=>"110111111",
  48346=>"011110010",
  48347=>"000100000",
  48348=>"100110101",
  48349=>"010100100",
  48350=>"000100101",
  48351=>"000010101",
  48352=>"011011000",
  48353=>"110000011",
  48354=>"110011110",
  48355=>"110011010",
  48356=>"001001001",
  48357=>"101010001",
  48358=>"101100010",
  48359=>"111010010",
  48360=>"111111111",
  48361=>"000101101",
  48362=>"000011000",
  48363=>"000100101",
  48364=>"110110110",
  48365=>"011001001",
  48366=>"011110111",
  48367=>"111000100",
  48368=>"000110110",
  48369=>"100000010",
  48370=>"111100101",
  48371=>"010101000",
  48372=>"010010100",
  48373=>"100011110",
  48374=>"000110111",
  48375=>"111111110",
  48376=>"110011010",
  48377=>"010111111",
  48378=>"001111010",
  48379=>"000010011",
  48380=>"001100111",
  48381=>"010100010",
  48382=>"001100011",
  48383=>"011001110",
  48384=>"010011011",
  48385=>"010001011",
  48386=>"110010000",
  48387=>"011010010",
  48388=>"111100010",
  48389=>"100111001",
  48390=>"001000000",
  48391=>"110110010",
  48392=>"011111011",
  48393=>"111110100",
  48394=>"010101110",
  48395=>"000101001",
  48396=>"110000000",
  48397=>"000010000",
  48398=>"000100111",
  48399=>"100000111",
  48400=>"100100010",
  48401=>"111101010",
  48402=>"001000110",
  48403=>"101101101",
  48404=>"010000100",
  48405=>"101110111",
  48406=>"100101100",
  48407=>"110000111",
  48408=>"011001010",
  48409=>"100001000",
  48410=>"000010000",
  48411=>"101000011",
  48412=>"010001110",
  48413=>"100100110",
  48414=>"001101010",
  48415=>"111111110",
  48416=>"110100000",
  48417=>"011010000",
  48418=>"111111101",
  48419=>"000001010",
  48420=>"101100010",
  48421=>"100100100",
  48422=>"111011110",
  48423=>"000110111",
  48424=>"101111011",
  48425=>"111110001",
  48426=>"011001001",
  48427=>"000100000",
  48428=>"111000110",
  48429=>"010010110",
  48430=>"101100000",
  48431=>"001111101",
  48432=>"100100011",
  48433=>"111101010",
  48434=>"000011001",
  48435=>"111111110",
  48436=>"111101000",
  48437=>"100010011",
  48438=>"101011100",
  48439=>"101101010",
  48440=>"000010111",
  48441=>"101111101",
  48442=>"010011111",
  48443=>"011101101",
  48444=>"100111101",
  48445=>"011101010",
  48446=>"101111001",
  48447=>"010110100",
  48448=>"011110111",
  48449=>"010110000",
  48450=>"110111110",
  48451=>"111100001",
  48452=>"110000111",
  48453=>"010010001",
  48454=>"010110010",
  48455=>"000001000",
  48456=>"101101000",
  48457=>"010010000",
  48458=>"111110000",
  48459=>"011001101",
  48460=>"000011111",
  48461=>"100110100",
  48462=>"100101100",
  48463=>"000000010",
  48464=>"101111001",
  48465=>"011000001",
  48466=>"000000000",
  48467=>"010000000",
  48468=>"010110101",
  48469=>"101111110",
  48470=>"001100100",
  48471=>"011010101",
  48472=>"111100101",
  48473=>"101100010",
  48474=>"011111110",
  48475=>"100111000",
  48476=>"001001101",
  48477=>"101010011",
  48478=>"101101111",
  48479=>"110011111",
  48480=>"001110011",
  48481=>"101101110",
  48482=>"010101010",
  48483=>"110101110",
  48484=>"100110100",
  48485=>"010001101",
  48486=>"000101100",
  48487=>"011111100",
  48488=>"110000010",
  48489=>"001110001",
  48490=>"011001011",
  48491=>"101101100",
  48492=>"110001010",
  48493=>"100000101",
  48494=>"100101101",
  48495=>"110110100",
  48496=>"000110110",
  48497=>"011000001",
  48498=>"001010110",
  48499=>"110101111",
  48500=>"011101000",
  48501=>"101110010",
  48502=>"011010101",
  48503=>"111010100",
  48504=>"111101100",
  48505=>"110110110",
  48506=>"010101110",
  48507=>"111000101",
  48508=>"011111000",
  48509=>"110001000",
  48510=>"010111010",
  48511=>"111001000",
  48512=>"001001011",
  48513=>"001001110",
  48514=>"101001111",
  48515=>"000101001",
  48516=>"110110101",
  48517=>"001110010",
  48518=>"111100010",
  48519=>"101101110",
  48520=>"101111010",
  48521=>"111110110",
  48522=>"111110100",
  48523=>"001010110",
  48524=>"101010000",
  48525=>"110111100",
  48526=>"101101100",
  48527=>"000001100",
  48528=>"010100101",
  48529=>"100011111",
  48530=>"100101011",
  48531=>"111001110",
  48532=>"110100000",
  48533=>"100111110",
  48534=>"011001011",
  48535=>"101100000",
  48536=>"000110000",
  48537=>"000111100",
  48538=>"000010111",
  48539=>"010001011",
  48540=>"000111100",
  48541=>"000110110",
  48542=>"010001101",
  48543=>"000001011",
  48544=>"111010111",
  48545=>"100000010",
  48546=>"010010110",
  48547=>"100001101",
  48548=>"010111100",
  48549=>"100001101",
  48550=>"100111000",
  48551=>"001100000",
  48552=>"100001010",
  48553=>"011101011",
  48554=>"001001100",
  48555=>"000101010",
  48556=>"110111011",
  48557=>"011011000",
  48558=>"000010000",
  48559=>"001001101",
  48560=>"010000100",
  48561=>"110001110",
  48562=>"110001011",
  48563=>"110101101",
  48564=>"001000100",
  48565=>"001001001",
  48566=>"011011001",
  48567=>"100100001",
  48568=>"000000100",
  48569=>"111100001",
  48570=>"000000011",
  48571=>"100010010",
  48572=>"111011001",
  48573=>"110110111",
  48574=>"000101100",
  48575=>"011000000",
  48576=>"001011011",
  48577=>"000100000",
  48578=>"000101011",
  48579=>"101111001",
  48580=>"100111010",
  48581=>"101011101",
  48582=>"101011110",
  48583=>"011010000",
  48584=>"001101111",
  48585=>"000011111",
  48586=>"100011110",
  48587=>"101101100",
  48588=>"011011010",
  48589=>"111001000",
  48590=>"001101110",
  48591=>"110111110",
  48592=>"000111010",
  48593=>"011100110",
  48594=>"110001101",
  48595=>"011110111",
  48596=>"111010101",
  48597=>"000011010",
  48598=>"000001000",
  48599=>"010000000",
  48600=>"111011001",
  48601=>"010001010",
  48602=>"010100101",
  48603=>"110010011",
  48604=>"001100110",
  48605=>"001111000",
  48606=>"000000110",
  48607=>"110010001",
  48608=>"000111110",
  48609=>"111111010",
  48610=>"101100100",
  48611=>"011100001",
  48612=>"111100100",
  48613=>"000011011",
  48614=>"011010000",
  48615=>"010000100",
  48616=>"111101111",
  48617=>"001000011",
  48618=>"010111011",
  48619=>"111111001",
  48620=>"001110101",
  48621=>"111010011",
  48622=>"111110110",
  48623=>"101001000",
  48624=>"011100010",
  48625=>"011011111",
  48626=>"111101110",
  48627=>"011101100",
  48628=>"011111011",
  48629=>"010100000",
  48630=>"101011010",
  48631=>"101101101",
  48632=>"000010111",
  48633=>"111100110",
  48634=>"111101000",
  48635=>"001110111",
  48636=>"100101000",
  48637=>"111101000",
  48638=>"011110001",
  48639=>"011110100",
  48640=>"110100111",
  48641=>"011110011",
  48642=>"010010011",
  48643=>"010100000",
  48644=>"000011101",
  48645=>"011100010",
  48646=>"010001010",
  48647=>"010001001",
  48648=>"000000000",
  48649=>"001101100",
  48650=>"010100111",
  48651=>"001010100",
  48652=>"101011000",
  48653=>"111001111",
  48654=>"100001011",
  48655=>"000100000",
  48656=>"000101111",
  48657=>"001000111",
  48658=>"110001011",
  48659=>"100111100",
  48660=>"000111010",
  48661=>"101011100",
  48662=>"010010110",
  48663=>"000011100",
  48664=>"110001100",
  48665=>"111010000",
  48666=>"100111001",
  48667=>"100011000",
  48668=>"100010010",
  48669=>"000011100",
  48670=>"011011111",
  48671=>"100100000",
  48672=>"111111011",
  48673=>"101011111",
  48674=>"101100011",
  48675=>"001100011",
  48676=>"101000011",
  48677=>"001111111",
  48678=>"001100100",
  48679=>"010010100",
  48680=>"101110000",
  48681=>"011000001",
  48682=>"110101001",
  48683=>"111110101",
  48684=>"111111101",
  48685=>"011001001",
  48686=>"001111110",
  48687=>"101000100",
  48688=>"010010000",
  48689=>"000011000",
  48690=>"111001101",
  48691=>"101011101",
  48692=>"101000111",
  48693=>"010100111",
  48694=>"001000000",
  48695=>"010110101",
  48696=>"100101110",
  48697=>"001101110",
  48698=>"111110111",
  48699=>"000000101",
  48700=>"101101010",
  48701=>"001011010",
  48702=>"010110001",
  48703=>"101011001",
  48704=>"101001101",
  48705=>"101000000",
  48706=>"100011000",
  48707=>"111111011",
  48708=>"000000100",
  48709=>"100111101",
  48710=>"000101000",
  48711=>"110010010",
  48712=>"110001101",
  48713=>"000111001",
  48714=>"100101001",
  48715=>"010100000",
  48716=>"110111111",
  48717=>"010011001",
  48718=>"010101111",
  48719=>"100001111",
  48720=>"100110011",
  48721=>"101111101",
  48722=>"101111111",
  48723=>"000100011",
  48724=>"101010011",
  48725=>"110110010",
  48726=>"101110010",
  48727=>"000010100",
  48728=>"001101110",
  48729=>"000011011",
  48730=>"011101100",
  48731=>"111011100",
  48732=>"110100100",
  48733=>"110011110",
  48734=>"001001000",
  48735=>"000010110",
  48736=>"110001011",
  48737=>"000011100",
  48738=>"001111111",
  48739=>"100001011",
  48740=>"010100000",
  48741=>"000011100",
  48742=>"110001000",
  48743=>"011101001",
  48744=>"100110010",
  48745=>"111111010",
  48746=>"111001011",
  48747=>"010110100",
  48748=>"010001110",
  48749=>"111011111",
  48750=>"100100111",
  48751=>"010011111",
  48752=>"011101100",
  48753=>"000010010",
  48754=>"110110101",
  48755=>"111110011",
  48756=>"100110100",
  48757=>"111010000",
  48758=>"011000000",
  48759=>"101101111",
  48760=>"101010111",
  48761=>"001101000",
  48762=>"110100011",
  48763=>"011100100",
  48764=>"100011001",
  48765=>"111111100",
  48766=>"010100001",
  48767=>"001100101",
  48768=>"000001010",
  48769=>"001011000",
  48770=>"110100000",
  48771=>"001101010",
  48772=>"101010000",
  48773=>"011010100",
  48774=>"101010011",
  48775=>"111010001",
  48776=>"000110111",
  48777=>"100000011",
  48778=>"011110011",
  48779=>"110100110",
  48780=>"101000010",
  48781=>"011011110",
  48782=>"000001000",
  48783=>"111110001",
  48784=>"101110100",
  48785=>"011100001",
  48786=>"101001110",
  48787=>"000101000",
  48788=>"110100101",
  48789=>"101100101",
  48790=>"000001001",
  48791=>"000101010",
  48792=>"010010111",
  48793=>"011101000",
  48794=>"010011011",
  48795=>"111011100",
  48796=>"011101111",
  48797=>"100101101",
  48798=>"000001101",
  48799=>"011101011",
  48800=>"011011000",
  48801=>"000111111",
  48802=>"000100110",
  48803=>"001101110",
  48804=>"010011110",
  48805=>"000110011",
  48806=>"001011000",
  48807=>"111000000",
  48808=>"001000000",
  48809=>"000010110",
  48810=>"101101101",
  48811=>"011011010",
  48812=>"001110111",
  48813=>"011111010",
  48814=>"101100011",
  48815=>"111101111",
  48816=>"100010001",
  48817=>"100000001",
  48818=>"100010000",
  48819=>"010101001",
  48820=>"001000101",
  48821=>"011100010",
  48822=>"010010000",
  48823=>"011101000",
  48824=>"101101100",
  48825=>"100011101",
  48826=>"111110000",
  48827=>"110010110",
  48828=>"100101101",
  48829=>"101100010",
  48830=>"111011001",
  48831=>"000110010",
  48832=>"010100000",
  48833=>"100000100",
  48834=>"010100000",
  48835=>"101001101",
  48836=>"111000000",
  48837=>"101111010",
  48838=>"110001000",
  48839=>"000010001",
  48840=>"010111000",
  48841=>"011001110",
  48842=>"100100000",
  48843=>"001110001",
  48844=>"110101101",
  48845=>"001101001",
  48846=>"101000101",
  48847=>"000100010",
  48848=>"010111110",
  48849=>"000111110",
  48850=>"101110000",
  48851=>"000011100",
  48852=>"010000100",
  48853=>"001110000",
  48854=>"011010101",
  48855=>"000001111",
  48856=>"100100111",
  48857=>"000010100",
  48858=>"110001111",
  48859=>"000001001",
  48860=>"101001100",
  48861=>"001001001",
  48862=>"011000011",
  48863=>"011001110",
  48864=>"111010101",
  48865=>"011010011",
  48866=>"011111111",
  48867=>"111011111",
  48868=>"000100000",
  48869=>"010011010",
  48870=>"010000111",
  48871=>"000110000",
  48872=>"111010011",
  48873=>"011110111",
  48874=>"010011101",
  48875=>"011111001",
  48876=>"011111000",
  48877=>"001010111",
  48878=>"100010111",
  48879=>"101010000",
  48880=>"111000001",
  48881=>"000011010",
  48882=>"010010000",
  48883=>"101111111",
  48884=>"110000100",
  48885=>"010010011",
  48886=>"101110110",
  48887=>"101111101",
  48888=>"111010010",
  48889=>"000110101",
  48890=>"010110000",
  48891=>"100011010",
  48892=>"000000001",
  48893=>"000000000",
  48894=>"101001011",
  48895=>"000010000",
  48896=>"111100100",
  48897=>"100100000",
  48898=>"010011111",
  48899=>"111001010",
  48900=>"011110011",
  48901=>"000101000",
  48902=>"010101100",
  48903=>"000101001",
  48904=>"100000010",
  48905=>"011110110",
  48906=>"111010111",
  48907=>"001111110",
  48908=>"100001111",
  48909=>"011111011",
  48910=>"100010111",
  48911=>"111000101",
  48912=>"100001001",
  48913=>"111001101",
  48914=>"100001100",
  48915=>"011110011",
  48916=>"001100000",
  48917=>"011001111",
  48918=>"010101000",
  48919=>"101011101",
  48920=>"010111000",
  48921=>"100010000",
  48922=>"010100001",
  48923=>"101100110",
  48924=>"111000001",
  48925=>"110100101",
  48926=>"001000110",
  48927=>"100100111",
  48928=>"100111111",
  48929=>"001100100",
  48930=>"110011010",
  48931=>"101110100",
  48932=>"001000011",
  48933=>"000110101",
  48934=>"000101100",
  48935=>"011100101",
  48936=>"100010111",
  48937=>"100011101",
  48938=>"000100110",
  48939=>"101010001",
  48940=>"010101010",
  48941=>"001010000",
  48942=>"100000111",
  48943=>"000001110",
  48944=>"011000001",
  48945=>"110001010",
  48946=>"010011111",
  48947=>"101101101",
  48948=>"111100001",
  48949=>"110001010",
  48950=>"100110010",
  48951=>"100100011",
  48952=>"110110000",
  48953=>"101000111",
  48954=>"111011100",
  48955=>"011101010",
  48956=>"010011000",
  48957=>"000000100",
  48958=>"100001100",
  48959=>"000110001",
  48960=>"000011101",
  48961=>"010011111",
  48962=>"010001011",
  48963=>"001000001",
  48964=>"111111101",
  48965=>"111000111",
  48966=>"110111001",
  48967=>"000000111",
  48968=>"111001000",
  48969=>"101001101",
  48970=>"011100001",
  48971=>"100010100",
  48972=>"100010010",
  48973=>"100001001",
  48974=>"100000110",
  48975=>"100001110",
  48976=>"010111100",
  48977=>"110000101",
  48978=>"100000111",
  48979=>"100001011",
  48980=>"011011000",
  48981=>"101001101",
  48982=>"000100101",
  48983=>"110111011",
  48984=>"000000111",
  48985=>"100001111",
  48986=>"010111001",
  48987=>"110111101",
  48988=>"000100100",
  48989=>"110010111",
  48990=>"011111011",
  48991=>"110110001",
  48992=>"101011000",
  48993=>"000010000",
  48994=>"101100100",
  48995=>"101111011",
  48996=>"100110111",
  48997=>"011010001",
  48998=>"100100110",
  48999=>"010110000",
  49000=>"001001001",
  49001=>"010100100",
  49002=>"000010000",
  49003=>"010000001",
  49004=>"000110010",
  49005=>"101000011",
  49006=>"111111010",
  49007=>"110011111",
  49008=>"100010101",
  49009=>"111111101",
  49010=>"100111001",
  49011=>"111111111",
  49012=>"011101000",
  49013=>"010111110",
  49014=>"110110100",
  49015=>"011011010",
  49016=>"100001000",
  49017=>"000001110",
  49018=>"000110111",
  49019=>"011011010",
  49020=>"000000101",
  49021=>"110101010",
  49022=>"000010011",
  49023=>"001100101",
  49024=>"011010111",
  49025=>"010100000",
  49026=>"101001010",
  49027=>"010111011",
  49028=>"101001001",
  49029=>"000010101",
  49030=>"101111111",
  49031=>"110011010",
  49032=>"100111011",
  49033=>"101011100",
  49034=>"001001010",
  49035=>"101111010",
  49036=>"111100001",
  49037=>"100010000",
  49038=>"010100010",
  49039=>"001111101",
  49040=>"111101011",
  49041=>"111110111",
  49042=>"010000110",
  49043=>"101110111",
  49044=>"110001010",
  49045=>"000101111",
  49046=>"010001010",
  49047=>"011101101",
  49048=>"000111110",
  49049=>"110111000",
  49050=>"000001000",
  49051=>"111000001",
  49052=>"001100111",
  49053=>"110101111",
  49054=>"110100100",
  49055=>"111101010",
  49056=>"111000101",
  49057=>"101110111",
  49058=>"010001000",
  49059=>"001010101",
  49060=>"011010001",
  49061=>"111110110",
  49062=>"010011010",
  49063=>"111000001",
  49064=>"010001110",
  49065=>"111001000",
  49066=>"111001110",
  49067=>"000010011",
  49068=>"110010100",
  49069=>"111000111",
  49070=>"001110110",
  49071=>"110011010",
  49072=>"010010011",
  49073=>"110001000",
  49074=>"000110110",
  49075=>"101101010",
  49076=>"101011010",
  49077=>"100100100",
  49078=>"010101001",
  49079=>"111101111",
  49080=>"101111110",
  49081=>"000110001",
  49082=>"110100101",
  49083=>"000000110",
  49084=>"110101010",
  49085=>"001000111",
  49086=>"100011111",
  49087=>"000100000",
  49088=>"100111101",
  49089=>"010001111",
  49090=>"010100000",
  49091=>"001111111",
  49092=>"001000111",
  49093=>"101001111",
  49094=>"101101011",
  49095=>"010101101",
  49096=>"110000000",
  49097=>"101111110",
  49098=>"000000110",
  49099=>"100001010",
  49100=>"000001011",
  49101=>"011101101",
  49102=>"111101100",
  49103=>"111110010",
  49104=>"010111111",
  49105=>"001111000",
  49106=>"010001001",
  49107=>"000100100",
  49108=>"010010000",
  49109=>"011100111",
  49110=>"000010111",
  49111=>"100101000",
  49112=>"100010000",
  49113=>"111010001",
  49114=>"110111111",
  49115=>"100001100",
  49116=>"000110101",
  49117=>"100101110",
  49118=>"111000111",
  49119=>"000111011",
  49120=>"011000000",
  49121=>"001011001",
  49122=>"111000100",
  49123=>"000111110",
  49124=>"110010001",
  49125=>"110101000",
  49126=>"110000001",
  49127=>"110010010",
  49128=>"010000000",
  49129=>"010000011",
  49130=>"111110010",
  49131=>"101101110",
  49132=>"111110000",
  49133=>"111101010",
  49134=>"000000011",
  49135=>"011101010",
  49136=>"000011001",
  49137=>"001010100",
  49138=>"000001001",
  49139=>"101111101",
  49140=>"000011100",
  49141=>"100001011",
  49142=>"001111100",
  49143=>"000010101",
  49144=>"011000110",
  49145=>"100000101",
  49146=>"010100100",
  49147=>"101100110",
  49148=>"000010010",
  49149=>"101111111",
  49150=>"011011000",
  49151=>"101001011",
  49152=>"111010101",
  49153=>"010000100",
  49154=>"111111010",
  49155=>"001001100",
  49156=>"100010100",
  49157=>"011010000",
  49158=>"110011101",
  49159=>"110001011",
  49160=>"111111110",
  49161=>"011110100",
  49162=>"010101000",
  49163=>"111000101",
  49164=>"111111110",
  49165=>"101010011",
  49166=>"011011011",
  49167=>"111100010",
  49168=>"100101110",
  49169=>"111111001",
  49170=>"111001001",
  49171=>"110101100",
  49172=>"111111001",
  49173=>"111100010",
  49174=>"000011010",
  49175=>"001111111",
  49176=>"111001000",
  49177=>"110011010",
  49178=>"100000110",
  49179=>"001101100",
  49180=>"010000101",
  49181=>"011110111",
  49182=>"001101101",
  49183=>"010100110",
  49184=>"111100110",
  49185=>"110101010",
  49186=>"100110000",
  49187=>"100101000",
  49188=>"000101111",
  49189=>"011010100",
  49190=>"011101110",
  49191=>"110111100",
  49192=>"000010000",
  49193=>"101101010",
  49194=>"110001010",
  49195=>"001011100",
  49196=>"110100011",
  49197=>"011110110",
  49198=>"001100110",
  49199=>"001000100",
  49200=>"011001100",
  49201=>"100000101",
  49202=>"010000111",
  49203=>"011001001",
  49204=>"001101100",
  49205=>"101000011",
  49206=>"111000110",
  49207=>"000001111",
  49208=>"010100001",
  49209=>"111001001",
  49210=>"000110001",
  49211=>"011001000",
  49212=>"110100011",
  49213=>"010100000",
  49214=>"111101101",
  49215=>"000001100",
  49216=>"001101100",
  49217=>"000100001",
  49218=>"000001000",
  49219=>"010011010",
  49220=>"000010001",
  49221=>"110100101",
  49222=>"101101000",
  49223=>"111110101",
  49224=>"100000001",
  49225=>"111011110",
  49226=>"010100001",
  49227=>"000000101",
  49228=>"111101100",
  49229=>"011000110",
  49230=>"111110100",
  49231=>"011001101",
  49232=>"111111100",
  49233=>"100000010",
  49234=>"110110101",
  49235=>"001110111",
  49236=>"101101011",
  49237=>"011000000",
  49238=>"110010011",
  49239=>"101011101",
  49240=>"010011100",
  49241=>"100001000",
  49242=>"111100001",
  49243=>"100010110",
  49244=>"010000000",
  49245=>"000111000",
  49246=>"000011001",
  49247=>"011110001",
  49248=>"000011010",
  49249=>"101111111",
  49250=>"000011111",
  49251=>"010101000",
  49252=>"000101000",
  49253=>"110101101",
  49254=>"110110111",
  49255=>"100110111",
  49256=>"010111110",
  49257=>"100000000",
  49258=>"110001011",
  49259=>"111111101",
  49260=>"110100010",
  49261=>"001010011",
  49262=>"111110101",
  49263=>"001011110",
  49264=>"110000110",
  49265=>"011011100",
  49266=>"101111001",
  49267=>"010010001",
  49268=>"111101010",
  49269=>"001101011",
  49270=>"001000110",
  49271=>"000110101",
  49272=>"100000011",
  49273=>"011111000",
  49274=>"100011100",
  49275=>"101011110",
  49276=>"000100010",
  49277=>"000000001",
  49278=>"101101011",
  49279=>"001101101",
  49280=>"011011101",
  49281=>"111000001",
  49282=>"000000111",
  49283=>"101001010",
  49284=>"001100111",
  49285=>"001111111",
  49286=>"011100101",
  49287=>"100000101",
  49288=>"010100111",
  49289=>"111011010",
  49290=>"110101101",
  49291=>"000101101",
  49292=>"110100110",
  49293=>"101100001",
  49294=>"100100111",
  49295=>"111101000",
  49296=>"100110100",
  49297=>"011011101",
  49298=>"000111000",
  49299=>"011001100",
  49300=>"111000111",
  49301=>"000100010",
  49302=>"001111001",
  49303=>"101010011",
  49304=>"000000100",
  49305=>"100101000",
  49306=>"101001100",
  49307=>"010000000",
  49308=>"101111111",
  49309=>"111101010",
  49310=>"111010000",
  49311=>"101101101",
  49312=>"011110111",
  49313=>"001100000",
  49314=>"100011010",
  49315=>"100100000",
  49316=>"110101111",
  49317=>"010011110",
  49318=>"011111110",
  49319=>"001011100",
  49320=>"000001101",
  49321=>"001011001",
  49322=>"011100010",
  49323=>"001110100",
  49324=>"110001010",
  49325=>"011001010",
  49326=>"011110110",
  49327=>"100101011",
  49328=>"100010110",
  49329=>"110011010",
  49330=>"001110101",
  49331=>"000000010",
  49332=>"110010010",
  49333=>"110001010",
  49334=>"011000100",
  49335=>"011111000",
  49336=>"000001110",
  49337=>"111100100",
  49338=>"001000000",
  49339=>"000001010",
  49340=>"111101000",
  49341=>"111001000",
  49342=>"110111110",
  49343=>"001111001",
  49344=>"101111011",
  49345=>"000011111",
  49346=>"100110110",
  49347=>"011001110",
  49348=>"110010000",
  49349=>"001100100",
  49350=>"011001001",
  49351=>"011100111",
  49352=>"010010011",
  49353=>"101111111",
  49354=>"000101110",
  49355=>"101011110",
  49356=>"101010001",
  49357=>"101111100",
  49358=>"011000011",
  49359=>"001000011",
  49360=>"001011110",
  49361=>"100110100",
  49362=>"110110101",
  49363=>"111101001",
  49364=>"100001010",
  49365=>"101001011",
  49366=>"000101010",
  49367=>"000101001",
  49368=>"100001001",
  49369=>"111010010",
  49370=>"000000101",
  49371=>"101000000",
  49372=>"001001000",
  49373=>"010000111",
  49374=>"101001011",
  49375=>"000110101",
  49376=>"100101110",
  49377=>"000101110",
  49378=>"011000010",
  49379=>"100010111",
  49380=>"010011110",
  49381=>"101110111",
  49382=>"101100011",
  49383=>"010001111",
  49384=>"011001001",
  49385=>"100001000",
  49386=>"001011001",
  49387=>"011101001",
  49388=>"011110110",
  49389=>"000011111",
  49390=>"100001001",
  49391=>"010001100",
  49392=>"010010101",
  49393=>"100011100",
  49394=>"000010011",
  49395=>"010011001",
  49396=>"011000111",
  49397=>"000110010",
  49398=>"000001111",
  49399=>"101101111",
  49400=>"000001010",
  49401=>"110110100",
  49402=>"100010111",
  49403=>"100101101",
  49404=>"110000000",
  49405=>"101011000",
  49406=>"011111000",
  49407=>"101111000",
  49408=>"111001111",
  49409=>"111001100",
  49410=>"000101111",
  49411=>"000100001",
  49412=>"010101111",
  49413=>"001010010",
  49414=>"100111011",
  49415=>"000010000",
  49416=>"100101111",
  49417=>"111010001",
  49418=>"100111011",
  49419=>"010110111",
  49420=>"000100100",
  49421=>"111101100",
  49422=>"110001111",
  49423=>"010001011",
  49424=>"110101001",
  49425=>"100011000",
  49426=>"010101101",
  49427=>"011000000",
  49428=>"101101001",
  49429=>"010011010",
  49430=>"000110111",
  49431=>"111110011",
  49432=>"010011001",
  49433=>"101000001",
  49434=>"110110000",
  49435=>"111001001",
  49436=>"001001000",
  49437=>"010110111",
  49438=>"100010000",
  49439=>"000110000",
  49440=>"001000101",
  49441=>"111111010",
  49442=>"010011111",
  49443=>"001011000",
  49444=>"010110011",
  49445=>"111000011",
  49446=>"000000101",
  49447=>"101101000",
  49448=>"010101000",
  49449=>"111001010",
  49450=>"100101100",
  49451=>"010111010",
  49452=>"001100001",
  49453=>"010111101",
  49454=>"011010101",
  49455=>"111101011",
  49456=>"100100111",
  49457=>"011110101",
  49458=>"110100000",
  49459=>"000001001",
  49460=>"010101010",
  49461=>"101100111",
  49462=>"111001100",
  49463=>"100110000",
  49464=>"111001101",
  49465=>"001111111",
  49466=>"111011100",
  49467=>"001011010",
  49468=>"111101101",
  49469=>"111111010",
  49470=>"110001000",
  49471=>"110000110",
  49472=>"010100111",
  49473=>"001000001",
  49474=>"011110110",
  49475=>"011111111",
  49476=>"101101001",
  49477=>"101010101",
  49478=>"001100010",
  49479=>"111010001",
  49480=>"001011000",
  49481=>"100101010",
  49482=>"000111101",
  49483=>"100000100",
  49484=>"110100001",
  49485=>"101001011",
  49486=>"101101110",
  49487=>"110100110",
  49488=>"100001101",
  49489=>"101000100",
  49490=>"110101000",
  49491=>"101100100",
  49492=>"101110111",
  49493=>"001100010",
  49494=>"101111100",
  49495=>"000110010",
  49496=>"110010100",
  49497=>"001101101",
  49498=>"101000010",
  49499=>"001100001",
  49500=>"000111010",
  49501=>"000111110",
  49502=>"000011011",
  49503=>"111100111",
  49504=>"100111011",
  49505=>"011011000",
  49506=>"101110101",
  49507=>"101111111",
  49508=>"010010101",
  49509=>"000110011",
  49510=>"100010001",
  49511=>"000110010",
  49512=>"010001010",
  49513=>"101011001",
  49514=>"001010101",
  49515=>"001010111",
  49516=>"000010010",
  49517=>"101110001",
  49518=>"110100010",
  49519=>"100000110",
  49520=>"000111000",
  49521=>"110011001",
  49522=>"101010000",
  49523=>"110111110",
  49524=>"011001111",
  49525=>"010011000",
  49526=>"111111111",
  49527=>"001111010",
  49528=>"010111001",
  49529=>"010110010",
  49530=>"100001011",
  49531=>"001010000",
  49532=>"010011001",
  49533=>"111110110",
  49534=>"010111100",
  49535=>"100110001",
  49536=>"000101100",
  49537=>"110101011",
  49538=>"001100110",
  49539=>"110101110",
  49540=>"110001001",
  49541=>"001010000",
  49542=>"010010110",
  49543=>"110101111",
  49544=>"101000011",
  49545=>"011101101",
  49546=>"000011010",
  49547=>"110101101",
  49548=>"111010000",
  49549=>"101101100",
  49550=>"100111101",
  49551=>"010101010",
  49552=>"010000010",
  49553=>"111101111",
  49554=>"010001010",
  49555=>"111000011",
  49556=>"110111010",
  49557=>"100000010",
  49558=>"100100001",
  49559=>"111010101",
  49560=>"101111100",
  49561=>"101100100",
  49562=>"101010001",
  49563=>"011000000",
  49564=>"100001100",
  49565=>"100001100",
  49566=>"101101110",
  49567=>"110010011",
  49568=>"101100111",
  49569=>"111110110",
  49570=>"001011011",
  49571=>"001110001",
  49572=>"111010011",
  49573=>"000100101",
  49574=>"011001111",
  49575=>"100111101",
  49576=>"000011001",
  49577=>"000010011",
  49578=>"001111001",
  49579=>"111000001",
  49580=>"010100100",
  49581=>"010111011",
  49582=>"110000001",
  49583=>"000100010",
  49584=>"111101101",
  49585=>"110110111",
  49586=>"100101101",
  49587=>"011000011",
  49588=>"011010000",
  49589=>"011110000",
  49590=>"100111011",
  49591=>"011000000",
  49592=>"010000010",
  49593=>"001000010",
  49594=>"011011000",
  49595=>"011110010",
  49596=>"110011101",
  49597=>"010010010",
  49598=>"110000101",
  49599=>"010111011",
  49600=>"101001110",
  49601=>"000000000",
  49602=>"100111110",
  49603=>"011110101",
  49604=>"000100010",
  49605=>"111011000",
  49606=>"011000011",
  49607=>"110100001",
  49608=>"100011000",
  49609=>"001101011",
  49610=>"111100111",
  49611=>"111010010",
  49612=>"010111010",
  49613=>"111101001",
  49614=>"110010010",
  49615=>"101101011",
  49616=>"100110111",
  49617=>"111000111",
  49618=>"011101001",
  49619=>"001001101",
  49620=>"100011110",
  49621=>"010111110",
  49622=>"001000110",
  49623=>"111100101",
  49624=>"101001001",
  49625=>"010001101",
  49626=>"000101111",
  49627=>"100010111",
  49628=>"111011101",
  49629=>"100101001",
  49630=>"111110111",
  49631=>"011101111",
  49632=>"111100101",
  49633=>"001101110",
  49634=>"100110111",
  49635=>"000111110",
  49636=>"100011000",
  49637=>"101000000",
  49638=>"011110010",
  49639=>"111011111",
  49640=>"000010001",
  49641=>"011110100",
  49642=>"010010111",
  49643=>"101011001",
  49644=>"111000110",
  49645=>"011010000",
  49646=>"111100000",
  49647=>"011000011",
  49648=>"110110101",
  49649=>"011011011",
  49650=>"000000010",
  49651=>"110001110",
  49652=>"100100101",
  49653=>"010100111",
  49654=>"001100101",
  49655=>"101110011",
  49656=>"100011110",
  49657=>"100010010",
  49658=>"111001111",
  49659=>"100011011",
  49660=>"101111001",
  49661=>"100011010",
  49662=>"011100010",
  49663=>"100010000",
  49664=>"011110010",
  49665=>"000001000",
  49666=>"101101110",
  49667=>"011110101",
  49668=>"111100001",
  49669=>"110100111",
  49670=>"100101111",
  49671=>"010001101",
  49672=>"000101111",
  49673=>"000111100",
  49674=>"110000001",
  49675=>"001000010",
  49676=>"100110100",
  49677=>"000111110",
  49678=>"110000000",
  49679=>"000001011",
  49680=>"111101110",
  49681=>"110110000",
  49682=>"100011000",
  49683=>"010111010",
  49684=>"010111110",
  49685=>"100010010",
  49686=>"011001011",
  49687=>"000110111",
  49688=>"001001100",
  49689=>"011101110",
  49690=>"010101010",
  49691=>"011000111",
  49692=>"100110100",
  49693=>"111000000",
  49694=>"111110100",
  49695=>"010101101",
  49696=>"100000100",
  49697=>"010101001",
  49698=>"101101010",
  49699=>"111100001",
  49700=>"101111111",
  49701=>"110100101",
  49702=>"010000001",
  49703=>"100110101",
  49704=>"000001110",
  49705=>"101110101",
  49706=>"101110111",
  49707=>"100011000",
  49708=>"011110001",
  49709=>"110011000",
  49710=>"011011111",
  49711=>"111110101",
  49712=>"000011011",
  49713=>"110101011",
  49714=>"101111010",
  49715=>"101101101",
  49716=>"100000111",
  49717=>"100010010",
  49718=>"001110111",
  49719=>"011100010",
  49720=>"110010001",
  49721=>"111101011",
  49722=>"000010010",
  49723=>"100111011",
  49724=>"011000100",
  49725=>"110011111",
  49726=>"001011101",
  49727=>"110010111",
  49728=>"111101001",
  49729=>"001001110",
  49730=>"101000100",
  49731=>"000111101",
  49732=>"111110111",
  49733=>"111110110",
  49734=>"110100111",
  49735=>"001100111",
  49736=>"001110011",
  49737=>"001101011",
  49738=>"101010011",
  49739=>"100100011",
  49740=>"000010110",
  49741=>"110100100",
  49742=>"001101110",
  49743=>"011000100",
  49744=>"001111101",
  49745=>"101001111",
  49746=>"111111101",
  49747=>"010011001",
  49748=>"111011111",
  49749=>"001000001",
  49750=>"101001101",
  49751=>"000001011",
  49752=>"100110100",
  49753=>"000001110",
  49754=>"101001000",
  49755=>"001100000",
  49756=>"101110010",
  49757=>"101110000",
  49758=>"000110001",
  49759=>"100110001",
  49760=>"000001001",
  49761=>"100111000",
  49762=>"011101011",
  49763=>"000011001",
  49764=>"111000101",
  49765=>"101010111",
  49766=>"111101001",
  49767=>"011000001",
  49768=>"011110111",
  49769=>"000111110",
  49770=>"000111101",
  49771=>"100100001",
  49772=>"100100101",
  49773=>"110101001",
  49774=>"101111010",
  49775=>"110001001",
  49776=>"000010011",
  49777=>"001110110",
  49778=>"000110010",
  49779=>"101101001",
  49780=>"011111111",
  49781=>"100010001",
  49782=>"111111100",
  49783=>"000101001",
  49784=>"111101011",
  49785=>"100111011",
  49786=>"101001011",
  49787=>"010001100",
  49788=>"000010000",
  49789=>"011111011",
  49790=>"111100110",
  49791=>"000111111",
  49792=>"000011100",
  49793=>"101011001",
  49794=>"100100011",
  49795=>"001010110",
  49796=>"000010100",
  49797=>"000100010",
  49798=>"001010000",
  49799=>"000100000",
  49800=>"100000100",
  49801=>"100110100",
  49802=>"010000010",
  49803=>"000100001",
  49804=>"001010111",
  49805=>"011011101",
  49806=>"011110100",
  49807=>"011101111",
  49808=>"110111011",
  49809=>"110111111",
  49810=>"000101010",
  49811=>"001000000",
  49812=>"010011000",
  49813=>"111001011",
  49814=>"001010010",
  49815=>"101011000",
  49816=>"110110010",
  49817=>"101000001",
  49818=>"100100101",
  49819=>"101101010",
  49820=>"111110100",
  49821=>"110000001",
  49822=>"001100100",
  49823=>"000010011",
  49824=>"100110011",
  49825=>"100000011",
  49826=>"111001111",
  49827=>"000100010",
  49828=>"000100110",
  49829=>"000001010",
  49830=>"001100100",
  49831=>"100000011",
  49832=>"010011000",
  49833=>"011111001",
  49834=>"010010011",
  49835=>"011010001",
  49836=>"010011010",
  49837=>"000000011",
  49838=>"111101100",
  49839=>"011011000",
  49840=>"000000010",
  49841=>"100101011",
  49842=>"110101010",
  49843=>"111000011",
  49844=>"111101010",
  49845=>"010010001",
  49846=>"001100000",
  49847=>"101010100",
  49848=>"110110011",
  49849=>"100101001",
  49850=>"100111000",
  49851=>"101010100",
  49852=>"111000000",
  49853=>"011001101",
  49854=>"000100111",
  49855=>"100110101",
  49856=>"101100001",
  49857=>"010100110",
  49858=>"001110010",
  49859=>"101001110",
  49860=>"010000110",
  49861=>"010110011",
  49862=>"000011010",
  49863=>"111101011",
  49864=>"101001011",
  49865=>"001011100",
  49866=>"100101110",
  49867=>"001011110",
  49868=>"000110011",
  49869=>"110000010",
  49870=>"101111101",
  49871=>"000011000",
  49872=>"011111101",
  49873=>"011100110",
  49874=>"100001110",
  49875=>"001011000",
  49876=>"000101101",
  49877=>"001111011",
  49878=>"101111011",
  49879=>"100110101",
  49880=>"101111101",
  49881=>"110111110",
  49882=>"010100111",
  49883=>"000000101",
  49884=>"000011110",
  49885=>"010101111",
  49886=>"011001000",
  49887=>"101110101",
  49888=>"110001011",
  49889=>"011101000",
  49890=>"000011011",
  49891=>"001001000",
  49892=>"000011011",
  49893=>"111000110",
  49894=>"011101101",
  49895=>"001010011",
  49896=>"000110111",
  49897=>"000100111",
  49898=>"000101011",
  49899=>"110001100",
  49900=>"000000001",
  49901=>"110111110",
  49902=>"101011001",
  49903=>"101010011",
  49904=>"111111011",
  49905=>"110000111",
  49906=>"011011001",
  49907=>"001110010",
  49908=>"101001001",
  49909=>"011100110",
  49910=>"110001111",
  49911=>"010010010",
  49912=>"011010111",
  49913=>"110100010",
  49914=>"101111001",
  49915=>"010101001",
  49916=>"110001000",
  49917=>"111100101",
  49918=>"100011001",
  49919=>"010101000",
  49920=>"011010100",
  49921=>"111111111",
  49922=>"110111011",
  49923=>"000100111",
  49924=>"001111000",
  49925=>"001000000",
  49926=>"110100011",
  49927=>"011000110",
  49928=>"100011111",
  49929=>"001111111",
  49930=>"011100101",
  49931=>"100111001",
  49932=>"010000000",
  49933=>"101101011",
  49934=>"111001101",
  49935=>"011111010",
  49936=>"000100010",
  49937=>"110101110",
  49938=>"100111000",
  49939=>"010010011",
  49940=>"101101000",
  49941=>"000010010",
  49942=>"011000100",
  49943=>"010101000",
  49944=>"101101101",
  49945=>"011001111",
  49946=>"000010011",
  49947=>"101100000",
  49948=>"111101000",
  49949=>"001010100",
  49950=>"111101000",
  49951=>"000110000",
  49952=>"011000010",
  49953=>"010000000",
  49954=>"101001000",
  49955=>"111001111",
  49956=>"010001010",
  49957=>"000001100",
  49958=>"000110110",
  49959=>"111001101",
  49960=>"011001111",
  49961=>"010100100",
  49962=>"110100110",
  49963=>"101100111",
  49964=>"001000010",
  49965=>"111010111",
  49966=>"100000110",
  49967=>"100110100",
  49968=>"110011100",
  49969=>"011101111",
  49970=>"001101101",
  49971=>"111000000",
  49972=>"001101000",
  49973=>"010000110",
  49974=>"110001000",
  49975=>"101001100",
  49976=>"100010000",
  49977=>"010001010",
  49978=>"001011110",
  49979=>"110101010",
  49980=>"001101001",
  49981=>"001001111",
  49982=>"110100101",
  49983=>"100010101",
  49984=>"011110111",
  49985=>"001001010",
  49986=>"110000100",
  49987=>"011100101",
  49988=>"111100011",
  49989=>"011000011",
  49990=>"001001101",
  49991=>"111001110",
  49992=>"000101001",
  49993=>"110011000",
  49994=>"001100111",
  49995=>"101001000",
  49996=>"111101110",
  49997=>"111111110",
  49998=>"111100000",
  49999=>"011010101",
  50000=>"110100100",
  50001=>"101101110",
  50002=>"111101001",
  50003=>"110011111",
  50004=>"101100100",
  50005=>"011001011",
  50006=>"000000100",
  50007=>"010101100",
  50008=>"111000010",
  50009=>"110100011",
  50010=>"101100101",
  50011=>"000101000",
  50012=>"001100100",
  50013=>"001101100",
  50014=>"010100000",
  50015=>"010001100",
  50016=>"100011111",
  50017=>"000101000",
  50018=>"101000100",
  50019=>"111111010",
  50020=>"011101010",
  50021=>"110011110",
  50022=>"101001101",
  50023=>"011110010",
  50024=>"110110011",
  50025=>"100101010",
  50026=>"000111000",
  50027=>"001111100",
  50028=>"001110111",
  50029=>"001001110",
  50030=>"001101110",
  50031=>"010000010",
  50032=>"100001111",
  50033=>"111111010",
  50034=>"010110010",
  50035=>"110000111",
  50036=>"001001000",
  50037=>"010011000",
  50038=>"100000011",
  50039=>"011000101",
  50040=>"101100010",
  50041=>"111100100",
  50042=>"001111101",
  50043=>"011000000",
  50044=>"111100110",
  50045=>"000001010",
  50046=>"100110101",
  50047=>"101010000",
  50048=>"000011000",
  50049=>"110111000",
  50050=>"101111000",
  50051=>"001010001",
  50052=>"000011010",
  50053=>"001111001",
  50054=>"000111100",
  50055=>"111000001",
  50056=>"001101011",
  50057=>"000111000",
  50058=>"010111010",
  50059=>"001001110",
  50060=>"100001010",
  50061=>"011001001",
  50062=>"011110111",
  50063=>"111111101",
  50064=>"010000110",
  50065=>"011011010",
  50066=>"110100011",
  50067=>"110011100",
  50068=>"010001000",
  50069=>"110010111",
  50070=>"101011101",
  50071=>"011011101",
  50072=>"000101101",
  50073=>"100001110",
  50074=>"111010000",
  50075=>"110111101",
  50076=>"001011100",
  50077=>"011101101",
  50078=>"010011111",
  50079=>"001101101",
  50080=>"101101111",
  50081=>"111101100",
  50082=>"010000101",
  50083=>"100000101",
  50084=>"001001111",
  50085=>"010100100",
  50086=>"001111110",
  50087=>"011111101",
  50088=>"001011101",
  50089=>"100000110",
  50090=>"110011111",
  50091=>"101100101",
  50092=>"001101011",
  50093=>"111010011",
  50094=>"010110101",
  50095=>"101101001",
  50096=>"000100101",
  50097=>"110110101",
  50098=>"000110100",
  50099=>"010011011",
  50100=>"100011100",
  50101=>"101111111",
  50102=>"101110000",
  50103=>"000001010",
  50104=>"101001110",
  50105=>"001110111",
  50106=>"001000000",
  50107=>"010101010",
  50108=>"001110111",
  50109=>"001101100",
  50110=>"100100001",
  50111=>"110101101",
  50112=>"100100001",
  50113=>"011011111",
  50114=>"111000001",
  50115=>"111110000",
  50116=>"100010110",
  50117=>"111000110",
  50118=>"000010010",
  50119=>"010000100",
  50120=>"101001000",
  50121=>"111100000",
  50122=>"101101110",
  50123=>"001000011",
  50124=>"111100000",
  50125=>"001110000",
  50126=>"010101100",
  50127=>"001100111",
  50128=>"011110101",
  50129=>"101011101",
  50130=>"000110110",
  50131=>"011000001",
  50132=>"010000010",
  50133=>"100110111",
  50134=>"000110000",
  50135=>"000010010",
  50136=>"110111011",
  50137=>"100001101",
  50138=>"101000011",
  50139=>"101100010",
  50140=>"100011000",
  50141=>"001101000",
  50142=>"011100100",
  50143=>"100100100",
  50144=>"100110000",
  50145=>"001010011",
  50146=>"011010010",
  50147=>"100011110",
  50148=>"001110011",
  50149=>"110101111",
  50150=>"010001111",
  50151=>"111000111",
  50152=>"001110100",
  50153=>"101010101",
  50154=>"111000010",
  50155=>"110100010",
  50156=>"000100010",
  50157=>"111111000",
  50158=>"100010110",
  50159=>"111001001",
  50160=>"101001110",
  50161=>"000011000",
  50162=>"001000011",
  50163=>"101010000",
  50164=>"110000100",
  50165=>"010011001",
  50166=>"110100010",
  50167=>"000010100",
  50168=>"011010100",
  50169=>"001110001",
  50170=>"010110000",
  50171=>"010110100",
  50172=>"010001100",
  50173=>"000111001",
  50174=>"101011111",
  50175=>"001011111",
  50176=>"011100000",
  50177=>"100000010",
  50178=>"010111101",
  50179=>"010110110",
  50180=>"000001010",
  50181=>"111000110",
  50182=>"100001010",
  50183=>"000010000",
  50184=>"000110110",
  50185=>"111001010",
  50186=>"011100101",
  50187=>"001110101",
  50188=>"111111110",
  50189=>"101100011",
  50190=>"001010001",
  50191=>"110011010",
  50192=>"100110000",
  50193=>"110001000",
  50194=>"011000010",
  50195=>"111011001",
  50196=>"111011011",
  50197=>"110001101",
  50198=>"000010101",
  50199=>"100000001",
  50200=>"000100110",
  50201=>"000001110",
  50202=>"001000010",
  50203=>"101000111",
  50204=>"010000101",
  50205=>"000000101",
  50206=>"010100011",
  50207=>"110011000",
  50208=>"101011011",
  50209=>"110010010",
  50210=>"100111100",
  50211=>"111101000",
  50212=>"101001101",
  50213=>"110010000",
  50214=>"000001100",
  50215=>"001010000",
  50216=>"010100111",
  50217=>"000000110",
  50218=>"100101001",
  50219=>"010110111",
  50220=>"100100101",
  50221=>"000111010",
  50222=>"110001010",
  50223=>"101000000",
  50224=>"101111101",
  50225=>"000001110",
  50226=>"001110111",
  50227=>"101101000",
  50228=>"000110100",
  50229=>"110100100",
  50230=>"110100001",
  50231=>"010110010",
  50232=>"101000101",
  50233=>"111010001",
  50234=>"111001011",
  50235=>"110011111",
  50236=>"001001000",
  50237=>"100000010",
  50238=>"001101000",
  50239=>"110111101",
  50240=>"110101011",
  50241=>"001000001",
  50242=>"110010010",
  50243=>"101110100",
  50244=>"010011101",
  50245=>"000000001",
  50246=>"110111001",
  50247=>"010101101",
  50248=>"101010110",
  50249=>"010000111",
  50250=>"000001010",
  50251=>"111000101",
  50252=>"010000111",
  50253=>"011001000",
  50254=>"011000000",
  50255=>"101101010",
  50256=>"101100111",
  50257=>"111101111",
  50258=>"000010110",
  50259=>"000000010",
  50260=>"001110110",
  50261=>"111110100",
  50262=>"001110100",
  50263=>"010111001",
  50264=>"001101111",
  50265=>"110111111",
  50266=>"101011000",
  50267=>"110000010",
  50268=>"111010101",
  50269=>"101000000",
  50270=>"100001010",
  50271=>"101000101",
  50272=>"010000001",
  50273=>"001110101",
  50274=>"111100100",
  50275=>"010000010",
  50276=>"110100010",
  50277=>"100001101",
  50278=>"100000100",
  50279=>"110110100",
  50280=>"011000100",
  50281=>"101011111",
  50282=>"110010111",
  50283=>"101110110",
  50284=>"111001111",
  50285=>"000000111",
  50286=>"101010010",
  50287=>"000101000",
  50288=>"101111101",
  50289=>"011101110",
  50290=>"111100110",
  50291=>"110110000",
  50292=>"100100110",
  50293=>"010101001",
  50294=>"000011110",
  50295=>"001000110",
  50296=>"010111111",
  50297=>"110111001",
  50298=>"110010100",
  50299=>"100000011",
  50300=>"000001011",
  50301=>"101010100",
  50302=>"001110000",
  50303=>"010011010",
  50304=>"001110000",
  50305=>"110000110",
  50306=>"110000001",
  50307=>"011011011",
  50308=>"011101111",
  50309=>"101010010",
  50310=>"001000110",
  50311=>"011100011",
  50312=>"001000101",
  50313=>"011001000",
  50314=>"011011000",
  50315=>"000000011",
  50316=>"101001111",
  50317=>"001100110",
  50318=>"110111111",
  50319=>"000101101",
  50320=>"101011010",
  50321=>"101111110",
  50322=>"000100000",
  50323=>"111100101",
  50324=>"000100100",
  50325=>"011100111",
  50326=>"000101001",
  50327=>"110001100",
  50328=>"010000000",
  50329=>"010011011",
  50330=>"011111110",
  50331=>"110010101",
  50332=>"101111111",
  50333=>"100000011",
  50334=>"011010010",
  50335=>"101001101",
  50336=>"100001111",
  50337=>"100100000",
  50338=>"101000101",
  50339=>"100011101",
  50340=>"010101001",
  50341=>"101100101",
  50342=>"101011001",
  50343=>"011100101",
  50344=>"011010110",
  50345=>"011011111",
  50346=>"100101001",
  50347=>"110100000",
  50348=>"101010111",
  50349=>"111001110",
  50350=>"101010101",
  50351=>"111101110",
  50352=>"010001001",
  50353=>"001011110",
  50354=>"001000001",
  50355=>"100000010",
  50356=>"000101100",
  50357=>"000101110",
  50358=>"011011100",
  50359=>"011111101",
  50360=>"001011010",
  50361=>"110011101",
  50362=>"100000110",
  50363=>"001110111",
  50364=>"001100101",
  50365=>"100100110",
  50366=>"001110011",
  50367=>"001011011",
  50368=>"010010010",
  50369=>"001010011",
  50370=>"100011001",
  50371=>"001001011",
  50372=>"010111101",
  50373=>"110101010",
  50374=>"100011110",
  50375=>"111000010",
  50376=>"010111110",
  50377=>"000101000",
  50378=>"111101001",
  50379=>"101110000",
  50380=>"101011000",
  50381=>"111000000",
  50382=>"000000001",
  50383=>"100001100",
  50384=>"011110011",
  50385=>"111111001",
  50386=>"110010110",
  50387=>"011000000",
  50388=>"111001001",
  50389=>"101101111",
  50390=>"001000011",
  50391=>"101110110",
  50392=>"010011000",
  50393=>"111010101",
  50394=>"011101011",
  50395=>"010111101",
  50396=>"101011001",
  50397=>"100101010",
  50398=>"000101011",
  50399=>"011011001",
  50400=>"101101110",
  50401=>"110100111",
  50402=>"011111001",
  50403=>"101111110",
  50404=>"010000110",
  50405=>"111101111",
  50406=>"011101011",
  50407=>"110001000",
  50408=>"100111111",
  50409=>"001000110",
  50410=>"100000100",
  50411=>"101101111",
  50412=>"100000001",
  50413=>"001110100",
  50414=>"101100010",
  50415=>"110011001",
  50416=>"110110100",
  50417=>"110011111",
  50418=>"000110100",
  50419=>"100011010",
  50420=>"001001100",
  50421=>"110001110",
  50422=>"011001101",
  50423=>"011100010",
  50424=>"010000000",
  50425=>"000001111",
  50426=>"111101000",
  50427=>"000100101",
  50428=>"011010011",
  50429=>"011010000",
  50430=>"010111100",
  50431=>"111001011",
  50432=>"100000001",
  50433=>"111110010",
  50434=>"111000111",
  50435=>"101110111",
  50436=>"111100000",
  50437=>"111111110",
  50438=>"001000001",
  50439=>"001110011",
  50440=>"011110011",
  50441=>"000010110",
  50442=>"111100100",
  50443=>"011100100",
  50444=>"011101100",
  50445=>"010100100",
  50446=>"101100001",
  50447=>"111101010",
  50448=>"000111010",
  50449=>"011111001",
  50450=>"110011001",
  50451=>"111100111",
  50452=>"111000100",
  50453=>"010100111",
  50454=>"010110100",
  50455=>"100111000",
  50456=>"010101110",
  50457=>"101110111",
  50458=>"010010100",
  50459=>"000110101",
  50460=>"100101110",
  50461=>"110101100",
  50462=>"011010100",
  50463=>"010000010",
  50464=>"100010010",
  50465=>"011111101",
  50466=>"101001100",
  50467=>"101001111",
  50468=>"010001011",
  50469=>"010010110",
  50470=>"001000010",
  50471=>"101011000",
  50472=>"010011000",
  50473=>"101010100",
  50474=>"100001000",
  50475=>"011010010",
  50476=>"101000101",
  50477=>"100000000",
  50478=>"010101111",
  50479=>"110011111",
  50480=>"100100111",
  50481=>"001110101",
  50482=>"100010101",
  50483=>"111010001",
  50484=>"000001101",
  50485=>"000000110",
  50486=>"100010011",
  50487=>"110001101",
  50488=>"100000011",
  50489=>"010001100",
  50490=>"110101000",
  50491=>"101001110",
  50492=>"110111100",
  50493=>"110111001",
  50494=>"110011101",
  50495=>"110110101",
  50496=>"101111010",
  50497=>"110111110",
  50498=>"011001000",
  50499=>"000011111",
  50500=>"010110010",
  50501=>"010101100",
  50502=>"000010011",
  50503=>"011111001",
  50504=>"110100100",
  50505=>"101010100",
  50506=>"110111111",
  50507=>"010111100",
  50508=>"001101000",
  50509=>"001100001",
  50510=>"111101110",
  50511=>"111101001",
  50512=>"110010101",
  50513=>"001100110",
  50514=>"010110000",
  50515=>"010110011",
  50516=>"111100110",
  50517=>"100010010",
  50518=>"111001100",
  50519=>"000110110",
  50520=>"000111101",
  50521=>"000000011",
  50522=>"111011100",
  50523=>"110000110",
  50524=>"110001110",
  50525=>"111111100",
  50526=>"010100110",
  50527=>"110000010",
  50528=>"111000000",
  50529=>"111111010",
  50530=>"000000000",
  50531=>"100101110",
  50532=>"000100010",
  50533=>"101101011",
  50534=>"000110111",
  50535=>"101110101",
  50536=>"101111101",
  50537=>"110111110",
  50538=>"100000010",
  50539=>"111001101",
  50540=>"101111111",
  50541=>"001100110",
  50542=>"010011110",
  50543=>"011101110",
  50544=>"010100111",
  50545=>"110011011",
  50546=>"011000101",
  50547=>"011100101",
  50548=>"001100101",
  50549=>"001110010",
  50550=>"101011011",
  50551=>"000100010",
  50552=>"000000111",
  50553=>"101100001",
  50554=>"011011011",
  50555=>"000101011",
  50556=>"111000101",
  50557=>"110111011",
  50558=>"101101000",
  50559=>"011000010",
  50560=>"111010011",
  50561=>"100011110",
  50562=>"001011010",
  50563=>"001101000",
  50564=>"001000011",
  50565=>"010000011",
  50566=>"111000010",
  50567=>"100001000",
  50568=>"010101011",
  50569=>"111111001",
  50570=>"001111000",
  50571=>"101001011",
  50572=>"000111000",
  50573=>"101110000",
  50574=>"001001001",
  50575=>"110101010",
  50576=>"100100010",
  50577=>"000111011",
  50578=>"111001101",
  50579=>"101111111",
  50580=>"001000111",
  50581=>"011000111",
  50582=>"010011100",
  50583=>"000000110",
  50584=>"100111000",
  50585=>"001110010",
  50586=>"100011010",
  50587=>"111000001",
  50588=>"110000111",
  50589=>"001000100",
  50590=>"111111110",
  50591=>"101100010",
  50592=>"000010010",
  50593=>"011001000",
  50594=>"101000101",
  50595=>"000101110",
  50596=>"010011000",
  50597=>"100001111",
  50598=>"001000010",
  50599=>"010110100",
  50600=>"001100001",
  50601=>"101100101",
  50602=>"111000010",
  50603=>"010000010",
  50604=>"001011110",
  50605=>"110100000",
  50606=>"101100100",
  50607=>"000100010",
  50608=>"000101110",
  50609=>"000110010",
  50610=>"001111001",
  50611=>"101001011",
  50612=>"011011001",
  50613=>"111010110",
  50614=>"101101001",
  50615=>"010010111",
  50616=>"000001011",
  50617=>"010000101",
  50618=>"101011110",
  50619=>"110100111",
  50620=>"010010100",
  50621=>"001100111",
  50622=>"000101101",
  50623=>"100000010",
  50624=>"010001111",
  50625=>"110000110",
  50626=>"100000001",
  50627=>"101110010",
  50628=>"010111001",
  50629=>"101010001",
  50630=>"010001110",
  50631=>"100100101",
  50632=>"100110000",
  50633=>"000110000",
  50634=>"010110011",
  50635=>"101001011",
  50636=>"111000101",
  50637=>"000111100",
  50638=>"111100010",
  50639=>"100100000",
  50640=>"011000110",
  50641=>"011111111",
  50642=>"000011011",
  50643=>"011000000",
  50644=>"010011010",
  50645=>"100100000",
  50646=>"001110100",
  50647=>"001000110",
  50648=>"110111001",
  50649=>"101110111",
  50650=>"001101111",
  50651=>"011101000",
  50652=>"111011110",
  50653=>"101100001",
  50654=>"010100010",
  50655=>"111000000",
  50656=>"001001000",
  50657=>"010000110",
  50658=>"101101000",
  50659=>"111101110",
  50660=>"111011001",
  50661=>"001001010",
  50662=>"111010110",
  50663=>"001100100",
  50664=>"011001101",
  50665=>"110111010",
  50666=>"001010110",
  50667=>"000000110",
  50668=>"001110110",
  50669=>"101100100",
  50670=>"101001100",
  50671=>"011111011",
  50672=>"101101101",
  50673=>"110110010",
  50674=>"011100011",
  50675=>"001001101",
  50676=>"110011111",
  50677=>"110010100",
  50678=>"110100011",
  50679=>"011000010",
  50680=>"000000111",
  50681=>"001011001",
  50682=>"110010110",
  50683=>"001001110",
  50684=>"011011101",
  50685=>"011000010",
  50686=>"010000101",
  50687=>"101011111",
  50688=>"011101110",
  50689=>"010011101",
  50690=>"000101100",
  50691=>"010101010",
  50692=>"010011111",
  50693=>"111010110",
  50694=>"000111101",
  50695=>"111110111",
  50696=>"101110000",
  50697=>"111100111",
  50698=>"110101101",
  50699=>"100011001",
  50700=>"111001000",
  50701=>"011001000",
  50702=>"010100010",
  50703=>"100010011",
  50704=>"110101110",
  50705=>"011100111",
  50706=>"000000100",
  50707=>"010010010",
  50708=>"000101000",
  50709=>"001100010",
  50710=>"000010000",
  50711=>"011110110",
  50712=>"101110111",
  50713=>"110011100",
  50714=>"000011001",
  50715=>"101101111",
  50716=>"100000011",
  50717=>"000011101",
  50718=>"110101011",
  50719=>"010101010",
  50720=>"001000001",
  50721=>"100001011",
  50722=>"101100111",
  50723=>"110000000",
  50724=>"001000010",
  50725=>"111110000",
  50726=>"000110100",
  50727=>"100000110",
  50728=>"110011001",
  50729=>"010010100",
  50730=>"100110011",
  50731=>"110010010",
  50732=>"011100011",
  50733=>"000110110",
  50734=>"010001111",
  50735=>"111110011",
  50736=>"101111111",
  50737=>"110100001",
  50738=>"100100011",
  50739=>"111001010",
  50740=>"100100010",
  50741=>"111010000",
  50742=>"110000001",
  50743=>"010111101",
  50744=>"000010000",
  50745=>"111100111",
  50746=>"101010101",
  50747=>"110001110",
  50748=>"001010110",
  50749=>"101011110",
  50750=>"000100110",
  50751=>"000000110",
  50752=>"111011001",
  50753=>"001000011",
  50754=>"010100101",
  50755=>"010011101",
  50756=>"111110000",
  50757=>"100111010",
  50758=>"100000100",
  50759=>"000010001",
  50760=>"000010010",
  50761=>"011001010",
  50762=>"100011100",
  50763=>"101101111",
  50764=>"011011000",
  50765=>"101000110",
  50766=>"010110000",
  50767=>"101101010",
  50768=>"011010111",
  50769=>"101111000",
  50770=>"000100101",
  50771=>"010110011",
  50772=>"000001100",
  50773=>"110111001",
  50774=>"100001100",
  50775=>"101111011",
  50776=>"100101100",
  50777=>"011001010",
  50778=>"100001010",
  50779=>"111010101",
  50780=>"100001100",
  50781=>"101100100",
  50782=>"111100101",
  50783=>"000110110",
  50784=>"111100000",
  50785=>"001111011",
  50786=>"001001100",
  50787=>"100000011",
  50788=>"010110110",
  50789=>"011100011",
  50790=>"000000001",
  50791=>"111010010",
  50792=>"101010101",
  50793=>"100111100",
  50794=>"011100010",
  50795=>"100100000",
  50796=>"101101011",
  50797=>"111110011",
  50798=>"111000000",
  50799=>"111101010",
  50800=>"111110010",
  50801=>"000010111",
  50802=>"111010100",
  50803=>"100100111",
  50804=>"001011010",
  50805=>"110110011",
  50806=>"011110110",
  50807=>"000010100",
  50808=>"010111101",
  50809=>"001101100",
  50810=>"101001100",
  50811=>"001011111",
  50812=>"001101000",
  50813=>"110010011",
  50814=>"111111110",
  50815=>"101000000",
  50816=>"010010111",
  50817=>"011000100",
  50818=>"010101010",
  50819=>"000110111",
  50820=>"110100110",
  50821=>"001110101",
  50822=>"000001110",
  50823=>"000001010",
  50824=>"001111010",
  50825=>"000110110",
  50826=>"100111001",
  50827=>"011010111",
  50828=>"100000101",
  50829=>"111000001",
  50830=>"001101110",
  50831=>"100001111",
  50832=>"101001000",
  50833=>"011010010",
  50834=>"101101001",
  50835=>"010011001",
  50836=>"010111001",
  50837=>"011100100",
  50838=>"000010000",
  50839=>"100111100",
  50840=>"111111010",
  50841=>"000110010",
  50842=>"111110101",
  50843=>"100111101",
  50844=>"001011100",
  50845=>"000110001",
  50846=>"000010000",
  50847=>"000011100",
  50848=>"010000011",
  50849=>"000000011",
  50850=>"000001000",
  50851=>"110100000",
  50852=>"010010101",
  50853=>"110010011",
  50854=>"101101000",
  50855=>"000110000",
  50856=>"111010111",
  50857=>"011110110",
  50858=>"110101101",
  50859=>"000010100",
  50860=>"111100111",
  50861=>"110010000",
  50862=>"111111000",
  50863=>"110010000",
  50864=>"100101011",
  50865=>"010110001",
  50866=>"111001000",
  50867=>"111101100",
  50868=>"101010101",
  50869=>"110001111",
  50870=>"011110001",
  50871=>"001010001",
  50872=>"010011010",
  50873=>"011000001",
  50874=>"110110100",
  50875=>"110110111",
  50876=>"111101011",
  50877=>"101111111",
  50878=>"000001110",
  50879=>"111111110",
  50880=>"110100110",
  50881=>"011110100",
  50882=>"010110111",
  50883=>"010111101",
  50884=>"101011101",
  50885=>"001001100",
  50886=>"100110101",
  50887=>"000000011",
  50888=>"001100010",
  50889=>"111000001",
  50890=>"100111100",
  50891=>"001110111",
  50892=>"101011010",
  50893=>"001001000",
  50894=>"001001000",
  50895=>"100100110",
  50896=>"010001010",
  50897=>"100011011",
  50898=>"100000111",
  50899=>"100110101",
  50900=>"101110000",
  50901=>"001100110",
  50902=>"001100110",
  50903=>"010100010",
  50904=>"100111111",
  50905=>"100001101",
  50906=>"001000101",
  50907=>"110101000",
  50908=>"101011011",
  50909=>"110100111",
  50910=>"101111011",
  50911=>"110110010",
  50912=>"100111110",
  50913=>"001100110",
  50914=>"011000000",
  50915=>"100100111",
  50916=>"111011111",
  50917=>"001011000",
  50918=>"111000000",
  50919=>"000010110",
  50920=>"110101000",
  50921=>"111010100",
  50922=>"011111011",
  50923=>"000000110",
  50924=>"011110011",
  50925=>"000101100",
  50926=>"000011100",
  50927=>"010010000",
  50928=>"111000111",
  50929=>"011001000",
  50930=>"000000010",
  50931=>"110100110",
  50932=>"110001001",
  50933=>"010110001",
  50934=>"000010011",
  50935=>"101110000",
  50936=>"111110001",
  50937=>"100001111",
  50938=>"100010010",
  50939=>"000111111",
  50940=>"001011110",
  50941=>"001101011",
  50942=>"011101001",
  50943=>"010000010",
  50944=>"111011101",
  50945=>"000111110",
  50946=>"011110001",
  50947=>"111111110",
  50948=>"000101100",
  50949=>"110101100",
  50950=>"000100001",
  50951=>"000000110",
  50952=>"111000001",
  50953=>"011111011",
  50954=>"010100100",
  50955=>"000010000",
  50956=>"011110100",
  50957=>"000000000",
  50958=>"111111011",
  50959=>"001110100",
  50960=>"001100010",
  50961=>"101101001",
  50962=>"010101110",
  50963=>"011011010",
  50964=>"000110101",
  50965=>"111001111",
  50966=>"001010000",
  50967=>"101011011",
  50968=>"111001001",
  50969=>"111000111",
  50970=>"010011000",
  50971=>"111110110",
  50972=>"011001010",
  50973=>"111111101",
  50974=>"101110101",
  50975=>"011101000",
  50976=>"111100100",
  50977=>"001010111",
  50978=>"100101100",
  50979=>"101100111",
  50980=>"010001100",
  50981=>"111110101",
  50982=>"110110010",
  50983=>"000011011",
  50984=>"110010101",
  50985=>"010010001",
  50986=>"111110011",
  50987=>"101101000",
  50988=>"011010011",
  50989=>"000000000",
  50990=>"010111111",
  50991=>"010111010",
  50992=>"001011000",
  50993=>"001000101",
  50994=>"010011111",
  50995=>"010100000",
  50996=>"010110000",
  50997=>"111101101",
  50998=>"111011100",
  50999=>"111111011",
  51000=>"001111011",
  51001=>"100100100",
  51002=>"011110011",
  51003=>"111100011",
  51004=>"100101110",
  51005=>"100010000",
  51006=>"111001010",
  51007=>"001000100",
  51008=>"011110001",
  51009=>"110111111",
  51010=>"000001100",
  51011=>"110100110",
  51012=>"110101011",
  51013=>"100011101",
  51014=>"111101110",
  51015=>"101101000",
  51016=>"101000010",
  51017=>"101111100",
  51018=>"011001000",
  51019=>"000000011",
  51020=>"100110001",
  51021=>"010011000",
  51022=>"111110011",
  51023=>"101011000",
  51024=>"110100100",
  51025=>"110000011",
  51026=>"011001101",
  51027=>"010110010",
  51028=>"001100011",
  51029=>"011011101",
  51030=>"100110101",
  51031=>"100001000",
  51032=>"001000010",
  51033=>"110011100",
  51034=>"000001000",
  51035=>"110000100",
  51036=>"011001100",
  51037=>"111101011",
  51038=>"110011010",
  51039=>"111101111",
  51040=>"001111011",
  51041=>"001001001",
  51042=>"101100111",
  51043=>"101111010",
  51044=>"100101101",
  51045=>"000001100",
  51046=>"001100100",
  51047=>"011001101",
  51048=>"001111001",
  51049=>"101001001",
  51050=>"000101000",
  51051=>"101100001",
  51052=>"001101010",
  51053=>"001101001",
  51054=>"000101111",
  51055=>"110101011",
  51056=>"000100001",
  51057=>"100101101",
  51058=>"110001110",
  51059=>"101111101",
  51060=>"010011101",
  51061=>"000111010",
  51062=>"100001110",
  51063=>"110101100",
  51064=>"010101101",
  51065=>"101000101",
  51066=>"010110100",
  51067=>"010110010",
  51068=>"110111111",
  51069=>"101001101",
  51070=>"011000100",
  51071=>"011001110",
  51072=>"000000001",
  51073=>"111001110",
  51074=>"011110100",
  51075=>"010001111",
  51076=>"011010011",
  51077=>"111000110",
  51078=>"100110011",
  51079=>"110001000",
  51080=>"111110111",
  51081=>"111001111",
  51082=>"101011001",
  51083=>"100101101",
  51084=>"110101011",
  51085=>"011100001",
  51086=>"111000001",
  51087=>"010111100",
  51088=>"100101100",
  51089=>"111100001",
  51090=>"111111001",
  51091=>"001110011",
  51092=>"011000110",
  51093=>"100111110",
  51094=>"010100100",
  51095=>"100001000",
  51096=>"111110001",
  51097=>"000000101",
  51098=>"011011001",
  51099=>"010000001",
  51100=>"000100001",
  51101=>"110010101",
  51102=>"010011100",
  51103=>"100101000",
  51104=>"101100000",
  51105=>"000010100",
  51106=>"100111011",
  51107=>"101010001",
  51108=>"000110100",
  51109=>"110000000",
  51110=>"001100110",
  51111=>"010001010",
  51112=>"000010000",
  51113=>"010011010",
  51114=>"001110101",
  51115=>"100110000",
  51116=>"101000000",
  51117=>"111000110",
  51118=>"010101000",
  51119=>"011001110",
  51120=>"011000100",
  51121=>"001000001",
  51122=>"101000100",
  51123=>"110111010",
  51124=>"011101111",
  51125=>"011110100",
  51126=>"110000001",
  51127=>"101011101",
  51128=>"100000000",
  51129=>"010010110",
  51130=>"100101100",
  51131=>"111101010",
  51132=>"110110101",
  51133=>"001001101",
  51134=>"011110001",
  51135=>"001010000",
  51136=>"101001110",
  51137=>"010000000",
  51138=>"111111010",
  51139=>"110100011",
  51140=>"111010000",
  51141=>"100011100",
  51142=>"011001100",
  51143=>"101010100",
  51144=>"110000100",
  51145=>"010110000",
  51146=>"110111101",
  51147=>"111000010",
  51148=>"000000000",
  51149=>"010100010",
  51150=>"111110011",
  51151=>"110010101",
  51152=>"101110001",
  51153=>"100000011",
  51154=>"001111010",
  51155=>"110001000",
  51156=>"111111111",
  51157=>"011000101",
  51158=>"001010100",
  51159=>"001101110",
  51160=>"101111110",
  51161=>"110111001",
  51162=>"011100111",
  51163=>"000000000",
  51164=>"010001111",
  51165=>"100111010",
  51166=>"111000000",
  51167=>"001000111",
  51168=>"111111110",
  51169=>"101110101",
  51170=>"000110101",
  51171=>"000000111",
  51172=>"011001101",
  51173=>"001000000",
  51174=>"110011111",
  51175=>"010110011",
  51176=>"000010111",
  51177=>"001010100",
  51178=>"011011110",
  51179=>"101001000",
  51180=>"111111111",
  51181=>"100011101",
  51182=>"010110011",
  51183=>"000111000",
  51184=>"111101110",
  51185=>"101111110",
  51186=>"000000000",
  51187=>"100000111",
  51188=>"110111101",
  51189=>"000001010",
  51190=>"000100000",
  51191=>"000011010",
  51192=>"111101000",
  51193=>"101111101",
  51194=>"110010010",
  51195=>"111010111",
  51196=>"111100101",
  51197=>"010011110",
  51198=>"110010101",
  51199=>"001010011",
  51200=>"001010100",
  51201=>"010100100",
  51202=>"100010010",
  51203=>"010000100",
  51204=>"010001100",
  51205=>"101111000",
  51206=>"101001001",
  51207=>"000110000",
  51208=>"101101001",
  51209=>"000101111",
  51210=>"100101101",
  51211=>"000010110",
  51212=>"101000100",
  51213=>"111110000",
  51214=>"000101100",
  51215=>"000100011",
  51216=>"001011100",
  51217=>"000011101",
  51218=>"000110101",
  51219=>"100010001",
  51220=>"000101110",
  51221=>"000101000",
  51222=>"000011000",
  51223=>"111101001",
  51224=>"110110011",
  51225=>"010000100",
  51226=>"101010000",
  51227=>"111101001",
  51228=>"110010101",
  51229=>"101110101",
  51230=>"000111111",
  51231=>"110001100",
  51232=>"001011011",
  51233=>"101111001",
  51234=>"000110100",
  51235=>"111011000",
  51236=>"011101010",
  51237=>"000100000",
  51238=>"000100100",
  51239=>"111001110",
  51240=>"110011011",
  51241=>"010101001",
  51242=>"111000001",
  51243=>"101110011",
  51244=>"101010101",
  51245=>"110001110",
  51246=>"001001001",
  51247=>"001001100",
  51248=>"011000001",
  51249=>"000010010",
  51250=>"001000101",
  51251=>"011101101",
  51252=>"010110100",
  51253=>"010100100",
  51254=>"111100001",
  51255=>"001001000",
  51256=>"001100101",
  51257=>"101111001",
  51258=>"100100101",
  51259=>"001111000",
  51260=>"111001101",
  51261=>"110000100",
  51262=>"011010101",
  51263=>"100000101",
  51264=>"101110000",
  51265=>"000100000",
  51266=>"100100101",
  51267=>"001100111",
  51268=>"010000001",
  51269=>"111111001",
  51270=>"100001101",
  51271=>"110101001",
  51272=>"001001100",
  51273=>"000011111",
  51274=>"010111011",
  51275=>"110101001",
  51276=>"000001111",
  51277=>"111110110",
  51278=>"011000001",
  51279=>"100100110",
  51280=>"110011101",
  51281=>"110011001",
  51282=>"101001110",
  51283=>"010000011",
  51284=>"101010100",
  51285=>"100011001",
  51286=>"010010111",
  51287=>"010111100",
  51288=>"000011110",
  51289=>"000000111",
  51290=>"110010110",
  51291=>"000001110",
  51292=>"000110011",
  51293=>"000010101",
  51294=>"010111011",
  51295=>"001110111",
  51296=>"110001001",
  51297=>"100000000",
  51298=>"101110000",
  51299=>"011000001",
  51300=>"010100101",
  51301=>"101010011",
  51302=>"011001011",
  51303=>"000001000",
  51304=>"100011000",
  51305=>"000000110",
  51306=>"111101100",
  51307=>"110101111",
  51308=>"110011011",
  51309=>"011111101",
  51310=>"111100001",
  51311=>"110011100",
  51312=>"000100011",
  51313=>"101101000",
  51314=>"011110010",
  51315=>"110001111",
  51316=>"011110101",
  51317=>"111101100",
  51318=>"000011101",
  51319=>"000100001",
  51320=>"100011010",
  51321=>"100100110",
  51322=>"101111000",
  51323=>"110100000",
  51324=>"010000001",
  51325=>"000001011",
  51326=>"110101110",
  51327=>"011110111",
  51328=>"000000001",
  51329=>"001001001",
  51330=>"101000110",
  51331=>"000010011",
  51332=>"101010010",
  51333=>"101111001",
  51334=>"111000000",
  51335=>"001100111",
  51336=>"111111111",
  51337=>"001001101",
  51338=>"000010011",
  51339=>"000011111",
  51340=>"110110000",
  51341=>"100101110",
  51342=>"011110101",
  51343=>"101010000",
  51344=>"010110001",
  51345=>"101001001",
  51346=>"001011101",
  51347=>"011000010",
  51348=>"010100111",
  51349=>"010110110",
  51350=>"010010010",
  51351=>"101111000",
  51352=>"010000111",
  51353=>"111000100",
  51354=>"110110101",
  51355=>"011001111",
  51356=>"101100101",
  51357=>"001111110",
  51358=>"000101110",
  51359=>"101000101",
  51360=>"011101111",
  51361=>"000000101",
  51362=>"010100101",
  51363=>"101001011",
  51364=>"000101011",
  51365=>"100111101",
  51366=>"110010010",
  51367=>"000001101",
  51368=>"011001010",
  51369=>"011101010",
  51370=>"001001110",
  51371=>"000011111",
  51372=>"001100001",
  51373=>"101101111",
  51374=>"110010100",
  51375=>"010000010",
  51376=>"000011011",
  51377=>"011100100",
  51378=>"010001100",
  51379=>"101011101",
  51380=>"001000110",
  51381=>"011010000",
  51382=>"011000011",
  51383=>"000101011",
  51384=>"001100110",
  51385=>"000110111",
  51386=>"101110110",
  51387=>"100000001",
  51388=>"101101101",
  51389=>"011000001",
  51390=>"010100110",
  51391=>"011001110",
  51392=>"111010001",
  51393=>"011001110",
  51394=>"011000111",
  51395=>"110100011",
  51396=>"000011001",
  51397=>"111001110",
  51398=>"001100111",
  51399=>"001110111",
  51400=>"101011010",
  51401=>"111110100",
  51402=>"010111110",
  51403=>"010100100",
  51404=>"110101101",
  51405=>"010111110",
  51406=>"011110010",
  51407=>"101000001",
  51408=>"111001100",
  51409=>"000110011",
  51410=>"000000010",
  51411=>"001110111",
  51412=>"010111011",
  51413=>"011011100",
  51414=>"100000100",
  51415=>"100001001",
  51416=>"101000010",
  51417=>"111111000",
  51418=>"110000001",
  51419=>"111110001",
  51420=>"001001000",
  51421=>"000110111",
  51422=>"110010001",
  51423=>"001000110",
  51424=>"010101010",
  51425=>"111011001",
  51426=>"000010010",
  51427=>"010000000",
  51428=>"100011010",
  51429=>"100111110",
  51430=>"100001000",
  51431=>"000100100",
  51432=>"101000101",
  51433=>"011111101",
  51434=>"100010000",
  51435=>"101111101",
  51436=>"010101011",
  51437=>"111110010",
  51438=>"000111110",
  51439=>"010000000",
  51440=>"100000001",
  51441=>"000011110",
  51442=>"110111101",
  51443=>"110000110",
  51444=>"110100010",
  51445=>"101010010",
  51446=>"100110101",
  51447=>"010010100",
  51448=>"101110011",
  51449=>"000001111",
  51450=>"011111100",
  51451=>"100011101",
  51452=>"011011111",
  51453=>"011010010",
  51454=>"100001101",
  51455=>"101000001",
  51456=>"111101000",
  51457=>"100101001",
  51458=>"001111100",
  51459=>"000100110",
  51460=>"000101001",
  51461=>"011111111",
  51462=>"001001001",
  51463=>"101100000",
  51464=>"011111111",
  51465=>"001110010",
  51466=>"111101101",
  51467=>"000101001",
  51468=>"010010101",
  51469=>"101000100",
  51470=>"011011010",
  51471=>"010010000",
  51472=>"001111110",
  51473=>"110010110",
  51474=>"000110010",
  51475=>"111101001",
  51476=>"011000001",
  51477=>"111100011",
  51478=>"101111011",
  51479=>"111000100",
  51480=>"100100011",
  51481=>"011001111",
  51482=>"001111111",
  51483=>"111010100",
  51484=>"011100011",
  51485=>"000101000",
  51486=>"100001011",
  51487=>"001000001",
  51488=>"100110101",
  51489=>"100101001",
  51490=>"010110001",
  51491=>"111011010",
  51492=>"110000100",
  51493=>"110011001",
  51494=>"010011110",
  51495=>"100111000",
  51496=>"100011111",
  51497=>"110011010",
  51498=>"100001010",
  51499=>"010000101",
  51500=>"111101111",
  51501=>"000101011",
  51502=>"000000010",
  51503=>"110111010",
  51504=>"100110111",
  51505=>"110010111",
  51506=>"001011100",
  51507=>"010000101",
  51508=>"110000111",
  51509=>"001111101",
  51510=>"010101110",
  51511=>"010010100",
  51512=>"010001111",
  51513=>"110111110",
  51514=>"110111111",
  51515=>"111011110",
  51516=>"011011000",
  51517=>"000111101",
  51518=>"110110111",
  51519=>"111101110",
  51520=>"010001100",
  51521=>"111011110",
  51522=>"100011100",
  51523=>"011111001",
  51524=>"101011000",
  51525=>"010100111",
  51526=>"110100000",
  51527=>"100000010",
  51528=>"101000011",
  51529=>"000001011",
  51530=>"100101000",
  51531=>"100000100",
  51532=>"001110110",
  51533=>"100010101",
  51534=>"110001011",
  51535=>"111010101",
  51536=>"011000010",
  51537=>"011110101",
  51538=>"010000101",
  51539=>"101101110",
  51540=>"100110111",
  51541=>"100111010",
  51542=>"011110100",
  51543=>"110011000",
  51544=>"011110100",
  51545=>"000001000",
  51546=>"001111110",
  51547=>"001111000",
  51548=>"110100101",
  51549=>"111011001",
  51550=>"101101001",
  51551=>"111101101",
  51552=>"000111101",
  51553=>"001001110",
  51554=>"110001000",
  51555=>"100111100",
  51556=>"010000101",
  51557=>"110011111",
  51558=>"101110001",
  51559=>"100011111",
  51560=>"110110111",
  51561=>"001111111",
  51562=>"000010001",
  51563=>"000000010",
  51564=>"000011111",
  51565=>"111011010",
  51566=>"010001100",
  51567=>"001110010",
  51568=>"101010110",
  51569=>"000100010",
  51570=>"000011100",
  51571=>"110101110",
  51572=>"110000001",
  51573=>"011001010",
  51574=>"101010001",
  51575=>"000000100",
  51576=>"001000000",
  51577=>"001011101",
  51578=>"010110000",
  51579=>"000101000",
  51580=>"111101111",
  51581=>"000011111",
  51582=>"001111010",
  51583=>"110010111",
  51584=>"100011000",
  51585=>"010110001",
  51586=>"001001100",
  51587=>"111111101",
  51588=>"011100111",
  51589=>"011010100",
  51590=>"010110001",
  51591=>"110101001",
  51592=>"011000000",
  51593=>"010001111",
  51594=>"111111100",
  51595=>"100011011",
  51596=>"110010100",
  51597=>"011101010",
  51598=>"010001000",
  51599=>"001010001",
  51600=>"111101111",
  51601=>"000110000",
  51602=>"101110011",
  51603=>"000011000",
  51604=>"101110000",
  51605=>"010000000",
  51606=>"001010011",
  51607=>"000011000",
  51608=>"001110101",
  51609=>"001110111",
  51610=>"101101100",
  51611=>"001010011",
  51612=>"100011011",
  51613=>"001111000",
  51614=>"010100001",
  51615=>"111000101",
  51616=>"011011111",
  51617=>"110110010",
  51618=>"001010100",
  51619=>"110101000",
  51620=>"001111000",
  51621=>"000110111",
  51622=>"001000111",
  51623=>"111100111",
  51624=>"100111110",
  51625=>"010110110",
  51626=>"100100110",
  51627=>"010010011",
  51628=>"101110100",
  51629=>"010111001",
  51630=>"011100100",
  51631=>"000101111",
  51632=>"010000101",
  51633=>"100110100",
  51634=>"010101101",
  51635=>"111011001",
  51636=>"001010001",
  51637=>"111101011",
  51638=>"101111110",
  51639=>"010100100",
  51640=>"111011001",
  51641=>"100100110",
  51642=>"001101000",
  51643=>"110010111",
  51644=>"111111101",
  51645=>"011100111",
  51646=>"100111101",
  51647=>"100010101",
  51648=>"000010000",
  51649=>"000101111",
  51650=>"110011100",
  51651=>"011000000",
  51652=>"111111110",
  51653=>"101001110",
  51654=>"110010101",
  51655=>"010000000",
  51656=>"100101010",
  51657=>"111101001",
  51658=>"001010000",
  51659=>"101011010",
  51660=>"101010011",
  51661=>"110000010",
  51662=>"100000000",
  51663=>"011010011",
  51664=>"110000111",
  51665=>"000010011",
  51666=>"100011110",
  51667=>"100111100",
  51668=>"010110110",
  51669=>"000101000",
  51670=>"100000001",
  51671=>"001001110",
  51672=>"001010110",
  51673=>"001010100",
  51674=>"110110101",
  51675=>"000100011",
  51676=>"111101111",
  51677=>"000101011",
  51678=>"100000100",
  51679=>"110111001",
  51680=>"010101001",
  51681=>"111101110",
  51682=>"111001010",
  51683=>"101100101",
  51684=>"100101010",
  51685=>"101010100",
  51686=>"001010111",
  51687=>"001110101",
  51688=>"110101000",
  51689=>"101111000",
  51690=>"001100100",
  51691=>"101000101",
  51692=>"010110001",
  51693=>"110010010",
  51694=>"101001010",
  51695=>"111011011",
  51696=>"100101111",
  51697=>"101001100",
  51698=>"001110100",
  51699=>"101100010",
  51700=>"101101011",
  51701=>"100011000",
  51702=>"100101010",
  51703=>"111110011",
  51704=>"010000000",
  51705=>"100011011",
  51706=>"001011011",
  51707=>"110010000",
  51708=>"100001101",
  51709=>"010111111",
  51710=>"011101100",
  51711=>"110011000",
  51712=>"100001111",
  51713=>"001110001",
  51714=>"100010101",
  51715=>"010100110",
  51716=>"110001000",
  51717=>"101101111",
  51718=>"100011100",
  51719=>"000101111",
  51720=>"100000011",
  51721=>"000101011",
  51722=>"110011001",
  51723=>"111100110",
  51724=>"011110011",
  51725=>"011110111",
  51726=>"111111100",
  51727=>"101011101",
  51728=>"110010111",
  51729=>"111101110",
  51730=>"001011010",
  51731=>"111001110",
  51732=>"001000110",
  51733=>"000000000",
  51734=>"011011000",
  51735=>"101000000",
  51736=>"000001010",
  51737=>"011010000",
  51738=>"000100011",
  51739=>"011101000",
  51740=>"111001111",
  51741=>"111100111",
  51742=>"000100101",
  51743=>"100011010",
  51744=>"100010000",
  51745=>"000010111",
  51746=>"010101001",
  51747=>"101000011",
  51748=>"111011110",
  51749=>"010100111",
  51750=>"010011111",
  51751=>"001111000",
  51752=>"010011001",
  51753=>"001111001",
  51754=>"111111110",
  51755=>"001000010",
  51756=>"011011111",
  51757=>"111111011",
  51758=>"011101110",
  51759=>"110101101",
  51760=>"000010111",
  51761=>"101000100",
  51762=>"110010000",
  51763=>"010100100",
  51764=>"000010111",
  51765=>"110001100",
  51766=>"011101111",
  51767=>"011111111",
  51768=>"111110101",
  51769=>"100100010",
  51770=>"111010100",
  51771=>"101010011",
  51772=>"101011110",
  51773=>"111000000",
  51774=>"001000010",
  51775=>"001000010",
  51776=>"101111000",
  51777=>"111110000",
  51778=>"100010101",
  51779=>"001001010",
  51780=>"100100000",
  51781=>"111101000",
  51782=>"000001110",
  51783=>"010010101",
  51784=>"011100000",
  51785=>"001011000",
  51786=>"101111011",
  51787=>"010101110",
  51788=>"001100010",
  51789=>"110010100",
  51790=>"100011111",
  51791=>"001101111",
  51792=>"110110111",
  51793=>"010101110",
  51794=>"101001001",
  51795=>"111001000",
  51796=>"000010111",
  51797=>"000101010",
  51798=>"010010000",
  51799=>"101011111",
  51800=>"101111111",
  51801=>"011101110",
  51802=>"010101010",
  51803=>"000100001",
  51804=>"110100011",
  51805=>"000001010",
  51806=>"100111000",
  51807=>"000010100",
  51808=>"010100101",
  51809=>"001111110",
  51810=>"010101010",
  51811=>"000101000",
  51812=>"011001001",
  51813=>"011111101",
  51814=>"011100011",
  51815=>"110111110",
  51816=>"110010001",
  51817=>"101110100",
  51818=>"100110011",
  51819=>"110010001",
  51820=>"000000101",
  51821=>"111010010",
  51822=>"111001010",
  51823=>"000010111",
  51824=>"101000000",
  51825=>"101010011",
  51826=>"001101110",
  51827=>"000101100",
  51828=>"010000111",
  51829=>"000001010",
  51830=>"111010110",
  51831=>"100000000",
  51832=>"101010010",
  51833=>"110110000",
  51834=>"101010100",
  51835=>"101110101",
  51836=>"101001010",
  51837=>"101011111",
  51838=>"101011111",
  51839=>"010100010",
  51840=>"100111100",
  51841=>"111110111",
  51842=>"011010010",
  51843=>"101001010",
  51844=>"000110010",
  51845=>"000001111",
  51846=>"110011111",
  51847=>"000011100",
  51848=>"010000111",
  51849=>"011101000",
  51850=>"010110001",
  51851=>"110001000",
  51852=>"011011100",
  51853=>"010110111",
  51854=>"111111111",
  51855=>"010101000",
  51856=>"001011100",
  51857=>"100100011",
  51858=>"100110100",
  51859=>"011111100",
  51860=>"001111101",
  51861=>"100101001",
  51862=>"001111001",
  51863=>"100010101",
  51864=>"100001011",
  51865=>"110000011",
  51866=>"000110100",
  51867=>"110100110",
  51868=>"011011001",
  51869=>"001011101",
  51870=>"010011111",
  51871=>"000110000",
  51872=>"110001000",
  51873=>"000000000",
  51874=>"011110110",
  51875=>"010111100",
  51876=>"111001101",
  51877=>"010110000",
  51878=>"101001000",
  51879=>"001011111",
  51880=>"100011111",
  51881=>"101100001",
  51882=>"111011001",
  51883=>"100111110",
  51884=>"101010000",
  51885=>"011011100",
  51886=>"101101100",
  51887=>"000011001",
  51888=>"100011011",
  51889=>"110111101",
  51890=>"010100111",
  51891=>"000100110",
  51892=>"111101111",
  51893=>"011111110",
  51894=>"000100111",
  51895=>"010011001",
  51896=>"011010010",
  51897=>"111011011",
  51898=>"111101100",
  51899=>"100110101",
  51900=>"001000000",
  51901=>"100010110",
  51902=>"001001111",
  51903=>"110111011",
  51904=>"100001001",
  51905=>"000110011",
  51906=>"000111000",
  51907=>"000111001",
  51908=>"110101010",
  51909=>"110010110",
  51910=>"110001110",
  51911=>"101110100",
  51912=>"000001111",
  51913=>"101110011",
  51914=>"101001111",
  51915=>"001010101",
  51916=>"010010110",
  51917=>"010001101",
  51918=>"101100010",
  51919=>"100000010",
  51920=>"101111001",
  51921=>"000000101",
  51922=>"111100011",
  51923=>"101101110",
  51924=>"001010110",
  51925=>"010011010",
  51926=>"100111011",
  51927=>"101011000",
  51928=>"110010011",
  51929=>"011100100",
  51930=>"000001111",
  51931=>"011100010",
  51932=>"011100011",
  51933=>"111001000",
  51934=>"011101010",
  51935=>"011111110",
  51936=>"001010010",
  51937=>"001000011",
  51938=>"100010010",
  51939=>"100100111",
  51940=>"011100001",
  51941=>"110111011",
  51942=>"110110110",
  51943=>"011010000",
  51944=>"001110110",
  51945=>"001111111",
  51946=>"111011110",
  51947=>"111011010",
  51948=>"101101011",
  51949=>"010011100",
  51950=>"110011111",
  51951=>"101111100",
  51952=>"100011100",
  51953=>"110110011",
  51954=>"111001010",
  51955=>"110001011",
  51956=>"111101111",
  51957=>"100011111",
  51958=>"111100000",
  51959=>"110111101",
  51960=>"010010100",
  51961=>"011000100",
  51962=>"001000011",
  51963=>"000001011",
  51964=>"011111010",
  51965=>"111101100",
  51966=>"011100001",
  51967=>"111101111",
  51968=>"101110010",
  51969=>"001011101",
  51970=>"010001101",
  51971=>"100000000",
  51972=>"110010101",
  51973=>"100101100",
  51974=>"110111001",
  51975=>"011101000",
  51976=>"000100111",
  51977=>"110111100",
  51978=>"010111001",
  51979=>"000101011",
  51980=>"111000011",
  51981=>"100101010",
  51982=>"111000100",
  51983=>"110000100",
  51984=>"111111100",
  51985=>"000101000",
  51986=>"100011000",
  51987=>"010100001",
  51988=>"010100100",
  51989=>"111000100",
  51990=>"110101011",
  51991=>"100100010",
  51992=>"011010010",
  51993=>"011000100",
  51994=>"111010110",
  51995=>"011111101",
  51996=>"110001110",
  51997=>"010100001",
  51998=>"000011111",
  51999=>"100001100",
  52000=>"101110111",
  52001=>"110111100",
  52002=>"001000010",
  52003=>"000001101",
  52004=>"011000110",
  52005=>"010100101",
  52006=>"111110010",
  52007=>"010001010",
  52008=>"101111001",
  52009=>"110101001",
  52010=>"111110111",
  52011=>"000011000",
  52012=>"111100111",
  52013=>"001000111",
  52014=>"011111010",
  52015=>"101001010",
  52016=>"001000011",
  52017=>"000001000",
  52018=>"111001101",
  52019=>"100110101",
  52020=>"001011010",
  52021=>"010111010",
  52022=>"000100010",
  52023=>"100110111",
  52024=>"111010011",
  52025=>"111110010",
  52026=>"101100111",
  52027=>"111110010",
  52028=>"000100000",
  52029=>"000010001",
  52030=>"000010011",
  52031=>"010100111",
  52032=>"100000010",
  52033=>"001101011",
  52034=>"010110000",
  52035=>"000010110",
  52036=>"100100001",
  52037=>"100101101",
  52038=>"110000000",
  52039=>"101000011",
  52040=>"101101110",
  52041=>"110110010",
  52042=>"111101111",
  52043=>"001101010",
  52044=>"010111000",
  52045=>"011001000",
  52046=>"101000010",
  52047=>"010010001",
  52048=>"001010001",
  52049=>"100000010",
  52050=>"100111010",
  52051=>"000101001",
  52052=>"111010110",
  52053=>"001111100",
  52054=>"011010100",
  52055=>"011000110",
  52056=>"100010011",
  52057=>"010011001",
  52058=>"100110111",
  52059=>"001100111",
  52060=>"111100001",
  52061=>"110111011",
  52062=>"101010001",
  52063=>"000000111",
  52064=>"111111000",
  52065=>"011001100",
  52066=>"101111011",
  52067=>"001101100",
  52068=>"001101011",
  52069=>"011110101",
  52070=>"001011101",
  52071=>"111101100",
  52072=>"011110101",
  52073=>"010000111",
  52074=>"000111100",
  52075=>"000111111",
  52076=>"101101111",
  52077=>"000111110",
  52078=>"101010100",
  52079=>"111010010",
  52080=>"010010000",
  52081=>"001100111",
  52082=>"100010000",
  52083=>"111010010",
  52084=>"101110001",
  52085=>"010010000",
  52086=>"111110111",
  52087=>"001000001",
  52088=>"010010011",
  52089=>"100111111",
  52090=>"100000001",
  52091=>"010000100",
  52092=>"100110100",
  52093=>"010110001",
  52094=>"000011001",
  52095=>"110111000",
  52096=>"111101110",
  52097=>"010110010",
  52098=>"000001000",
  52099=>"000110010",
  52100=>"000110111",
  52101=>"011100101",
  52102=>"011011101",
  52103=>"100101110",
  52104=>"011110011",
  52105=>"001100010",
  52106=>"001100010",
  52107=>"000010000",
  52108=>"011111110",
  52109=>"111010110",
  52110=>"100101011",
  52111=>"110001111",
  52112=>"010010010",
  52113=>"101101011",
  52114=>"000100100",
  52115=>"110101100",
  52116=>"111110110",
  52117=>"100100011",
  52118=>"011001001",
  52119=>"011000000",
  52120=>"100110100",
  52121=>"000110101",
  52122=>"111000000",
  52123=>"111111001",
  52124=>"000111000",
  52125=>"000010110",
  52126=>"011111000",
  52127=>"000111011",
  52128=>"111101001",
  52129=>"100110001",
  52130=>"101101000",
  52131=>"101011111",
  52132=>"010100010",
  52133=>"001101100",
  52134=>"011100110",
  52135=>"011001000",
  52136=>"000010111",
  52137=>"010100011",
  52138=>"110101110",
  52139=>"111101111",
  52140=>"010001001",
  52141=>"111011101",
  52142=>"110100010",
  52143=>"101011010",
  52144=>"011100011",
  52145=>"111001001",
  52146=>"000101110",
  52147=>"000111110",
  52148=>"101010001",
  52149=>"011010110",
  52150=>"110000001",
  52151=>"011001010",
  52152=>"101010100",
  52153=>"001100110",
  52154=>"010010100",
  52155=>"101000011",
  52156=>"001010011",
  52157=>"110010110",
  52158=>"110110111",
  52159=>"001100111",
  52160=>"110010111",
  52161=>"101111110",
  52162=>"010100010",
  52163=>"000001110",
  52164=>"101000010",
  52165=>"111111111",
  52166=>"011110110",
  52167=>"101000010",
  52168=>"000001011",
  52169=>"110110011",
  52170=>"001000000",
  52171=>"001000110",
  52172=>"010010110",
  52173=>"111000000",
  52174=>"111100011",
  52175=>"100010110",
  52176=>"011001011",
  52177=>"110001100",
  52178=>"101001011",
  52179=>"000100010",
  52180=>"000111110",
  52181=>"111111110",
  52182=>"111000101",
  52183=>"101011000",
  52184=>"000011110",
  52185=>"100110110",
  52186=>"110000100",
  52187=>"110100010",
  52188=>"100100110",
  52189=>"100001100",
  52190=>"101010010",
  52191=>"111110100",
  52192=>"100111001",
  52193=>"110111101",
  52194=>"011010010",
  52195=>"100010110",
  52196=>"010010110",
  52197=>"100000011",
  52198=>"110111101",
  52199=>"000100001",
  52200=>"000011101",
  52201=>"000010110",
  52202=>"010011111",
  52203=>"000110000",
  52204=>"101111111",
  52205=>"001001001",
  52206=>"000101001",
  52207=>"110011101",
  52208=>"000010111",
  52209=>"100101000",
  52210=>"011101000",
  52211=>"101111000",
  52212=>"110110001",
  52213=>"001000011",
  52214=>"110110000",
  52215=>"101001010",
  52216=>"001100110",
  52217=>"111100110",
  52218=>"110011110",
  52219=>"110110010",
  52220=>"101101111",
  52221=>"111100011",
  52222=>"010010001",
  52223=>"011110111",
  52224=>"110000100",
  52225=>"010011101",
  52226=>"100110010",
  52227=>"000101001",
  52228=>"000111111",
  52229=>"001010110",
  52230=>"111100110",
  52231=>"111111111",
  52232=>"110100110",
  52233=>"101001111",
  52234=>"000011011",
  52235=>"010000100",
  52236=>"111011111",
  52237=>"011110100",
  52238=>"001000011",
  52239=>"000000001",
  52240=>"101101110",
  52241=>"101111011",
  52242=>"101111111",
  52243=>"100110100",
  52244=>"011100010",
  52245=>"101100010",
  52246=>"010010001",
  52247=>"111110100",
  52248=>"110000011",
  52249=>"100000001",
  52250=>"010000110",
  52251=>"111111010",
  52252=>"100000101",
  52253=>"100011011",
  52254=>"111100001",
  52255=>"101111011",
  52256=>"111010001",
  52257=>"011001111",
  52258=>"011010111",
  52259=>"111000010",
  52260=>"111101101",
  52261=>"101101011",
  52262=>"110000000",
  52263=>"111001001",
  52264=>"001001100",
  52265=>"111101011",
  52266=>"001011010",
  52267=>"001010111",
  52268=>"111000001",
  52269=>"001101111",
  52270=>"101010011",
  52271=>"011010111",
  52272=>"111101001",
  52273=>"011100111",
  52274=>"111000100",
  52275=>"000110011",
  52276=>"101100101",
  52277=>"110100010",
  52278=>"010110111",
  52279=>"111110100",
  52280=>"111010001",
  52281=>"101100011",
  52282=>"011010001",
  52283=>"001001001",
  52284=>"011001001",
  52285=>"001010001",
  52286=>"111001000",
  52287=>"011011111",
  52288=>"011010110",
  52289=>"111100100",
  52290=>"011111100",
  52291=>"001101100",
  52292=>"000001100",
  52293=>"011100000",
  52294=>"111011100",
  52295=>"101100010",
  52296=>"011010101",
  52297=>"011100100",
  52298=>"001111110",
  52299=>"101001110",
  52300=>"100010011",
  52301=>"110101000",
  52302=>"010011011",
  52303=>"001111101",
  52304=>"001000111",
  52305=>"001011111",
  52306=>"010010110",
  52307=>"000001110",
  52308=>"011100100",
  52309=>"101010101",
  52310=>"110110100",
  52311=>"111111001",
  52312=>"000100000",
  52313=>"110111111",
  52314=>"101111110",
  52315=>"000000000",
  52316=>"001001111",
  52317=>"010011000",
  52318=>"000000000",
  52319=>"010101110",
  52320=>"110010111",
  52321=>"011010100",
  52322=>"011100001",
  52323=>"010001000",
  52324=>"100000000",
  52325=>"011110011",
  52326=>"110110111",
  52327=>"011111111",
  52328=>"111001111",
  52329=>"100110100",
  52330=>"110000001",
  52331=>"011011011",
  52332=>"101001111",
  52333=>"101001110",
  52334=>"011111100",
  52335=>"000001111",
  52336=>"100001101",
  52337=>"110101010",
  52338=>"011111000",
  52339=>"110000001",
  52340=>"111111101",
  52341=>"001000111",
  52342=>"101110000",
  52343=>"000101111",
  52344=>"110111110",
  52345=>"000110010",
  52346=>"011101000",
  52347=>"110110011",
  52348=>"100110100",
  52349=>"000100000",
  52350=>"011011111",
  52351=>"110010011",
  52352=>"101110001",
  52353=>"110010100",
  52354=>"011111111",
  52355=>"000111101",
  52356=>"100111100",
  52357=>"111100111",
  52358=>"011011000",
  52359=>"001100100",
  52360=>"000111000",
  52361=>"110111011",
  52362=>"100011111",
  52363=>"111101000",
  52364=>"100000001",
  52365=>"101000001",
  52366=>"001001001",
  52367=>"101100001",
  52368=>"001000011",
  52369=>"011010001",
  52370=>"001000000",
  52371=>"001000010",
  52372=>"011001000",
  52373=>"100010110",
  52374=>"111001111",
  52375=>"111001001",
  52376=>"111011000",
  52377=>"100100001",
  52378=>"010010000",
  52379=>"001110111",
  52380=>"111101011",
  52381=>"000000000",
  52382=>"001101001",
  52383=>"100110001",
  52384=>"101011001",
  52385=>"110010101",
  52386=>"111011100",
  52387=>"001000111",
  52388=>"110011111",
  52389=>"110000000",
  52390=>"101000001",
  52391=>"110101100",
  52392=>"110111100",
  52393=>"001101011",
  52394=>"010110100",
  52395=>"000110101",
  52396=>"101011100",
  52397=>"101000110",
  52398=>"110000010",
  52399=>"011011111",
  52400=>"111111000",
  52401=>"000001101",
  52402=>"111100000",
  52403=>"000111010",
  52404=>"001011010",
  52405=>"100001010",
  52406=>"101111101",
  52407=>"100011110",
  52408=>"101110000",
  52409=>"010001101",
  52410=>"111110011",
  52411=>"110000000",
  52412=>"010111100",
  52413=>"011000101",
  52414=>"011101000",
  52415=>"000111101",
  52416=>"101101101",
  52417=>"010011011",
  52418=>"011111101",
  52419=>"111011011",
  52420=>"111111100",
  52421=>"110011001",
  52422=>"111001001",
  52423=>"110110111",
  52424=>"101010111",
  52425=>"111111111",
  52426=>"110000000",
  52427=>"010011111",
  52428=>"000100111",
  52429=>"001011001",
  52430=>"111000101",
  52431=>"001001101",
  52432=>"101001001",
  52433=>"011010011",
  52434=>"011011010",
  52435=>"001001110",
  52436=>"101110100",
  52437=>"000111011",
  52438=>"000111101",
  52439=>"101011111",
  52440=>"001000011",
  52441=>"100101111",
  52442=>"010000100",
  52443=>"101111110",
  52444=>"101001110",
  52445=>"100010010",
  52446=>"010111000",
  52447=>"010011011",
  52448=>"001000010",
  52449=>"000011011",
  52450=>"110001110",
  52451=>"111111011",
  52452=>"101011011",
  52453=>"101000101",
  52454=>"001100001",
  52455=>"110111010",
  52456=>"111011111",
  52457=>"001111011",
  52458=>"011111011",
  52459=>"110001111",
  52460=>"000011000",
  52461=>"111101010",
  52462=>"001111110",
  52463=>"011010101",
  52464=>"110001001",
  52465=>"111011000",
  52466=>"101110111",
  52467=>"100101110",
  52468=>"110111101",
  52469=>"001000111",
  52470=>"011000000",
  52471=>"101111010",
  52472=>"000110001",
  52473=>"010000000",
  52474=>"001101101",
  52475=>"000011001",
  52476=>"011100000",
  52477=>"001110001",
  52478=>"011110111",
  52479=>"011100110",
  52480=>"111100110",
  52481=>"100100100",
  52482=>"110100100",
  52483=>"110000010",
  52484=>"000000011",
  52485=>"111101010",
  52486=>"000101011",
  52487=>"011000000",
  52488=>"110111101",
  52489=>"101111110",
  52490=>"011011000",
  52491=>"110101100",
  52492=>"001010111",
  52493=>"010100000",
  52494=>"101011100",
  52495=>"101001010",
  52496=>"001010100",
  52497=>"001100011",
  52498=>"100000110",
  52499=>"110000101",
  52500=>"000011001",
  52501=>"001001000",
  52502=>"001111111",
  52503=>"010010001",
  52504=>"111110111",
  52505=>"111101101",
  52506=>"000100011",
  52507=>"111010101",
  52508=>"011111011",
  52509=>"101001100",
  52510=>"101001110",
  52511=>"111011100",
  52512=>"101011000",
  52513=>"100000011",
  52514=>"101010101",
  52515=>"101111101",
  52516=>"100100100",
  52517=>"000000000",
  52518=>"001010011",
  52519=>"011010010",
  52520=>"000110110",
  52521=>"001110001",
  52522=>"010001001",
  52523=>"011000111",
  52524=>"110011001",
  52525=>"000100100",
  52526=>"111111111",
  52527=>"001100000",
  52528=>"001000000",
  52529=>"100101110",
  52530=>"110111011",
  52531=>"100101111",
  52532=>"010100011",
  52533=>"011111000",
  52534=>"100110111",
  52535=>"100110010",
  52536=>"110100110",
  52537=>"001100111",
  52538=>"000001011",
  52539=>"000111000",
  52540=>"110010010",
  52541=>"001111100",
  52542=>"000110110",
  52543=>"101000000",
  52544=>"000101001",
  52545=>"011000111",
  52546=>"111011111",
  52547=>"011100011",
  52548=>"101001001",
  52549=>"010100011",
  52550=>"011110110",
  52551=>"000011101",
  52552=>"001100001",
  52553=>"111110010",
  52554=>"100000101",
  52555=>"000101100",
  52556=>"011001000",
  52557=>"000001011",
  52558=>"001001000",
  52559=>"100010100",
  52560=>"000101000",
  52561=>"111110001",
  52562=>"000000100",
  52563=>"010000010",
  52564=>"011001001",
  52565=>"101110010",
  52566=>"111110011",
  52567=>"000100111",
  52568=>"001010111",
  52569=>"101001101",
  52570=>"000111010",
  52571=>"010000111",
  52572=>"100001001",
  52573=>"100000111",
  52574=>"011100111",
  52575=>"111100011",
  52576=>"011011000",
  52577=>"011011101",
  52578=>"110101000",
  52579=>"110110011",
  52580=>"011000100",
  52581=>"001000001",
  52582=>"101110001",
  52583=>"010110010",
  52584=>"011000111",
  52585=>"101001011",
  52586=>"100101010",
  52587=>"110110011",
  52588=>"011101101",
  52589=>"101001100",
  52590=>"011000011",
  52591=>"101011101",
  52592=>"100110111",
  52593=>"101110111",
  52594=>"101111100",
  52595=>"011001001",
  52596=>"110110100",
  52597=>"011100001",
  52598=>"011111010",
  52599=>"010100101",
  52600=>"011000011",
  52601=>"001011100",
  52602=>"110101000",
  52603=>"000110010",
  52604=>"110101001",
  52605=>"110010001",
  52606=>"010011111",
  52607=>"000010100",
  52608=>"000000100",
  52609=>"111001110",
  52610=>"100100010",
  52611=>"001101011",
  52612=>"100001111",
  52613=>"000011111",
  52614=>"100001001",
  52615=>"000101000",
  52616=>"111101011",
  52617=>"110110010",
  52618=>"100001000",
  52619=>"101111111",
  52620=>"111001010",
  52621=>"011000100",
  52622=>"000101101",
  52623=>"000011100",
  52624=>"010110011",
  52625=>"000110011",
  52626=>"100010101",
  52627=>"110111101",
  52628=>"001111001",
  52629=>"101110100",
  52630=>"010001101",
  52631=>"000101000",
  52632=>"000110000",
  52633=>"010111001",
  52634=>"100010001",
  52635=>"001000100",
  52636=>"100110011",
  52637=>"110100000",
  52638=>"111101110",
  52639=>"010000100",
  52640=>"010011100",
  52641=>"011010000",
  52642=>"011000011",
  52643=>"010110011",
  52644=>"001001100",
  52645=>"100000100",
  52646=>"010011000",
  52647=>"010010101",
  52648=>"111110001",
  52649=>"001000000",
  52650=>"001011011",
  52651=>"010000101",
  52652=>"110000010",
  52653=>"111110011",
  52654=>"101111011",
  52655=>"010010001",
  52656=>"000111001",
  52657=>"011000000",
  52658=>"010001000",
  52659=>"110101001",
  52660=>"110100001",
  52661=>"011010010",
  52662=>"101011111",
  52663=>"011011110",
  52664=>"110110100",
  52665=>"011100000",
  52666=>"001011111",
  52667=>"100000111",
  52668=>"101100100",
  52669=>"001011010",
  52670=>"001100000",
  52671=>"010010110",
  52672=>"011110001",
  52673=>"001000011",
  52674=>"011111001",
  52675=>"100000111",
  52676=>"001000011",
  52677=>"101011001",
  52678=>"111101000",
  52679=>"000000110",
  52680=>"001110101",
  52681=>"000101010",
  52682=>"111000001",
  52683=>"001101011",
  52684=>"001000110",
  52685=>"101101100",
  52686=>"101111110",
  52687=>"111100010",
  52688=>"100100101",
  52689=>"011111010",
  52690=>"111111001",
  52691=>"011001000",
  52692=>"110110111",
  52693=>"111101010",
  52694=>"110000111",
  52695=>"010111001",
  52696=>"010110000",
  52697=>"001101011",
  52698=>"001011011",
  52699=>"011011001",
  52700=>"010001110",
  52701=>"011010010",
  52702=>"001110011",
  52703=>"100101100",
  52704=>"100011100",
  52705=>"000001101",
  52706=>"000001001",
  52707=>"001110011",
  52708=>"110001001",
  52709=>"110101001",
  52710=>"100010100",
  52711=>"110101101",
  52712=>"010010000",
  52713=>"000001100",
  52714=>"101000011",
  52715=>"010010000",
  52716=>"111111001",
  52717=>"111001001",
  52718=>"111100000",
  52719=>"111000101",
  52720=>"100101010",
  52721=>"001101001",
  52722=>"010010111",
  52723=>"011000001",
  52724=>"100111111",
  52725=>"000001000",
  52726=>"100011010",
  52727=>"111000101",
  52728=>"110111101",
  52729=>"011000011",
  52730=>"000010000",
  52731=>"000111001",
  52732=>"110001010",
  52733=>"000010100",
  52734=>"101011010",
  52735=>"011101110",
  52736=>"101000100",
  52737=>"000101000",
  52738=>"011001001",
  52739=>"011001011",
  52740=>"111111001",
  52741=>"100100101",
  52742=>"011000011",
  52743=>"111001100",
  52744=>"111110101",
  52745=>"111001001",
  52746=>"111000111",
  52747=>"100010101",
  52748=>"110110010",
  52749=>"111100100",
  52750=>"101101111",
  52751=>"001001111",
  52752=>"101101011",
  52753=>"110111001",
  52754=>"110101111",
  52755=>"001001101",
  52756=>"011101011",
  52757=>"111011000",
  52758=>"000001011",
  52759=>"010111111",
  52760=>"110111011",
  52761=>"011011001",
  52762=>"111000000",
  52763=>"001101110",
  52764=>"111001101",
  52765=>"110101110",
  52766=>"001011001",
  52767=>"000000000",
  52768=>"001011111",
  52769=>"111100111",
  52770=>"010010001",
  52771=>"110010000",
  52772=>"001111111",
  52773=>"000010011",
  52774=>"000101011",
  52775=>"001011111",
  52776=>"001110001",
  52777=>"011011000",
  52778=>"001110001",
  52779=>"001101001",
  52780=>"011010111",
  52781=>"101110000",
  52782=>"010011000",
  52783=>"101000011",
  52784=>"001111111",
  52785=>"101001011",
  52786=>"111011101",
  52787=>"100100000",
  52788=>"011111110",
  52789=>"001101000",
  52790=>"110001110",
  52791=>"110011111",
  52792=>"100000000",
  52793=>"110001010",
  52794=>"101100110",
  52795=>"111000001",
  52796=>"010111000",
  52797=>"011001111",
  52798=>"010101011",
  52799=>"110100101",
  52800=>"100101111",
  52801=>"001111000",
  52802=>"101100111",
  52803=>"110100100",
  52804=>"111100111",
  52805=>"011010000",
  52806=>"101100101",
  52807=>"101001011",
  52808=>"011111111",
  52809=>"100110111",
  52810=>"000101111",
  52811=>"000000001",
  52812=>"111001011",
  52813=>"000001001",
  52814=>"110001010",
  52815=>"100011101",
  52816=>"011001000",
  52817=>"010010101",
  52818=>"011001111",
  52819=>"111100011",
  52820=>"010111001",
  52821=>"010010110",
  52822=>"101001110",
  52823=>"001010000",
  52824=>"000111111",
  52825=>"101011111",
  52826=>"111101000",
  52827=>"111001010",
  52828=>"001000110",
  52829=>"000000010",
  52830=>"001000001",
  52831=>"011010001",
  52832=>"110101000",
  52833=>"001111011",
  52834=>"001000100",
  52835=>"010110011",
  52836=>"110011110",
  52837=>"110100101",
  52838=>"000000000",
  52839=>"000100001",
  52840=>"010100100",
  52841=>"111011110",
  52842=>"100011001",
  52843=>"010110100",
  52844=>"110111101",
  52845=>"011011110",
  52846=>"101001110",
  52847=>"000100101",
  52848=>"110100011",
  52849=>"100111101",
  52850=>"011000011",
  52851=>"011001001",
  52852=>"110011111",
  52853=>"101100111",
  52854=>"001110111",
  52855=>"001000110",
  52856=>"101010111",
  52857=>"011101100",
  52858=>"110001001",
  52859=>"110111111",
  52860=>"110100001",
  52861=>"101001001",
  52862=>"010101000",
  52863=>"110010110",
  52864=>"110001011",
  52865=>"100000101",
  52866=>"001001101",
  52867=>"000001111",
  52868=>"011011111",
  52869=>"101010111",
  52870=>"110010101",
  52871=>"110100100",
  52872=>"010010011",
  52873=>"011011001",
  52874=>"011100001",
  52875=>"110110111",
  52876=>"111001100",
  52877=>"111010111",
  52878=>"010000000",
  52879=>"001001001",
  52880=>"100101001",
  52881=>"000010011",
  52882=>"100110101",
  52883=>"100101101",
  52884=>"011010101",
  52885=>"101000001",
  52886=>"111111101",
  52887=>"101011011",
  52888=>"011000101",
  52889=>"111101010",
  52890=>"000010110",
  52891=>"100111010",
  52892=>"111001101",
  52893=>"011011001",
  52894=>"100010100",
  52895=>"011000100",
  52896=>"001010000",
  52897=>"011001100",
  52898=>"111100000",
  52899=>"100001100",
  52900=>"001101011",
  52901=>"111001111",
  52902=>"100010010",
  52903=>"001001100",
  52904=>"111010000",
  52905=>"110111000",
  52906=>"110011100",
  52907=>"101010100",
  52908=>"000110010",
  52909=>"110111001",
  52910=>"001111001",
  52911=>"100100000",
  52912=>"011011111",
  52913=>"011001010",
  52914=>"011010011",
  52915=>"011000010",
  52916=>"101001001",
  52917=>"111111010",
  52918=>"101011001",
  52919=>"011000000",
  52920=>"111110001",
  52921=>"001101100",
  52922=>"101111001",
  52923=>"000000111",
  52924=>"100100100",
  52925=>"011111011",
  52926=>"001100000",
  52927=>"001001111",
  52928=>"101011100",
  52929=>"110100110",
  52930=>"000110010",
  52931=>"001110111",
  52932=>"110100100",
  52933=>"010100100",
  52934=>"111000011",
  52935=>"011001011",
  52936=>"011010001",
  52937=>"011011001",
  52938=>"101010100",
  52939=>"111110101",
  52940=>"100000010",
  52941=>"110000010",
  52942=>"111101110",
  52943=>"011000110",
  52944=>"111111000",
  52945=>"101100100",
  52946=>"001110010",
  52947=>"101111110",
  52948=>"010000000",
  52949=>"011110011",
  52950=>"011101000",
  52951=>"010011000",
  52952=>"100000100",
  52953=>"111001110",
  52954=>"001110010",
  52955=>"001011011",
  52956=>"111100110",
  52957=>"110100000",
  52958=>"101001111",
  52959=>"111101111",
  52960=>"101110011",
  52961=>"100101001",
  52962=>"010001101",
  52963=>"111010010",
  52964=>"010100000",
  52965=>"111001100",
  52966=>"100010011",
  52967=>"111111111",
  52968=>"010000010",
  52969=>"101111000",
  52970=>"011111111",
  52971=>"001101111",
  52972=>"101110011",
  52973=>"110101011",
  52974=>"110110111",
  52975=>"011011001",
  52976=>"000101111",
  52977=>"101010011",
  52978=>"000101111",
  52979=>"001110000",
  52980=>"000110000",
  52981=>"110110111",
  52982=>"000010010",
  52983=>"001101101",
  52984=>"101111101",
  52985=>"001111001",
  52986=>"000110101",
  52987=>"101011001",
  52988=>"000100010",
  52989=>"000111000",
  52990=>"101111000",
  52991=>"011011011",
  52992=>"011001101",
  52993=>"001011111",
  52994=>"111000101",
  52995=>"111111000",
  52996=>"010111000",
  52997=>"011111011",
  52998=>"010101111",
  52999=>"110001011",
  53000=>"000000100",
  53001=>"010111010",
  53002=>"011001001",
  53003=>"011000001",
  53004=>"101010000",
  53005=>"111110101",
  53006=>"000100110",
  53007=>"111011010",
  53008=>"011001011",
  53009=>"001001100",
  53010=>"111011110",
  53011=>"101101111",
  53012=>"001110000",
  53013=>"101101000",
  53014=>"110100101",
  53015=>"011001111",
  53016=>"001011111",
  53017=>"111111011",
  53018=>"100010100",
  53019=>"110010111",
  53020=>"011111100",
  53021=>"000010011",
  53022=>"000111110",
  53023=>"000000101",
  53024=>"000110100",
  53025=>"111110111",
  53026=>"111110101",
  53027=>"011101111",
  53028=>"001010100",
  53029=>"011100010",
  53030=>"110000110",
  53031=>"110000100",
  53032=>"000000100",
  53033=>"111101101",
  53034=>"111010001",
  53035=>"001000101",
  53036=>"101000101",
  53037=>"001101000",
  53038=>"111001001",
  53039=>"001001010",
  53040=>"111011110",
  53041=>"101111001",
  53042=>"101110100",
  53043=>"000110000",
  53044=>"000010000",
  53045=>"100000010",
  53046=>"000011011",
  53047=>"011110110",
  53048=>"110111010",
  53049=>"101011010",
  53050=>"100110100",
  53051=>"101110111",
  53052=>"001011010",
  53053=>"101111000",
  53054=>"001101011",
  53055=>"110010000",
  53056=>"000011100",
  53057=>"011110000",
  53058=>"101010101",
  53059=>"001010110",
  53060=>"010001011",
  53061=>"011110010",
  53062=>"011011001",
  53063=>"101100010",
  53064=>"111110010",
  53065=>"100111111",
  53066=>"101011000",
  53067=>"001000010",
  53068=>"110000011",
  53069=>"111010011",
  53070=>"010000101",
  53071=>"010110111",
  53072=>"011010000",
  53073=>"110110010",
  53074=>"001001000",
  53075=>"111001011",
  53076=>"101110011",
  53077=>"110101100",
  53078=>"010000111",
  53079=>"110110101",
  53080=>"111100110",
  53081=>"011010100",
  53082=>"110000101",
  53083=>"000011101",
  53084=>"101001111",
  53085=>"000110111",
  53086=>"110110110",
  53087=>"100111011",
  53088=>"110111001",
  53089=>"011010001",
  53090=>"011000011",
  53091=>"101010011",
  53092=>"100000111",
  53093=>"101110000",
  53094=>"010000000",
  53095=>"110100101",
  53096=>"001011101",
  53097=>"110001011",
  53098=>"110111001",
  53099=>"000011110",
  53100=>"101001111",
  53101=>"001111111",
  53102=>"010000101",
  53103=>"010110100",
  53104=>"001000000",
  53105=>"111011111",
  53106=>"011001101",
  53107=>"011000011",
  53108=>"001011010",
  53109=>"001101111",
  53110=>"111011110",
  53111=>"111111000",
  53112=>"011011000",
  53113=>"111101110",
  53114=>"000100101",
  53115=>"000010010",
  53116=>"011011011",
  53117=>"111101010",
  53118=>"010001000",
  53119=>"110011000",
  53120=>"001001100",
  53121=>"101111011",
  53122=>"111100111",
  53123=>"110001110",
  53124=>"101110111",
  53125=>"001000111",
  53126=>"101111111",
  53127=>"110010100",
  53128=>"000010010",
  53129=>"010110001",
  53130=>"000010001",
  53131=>"000100111",
  53132=>"111010011",
  53133=>"101111011",
  53134=>"100010011",
  53135=>"100011111",
  53136=>"001110100",
  53137=>"110000110",
  53138=>"010110110",
  53139=>"000010000",
  53140=>"001111100",
  53141=>"111101000",
  53142=>"001111001",
  53143=>"001001111",
  53144=>"111101001",
  53145=>"011001000",
  53146=>"000010011",
  53147=>"001000101",
  53148=>"010011100",
  53149=>"000111110",
  53150=>"010011011",
  53151=>"011000010",
  53152=>"011011111",
  53153=>"001001001",
  53154=>"101111011",
  53155=>"100000000",
  53156=>"011011101",
  53157=>"010001100",
  53158=>"000000011",
  53159=>"101101111",
  53160=>"011110001",
  53161=>"111110001",
  53162=>"100011011",
  53163=>"101010010",
  53164=>"010100101",
  53165=>"100111101",
  53166=>"001010100",
  53167=>"010001100",
  53168=>"110110100",
  53169=>"000110110",
  53170=>"011001001",
  53171=>"000000111",
  53172=>"010101110",
  53173=>"000110110",
  53174=>"001001010",
  53175=>"001001111",
  53176=>"011100111",
  53177=>"001010101",
  53178=>"100111110",
  53179=>"111010000",
  53180=>"010011101",
  53181=>"111110100",
  53182=>"000111111",
  53183=>"100000000",
  53184=>"100000010",
  53185=>"110000101",
  53186=>"110100101",
  53187=>"010010101",
  53188=>"011011101",
  53189=>"111111101",
  53190=>"001101111",
  53191=>"001101001",
  53192=>"101100110",
  53193=>"110011001",
  53194=>"100100011",
  53195=>"000111001",
  53196=>"111000011",
  53197=>"110010000",
  53198=>"000110000",
  53199=>"110011100",
  53200=>"000000011",
  53201=>"011110101",
  53202=>"111101010",
  53203=>"011011111",
  53204=>"111101000",
  53205=>"101010111",
  53206=>"010001001",
  53207=>"101110001",
  53208=>"110000011",
  53209=>"001001011",
  53210=>"010110100",
  53211=>"100110101",
  53212=>"101111010",
  53213=>"100101100",
  53214=>"110111000",
  53215=>"011001010",
  53216=>"110110111",
  53217=>"100010010",
  53218=>"001110011",
  53219=>"101001001",
  53220=>"111001011",
  53221=>"001011101",
  53222=>"100010101",
  53223=>"001111100",
  53224=>"111101000",
  53225=>"010011010",
  53226=>"100011011",
  53227=>"110001110",
  53228=>"100010111",
  53229=>"001111011",
  53230=>"000100001",
  53231=>"010011110",
  53232=>"000100001",
  53233=>"001100000",
  53234=>"111010110",
  53235=>"011110011",
  53236=>"001100100",
  53237=>"111100000",
  53238=>"010101011",
  53239=>"111101111",
  53240=>"000110000",
  53241=>"100110100",
  53242=>"100001111",
  53243=>"010010100",
  53244=>"001001001",
  53245=>"100100100",
  53246=>"110001101",
  53247=>"111111010",
  53248=>"111011111",
  53249=>"110000100",
  53250=>"111000001",
  53251=>"111110000",
  53252=>"011000010",
  53253=>"000010100",
  53254=>"001110110",
  53255=>"100001100",
  53256=>"011000110",
  53257=>"100000100",
  53258=>"010010110",
  53259=>"001100111",
  53260=>"110000010",
  53261=>"100010110",
  53262=>"101010101",
  53263=>"001000001",
  53264=>"111010010",
  53265=>"101111000",
  53266=>"011001101",
  53267=>"000101111",
  53268=>"110001111",
  53269=>"111101101",
  53270=>"101100101",
  53271=>"110010110",
  53272=>"111001001",
  53273=>"110000011",
  53274=>"111011010",
  53275=>"111100011",
  53276=>"011100011",
  53277=>"011100101",
  53278=>"011101001",
  53279=>"100000101",
  53280=>"001010101",
  53281=>"000010011",
  53282=>"101100000",
  53283=>"101010111",
  53284=>"000011101",
  53285=>"100011111",
  53286=>"110100000",
  53287=>"001110010",
  53288=>"000111001",
  53289=>"100100110",
  53290=>"011001001",
  53291=>"000110000",
  53292=>"101100110",
  53293=>"110001100",
  53294=>"110001111",
  53295=>"001111010",
  53296=>"111101110",
  53297=>"101100011",
  53298=>"010101010",
  53299=>"010001000",
  53300=>"011000100",
  53301=>"011101011",
  53302=>"100110101",
  53303=>"011111101",
  53304=>"100000000",
  53305=>"101100011",
  53306=>"111000110",
  53307=>"010000100",
  53308=>"101101100",
  53309=>"111100000",
  53310=>"100111101",
  53311=>"011110011",
  53312=>"000101111",
  53313=>"000000000",
  53314=>"100110001",
  53315=>"100000101",
  53316=>"001000011",
  53317=>"110111010",
  53318=>"010111010",
  53319=>"101101101",
  53320=>"010000100",
  53321=>"111111011",
  53322=>"000010001",
  53323=>"110101100",
  53324=>"110000100",
  53325=>"001101110",
  53326=>"011111100",
  53327=>"111111010",
  53328=>"000001000",
  53329=>"000100111",
  53330=>"011101100",
  53331=>"100101001",
  53332=>"011011010",
  53333=>"100001000",
  53334=>"111101000",
  53335=>"101010011",
  53336=>"011011011",
  53337=>"001011101",
  53338=>"111101010",
  53339=>"000000100",
  53340=>"000010111",
  53341=>"010001010",
  53342=>"100100110",
  53343=>"001010011",
  53344=>"011111011",
  53345=>"001011000",
  53346=>"001100101",
  53347=>"000011111",
  53348=>"001001100",
  53349=>"110110100",
  53350=>"011100010",
  53351=>"001111110",
  53352=>"011100001",
  53353=>"000101001",
  53354=>"100001100",
  53355=>"110100001",
  53356=>"100110101",
  53357=>"011010111",
  53358=>"001101000",
  53359=>"001001000",
  53360=>"101010001",
  53361=>"011000000",
  53362=>"101010110",
  53363=>"011111011",
  53364=>"001000001",
  53365=>"010110010",
  53366=>"001110000",
  53367=>"010100111",
  53368=>"011000011",
  53369=>"001000001",
  53370=>"010001111",
  53371=>"111110001",
  53372=>"000011000",
  53373=>"110010000",
  53374=>"010011101",
  53375=>"000111001",
  53376=>"101011001",
  53377=>"110100101",
  53378=>"000101001",
  53379=>"000001111",
  53380=>"101000101",
  53381=>"101111010",
  53382=>"100111110",
  53383=>"111001001",
  53384=>"000110111",
  53385=>"110111000",
  53386=>"000011000",
  53387=>"010111001",
  53388=>"000010110",
  53389=>"100001011",
  53390=>"100101100",
  53391=>"100000110",
  53392=>"001000111",
  53393=>"110100111",
  53394=>"111001010",
  53395=>"010101100",
  53396=>"101011000",
  53397=>"101000101",
  53398=>"111001001",
  53399=>"010001101",
  53400=>"110101111",
  53401=>"010000111",
  53402=>"111111001",
  53403=>"110110101",
  53404=>"100001100",
  53405=>"101101111",
  53406=>"001011110",
  53407=>"101011100",
  53408=>"000101111",
  53409=>"011011101",
  53410=>"110011001",
  53411=>"110000000",
  53412=>"010011101",
  53413=>"111011110",
  53414=>"110010000",
  53415=>"100010010",
  53416=>"010101111",
  53417=>"010100110",
  53418=>"100001000",
  53419=>"100110101",
  53420=>"101001111",
  53421=>"111001010",
  53422=>"100111100",
  53423=>"010010111",
  53424=>"000001100",
  53425=>"101101010",
  53426=>"111001000",
  53427=>"101000000",
  53428=>"001000001",
  53429=>"101001111",
  53430=>"010000000",
  53431=>"011100011",
  53432=>"001001100",
  53433=>"010110101",
  53434=>"000010010",
  53435=>"001110000",
  53436=>"000100000",
  53437=>"000001111",
  53438=>"110100111",
  53439=>"100101011",
  53440=>"101110001",
  53441=>"010101001",
  53442=>"110011110",
  53443=>"000110101",
  53444=>"010111100",
  53445=>"001010100",
  53446=>"011001001",
  53447=>"000001010",
  53448=>"001010010",
  53449=>"110010000",
  53450=>"000010000",
  53451=>"010111000",
  53452=>"010111111",
  53453=>"001000011",
  53454=>"101110000",
  53455=>"110000011",
  53456=>"011010111",
  53457=>"100111010",
  53458=>"110010110",
  53459=>"101000001",
  53460=>"101010111",
  53461=>"111001110",
  53462=>"110110001",
  53463=>"101100010",
  53464=>"001000001",
  53465=>"110000000",
  53466=>"010000001",
  53467=>"110101110",
  53468=>"000110101",
  53469=>"000101100",
  53470=>"011000000",
  53471=>"000000100",
  53472=>"001100101",
  53473=>"101000111",
  53474=>"110101010",
  53475=>"110100101",
  53476=>"011000100",
  53477=>"010111000",
  53478=>"101100001",
  53479=>"110001000",
  53480=>"100010010",
  53481=>"011010100",
  53482=>"000100010",
  53483=>"001000100",
  53484=>"001001100",
  53485=>"001000101",
  53486=>"101000010",
  53487=>"000101010",
  53488=>"011110111",
  53489=>"001100000",
  53490=>"011000111",
  53491=>"001110010",
  53492=>"101000010",
  53493=>"101101011",
  53494=>"001011101",
  53495=>"010000000",
  53496=>"010100111",
  53497=>"010101111",
  53498=>"010111100",
  53499=>"001000100",
  53500=>"011111010",
  53501=>"101000001",
  53502=>"000000010",
  53503=>"111010001",
  53504=>"101001110",
  53505=>"011001010",
  53506=>"100011111",
  53507=>"000011111",
  53508=>"010000001",
  53509=>"110000000",
  53510=>"000110111",
  53511=>"111001110",
  53512=>"010110010",
  53513=>"011101110",
  53514=>"100110100",
  53515=>"110111111",
  53516=>"000010000",
  53517=>"110001100",
  53518=>"111000010",
  53519=>"011110010",
  53520=>"111011000",
  53521=>"100001001",
  53522=>"110111111",
  53523=>"110100101",
  53524=>"000001110",
  53525=>"011000011",
  53526=>"000000000",
  53527=>"011010101",
  53528=>"011100101",
  53529=>"011010101",
  53530=>"110000110",
  53531=>"010110010",
  53532=>"100101111",
  53533=>"010001000",
  53534=>"100101101",
  53535=>"000000100",
  53536=>"101000110",
  53537=>"111101100",
  53538=>"100001000",
  53539=>"111101111",
  53540=>"001111000",
  53541=>"000000000",
  53542=>"010010100",
  53543=>"101000111",
  53544=>"000001011",
  53545=>"100101111",
  53546=>"010001011",
  53547=>"001011000",
  53548=>"110101110",
  53549=>"110010001",
  53550=>"000001010",
  53551=>"001010110",
  53552=>"100111001",
  53553=>"110111000",
  53554=>"100000110",
  53555=>"110001000",
  53556=>"000000001",
  53557=>"100000111",
  53558=>"000101110",
  53559=>"110001111",
  53560=>"000110000",
  53561=>"101000100",
  53562=>"001111100",
  53563=>"111011011",
  53564=>"001111100",
  53565=>"110000010",
  53566=>"010000010",
  53567=>"001110111",
  53568=>"101101001",
  53569=>"111110001",
  53570=>"011110111",
  53571=>"111101000",
  53572=>"000110111",
  53573=>"110101111",
  53574=>"110000010",
  53575=>"000001000",
  53576=>"011011001",
  53577=>"111100011",
  53578=>"001100001",
  53579=>"101001000",
  53580=>"111111100",
  53581=>"000010110",
  53582=>"010101100",
  53583=>"111000101",
  53584=>"110111110",
  53585=>"111101010",
  53586=>"011000101",
  53587=>"101000000",
  53588=>"010100010",
  53589=>"000001110",
  53590=>"101011000",
  53591=>"110011101",
  53592=>"111001000",
  53593=>"010011111",
  53594=>"001011011",
  53595=>"000110100",
  53596=>"100110011",
  53597=>"001101100",
  53598=>"110010010",
  53599=>"000110011",
  53600=>"000000111",
  53601=>"010100100",
  53602=>"011110100",
  53603=>"001001000",
  53604=>"101110110",
  53605=>"011011000",
  53606=>"011100101",
  53607=>"010111101",
  53608=>"100001001",
  53609=>"011101011",
  53610=>"011100011",
  53611=>"100110101",
  53612=>"100011000",
  53613=>"010111110",
  53614=>"100100110",
  53615=>"010100101",
  53616=>"110011001",
  53617=>"101001011",
  53618=>"010110001",
  53619=>"001100000",
  53620=>"100111011",
  53621=>"111100001",
  53622=>"000000100",
  53623=>"001001010",
  53624=>"110010011",
  53625=>"011000000",
  53626=>"111000100",
  53627=>"110110001",
  53628=>"000110110",
  53629=>"101011111",
  53630=>"010001100",
  53631=>"101110011",
  53632=>"101111101",
  53633=>"001000011",
  53634=>"101001110",
  53635=>"100110110",
  53636=>"110011011",
  53637=>"000111011",
  53638=>"011110111",
  53639=>"000010101",
  53640=>"000011111",
  53641=>"011001100",
  53642=>"100110000",
  53643=>"011000001",
  53644=>"000100100",
  53645=>"001100101",
  53646=>"001101110",
  53647=>"111011000",
  53648=>"001110110",
  53649=>"000011111",
  53650=>"000110011",
  53651=>"000100001",
  53652=>"111000110",
  53653=>"001100101",
  53654=>"001111110",
  53655=>"000010111",
  53656=>"110101110",
  53657=>"100101111",
  53658=>"010110111",
  53659=>"011100101",
  53660=>"100110011",
  53661=>"100000001",
  53662=>"101100111",
  53663=>"111001101",
  53664=>"000111000",
  53665=>"110110000",
  53666=>"110011000",
  53667=>"000000110",
  53668=>"001010010",
  53669=>"100110000",
  53670=>"011000001",
  53671=>"111001111",
  53672=>"010010110",
  53673=>"011010011",
  53674=>"001001100",
  53675=>"000010100",
  53676=>"101000110",
  53677=>"000001111",
  53678=>"000110001",
  53679=>"110110111",
  53680=>"000000001",
  53681=>"110111010",
  53682=>"001010010",
  53683=>"111010100",
  53684=>"000000100",
  53685=>"000010100",
  53686=>"010011001",
  53687=>"111000111",
  53688=>"001110110",
  53689=>"110000001",
  53690=>"100100000",
  53691=>"010000110",
  53692=>"110100000",
  53693=>"010001001",
  53694=>"000110110",
  53695=>"010101000",
  53696=>"001010101",
  53697=>"001000011",
  53698=>"111101000",
  53699=>"100000110",
  53700=>"100011001",
  53701=>"010000101",
  53702=>"111100010",
  53703=>"001000001",
  53704=>"011110000",
  53705=>"101111110",
  53706=>"111001010",
  53707=>"011010010",
  53708=>"010110110",
  53709=>"000110001",
  53710=>"101110011",
  53711=>"010100000",
  53712=>"110001101",
  53713=>"011000011",
  53714=>"001010001",
  53715=>"101111011",
  53716=>"000110111",
  53717=>"100010101",
  53718=>"111101011",
  53719=>"100101101",
  53720=>"111000000",
  53721=>"000101111",
  53722=>"111001100",
  53723=>"000111000",
  53724=>"000001000",
  53725=>"111110101",
  53726=>"010110010",
  53727=>"011111101",
  53728=>"000010011",
  53729=>"001101111",
  53730=>"110110001",
  53731=>"001110011",
  53732=>"011100110",
  53733=>"010100100",
  53734=>"010011010",
  53735=>"011001000",
  53736=>"010111110",
  53737=>"011011101",
  53738=>"000110101",
  53739=>"000110100",
  53740=>"111110100",
  53741=>"011100000",
  53742=>"110100001",
  53743=>"111101001",
  53744=>"011011110",
  53745=>"010000000",
  53746=>"111000001",
  53747=>"111000011",
  53748=>"100110010",
  53749=>"011110011",
  53750=>"111011111",
  53751=>"010111010",
  53752=>"011001010",
  53753=>"011011011",
  53754=>"111100010",
  53755=>"101001111",
  53756=>"110100101",
  53757=>"100001100",
  53758=>"001000001",
  53759=>"000110001",
  53760=>"100001001",
  53761=>"000010101",
  53762=>"001100000",
  53763=>"011010000",
  53764=>"001001000",
  53765=>"101001001",
  53766=>"001011010",
  53767=>"000011011",
  53768=>"110000101",
  53769=>"111011101",
  53770=>"001100011",
  53771=>"110111100",
  53772=>"001110101",
  53773=>"110010100",
  53774=>"100000111",
  53775=>"010110010",
  53776=>"100100101",
  53777=>"111000111",
  53778=>"100111101",
  53779=>"000011110",
  53780=>"001100110",
  53781=>"000010000",
  53782=>"000100110",
  53783=>"011100000",
  53784=>"011100101",
  53785=>"000101100",
  53786=>"110001110",
  53787=>"110000010",
  53788=>"011011111",
  53789=>"000101100",
  53790=>"001101110",
  53791=>"101111111",
  53792=>"010001010",
  53793=>"000101010",
  53794=>"001001000",
  53795=>"010110100",
  53796=>"000100011",
  53797=>"100001111",
  53798=>"111010000",
  53799=>"100100110",
  53800=>"011111111",
  53801=>"011110010",
  53802=>"101010100",
  53803=>"101111001",
  53804=>"010000111",
  53805=>"000011000",
  53806=>"011101111",
  53807=>"001111011",
  53808=>"001111011",
  53809=>"111100101",
  53810=>"110101100",
  53811=>"000001110",
  53812=>"000000100",
  53813=>"000100100",
  53814=>"010101100",
  53815=>"110101100",
  53816=>"100011111",
  53817=>"111101011",
  53818=>"111101011",
  53819=>"001000000",
  53820=>"100111011",
  53821=>"111010011",
  53822=>"110011010",
  53823=>"000101010",
  53824=>"111111000",
  53825=>"111000001",
  53826=>"011001111",
  53827=>"010111000",
  53828=>"011000110",
  53829=>"100101111",
  53830=>"100010000",
  53831=>"111000110",
  53832=>"011111110",
  53833=>"100111110",
  53834=>"011000001",
  53835=>"011101111",
  53836=>"011110111",
  53837=>"010101110",
  53838=>"110100101",
  53839=>"000110001",
  53840=>"100000011",
  53841=>"001001100",
  53842=>"000111100",
  53843=>"001100110",
  53844=>"000001111",
  53845=>"001100101",
  53846=>"010100100",
  53847=>"010100001",
  53848=>"111000011",
  53849=>"011001000",
  53850=>"000100100",
  53851=>"000010100",
  53852=>"010010110",
  53853=>"101001000",
  53854=>"010000000",
  53855=>"101000100",
  53856=>"100000001",
  53857=>"001110001",
  53858=>"010100110",
  53859=>"101010100",
  53860=>"111100010",
  53861=>"011101101",
  53862=>"110011011",
  53863=>"001101101",
  53864=>"100010100",
  53865=>"001000011",
  53866=>"011100101",
  53867=>"011010111",
  53868=>"100000110",
  53869=>"011001011",
  53870=>"000011010",
  53871=>"001000011",
  53872=>"000010010",
  53873=>"100100110",
  53874=>"011110111",
  53875=>"110001101",
  53876=>"101001010",
  53877=>"101110110",
  53878=>"000100010",
  53879=>"000101000",
  53880=>"001010000",
  53881=>"001101000",
  53882=>"001101001",
  53883=>"011010000",
  53884=>"101110010",
  53885=>"110101010",
  53886=>"110101101",
  53887=>"111001111",
  53888=>"100010100",
  53889=>"100000111",
  53890=>"001000111",
  53891=>"100100010",
  53892=>"000101001",
  53893=>"011100100",
  53894=>"101000010",
  53895=>"100101101",
  53896=>"101011010",
  53897=>"000111000",
  53898=>"100110001",
  53899=>"101110101",
  53900=>"011011101",
  53901=>"011101101",
  53902=>"010100110",
  53903=>"100111011",
  53904=>"111101001",
  53905=>"001100111",
  53906=>"001000101",
  53907=>"101000011",
  53908=>"101001000",
  53909=>"000000111",
  53910=>"011000100",
  53911=>"010000011",
  53912=>"000011011",
  53913=>"100010010",
  53914=>"011101000",
  53915=>"101100110",
  53916=>"000011101",
  53917=>"001011001",
  53918=>"101100111",
  53919=>"111001111",
  53920=>"100001010",
  53921=>"101111010",
  53922=>"101101000",
  53923=>"101010100",
  53924=>"111101010",
  53925=>"001011000",
  53926=>"000001101",
  53927=>"001111001",
  53928=>"111001100",
  53929=>"110111101",
  53930=>"000100001",
  53931=>"010000110",
  53932=>"110110010",
  53933=>"000100111",
  53934=>"011111010",
  53935=>"001000101",
  53936=>"000011101",
  53937=>"101110111",
  53938=>"010011100",
  53939=>"000001100",
  53940=>"111011000",
  53941=>"101001000",
  53942=>"011011101",
  53943=>"000010101",
  53944=>"100000001",
  53945=>"100010110",
  53946=>"010011100",
  53947=>"000010101",
  53948=>"011100111",
  53949=>"001010100",
  53950=>"000000000",
  53951=>"100101100",
  53952=>"011000111",
  53953=>"011100111",
  53954=>"000000111",
  53955=>"111011101",
  53956=>"111100011",
  53957=>"110010000",
  53958=>"100010001",
  53959=>"111111010",
  53960=>"110011001",
  53961=>"111001011",
  53962=>"011011001",
  53963=>"000001101",
  53964=>"000111100",
  53965=>"000111100",
  53966=>"001111100",
  53967=>"110101111",
  53968=>"100000001",
  53969=>"001100000",
  53970=>"000000000",
  53971=>"000100001",
  53972=>"010000010",
  53973=>"000000110",
  53974=>"111111111",
  53975=>"010000110",
  53976=>"010000110",
  53977=>"110001001",
  53978=>"001000011",
  53979=>"000100100",
  53980=>"000111111",
  53981=>"100010111",
  53982=>"010100010",
  53983=>"011111100",
  53984=>"000000000",
  53985=>"110000000",
  53986=>"000111011",
  53987=>"000010101",
  53988=>"000001100",
  53989=>"110111011",
  53990=>"000100010",
  53991=>"100001001",
  53992=>"010101101",
  53993=>"110011011",
  53994=>"110001110",
  53995=>"000011100",
  53996=>"011101001",
  53997=>"100111000",
  53998=>"111001000",
  53999=>"101100000",
  54000=>"011101011",
  54001=>"101010101",
  54002=>"101000110",
  54003=>"001010001",
  54004=>"010110010",
  54005=>"100010000",
  54006=>"010101110",
  54007=>"111010111",
  54008=>"011010110",
  54009=>"010001001",
  54010=>"110100111",
  54011=>"110011001",
  54012=>"000000101",
  54013=>"011010111",
  54014=>"100010110",
  54015=>"110000111",
  54016=>"101000010",
  54017=>"010100100",
  54018=>"010000100",
  54019=>"001101010",
  54020=>"110111101",
  54021=>"000000111",
  54022=>"110010110",
  54023=>"111010010",
  54024=>"000100111",
  54025=>"011000010",
  54026=>"101101111",
  54027=>"010010001",
  54028=>"100001010",
  54029=>"110101101",
  54030=>"111010110",
  54031=>"001111000",
  54032=>"000111111",
  54033=>"001100100",
  54034=>"001110011",
  54035=>"011000001",
  54036=>"110101001",
  54037=>"110101111",
  54038=>"101101000",
  54039=>"110111100",
  54040=>"000001100",
  54041=>"000110111",
  54042=>"001111101",
  54043=>"101110101",
  54044=>"110010010",
  54045=>"101011000",
  54046=>"001111111",
  54047=>"011010010",
  54048=>"101101000",
  54049=>"110101111",
  54050=>"001010101",
  54051=>"011000010",
  54052=>"111010100",
  54053=>"100011010",
  54054=>"011011101",
  54055=>"101100001",
  54056=>"000001110",
  54057=>"111011000",
  54058=>"011011010",
  54059=>"101001111",
  54060=>"010000001",
  54061=>"011101010",
  54062=>"000100011",
  54063=>"111110101",
  54064=>"100000111",
  54065=>"010100110",
  54066=>"001010110",
  54067=>"001011001",
  54068=>"111010000",
  54069=>"000111111",
  54070=>"010110100",
  54071=>"100101000",
  54072=>"111010010",
  54073=>"000011001",
  54074=>"001010010",
  54075=>"110111001",
  54076=>"100010011",
  54077=>"101000011",
  54078=>"110100000",
  54079=>"010010110",
  54080=>"010111100",
  54081=>"111100001",
  54082=>"001011001",
  54083=>"111010100",
  54084=>"001110010",
  54085=>"111100100",
  54086=>"011011100",
  54087=>"011111011",
  54088=>"010111101",
  54089=>"011100000",
  54090=>"010001011",
  54091=>"110100101",
  54092=>"111111001",
  54093=>"000000110",
  54094=>"101011011",
  54095=>"000100110",
  54096=>"000011000",
  54097=>"000100010",
  54098=>"011000010",
  54099=>"000010110",
  54100=>"011101111",
  54101=>"011001101",
  54102=>"100001111",
  54103=>"101010101",
  54104=>"110110100",
  54105=>"100101000",
  54106=>"011111010",
  54107=>"111000010",
  54108=>"101001111",
  54109=>"110111010",
  54110=>"010111001",
  54111=>"100000000",
  54112=>"111101110",
  54113=>"111011001",
  54114=>"001001111",
  54115=>"110010000",
  54116=>"100101101",
  54117=>"110101110",
  54118=>"101110000",
  54119=>"001110101",
  54120=>"001000011",
  54121=>"100100110",
  54122=>"000100010",
  54123=>"111101101",
  54124=>"100001101",
  54125=>"111111000",
  54126=>"100111011",
  54127=>"000000011",
  54128=>"100101001",
  54129=>"000000010",
  54130=>"001011010",
  54131=>"101110100",
  54132=>"011010100",
  54133=>"110010110",
  54134=>"100100110",
  54135=>"011000010",
  54136=>"000011010",
  54137=>"010011011",
  54138=>"100000100",
  54139=>"001011001",
  54140=>"001000010",
  54141=>"111000111",
  54142=>"111010101",
  54143=>"110111111",
  54144=>"111011111",
  54145=>"111010000",
  54146=>"000010111",
  54147=>"001001100",
  54148=>"010111101",
  54149=>"011110000",
  54150=>"011101100",
  54151=>"000000111",
  54152=>"000001011",
  54153=>"011011010",
  54154=>"101111001",
  54155=>"001010001",
  54156=>"000110100",
  54157=>"000100100",
  54158=>"100111010",
  54159=>"001010111",
  54160=>"100010111",
  54161=>"111110001",
  54162=>"101010001",
  54163=>"010010011",
  54164=>"001000100",
  54165=>"100011000",
  54166=>"001100111",
  54167=>"011111010",
  54168=>"100100000",
  54169=>"110010101",
  54170=>"100100011",
  54171=>"100110010",
  54172=>"011110111",
  54173=>"100000110",
  54174=>"000100000",
  54175=>"010110100",
  54176=>"010000010",
  54177=>"001110011",
  54178=>"010101101",
  54179=>"110001100",
  54180=>"100000000",
  54181=>"101110011",
  54182=>"101101111",
  54183=>"101000101",
  54184=>"001100011",
  54185=>"100011011",
  54186=>"111101111",
  54187=>"110101101",
  54188=>"111001111",
  54189=>"011010011",
  54190=>"101101101",
  54191=>"010001011",
  54192=>"011010111",
  54193=>"001100111",
  54194=>"001010011",
  54195=>"100101000",
  54196=>"000110101",
  54197=>"110001110",
  54198=>"010000101",
  54199=>"000111110",
  54200=>"000110001",
  54201=>"100001111",
  54202=>"011100111",
  54203=>"010000110",
  54204=>"010110111",
  54205=>"111010001",
  54206=>"001011001",
  54207=>"010011111",
  54208=>"001110001",
  54209=>"000111010",
  54210=>"101001011",
  54211=>"010110000",
  54212=>"101010011",
  54213=>"011111110",
  54214=>"110011010",
  54215=>"101111111",
  54216=>"100100011",
  54217=>"000000000",
  54218=>"001011110",
  54219=>"100010011",
  54220=>"010101000",
  54221=>"110010000",
  54222=>"000011111",
  54223=>"110101110",
  54224=>"101100010",
  54225=>"100001000",
  54226=>"101101111",
  54227=>"111000000",
  54228=>"010100010",
  54229=>"100000100",
  54230=>"101100001",
  54231=>"000011000",
  54232=>"101001011",
  54233=>"000100101",
  54234=>"101111010",
  54235=>"111001100",
  54236=>"011000111",
  54237=>"101000000",
  54238=>"000101101",
  54239=>"010000010",
  54240=>"100110101",
  54241=>"011110110",
  54242=>"101110101",
  54243=>"110001000",
  54244=>"010010001",
  54245=>"100010101",
  54246=>"000111000",
  54247=>"100000110",
  54248=>"001000101",
  54249=>"100100100",
  54250=>"000001110",
  54251=>"011110111",
  54252=>"101001010",
  54253=>"000101111",
  54254=>"111100110",
  54255=>"101010000",
  54256=>"001011000",
  54257=>"100111001",
  54258=>"001101111",
  54259=>"101001001",
  54260=>"010010000",
  54261=>"010101111",
  54262=>"000101001",
  54263=>"000111010",
  54264=>"100100100",
  54265=>"111001111",
  54266=>"000001000",
  54267=>"010110010",
  54268=>"001100001",
  54269=>"000001001",
  54270=>"110011011",
  54271=>"100110011",
  54272=>"101001000",
  54273=>"011010010",
  54274=>"010100111",
  54275=>"001111110",
  54276=>"101110011",
  54277=>"001000101",
  54278=>"111101010",
  54279=>"000011100",
  54280=>"000000111",
  54281=>"001001111",
  54282=>"111011000",
  54283=>"100000011",
  54284=>"100010010",
  54285=>"011100000",
  54286=>"000000111",
  54287=>"010100000",
  54288=>"110111010",
  54289=>"011111110",
  54290=>"001111000",
  54291=>"111000101",
  54292=>"101101110",
  54293=>"011000100",
  54294=>"101110101",
  54295=>"111101000",
  54296=>"110010000",
  54297=>"110010100",
  54298=>"001110111",
  54299=>"101111101",
  54300=>"011011110",
  54301=>"111011111",
  54302=>"110000010",
  54303=>"110111001",
  54304=>"011011110",
  54305=>"110001000",
  54306=>"101101000",
  54307=>"010011110",
  54308=>"011111011",
  54309=>"010010001",
  54310=>"010101000",
  54311=>"000011000",
  54312=>"111111101",
  54313=>"001011010",
  54314=>"110011011",
  54315=>"110011101",
  54316=>"100011010",
  54317=>"111111011",
  54318=>"111111111",
  54319=>"111001000",
  54320=>"111001100",
  54321=>"110011101",
  54322=>"101111101",
  54323=>"000001000",
  54324=>"111000001",
  54325=>"001000101",
  54326=>"000001001",
  54327=>"101101100",
  54328=>"011101100",
  54329=>"010100000",
  54330=>"100101100",
  54331=>"111111111",
  54332=>"010111111",
  54333=>"100111011",
  54334=>"001010110",
  54335=>"110001011",
  54336=>"010010010",
  54337=>"110110100",
  54338=>"010001001",
  54339=>"010000001",
  54340=>"100001001",
  54341=>"110000011",
  54342=>"000110110",
  54343=>"100001010",
  54344=>"001101001",
  54345=>"111001101",
  54346=>"111111000",
  54347=>"000000110",
  54348=>"001000100",
  54349=>"001000100",
  54350=>"110011011",
  54351=>"111100010",
  54352=>"011100001",
  54353=>"111101010",
  54354=>"010011010",
  54355=>"011000010",
  54356=>"100000101",
  54357=>"100010010",
  54358=>"011001111",
  54359=>"100111011",
  54360=>"011010011",
  54361=>"111111000",
  54362=>"100000000",
  54363=>"100111111",
  54364=>"001111001",
  54365=>"000001111",
  54366=>"001011001",
  54367=>"000001000",
  54368=>"111110011",
  54369=>"100000010",
  54370=>"111110001",
  54371=>"111111000",
  54372=>"011010000",
  54373=>"001000010",
  54374=>"011110110",
  54375=>"001111010",
  54376=>"000100101",
  54377=>"010100100",
  54378=>"011011110",
  54379=>"001011101",
  54380=>"000110010",
  54381=>"101000110",
  54382=>"001111100",
  54383=>"111000011",
  54384=>"101001100",
  54385=>"101011100",
  54386=>"111001111",
  54387=>"000011011",
  54388=>"100100101",
  54389=>"011111001",
  54390=>"000110010",
  54391=>"101110110",
  54392=>"010110110",
  54393=>"001000111",
  54394=>"001000011",
  54395=>"011010111",
  54396=>"000011101",
  54397=>"011001101",
  54398=>"101100010",
  54399=>"110101010",
  54400=>"100110110",
  54401=>"111111110",
  54402=>"100011010",
  54403=>"111111001",
  54404=>"100110001",
  54405=>"010000010",
  54406=>"110101001",
  54407=>"001011010",
  54408=>"011000101",
  54409=>"011100111",
  54410=>"111010001",
  54411=>"000110000",
  54412=>"111110001",
  54413=>"100001001",
  54414=>"001000110",
  54415=>"000100110",
  54416=>"111100010",
  54417=>"000101100",
  54418=>"001000100",
  54419=>"011010111",
  54420=>"101001100",
  54421=>"010000001",
  54422=>"110111101",
  54423=>"101101001",
  54424=>"110011001",
  54425=>"100111110",
  54426=>"001000110",
  54427=>"010011001",
  54428=>"000001011",
  54429=>"100110111",
  54430=>"110000011",
  54431=>"001000100",
  54432=>"101001101",
  54433=>"001000010",
  54434=>"010000111",
  54435=>"101110101",
  54436=>"100011111",
  54437=>"011100101",
  54438=>"100011011",
  54439=>"011001010",
  54440=>"101111101",
  54441=>"110010101",
  54442=>"111010011",
  54443=>"100000101",
  54444=>"011011000",
  54445=>"000010000",
  54446=>"100001001",
  54447=>"000001111",
  54448=>"011000000",
  54449=>"110001001",
  54450=>"101111110",
  54451=>"101011001",
  54452=>"110101101",
  54453=>"010100101",
  54454=>"101100101",
  54455=>"010001111",
  54456=>"100110001",
  54457=>"100111000",
  54458=>"001010011",
  54459=>"110101111",
  54460=>"101010001",
  54461=>"010110101",
  54462=>"011100001",
  54463=>"110000010",
  54464=>"010101001",
  54465=>"010000000",
  54466=>"111110111",
  54467=>"100010000",
  54468=>"100110111",
  54469=>"000111000",
  54470=>"000010011",
  54471=>"010110010",
  54472=>"000110000",
  54473=>"100110011",
  54474=>"000000000",
  54475=>"101100001",
  54476=>"010001100",
  54477=>"100110111",
  54478=>"010010101",
  54479=>"100111000",
  54480=>"111011010",
  54481=>"111111110",
  54482=>"100101000",
  54483=>"110100001",
  54484=>"110001001",
  54485=>"110011010",
  54486=>"011000100",
  54487=>"111010111",
  54488=>"101001101",
  54489=>"100011100",
  54490=>"001001010",
  54491=>"110101011",
  54492=>"011100100",
  54493=>"101001110",
  54494=>"000101010",
  54495=>"001110001",
  54496=>"001111000",
  54497=>"111001011",
  54498=>"011010111",
  54499=>"111100110",
  54500=>"010010011",
  54501=>"101101000",
  54502=>"111111111",
  54503=>"010011001",
  54504=>"111101101",
  54505=>"100111110",
  54506=>"011111010",
  54507=>"101110011",
  54508=>"100100001",
  54509=>"011100111",
  54510=>"011111101",
  54511=>"101000110",
  54512=>"000100110",
  54513=>"100011001",
  54514=>"001100111",
  54515=>"100000100",
  54516=>"110011000",
  54517=>"000110110",
  54518=>"101000101",
  54519=>"001101001",
  54520=>"111010101",
  54521=>"111111111",
  54522=>"100010000",
  54523=>"011100111",
  54524=>"000011111",
  54525=>"100101010",
  54526=>"010101100",
  54527=>"001100001",
  54528=>"101011100",
  54529=>"000010111",
  54530=>"001101100",
  54531=>"010100110",
  54532=>"010011000",
  54533=>"110101001",
  54534=>"010001101",
  54535=>"010001111",
  54536=>"011100111",
  54537=>"011111001",
  54538=>"111001001",
  54539=>"010000010",
  54540=>"111110000",
  54541=>"010000010",
  54542=>"101001111",
  54543=>"111010101",
  54544=>"000010110",
  54545=>"110000111",
  54546=>"111000100",
  54547=>"100101011",
  54548=>"000000000",
  54549=>"110101101",
  54550=>"000010000",
  54551=>"011100010",
  54552=>"011110000",
  54553=>"101101111",
  54554=>"000000001",
  54555=>"000100001",
  54556=>"110000011",
  54557=>"111111101",
  54558=>"111100000",
  54559=>"101100110",
  54560=>"010110010",
  54561=>"000000011",
  54562=>"111101111",
  54563=>"110010111",
  54564=>"000000111",
  54565=>"101101001",
  54566=>"111111000",
  54567=>"000011110",
  54568=>"000100001",
  54569=>"001000101",
  54570=>"000000011",
  54571=>"011010011",
  54572=>"111000101",
  54573=>"000011010",
  54574=>"111111111",
  54575=>"110010010",
  54576=>"111011110",
  54577=>"010110101",
  54578=>"110000011",
  54579=>"101010110",
  54580=>"110100001",
  54581=>"111011010",
  54582=>"001000101",
  54583=>"101010111",
  54584=>"111101000",
  54585=>"100000100",
  54586=>"111100000",
  54587=>"111010011",
  54588=>"000001111",
  54589=>"101000000",
  54590=>"011111100",
  54591=>"111110111",
  54592=>"000111100",
  54593=>"101000001",
  54594=>"101010100",
  54595=>"011000100",
  54596=>"110111000",
  54597=>"111001001",
  54598=>"100110110",
  54599=>"110100010",
  54600=>"100111100",
  54601=>"110001000",
  54602=>"100111011",
  54603=>"001110010",
  54604=>"101110001",
  54605=>"000010100",
  54606=>"110110101",
  54607=>"101011111",
  54608=>"101110111",
  54609=>"110100101",
  54610=>"010100010",
  54611=>"000001100",
  54612=>"110101100",
  54613=>"101000101",
  54614=>"011110011",
  54615=>"111010001",
  54616=>"110011101",
  54617=>"000101101",
  54618=>"110110011",
  54619=>"111011101",
  54620=>"010010011",
  54621=>"010101010",
  54622=>"000010110",
  54623=>"110011010",
  54624=>"000000000",
  54625=>"000110000",
  54626=>"001110101",
  54627=>"111110001",
  54628=>"010001000",
  54629=>"000010000",
  54630=>"011010000",
  54631=>"000100010",
  54632=>"100000010",
  54633=>"100011110",
  54634=>"110111011",
  54635=>"111110101",
  54636=>"111101010",
  54637=>"111101011",
  54638=>"100100111",
  54639=>"111000111",
  54640=>"000001000",
  54641=>"101100000",
  54642=>"010011111",
  54643=>"011011101",
  54644=>"001100111",
  54645=>"111011010",
  54646=>"110100000",
  54647=>"010000010",
  54648=>"000110100",
  54649=>"000111100",
  54650=>"011011101",
  54651=>"001000000",
  54652=>"000010010",
  54653=>"101110011",
  54654=>"100110001",
  54655=>"000001110",
  54656=>"111101011",
  54657=>"010011000",
  54658=>"110011110",
  54659=>"011011001",
  54660=>"011111100",
  54661=>"011001111",
  54662=>"100100111",
  54663=>"000011101",
  54664=>"000011011",
  54665=>"001101001",
  54666=>"010101001",
  54667=>"100000100",
  54668=>"000000100",
  54669=>"000110010",
  54670=>"111111100",
  54671=>"100110101",
  54672=>"111000101",
  54673=>"101000101",
  54674=>"101110101",
  54675=>"000100101",
  54676=>"011010111",
  54677=>"111101010",
  54678=>"000110000",
  54679=>"010111100",
  54680=>"111100011",
  54681=>"001101001",
  54682=>"110110110",
  54683=>"110011000",
  54684=>"010010001",
  54685=>"000100001",
  54686=>"111100111",
  54687=>"111000000",
  54688=>"110011111",
  54689=>"001000000",
  54690=>"101111000",
  54691=>"110100000",
  54692=>"101111110",
  54693=>"000101111",
  54694=>"011110000",
  54695=>"111111100",
  54696=>"100010100",
  54697=>"000101000",
  54698=>"110000100",
  54699=>"000110110",
  54700=>"111001011",
  54701=>"101000101",
  54702=>"000000100",
  54703=>"011011101",
  54704=>"111100010",
  54705=>"111111110",
  54706=>"000010000",
  54707=>"010110000",
  54708=>"101001110",
  54709=>"111000001",
  54710=>"111111000",
  54711=>"101110110",
  54712=>"010011010",
  54713=>"001000001",
  54714=>"100011110",
  54715=>"100000001",
  54716=>"000010100",
  54717=>"000001110",
  54718=>"001000100",
  54719=>"111001111",
  54720=>"011010000",
  54721=>"011000001",
  54722=>"100100010",
  54723=>"000011011",
  54724=>"111111111",
  54725=>"100111111",
  54726=>"111001000",
  54727=>"000111100",
  54728=>"110011000",
  54729=>"001101001",
  54730=>"110101101",
  54731=>"111100100",
  54732=>"010110000",
  54733=>"011011001",
  54734=>"011001001",
  54735=>"111100010",
  54736=>"001110100",
  54737=>"011010001",
  54738=>"111001001",
  54739=>"001100100",
  54740=>"111001100",
  54741=>"100011000",
  54742=>"010100111",
  54743=>"001101000",
  54744=>"111111001",
  54745=>"010011010",
  54746=>"010110101",
  54747=>"000100011",
  54748=>"001001100",
  54749=>"100111011",
  54750=>"101010010",
  54751=>"010000111",
  54752=>"001110110",
  54753=>"111001110",
  54754=>"101111010",
  54755=>"010111001",
  54756=>"100110010",
  54757=>"010100111",
  54758=>"001010010",
  54759=>"101110010",
  54760=>"001101000",
  54761=>"111010100",
  54762=>"001000011",
  54763=>"011001000",
  54764=>"000001101",
  54765=>"001011000",
  54766=>"001010101",
  54767=>"010101001",
  54768=>"100111110",
  54769=>"000001000",
  54770=>"101011111",
  54771=>"110011101",
  54772=>"011101000",
  54773=>"111101000",
  54774=>"110011111",
  54775=>"101111101",
  54776=>"000000110",
  54777=>"101010011",
  54778=>"001101010",
  54779=>"010010111",
  54780=>"001100001",
  54781=>"111100010",
  54782=>"000111111",
  54783=>"001010101",
  54784=>"101101011",
  54785=>"101100110",
  54786=>"110011011",
  54787=>"010100111",
  54788=>"100011011",
  54789=>"001110110",
  54790=>"011000011",
  54791=>"101111001",
  54792=>"101110011",
  54793=>"111111110",
  54794=>"101001111",
  54795=>"100000011",
  54796=>"100001001",
  54797=>"100011011",
  54798=>"011101110",
  54799=>"110111011",
  54800=>"101001100",
  54801=>"110011010",
  54802=>"011001100",
  54803=>"100000010",
  54804=>"000110101",
  54805=>"111100000",
  54806=>"010111111",
  54807=>"010110010",
  54808=>"111000001",
  54809=>"110010101",
  54810=>"000011011",
  54811=>"100111001",
  54812=>"101110100",
  54813=>"010001100",
  54814=>"100010010",
  54815=>"010101110",
  54816=>"000011001",
  54817=>"000111001",
  54818=>"000001101",
  54819=>"010011100",
  54820=>"111011111",
  54821=>"111111100",
  54822=>"011110000",
  54823=>"111000110",
  54824=>"000000011",
  54825=>"111111111",
  54826=>"010110010",
  54827=>"100011110",
  54828=>"011100110",
  54829=>"111011010",
  54830=>"010111001",
  54831=>"110111111",
  54832=>"001010100",
  54833=>"000110101",
  54834=>"001101011",
  54835=>"110111111",
  54836=>"011001110",
  54837=>"111110110",
  54838=>"010011111",
  54839=>"000000101",
  54840=>"111010010",
  54841=>"001000110",
  54842=>"100001010",
  54843=>"101001100",
  54844=>"101101100",
  54845=>"010000111",
  54846=>"100001001",
  54847=>"111010111",
  54848=>"111010101",
  54849=>"111011010",
  54850=>"101101001",
  54851=>"100011000",
  54852=>"110100001",
  54853=>"011110100",
  54854=>"010001011",
  54855=>"111001011",
  54856=>"100110001",
  54857=>"000011110",
  54858=>"111000100",
  54859=>"110011100",
  54860=>"001011001",
  54861=>"000010011",
  54862=>"110100101",
  54863=>"000011000",
  54864=>"011101110",
  54865=>"111010000",
  54866=>"100110101",
  54867=>"001100011",
  54868=>"110100111",
  54869=>"000101110",
  54870=>"100011000",
  54871=>"000110010",
  54872=>"000000000",
  54873=>"110000110",
  54874=>"110001101",
  54875=>"110111010",
  54876=>"110010001",
  54877=>"111010111",
  54878=>"100011110",
  54879=>"111001101",
  54880=>"101101011",
  54881=>"010000111",
  54882=>"000101110",
  54883=>"100001010",
  54884=>"101110001",
  54885=>"000011010",
  54886=>"001100111",
  54887=>"000110001",
  54888=>"111111000",
  54889=>"111001111",
  54890=>"001000101",
  54891=>"111110101",
  54892=>"110001011",
  54893=>"100010000",
  54894=>"010100001",
  54895=>"000000011",
  54896=>"110101110",
  54897=>"000001001",
  54898=>"111100101",
  54899=>"110101000",
  54900=>"001101010",
  54901=>"101001001",
  54902=>"111111111",
  54903=>"111111110",
  54904=>"011100110",
  54905=>"011001111",
  54906=>"011001100",
  54907=>"011110110",
  54908=>"111101001",
  54909=>"111000001",
  54910=>"101011111",
  54911=>"101011011",
  54912=>"011110000",
  54913=>"110001011",
  54914=>"110011010",
  54915=>"101001011",
  54916=>"111101111",
  54917=>"001010011",
  54918=>"101011111",
  54919=>"100010010",
  54920=>"100110011",
  54921=>"101101001",
  54922=>"100111001",
  54923=>"000110110",
  54924=>"111101100",
  54925=>"101001111",
  54926=>"011011001",
  54927=>"110010101",
  54928=>"111110110",
  54929=>"000101011",
  54930=>"000000001",
  54931=>"100010011",
  54932=>"100100111",
  54933=>"101111111",
  54934=>"101111111",
  54935=>"100000101",
  54936=>"011011101",
  54937=>"010001010",
  54938=>"010111001",
  54939=>"100110001",
  54940=>"011100001",
  54941=>"001110100",
  54942=>"001000110",
  54943=>"100100000",
  54944=>"100001000",
  54945=>"101010011",
  54946=>"001001110",
  54947=>"100001110",
  54948=>"111111101",
  54949=>"101010011",
  54950=>"111001000",
  54951=>"011101000",
  54952=>"101100010",
  54953=>"100110010",
  54954=>"000000101",
  54955=>"101011000",
  54956=>"110000101",
  54957=>"101010001",
  54958=>"000110110",
  54959=>"100101100",
  54960=>"100101101",
  54961=>"011001000",
  54962=>"000011101",
  54963=>"100100000",
  54964=>"110000000",
  54965=>"001111000",
  54966=>"111100100",
  54967=>"000000011",
  54968=>"001110010",
  54969=>"110010110",
  54970=>"101011100",
  54971=>"000000000",
  54972=>"111101100",
  54973=>"010100010",
  54974=>"010010001",
  54975=>"110111100",
  54976=>"001110100",
  54977=>"000011001",
  54978=>"111101101",
  54979=>"111110001",
  54980=>"011110001",
  54981=>"101000011",
  54982=>"111111101",
  54983=>"110111111",
  54984=>"111100100",
  54985=>"110011101",
  54986=>"011000000",
  54987=>"110111000",
  54988=>"101001000",
  54989=>"001101101",
  54990=>"001000011",
  54991=>"000110001",
  54992=>"101000000",
  54993=>"011010000",
  54994=>"100001111",
  54995=>"101001001",
  54996=>"000010000",
  54997=>"001101000",
  54998=>"100010100",
  54999=>"110011100",
  55000=>"111000110",
  55001=>"001111101",
  55002=>"011111010",
  55003=>"101000001",
  55004=>"011101101",
  55005=>"010000100",
  55006=>"001110100",
  55007=>"101111001",
  55008=>"110000100",
  55009=>"000001001",
  55010=>"111111101",
  55011=>"001001001",
  55012=>"000101010",
  55013=>"100011100",
  55014=>"100011111",
  55015=>"011100011",
  55016=>"011001110",
  55017=>"111110011",
  55018=>"110111111",
  55019=>"101000100",
  55020=>"110000000",
  55021=>"000101111",
  55022=>"100100001",
  55023=>"000001000",
  55024=>"000111100",
  55025=>"000110000",
  55026=>"011000001",
  55027=>"011010101",
  55028=>"110000011",
  55029=>"100010010",
  55030=>"101001010",
  55031=>"001001011",
  55032=>"011011101",
  55033=>"111011111",
  55034=>"101110100",
  55035=>"111001010",
  55036=>"011110010",
  55037=>"100110011",
  55038=>"001110101",
  55039=>"010011110",
  55040=>"100101110",
  55041=>"100101111",
  55042=>"000011101",
  55043=>"110011100",
  55044=>"100110011",
  55045=>"000101011",
  55046=>"110111111",
  55047=>"000110010",
  55048=>"101000101",
  55049=>"101000011",
  55050=>"011111110",
  55051=>"000010111",
  55052=>"001100010",
  55053=>"001011111",
  55054=>"000100001",
  55055=>"100100101",
  55056=>"110111110",
  55057=>"011101110",
  55058=>"000001000",
  55059=>"101000100",
  55060=>"111110000",
  55061=>"110010111",
  55062=>"100010110",
  55063=>"010110100",
  55064=>"100100101",
  55065=>"001011100",
  55066=>"100001001",
  55067=>"010101010",
  55068=>"000001101",
  55069=>"111111000",
  55070=>"010100001",
  55071=>"110101010",
  55072=>"001001101",
  55073=>"101000101",
  55074=>"100001111",
  55075=>"111101000",
  55076=>"110010101",
  55077=>"111001011",
  55078=>"011010111",
  55079=>"100101110",
  55080=>"011110101",
  55081=>"000010011",
  55082=>"001110000",
  55083=>"100001111",
  55084=>"001001110",
  55085=>"000010010",
  55086=>"100100011",
  55087=>"100010011",
  55088=>"100101011",
  55089=>"101010110",
  55090=>"010111010",
  55091=>"000010010",
  55092=>"010011010",
  55093=>"001011010",
  55094=>"000100110",
  55095=>"001101110",
  55096=>"010111011",
  55097=>"000010000",
  55098=>"011101000",
  55099=>"001110101",
  55100=>"111010111",
  55101=>"001111111",
  55102=>"011000010",
  55103=>"001000011",
  55104=>"000110100",
  55105=>"000110100",
  55106=>"110011100",
  55107=>"111010110",
  55108=>"011010110",
  55109=>"001110111",
  55110=>"110011001",
  55111=>"110100000",
  55112=>"001000011",
  55113=>"011000011",
  55114=>"011100011",
  55115=>"101101110",
  55116=>"111001100",
  55117=>"000111110",
  55118=>"000110010",
  55119=>"100000000",
  55120=>"011011001",
  55121=>"010010000",
  55122=>"001101000",
  55123=>"111110001",
  55124=>"100110100",
  55125=>"101101101",
  55126=>"101110011",
  55127=>"011010000",
  55128=>"111011011",
  55129=>"101011001",
  55130=>"000010011",
  55131=>"110101101",
  55132=>"000101010",
  55133=>"111001100",
  55134=>"110001110",
  55135=>"100001010",
  55136=>"111001101",
  55137=>"111110100",
  55138=>"110100000",
  55139=>"011010111",
  55140=>"001010111",
  55141=>"110001010",
  55142=>"010010110",
  55143=>"111000100",
  55144=>"000001000",
  55145=>"001001000",
  55146=>"110110100",
  55147=>"001000110",
  55148=>"001111100",
  55149=>"100010000",
  55150=>"001111011",
  55151=>"011011011",
  55152=>"011000101",
  55153=>"011010111",
  55154=>"011010101",
  55155=>"111000010",
  55156=>"000101111",
  55157=>"000000110",
  55158=>"001001111",
  55159=>"010101001",
  55160=>"001111000",
  55161=>"001001000",
  55162=>"001001110",
  55163=>"111001111",
  55164=>"000000001",
  55165=>"000011110",
  55166=>"001101001",
  55167=>"101010001",
  55168=>"001011010",
  55169=>"010000001",
  55170=>"010000110",
  55171=>"000101000",
  55172=>"110101000",
  55173=>"010010010",
  55174=>"110110010",
  55175=>"001011111",
  55176=>"010101000",
  55177=>"010100111",
  55178=>"110000010",
  55179=>"011101000",
  55180=>"101110100",
  55181=>"101101101",
  55182=>"110110110",
  55183=>"111111100",
  55184=>"001011101",
  55185=>"100010101",
  55186=>"001101101",
  55187=>"111111111",
  55188=>"000000000",
  55189=>"101110000",
  55190=>"110001000",
  55191=>"010001010",
  55192=>"100111000",
  55193=>"010111100",
  55194=>"100010101",
  55195=>"000000110",
  55196=>"111110101",
  55197=>"111000100",
  55198=>"100001000",
  55199=>"100110001",
  55200=>"010000100",
  55201=>"010111011",
  55202=>"100010011",
  55203=>"001001110",
  55204=>"110000011",
  55205=>"111110111",
  55206=>"111101010",
  55207=>"000010100",
  55208=>"001000100",
  55209=>"111101111",
  55210=>"101001011",
  55211=>"010011001",
  55212=>"000100100",
  55213=>"010010111",
  55214=>"111100110",
  55215=>"010111111",
  55216=>"000111111",
  55217=>"110110000",
  55218=>"101101101",
  55219=>"000001011",
  55220=>"000100101",
  55221=>"111000011",
  55222=>"101111001",
  55223=>"101011110",
  55224=>"100001011",
  55225=>"011110001",
  55226=>"100101000",
  55227=>"001001100",
  55228=>"111110100",
  55229=>"111101111",
  55230=>"000101000",
  55231=>"010110010",
  55232=>"110111110",
  55233=>"000010010",
  55234=>"101101110",
  55235=>"001000010",
  55236=>"001010110",
  55237=>"111111100",
  55238=>"010010101",
  55239=>"111111000",
  55240=>"010100001",
  55241=>"001001101",
  55242=>"001100010",
  55243=>"001010100",
  55244=>"111111100",
  55245=>"011011011",
  55246=>"110010100",
  55247=>"110011011",
  55248=>"101111100",
  55249=>"111001001",
  55250=>"111011111",
  55251=>"010000110",
  55252=>"101110101",
  55253=>"110010011",
  55254=>"100110110",
  55255=>"010000000",
  55256=>"110100111",
  55257=>"001100011",
  55258=>"101000011",
  55259=>"001111110",
  55260=>"110110010",
  55261=>"101010111",
  55262=>"000000000",
  55263=>"100011011",
  55264=>"101011110",
  55265=>"011000100",
  55266=>"010100110",
  55267=>"101011100",
  55268=>"010100001",
  55269=>"100011111",
  55270=>"101101001",
  55271=>"001001101",
  55272=>"010101100",
  55273=>"011000000",
  55274=>"111111000",
  55275=>"001000100",
  55276=>"001100010",
  55277=>"110110001",
  55278=>"100101010",
  55279=>"010100011",
  55280=>"101110010",
  55281=>"000011101",
  55282=>"000010000",
  55283=>"110101000",
  55284=>"000101010",
  55285=>"000100010",
  55286=>"101110001",
  55287=>"101110000",
  55288=>"110010111",
  55289=>"101111111",
  55290=>"110001000",
  55291=>"011111100",
  55292=>"100010110",
  55293=>"101011000",
  55294=>"101010001",
  55295=>"110101011",
  55296=>"010000010",
  55297=>"100001100",
  55298=>"000011010",
  55299=>"111000011",
  55300=>"110100000",
  55301=>"001000100",
  55302=>"010111110",
  55303=>"101010011",
  55304=>"100101111",
  55305=>"100110111",
  55306=>"101101011",
  55307=>"100011001",
  55308=>"110101011",
  55309=>"011010100",
  55310=>"110010010",
  55311=>"001100000",
  55312=>"100010011",
  55313=>"001110010",
  55314=>"001100001",
  55315=>"101001010",
  55316=>"010000100",
  55317=>"010010011",
  55318=>"001110111",
  55319=>"001111000",
  55320=>"010101101",
  55321=>"101011010",
  55322=>"001011011",
  55323=>"110100000",
  55324=>"001100011",
  55325=>"011001011",
  55326=>"010100001",
  55327=>"100001100",
  55328=>"110111000",
  55329=>"001000101",
  55330=>"101000100",
  55331=>"110111101",
  55332=>"111110111",
  55333=>"001000100",
  55334=>"010000111",
  55335=>"010001111",
  55336=>"000111111",
  55337=>"000001110",
  55338=>"100111100",
  55339=>"010100010",
  55340=>"001010011",
  55341=>"011010001",
  55342=>"000000100",
  55343=>"110111110",
  55344=>"110111001",
  55345=>"011000000",
  55346=>"011010011",
  55347=>"001000111",
  55348=>"001011001",
  55349=>"010111011",
  55350=>"101010000",
  55351=>"110100101",
  55352=>"001100100",
  55353=>"101010001",
  55354=>"001111101",
  55355=>"111110101",
  55356=>"011110000",
  55357=>"101111000",
  55358=>"100001010",
  55359=>"111111100",
  55360=>"110001001",
  55361=>"001101100",
  55362=>"111000100",
  55363=>"000000110",
  55364=>"101010011",
  55365=>"001001000",
  55366=>"110101000",
  55367=>"111000101",
  55368=>"010111110",
  55369=>"010000100",
  55370=>"111000000",
  55371=>"011110011",
  55372=>"000010001",
  55373=>"000101000",
  55374=>"000000100",
  55375=>"011110100",
  55376=>"110101010",
  55377=>"001001110",
  55378=>"011110100",
  55379=>"000000110",
  55380=>"100100001",
  55381=>"110001100",
  55382=>"000000110",
  55383=>"110000001",
  55384=>"100000001",
  55385=>"000100111",
  55386=>"001000011",
  55387=>"101110100",
  55388=>"011011001",
  55389=>"001000100",
  55390=>"010011000",
  55391=>"001000101",
  55392=>"010001101",
  55393=>"100000110",
  55394=>"111011100",
  55395=>"000100010",
  55396=>"111111000",
  55397=>"101110010",
  55398=>"111111010",
  55399=>"111111110",
  55400=>"000010001",
  55401=>"111100001",
  55402=>"000000010",
  55403=>"110010010",
  55404=>"111000101",
  55405=>"011011000",
  55406=>"000000010",
  55407=>"100110001",
  55408=>"001101000",
  55409=>"011010100",
  55410=>"011011011",
  55411=>"111001100",
  55412=>"011100110",
  55413=>"001001000",
  55414=>"111101101",
  55415=>"000101001",
  55416=>"100101001",
  55417=>"001001001",
  55418=>"010110101",
  55419=>"111011100",
  55420=>"001101100",
  55421=>"100001001",
  55422=>"100001000",
  55423=>"001011110",
  55424=>"100011000",
  55425=>"011111101",
  55426=>"000001000",
  55427=>"110110000",
  55428=>"001001001",
  55429=>"000100010",
  55430=>"001111110",
  55431=>"011101000",
  55432=>"000001000",
  55433=>"010000000",
  55434=>"011001011",
  55435=>"010010111",
  55436=>"111100101",
  55437=>"011100010",
  55438=>"110001000",
  55439=>"100110010",
  55440=>"111001111",
  55441=>"010010010",
  55442=>"001100011",
  55443=>"001111101",
  55444=>"101111111",
  55445=>"111011111",
  55446=>"111111111",
  55447=>"111011000",
  55448=>"111110010",
  55449=>"111010000",
  55450=>"011111101",
  55451=>"001101010",
  55452=>"000111000",
  55453=>"111011011",
  55454=>"101010000",
  55455=>"101010111",
  55456=>"010111011",
  55457=>"010111000",
  55458=>"010001010",
  55459=>"101111100",
  55460=>"110010111",
  55461=>"010001110",
  55462=>"000111100",
  55463=>"001111001",
  55464=>"110000110",
  55465=>"110110111",
  55466=>"101111111",
  55467=>"011101011",
  55468=>"011010110",
  55469=>"011100100",
  55470=>"011111110",
  55471=>"011011101",
  55472=>"100101111",
  55473=>"100111111",
  55474=>"001010010",
  55475=>"101000000",
  55476=>"111100100",
  55477=>"111000111",
  55478=>"011001110",
  55479=>"010011010",
  55480=>"011101011",
  55481=>"000000101",
  55482=>"100101001",
  55483=>"110010000",
  55484=>"111100101",
  55485=>"000100100",
  55486=>"101100111",
  55487=>"111010000",
  55488=>"100000111",
  55489=>"011101111",
  55490=>"111110001",
  55491=>"001011001",
  55492=>"011000111",
  55493=>"001100110",
  55494=>"000111100",
  55495=>"100110010",
  55496=>"000010100",
  55497=>"010001111",
  55498=>"011001111",
  55499=>"100011010",
  55500=>"010010000",
  55501=>"010000100",
  55502=>"100110111",
  55503=>"011000101",
  55504=>"011101001",
  55505=>"000011101",
  55506=>"011000001",
  55507=>"001111101",
  55508=>"100000110",
  55509=>"000010100",
  55510=>"101001000",
  55511=>"000011101",
  55512=>"010100000",
  55513=>"001001100",
  55514=>"100001110",
  55515=>"001011111",
  55516=>"011111001",
  55517=>"101001100",
  55518=>"101010100",
  55519=>"011100100",
  55520=>"111111011",
  55521=>"010010010",
  55522=>"010001011",
  55523=>"010100001",
  55524=>"011110011",
  55525=>"011110110",
  55526=>"100001000",
  55527=>"010011110",
  55528=>"011001110",
  55529=>"100010001",
  55530=>"000010111",
  55531=>"101011011",
  55532=>"100101001",
  55533=>"010000010",
  55534=>"011000011",
  55535=>"110001100",
  55536=>"101011011",
  55537=>"100110100",
  55538=>"000100010",
  55539=>"110101111",
  55540=>"110011001",
  55541=>"000101001",
  55542=>"011100000",
  55543=>"110011101",
  55544=>"100100101",
  55545=>"111101111",
  55546=>"010111100",
  55547=>"001001010",
  55548=>"010000110",
  55549=>"111111100",
  55550=>"101011110",
  55551=>"111111110",
  55552=>"111111101",
  55553=>"101010001",
  55554=>"110011001",
  55555=>"111101101",
  55556=>"001010001",
  55557=>"001101001",
  55558=>"101001000",
  55559=>"010111111",
  55560=>"111001110",
  55561=>"000011111",
  55562=>"101101000",
  55563=>"100000010",
  55564=>"000010000",
  55565=>"011101110",
  55566=>"000101100",
  55567=>"111010011",
  55568=>"010110010",
  55569=>"000110110",
  55570=>"111001000",
  55571=>"000011110",
  55572=>"101010000",
  55573=>"100011001",
  55574=>"000100100",
  55575=>"001010011",
  55576=>"001111001",
  55577=>"001011000",
  55578=>"111011001",
  55579=>"000111111",
  55580=>"010011100",
  55581=>"100000101",
  55582=>"100011100",
  55583=>"000001011",
  55584=>"101111011",
  55585=>"001100010",
  55586=>"111011010",
  55587=>"010111110",
  55588=>"011110100",
  55589=>"110001111",
  55590=>"110010010",
  55591=>"011000111",
  55592=>"010100011",
  55593=>"110101011",
  55594=>"101111111",
  55595=>"010111000",
  55596=>"111000001",
  55597=>"101101110",
  55598=>"001011111",
  55599=>"100111110",
  55600=>"100100000",
  55601=>"001010000",
  55602=>"111001001",
  55603=>"010011000",
  55604=>"111000100",
  55605=>"011000111",
  55606=>"100001000",
  55607=>"111111011",
  55608=>"010111011",
  55609=>"010011001",
  55610=>"100010011",
  55611=>"110000100",
  55612=>"110010111",
  55613=>"010010100",
  55614=>"101011011",
  55615=>"110101100",
  55616=>"000100110",
  55617=>"000010000",
  55618=>"001010011",
  55619=>"110010100",
  55620=>"001000111",
  55621=>"110010000",
  55622=>"101010001",
  55623=>"000100110",
  55624=>"100101101",
  55625=>"001010000",
  55626=>"100011011",
  55627=>"001101111",
  55628=>"110101111",
  55629=>"101111000",
  55630=>"000010110",
  55631=>"110011100",
  55632=>"111011111",
  55633=>"101000000",
  55634=>"111100111",
  55635=>"101101111",
  55636=>"100001011",
  55637=>"000000011",
  55638=>"110011011",
  55639=>"100111000",
  55640=>"101110110",
  55641=>"110000100",
  55642=>"011011001",
  55643=>"001000011",
  55644=>"010110001",
  55645=>"010001000",
  55646=>"010110111",
  55647=>"000101000",
  55648=>"000010101",
  55649=>"010111011",
  55650=>"001011000",
  55651=>"001011001",
  55652=>"010001000",
  55653=>"000111111",
  55654=>"101110000",
  55655=>"001111110",
  55656=>"110000000",
  55657=>"110101100",
  55658=>"011110011",
  55659=>"110111111",
  55660=>"010000101",
  55661=>"100111000",
  55662=>"000001110",
  55663=>"011101110",
  55664=>"010100110",
  55665=>"000111101",
  55666=>"111001001",
  55667=>"111010011",
  55668=>"000011111",
  55669=>"001101111",
  55670=>"011010110",
  55671=>"001101001",
  55672=>"010101010",
  55673=>"011011010",
  55674=>"110100001",
  55675=>"000101001",
  55676=>"011000000",
  55677=>"100010000",
  55678=>"110011010",
  55679=>"011010000",
  55680=>"001101101",
  55681=>"110000110",
  55682=>"111101001",
  55683=>"001110001",
  55684=>"000101000",
  55685=>"001011011",
  55686=>"100110001",
  55687=>"000000000",
  55688=>"101010010",
  55689=>"011110111",
  55690=>"001010011",
  55691=>"111010001",
  55692=>"001000000",
  55693=>"000100100",
  55694=>"111001000",
  55695=>"011010101",
  55696=>"010010011",
  55697=>"101100101",
  55698=>"010000001",
  55699=>"010001001",
  55700=>"011010010",
  55701=>"100110110",
  55702=>"101111111",
  55703=>"100110011",
  55704=>"110011100",
  55705=>"100010111",
  55706=>"111011001",
  55707=>"001010011",
  55708=>"111011111",
  55709=>"011001100",
  55710=>"110010100",
  55711=>"000101110",
  55712=>"110110011",
  55713=>"101101011",
  55714=>"001000000",
  55715=>"010111101",
  55716=>"000101101",
  55717=>"000011101",
  55718=>"110011110",
  55719=>"011011000",
  55720=>"010100001",
  55721=>"101101101",
  55722=>"100001100",
  55723=>"111111011",
  55724=>"100011011",
  55725=>"100000111",
  55726=>"001100000",
  55727=>"000010000",
  55728=>"100001010",
  55729=>"111010000",
  55730=>"110010010",
  55731=>"100111100",
  55732=>"001000000",
  55733=>"000110011",
  55734=>"101111000",
  55735=>"101010000",
  55736=>"001010111",
  55737=>"101100001",
  55738=>"000001000",
  55739=>"001100100",
  55740=>"110010110",
  55741=>"100101011",
  55742=>"011100101",
  55743=>"011001011",
  55744=>"000100110",
  55745=>"000001000",
  55746=>"000110000",
  55747=>"000111001",
  55748=>"101111101",
  55749=>"101100001",
  55750=>"010110110",
  55751=>"011101000",
  55752=>"011110110",
  55753=>"010100011",
  55754=>"101110111",
  55755=>"001001001",
  55756=>"010110011",
  55757=>"000010111",
  55758=>"001010100",
  55759=>"100010100",
  55760=>"111011110",
  55761=>"111101001",
  55762=>"101110000",
  55763=>"010011101",
  55764=>"101110110",
  55765=>"100010000",
  55766=>"111010110",
  55767=>"111001001",
  55768=>"000110001",
  55769=>"100010101",
  55770=>"000000111",
  55771=>"001111001",
  55772=>"010001100",
  55773=>"101000100",
  55774=>"100010000",
  55775=>"010001011",
  55776=>"100000110",
  55777=>"001000111",
  55778=>"111100000",
  55779=>"101010010",
  55780=>"110000001",
  55781=>"010010010",
  55782=>"110010000",
  55783=>"010100100",
  55784=>"000110010",
  55785=>"101111001",
  55786=>"101100111",
  55787=>"111010111",
  55788=>"100111101",
  55789=>"011000110",
  55790=>"010100111",
  55791=>"001011101",
  55792=>"111000000",
  55793=>"010101010",
  55794=>"011011010",
  55795=>"001010100",
  55796=>"110100101",
  55797=>"110101111",
  55798=>"110011101",
  55799=>"110011100",
  55800=>"010100000",
  55801=>"011101010",
  55802=>"101101111",
  55803=>"101011001",
  55804=>"000001001",
  55805=>"000111111",
  55806=>"010101000",
  55807=>"011100011",
  55808=>"000100110",
  55809=>"000111000",
  55810=>"011111111",
  55811=>"011110000",
  55812=>"110001100",
  55813=>"011011010",
  55814=>"100110011",
  55815=>"110010100",
  55816=>"010100111",
  55817=>"011101111",
  55818=>"100110100",
  55819=>"010001100",
  55820=>"110100010",
  55821=>"010110100",
  55822=>"001000111",
  55823=>"110111001",
  55824=>"011110110",
  55825=>"001110001",
  55826=>"111101111",
  55827=>"100101111",
  55828=>"110001110",
  55829=>"001110111",
  55830=>"100101000",
  55831=>"011101011",
  55832=>"100000100",
  55833=>"000011010",
  55834=>"000001000",
  55835=>"101110101",
  55836=>"100110010",
  55837=>"100000000",
  55838=>"101101111",
  55839=>"111100101",
  55840=>"100001000",
  55841=>"000101001",
  55842=>"001110101",
  55843=>"001110010",
  55844=>"110001000",
  55845=>"011001101",
  55846=>"000000001",
  55847=>"001001100",
  55848=>"110000000",
  55849=>"000110110",
  55850=>"110101111",
  55851=>"010010110",
  55852=>"101001010",
  55853=>"100000101",
  55854=>"000011100",
  55855=>"000100000",
  55856=>"010111110",
  55857=>"110001011",
  55858=>"011001111",
  55859=>"000011101",
  55860=>"000110000",
  55861=>"100000000",
  55862=>"010011111",
  55863=>"001111011",
  55864=>"010111001",
  55865=>"010100000",
  55866=>"011100001",
  55867=>"000010000",
  55868=>"000111000",
  55869=>"110110101",
  55870=>"111101011",
  55871=>"011010101",
  55872=>"110111010",
  55873=>"101011101",
  55874=>"100011101",
  55875=>"001101011",
  55876=>"000111111",
  55877=>"000001001",
  55878=>"110010110",
  55879=>"000000100",
  55880=>"001110100",
  55881=>"111000010",
  55882=>"000100110",
  55883=>"000011001",
  55884=>"101000100",
  55885=>"001011100",
  55886=>"001000000",
  55887=>"010111011",
  55888=>"110110111",
  55889=>"001001000",
  55890=>"111001110",
  55891=>"101110111",
  55892=>"101010011",
  55893=>"001011001",
  55894=>"111000100",
  55895=>"110111001",
  55896=>"000110101",
  55897=>"110101101",
  55898=>"101110000",
  55899=>"100011111",
  55900=>"110101100",
  55901=>"111000100",
  55902=>"000101111",
  55903=>"100110011",
  55904=>"101001100",
  55905=>"000000110",
  55906=>"010010000",
  55907=>"110001101",
  55908=>"011010110",
  55909=>"010100101",
  55910=>"010011010",
  55911=>"101100111",
  55912=>"111010100",
  55913=>"100100011",
  55914=>"100000111",
  55915=>"111100111",
  55916=>"100001110",
  55917=>"000000001",
  55918=>"010011101",
  55919=>"100100010",
  55920=>"100110100",
  55921=>"001110010",
  55922=>"100101110",
  55923=>"011000100",
  55924=>"100000100",
  55925=>"001000110",
  55926=>"111100111",
  55927=>"110000111",
  55928=>"101010100",
  55929=>"100010100",
  55930=>"000010001",
  55931=>"001000100",
  55932=>"001001110",
  55933=>"101011011",
  55934=>"101000011",
  55935=>"010111001",
  55936=>"110001011",
  55937=>"101111010",
  55938=>"110001100",
  55939=>"101100111",
  55940=>"110000000",
  55941=>"100011000",
  55942=>"000111000",
  55943=>"111010101",
  55944=>"001100100",
  55945=>"110011110",
  55946=>"010000111",
  55947=>"000111001",
  55948=>"011000010",
  55949=>"000100010",
  55950=>"111111111",
  55951=>"000110101",
  55952=>"001001010",
  55953=>"001110000",
  55954=>"011111010",
  55955=>"101000010",
  55956=>"110100111",
  55957=>"100111111",
  55958=>"010101011",
  55959=>"010000000",
  55960=>"100110010",
  55961=>"001011100",
  55962=>"011001110",
  55963=>"001011101",
  55964=>"011000000",
  55965=>"101101111",
  55966=>"111000011",
  55967=>"000100111",
  55968=>"000100001",
  55969=>"110101110",
  55970=>"110111011",
  55971=>"001011001",
  55972=>"101001100",
  55973=>"010111100",
  55974=>"000011010",
  55975=>"100110101",
  55976=>"011001010",
  55977=>"101010001",
  55978=>"001000101",
  55979=>"011111111",
  55980=>"110001111",
  55981=>"001000110",
  55982=>"100100101",
  55983=>"011110111",
  55984=>"010011100",
  55985=>"010011111",
  55986=>"100110011",
  55987=>"000100110",
  55988=>"100000011",
  55989=>"111100000",
  55990=>"001100001",
  55991=>"010011010",
  55992=>"001000001",
  55993=>"101100111",
  55994=>"101101110",
  55995=>"010101111",
  55996=>"011101111",
  55997=>"001101010",
  55998=>"001011100",
  55999=>"001100101",
  56000=>"100001001",
  56001=>"110010110",
  56002=>"111111011",
  56003=>"110000100",
  56004=>"110010011",
  56005=>"100110001",
  56006=>"011011001",
  56007=>"101110110",
  56008=>"111001101",
  56009=>"100100101",
  56010=>"010100101",
  56011=>"000000100",
  56012=>"111011100",
  56013=>"111010101",
  56014=>"101000100",
  56015=>"101011110",
  56016=>"001101011",
  56017=>"100000100",
  56018=>"001010010",
  56019=>"000001001",
  56020=>"101000000",
  56021=>"100000110",
  56022=>"100100011",
  56023=>"111110100",
  56024=>"001101010",
  56025=>"000100110",
  56026=>"001110111",
  56027=>"001010000",
  56028=>"001010011",
  56029=>"000101000",
  56030=>"100100010",
  56031=>"010011011",
  56032=>"100011100",
  56033=>"010000110",
  56034=>"101100010",
  56035=>"000110110",
  56036=>"100110101",
  56037=>"010111110",
  56038=>"010000111",
  56039=>"011000101",
  56040=>"000101001",
  56041=>"011101001",
  56042=>"000000010",
  56043=>"010010001",
  56044=>"010111011",
  56045=>"110001111",
  56046=>"111000000",
  56047=>"100110100",
  56048=>"101101111",
  56049=>"101111011",
  56050=>"000011001",
  56051=>"000110100",
  56052=>"011000001",
  56053=>"111000101",
  56054=>"000010010",
  56055=>"001000110",
  56056=>"111100110",
  56057=>"011000001",
  56058=>"100100001",
  56059=>"011010111",
  56060=>"001010110",
  56061=>"110101101",
  56062=>"001001101",
  56063=>"010011101",
  56064=>"000010110",
  56065=>"010011100",
  56066=>"110010110",
  56067=>"111011101",
  56068=>"110001101",
  56069=>"001100000",
  56070=>"101000101",
  56071=>"010111010",
  56072=>"000111111",
  56073=>"010110010",
  56074=>"001011000",
  56075=>"010011000",
  56076=>"001101110",
  56077=>"011101000",
  56078=>"011000101",
  56079=>"010101111",
  56080=>"011101011",
  56081=>"001000000",
  56082=>"011001101",
  56083=>"011001111",
  56084=>"001010001",
  56085=>"001110101",
  56086=>"011101001",
  56087=>"101110001",
  56088=>"010100010",
  56089=>"110010001",
  56090=>"101110110",
  56091=>"101010010",
  56092=>"100001110",
  56093=>"011011000",
  56094=>"111100110",
  56095=>"101000010",
  56096=>"001100111",
  56097=>"010000101",
  56098=>"110111100",
  56099=>"000111010",
  56100=>"101100111",
  56101=>"101001101",
  56102=>"101110001",
  56103=>"010000000",
  56104=>"010011001",
  56105=>"110000000",
  56106=>"011111010",
  56107=>"110000011",
  56108=>"110111000",
  56109=>"101110001",
  56110=>"111101110",
  56111=>"100101011",
  56112=>"001010101",
  56113=>"000101110",
  56114=>"011111101",
  56115=>"111011000",
  56116=>"111010010",
  56117=>"000011101",
  56118=>"100010001",
  56119=>"101101111",
  56120=>"010111110",
  56121=>"111000011",
  56122=>"110111001",
  56123=>"011100110",
  56124=>"111101110",
  56125=>"101111111",
  56126=>"010001111",
  56127=>"011000000",
  56128=>"111110100",
  56129=>"111000001",
  56130=>"010000100",
  56131=>"000000000",
  56132=>"001011101",
  56133=>"011011101",
  56134=>"100001110",
  56135=>"000111101",
  56136=>"011100000",
  56137=>"110010111",
  56138=>"011010101",
  56139=>"001101110",
  56140=>"000000110",
  56141=>"000001001",
  56142=>"000000100",
  56143=>"100100000",
  56144=>"101100110",
  56145=>"001010011",
  56146=>"000000110",
  56147=>"001111000",
  56148=>"001101111",
  56149=>"110101111",
  56150=>"101001101",
  56151=>"111111010",
  56152=>"111101011",
  56153=>"000101101",
  56154=>"100010011",
  56155=>"001000000",
  56156=>"010111001",
  56157=>"000110000",
  56158=>"001001110",
  56159=>"000101111",
  56160=>"010110000",
  56161=>"110110011",
  56162=>"010010100",
  56163=>"011011011",
  56164=>"010101110",
  56165=>"000101101",
  56166=>"001011011",
  56167=>"000100101",
  56168=>"111011011",
  56169=>"000100110",
  56170=>"111011110",
  56171=>"011001101",
  56172=>"111100101",
  56173=>"011001001",
  56174=>"000001000",
  56175=>"100010000",
  56176=>"100100001",
  56177=>"111011100",
  56178=>"100100001",
  56179=>"000110000",
  56180=>"011100110",
  56181=>"100100010",
  56182=>"101110110",
  56183=>"010100101",
  56184=>"000011111",
  56185=>"001011000",
  56186=>"101111101",
  56187=>"110010100",
  56188=>"001000010",
  56189=>"101000000",
  56190=>"111100010",
  56191=>"010011010",
  56192=>"101011011",
  56193=>"001101010",
  56194=>"110000111",
  56195=>"111110000",
  56196=>"000100100",
  56197=>"110100011",
  56198=>"000100011",
  56199=>"001101100",
  56200=>"000110100",
  56201=>"001110001",
  56202=>"000111110",
  56203=>"100100000",
  56204=>"001110100",
  56205=>"100011111",
  56206=>"100111010",
  56207=>"100101000",
  56208=>"101100000",
  56209=>"001000010",
  56210=>"100010111",
  56211=>"110100000",
  56212=>"001010010",
  56213=>"110111101",
  56214=>"010101011",
  56215=>"101100110",
  56216=>"001011111",
  56217=>"011111011",
  56218=>"111101100",
  56219=>"100100110",
  56220=>"011110111",
  56221=>"010001100",
  56222=>"010100111",
  56223=>"000001001",
  56224=>"010100000",
  56225=>"001010110",
  56226=>"001011111",
  56227=>"011101001",
  56228=>"001000011",
  56229=>"110100111",
  56230=>"000101111",
  56231=>"001000011",
  56232=>"000110100",
  56233=>"011000111",
  56234=>"110010001",
  56235=>"111101001",
  56236=>"000001011",
  56237=>"101101001",
  56238=>"000011110",
  56239=>"010110101",
  56240=>"110101111",
  56241=>"000111011",
  56242=>"000011111",
  56243=>"010101001",
  56244=>"011000001",
  56245=>"001110011",
  56246=>"001000001",
  56247=>"010011000",
  56248=>"000100000",
  56249=>"001000000",
  56250=>"011000000",
  56251=>"000111100",
  56252=>"000001000",
  56253=>"100011111",
  56254=>"111001011",
  56255=>"001010100",
  56256=>"111010010",
  56257=>"000111001",
  56258=>"111111011",
  56259=>"011110111",
  56260=>"111111000",
  56261=>"001001111",
  56262=>"110100001",
  56263=>"111111111",
  56264=>"010101001",
  56265=>"010100000",
  56266=>"011001110",
  56267=>"110010110",
  56268=>"110110101",
  56269=>"001010000",
  56270=>"010111101",
  56271=>"100010101",
  56272=>"100101110",
  56273=>"011000000",
  56274=>"000100000",
  56275=>"010010001",
  56276=>"111010101",
  56277=>"010011001",
  56278=>"111111101",
  56279=>"001001011",
  56280=>"101010111",
  56281=>"000111111",
  56282=>"101010100",
  56283=>"100001010",
  56284=>"111111111",
  56285=>"101010011",
  56286=>"010101111",
  56287=>"101010101",
  56288=>"001111110",
  56289=>"111100111",
  56290=>"011001100",
  56291=>"101101000",
  56292=>"110101111",
  56293=>"101110010",
  56294=>"100000000",
  56295=>"100000010",
  56296=>"000000110",
  56297=>"001110111",
  56298=>"101000100",
  56299=>"000011111",
  56300=>"011011111",
  56301=>"100001011",
  56302=>"000111000",
  56303=>"111101100",
  56304=>"101110101",
  56305=>"101010001",
  56306=>"100101101",
  56307=>"010100010",
  56308=>"010101111",
  56309=>"100111111",
  56310=>"110111000",
  56311=>"010001100",
  56312=>"111111101",
  56313=>"000001101",
  56314=>"000001010",
  56315=>"010011000",
  56316=>"111110001",
  56317=>"010111100",
  56318=>"100111111",
  56319=>"110010110",
  56320=>"010011011",
  56321=>"111000000",
  56322=>"111111111",
  56323=>"010011101",
  56324=>"000001000",
  56325=>"100110011",
  56326=>"000001000",
  56327=>"000000000",
  56328=>"011001001",
  56329=>"010100001",
  56330=>"110000111",
  56331=>"110000101",
  56332=>"000010010",
  56333=>"111111100",
  56334=>"000100000",
  56335=>"011110101",
  56336=>"011101010",
  56337=>"010001010",
  56338=>"101011111",
  56339=>"101100011",
  56340=>"101111010",
  56341=>"001001111",
  56342=>"111110000",
  56343=>"001111110",
  56344=>"100011110",
  56345=>"001100110",
  56346=>"000101011",
  56347=>"101001010",
  56348=>"010001001",
  56349=>"110110010",
  56350=>"110011100",
  56351=>"101010001",
  56352=>"101010010",
  56353=>"110001111",
  56354=>"111100100",
  56355=>"100100010",
  56356=>"110111000",
  56357=>"111100110",
  56358=>"100101111",
  56359=>"010100100",
  56360=>"100001110",
  56361=>"000010110",
  56362=>"010001110",
  56363=>"111011010",
  56364=>"000000010",
  56365=>"100011001",
  56366=>"110111010",
  56367=>"011101110",
  56368=>"101000010",
  56369=>"000111011",
  56370=>"000010000",
  56371=>"110010100",
  56372=>"111111111",
  56373=>"000000100",
  56374=>"000100101",
  56375=>"111100000",
  56376=>"001110001",
  56377=>"101100010",
  56378=>"000010110",
  56379=>"100011000",
  56380=>"010000000",
  56381=>"010010010",
  56382=>"110011100",
  56383=>"100111000",
  56384=>"101110001",
  56385=>"110000010",
  56386=>"100111001",
  56387=>"011110000",
  56388=>"010101000",
  56389=>"011010011",
  56390=>"011101110",
  56391=>"010011010",
  56392=>"001100100",
  56393=>"111010011",
  56394=>"110110001",
  56395=>"011011010",
  56396=>"101111101",
  56397=>"110101101",
  56398=>"001111001",
  56399=>"000110010",
  56400=>"111011100",
  56401=>"000111010",
  56402=>"110001011",
  56403=>"100000011",
  56404=>"000011100",
  56405=>"000001011",
  56406=>"001100001",
  56407=>"010000111",
  56408=>"000111010",
  56409=>"100111111",
  56410=>"100000001",
  56411=>"111100101",
  56412=>"000001101",
  56413=>"101010101",
  56414=>"010100101",
  56415=>"101010101",
  56416=>"110100110",
  56417=>"000000100",
  56418=>"100110000",
  56419=>"100000100",
  56420=>"111000101",
  56421=>"011111110",
  56422=>"010011010",
  56423=>"101110100",
  56424=>"000011010",
  56425=>"100111011",
  56426=>"000000100",
  56427=>"110001100",
  56428=>"001100110",
  56429=>"100010101",
  56430=>"010110001",
  56431=>"111100110",
  56432=>"000001010",
  56433=>"010000110",
  56434=>"011100000",
  56435=>"100001101",
  56436=>"110010110",
  56437=>"001001001",
  56438=>"011110101",
  56439=>"101010010",
  56440=>"110111000",
  56441=>"010100111",
  56442=>"111111011",
  56443=>"010000011",
  56444=>"100011001",
  56445=>"001011100",
  56446=>"110111111",
  56447=>"000001000",
  56448=>"010000100",
  56449=>"000101100",
  56450=>"010111011",
  56451=>"100101000",
  56452=>"000111000",
  56453=>"100011111",
  56454=>"011011001",
  56455=>"000010100",
  56456=>"011111010",
  56457=>"000111011",
  56458=>"011000100",
  56459=>"101100101",
  56460=>"000101110",
  56461=>"110001010",
  56462=>"010100010",
  56463=>"100111010",
  56464=>"010100111",
  56465=>"110100101",
  56466=>"010011001",
  56467=>"011010001",
  56468=>"100110001",
  56469=>"010111001",
  56470=>"001010000",
  56471=>"011001001",
  56472=>"000101001",
  56473=>"110001101",
  56474=>"110111100",
  56475=>"000101000",
  56476=>"000101001",
  56477=>"100111101",
  56478=>"011010110",
  56479=>"011010110",
  56480=>"010010101",
  56481=>"111010100",
  56482=>"111100001",
  56483=>"011000111",
  56484=>"101111110",
  56485=>"110110100",
  56486=>"101100100",
  56487=>"111111111",
  56488=>"001100000",
  56489=>"010110010",
  56490=>"000111001",
  56491=>"000011101",
  56492=>"101001010",
  56493=>"101011000",
  56494=>"110100001",
  56495=>"111011010",
  56496=>"111101100",
  56497=>"111001001",
  56498=>"001011100",
  56499=>"101110011",
  56500=>"000110111",
  56501=>"000010000",
  56502=>"001111101",
  56503=>"111001011",
  56504=>"110001110",
  56505=>"101000100",
  56506=>"001110000",
  56507=>"100000000",
  56508=>"100011011",
  56509=>"110111011",
  56510=>"011101011",
  56511=>"000010100",
  56512=>"001010110",
  56513=>"011110101",
  56514=>"111111101",
  56515=>"101000001",
  56516=>"010000000",
  56517=>"101111001",
  56518=>"010111111",
  56519=>"101101011",
  56520=>"011100111",
  56521=>"001101100",
  56522=>"010110101",
  56523=>"110110011",
  56524=>"000010101",
  56525=>"001011010",
  56526=>"110001010",
  56527=>"001110011",
  56528=>"000011100",
  56529=>"110001011",
  56530=>"100010001",
  56531=>"010001100",
  56532=>"101001000",
  56533=>"101001000",
  56534=>"001010101",
  56535=>"010010011",
  56536=>"001100000",
  56537=>"010111100",
  56538=>"111100101",
  56539=>"001000111",
  56540=>"101010000",
  56541=>"110110000",
  56542=>"011100100",
  56543=>"111100101",
  56544=>"010001000",
  56545=>"010110011",
  56546=>"110101000",
  56547=>"101100110",
  56548=>"010101111",
  56549=>"101110001",
  56550=>"010000100",
  56551=>"010100110",
  56552=>"110010111",
  56553=>"100101110",
  56554=>"100001100",
  56555=>"101000111",
  56556=>"100101111",
  56557=>"100101110",
  56558=>"101000111",
  56559=>"000001011",
  56560=>"110101010",
  56561=>"111010110",
  56562=>"011000100",
  56563=>"010011011",
  56564=>"011101111",
  56565=>"101111100",
  56566=>"101011011",
  56567=>"100100100",
  56568=>"110001000",
  56569=>"011011001",
  56570=>"000000001",
  56571=>"100011100",
  56572=>"110110000",
  56573=>"100011110",
  56574=>"010000100",
  56575=>"001010000",
  56576=>"111110010",
  56577=>"110101011",
  56578=>"110111110",
  56579=>"101010111",
  56580=>"011011011",
  56581=>"110001100",
  56582=>"010011111",
  56583=>"001000100",
  56584=>"001001010",
  56585=>"001111011",
  56586=>"111001101",
  56587=>"000011011",
  56588=>"100111100",
  56589=>"000110100",
  56590=>"101101111",
  56591=>"000000101",
  56592=>"011101111",
  56593=>"110000110",
  56594=>"101010011",
  56595=>"111011101",
  56596=>"101110111",
  56597=>"000110110",
  56598=>"000111000",
  56599=>"111111001",
  56600=>"100000101",
  56601=>"011011001",
  56602=>"011011001",
  56603=>"010110110",
  56604=>"000100111",
  56605=>"100001000",
  56606=>"111011110",
  56607=>"111100001",
  56608=>"000010001",
  56609=>"110100001",
  56610=>"101110111",
  56611=>"110100000",
  56612=>"011100011",
  56613=>"111101011",
  56614=>"000100000",
  56615=>"101001100",
  56616=>"011111101",
  56617=>"111010111",
  56618=>"111011010",
  56619=>"010000011",
  56620=>"101100100",
  56621=>"001001100",
  56622=>"000111001",
  56623=>"001000011",
  56624=>"001100110",
  56625=>"101011010",
  56626=>"010000001",
  56627=>"111001000",
  56628=>"010011010",
  56629=>"001100111",
  56630=>"010110000",
  56631=>"010011000",
  56632=>"101111100",
  56633=>"011111000",
  56634=>"001100010",
  56635=>"010100000",
  56636=>"010011010",
  56637=>"001110101",
  56638=>"010001000",
  56639=>"011001011",
  56640=>"011111010",
  56641=>"010111110",
  56642=>"100110000",
  56643=>"100101011",
  56644=>"011100000",
  56645=>"010010101",
  56646=>"110011001",
  56647=>"100010101",
  56648=>"011011000",
  56649=>"011010010",
  56650=>"000101111",
  56651=>"010010011",
  56652=>"111101110",
  56653=>"100000101",
  56654=>"010110101",
  56655=>"001111111",
  56656=>"101001101",
  56657=>"011001111",
  56658=>"111111011",
  56659=>"111101000",
  56660=>"010000000",
  56661=>"100010100",
  56662=>"111111100",
  56663=>"110110000",
  56664=>"101011100",
  56665=>"101110001",
  56666=>"100001011",
  56667=>"100000111",
  56668=>"101000011",
  56669=>"110110000",
  56670=>"000011010",
  56671=>"001000010",
  56672=>"101011010",
  56673=>"111001100",
  56674=>"100111110",
  56675=>"010000000",
  56676=>"111101011",
  56677=>"011100101",
  56678=>"101000011",
  56679=>"010001000",
  56680=>"101110101",
  56681=>"111110010",
  56682=>"100010011",
  56683=>"101000011",
  56684=>"101001010",
  56685=>"000111110",
  56686=>"100110100",
  56687=>"100110110",
  56688=>"110100010",
  56689=>"110011000",
  56690=>"010110101",
  56691=>"111101001",
  56692=>"111001010",
  56693=>"110111000",
  56694=>"100000011",
  56695=>"111101111",
  56696=>"000111111",
  56697=>"110001111",
  56698=>"110010001",
  56699=>"110000110",
  56700=>"111111000",
  56701=>"000000000",
  56702=>"110001110",
  56703=>"110110111",
  56704=>"110000001",
  56705=>"101100111",
  56706=>"110001000",
  56707=>"000001010",
  56708=>"110111000",
  56709=>"101010011",
  56710=>"000000011",
  56711=>"010110101",
  56712=>"010100100",
  56713=>"011110001",
  56714=>"110010001",
  56715=>"000111001",
  56716=>"000001000",
  56717=>"001110110",
  56718=>"110101101",
  56719=>"001001001",
  56720=>"010000111",
  56721=>"010010101",
  56722=>"100110101",
  56723=>"010011001",
  56724=>"101111011",
  56725=>"110101110",
  56726=>"000110101",
  56727=>"111111111",
  56728=>"000101011",
  56729=>"011110001",
  56730=>"010011011",
  56731=>"011111111",
  56732=>"011001000",
  56733=>"011001010",
  56734=>"110101110",
  56735=>"000000010",
  56736=>"101010010",
  56737=>"101101011",
  56738=>"100100100",
  56739=>"010011111",
  56740=>"101011111",
  56741=>"010000100",
  56742=>"100010110",
  56743=>"110010111",
  56744=>"010100001",
  56745=>"010000000",
  56746=>"010000010",
  56747=>"010001101",
  56748=>"001100011",
  56749=>"010000111",
  56750=>"101110111",
  56751=>"001111111",
  56752=>"010101011",
  56753=>"000000101",
  56754=>"001011011",
  56755=>"111111111",
  56756=>"000100000",
  56757=>"111101001",
  56758=>"101001001",
  56759=>"110011110",
  56760=>"011110011",
  56761=>"001100111",
  56762=>"010000100",
  56763=>"010010000",
  56764=>"111011000",
  56765=>"110000100",
  56766=>"000101110",
  56767=>"101010101",
  56768=>"101011001",
  56769=>"100100101",
  56770=>"101111101",
  56771=>"110101101",
  56772=>"001010111",
  56773=>"001011111",
  56774=>"111001110",
  56775=>"100111101",
  56776=>"011010011",
  56777=>"011100100",
  56778=>"111101011",
  56779=>"111000010",
  56780=>"111010111",
  56781=>"000101111",
  56782=>"100100001",
  56783=>"100100110",
  56784=>"001100010",
  56785=>"110010000",
  56786=>"001100101",
  56787=>"110101101",
  56788=>"001011100",
  56789=>"010100011",
  56790=>"100010010",
  56791=>"000110000",
  56792=>"010100100",
  56793=>"010010001",
  56794=>"000101111",
  56795=>"101011011",
  56796=>"000010011",
  56797=>"111000010",
  56798=>"001100001",
  56799=>"100001110",
  56800=>"100101111",
  56801=>"100011001",
  56802=>"010111000",
  56803=>"000101111",
  56804=>"101100000",
  56805=>"100110100",
  56806=>"000100000",
  56807=>"011111101",
  56808=>"000101011",
  56809=>"010000011",
  56810=>"111111101",
  56811=>"000110100",
  56812=>"100010001",
  56813=>"011010101",
  56814=>"010010001",
  56815=>"111000100",
  56816=>"000011110",
  56817=>"110100110",
  56818=>"110111101",
  56819=>"110001010",
  56820=>"100001011",
  56821=>"010110101",
  56822=>"011111000",
  56823=>"000100100",
  56824=>"110111000",
  56825=>"011010010",
  56826=>"101001011",
  56827=>"000101111",
  56828=>"110000000",
  56829=>"101000110",
  56830=>"010010111",
  56831=>"111000100",
  56832=>"111111100",
  56833=>"011110110",
  56834=>"001100010",
  56835=>"001101000",
  56836=>"011001100",
  56837=>"000001111",
  56838=>"010001001",
  56839=>"011101111",
  56840=>"110110110",
  56841=>"111010111",
  56842=>"000000000",
  56843=>"001011000",
  56844=>"101110110",
  56845=>"001001010",
  56846=>"010011010",
  56847=>"101001110",
  56848=>"111110011",
  56849=>"001000100",
  56850=>"101000010",
  56851=>"001000011",
  56852=>"111010111",
  56853=>"111100110",
  56854=>"010101001",
  56855=>"011000111",
  56856=>"001100001",
  56857=>"010100110",
  56858=>"111010001",
  56859=>"001101011",
  56860=>"001101001",
  56861=>"101010000",
  56862=>"110111011",
  56863=>"110000000",
  56864=>"000101011",
  56865=>"110011101",
  56866=>"101000110",
  56867=>"100101000",
  56868=>"011011110",
  56869=>"000011011",
  56870=>"110001101",
  56871=>"011111001",
  56872=>"111000110",
  56873=>"000001111",
  56874=>"011000110",
  56875=>"000001100",
  56876=>"011000000",
  56877=>"101111110",
  56878=>"101110000",
  56879=>"110000100",
  56880=>"001000011",
  56881=>"100001101",
  56882=>"000000101",
  56883=>"101110010",
  56884=>"100000101",
  56885=>"001001100",
  56886=>"001110001",
  56887=>"111101011",
  56888=>"001010110",
  56889=>"100010000",
  56890=>"111010010",
  56891=>"101101100",
  56892=>"101110011",
  56893=>"111001110",
  56894=>"011010000",
  56895=>"101011101",
  56896=>"010110010",
  56897=>"010110000",
  56898=>"101000000",
  56899=>"101000111",
  56900=>"100011100",
  56901=>"010011100",
  56902=>"000101011",
  56903=>"000001001",
  56904=>"000100001",
  56905=>"001010000",
  56906=>"101111010",
  56907=>"000101101",
  56908=>"101100111",
  56909=>"111000000",
  56910=>"001000000",
  56911=>"101001010",
  56912=>"011000010",
  56913=>"000000001",
  56914=>"111010110",
  56915=>"100011110",
  56916=>"010000000",
  56917=>"111000011",
  56918=>"011111111",
  56919=>"000001111",
  56920=>"000110001",
  56921=>"111011000",
  56922=>"101000011",
  56923=>"000111000",
  56924=>"111100010",
  56925=>"111000111",
  56926=>"001000110",
  56927=>"001111001",
  56928=>"010010011",
  56929=>"100010010",
  56930=>"101111101",
  56931=>"111100111",
  56932=>"111110100",
  56933=>"101100110",
  56934=>"000001010",
  56935=>"010010001",
  56936=>"000010011",
  56937=>"010100111",
  56938=>"111100110",
  56939=>"110000000",
  56940=>"111111000",
  56941=>"000101010",
  56942=>"101101001",
  56943=>"100111101",
  56944=>"000110101",
  56945=>"111001010",
  56946=>"100101100",
  56947=>"010011010",
  56948=>"110001111",
  56949=>"110000000",
  56950=>"000110010",
  56951=>"101111000",
  56952=>"111111110",
  56953=>"101101010",
  56954=>"110110011",
  56955=>"101110110",
  56956=>"101010110",
  56957=>"000000011",
  56958=>"101011011",
  56959=>"000001001",
  56960=>"010101110",
  56961=>"111100010",
  56962=>"001100011",
  56963=>"110000011",
  56964=>"110111100",
  56965=>"110110111",
  56966=>"010010001",
  56967=>"110000111",
  56968=>"100110111",
  56969=>"001101011",
  56970=>"111100010",
  56971=>"101110110",
  56972=>"001011000",
  56973=>"110000001",
  56974=>"010100110",
  56975=>"111101110",
  56976=>"000100010",
  56977=>"011100000",
  56978=>"101100100",
  56979=>"010101111",
  56980=>"000110011",
  56981=>"110110100",
  56982=>"110111011",
  56983=>"110011101",
  56984=>"011111100",
  56985=>"110010010",
  56986=>"011100011",
  56987=>"000001100",
  56988=>"000101000",
  56989=>"001000101",
  56990=>"011000001",
  56991=>"000110100",
  56992=>"110011010",
  56993=>"111111011",
  56994=>"011011011",
  56995=>"111100001",
  56996=>"010000010",
  56997=>"110110010",
  56998=>"011100111",
  56999=>"111110000",
  57000=>"110010000",
  57001=>"001100010",
  57002=>"110100100",
  57003=>"010000101",
  57004=>"011000010",
  57005=>"101000111",
  57006=>"100111000",
  57007=>"011001110",
  57008=>"110010011",
  57009=>"110001010",
  57010=>"000010000",
  57011=>"111011000",
  57012=>"000101001",
  57013=>"111111101",
  57014=>"101001100",
  57015=>"001000000",
  57016=>"100111011",
  57017=>"011111111",
  57018=>"101011110",
  57019=>"110100010",
  57020=>"111000001",
  57021=>"101110110",
  57022=>"000111111",
  57023=>"011110101",
  57024=>"101001010",
  57025=>"100111111",
  57026=>"000011010",
  57027=>"100101010",
  57028=>"011111001",
  57029=>"100011011",
  57030=>"010010000",
  57031=>"001101000",
  57032=>"010100001",
  57033=>"000100011",
  57034=>"110010010",
  57035=>"001100100",
  57036=>"101000101",
  57037=>"101000100",
  57038=>"110110100",
  57039=>"100001010",
  57040=>"100101111",
  57041=>"010101110",
  57042=>"011101001",
  57043=>"011001110",
  57044=>"001000110",
  57045=>"010101101",
  57046=>"100111001",
  57047=>"001010110",
  57048=>"000000110",
  57049=>"010001010",
  57050=>"101101101",
  57051=>"000111011",
  57052=>"111110001",
  57053=>"110110011",
  57054=>"010110111",
  57055=>"101110010",
  57056=>"010111001",
  57057=>"111001011",
  57058=>"111001011",
  57059=>"000000101",
  57060=>"010000110",
  57061=>"110100011",
  57062=>"010001010",
  57063=>"111110000",
  57064=>"110111110",
  57065=>"111101001",
  57066=>"011010100",
  57067=>"000100100",
  57068=>"111100001",
  57069=>"101011011",
  57070=>"011100011",
  57071=>"011110001",
  57072=>"111000001",
  57073=>"100010010",
  57074=>"010100011",
  57075=>"111011111",
  57076=>"011101011",
  57077=>"111001110",
  57078=>"111011010",
  57079=>"110101110",
  57080=>"100011110",
  57081=>"001110100",
  57082=>"000100110",
  57083=>"111010011",
  57084=>"011101111",
  57085=>"001110110",
  57086=>"110010011",
  57087=>"110011111",
  57088=>"011010100",
  57089=>"001101100",
  57090=>"101010111",
  57091=>"011001000",
  57092=>"101111011",
  57093=>"001000111",
  57094=>"000001011",
  57095=>"010101001",
  57096=>"011111110",
  57097=>"011101001",
  57098=>"001100001",
  57099=>"100001000",
  57100=>"110111111",
  57101=>"010011110",
  57102=>"000011011",
  57103=>"010010001",
  57104=>"001001011",
  57105=>"010011000",
  57106=>"100110011",
  57107=>"000000111",
  57108=>"010111101",
  57109=>"010101000",
  57110=>"010000001",
  57111=>"100010010",
  57112=>"100110000",
  57113=>"010111100",
  57114=>"011101011",
  57115=>"110100111",
  57116=>"010001111",
  57117=>"111110011",
  57118=>"011001000",
  57119=>"001011001",
  57120=>"111010001",
  57121=>"010100100",
  57122=>"010001011",
  57123=>"111100000",
  57124=>"010100111",
  57125=>"110011100",
  57126=>"001100000",
  57127=>"110011011",
  57128=>"110011011",
  57129=>"000111001",
  57130=>"010011011",
  57131=>"100100011",
  57132=>"001010011",
  57133=>"100110010",
  57134=>"110000000",
  57135=>"100000000",
  57136=>"011011101",
  57137=>"100100110",
  57138=>"010111000",
  57139=>"000100111",
  57140=>"100010111",
  57141=>"011000000",
  57142=>"010010111",
  57143=>"100101111",
  57144=>"011111111",
  57145=>"101101101",
  57146=>"011100010",
  57147=>"000110000",
  57148=>"001000101",
  57149=>"100000001",
  57150=>"010111101",
  57151=>"011000000",
  57152=>"010000011",
  57153=>"001110001",
  57154=>"100001011",
  57155=>"011101001",
  57156=>"111011011",
  57157=>"111110101",
  57158=>"000010100",
  57159=>"011000110",
  57160=>"100001011",
  57161=>"011100100",
  57162=>"001110001",
  57163=>"100011001",
  57164=>"001111100",
  57165=>"000001111",
  57166=>"010010110",
  57167=>"000001000",
  57168=>"111101111",
  57169=>"000110000",
  57170=>"001111000",
  57171=>"100000000",
  57172=>"011110011",
  57173=>"111111101",
  57174=>"001100110",
  57175=>"011101000",
  57176=>"101010001",
  57177=>"110100001",
  57178=>"000100011",
  57179=>"100101011",
  57180=>"110100111",
  57181=>"001111001",
  57182=>"011010000",
  57183=>"111111111",
  57184=>"001110110",
  57185=>"011011100",
  57186=>"011001011",
  57187=>"010011110",
  57188=>"011100000",
  57189=>"000101010",
  57190=>"011111011",
  57191=>"111101111",
  57192=>"100100001",
  57193=>"011011011",
  57194=>"011110000",
  57195=>"000101111",
  57196=>"001111101",
  57197=>"010010101",
  57198=>"010100011",
  57199=>"010001001",
  57200=>"111101110",
  57201=>"000100010",
  57202=>"111010111",
  57203=>"001101010",
  57204=>"111010010",
  57205=>"101011111",
  57206=>"001011001",
  57207=>"001000000",
  57208=>"011000001",
  57209=>"101110101",
  57210=>"000100110",
  57211=>"110111111",
  57212=>"100010010",
  57213=>"010010111",
  57214=>"000000101",
  57215=>"110010010",
  57216=>"100111111",
  57217=>"111000110",
  57218=>"111110110",
  57219=>"011001110",
  57220=>"001000011",
  57221=>"000101011",
  57222=>"011000010",
  57223=>"100011101",
  57224=>"000111101",
  57225=>"000110000",
  57226=>"011100010",
  57227=>"111111010",
  57228=>"101100101",
  57229=>"001000001",
  57230=>"000111111",
  57231=>"110100011",
  57232=>"111011000",
  57233=>"000011010",
  57234=>"001000010",
  57235=>"010101010",
  57236=>"010100100",
  57237=>"001110000",
  57238=>"110001011",
  57239=>"100101110",
  57240=>"010011010",
  57241=>"010100100",
  57242=>"110000101",
  57243=>"101100110",
  57244=>"001110100",
  57245=>"101001110",
  57246=>"011101010",
  57247=>"110101100",
  57248=>"000001100",
  57249=>"000110011",
  57250=>"001011010",
  57251=>"000001100",
  57252=>"100011001",
  57253=>"001000110",
  57254=>"001001110",
  57255=>"011011001",
  57256=>"100110011",
  57257=>"101011001",
  57258=>"111000001",
  57259=>"010100011",
  57260=>"000001010",
  57261=>"101111101",
  57262=>"110011000",
  57263=>"100111000",
  57264=>"000110100",
  57265=>"010101010",
  57266=>"100000100",
  57267=>"010101110",
  57268=>"111111011",
  57269=>"111111100",
  57270=>"100110000",
  57271=>"111001001",
  57272=>"100010010",
  57273=>"001001100",
  57274=>"100101110",
  57275=>"000101010",
  57276=>"110110101",
  57277=>"011011010",
  57278=>"001010100",
  57279=>"011111101",
  57280=>"001011111",
  57281=>"100110011",
  57282=>"110111110",
  57283=>"000101100",
  57284=>"101001000",
  57285=>"110001011",
  57286=>"011010110",
  57287=>"000111111",
  57288=>"101010011",
  57289=>"001000111",
  57290=>"100111000",
  57291=>"000110111",
  57292=>"001011110",
  57293=>"001000001",
  57294=>"101011111",
  57295=>"110101000",
  57296=>"001100000",
  57297=>"010110101",
  57298=>"010001011",
  57299=>"000101011",
  57300=>"100110101",
  57301=>"110111100",
  57302=>"100010100",
  57303=>"100100111",
  57304=>"001010011",
  57305=>"101110001",
  57306=>"011010000",
  57307=>"101101001",
  57308=>"100100000",
  57309=>"000001110",
  57310=>"000010011",
  57311=>"000011011",
  57312=>"111100001",
  57313=>"100101010",
  57314=>"100100101",
  57315=>"110100100",
  57316=>"101010010",
  57317=>"010000100",
  57318=>"000101010",
  57319=>"100000000",
  57320=>"001001010",
  57321=>"010001110",
  57322=>"100111000",
  57323=>"000000011",
  57324=>"101010111",
  57325=>"110001000",
  57326=>"001000001",
  57327=>"001001010",
  57328=>"111000100",
  57329=>"111010001",
  57330=>"011100110",
  57331=>"001100011",
  57332=>"000001101",
  57333=>"101111101",
  57334=>"110010000",
  57335=>"111000000",
  57336=>"101000001",
  57337=>"010010111",
  57338=>"101010011",
  57339=>"010110111",
  57340=>"000010000",
  57341=>"110110001",
  57342=>"001011010",
  57343=>"011011011",
  57344=>"101001110",
  57345=>"111101001",
  57346=>"111000111",
  57347=>"111111011",
  57348=>"100000111",
  57349=>"000001001",
  57350=>"000011000",
  57351=>"001111010",
  57352=>"110001001",
  57353=>"000110000",
  57354=>"110111011",
  57355=>"010100110",
  57356=>"001010000",
  57357=>"111000000",
  57358=>"011100010",
  57359=>"001010011",
  57360=>"010101000",
  57361=>"110100010",
  57362=>"010001111",
  57363=>"010100000",
  57364=>"111001101",
  57365=>"110110100",
  57366=>"011101001",
  57367=>"100000101",
  57368=>"011000100",
  57369=>"000010111",
  57370=>"001011011",
  57371=>"000000101",
  57372=>"000101010",
  57373=>"101001110",
  57374=>"100111111",
  57375=>"000110011",
  57376=>"010001000",
  57377=>"001101100",
  57378=>"111111110",
  57379=>"011100111",
  57380=>"100100001",
  57381=>"001010100",
  57382=>"010001010",
  57383=>"111001000",
  57384=>"110110111",
  57385=>"100000010",
  57386=>"011000111",
  57387=>"101110110",
  57388=>"101100000",
  57389=>"010110111",
  57390=>"000001011",
  57391=>"111111111",
  57392=>"110011111",
  57393=>"001000111",
  57394=>"110010101",
  57395=>"100110101",
  57396=>"110000101",
  57397=>"011101000",
  57398=>"010110000",
  57399=>"100011101",
  57400=>"100000001",
  57401=>"101111010",
  57402=>"110110010",
  57403=>"100101111",
  57404=>"100011011",
  57405=>"100110001",
  57406=>"001000100",
  57407=>"010010000",
  57408=>"100100111",
  57409=>"010000101",
  57410=>"011011001",
  57411=>"101110100",
  57412=>"100111011",
  57413=>"010010000",
  57414=>"010100100",
  57415=>"101001011",
  57416=>"001010000",
  57417=>"111111010",
  57418=>"100101001",
  57419=>"001111001",
  57420=>"001100000",
  57421=>"101000101",
  57422=>"000111101",
  57423=>"011000100",
  57424=>"010010011",
  57425=>"100001000",
  57426=>"110010010",
  57427=>"001000100",
  57428=>"011000000",
  57429=>"101001110",
  57430=>"111010100",
  57431=>"000011000",
  57432=>"001100000",
  57433=>"100111111",
  57434=>"110010000",
  57435=>"100101010",
  57436=>"001111111",
  57437=>"010001001",
  57438=>"001001010",
  57439=>"000000100",
  57440=>"010001000",
  57441=>"011110010",
  57442=>"001001100",
  57443=>"000100001",
  57444=>"011110000",
  57445=>"011010001",
  57446=>"110000001",
  57447=>"111110100",
  57448=>"000000010",
  57449=>"010100111",
  57450=>"000111100",
  57451=>"011001100",
  57452=>"001001101",
  57453=>"011101100",
  57454=>"011101000",
  57455=>"111100011",
  57456=>"111111000",
  57457=>"000000000",
  57458=>"101010011",
  57459=>"001000100",
  57460=>"111111010",
  57461=>"000111000",
  57462=>"010010101",
  57463=>"001010011",
  57464=>"011111101",
  57465=>"010111001",
  57466=>"010100100",
  57467=>"110111001",
  57468=>"000011011",
  57469=>"111001101",
  57470=>"010110011",
  57471=>"010001001",
  57472=>"001001000",
  57473=>"100110111",
  57474=>"010100000",
  57475=>"001010000",
  57476=>"101101101",
  57477=>"001001101",
  57478=>"001010100",
  57479=>"100011100",
  57480=>"110111011",
  57481=>"001110110",
  57482=>"000000100",
  57483=>"101000011",
  57484=>"001101001",
  57485=>"111111000",
  57486=>"001110011",
  57487=>"111111000",
  57488=>"010110011",
  57489=>"010010010",
  57490=>"110001110",
  57491=>"011011111",
  57492=>"011010100",
  57493=>"111111010",
  57494=>"101011101",
  57495=>"110100111",
  57496=>"000101101",
  57497=>"001011011",
  57498=>"111000100",
  57499=>"110110011",
  57500=>"101001101",
  57501=>"000000000",
  57502=>"000100000",
  57503=>"101011110",
  57504=>"111000110",
  57505=>"011000000",
  57506=>"000110101",
  57507=>"101100001",
  57508=>"001111001",
  57509=>"001110110",
  57510=>"100101111",
  57511=>"100010001",
  57512=>"111010001",
  57513=>"000011111",
  57514=>"010001010",
  57515=>"111110000",
  57516=>"100110110",
  57517=>"110010111",
  57518=>"100010101",
  57519=>"111110011",
  57520=>"011000010",
  57521=>"110000011",
  57522=>"000011010",
  57523=>"010000101",
  57524=>"001010111",
  57525=>"100100110",
  57526=>"101111000",
  57527=>"001101011",
  57528=>"100110001",
  57529=>"001101100",
  57530=>"100100101",
  57531=>"111111100",
  57532=>"001011010",
  57533=>"001100011",
  57534=>"110111001",
  57535=>"101001111",
  57536=>"010101011",
  57537=>"011111100",
  57538=>"111001100",
  57539=>"101011110",
  57540=>"110010111",
  57541=>"010101010",
  57542=>"001000111",
  57543=>"010100100",
  57544=>"001101000",
  57545=>"011010011",
  57546=>"111111011",
  57547=>"000000001",
  57548=>"110111100",
  57549=>"110110110",
  57550=>"001100010",
  57551=>"111001000",
  57552=>"000000111",
  57553=>"001000101",
  57554=>"100001110",
  57555=>"000000100",
  57556=>"100000001",
  57557=>"011000011",
  57558=>"011111111",
  57559=>"001001101",
  57560=>"101111000",
  57561=>"111110000",
  57562=>"000111001",
  57563=>"110111101",
  57564=>"001110100",
  57565=>"000011100",
  57566=>"011101100",
  57567=>"011000101",
  57568=>"100101110",
  57569=>"001100000",
  57570=>"001010011",
  57571=>"000000000",
  57572=>"110001010",
  57573=>"101101111",
  57574=>"000100011",
  57575=>"000010110",
  57576=>"000010010",
  57577=>"101001100",
  57578=>"010000001",
  57579=>"111000011",
  57580=>"111110001",
  57581=>"000101100",
  57582=>"110110111",
  57583=>"110000001",
  57584=>"100000101",
  57585=>"100101010",
  57586=>"100001110",
  57587=>"101100111",
  57588=>"010110010",
  57589=>"110011111",
  57590=>"011100110",
  57591=>"110100111",
  57592=>"010010001",
  57593=>"111100010",
  57594=>"111100001",
  57595=>"010100000",
  57596=>"010010110",
  57597=>"110111111",
  57598=>"110001000",
  57599=>"111110000",
  57600=>"001001000",
  57601=>"000100000",
  57602=>"010000001",
  57603=>"110111101",
  57604=>"010000100",
  57605=>"101001001",
  57606=>"000001101",
  57607=>"010100010",
  57608=>"000100000",
  57609=>"110100111",
  57610=>"101111011",
  57611=>"010100111",
  57612=>"000111011",
  57613=>"000100000",
  57614=>"001010000",
  57615=>"100111110",
  57616=>"101010110",
  57617=>"000011010",
  57618=>"100101011",
  57619=>"110101011",
  57620=>"000111010",
  57621=>"101101000",
  57622=>"111101111",
  57623=>"101011101",
  57624=>"001001000",
  57625=>"011001011",
  57626=>"010001110",
  57627=>"000011001",
  57628=>"100010010",
  57629=>"101010000",
  57630=>"110001100",
  57631=>"100101111",
  57632=>"011111000",
  57633=>"111111111",
  57634=>"010100111",
  57635=>"100000101",
  57636=>"100111011",
  57637=>"000111100",
  57638=>"000111001",
  57639=>"000010110",
  57640=>"101000011",
  57641=>"010100110",
  57642=>"000000010",
  57643=>"111101101",
  57644=>"101110100",
  57645=>"100010001",
  57646=>"110100010",
  57647=>"101101010",
  57648=>"111010111",
  57649=>"011110101",
  57650=>"111110110",
  57651=>"010011000",
  57652=>"110010011",
  57653=>"100100001",
  57654=>"010010101",
  57655=>"111001001",
  57656=>"111011100",
  57657=>"100000110",
  57658=>"111101111",
  57659=>"111100011",
  57660=>"011001010",
  57661=>"000101000",
  57662=>"011100001",
  57663=>"001110000",
  57664=>"011000001",
  57665=>"001010100",
  57666=>"000101011",
  57667=>"101000111",
  57668=>"000100110",
  57669=>"100001101",
  57670=>"101011010",
  57671=>"110101001",
  57672=>"110111000",
  57673=>"101011000",
  57674=>"100010100",
  57675=>"000100001",
  57676=>"010100011",
  57677=>"110010000",
  57678=>"111110011",
  57679=>"010001010",
  57680=>"011011100",
  57681=>"010001000",
  57682=>"001011000",
  57683=>"001111101",
  57684=>"011101111",
  57685=>"111000001",
  57686=>"011110000",
  57687=>"111001111",
  57688=>"110010010",
  57689=>"101011001",
  57690=>"001111010",
  57691=>"111001000",
  57692=>"111111000",
  57693=>"101111011",
  57694=>"111111100",
  57695=>"011000100",
  57696=>"001100011",
  57697=>"001001010",
  57698=>"000000010",
  57699=>"111000101",
  57700=>"100101000",
  57701=>"001011110",
  57702=>"110011100",
  57703=>"100011010",
  57704=>"100101010",
  57705=>"000000101",
  57706=>"111111001",
  57707=>"010000001",
  57708=>"000110100",
  57709=>"010101010",
  57710=>"100100100",
  57711=>"011100011",
  57712=>"001110011",
  57713=>"111111010",
  57714=>"111111011",
  57715=>"010101110",
  57716=>"100010110",
  57717=>"111000110",
  57718=>"001101001",
  57719=>"111001011",
  57720=>"111000010",
  57721=>"111111011",
  57722=>"010010101",
  57723=>"111000110",
  57724=>"011100011",
  57725=>"101001010",
  57726=>"011100110",
  57727=>"000010101",
  57728=>"000011100",
  57729=>"011101110",
  57730=>"010001100",
  57731=>"100001101",
  57732=>"100111110",
  57733=>"000101111",
  57734=>"011111000",
  57735=>"111110100",
  57736=>"001001100",
  57737=>"000110100",
  57738=>"110000001",
  57739=>"001010001",
  57740=>"000010001",
  57741=>"100011000",
  57742=>"101011010",
  57743=>"000101110",
  57744=>"011011111",
  57745=>"111101000",
  57746=>"110110010",
  57747=>"100011111",
  57748=>"011000110",
  57749=>"101101001",
  57750=>"101001000",
  57751=>"010100000",
  57752=>"101110010",
  57753=>"001011101",
  57754=>"100010110",
  57755=>"101010011",
  57756=>"011011110",
  57757=>"111000110",
  57758=>"101001001",
  57759=>"101000010",
  57760=>"110101000",
  57761=>"100110001",
  57762=>"110011100",
  57763=>"011110100",
  57764=>"111101101",
  57765=>"001010100",
  57766=>"001111001",
  57767=>"110101000",
  57768=>"000010000",
  57769=>"111001111",
  57770=>"111000000",
  57771=>"011000000",
  57772=>"100011101",
  57773=>"100100111",
  57774=>"001100100",
  57775=>"001011011",
  57776=>"010010100",
  57777=>"100110010",
  57778=>"000001100",
  57779=>"100110110",
  57780=>"101001110",
  57781=>"011100111",
  57782=>"000111110",
  57783=>"000001001",
  57784=>"110000001",
  57785=>"100011001",
  57786=>"100001010",
  57787=>"011110000",
  57788=>"101100001",
  57789=>"010010101",
  57790=>"111111111",
  57791=>"111001001",
  57792=>"110110011",
  57793=>"110101000",
  57794=>"010100110",
  57795=>"000010011",
  57796=>"101011111",
  57797=>"010010010",
  57798=>"000110011",
  57799=>"101111001",
  57800=>"001001111",
  57801=>"100011011",
  57802=>"010000100",
  57803=>"010001000",
  57804=>"101011111",
  57805=>"010110000",
  57806=>"010100001",
  57807=>"110100110",
  57808=>"100000100",
  57809=>"000110011",
  57810=>"110101100",
  57811=>"001101110",
  57812=>"000111010",
  57813=>"000001010",
  57814=>"000010000",
  57815=>"000000110",
  57816=>"011001001",
  57817=>"001111110",
  57818=>"111001000",
  57819=>"101111110",
  57820=>"101101010",
  57821=>"101101111",
  57822=>"000011010",
  57823=>"001011011",
  57824=>"111000000",
  57825=>"111100011",
  57826=>"101000000",
  57827=>"110111110",
  57828=>"010101100",
  57829=>"101101110",
  57830=>"111110010",
  57831=>"001011110",
  57832=>"101110110",
  57833=>"101111110",
  57834=>"001000110",
  57835=>"001101110",
  57836=>"100101111",
  57837=>"000100101",
  57838=>"000011011",
  57839=>"100110000",
  57840=>"101010110",
  57841=>"111110110",
  57842=>"111110011",
  57843=>"010001010",
  57844=>"000100010",
  57845=>"011011001",
  57846=>"001011111",
  57847=>"011000110",
  57848=>"000010001",
  57849=>"001110110",
  57850=>"000000110",
  57851=>"011111111",
  57852=>"001101100",
  57853=>"110010001",
  57854=>"100001111",
  57855=>"111111010",
  57856=>"100100110",
  57857=>"010110000",
  57858=>"011111010",
  57859=>"000001111",
  57860=>"110100111",
  57861=>"101001010",
  57862=>"110011001",
  57863=>"111101111",
  57864=>"000001110",
  57865=>"111011011",
  57866=>"111110000",
  57867=>"000000100",
  57868=>"100011010",
  57869=>"000101011",
  57870=>"101010000",
  57871=>"101011001",
  57872=>"011111110",
  57873=>"000010011",
  57874=>"001001001",
  57875=>"100111011",
  57876=>"011001001",
  57877=>"001010000",
  57878=>"000001111",
  57879=>"011011101",
  57880=>"100000100",
  57881=>"110101001",
  57882=>"000010010",
  57883=>"110000000",
  57884=>"011010110",
  57885=>"011000111",
  57886=>"001010000",
  57887=>"011011100",
  57888=>"111011110",
  57889=>"111011011",
  57890=>"001000010",
  57891=>"101100110",
  57892=>"101101111",
  57893=>"011000110",
  57894=>"001010010",
  57895=>"110101101",
  57896=>"011100101",
  57897=>"001001000",
  57898=>"010101010",
  57899=>"001110101",
  57900=>"010100001",
  57901=>"101110000",
  57902=>"111010111",
  57903=>"010110100",
  57904=>"000001000",
  57905=>"001101100",
  57906=>"100100000",
  57907=>"000101111",
  57908=>"011001011",
  57909=>"000010000",
  57910=>"111011001",
  57911=>"100000001",
  57912=>"001100001",
  57913=>"000101100",
  57914=>"011111000",
  57915=>"110111011",
  57916=>"000011010",
  57917=>"001100101",
  57918=>"010001111",
  57919=>"000111001",
  57920=>"010110011",
  57921=>"001000011",
  57922=>"000100000",
  57923=>"101000110",
  57924=>"001111110",
  57925=>"001110011",
  57926=>"101011111",
  57927=>"110100111",
  57928=>"110110010",
  57929=>"011110011",
  57930=>"101110010",
  57931=>"100010100",
  57932=>"001011111",
  57933=>"101011111",
  57934=>"001000110",
  57935=>"100111101",
  57936=>"011010000",
  57937=>"000000010",
  57938=>"000010110",
  57939=>"100110101",
  57940=>"111000000",
  57941=>"110010101",
  57942=>"111100101",
  57943=>"110010010",
  57944=>"000101001",
  57945=>"110011011",
  57946=>"001000110",
  57947=>"011100101",
  57948=>"000001100",
  57949=>"000011011",
  57950=>"101111010",
  57951=>"111000000",
  57952=>"110001000",
  57953=>"000000001",
  57954=>"101110111",
  57955=>"111111000",
  57956=>"101010000",
  57957=>"100010111",
  57958=>"000010000",
  57959=>"101101101",
  57960=>"001110110",
  57961=>"010100110",
  57962=>"000101000",
  57963=>"111111000",
  57964=>"100100101",
  57965=>"010011101",
  57966=>"101101010",
  57967=>"101011111",
  57968=>"111010011",
  57969=>"110100110",
  57970=>"000100000",
  57971=>"100111000",
  57972=>"100101100",
  57973=>"010001111",
  57974=>"100000011",
  57975=>"100011010",
  57976=>"000000010",
  57977=>"100000101",
  57978=>"111111111",
  57979=>"000000111",
  57980=>"111101110",
  57981=>"001000100",
  57982=>"010000001",
  57983=>"100100011",
  57984=>"000011100",
  57985=>"010000000",
  57986=>"011011000",
  57987=>"100000100",
  57988=>"110110111",
  57989=>"100010110",
  57990=>"101110100",
  57991=>"100011111",
  57992=>"100101111",
  57993=>"000000110",
  57994=>"011010011",
  57995=>"000101111",
  57996=>"010110000",
  57997=>"110110101",
  57998=>"110011111",
  57999=>"001011011",
  58000=>"101101111",
  58001=>"101010100",
  58002=>"010011011",
  58003=>"101000000",
  58004=>"011100101",
  58005=>"011100010",
  58006=>"010000110",
  58007=>"100101100",
  58008=>"100010010",
  58009=>"110111010",
  58010=>"010111011",
  58011=>"101101011",
  58012=>"000111111",
  58013=>"111101001",
  58014=>"101111111",
  58015=>"001101101",
  58016=>"110100000",
  58017=>"001111001",
  58018=>"001111110",
  58019=>"000101010",
  58020=>"000000100",
  58021=>"111010110",
  58022=>"111111010",
  58023=>"101110111",
  58024=>"001010100",
  58025=>"000011111",
  58026=>"100110100",
  58027=>"100011000",
  58028=>"001001010",
  58029=>"110100110",
  58030=>"001100101",
  58031=>"000011010",
  58032=>"100000111",
  58033=>"101010100",
  58034=>"111111001",
  58035=>"000011011",
  58036=>"100101000",
  58037=>"001110110",
  58038=>"100000110",
  58039=>"111111000",
  58040=>"110010100",
  58041=>"000000010",
  58042=>"111011100",
  58043=>"100111001",
  58044=>"001101111",
  58045=>"101000001",
  58046=>"100000110",
  58047=>"100111000",
  58048=>"011110000",
  58049=>"100101111",
  58050=>"111101000",
  58051=>"110110110",
  58052=>"100100011",
  58053=>"110011111",
  58054=>"010011111",
  58055=>"001011010",
  58056=>"001111000",
  58057=>"111101110",
  58058=>"001000101",
  58059=>"101101101",
  58060=>"001101011",
  58061=>"100111110",
  58062=>"110110101",
  58063=>"100010001",
  58064=>"011101000",
  58065=>"100111010",
  58066=>"100011000",
  58067=>"101100001",
  58068=>"100000000",
  58069=>"010110100",
  58070=>"110001000",
  58071=>"110101101",
  58072=>"011110101",
  58073=>"000011000",
  58074=>"101111000",
  58075=>"101011000",
  58076=>"000000100",
  58077=>"010100000",
  58078=>"011001010",
  58079=>"010101001",
  58080=>"110001010",
  58081=>"100001111",
  58082=>"010100000",
  58083=>"111100110",
  58084=>"010111000",
  58085=>"010000111",
  58086=>"011111001",
  58087=>"000010110",
  58088=>"110111100",
  58089=>"111101000",
  58090=>"100010111",
  58091=>"110100010",
  58092=>"111111101",
  58093=>"111000010",
  58094=>"010011001",
  58095=>"011001100",
  58096=>"001010001",
  58097=>"111100110",
  58098=>"111010101",
  58099=>"110111111",
  58100=>"101110101",
  58101=>"110001111",
  58102=>"010010111",
  58103=>"000110101",
  58104=>"010110111",
  58105=>"110010000",
  58106=>"101010001",
  58107=>"010011111",
  58108=>"000100110",
  58109=>"000011010",
  58110=>"000010000",
  58111=>"000101110",
  58112=>"111111000",
  58113=>"100010101",
  58114=>"001010010",
  58115=>"000001101",
  58116=>"101000000",
  58117=>"100001011",
  58118=>"011110100",
  58119=>"110010111",
  58120=>"111100000",
  58121=>"011111010",
  58122=>"000110100",
  58123=>"001101100",
  58124=>"111010100",
  58125=>"011100011",
  58126=>"101011110",
  58127=>"000101000",
  58128=>"001110011",
  58129=>"000010000",
  58130=>"111001001",
  58131=>"000110101",
  58132=>"110000000",
  58133=>"110100101",
  58134=>"101110100",
  58135=>"101111001",
  58136=>"000001100",
  58137=>"011111100",
  58138=>"001101011",
  58139=>"011000010",
  58140=>"011011000",
  58141=>"101011101",
  58142=>"011000101",
  58143=>"011100111",
  58144=>"111010111",
  58145=>"101111010",
  58146=>"111000100",
  58147=>"100111011",
  58148=>"110011000",
  58149=>"110000110",
  58150=>"000110010",
  58151=>"110111111",
  58152=>"111010111",
  58153=>"110101001",
  58154=>"001011000",
  58155=>"000111011",
  58156=>"101010110",
  58157=>"100001000",
  58158=>"010100100",
  58159=>"010011111",
  58160=>"010111111",
  58161=>"000000111",
  58162=>"000110101",
  58163=>"111000001",
  58164=>"111111101",
  58165=>"000011000",
  58166=>"000100011",
  58167=>"110110001",
  58168=>"000010110",
  58169=>"010100110",
  58170=>"000001001",
  58171=>"000001100",
  58172=>"110000000",
  58173=>"101011011",
  58174=>"010110001",
  58175=>"010001101",
  58176=>"100000011",
  58177=>"110111011",
  58178=>"101100111",
  58179=>"100100100",
  58180=>"011111000",
  58181=>"010100111",
  58182=>"000000101",
  58183=>"010001001",
  58184=>"101000000",
  58185=>"000111000",
  58186=>"110000000",
  58187=>"010100001",
  58188=>"100010000",
  58189=>"010000110",
  58190=>"101011001",
  58191=>"110111001",
  58192=>"111110101",
  58193=>"110110111",
  58194=>"000110000",
  58195=>"000011100",
  58196=>"001011011",
  58197=>"000111010",
  58198=>"000001001",
  58199=>"000011011",
  58200=>"100000111",
  58201=>"110000110",
  58202=>"101111011",
  58203=>"000000101",
  58204=>"100101001",
  58205=>"000101010",
  58206=>"010010110",
  58207=>"111101101",
  58208=>"100010000",
  58209=>"110000100",
  58210=>"111111000",
  58211=>"000001111",
  58212=>"110011010",
  58213=>"000110110",
  58214=>"001010110",
  58215=>"101001010",
  58216=>"010000111",
  58217=>"111011100",
  58218=>"100010001",
  58219=>"000010010",
  58220=>"000001111",
  58221=>"111000111",
  58222=>"100001110",
  58223=>"010101000",
  58224=>"110111111",
  58225=>"010001101",
  58226=>"011011011",
  58227=>"010111100",
  58228=>"100001010",
  58229=>"000001011",
  58230=>"111101110",
  58231=>"110111001",
  58232=>"001001010",
  58233=>"001001011",
  58234=>"110100101",
  58235=>"101001111",
  58236=>"000101010",
  58237=>"000010111",
  58238=>"000101110",
  58239=>"100011011",
  58240=>"000111010",
  58241=>"001010001",
  58242=>"000110100",
  58243=>"010100111",
  58244=>"111000001",
  58245=>"100010010",
  58246=>"111011010",
  58247=>"000010000",
  58248=>"001010001",
  58249=>"111000001",
  58250=>"000110000",
  58251=>"000111011",
  58252=>"000001111",
  58253=>"110001101",
  58254=>"010000010",
  58255=>"101111110",
  58256=>"101000100",
  58257=>"000000010",
  58258=>"100100100",
  58259=>"100111001",
  58260=>"010010100",
  58261=>"001011010",
  58262=>"101010001",
  58263=>"101011101",
  58264=>"101101111",
  58265=>"011111011",
  58266=>"010010100",
  58267=>"010101011",
  58268=>"000110010",
  58269=>"011001010",
  58270=>"100101000",
  58271=>"001000001",
  58272=>"000010010",
  58273=>"101011110",
  58274=>"010101011",
  58275=>"101010101",
  58276=>"111111111",
  58277=>"100010101",
  58278=>"011111100",
  58279=>"001000101",
  58280=>"110000111",
  58281=>"001000100",
  58282=>"100101111",
  58283=>"100111100",
  58284=>"011111110",
  58285=>"101010110",
  58286=>"001101010",
  58287=>"101101101",
  58288=>"000000100",
  58289=>"110011000",
  58290=>"111100001",
  58291=>"110010010",
  58292=>"101000110",
  58293=>"011000010",
  58294=>"001010001",
  58295=>"001100000",
  58296=>"101101011",
  58297=>"011101001",
  58298=>"101110111",
  58299=>"011101100",
  58300=>"001011001",
  58301=>"011110101",
  58302=>"111001011",
  58303=>"010110000",
  58304=>"101111010",
  58305=>"100010110",
  58306=>"010101111",
  58307=>"010011100",
  58308=>"111001100",
  58309=>"000010000",
  58310=>"001101010",
  58311=>"101100101",
  58312=>"000000110",
  58313=>"100001001",
  58314=>"100010110",
  58315=>"011000000",
  58316=>"000000010",
  58317=>"111111011",
  58318=>"010000100",
  58319=>"100011101",
  58320=>"000110011",
  58321=>"011101001",
  58322=>"000011000",
  58323=>"100101011",
  58324=>"000000010",
  58325=>"110101000",
  58326=>"011110000",
  58327=>"100010111",
  58328=>"000000101",
  58329=>"001111110",
  58330=>"110011100",
  58331=>"011000100",
  58332=>"100000001",
  58333=>"110000011",
  58334=>"110100110",
  58335=>"100100011",
  58336=>"011001100",
  58337=>"010100001",
  58338=>"010011010",
  58339=>"110100011",
  58340=>"010011000",
  58341=>"111110010",
  58342=>"101001000",
  58343=>"111011010",
  58344=>"001000110",
  58345=>"010011110",
  58346=>"000111100",
  58347=>"111010100",
  58348=>"010010111",
  58349=>"011000111",
  58350=>"000001001",
  58351=>"000101011",
  58352=>"000010010",
  58353=>"000001000",
  58354=>"011001110",
  58355=>"001100001",
  58356=>"001111010",
  58357=>"111010010",
  58358=>"000000100",
  58359=>"011110001",
  58360=>"011010010",
  58361=>"000111111",
  58362=>"100011010",
  58363=>"100111000",
  58364=>"100100101",
  58365=>"011010001",
  58366=>"011101100",
  58367=>"000110110",
  58368=>"000010010",
  58369=>"001010101",
  58370=>"101111111",
  58371=>"010011101",
  58372=>"101100111",
  58373=>"111011101",
  58374=>"000001011",
  58375=>"000100101",
  58376=>"111001001",
  58377=>"100110011",
  58378=>"001001000",
  58379=>"110111010",
  58380=>"001101100",
  58381=>"000100011",
  58382=>"010100100",
  58383=>"000001101",
  58384=>"110111100",
  58385=>"001000000",
  58386=>"110011000",
  58387=>"001011000",
  58388=>"101101111",
  58389=>"011101100",
  58390=>"100000011",
  58391=>"010111110",
  58392=>"101100001",
  58393=>"001001001",
  58394=>"000010101",
  58395=>"011001100",
  58396=>"011011011",
  58397=>"001100011",
  58398=>"100000100",
  58399=>"001100000",
  58400=>"100100101",
  58401=>"100100000",
  58402=>"001001000",
  58403=>"101101000",
  58404=>"011110110",
  58405=>"011111010",
  58406=>"010011011",
  58407=>"111011111",
  58408=>"111000100",
  58409=>"101111000",
  58410=>"101101100",
  58411=>"011010111",
  58412=>"001010011",
  58413=>"101010010",
  58414=>"100010001",
  58415=>"101001011",
  58416=>"111111001",
  58417=>"000011111",
  58418=>"111100101",
  58419=>"110010100",
  58420=>"110000000",
  58421=>"000111000",
  58422=>"101010100",
  58423=>"100110010",
  58424=>"001100111",
  58425=>"110101001",
  58426=>"100110011",
  58427=>"010101110",
  58428=>"000001100",
  58429=>"001001001",
  58430=>"111110000",
  58431=>"100001011",
  58432=>"111100001",
  58433=>"001000110",
  58434=>"101000000",
  58435=>"001011011",
  58436=>"100100111",
  58437=>"111111111",
  58438=>"101010100",
  58439=>"101000110",
  58440=>"001111011",
  58441=>"001001001",
  58442=>"001001000",
  58443=>"010011110",
  58444=>"000000101",
  58445=>"101011011",
  58446=>"001000100",
  58447=>"110000001",
  58448=>"100011000",
  58449=>"100000101",
  58450=>"001111111",
  58451=>"010110100",
  58452=>"100000000",
  58453=>"111101010",
  58454=>"010110101",
  58455=>"001011100",
  58456=>"111100010",
  58457=>"000111001",
  58458=>"000110111",
  58459=>"000001000",
  58460=>"001010000",
  58461=>"001010011",
  58462=>"000010000",
  58463=>"000011001",
  58464=>"000010010",
  58465=>"001010111",
  58466=>"000001111",
  58467=>"000100010",
  58468=>"100010011",
  58469=>"000010011",
  58470=>"101000010",
  58471=>"010010110",
  58472=>"111011011",
  58473=>"100110010",
  58474=>"011100000",
  58475=>"111100010",
  58476=>"000110001",
  58477=>"111001100",
  58478=>"110111010",
  58479=>"111101011",
  58480=>"000000011",
  58481=>"111100010",
  58482=>"101011111",
  58483=>"101000110",
  58484=>"111010011",
  58485=>"111011111",
  58486=>"001001010",
  58487=>"100011001",
  58488=>"000000100",
  58489=>"101111101",
  58490=>"000101110",
  58491=>"111000101",
  58492=>"101100101",
  58493=>"111101100",
  58494=>"011100111",
  58495=>"000101000",
  58496=>"000011001",
  58497=>"000011110",
  58498=>"000100101",
  58499=>"001100011",
  58500=>"010000001",
  58501=>"001101110",
  58502=>"100010000",
  58503=>"001011011",
  58504=>"100010110",
  58505=>"001010101",
  58506=>"101010010",
  58507=>"110001000",
  58508=>"111100010",
  58509=>"011001100",
  58510=>"010101110",
  58511=>"001111001",
  58512=>"111111100",
  58513=>"111100100",
  58514=>"100000111",
  58515=>"000011001",
  58516=>"101111010",
  58517=>"110010011",
  58518=>"001011111",
  58519=>"001001010",
  58520=>"010001111",
  58521=>"110000000",
  58522=>"010001111",
  58523=>"101000101",
  58524=>"010111101",
  58525=>"110110000",
  58526=>"101110001",
  58527=>"110001011",
  58528=>"110000000",
  58529=>"100011110",
  58530=>"001110000",
  58531=>"000110010",
  58532=>"110000110",
  58533=>"000110011",
  58534=>"101000000",
  58535=>"011101000",
  58536=>"101000001",
  58537=>"010001000",
  58538=>"110110100",
  58539=>"111101011",
  58540=>"010101100",
  58541=>"011010011",
  58542=>"000000111",
  58543=>"111000110",
  58544=>"001101011",
  58545=>"011110100",
  58546=>"000110110",
  58547=>"001100111",
  58548=>"101110101",
  58549=>"100010111",
  58550=>"001010000",
  58551=>"100000101",
  58552=>"110110111",
  58553=>"001001000",
  58554=>"000000101",
  58555=>"110100011",
  58556=>"111001100",
  58557=>"100101101",
  58558=>"001011010",
  58559=>"110001111",
  58560=>"000110001",
  58561=>"100110010",
  58562=>"001011000",
  58563=>"000011000",
  58564=>"111111000",
  58565=>"000111111",
  58566=>"001001000",
  58567=>"111000111",
  58568=>"101010000",
  58569=>"111010010",
  58570=>"100100111",
  58571=>"100111001",
  58572=>"111100010",
  58573=>"110010010",
  58574=>"001111001",
  58575=>"101000000",
  58576=>"011101100",
  58577=>"101001100",
  58578=>"000101101",
  58579=>"101110101",
  58580=>"100110100",
  58581=>"010101011",
  58582=>"100001100",
  58583=>"001010010",
  58584=>"010101001",
  58585=>"111110110",
  58586=>"010101100",
  58587=>"101110011",
  58588=>"110101010",
  58589=>"110001101",
  58590=>"010010110",
  58591=>"111011001",
  58592=>"011001111",
  58593=>"001011010",
  58594=>"010110111",
  58595=>"010001100",
  58596=>"100111000",
  58597=>"010100110",
  58598=>"000101101",
  58599=>"101101011",
  58600=>"111000110",
  58601=>"110011001",
  58602=>"000011110",
  58603=>"000101111",
  58604=>"010111011",
  58605=>"100100001",
  58606=>"000000100",
  58607=>"010101001",
  58608=>"000111111",
  58609=>"010010010",
  58610=>"000100001",
  58611=>"000101001",
  58612=>"100101001",
  58613=>"111100001",
  58614=>"000001100",
  58615=>"000110000",
  58616=>"001100001",
  58617=>"101010011",
  58618=>"100011000",
  58619=>"010011110",
  58620=>"000111100",
  58621=>"011110011",
  58622=>"111000001",
  58623=>"001110110",
  58624=>"111110101",
  58625=>"100110001",
  58626=>"010110101",
  58627=>"101011010",
  58628=>"000001111",
  58629=>"111001011",
  58630=>"101100011",
  58631=>"000111001",
  58632=>"001001101",
  58633=>"111010110",
  58634=>"111010110",
  58635=>"010011001",
  58636=>"110111001",
  58637=>"100001111",
  58638=>"011000000",
  58639=>"000100111",
  58640=>"100001000",
  58641=>"001101111",
  58642=>"111110101",
  58643=>"111110110",
  58644=>"000101101",
  58645=>"111000001",
  58646=>"100011101",
  58647=>"001011101",
  58648=>"110111100",
  58649=>"010000000",
  58650=>"001100011",
  58651=>"110101101",
  58652=>"001010000",
  58653=>"101000100",
  58654=>"011110001",
  58655=>"100000100",
  58656=>"000101100",
  58657=>"000001000",
  58658=>"101000010",
  58659=>"100011010",
  58660=>"001110100",
  58661=>"001110101",
  58662=>"101110010",
  58663=>"001110000",
  58664=>"010001001",
  58665=>"011001101",
  58666=>"001000111",
  58667=>"000010000",
  58668=>"111000100",
  58669=>"001011110",
  58670=>"011101001",
  58671=>"110000010",
  58672=>"001110100",
  58673=>"011001010",
  58674=>"000111110",
  58675=>"010010110",
  58676=>"010010100",
  58677=>"110110010",
  58678=>"011110110",
  58679=>"011011010",
  58680=>"000000001",
  58681=>"010010101",
  58682=>"101100101",
  58683=>"010010111",
  58684=>"101111010",
  58685=>"000001001",
  58686=>"100111011",
  58687=>"011111110",
  58688=>"011100101",
  58689=>"000000011",
  58690=>"011100000",
  58691=>"011001000",
  58692=>"111011011",
  58693=>"110000111",
  58694=>"000001001",
  58695=>"000011111",
  58696=>"000110001",
  58697=>"000101001",
  58698=>"110110100",
  58699=>"101111000",
  58700=>"100000001",
  58701=>"001101100",
  58702=>"101111110",
  58703=>"000110101",
  58704=>"011011100",
  58705=>"100010100",
  58706=>"101101011",
  58707=>"001111000",
  58708=>"011101100",
  58709=>"111100001",
  58710=>"001000000",
  58711=>"010101011",
  58712=>"100001000",
  58713=>"010000101",
  58714=>"001010001",
  58715=>"010010100",
  58716=>"101111111",
  58717=>"110010010",
  58718=>"111000000",
  58719=>"110101110",
  58720=>"000000010",
  58721=>"111100110",
  58722=>"001010100",
  58723=>"000000111",
  58724=>"101110111",
  58725=>"100000010",
  58726=>"100001010",
  58727=>"111111101",
  58728=>"100101100",
  58729=>"001000101",
  58730=>"101100001",
  58731=>"010010000",
  58732=>"001010011",
  58733=>"111001110",
  58734=>"000110011",
  58735=>"001000111",
  58736=>"011001101",
  58737=>"111100001",
  58738=>"101011011",
  58739=>"011001100",
  58740=>"000010010",
  58741=>"000011100",
  58742=>"100011011",
  58743=>"110111100",
  58744=>"000111110",
  58745=>"111100101",
  58746=>"101100110",
  58747=>"010110111",
  58748=>"100111111",
  58749=>"111011011",
  58750=>"001010000",
  58751=>"101000101",
  58752=>"111101010",
  58753=>"001000100",
  58754=>"010000011",
  58755=>"000110101",
  58756=>"001011011",
  58757=>"000101110",
  58758=>"011111011",
  58759=>"000111000",
  58760=>"100100110",
  58761=>"110101100",
  58762=>"100001111",
  58763=>"001000110",
  58764=>"000001100",
  58765=>"000010000",
  58766=>"010010000",
  58767=>"000101111",
  58768=>"100100100",
  58769=>"111010001",
  58770=>"001110000",
  58771=>"011100101",
  58772=>"011010100",
  58773=>"101111111",
  58774=>"111101010",
  58775=>"111010100",
  58776=>"010101000",
  58777=>"010101101",
  58778=>"001000101",
  58779=>"011011110",
  58780=>"010100100",
  58781=>"111100001",
  58782=>"010011001",
  58783=>"111111011",
  58784=>"000110000",
  58785=>"001000101",
  58786=>"001011110",
  58787=>"010000010",
  58788=>"001010000",
  58789=>"010001100",
  58790=>"000100110",
  58791=>"010000100",
  58792=>"011101101",
  58793=>"100011110",
  58794=>"100011000",
  58795=>"011100100",
  58796=>"000011000",
  58797=>"111011010",
  58798=>"111101001",
  58799=>"011110011",
  58800=>"000011110",
  58801=>"100001111",
  58802=>"000111101",
  58803=>"000000001",
  58804=>"111011000",
  58805=>"110100001",
  58806=>"100100000",
  58807=>"001000100",
  58808=>"000000101",
  58809=>"011100000",
  58810=>"000110100",
  58811=>"001010111",
  58812=>"000111100",
  58813=>"100011011",
  58814=>"001010110",
  58815=>"011110111",
  58816=>"101101001",
  58817=>"010111100",
  58818=>"100001011",
  58819=>"010101000",
  58820=>"000101000",
  58821=>"011011111",
  58822=>"100000110",
  58823=>"001101101",
  58824=>"010101000",
  58825=>"110111111",
  58826=>"011010110",
  58827=>"111100100",
  58828=>"010010101",
  58829=>"101001110",
  58830=>"100110100",
  58831=>"001101110",
  58832=>"011001110",
  58833=>"000100101",
  58834=>"101011001",
  58835=>"001101001",
  58836=>"000010101",
  58837=>"111111000",
  58838=>"111011001",
  58839=>"010010011",
  58840=>"110000000",
  58841=>"101001100",
  58842=>"111011010",
  58843=>"000110001",
  58844=>"100001000",
  58845=>"100011001",
  58846=>"110110011",
  58847=>"010110110",
  58848=>"111100010",
  58849=>"011100100",
  58850=>"111001101",
  58851=>"100010010",
  58852=>"011111010",
  58853=>"111111000",
  58854=>"010100010",
  58855=>"111000000",
  58856=>"000001111",
  58857=>"100010001",
  58858=>"000110000",
  58859=>"011110011",
  58860=>"000001000",
  58861=>"111101001",
  58862=>"010111000",
  58863=>"110011000",
  58864=>"100010110",
  58865=>"000001001",
  58866=>"110000100",
  58867=>"100101001",
  58868=>"011101100",
  58869=>"100101000",
  58870=>"010111011",
  58871=>"110101110",
  58872=>"011010001",
  58873=>"111001010",
  58874=>"010111110",
  58875=>"100111011",
  58876=>"000001010",
  58877=>"101001001",
  58878=>"010011010",
  58879=>"000001011",
  58880=>"010100011",
  58881=>"001110010",
  58882=>"101010100",
  58883=>"011000111",
  58884=>"001101000",
  58885=>"100000001",
  58886=>"100110111",
  58887=>"100010000",
  58888=>"000111111",
  58889=>"010101001",
  58890=>"100001111",
  58891=>"010011100",
  58892=>"101101000",
  58893=>"111101010",
  58894=>"111101010",
  58895=>"111001101",
  58896=>"101110011",
  58897=>"100010011",
  58898=>"101001100",
  58899=>"110011100",
  58900=>"010001111",
  58901=>"110110000",
  58902=>"110000101",
  58903=>"001100111",
  58904=>"110000111",
  58905=>"101001101",
  58906=>"101001000",
  58907=>"000000100",
  58908=>"100111101",
  58909=>"000000011",
  58910=>"010010101",
  58911=>"100000100",
  58912=>"010001011",
  58913=>"101000010",
  58914=>"000100101",
  58915=>"101101100",
  58916=>"110010111",
  58917=>"000001110",
  58918=>"011001010",
  58919=>"011101110",
  58920=>"011110000",
  58921=>"010011110",
  58922=>"111011000",
  58923=>"101011001",
  58924=>"010010111",
  58925=>"011100100",
  58926=>"000000001",
  58927=>"010111000",
  58928=>"010110101",
  58929=>"100111100",
  58930=>"011111101",
  58931=>"101001000",
  58932=>"101001100",
  58933=>"111111000",
  58934=>"011000001",
  58935=>"010010001",
  58936=>"111001011",
  58937=>"110100110",
  58938=>"001101010",
  58939=>"101000000",
  58940=>"110000101",
  58941=>"100001010",
  58942=>"100010100",
  58943=>"111000011",
  58944=>"111111110",
  58945=>"010010001",
  58946=>"110111000",
  58947=>"101001000",
  58948=>"010010000",
  58949=>"000000110",
  58950=>"000011000",
  58951=>"111010110",
  58952=>"110101000",
  58953=>"001000111",
  58954=>"100001110",
  58955=>"101101010",
  58956=>"101101110",
  58957=>"110101101",
  58958=>"111111101",
  58959=>"001101111",
  58960=>"101100011",
  58961=>"010000100",
  58962=>"001100011",
  58963=>"001100010",
  58964=>"110010001",
  58965=>"000100100",
  58966=>"100010000",
  58967=>"100100001",
  58968=>"011001001",
  58969=>"111000101",
  58970=>"110000000",
  58971=>"001010001",
  58972=>"001000100",
  58973=>"110011110",
  58974=>"001000000",
  58975=>"111001000",
  58976=>"111110101",
  58977=>"100000111",
  58978=>"011010100",
  58979=>"001011100",
  58980=>"001001101",
  58981=>"100000100",
  58982=>"000110000",
  58983=>"101001010",
  58984=>"000010011",
  58985=>"000100100",
  58986=>"010111110",
  58987=>"101111000",
  58988=>"000000011",
  58989=>"110111110",
  58990=>"011001101",
  58991=>"100001010",
  58992=>"011001001",
  58993=>"010000100",
  58994=>"001100100",
  58995=>"011011100",
  58996=>"101010101",
  58997=>"001110000",
  58998=>"001111100",
  58999=>"011001100",
  59000=>"010111001",
  59001=>"000010001",
  59002=>"100000110",
  59003=>"011100011",
  59004=>"101100100",
  59005=>"011011110",
  59006=>"010101111",
  59007=>"101111110",
  59008=>"101000111",
  59009=>"111100100",
  59010=>"110110100",
  59011=>"001000001",
  59012=>"000010111",
  59013=>"101000101",
  59014=>"101101011",
  59015=>"010001000",
  59016=>"101100011",
  59017=>"110000001",
  59018=>"110100111",
  59019=>"001100110",
  59020=>"100010101",
  59021=>"110111100",
  59022=>"101111100",
  59023=>"101110101",
  59024=>"100100101",
  59025=>"100011100",
  59026=>"111111111",
  59027=>"111110000",
  59028=>"000000001",
  59029=>"100100101",
  59030=>"000100111",
  59031=>"101111010",
  59032=>"101000000",
  59033=>"111110110",
  59034=>"110111000",
  59035=>"010100111",
  59036=>"101000011",
  59037=>"100100000",
  59038=>"101110001",
  59039=>"110111100",
  59040=>"001000000",
  59041=>"101000101",
  59042=>"001110111",
  59043=>"001110010",
  59044=>"100011101",
  59045=>"000100001",
  59046=>"010100110",
  59047=>"000010110",
  59048=>"011011110",
  59049=>"101110011",
  59050=>"111001010",
  59051=>"100000011",
  59052=>"000001111",
  59053=>"010011100",
  59054=>"010101010",
  59055=>"001000010",
  59056=>"000111011",
  59057=>"001010101",
  59058=>"110100101",
  59059=>"000001000",
  59060=>"001000110",
  59061=>"011100100",
  59062=>"001001011",
  59063=>"100110110",
  59064=>"011010000",
  59065=>"001111010",
  59066=>"101111110",
  59067=>"111111100",
  59068=>"001111111",
  59069=>"100100100",
  59070=>"011100100",
  59071=>"011001101",
  59072=>"110001100",
  59073=>"111001001",
  59074=>"100001110",
  59075=>"110100000",
  59076=>"000100011",
  59077=>"101101110",
  59078=>"110101011",
  59079=>"011111000",
  59080=>"011100101",
  59081=>"111011010",
  59082=>"110100111",
  59083=>"110001111",
  59084=>"000000100",
  59085=>"110110000",
  59086=>"110000101",
  59087=>"001101010",
  59088=>"100011010",
  59089=>"010000110",
  59090=>"100011101",
  59091=>"110100000",
  59092=>"111011100",
  59093=>"111100011",
  59094=>"101000101",
  59095=>"110111111",
  59096=>"000000001",
  59097=>"010111100",
  59098=>"000001000",
  59099=>"111011100",
  59100=>"001100000",
  59101=>"110010001",
  59102=>"111000100",
  59103=>"100101100",
  59104=>"001010110",
  59105=>"000000100",
  59106=>"001011010",
  59107=>"110010101",
  59108=>"000001100",
  59109=>"101001001",
  59110=>"010011010",
  59111=>"111010100",
  59112=>"100111101",
  59113=>"111011110",
  59114=>"010001011",
  59115=>"010010110",
  59116=>"000001010",
  59117=>"101111110",
  59118=>"111001100",
  59119=>"111011101",
  59120=>"111101110",
  59121=>"011011001",
  59122=>"110011111",
  59123=>"111010110",
  59124=>"100111111",
  59125=>"111101110",
  59126=>"001100110",
  59127=>"110100111",
  59128=>"110000011",
  59129=>"000101100",
  59130=>"010001001",
  59131=>"101001011",
  59132=>"110110000",
  59133=>"001100111",
  59134=>"011010010",
  59135=>"001011110",
  59136=>"001000010",
  59137=>"001011100",
  59138=>"100000110",
  59139=>"101001010",
  59140=>"000001010",
  59141=>"100000001",
  59142=>"000101110",
  59143=>"110100001",
  59144=>"011100001",
  59145=>"010100001",
  59146=>"010100000",
  59147=>"101010011",
  59148=>"000000101",
  59149=>"101011111",
  59150=>"000000110",
  59151=>"010000110",
  59152=>"010010000",
  59153=>"001000100",
  59154=>"100010010",
  59155=>"101111010",
  59156=>"001001010",
  59157=>"011110100",
  59158=>"110000000",
  59159=>"001001010",
  59160=>"110000010",
  59161=>"000001101",
  59162=>"111000010",
  59163=>"100001110",
  59164=>"001010000",
  59165=>"010111110",
  59166=>"100000001",
  59167=>"010000100",
  59168=>"010100111",
  59169=>"101111001",
  59170=>"101011011",
  59171=>"000110010",
  59172=>"010011001",
  59173=>"111101100",
  59174=>"010101101",
  59175=>"111111100",
  59176=>"000100110",
  59177=>"111000011",
  59178=>"011010010",
  59179=>"000101001",
  59180=>"011100001",
  59181=>"000111011",
  59182=>"111101100",
  59183=>"111110010",
  59184=>"000011110",
  59185=>"000010101",
  59186=>"101111000",
  59187=>"010011100",
  59188=>"100110010",
  59189=>"010000100",
  59190=>"100010100",
  59191=>"000000100",
  59192=>"001010010",
  59193=>"111110010",
  59194=>"010111000",
  59195=>"100001100",
  59196=>"111010011",
  59197=>"000000101",
  59198=>"000111101",
  59199=>"111011110",
  59200=>"010000111",
  59201=>"111001111",
  59202=>"011011110",
  59203=>"000011100",
  59204=>"111001101",
  59205=>"011101100",
  59206=>"001000100",
  59207=>"010101100",
  59208=>"001010011",
  59209=>"000111111",
  59210=>"000111111",
  59211=>"100010101",
  59212=>"000111010",
  59213=>"101110110",
  59214=>"001000011",
  59215=>"001011111",
  59216=>"110000010",
  59217=>"110111110",
  59218=>"011000011",
  59219=>"011010001",
  59220=>"111000001",
  59221=>"100000110",
  59222=>"001100000",
  59223=>"011010111",
  59224=>"001101001",
  59225=>"111111110",
  59226=>"111010010",
  59227=>"000010111",
  59228=>"101101001",
  59229=>"001000110",
  59230=>"011001010",
  59231=>"010110011",
  59232=>"111011000",
  59233=>"110011010",
  59234=>"001001000",
  59235=>"111011101",
  59236=>"101110010",
  59237=>"100110001",
  59238=>"001011010",
  59239=>"011001100",
  59240=>"001001111",
  59241=>"101001011",
  59242=>"100010110",
  59243=>"101110000",
  59244=>"110111000",
  59245=>"010101110",
  59246=>"101010101",
  59247=>"000100111",
  59248=>"010110111",
  59249=>"001011111",
  59250=>"110100111",
  59251=>"000010001",
  59252=>"001011110",
  59253=>"110000101",
  59254=>"000101010",
  59255=>"011000110",
  59256=>"100001000",
  59257=>"001000001",
  59258=>"000110011",
  59259=>"100011100",
  59260=>"000010000",
  59261=>"001000001",
  59262=>"110110111",
  59263=>"101110110",
  59264=>"010100100",
  59265=>"010001000",
  59266=>"110000100",
  59267=>"111000010",
  59268=>"111110111",
  59269=>"101001100",
  59270=>"010110000",
  59271=>"000101101",
  59272=>"011111101",
  59273=>"111111100",
  59274=>"010011010",
  59275=>"010100101",
  59276=>"001000011",
  59277=>"110011101",
  59278=>"100101001",
  59279=>"001000110",
  59280=>"010111101",
  59281=>"101010111",
  59282=>"011110110",
  59283=>"011011111",
  59284=>"000010111",
  59285=>"100011011",
  59286=>"010111001",
  59287=>"111001000",
  59288=>"000001101",
  59289=>"111000101",
  59290=>"001011111",
  59291=>"001101011",
  59292=>"010100000",
  59293=>"011001000",
  59294=>"100000000",
  59295=>"010011101",
  59296=>"111100101",
  59297=>"110100011",
  59298=>"110101101",
  59299=>"010011110",
  59300=>"001010110",
  59301=>"110000111",
  59302=>"001101100",
  59303=>"000001001",
  59304=>"010111001",
  59305=>"011110101",
  59306=>"100011110",
  59307=>"010101111",
  59308=>"000000111",
  59309=>"000110100",
  59310=>"111111110",
  59311=>"111100001",
  59312=>"010011101",
  59313=>"110101111",
  59314=>"000111100",
  59315=>"101001101",
  59316=>"111110100",
  59317=>"010000011",
  59318=>"011110111",
  59319=>"111101011",
  59320=>"110001101",
  59321=>"111000111",
  59322=>"110011010",
  59323=>"000011100",
  59324=>"011000110",
  59325=>"000101000",
  59326=>"000000000",
  59327=>"010000100",
  59328=>"000001101",
  59329=>"110111110",
  59330=>"100010110",
  59331=>"110010101",
  59332=>"011010001",
  59333=>"111110011",
  59334=>"011000001",
  59335=>"110110011",
  59336=>"000011011",
  59337=>"111000000",
  59338=>"010010111",
  59339=>"111000001",
  59340=>"111001011",
  59341=>"010001100",
  59342=>"010000010",
  59343=>"011010101",
  59344=>"100000010",
  59345=>"001111000",
  59346=>"011001110",
  59347=>"100011100",
  59348=>"111001110",
  59349=>"111010101",
  59350=>"010111011",
  59351=>"000100001",
  59352=>"000110111",
  59353=>"100110101",
  59354=>"010111001",
  59355=>"010100000",
  59356=>"111111001",
  59357=>"011110000",
  59358=>"111010111",
  59359=>"111100011",
  59360=>"001101100",
  59361=>"001011001",
  59362=>"000010110",
  59363=>"000000000",
  59364=>"110010100",
  59365=>"111110111",
  59366=>"110000011",
  59367=>"010110010",
  59368=>"000101011",
  59369=>"101011010",
  59370=>"111000110",
  59371=>"001110111",
  59372=>"110111010",
  59373=>"001011111",
  59374=>"010111000",
  59375=>"100010001",
  59376=>"001101111",
  59377=>"011100110",
  59378=>"101001011",
  59379=>"100010100",
  59380=>"100111011",
  59381=>"010111000",
  59382=>"010101110",
  59383=>"010100111",
  59384=>"000000001",
  59385=>"011000010",
  59386=>"010011100",
  59387=>"100010111",
  59388=>"100110010",
  59389=>"101000100",
  59390=>"011000001",
  59391=>"101010111",
  59392=>"101011100",
  59393=>"100111110",
  59394=>"000010100",
  59395=>"000100000",
  59396=>"001010111",
  59397=>"001110110",
  59398=>"001111010",
  59399=>"010111000",
  59400=>"111100000",
  59401=>"111101010",
  59402=>"011011100",
  59403=>"000010100",
  59404=>"011011001",
  59405=>"101111100",
  59406=>"110110010",
  59407=>"011001010",
  59408=>"010100101",
  59409=>"001001101",
  59410=>"011000101",
  59411=>"010111110",
  59412=>"100110111",
  59413=>"000011111",
  59414=>"010100011",
  59415=>"110011010",
  59416=>"110101101",
  59417=>"010000111",
  59418=>"100000100",
  59419=>"110101001",
  59420=>"110000010",
  59421=>"100110000",
  59422=>"100111110",
  59423=>"010000010",
  59424=>"110100101",
  59425=>"101000100",
  59426=>"011101010",
  59427=>"001111100",
  59428=>"000101100",
  59429=>"010000011",
  59430=>"011101011",
  59431=>"010111111",
  59432=>"111111011",
  59433=>"001101111",
  59434=>"001001010",
  59435=>"001000001",
  59436=>"011010010",
  59437=>"100110110",
  59438=>"100010101",
  59439=>"000001010",
  59440=>"010101100",
  59441=>"110000000",
  59442=>"111111111",
  59443=>"101000010",
  59444=>"010110101",
  59445=>"100001110",
  59446=>"110100011",
  59447=>"001100100",
  59448=>"010001011",
  59449=>"011101010",
  59450=>"111000011",
  59451=>"110011111",
  59452=>"001100000",
  59453=>"011001011",
  59454=>"111010110",
  59455=>"001001101",
  59456=>"111000100",
  59457=>"111001011",
  59458=>"100111000",
  59459=>"010100010",
  59460=>"001110100",
  59461=>"101001110",
  59462=>"001001100",
  59463=>"111100001",
  59464=>"111110111",
  59465=>"000100111",
  59466=>"111100100",
  59467=>"000100101",
  59468=>"110001100",
  59469=>"000110011",
  59470=>"110111010",
  59471=>"110010110",
  59472=>"111111111",
  59473=>"000011011",
  59474=>"000111100",
  59475=>"100010110",
  59476=>"101011000",
  59477=>"010100011",
  59478=>"100000100",
  59479=>"111110000",
  59480=>"000010010",
  59481=>"111100110",
  59482=>"101111001",
  59483=>"111010000",
  59484=>"010100111",
  59485=>"101001101",
  59486=>"111010010",
  59487=>"101111010",
  59488=>"000001101",
  59489=>"010010000",
  59490=>"101010000",
  59491=>"101110100",
  59492=>"110000101",
  59493=>"110100110",
  59494=>"010001101",
  59495=>"011000011",
  59496=>"101010010",
  59497=>"110111010",
  59498=>"010110000",
  59499=>"100110000",
  59500=>"010101100",
  59501=>"100010000",
  59502=>"110011000",
  59503=>"011010111",
  59504=>"110111010",
  59505=>"011000011",
  59506=>"111110000",
  59507=>"000001100",
  59508=>"001101110",
  59509=>"011100110",
  59510=>"100011000",
  59511=>"000010001",
  59512=>"000001011",
  59513=>"011000011",
  59514=>"110111000",
  59515=>"011011001",
  59516=>"001110101",
  59517=>"101100110",
  59518=>"111000101",
  59519=>"100100001",
  59520=>"110100011",
  59521=>"010000111",
  59522=>"100110100",
  59523=>"111110000",
  59524=>"111110000",
  59525=>"111000100",
  59526=>"111011011",
  59527=>"010101000",
  59528=>"000100100",
  59529=>"110110100",
  59530=>"101101000",
  59531=>"110100000",
  59532=>"100110001",
  59533=>"010000001",
  59534=>"000010011",
  59535=>"001010111",
  59536=>"110001111",
  59537=>"111101111",
  59538=>"010011010",
  59539=>"110000010",
  59540=>"010110000",
  59541=>"000101101",
  59542=>"111101001",
  59543=>"010010110",
  59544=>"010011110",
  59545=>"000111001",
  59546=>"010011011",
  59547=>"100001111",
  59548=>"000001110",
  59549=>"001011000",
  59550=>"111010011",
  59551=>"010111101",
  59552=>"011100101",
  59553=>"011011001",
  59554=>"011111011",
  59555=>"001111111",
  59556=>"010000001",
  59557=>"011010110",
  59558=>"111010011",
  59559=>"111110000",
  59560=>"011000100",
  59561=>"011010000",
  59562=>"000001010",
  59563=>"101100001",
  59564=>"100010000",
  59565=>"100010000",
  59566=>"100010000",
  59567=>"101101000",
  59568=>"110101100",
  59569=>"011110010",
  59570=>"000011001",
  59571=>"010001001",
  59572=>"101000001",
  59573=>"001111010",
  59574=>"101100101",
  59575=>"010010111",
  59576=>"110000111",
  59577=>"001100010",
  59578=>"100111011",
  59579=>"100101110",
  59580=>"000010011",
  59581=>"110111010",
  59582=>"110100000",
  59583=>"010011100",
  59584=>"101101001",
  59585=>"101101011",
  59586=>"101101010",
  59587=>"111101101",
  59588=>"101011011",
  59589=>"011100101",
  59590=>"000111010",
  59591=>"000010010",
  59592=>"000000100",
  59593=>"011101001",
  59594=>"000000010",
  59595=>"011110110",
  59596=>"111011111",
  59597=>"111000101",
  59598=>"001000000",
  59599=>"011111101",
  59600=>"010111101",
  59601=>"011011100",
  59602=>"010000001",
  59603=>"011011111",
  59604=>"111101001",
  59605=>"100111000",
  59606=>"010111111",
  59607=>"110100000",
  59608=>"001100100",
  59609=>"100100001",
  59610=>"001100111",
  59611=>"100001001",
  59612=>"111111110",
  59613=>"010110100",
  59614=>"100010100",
  59615=>"010000100",
  59616=>"101101100",
  59617=>"010010110",
  59618=>"100010110",
  59619=>"011101011",
  59620=>"011110111",
  59621=>"100101010",
  59622=>"001010000",
  59623=>"111111001",
  59624=>"110000010",
  59625=>"001110101",
  59626=>"010100101",
  59627=>"000101100",
  59628=>"010100001",
  59629=>"110101101",
  59630=>"000001001",
  59631=>"000100111",
  59632=>"100111010",
  59633=>"011011010",
  59634=>"101001110",
  59635=>"001100100",
  59636=>"111011110",
  59637=>"010110001",
  59638=>"101110101",
  59639=>"001010001",
  59640=>"011101111",
  59641=>"010110001",
  59642=>"000000010",
  59643=>"101110000",
  59644=>"011010100",
  59645=>"111110001",
  59646=>"111101001",
  59647=>"000101011",
  59648=>"101101101",
  59649=>"100110011",
  59650=>"011101011",
  59651=>"111100100",
  59652=>"011111101",
  59653=>"110010000",
  59654=>"110111100",
  59655=>"111011100",
  59656=>"000000111",
  59657=>"100001011",
  59658=>"001000001",
  59659=>"010100011",
  59660=>"011101101",
  59661=>"101000110",
  59662=>"001000011",
  59663=>"001000000",
  59664=>"011001110",
  59665=>"100010011",
  59666=>"111110100",
  59667=>"101010110",
  59668=>"111110010",
  59669=>"000000111",
  59670=>"111101000",
  59671=>"000110011",
  59672=>"111100100",
  59673=>"111100101",
  59674=>"001100101",
  59675=>"111111011",
  59676=>"001000001",
  59677=>"111000000",
  59678=>"001100111",
  59679=>"111001000",
  59680=>"111000000",
  59681=>"111010110",
  59682=>"011010101",
  59683=>"110001100",
  59684=>"001010001",
  59685=>"000100000",
  59686=>"011000001",
  59687=>"101100110",
  59688=>"010100001",
  59689=>"111011100",
  59690=>"001111110",
  59691=>"111011010",
  59692=>"111000110",
  59693=>"010110010",
  59694=>"111111001",
  59695=>"100001000",
  59696=>"010001010",
  59697=>"111101001",
  59698=>"100000100",
  59699=>"011100001",
  59700=>"010000110",
  59701=>"101110100",
  59702=>"011101101",
  59703=>"000111110",
  59704=>"011000001",
  59705=>"111100001",
  59706=>"010111011",
  59707=>"100100111",
  59708=>"111001010",
  59709=>"001100110",
  59710=>"001011010",
  59711=>"010100100",
  59712=>"101001000",
  59713=>"110110110",
  59714=>"111011001",
  59715=>"101101100",
  59716=>"000101101",
  59717=>"110100111",
  59718=>"111110000",
  59719=>"000011111",
  59720=>"101001000",
  59721=>"001111110",
  59722=>"101011001",
  59723=>"011110010",
  59724=>"010010011",
  59725=>"011011111",
  59726=>"000100010",
  59727=>"001100110",
  59728=>"000011110",
  59729=>"110000110",
  59730=>"000011001",
  59731=>"000101110",
  59732=>"110111010",
  59733=>"011010100",
  59734=>"101010011",
  59735=>"001100100",
  59736=>"101101111",
  59737=>"101000010",
  59738=>"001000100",
  59739=>"011011010",
  59740=>"101100001",
  59741=>"000111101",
  59742=>"100001111",
  59743=>"111011001",
  59744=>"110101001",
  59745=>"110110110",
  59746=>"111111001",
  59747=>"110110010",
  59748=>"100101100",
  59749=>"001000000",
  59750=>"011100100",
  59751=>"111101000",
  59752=>"100101111",
  59753=>"001011100",
  59754=>"000001111",
  59755=>"110010011",
  59756=>"111011000",
  59757=>"100101001",
  59758=>"111111101",
  59759=>"010011110",
  59760=>"001001111",
  59761=>"010110100",
  59762=>"001011110",
  59763=>"000110010",
  59764=>"010010011",
  59765=>"100010000",
  59766=>"101100101",
  59767=>"011110110",
  59768=>"000001101",
  59769=>"010000111",
  59770=>"111000010",
  59771=>"111011011",
  59772=>"000111111",
  59773=>"011111001",
  59774=>"111000100",
  59775=>"001000001",
  59776=>"101000111",
  59777=>"100001100",
  59778=>"000110010",
  59779=>"011110010",
  59780=>"110111111",
  59781=>"010110100",
  59782=>"111101000",
  59783=>"010000001",
  59784=>"101010001",
  59785=>"101101010",
  59786=>"010001001",
  59787=>"010111110",
  59788=>"101011110",
  59789=>"111111000",
  59790=>"100110011",
  59791=>"000010110",
  59792=>"111010110",
  59793=>"111011001",
  59794=>"111011001",
  59795=>"100010100",
  59796=>"011010110",
  59797=>"101010110",
  59798=>"000100000",
  59799=>"100100010",
  59800=>"000000110",
  59801=>"101100000",
  59802=>"010100001",
  59803=>"011111110",
  59804=>"011010011",
  59805=>"011101101",
  59806=>"000011101",
  59807=>"001110011",
  59808=>"100010000",
  59809=>"011000000",
  59810=>"011110111",
  59811=>"111000101",
  59812=>"011001100",
  59813=>"101101010",
  59814=>"100011110",
  59815=>"100100111",
  59816=>"001111011",
  59817=>"101111001",
  59818=>"010010001",
  59819=>"110001101",
  59820=>"001001111",
  59821=>"111100101",
  59822=>"110001100",
  59823=>"101111001",
  59824=>"101101111",
  59825=>"101000011",
  59826=>"110001110",
  59827=>"101011011",
  59828=>"101101011",
  59829=>"110000110",
  59830=>"100010010",
  59831=>"011010100",
  59832=>"000101011",
  59833=>"000100001",
  59834=>"010000010",
  59835=>"100001000",
  59836=>"110001011",
  59837=>"110001111",
  59838=>"010000001",
  59839=>"011000111",
  59840=>"001011001",
  59841=>"011110101",
  59842=>"101100111",
  59843=>"000111001",
  59844=>"111001011",
  59845=>"111110000",
  59846=>"110111111",
  59847=>"011011100",
  59848=>"110001000",
  59849=>"010111111",
  59850=>"000100001",
  59851=>"000001100",
  59852=>"000001101",
  59853=>"110101110",
  59854=>"101011011",
  59855=>"011111000",
  59856=>"001111011",
  59857=>"001011010",
  59858=>"000000110",
  59859=>"000000110",
  59860=>"101000001",
  59861=>"101011001",
  59862=>"111101001",
  59863=>"111000110",
  59864=>"010111010",
  59865=>"100100001",
  59866=>"010001010",
  59867=>"011010101",
  59868=>"101000110",
  59869=>"001101010",
  59870=>"011010101",
  59871=>"000010010",
  59872=>"011110110",
  59873=>"111111010",
  59874=>"011111000",
  59875=>"100101111",
  59876=>"010001111",
  59877=>"101110000",
  59878=>"101111100",
  59879=>"101001011",
  59880=>"011000111",
  59881=>"010110011",
  59882=>"100100110",
  59883=>"011001001",
  59884=>"011101010",
  59885=>"101001101",
  59886=>"000010010",
  59887=>"111101001",
  59888=>"001010000",
  59889=>"111101100",
  59890=>"000100010",
  59891=>"100101111",
  59892=>"101001111",
  59893=>"110110001",
  59894=>"010111110",
  59895=>"101001001",
  59896=>"101110110",
  59897=>"011001110",
  59898=>"011100010",
  59899=>"011010100",
  59900=>"100010110",
  59901=>"011101111",
  59902=>"111000101",
  59903=>"010010010",
  59904=>"111100110",
  59905=>"101111011",
  59906=>"111001110",
  59907=>"101010010",
  59908=>"101100011",
  59909=>"001111001",
  59910=>"100110100",
  59911=>"111000000",
  59912=>"010110001",
  59913=>"000100000",
  59914=>"000101100",
  59915=>"000110111",
  59916=>"000000001",
  59917=>"100010010",
  59918=>"001000111",
  59919=>"110110101",
  59920=>"001101101",
  59921=>"011111111",
  59922=>"100000110",
  59923=>"100100001",
  59924=>"111100010",
  59925=>"101011001",
  59926=>"001100101",
  59927=>"010100111",
  59928=>"100010111",
  59929=>"101111100",
  59930=>"111010100",
  59931=>"000110001",
  59932=>"011001000",
  59933=>"110000111",
  59934=>"111111011",
  59935=>"011001010",
  59936=>"111011010",
  59937=>"101100000",
  59938=>"100110101",
  59939=>"110100001",
  59940=>"111110100",
  59941=>"100001010",
  59942=>"111110000",
  59943=>"011011100",
  59944=>"010011111",
  59945=>"000111010",
  59946=>"011100001",
  59947=>"001001111",
  59948=>"010101111",
  59949=>"111101111",
  59950=>"000111110",
  59951=>"110011111",
  59952=>"001010110",
  59953=>"110011011",
  59954=>"101111100",
  59955=>"110000100",
  59956=>"100001111",
  59957=>"110010010",
  59958=>"011000110",
  59959=>"111001110",
  59960=>"001111110",
  59961=>"000101010",
  59962=>"001100111",
  59963=>"010010100",
  59964=>"000100001",
  59965=>"100010011",
  59966=>"100000111",
  59967=>"110000010",
  59968=>"111011011",
  59969=>"010111010",
  59970=>"011001011",
  59971=>"111000000",
  59972=>"011011111",
  59973=>"010010001",
  59974=>"000011010",
  59975=>"111111111",
  59976=>"111011101",
  59977=>"111100110",
  59978=>"110011011",
  59979=>"001111101",
  59980=>"010010100",
  59981=>"100101001",
  59982=>"110110010",
  59983=>"000010100",
  59984=>"110011011",
  59985=>"010101001",
  59986=>"011101001",
  59987=>"011011110",
  59988=>"000000001",
  59989=>"001110001",
  59990=>"110101010",
  59991=>"111001110",
  59992=>"000101100",
  59993=>"000001010",
  59994=>"101001011",
  59995=>"111101100",
  59996=>"011111111",
  59997=>"001101000",
  59998=>"001101100",
  59999=>"010011101",
  60000=>"001011101",
  60001=>"111100001",
  60002=>"111111010",
  60003=>"010011010",
  60004=>"011010111",
  60005=>"101111110",
  60006=>"110011100",
  60007=>"000000001",
  60008=>"010010000",
  60009=>"011110101",
  60010=>"010110001",
  60011=>"000001101",
  60012=>"001011101",
  60013=>"001000100",
  60014=>"001010000",
  60015=>"010111100",
  60016=>"101001010",
  60017=>"111110100",
  60018=>"110111011",
  60019=>"111000010",
  60020=>"011001001",
  60021=>"110100000",
  60022=>"111110111",
  60023=>"101000011",
  60024=>"011000001",
  60025=>"101101111",
  60026=>"001111010",
  60027=>"000111111",
  60028=>"100110010",
  60029=>"100100000",
  60030=>"000000000",
  60031=>"110100111",
  60032=>"101000011",
  60033=>"101100101",
  60034=>"011011011",
  60035=>"011010010",
  60036=>"001010010",
  60037=>"001010101",
  60038=>"111000010",
  60039=>"111110110",
  60040=>"111100101",
  60041=>"111011101",
  60042=>"000000011",
  60043=>"011110011",
  60044=>"001110111",
  60045=>"010011001",
  60046=>"111110011",
  60047=>"110010010",
  60048=>"111100100",
  60049=>"011111001",
  60050=>"000000111",
  60051=>"111111101",
  60052=>"111010101",
  60053=>"011000100",
  60054=>"101111000",
  60055=>"011110110",
  60056=>"001010100",
  60057=>"011101111",
  60058=>"011110000",
  60059=>"101100110",
  60060=>"100111000",
  60061=>"011011011",
  60062=>"010100100",
  60063=>"011010011",
  60064=>"000011001",
  60065=>"000001100",
  60066=>"011101001",
  60067=>"110111111",
  60068=>"011001001",
  60069=>"001111101",
  60070=>"111000011",
  60071=>"011100100",
  60072=>"111010001",
  60073=>"001010110",
  60074=>"000011100",
  60075=>"101110000",
  60076=>"100111010",
  60077=>"110000101",
  60078=>"100110110",
  60079=>"111001101",
  60080=>"111101111",
  60081=>"000000010",
  60082=>"111110011",
  60083=>"011000111",
  60084=>"101010110",
  60085=>"000011000",
  60086=>"010111011",
  60087=>"011100010",
  60088=>"110000001",
  60089=>"000010100",
  60090=>"011000111",
  60091=>"001101101",
  60092=>"110000100",
  60093=>"011001001",
  60094=>"100000001",
  60095=>"101100100",
  60096=>"001001111",
  60097=>"010110100",
  60098=>"000111101",
  60099=>"010111001",
  60100=>"110000100",
  60101=>"110101011",
  60102=>"111011100",
  60103=>"000000101",
  60104=>"011011111",
  60105=>"111010110",
  60106=>"011110110",
  60107=>"110110100",
  60108=>"011100000",
  60109=>"101110100",
  60110=>"000001101",
  60111=>"001001111",
  60112=>"100101100",
  60113=>"111101110",
  60114=>"111111001",
  60115=>"001110000",
  60116=>"100001100",
  60117=>"001010000",
  60118=>"111111010",
  60119=>"101010001",
  60120=>"011001011",
  60121=>"100100110",
  60122=>"111001101",
  60123=>"110001010",
  60124=>"011100010",
  60125=>"111100000",
  60126=>"000010000",
  60127=>"001100001",
  60128=>"011000011",
  60129=>"100110111",
  60130=>"000000010",
  60131=>"101010001",
  60132=>"010011001",
  60133=>"011011010",
  60134=>"011000111",
  60135=>"010100001",
  60136=>"000001000",
  60137=>"111110101",
  60138=>"100100101",
  60139=>"100011101",
  60140=>"100000010",
  60141=>"110001111",
  60142=>"000010110",
  60143=>"001011111",
  60144=>"101111101",
  60145=>"000001001",
  60146=>"110110000",
  60147=>"011000100",
  60148=>"000110001",
  60149=>"100010000",
  60150=>"110110110",
  60151=>"011000101",
  60152=>"001000010",
  60153=>"001111011",
  60154=>"010010100",
  60155=>"110101101",
  60156=>"110011101",
  60157=>"000101011",
  60158=>"001010000",
  60159=>"011001101",
  60160=>"101011010",
  60161=>"000111001",
  60162=>"110001000",
  60163=>"101001000",
  60164=>"100101000",
  60165=>"011100011",
  60166=>"001000011",
  60167=>"011101111",
  60168=>"101100001",
  60169=>"111111110",
  60170=>"110011001",
  60171=>"011100000",
  60172=>"100101011",
  60173=>"110101110",
  60174=>"110010000",
  60175=>"000101111",
  60176=>"100000101",
  60177=>"001011011",
  60178=>"010101011",
  60179=>"111110000",
  60180=>"110110111",
  60181=>"001011001",
  60182=>"111111100",
  60183=>"111000011",
  60184=>"111101011",
  60185=>"000111110",
  60186=>"000000111",
  60187=>"100100110",
  60188=>"000000000",
  60189=>"000011110",
  60190=>"000100000",
  60191=>"111000000",
  60192=>"111011010",
  60193=>"010011011",
  60194=>"111010010",
  60195=>"001000101",
  60196=>"001000001",
  60197=>"011111110",
  60198=>"111010000",
  60199=>"010000111",
  60200=>"011011000",
  60201=>"101011100",
  60202=>"011010111",
  60203=>"110111110",
  60204=>"001101101",
  60205=>"100001010",
  60206=>"000110001",
  60207=>"101101010",
  60208=>"000001100",
  60209=>"000111111",
  60210=>"110111100",
  60211=>"010000101",
  60212=>"111100010",
  60213=>"111010010",
  60214=>"110001111",
  60215=>"110100000",
  60216=>"000101110",
  60217=>"111111011",
  60218=>"001111000",
  60219=>"001111100",
  60220=>"011100101",
  60221=>"101001100",
  60222=>"111111001",
  60223=>"000011111",
  60224=>"010100101",
  60225=>"000111111",
  60226=>"000001011",
  60227=>"100100101",
  60228=>"010011010",
  60229=>"000110010",
  60230=>"011001111",
  60231=>"110011111",
  60232=>"000000101",
  60233=>"110011101",
  60234=>"010100111",
  60235=>"001111000",
  60236=>"011000011",
  60237=>"100100011",
  60238=>"000011100",
  60239=>"111011110",
  60240=>"001100010",
  60241=>"010100000",
  60242=>"011100001",
  60243=>"000000000",
  60244=>"101101101",
  60245=>"010010010",
  60246=>"000111101",
  60247=>"110011000",
  60248=>"011110100",
  60249=>"000011100",
  60250=>"010110011",
  60251=>"101001100",
  60252=>"111101001",
  60253=>"110000111",
  60254=>"011011010",
  60255=>"011101001",
  60256=>"001100001",
  60257=>"011100011",
  60258=>"001010111",
  60259=>"000101011",
  60260=>"110001010",
  60261=>"101000110",
  60262=>"111011000",
  60263=>"100100100",
  60264=>"111110011",
  60265=>"011000010",
  60266=>"011011000",
  60267=>"100110101",
  60268=>"101110001",
  60269=>"111011110",
  60270=>"100110011",
  60271=>"000101101",
  60272=>"101100000",
  60273=>"001011111",
  60274=>"011011011",
  60275=>"101001010",
  60276=>"110001110",
  60277=>"100000110",
  60278=>"000111001",
  60279=>"011000101",
  60280=>"000111101",
  60281=>"000110110",
  60282=>"011110001",
  60283=>"011010110",
  60284=>"000111000",
  60285=>"110100010",
  60286=>"000101111",
  60287=>"100111010",
  60288=>"010000101",
  60289=>"100111110",
  60290=>"111100001",
  60291=>"101101000",
  60292=>"100011111",
  60293=>"010010001",
  60294=>"101011010",
  60295=>"101100110",
  60296=>"111111000",
  60297=>"100110000",
  60298=>"000000001",
  60299=>"011001001",
  60300=>"101100001",
  60301=>"110111011",
  60302=>"011101000",
  60303=>"010000100",
  60304=>"001110001",
  60305=>"111110110",
  60306=>"101100000",
  60307=>"101100001",
  60308=>"101000100",
  60309=>"110010111",
  60310=>"011111111",
  60311=>"101010000",
  60312=>"101111100",
  60313=>"010001011",
  60314=>"001101011",
  60315=>"010100010",
  60316=>"000000000",
  60317=>"010001111",
  60318=>"100000000",
  60319=>"110111000",
  60320=>"111111111",
  60321=>"110110101",
  60322=>"111011010",
  60323=>"111000111",
  60324=>"011111100",
  60325=>"110010110",
  60326=>"001010011",
  60327=>"010100111",
  60328=>"001101011",
  60329=>"000101011",
  60330=>"111000100",
  60331=>"010001000",
  60332=>"101110001",
  60333=>"000100000",
  60334=>"100000100",
  60335=>"000001000",
  60336=>"001110011",
  60337=>"011111101",
  60338=>"110000101",
  60339=>"011100001",
  60340=>"100111101",
  60341=>"011011011",
  60342=>"100101110",
  60343=>"100001110",
  60344=>"000010011",
  60345=>"000011000",
  60346=>"000011101",
  60347=>"011001101",
  60348=>"101111100",
  60349=>"000011101",
  60350=>"011111001",
  60351=>"010110010",
  60352=>"001001010",
  60353=>"010011001",
  60354=>"101001000",
  60355=>"111011100",
  60356=>"010101100",
  60357=>"101010001",
  60358=>"100100100",
  60359=>"010100100",
  60360=>"000110000",
  60361=>"011010000",
  60362=>"000010101",
  60363=>"001110001",
  60364=>"000000001",
  60365=>"000000110",
  60366=>"100100100",
  60367=>"111110000",
  60368=>"000000001",
  60369=>"101101010",
  60370=>"100000110",
  60371=>"100010111",
  60372=>"001011111",
  60373=>"101110101",
  60374=>"110111010",
  60375=>"011101111",
  60376=>"000000101",
  60377=>"001110110",
  60378=>"110111100",
  60379=>"001010001",
  60380=>"101001111",
  60381=>"010010000",
  60382=>"110001011",
  60383=>"111011111",
  60384=>"011100101",
  60385=>"010011111",
  60386=>"101100111",
  60387=>"011011101",
  60388=>"000010011",
  60389=>"111101010",
  60390=>"110001000",
  60391=>"101110111",
  60392=>"011111110",
  60393=>"110111100",
  60394=>"001101110",
  60395=>"111011111",
  60396=>"100110111",
  60397=>"111110010",
  60398=>"100111100",
  60399=>"110011101",
  60400=>"110001111",
  60401=>"101011011",
  60402=>"100011100",
  60403=>"011100011",
  60404=>"110101000",
  60405=>"111100110",
  60406=>"110001010",
  60407=>"100010001",
  60408=>"110110101",
  60409=>"100110110",
  60410=>"101100111",
  60411=>"111100000",
  60412=>"111011111",
  60413=>"110100101",
  60414=>"111100011",
  60415=>"101111001",
  60416=>"010011110",
  60417=>"000011010",
  60418=>"110010000",
  60419=>"110010100",
  60420=>"001101101",
  60421=>"010110001",
  60422=>"001110110",
  60423=>"001001110",
  60424=>"000010000",
  60425=>"100010101",
  60426=>"001100010",
  60427=>"111000001",
  60428=>"100101111",
  60429=>"011000110",
  60430=>"111110111",
  60431=>"100101111",
  60432=>"111001001",
  60433=>"100110111",
  60434=>"011111100",
  60435=>"101111100",
  60436=>"011101000",
  60437=>"110011010",
  60438=>"011001011",
  60439=>"101011100",
  60440=>"000111101",
  60441=>"000111110",
  60442=>"000100101",
  60443=>"001100101",
  60444=>"110000101",
  60445=>"111010011",
  60446=>"100010001",
  60447=>"100110101",
  60448=>"111010010",
  60449=>"110010000",
  60450=>"110000100",
  60451=>"010110100",
  60452=>"001111100",
  60453=>"010000101",
  60454=>"011001111",
  60455=>"111000100",
  60456=>"010101011",
  60457=>"101011110",
  60458=>"100001100",
  60459=>"100110010",
  60460=>"110100101",
  60461=>"001101100",
  60462=>"111111111",
  60463=>"100011010",
  60464=>"101010100",
  60465=>"110000101",
  60466=>"111011011",
  60467=>"100011111",
  60468=>"111111110",
  60469=>"000011101",
  60470=>"100100001",
  60471=>"101111010",
  60472=>"111010010",
  60473=>"010110101",
  60474=>"011110110",
  60475=>"001111011",
  60476=>"000100110",
  60477=>"011110110",
  60478=>"110010001",
  60479=>"111110110",
  60480=>"000010010",
  60481=>"000101111",
  60482=>"111100111",
  60483=>"000111000",
  60484=>"001010000",
  60485=>"001010001",
  60486=>"010000100",
  60487=>"110100100",
  60488=>"110010000",
  60489=>"110010101",
  60490=>"110100100",
  60491=>"011001111",
  60492=>"001011101",
  60493=>"011001101",
  60494=>"101001111",
  60495=>"011111100",
  60496=>"001101110",
  60497=>"011111111",
  60498=>"001000000",
  60499=>"110000111",
  60500=>"100000001",
  60501=>"000010111",
  60502=>"001011000",
  60503=>"101111010",
  60504=>"000101000",
  60505=>"000100100",
  60506=>"010111000",
  60507=>"100010011",
  60508=>"010010010",
  60509=>"101111110",
  60510=>"110111010",
  60511=>"001001010",
  60512=>"100101000",
  60513=>"101001100",
  60514=>"011111010",
  60515=>"101110000",
  60516=>"100000101",
  60517=>"011011000",
  60518=>"000011010",
  60519=>"111110110",
  60520=>"110000010",
  60521=>"100000110",
  60522=>"001101011",
  60523=>"001111001",
  60524=>"001100111",
  60525=>"100111110",
  60526=>"100010000",
  60527=>"111011000",
  60528=>"000111011",
  60529=>"001101110",
  60530=>"111000110",
  60531=>"101011000",
  60532=>"000101001",
  60533=>"010000010",
  60534=>"010001101",
  60535=>"011111110",
  60536=>"000101010",
  60537=>"010011100",
  60538=>"010010100",
  60539=>"001100110",
  60540=>"000101011",
  60541=>"111100001",
  60542=>"001011000",
  60543=>"011101110",
  60544=>"110011111",
  60545=>"010100011",
  60546=>"011001011",
  60547=>"011001111",
  60548=>"100001110",
  60549=>"101101011",
  60550=>"000101110",
  60551=>"111010000",
  60552=>"010110001",
  60553=>"011111001",
  60554=>"101110100",
  60555=>"110010001",
  60556=>"001010111",
  60557=>"111111011",
  60558=>"101100011",
  60559=>"010000011",
  60560=>"110100011",
  60561=>"110111001",
  60562=>"101010101",
  60563=>"101010100",
  60564=>"111011110",
  60565=>"100111110",
  60566=>"001011101",
  60567=>"100011101",
  60568=>"111101011",
  60569=>"000111011",
  60570=>"001101101",
  60571=>"011011001",
  60572=>"010111110",
  60573=>"011110000",
  60574=>"000110011",
  60575=>"100100110",
  60576=>"011100100",
  60577=>"110111010",
  60578=>"110010101",
  60579=>"000010001",
  60580=>"111110011",
  60581=>"100010000",
  60582=>"000001101",
  60583=>"110000011",
  60584=>"001110010",
  60585=>"101111010",
  60586=>"001100011",
  60587=>"001111110",
  60588=>"010100111",
  60589=>"111111111",
  60590=>"011010111",
  60591=>"010100010",
  60592=>"111100000",
  60593=>"011110011",
  60594=>"011011011",
  60595=>"000111010",
  60596=>"110111011",
  60597=>"101011011",
  60598=>"000110000",
  60599=>"001101101",
  60600=>"101111101",
  60601=>"000010100",
  60602=>"010101110",
  60603=>"100111010",
  60604=>"000101010",
  60605=>"101111101",
  60606=>"010100000",
  60607=>"101010110",
  60608=>"111100111",
  60609=>"010100111",
  60610=>"001110101",
  60611=>"110111100",
  60612=>"101000011",
  60613=>"111001101",
  60614=>"101111110",
  60615=>"111101111",
  60616=>"011100001",
  60617=>"100000010",
  60618=>"011110001",
  60619=>"101101010",
  60620=>"100001001",
  60621=>"101101110",
  60622=>"101011001",
  60623=>"101101011",
  60624=>"000001011",
  60625=>"101101111",
  60626=>"000001111",
  60627=>"001010110",
  60628=>"011100001",
  60629=>"011111111",
  60630=>"011000101",
  60631=>"110001100",
  60632=>"010010110",
  60633=>"001010100",
  60634=>"100010000",
  60635=>"010100001",
  60636=>"010001001",
  60637=>"001111101",
  60638=>"111001111",
  60639=>"110100011",
  60640=>"001100101",
  60641=>"011111101",
  60642=>"010010011",
  60643=>"110001010",
  60644=>"000000100",
  60645=>"010110011",
  60646=>"000010100",
  60647=>"001100001",
  60648=>"011011111",
  60649=>"100001111",
  60650=>"001000001",
  60651=>"100011111",
  60652=>"010100010",
  60653=>"011101110",
  60654=>"101100111",
  60655=>"011110000",
  60656=>"110111111",
  60657=>"001101111",
  60658=>"111010011",
  60659=>"100001001",
  60660=>"100110011",
  60661=>"101110010",
  60662=>"011010010",
  60663=>"000011011",
  60664=>"111101000",
  60665=>"000010001",
  60666=>"111101001",
  60667=>"000001110",
  60668=>"010000101",
  60669=>"111101101",
  60670=>"111010010",
  60671=>"100100010",
  60672=>"111000100",
  60673=>"011100101",
  60674=>"110011100",
  60675=>"111101100",
  60676=>"100010111",
  60677=>"001101000",
  60678=>"101111110",
  60679=>"101110101",
  60680=>"001111000",
  60681=>"101001101",
  60682=>"010100010",
  60683=>"011010100",
  60684=>"110011110",
  60685=>"100010000",
  60686=>"110000001",
  60687=>"000001111",
  60688=>"100111001",
  60689=>"010111011",
  60690=>"110011101",
  60691=>"100001001",
  60692=>"001110111",
  60693=>"111011100",
  60694=>"011100000",
  60695=>"110011010",
  60696=>"001010100",
  60697=>"010100110",
  60698=>"101111001",
  60699=>"101110010",
  60700=>"111101011",
  60701=>"011101000",
  60702=>"101111110",
  60703=>"100011111",
  60704=>"011110011",
  60705=>"111001101",
  60706=>"111111011",
  60707=>"010011111",
  60708=>"010101000",
  60709=>"001110010",
  60710=>"010101000",
  60711=>"000010111",
  60712=>"010100100",
  60713=>"001011011",
  60714=>"011101100",
  60715=>"011111111",
  60716=>"110011111",
  60717=>"000000110",
  60718=>"111000000",
  60719=>"001100001",
  60720=>"111101100",
  60721=>"101011100",
  60722=>"001001001",
  60723=>"011001101",
  60724=>"110110100",
  60725=>"011100101",
  60726=>"000011011",
  60727=>"011101001",
  60728=>"011001011",
  60729=>"000111100",
  60730=>"100000001",
  60731=>"011111100",
  60732=>"000010000",
  60733=>"001111100",
  60734=>"111010101",
  60735=>"010100101",
  60736=>"010110100",
  60737=>"110100011",
  60738=>"101111111",
  60739=>"110101110",
  60740=>"011010101",
  60741=>"110010001",
  60742=>"011110000",
  60743=>"100001111",
  60744=>"101101010",
  60745=>"011000101",
  60746=>"000011100",
  60747=>"111010100",
  60748=>"110010010",
  60749=>"110110000",
  60750=>"001010010",
  60751=>"010110011",
  60752=>"000000101",
  60753=>"010000011",
  60754=>"011101000",
  60755=>"000101010",
  60756=>"010011000",
  60757=>"000011000",
  60758=>"100000100",
  60759=>"111111110",
  60760=>"101000001",
  60761=>"000111110",
  60762=>"110100011",
  60763=>"011101010",
  60764=>"001000011",
  60765=>"111100001",
  60766=>"010011100",
  60767=>"111111110",
  60768=>"000110101",
  60769=>"011110111",
  60770=>"110101101",
  60771=>"101011110",
  60772=>"111010010",
  60773=>"011000101",
  60774=>"011110010",
  60775=>"101010100",
  60776=>"001000111",
  60777=>"001101101",
  60778=>"110010110",
  60779=>"010010011",
  60780=>"110010011",
  60781=>"101001100",
  60782=>"011000011",
  60783=>"011100010",
  60784=>"011111101",
  60785=>"111111011",
  60786=>"100100100",
  60787=>"001001100",
  60788=>"100111001",
  60789=>"010000111",
  60790=>"110001000",
  60791=>"111110000",
  60792=>"001111010",
  60793=>"100100000",
  60794=>"100000101",
  60795=>"000001000",
  60796=>"010011110",
  60797=>"100111111",
  60798=>"011110101",
  60799=>"110010110",
  60800=>"111111111",
  60801=>"001010100",
  60802=>"101110110",
  60803=>"101110100",
  60804=>"101110001",
  60805=>"101001111",
  60806=>"011011001",
  60807=>"000100010",
  60808=>"000111001",
  60809=>"110001100",
  60810=>"100000111",
  60811=>"111110110",
  60812=>"000110110",
  60813=>"111001101",
  60814=>"011011111",
  60815=>"000000011",
  60816=>"011100111",
  60817=>"000000100",
  60818=>"111001001",
  60819=>"010101000",
  60820=>"110101101",
  60821=>"110000101",
  60822=>"010111000",
  60823=>"010001100",
  60824=>"110110011",
  60825=>"001111000",
  60826=>"011001111",
  60827=>"100111111",
  60828=>"011000001",
  60829=>"101011111",
  60830=>"000100100",
  60831=>"111011001",
  60832=>"010111000",
  60833=>"111001110",
  60834=>"110110001",
  60835=>"000000000",
  60836=>"110100000",
  60837=>"110110001",
  60838=>"010010011",
  60839=>"111011000",
  60840=>"110010011",
  60841=>"011011000",
  60842=>"001001011",
  60843=>"100110001",
  60844=>"001111111",
  60845=>"000011010",
  60846=>"011111001",
  60847=>"000010101",
  60848=>"011101001",
  60849=>"011011010",
  60850=>"011000001",
  60851=>"100101101",
  60852=>"000011101",
  60853=>"011111001",
  60854=>"001000011",
  60855=>"001010011",
  60856=>"111011110",
  60857=>"001100110",
  60858=>"100011010",
  60859=>"001111111",
  60860=>"110110011",
  60861=>"100100111",
  60862=>"011110111",
  60863=>"010100001",
  60864=>"010011000",
  60865=>"100011001",
  60866=>"101010001",
  60867=>"001110110",
  60868=>"111111101",
  60869=>"111000010",
  60870=>"111011111",
  60871=>"000010111",
  60872=>"110001110",
  60873=>"100111011",
  60874=>"101010101",
  60875=>"110110100",
  60876=>"101001011",
  60877=>"010011100",
  60878=>"110100011",
  60879=>"000101000",
  60880=>"110010010",
  60881=>"110011000",
  60882=>"111011001",
  60883=>"011110110",
  60884=>"000001100",
  60885=>"111101101",
  60886=>"010001010",
  60887=>"100110110",
  60888=>"101010111",
  60889=>"101001101",
  60890=>"010011101",
  60891=>"001000000",
  60892=>"111001000",
  60893=>"110010101",
  60894=>"100000001",
  60895=>"001000010",
  60896=>"111110101",
  60897=>"111110111",
  60898=>"001000010",
  60899=>"010101001",
  60900=>"111110110",
  60901=>"100000010",
  60902=>"001100111",
  60903=>"111101000",
  60904=>"111110101",
  60905=>"100011111",
  60906=>"111111101",
  60907=>"000010001",
  60908=>"110101001",
  60909=>"100010011",
  60910=>"101110100",
  60911=>"111110100",
  60912=>"101010001",
  60913=>"111001111",
  60914=>"010010101",
  60915=>"100010010",
  60916=>"101110011",
  60917=>"100100111",
  60918=>"000000010",
  60919=>"111110001",
  60920=>"000100001",
  60921=>"000001000",
  60922=>"111001011",
  60923=>"011101010",
  60924=>"000010010",
  60925=>"001000001",
  60926=>"011111011",
  60927=>"001111111",
  60928=>"100011001",
  60929=>"110001110",
  60930=>"100010101",
  60931=>"000111110",
  60932=>"000011000",
  60933=>"001011000",
  60934=>"011001011",
  60935=>"110010010",
  60936=>"000001011",
  60937=>"101111111",
  60938=>"111011010",
  60939=>"100100011",
  60940=>"011101000",
  60941=>"101111011",
  60942=>"100100011",
  60943=>"110110001",
  60944=>"110110101",
  60945=>"001111110",
  60946=>"001011100",
  60947=>"101101100",
  60948=>"011011101",
  60949=>"111001000",
  60950=>"111010001",
  60951=>"111010111",
  60952=>"111101010",
  60953=>"011111010",
  60954=>"111010001",
  60955=>"011010001",
  60956=>"001010101",
  60957=>"011111101",
  60958=>"011111000",
  60959=>"100101010",
  60960=>"000110011",
  60961=>"100001000",
  60962=>"111111110",
  60963=>"010001111",
  60964=>"110110101",
  60965=>"001111001",
  60966=>"000001111",
  60967=>"000000010",
  60968=>"010010010",
  60969=>"000101111",
  60970=>"001010011",
  60971=>"101110110",
  60972=>"000000111",
  60973=>"010010110",
  60974=>"000100111",
  60975=>"111011001",
  60976=>"110011011",
  60977=>"110101101",
  60978=>"111111010",
  60979=>"101000110",
  60980=>"100010000",
  60981=>"011010001",
  60982=>"101000101",
  60983=>"000011100",
  60984=>"111011110",
  60985=>"111000010",
  60986=>"111000101",
  60987=>"111110010",
  60988=>"101001110",
  60989=>"111001001",
  60990=>"000011010",
  60991=>"000111010",
  60992=>"001101111",
  60993=>"010111110",
  60994=>"100010101",
  60995=>"111100111",
  60996=>"000000101",
  60997=>"001111100",
  60998=>"101111111",
  60999=>"100111000",
  61000=>"011101111",
  61001=>"110000100",
  61002=>"111000000",
  61003=>"000001000",
  61004=>"111110111",
  61005=>"011001011",
  61006=>"101100110",
  61007=>"111101100",
  61008=>"111000000",
  61009=>"110100110",
  61010=>"111010101",
  61011=>"010011100",
  61012=>"111110101",
  61013=>"101000100",
  61014=>"010010011",
  61015=>"010011101",
  61016=>"011111011",
  61017=>"100111011",
  61018=>"001000000",
  61019=>"000101000",
  61020=>"001001000",
  61021=>"000000111",
  61022=>"110110101",
  61023=>"011010000",
  61024=>"101011010",
  61025=>"111001011",
  61026=>"100111101",
  61027=>"101000111",
  61028=>"001110001",
  61029=>"010101111",
  61030=>"001011100",
  61031=>"011011101",
  61032=>"011010001",
  61033=>"100111110",
  61034=>"010101001",
  61035=>"000001110",
  61036=>"010010010",
  61037=>"001011101",
  61038=>"011010001",
  61039=>"110110011",
  61040=>"111110110",
  61041=>"101100000",
  61042=>"100001011",
  61043=>"001010111",
  61044=>"010010101",
  61045=>"111100110",
  61046=>"110110000",
  61047=>"101101110",
  61048=>"010111000",
  61049=>"111100100",
  61050=>"110011101",
  61051=>"110100011",
  61052=>"100101111",
  61053=>"101100001",
  61054=>"101001111",
  61055=>"011111010",
  61056=>"100111110",
  61057=>"011100110",
  61058=>"011011011",
  61059=>"011001100",
  61060=>"100101101",
  61061=>"101110111",
  61062=>"100001011",
  61063=>"010100101",
  61064=>"011001111",
  61065=>"000111010",
  61066=>"011110100",
  61067=>"000111110",
  61068=>"011010000",
  61069=>"010010110",
  61070=>"010000101",
  61071=>"111100110",
  61072=>"011011010",
  61073=>"110111000",
  61074=>"111001100",
  61075=>"010010100",
  61076=>"110001001",
  61077=>"001011010",
  61078=>"111110010",
  61079=>"010101100",
  61080=>"110010001",
  61081=>"001100010",
  61082=>"100011100",
  61083=>"101110000",
  61084=>"000111111",
  61085=>"111100111",
  61086=>"111001101",
  61087=>"101100001",
  61088=>"010001000",
  61089=>"011111111",
  61090=>"110001101",
  61091=>"100111101",
  61092=>"101101100",
  61093=>"010010011",
  61094=>"011110110",
  61095=>"000010010",
  61096=>"111101110",
  61097=>"111001010",
  61098=>"001011001",
  61099=>"111001111",
  61100=>"000000000",
  61101=>"110011101",
  61102=>"111100111",
  61103=>"011001010",
  61104=>"111010100",
  61105=>"010110111",
  61106=>"110000000",
  61107=>"111011101",
  61108=>"111111000",
  61109=>"011111001",
  61110=>"010001000",
  61111=>"010110101",
  61112=>"000110100",
  61113=>"001000010",
  61114=>"011111111",
  61115=>"001110001",
  61116=>"101010110",
  61117=>"101011001",
  61118=>"101000101",
  61119=>"100000001",
  61120=>"001110101",
  61121=>"100000010",
  61122=>"001111000",
  61123=>"100010000",
  61124=>"101111101",
  61125=>"001101001",
  61126=>"011000101",
  61127=>"010101110",
  61128=>"111000010",
  61129=>"001100010",
  61130=>"001010101",
  61131=>"101111101",
  61132=>"010010111",
  61133=>"000101111",
  61134=>"010100110",
  61135=>"010000000",
  61136=>"101000101",
  61137=>"010011001",
  61138=>"011000100",
  61139=>"100010001",
  61140=>"001111101",
  61141=>"101000111",
  61142=>"011010011",
  61143=>"110101111",
  61144=>"010111010",
  61145=>"011111000",
  61146=>"011001101",
  61147=>"010110010",
  61148=>"101101111",
  61149=>"001110011",
  61150=>"001100010",
  61151=>"101110111",
  61152=>"111101110",
  61153=>"100000001",
  61154=>"101100111",
  61155=>"000010110",
  61156=>"111100111",
  61157=>"000011011",
  61158=>"001100110",
  61159=>"110101101",
  61160=>"111101000",
  61161=>"001010110",
  61162=>"000010011",
  61163=>"101111010",
  61164=>"101110111",
  61165=>"101001111",
  61166=>"010001010",
  61167=>"100110011",
  61168=>"110101100",
  61169=>"101100101",
  61170=>"111011000",
  61171=>"110100010",
  61172=>"111110001",
  61173=>"100010010",
  61174=>"100010001",
  61175=>"111001000",
  61176=>"010011000",
  61177=>"001001101",
  61178=>"110100011",
  61179=>"100001000",
  61180=>"111011011",
  61181=>"100101011",
  61182=>"010111111",
  61183=>"101000101",
  61184=>"101001011",
  61185=>"101100010",
  61186=>"010100011",
  61187=>"101010000",
  61188=>"111101101",
  61189=>"001010001",
  61190=>"110101110",
  61191=>"110011110",
  61192=>"000101101",
  61193=>"110101000",
  61194=>"101111000",
  61195=>"001000100",
  61196=>"011110101",
  61197=>"101001111",
  61198=>"100010111",
  61199=>"011011010",
  61200=>"011000010",
  61201=>"010000001",
  61202=>"101001111",
  61203=>"110100001",
  61204=>"100100100",
  61205=>"011011110",
  61206=>"101111011",
  61207=>"001010011",
  61208=>"000110101",
  61209=>"001010000",
  61210=>"111010011",
  61211=>"101010111",
  61212=>"010010000",
  61213=>"101000000",
  61214=>"010011101",
  61215=>"100101111",
  61216=>"100001101",
  61217=>"000110111",
  61218=>"011010000",
  61219=>"011010010",
  61220=>"010110011",
  61221=>"000100111",
  61222=>"101011000",
  61223=>"010001101",
  61224=>"000111010",
  61225=>"001100100",
  61226=>"001111001",
  61227=>"110001100",
  61228=>"101110101",
  61229=>"111001110",
  61230=>"110110100",
  61231=>"010100011",
  61232=>"000000110",
  61233=>"110100011",
  61234=>"011101011",
  61235=>"001100100",
  61236=>"110001001",
  61237=>"011010010",
  61238=>"110100010",
  61239=>"111011001",
  61240=>"111111101",
  61241=>"100001000",
  61242=>"011001001",
  61243=>"001000000",
  61244=>"110011011",
  61245=>"100001010",
  61246=>"100010110",
  61247=>"011000000",
  61248=>"001000000",
  61249=>"100100011",
  61250=>"111110010",
  61251=>"101011111",
  61252=>"010110110",
  61253=>"000001001",
  61254=>"101001000",
  61255=>"101101110",
  61256=>"011011111",
  61257=>"111000110",
  61258=>"110000010",
  61259=>"110010100",
  61260=>"110001010",
  61261=>"011111111",
  61262=>"110000001",
  61263=>"100100010",
  61264=>"100101111",
  61265=>"101101000",
  61266=>"110111110",
  61267=>"110100001",
  61268=>"110011101",
  61269=>"001111001",
  61270=>"010001000",
  61271=>"000101110",
  61272=>"011111101",
  61273=>"100000110",
  61274=>"001100101",
  61275=>"010101011",
  61276=>"010011000",
  61277=>"010100011",
  61278=>"111111111",
  61279=>"011101101",
  61280=>"000110110",
  61281=>"001100110",
  61282=>"101111101",
  61283=>"011000110",
  61284=>"110110110",
  61285=>"001010000",
  61286=>"011100110",
  61287=>"000101111",
  61288=>"000000011",
  61289=>"101100011",
  61290=>"010001111",
  61291=>"000010001",
  61292=>"010000000",
  61293=>"000000000",
  61294=>"011101000",
  61295=>"010111000",
  61296=>"111101001",
  61297=>"011010011",
  61298=>"110100111",
  61299=>"101010110",
  61300=>"111000110",
  61301=>"001011011",
  61302=>"111111110",
  61303=>"111001000",
  61304=>"101110110",
  61305=>"001011110",
  61306=>"101111101",
  61307=>"100111100",
  61308=>"110011101",
  61309=>"010000000",
  61310=>"100111010",
  61311=>"111111110",
  61312=>"001110101",
  61313=>"101111001",
  61314=>"100101111",
  61315=>"000111101",
  61316=>"011110001",
  61317=>"001101010",
  61318=>"111001110",
  61319=>"010110001",
  61320=>"110011111",
  61321=>"110100011",
  61322=>"011101011",
  61323=>"001110010",
  61324=>"100000111",
  61325=>"001110000",
  61326=>"001111111",
  61327=>"111001000",
  61328=>"000010010",
  61329=>"110001110",
  61330=>"101001111",
  61331=>"100111000",
  61332=>"001001101",
  61333=>"101100110",
  61334=>"010111000",
  61335=>"101010101",
  61336=>"100010011",
  61337=>"000010111",
  61338=>"110000110",
  61339=>"011101110",
  61340=>"010001100",
  61341=>"111101100",
  61342=>"001000101",
  61343=>"110000000",
  61344=>"111010100",
  61345=>"111010101",
  61346=>"101111011",
  61347=>"011011110",
  61348=>"000001001",
  61349=>"001111111",
  61350=>"010010111",
  61351=>"000100111",
  61352=>"111100101",
  61353=>"001110110",
  61354=>"101100011",
  61355=>"010100110",
  61356=>"101101000",
  61357=>"101100110",
  61358=>"110001111",
  61359=>"101000000",
  61360=>"000101010",
  61361=>"100000010",
  61362=>"100100111",
  61363=>"101100010",
  61364=>"010011110",
  61365=>"111110101",
  61366=>"010011111",
  61367=>"100110111",
  61368=>"101100100",
  61369=>"000100010",
  61370=>"100000111",
  61371=>"111010000",
  61372=>"101101010",
  61373=>"111110100",
  61374=>"100100010",
  61375=>"011000000",
  61376=>"001011011",
  61377=>"111100101",
  61378=>"111101100",
  61379=>"010101111",
  61380=>"000011000",
  61381=>"010011101",
  61382=>"111111101",
  61383=>"110000011",
  61384=>"011011111",
  61385=>"010011100",
  61386=>"010100100",
  61387=>"111110110",
  61388=>"101010010",
  61389=>"111110001",
  61390=>"001111010",
  61391=>"000011000",
  61392=>"110101100",
  61393=>"000100110",
  61394=>"000101011",
  61395=>"111000111",
  61396=>"011111000",
  61397=>"110100111",
  61398=>"010111110",
  61399=>"111111110",
  61400=>"010100110",
  61401=>"001111100",
  61402=>"100101110",
  61403=>"001000111",
  61404=>"011110010",
  61405=>"101001000",
  61406=>"101100110",
  61407=>"100110001",
  61408=>"111110011",
  61409=>"000000011",
  61410=>"001011110",
  61411=>"101110110",
  61412=>"010000011",
  61413=>"110110000",
  61414=>"101000010",
  61415=>"001001101",
  61416=>"010001000",
  61417=>"100100100",
  61418=>"000001011",
  61419=>"000000111",
  61420=>"001001000",
  61421=>"001101111",
  61422=>"100000100",
  61423=>"110001011",
  61424=>"011001100",
  61425=>"001010100",
  61426=>"111011110",
  61427=>"011111001",
  61428=>"010000001",
  61429=>"001110001",
  61430=>"010110010",
  61431=>"110100101",
  61432=>"111110100",
  61433=>"110100010",
  61434=>"101111111",
  61435=>"110011000",
  61436=>"010010111",
  61437=>"111001111",
  61438=>"110011010",
  61439=>"100100010",
  61440=>"100100100",
  61441=>"000110001",
  61442=>"111011110",
  61443=>"110011111",
  61444=>"110001101",
  61445=>"011101000",
  61446=>"101101100",
  61447=>"000000100",
  61448=>"010111110",
  61449=>"101001001",
  61450=>"111000111",
  61451=>"101011101",
  61452=>"101101000",
  61453=>"001000001",
  61454=>"110101100",
  61455=>"001011110",
  61456=>"110010010",
  61457=>"111100011",
  61458=>"101110001",
  61459=>"010010100",
  61460=>"011101010",
  61461=>"101000010",
  61462=>"000010000",
  61463=>"100101111",
  61464=>"001000000",
  61465=>"110101001",
  61466=>"011000000",
  61467=>"000000011",
  61468=>"000010010",
  61469=>"011111100",
  61470=>"110111001",
  61471=>"101101111",
  61472=>"011010000",
  61473=>"111011101",
  61474=>"011011100",
  61475=>"000001010",
  61476=>"110111000",
  61477=>"111010011",
  61478=>"000110001",
  61479=>"110100100",
  61480=>"100001101",
  61481=>"111110101",
  61482=>"000101110",
  61483=>"010001000",
  61484=>"000111011",
  61485=>"011010010",
  61486=>"010011100",
  61487=>"111011011",
  61488=>"000110100",
  61489=>"101111100",
  61490=>"010111010",
  61491=>"000111000",
  61492=>"000101110",
  61493=>"111110101",
  61494=>"010001010",
  61495=>"100111101",
  61496=>"001001010",
  61497=>"101011001",
  61498=>"101101010",
  61499=>"110111010",
  61500=>"001010000",
  61501=>"100101101",
  61502=>"001011000",
  61503=>"010010000",
  61504=>"000001100",
  61505=>"010010110",
  61506=>"101001000",
  61507=>"001010101",
  61508=>"100100110",
  61509=>"101101100",
  61510=>"001011001",
  61511=>"111111100",
  61512=>"010011110",
  61513=>"100001111",
  61514=>"100000010",
  61515=>"100100100",
  61516=>"101100001",
  61517=>"001110000",
  61518=>"100111011",
  61519=>"001001000",
  61520=>"110010100",
  61521=>"000101101",
  61522=>"000111100",
  61523=>"000011101",
  61524=>"011011110",
  61525=>"001101011",
  61526=>"101010100",
  61527=>"000000111",
  61528=>"111111001",
  61529=>"000100100",
  61530=>"010100100",
  61531=>"101111100",
  61532=>"011110010",
  61533=>"011010100",
  61534=>"110000001",
  61535=>"000011101",
  61536=>"010111001",
  61537=>"001111101",
  61538=>"011010111",
  61539=>"001001011",
  61540=>"000010010",
  61541=>"010111110",
  61542=>"000111010",
  61543=>"000000101",
  61544=>"111011110",
  61545=>"000111010",
  61546=>"110100001",
  61547=>"010011101",
  61548=>"010101001",
  61549=>"100011011",
  61550=>"010100110",
  61551=>"000011110",
  61552=>"100010000",
  61553=>"101111100",
  61554=>"001000000",
  61555=>"010110110",
  61556=>"110011001",
  61557=>"000001001",
  61558=>"111111110",
  61559=>"101110001",
  61560=>"100001001",
  61561=>"100001011",
  61562=>"110100000",
  61563=>"100101111",
  61564=>"110111101",
  61565=>"101100111",
  61566=>"100100010",
  61567=>"001001000",
  61568=>"001001111",
  61569=>"001110110",
  61570=>"011110010",
  61571=>"001100000",
  61572=>"101001001",
  61573=>"000000010",
  61574=>"000110101",
  61575=>"100101100",
  61576=>"101011000",
  61577=>"100011000",
  61578=>"011010111",
  61579=>"100001111",
  61580=>"111100011",
  61581=>"110000011",
  61582=>"011001101",
  61583=>"000101101",
  61584=>"100111000",
  61585=>"001000001",
  61586=>"011010010",
  61587=>"001111101",
  61588=>"101111010",
  61589=>"100101111",
  61590=>"011101010",
  61591=>"100111100",
  61592=>"010100101",
  61593=>"110000110",
  61594=>"001010100",
  61595=>"101010010",
  61596=>"100000000",
  61597=>"000000000",
  61598=>"101010100",
  61599=>"101000010",
  61600=>"101100001",
  61601=>"010110100",
  61602=>"110011011",
  61603=>"001111110",
  61604=>"111101101",
  61605=>"010100110",
  61606=>"110001000",
  61607=>"111111011",
  61608=>"110011111",
  61609=>"011100111",
  61610=>"011111000",
  61611=>"001000000",
  61612=>"001010100",
  61613=>"001011011",
  61614=>"111011011",
  61615=>"010111010",
  61616=>"010100101",
  61617=>"111101001",
  61618=>"001010001",
  61619=>"111111110",
  61620=>"111100101",
  61621=>"001110111",
  61622=>"110111101",
  61623=>"101010010",
  61624=>"011010111",
  61625=>"000110000",
  61626=>"110100010",
  61627=>"010111001",
  61628=>"000000101",
  61629=>"000101110",
  61630=>"000011111",
  61631=>"010110111",
  61632=>"011111001",
  61633=>"101011001",
  61634=>"010011010",
  61635=>"011110010",
  61636=>"011010010",
  61637=>"010001101",
  61638=>"000101111",
  61639=>"000110011",
  61640=>"101101111",
  61641=>"111001101",
  61642=>"100000111",
  61643=>"101000010",
  61644=>"110001010",
  61645=>"110000101",
  61646=>"101111111",
  61647=>"111000011",
  61648=>"001111111",
  61649=>"001111111",
  61650=>"000011000",
  61651=>"110100000",
  61652=>"101001001",
  61653=>"011110000",
  61654=>"100010100",
  61655=>"100001101",
  61656=>"001000000",
  61657=>"100010110",
  61658=>"000001001",
  61659=>"000000001",
  61660=>"100101000",
  61661=>"010100111",
  61662=>"000110001",
  61663=>"000111111",
  61664=>"100111000",
  61665=>"110000100",
  61666=>"111111111",
  61667=>"011011001",
  61668=>"001011001",
  61669=>"111111011",
  61670=>"100101000",
  61671=>"010111111",
  61672=>"101110000",
  61673=>"011111000",
  61674=>"011001110",
  61675=>"100001110",
  61676=>"011000010",
  61677=>"011010000",
  61678=>"010010011",
  61679=>"010010000",
  61680=>"000000010",
  61681=>"000100011",
  61682=>"001100011",
  61683=>"000110011",
  61684=>"000010110",
  61685=>"001000100",
  61686=>"101110100",
  61687=>"111010000",
  61688=>"001100101",
  61689=>"111111100",
  61690=>"111110100",
  61691=>"011111000",
  61692=>"101011100",
  61693=>"101110110",
  61694=>"000010000",
  61695=>"010011100",
  61696=>"100110011",
  61697=>"001111010",
  61698=>"011111001",
  61699=>"001110100",
  61700=>"111100001",
  61701=>"001101011",
  61702=>"001100011",
  61703=>"110100101",
  61704=>"111111110",
  61705=>"010010000",
  61706=>"000011100",
  61707=>"101010010",
  61708=>"111000000",
  61709=>"100010010",
  61710=>"001101001",
  61711=>"111010110",
  61712=>"000001000",
  61713=>"010101011",
  61714=>"000010100",
  61715=>"111000110",
  61716=>"011101001",
  61717=>"110100010",
  61718=>"101100101",
  61719=>"110001000",
  61720=>"111001001",
  61721=>"100101011",
  61722=>"000100110",
  61723=>"110100010",
  61724=>"100110010",
  61725=>"101110100",
  61726=>"100010111",
  61727=>"100001111",
  61728=>"110000001",
  61729=>"000100010",
  61730=>"000000010",
  61731=>"011100110",
  61732=>"011011010",
  61733=>"010100000",
  61734=>"110011111",
  61735=>"001011111",
  61736=>"100000100",
  61737=>"100000110",
  61738=>"010001001",
  61739=>"001101000",
  61740=>"100111001",
  61741=>"110110000",
  61742=>"011111011",
  61743=>"010010100",
  61744=>"110111101",
  61745=>"000001001",
  61746=>"111110111",
  61747=>"110100010",
  61748=>"011010000",
  61749=>"001011000",
  61750=>"010001000",
  61751=>"011001000",
  61752=>"000000000",
  61753=>"100101100",
  61754=>"101100100",
  61755=>"101111101",
  61756=>"110110110",
  61757=>"100101000",
  61758=>"110101010",
  61759=>"010101110",
  61760=>"110011100",
  61761=>"010111000",
  61762=>"101011001",
  61763=>"011010111",
  61764=>"110100111",
  61765=>"110111110",
  61766=>"000101011",
  61767=>"111110100",
  61768=>"000100001",
  61769=>"111101010",
  61770=>"001111000",
  61771=>"000000001",
  61772=>"011001101",
  61773=>"000111100",
  61774=>"101100111",
  61775=>"000011010",
  61776=>"111100011",
  61777=>"101010001",
  61778=>"000000010",
  61779=>"001110011",
  61780=>"100001000",
  61781=>"101001100",
  61782=>"110110010",
  61783=>"011011101",
  61784=>"110100110",
  61785=>"000110001",
  61786=>"000110100",
  61787=>"010001101",
  61788=>"110000001",
  61789=>"100000100",
  61790=>"000110110",
  61791=>"110110011",
  61792=>"001011000",
  61793=>"000111000",
  61794=>"110110101",
  61795=>"011100110",
  61796=>"000011111",
  61797=>"110101111",
  61798=>"010011011",
  61799=>"000001011",
  61800=>"010100111",
  61801=>"010101101",
  61802=>"101110101",
  61803=>"001010111",
  61804=>"101011101",
  61805=>"000011000",
  61806=>"110001010",
  61807=>"101001010",
  61808=>"111011101",
  61809=>"000010110",
  61810=>"011110001",
  61811=>"101110110",
  61812=>"100110000",
  61813=>"111101101",
  61814=>"011101101",
  61815=>"110101001",
  61816=>"001101100",
  61817=>"001000111",
  61818=>"101101011",
  61819=>"100110001",
  61820=>"000010110",
  61821=>"010111101",
  61822=>"001001111",
  61823=>"100101000",
  61824=>"110111010",
  61825=>"111000100",
  61826=>"101111110",
  61827=>"101101101",
  61828=>"100010110",
  61829=>"001101011",
  61830=>"011001010",
  61831=>"110000101",
  61832=>"111010100",
  61833=>"110110000",
  61834=>"111101001",
  61835=>"001000100",
  61836=>"101101110",
  61837=>"010011110",
  61838=>"010010010",
  61839=>"111000110",
  61840=>"111001000",
  61841=>"011100100",
  61842=>"011110111",
  61843=>"101000100",
  61844=>"111101011",
  61845=>"011011010",
  61846=>"110111011",
  61847=>"000011100",
  61848=>"100101101",
  61849=>"010111110",
  61850=>"100001001",
  61851=>"001101111",
  61852=>"100010111",
  61853=>"111011010",
  61854=>"101000000",
  61855=>"110101101",
  61856=>"110001000",
  61857=>"111101100",
  61858=>"111010001",
  61859=>"011111100",
  61860=>"101001000",
  61861=>"111000100",
  61862=>"010010001",
  61863=>"110001110",
  61864=>"110110001",
  61865=>"000001011",
  61866=>"110011110",
  61867=>"111101000",
  61868=>"011011010",
  61869=>"001011011",
  61870=>"010000100",
  61871=>"101110111",
  61872=>"111101000",
  61873=>"000110011",
  61874=>"011101001",
  61875=>"010010000",
  61876=>"011000111",
  61877=>"100000000",
  61878=>"000111011",
  61879=>"011111001",
  61880=>"000100001",
  61881=>"010110110",
  61882=>"111011000",
  61883=>"111011101",
  61884=>"110101111",
  61885=>"010001001",
  61886=>"110001110",
  61887=>"111000111",
  61888=>"000011011",
  61889=>"000110111",
  61890=>"010000010",
  61891=>"100111111",
  61892=>"000101010",
  61893=>"110010101",
  61894=>"010001111",
  61895=>"111011110",
  61896=>"110001111",
  61897=>"110011100",
  61898=>"011100001",
  61899=>"110111100",
  61900=>"110011111",
  61901=>"011010011",
  61902=>"000010110",
  61903=>"101110101",
  61904=>"111010110",
  61905=>"010001111",
  61906=>"100011111",
  61907=>"011100101",
  61908=>"000001110",
  61909=>"001100100",
  61910=>"001000001",
  61911=>"011011001",
  61912=>"010110100",
  61913=>"101011101",
  61914=>"001011011",
  61915=>"010010110",
  61916=>"001101101",
  61917=>"001000011",
  61918=>"101100010",
  61919=>"110001110",
  61920=>"100110110",
  61921=>"111010100",
  61922=>"010111111",
  61923=>"001100111",
  61924=>"000000000",
  61925=>"001110011",
  61926=>"111101100",
  61927=>"010000100",
  61928=>"111100011",
  61929=>"010011110",
  61930=>"110100100",
  61931=>"001110011",
  61932=>"100010000",
  61933=>"011000100",
  61934=>"101011001",
  61935=>"101010001",
  61936=>"100111101",
  61937=>"010010000",
  61938=>"000100110",
  61939=>"101110011",
  61940=>"010010001",
  61941=>"000110011",
  61942=>"110000110",
  61943=>"001110110",
  61944=>"010010010",
  61945=>"011111000",
  61946=>"110010110",
  61947=>"110110011",
  61948=>"101111100",
  61949=>"000100100",
  61950=>"001101111",
  61951=>"101001000",
  61952=>"100101010",
  61953=>"011001011",
  61954=>"001000111",
  61955=>"000010010",
  61956=>"101000100",
  61957=>"101100000",
  61958=>"010011001",
  61959=>"101001100",
  61960=>"000010000",
  61961=>"110000101",
  61962=>"001010100",
  61963=>"111111000",
  61964=>"111100100",
  61965=>"111101111",
  61966=>"101001111",
  61967=>"100111001",
  61968=>"110110100",
  61969=>"110011011",
  61970=>"000110110",
  61971=>"100110011",
  61972=>"100011011",
  61973=>"010111111",
  61974=>"110100010",
  61975=>"001111010",
  61976=>"111011001",
  61977=>"010010111",
  61978=>"010011111",
  61979=>"110110101",
  61980=>"111010111",
  61981=>"110011001",
  61982=>"111111110",
  61983=>"000010101",
  61984=>"101000000",
  61985=>"010110001",
  61986=>"111111000",
  61987=>"001011111",
  61988=>"100101011",
  61989=>"011101000",
  61990=>"001100110",
  61991=>"101100100",
  61992=>"100000101",
  61993=>"101001110",
  61994=>"010000001",
  61995=>"110111010",
  61996=>"011110110",
  61997=>"110001010",
  61998=>"010000101",
  61999=>"001100001",
  62000=>"000110100",
  62001=>"101011101",
  62002=>"101000111",
  62003=>"101001101",
  62004=>"101010000",
  62005=>"011011000",
  62006=>"011111001",
  62007=>"111111001",
  62008=>"011011101",
  62009=>"011111000",
  62010=>"000100111",
  62011=>"010100110",
  62012=>"101011011",
  62013=>"111000010",
  62014=>"100000000",
  62015=>"000011000",
  62016=>"100111100",
  62017=>"001000011",
  62018=>"110010000",
  62019=>"111011001",
  62020=>"001000001",
  62021=>"111111110",
  62022=>"000010000",
  62023=>"100111001",
  62024=>"101110000",
  62025=>"000110000",
  62026=>"100101111",
  62027=>"101001011",
  62028=>"101110000",
  62029=>"000110100",
  62030=>"101110001",
  62031=>"010100100",
  62032=>"010011001",
  62033=>"010110100",
  62034=>"100010111",
  62035=>"001100110",
  62036=>"110000011",
  62037=>"110100010",
  62038=>"111000010",
  62039=>"111111111",
  62040=>"101010010",
  62041=>"000011101",
  62042=>"100010011",
  62043=>"111101011",
  62044=>"011111111",
  62045=>"001001010",
  62046=>"000001110",
  62047=>"001110001",
  62048=>"000010111",
  62049=>"111101000",
  62050=>"111101101",
  62051=>"000011111",
  62052=>"001000110",
  62053=>"001011111",
  62054=>"111100100",
  62055=>"111000001",
  62056=>"011001011",
  62057=>"111100110",
  62058=>"010000011",
  62059=>"111001110",
  62060=>"011100010",
  62061=>"010111100",
  62062=>"001001000",
  62063=>"001001000",
  62064=>"100010000",
  62065=>"000010000",
  62066=>"000001010",
  62067=>"101110100",
  62068=>"111111101",
  62069=>"001100000",
  62070=>"010001001",
  62071=>"101110110",
  62072=>"010000011",
  62073=>"000000011",
  62074=>"000110110",
  62075=>"000101101",
  62076=>"001111010",
  62077=>"000011000",
  62078=>"110100101",
  62079=>"111100010",
  62080=>"001111111",
  62081=>"110101110",
  62082=>"010101001",
  62083=>"101100011",
  62084=>"010100001",
  62085=>"100001000",
  62086=>"011001000",
  62087=>"000010111",
  62088=>"011110110",
  62089=>"110100100",
  62090=>"000010111",
  62091=>"111010000",
  62092=>"001011000",
  62093=>"010000110",
  62094=>"110111000",
  62095=>"101111000",
  62096=>"001011101",
  62097=>"001000011",
  62098=>"111000111",
  62099=>"000011100",
  62100=>"111011001",
  62101=>"010010111",
  62102=>"001010011",
  62103=>"010001111",
  62104=>"110011100",
  62105=>"110000001",
  62106=>"000000011",
  62107=>"010100010",
  62108=>"000000000",
  62109=>"111011101",
  62110=>"111111011",
  62111=>"010000100",
  62112=>"001110110",
  62113=>"010011100",
  62114=>"100111100",
  62115=>"110001110",
  62116=>"110101001",
  62117=>"110111001",
  62118=>"001011001",
  62119=>"111000000",
  62120=>"001011011",
  62121=>"101101001",
  62122=>"110111000",
  62123=>"000100000",
  62124=>"000000010",
  62125=>"011101100",
  62126=>"011111001",
  62127=>"110010011",
  62128=>"111000100",
  62129=>"011100110",
  62130=>"101100110",
  62131=>"010101101",
  62132=>"110011100",
  62133=>"100001110",
  62134=>"111111110",
  62135=>"101110111",
  62136=>"100100111",
  62137=>"111010010",
  62138=>"110110100",
  62139=>"100111110",
  62140=>"000011101",
  62141=>"001010010",
  62142=>"100011000",
  62143=>"111100101",
  62144=>"011110100",
  62145=>"110111010",
  62146=>"100000100",
  62147=>"111101000",
  62148=>"001001100",
  62149=>"111110101",
  62150=>"011111001",
  62151=>"111001100",
  62152=>"011101111",
  62153=>"111111010",
  62154=>"110100101",
  62155=>"001110000",
  62156=>"010110001",
  62157=>"100001001",
  62158=>"110010101",
  62159=>"010111101",
  62160=>"111101110",
  62161=>"100110000",
  62162=>"010011000",
  62163=>"001110011",
  62164=>"011101000",
  62165=>"001110110",
  62166=>"100010010",
  62167=>"100111101",
  62168=>"111101011",
  62169=>"010011100",
  62170=>"110101110",
  62171=>"010000000",
  62172=>"000011100",
  62173=>"000111110",
  62174=>"001010101",
  62175=>"010011000",
  62176=>"001001100",
  62177=>"101110111",
  62178=>"110011101",
  62179=>"111010000",
  62180=>"111011111",
  62181=>"111110100",
  62182=>"101011000",
  62183=>"001000001",
  62184=>"100110111",
  62185=>"000101001",
  62186=>"001101110",
  62187=>"010110010",
  62188=>"011010000",
  62189=>"110001010",
  62190=>"001001001",
  62191=>"000101011",
  62192=>"111011101",
  62193=>"000101010",
  62194=>"110001100",
  62195=>"110000110",
  62196=>"111011100",
  62197=>"011011100",
  62198=>"000010110",
  62199=>"000010101",
  62200=>"110111110",
  62201=>"100110000",
  62202=>"111100000",
  62203=>"000011011",
  62204=>"110001000",
  62205=>"101111101",
  62206=>"100001000",
  62207=>"001100010",
  62208=>"000101101",
  62209=>"010011011",
  62210=>"000101110",
  62211=>"000100001",
  62212=>"001111010",
  62213=>"100110110",
  62214=>"110010011",
  62215=>"110010011",
  62216=>"100010000",
  62217=>"001101101",
  62218=>"001101000",
  62219=>"011110010",
  62220=>"101010100",
  62221=>"100101101",
  62222=>"000000000",
  62223=>"100000111",
  62224=>"110100011",
  62225=>"010000101",
  62226=>"110011010",
  62227=>"001000100",
  62228=>"010110110",
  62229=>"001001010",
  62230=>"010101100",
  62231=>"001100111",
  62232=>"001110011",
  62233=>"101010000",
  62234=>"001011011",
  62235=>"011010000",
  62236=>"100100101",
  62237=>"000000111",
  62238=>"111101001",
  62239=>"110101101",
  62240=>"001000011",
  62241=>"101101001",
  62242=>"110111101",
  62243=>"000001001",
  62244=>"000011110",
  62245=>"001001010",
  62246=>"000110001",
  62247=>"000001110",
  62248=>"101110100",
  62249=>"010111011",
  62250=>"111100111",
  62251=>"010111101",
  62252=>"101011100",
  62253=>"010001110",
  62254=>"100001100",
  62255=>"110111100",
  62256=>"011000100",
  62257=>"000100111",
  62258=>"110100010",
  62259=>"011011101",
  62260=>"111001000",
  62261=>"001010111",
  62262=>"101001010",
  62263=>"111110011",
  62264=>"011001010",
  62265=>"100010100",
  62266=>"101000111",
  62267=>"100011100",
  62268=>"101110000",
  62269=>"101100101",
  62270=>"110001110",
  62271=>"110101100",
  62272=>"101110000",
  62273=>"011110001",
  62274=>"111000101",
  62275=>"011010100",
  62276=>"011010111",
  62277=>"011110111",
  62278=>"010110101",
  62279=>"101000110",
  62280=>"001101000",
  62281=>"000001101",
  62282=>"110010011",
  62283=>"110111100",
  62284=>"000001110",
  62285=>"000000100",
  62286=>"111101100",
  62287=>"011100011",
  62288=>"100100010",
  62289=>"001111101",
  62290=>"111001100",
  62291=>"001000000",
  62292=>"000001010",
  62293=>"110100101",
  62294=>"001000000",
  62295=>"000001110",
  62296=>"000101110",
  62297=>"010001010",
  62298=>"000111010",
  62299=>"101100011",
  62300=>"110110000",
  62301=>"100000100",
  62302=>"001100011",
  62303=>"110011111",
  62304=>"110110001",
  62305=>"011001010",
  62306=>"111111001",
  62307=>"001010000",
  62308=>"010011100",
  62309=>"111111110",
  62310=>"110100101",
  62311=>"000011111",
  62312=>"110111111",
  62313=>"111111101",
  62314=>"011100011",
  62315=>"011001001",
  62316=>"110101000",
  62317=>"110010111",
  62318=>"000001101",
  62319=>"000101111",
  62320=>"100111011",
  62321=>"011111010",
  62322=>"111100101",
  62323=>"010000100",
  62324=>"111111111",
  62325=>"111110111",
  62326=>"010100100",
  62327=>"000010101",
  62328=>"011101111",
  62329=>"111011111",
  62330=>"010011101",
  62331=>"110101000",
  62332=>"111000101",
  62333=>"001110110",
  62334=>"110000001",
  62335=>"000011101",
  62336=>"010110001",
  62337=>"111110111",
  62338=>"001110101",
  62339=>"101001010",
  62340=>"000010000",
  62341=>"000001000",
  62342=>"001111001",
  62343=>"000111001",
  62344=>"011000101",
  62345=>"001110101",
  62346=>"111011111",
  62347=>"001001110",
  62348=>"001110100",
  62349=>"110100011",
  62350=>"101001101",
  62351=>"000101101",
  62352=>"111001100",
  62353=>"001110110",
  62354=>"110000000",
  62355=>"110000000",
  62356=>"111111111",
  62357=>"110011001",
  62358=>"111101111",
  62359=>"010010100",
  62360=>"010110011",
  62361=>"101111100",
  62362=>"011011111",
  62363=>"001011111",
  62364=>"110110000",
  62365=>"010000011",
  62366=>"100001011",
  62367=>"001100110",
  62368=>"000100010",
  62369=>"111000011",
  62370=>"010011111",
  62371=>"001001001",
  62372=>"000111011",
  62373=>"010100001",
  62374=>"011011110",
  62375=>"100001100",
  62376=>"001111001",
  62377=>"011011010",
  62378=>"010101011",
  62379=>"100000101",
  62380=>"000100101",
  62381=>"111101011",
  62382=>"101111110",
  62383=>"100110001",
  62384=>"001011001",
  62385=>"101101010",
  62386=>"000101010",
  62387=>"001001100",
  62388=>"111001101",
  62389=>"000011100",
  62390=>"111000000",
  62391=>"011010110",
  62392=>"001010110",
  62393=>"111110110",
  62394=>"100000101",
  62395=>"001111010",
  62396=>"000000011",
  62397=>"000100001",
  62398=>"111010111",
  62399=>"111000111",
  62400=>"010001111",
  62401=>"011101111",
  62402=>"111000111",
  62403=>"010100001",
  62404=>"001101101",
  62405=>"111100000",
  62406=>"100010101",
  62407=>"000100001",
  62408=>"111100111",
  62409=>"101000011",
  62410=>"000111110",
  62411=>"001110010",
  62412=>"000110101",
  62413=>"100010111",
  62414=>"011001101",
  62415=>"000001101",
  62416=>"011010111",
  62417=>"101101011",
  62418=>"111011100",
  62419=>"001000101",
  62420=>"110110011",
  62421=>"011000000",
  62422=>"011101001",
  62423=>"101011001",
  62424=>"000010101",
  62425=>"011011110",
  62426=>"111000000",
  62427=>"100001100",
  62428=>"101100010",
  62429=>"011001111",
  62430=>"100101000",
  62431=>"011110000",
  62432=>"110111111",
  62433=>"000101000",
  62434=>"100010001",
  62435=>"010011011",
  62436=>"001101100",
  62437=>"000101110",
  62438=>"101101110",
  62439=>"101001100",
  62440=>"000000010",
  62441=>"011011001",
  62442=>"101111000",
  62443=>"010001100",
  62444=>"011110101",
  62445=>"000101111",
  62446=>"001000000",
  62447=>"100100001",
  62448=>"000001001",
  62449=>"110001110",
  62450=>"101101101",
  62451=>"110110000",
  62452=>"100100010",
  62453=>"001001000",
  62454=>"101100100",
  62455=>"110001101",
  62456=>"100101011",
  62457=>"011000101",
  62458=>"010011100",
  62459=>"010000101",
  62460=>"100100010",
  62461=>"011011000",
  62462=>"101010000",
  62463=>"111010001",
  62464=>"010100000",
  62465=>"010011110",
  62466=>"011101000",
  62467=>"111000100",
  62468=>"011010101",
  62469=>"000100011",
  62470=>"000110000",
  62471=>"011111100",
  62472=>"111101010",
  62473=>"110110000",
  62474=>"010100010",
  62475=>"000100100",
  62476=>"110111100",
  62477=>"011100100",
  62478=>"100010011",
  62479=>"101110011",
  62480=>"110111111",
  62481=>"011100111",
  62482=>"001011111",
  62483=>"011000000",
  62484=>"111101100",
  62485=>"110101000",
  62486=>"111111011",
  62487=>"010111100",
  62488=>"111010101",
  62489=>"010101110",
  62490=>"111010100",
  62491=>"010110010",
  62492=>"111000010",
  62493=>"110111101",
  62494=>"010001111",
  62495=>"100111011",
  62496=>"101100100",
  62497=>"111110100",
  62498=>"100100101",
  62499=>"111100110",
  62500=>"111000100",
  62501=>"000000110",
  62502=>"000100100",
  62503=>"001100001",
  62504=>"100000010",
  62505=>"110001011",
  62506=>"010011100",
  62507=>"011001010",
  62508=>"100001100",
  62509=>"000111101",
  62510=>"111101101",
  62511=>"100101011",
  62512=>"110111111",
  62513=>"101111101",
  62514=>"001011011",
  62515=>"011000100",
  62516=>"110011110",
  62517=>"101001000",
  62518=>"011001010",
  62519=>"000110110",
  62520=>"000001100",
  62521=>"000110100",
  62522=>"101111100",
  62523=>"010110011",
  62524=>"011000000",
  62525=>"010111000",
  62526=>"000100111",
  62527=>"000000101",
  62528=>"111111000",
  62529=>"110010101",
  62530=>"101100110",
  62531=>"000101011",
  62532=>"000001100",
  62533=>"011111100",
  62534=>"101001001",
  62535=>"001110110",
  62536=>"000100101",
  62537=>"101000000",
  62538=>"111000101",
  62539=>"000011110",
  62540=>"001110110",
  62541=>"001100011",
  62542=>"011011100",
  62543=>"100000100",
  62544=>"100000100",
  62545=>"000010010",
  62546=>"011001000",
  62547=>"101101100",
  62548=>"110111010",
  62549=>"110010101",
  62550=>"111010100",
  62551=>"101100001",
  62552=>"100000000",
  62553=>"001101100",
  62554=>"111101001",
  62555=>"000011110",
  62556=>"000011010",
  62557=>"100100100",
  62558=>"100010000",
  62559=>"000001110",
  62560=>"100001001",
  62561=>"110101111",
  62562=>"011001111",
  62563=>"001010011",
  62564=>"101100100",
  62565=>"011001100",
  62566=>"111000111",
  62567=>"111011100",
  62568=>"001111111",
  62569=>"110111100",
  62570=>"100100101",
  62571=>"000011100",
  62572=>"011011000",
  62573=>"101100000",
  62574=>"100101010",
  62575=>"010000001",
  62576=>"000001101",
  62577=>"000000101",
  62578=>"000011101",
  62579=>"111011100",
  62580=>"000101011",
  62581=>"000010011",
  62582=>"111001111",
  62583=>"101100001",
  62584=>"110100100",
  62585=>"110111011",
  62586=>"010110111",
  62587=>"110001001",
  62588=>"010010100",
  62589=>"001101000",
  62590=>"110011000",
  62591=>"011010101",
  62592=>"110101100",
  62593=>"000001011",
  62594=>"000100010",
  62595=>"101000011",
  62596=>"101000000",
  62597=>"011100011",
  62598=>"000111001",
  62599=>"011010011",
  62600=>"011011011",
  62601=>"011101011",
  62602=>"111101010",
  62603=>"111011101",
  62604=>"010011111",
  62605=>"111010001",
  62606=>"100111101",
  62607=>"111000000",
  62608=>"000001100",
  62609=>"111000100",
  62610=>"010111110",
  62611=>"001101010",
  62612=>"110010110",
  62613=>"100110010",
  62614=>"101001110",
  62615=>"100111001",
  62616=>"101101011",
  62617=>"100100001",
  62618=>"011101101",
  62619=>"001110001",
  62620=>"000110111",
  62621=>"010100111",
  62622=>"101000001",
  62623=>"110001011",
  62624=>"110011110",
  62625=>"001110101",
  62626=>"001001001",
  62627=>"101000110",
  62628=>"011101011",
  62629=>"000111100",
  62630=>"011010101",
  62631=>"111101111",
  62632=>"111101101",
  62633=>"011001001",
  62634=>"111100101",
  62635=>"000000111",
  62636=>"101000000",
  62637=>"001110011",
  62638=>"000110010",
  62639=>"010100011",
  62640=>"101000110",
  62641=>"111110100",
  62642=>"000111111",
  62643=>"000000000",
  62644=>"000100111",
  62645=>"001010000",
  62646=>"011101101",
  62647=>"010100000",
  62648=>"000100110",
  62649=>"101000101",
  62650=>"100001000",
  62651=>"000010010",
  62652=>"110110000",
  62653=>"101010010",
  62654=>"101011111",
  62655=>"100010011",
  62656=>"110110011",
  62657=>"110111011",
  62658=>"001011001",
  62659=>"000000011",
  62660=>"111010111",
  62661=>"000011110",
  62662=>"101011101",
  62663=>"010001000",
  62664=>"110100111",
  62665=>"011101011",
  62666=>"001010110",
  62667=>"000100111",
  62668=>"011010111",
  62669=>"100000111",
  62670=>"101000000",
  62671=>"110101001",
  62672=>"110000110",
  62673=>"101101000",
  62674=>"100101101",
  62675=>"000111000",
  62676=>"110110000",
  62677=>"000011010",
  62678=>"010010010",
  62679=>"001110111",
  62680=>"000101111",
  62681=>"111100110",
  62682=>"001100000",
  62683=>"001001100",
  62684=>"001011110",
  62685=>"000011000",
  62686=>"011001011",
  62687=>"011001000",
  62688=>"101100100",
  62689=>"010011100",
  62690=>"101100010",
  62691=>"111000001",
  62692=>"110001001",
  62693=>"001001110",
  62694=>"001101110",
  62695=>"111111101",
  62696=>"111010000",
  62697=>"010101111",
  62698=>"000100011",
  62699=>"111011000",
  62700=>"001111001",
  62701=>"111011001",
  62702=>"001011000",
  62703=>"000000100",
  62704=>"100110001",
  62705=>"000111111",
  62706=>"010001000",
  62707=>"000000110",
  62708=>"101001011",
  62709=>"110011110",
  62710=>"001100110",
  62711=>"101110110",
  62712=>"000101100",
  62713=>"100000110",
  62714=>"110000000",
  62715=>"001010010",
  62716=>"110010011",
  62717=>"011011011",
  62718=>"011010011",
  62719=>"001000001",
  62720=>"111110011",
  62721=>"101010010",
  62722=>"010010110",
  62723=>"001100010",
  62724=>"110110000",
  62725=>"100100001",
  62726=>"001010100",
  62727=>"011101101",
  62728=>"000111110",
  62729=>"111100111",
  62730=>"101011000",
  62731=>"110000110",
  62732=>"010000110",
  62733=>"011100110",
  62734=>"011011011",
  62735=>"001010010",
  62736=>"011110001",
  62737=>"011100101",
  62738=>"000001101",
  62739=>"001110001",
  62740=>"000110000",
  62741=>"011100000",
  62742=>"000011000",
  62743=>"000011110",
  62744=>"111000101",
  62745=>"110001010",
  62746=>"111010000",
  62747=>"011000001",
  62748=>"001110110",
  62749=>"001001111",
  62750=>"011010100",
  62751=>"010110100",
  62752=>"001000000",
  62753=>"111111011",
  62754=>"101000010",
  62755=>"001001111",
  62756=>"101010011",
  62757=>"010111110",
  62758=>"111000010",
  62759=>"000010000",
  62760=>"101001000",
  62761=>"110001100",
  62762=>"100000000",
  62763=>"010110111",
  62764=>"010010010",
  62765=>"000100111",
  62766=>"111100101",
  62767=>"000110010",
  62768=>"000111100",
  62769=>"011110001",
  62770=>"110111111",
  62771=>"011100111",
  62772=>"111111011",
  62773=>"101110101",
  62774=>"001011001",
  62775=>"010101110",
  62776=>"111111100",
  62777=>"001001010",
  62778=>"010100000",
  62779=>"011001100",
  62780=>"100000110",
  62781=>"111111111",
  62782=>"111011100",
  62783=>"110001000",
  62784=>"111100110",
  62785=>"111111111",
  62786=>"000100001",
  62787=>"010110000",
  62788=>"000011010",
  62789=>"101001101",
  62790=>"100010101",
  62791=>"100111111",
  62792=>"100010000",
  62793=>"110101010",
  62794=>"011001100",
  62795=>"001111111",
  62796=>"011000010",
  62797=>"011101011",
  62798=>"101111111",
  62799=>"100001010",
  62800=>"100100111",
  62801=>"000110111",
  62802=>"000111111",
  62803=>"101001111",
  62804=>"111111111",
  62805=>"000101000",
  62806=>"101100001",
  62807=>"010010101",
  62808=>"101001101",
  62809=>"001111010",
  62810=>"100000100",
  62811=>"100100011",
  62812=>"001111101",
  62813=>"001101001",
  62814=>"000011111",
  62815=>"010101100",
  62816=>"111110000",
  62817=>"001000011",
  62818=>"101100111",
  62819=>"010000011",
  62820=>"010100111",
  62821=>"101100001",
  62822=>"111111100",
  62823=>"100000001",
  62824=>"111110111",
  62825=>"001000010",
  62826=>"010010100",
  62827=>"110110011",
  62828=>"001111101",
  62829=>"001000111",
  62830=>"100001011",
  62831=>"001011100",
  62832=>"100111001",
  62833=>"010011011",
  62834=>"001101000",
  62835=>"100011100",
  62836=>"000110000",
  62837=>"110110010",
  62838=>"111110111",
  62839=>"000110100",
  62840=>"010001100",
  62841=>"110110001",
  62842=>"001010001",
  62843=>"100011100",
  62844=>"011110101",
  62845=>"110101011",
  62846=>"010010001",
  62847=>"111011101",
  62848=>"000011001",
  62849=>"011101001",
  62850=>"010010011",
  62851=>"110100100",
  62852=>"001110001",
  62853=>"111000001",
  62854=>"100110000",
  62855=>"111110101",
  62856=>"100111011",
  62857=>"000001110",
  62858=>"010010111",
  62859=>"101100101",
  62860=>"011001010",
  62861=>"101001111",
  62862=>"111110000",
  62863=>"101010011",
  62864=>"101000001",
  62865=>"111001010",
  62866=>"100111000",
  62867=>"000100001",
  62868=>"101001011",
  62869=>"110000010",
  62870=>"101001011",
  62871=>"101010100",
  62872=>"001101011",
  62873=>"101001100",
  62874=>"110110100",
  62875=>"100000100",
  62876=>"110110010",
  62877=>"010011011",
  62878=>"111111010",
  62879=>"010110111",
  62880=>"001000100",
  62881=>"000011111",
  62882=>"111100011",
  62883=>"011110001",
  62884=>"101111110",
  62885=>"011001001",
  62886=>"101111101",
  62887=>"111000111",
  62888=>"001111110",
  62889=>"100101110",
  62890=>"110101111",
  62891=>"010101100",
  62892=>"010010101",
  62893=>"010000010",
  62894=>"010110110",
  62895=>"000010111",
  62896=>"100100100",
  62897=>"010111011",
  62898=>"010111000",
  62899=>"111001100",
  62900=>"100110110",
  62901=>"101001110",
  62902=>"011000011",
  62903=>"011000010",
  62904=>"111000101",
  62905=>"010101101",
  62906=>"001100110",
  62907=>"010111011",
  62908=>"010000100",
  62909=>"011010010",
  62910=>"011101110",
  62911=>"000011100",
  62912=>"110001011",
  62913=>"111101111",
  62914=>"011111101",
  62915=>"110110111",
  62916=>"100100010",
  62917=>"110011111",
  62918=>"101000111",
  62919=>"011101001",
  62920=>"101010100",
  62921=>"101011111",
  62922=>"111111001",
  62923=>"011101111",
  62924=>"000110011",
  62925=>"001100111",
  62926=>"010011110",
  62927=>"101101110",
  62928=>"010000110",
  62929=>"110101101",
  62930=>"100100000",
  62931=>"000000000",
  62932=>"110010010",
  62933=>"010101010",
  62934=>"000000010",
  62935=>"001101011",
  62936=>"010111010",
  62937=>"000000001",
  62938=>"101000110",
  62939=>"011101100",
  62940=>"101111100",
  62941=>"111101101",
  62942=>"111000111",
  62943=>"011010000",
  62944=>"000001101",
  62945=>"110000100",
  62946=>"000111101",
  62947=>"011011010",
  62948=>"110100110",
  62949=>"111100100",
  62950=>"110111010",
  62951=>"100111100",
  62952=>"110011000",
  62953=>"000100010",
  62954=>"000000010",
  62955=>"010111101",
  62956=>"110100001",
  62957=>"100100011",
  62958=>"001110000",
  62959=>"001010111",
  62960=>"010000101",
  62961=>"111000111",
  62962=>"110000011",
  62963=>"100010001",
  62964=>"110101000",
  62965=>"001101100",
  62966=>"001110000",
  62967=>"010110110",
  62968=>"101101101",
  62969=>"100101101",
  62970=>"001111111",
  62971=>"101001100",
  62972=>"101111111",
  62973=>"001010100",
  62974=>"000011000",
  62975=>"110000010",
  62976=>"111111100",
  62977=>"000110000",
  62978=>"001101101",
  62979=>"001001001",
  62980=>"110101010",
  62981=>"100101001",
  62982=>"101100011",
  62983=>"010111010",
  62984=>"101010110",
  62985=>"011110000",
  62986=>"111111110",
  62987=>"011010010",
  62988=>"101101100",
  62989=>"001110100",
  62990=>"101100100",
  62991=>"111100111",
  62992=>"011101010",
  62993=>"110100100",
  62994=>"000010010",
  62995=>"100010001",
  62996=>"011000101",
  62997=>"010100000",
  62998=>"010011010",
  62999=>"101101010",
  63000=>"110000010",
  63001=>"001001110",
  63002=>"000010001",
  63003=>"110111001",
  63004=>"001100101",
  63005=>"000000010",
  63006=>"111010110",
  63007=>"000011011",
  63008=>"110110011",
  63009=>"101111000",
  63010=>"000000111",
  63011=>"000111011",
  63012=>"110111101",
  63013=>"011101110",
  63014=>"110101100",
  63015=>"111000100",
  63016=>"111010001",
  63017=>"000000000",
  63018=>"101111110",
  63019=>"100000010",
  63020=>"011010000",
  63021=>"110011110",
  63022=>"000101001",
  63023=>"000010010",
  63024=>"100010111",
  63025=>"111111101",
  63026=>"100111101",
  63027=>"010001111",
  63028=>"011100010",
  63029=>"010111010",
  63030=>"001100011",
  63031=>"011011010",
  63032=>"010010111",
  63033=>"111101100",
  63034=>"010101100",
  63035=>"101111111",
  63036=>"100010100",
  63037=>"100110100",
  63038=>"111111100",
  63039=>"000101011",
  63040=>"011110011",
  63041=>"011101110",
  63042=>"111010010",
  63043=>"010100100",
  63044=>"110111001",
  63045=>"101101000",
  63046=>"010110010",
  63047=>"111001011",
  63048=>"100000010",
  63049=>"011100101",
  63050=>"111000101",
  63051=>"111000100",
  63052=>"001111010",
  63053=>"101100110",
  63054=>"011000101",
  63055=>"111010010",
  63056=>"111000100",
  63057=>"100111010",
  63058=>"100100101",
  63059=>"111000101",
  63060=>"001110111",
  63061=>"101100010",
  63062=>"000001111",
  63063=>"010111111",
  63064=>"010001100",
  63065=>"110011010",
  63066=>"101111011",
  63067=>"000001111",
  63068=>"101011110",
  63069=>"001110100",
  63070=>"001101111",
  63071=>"001000001",
  63072=>"011001011",
  63073=>"110010011",
  63074=>"000110011",
  63075=>"110011000",
  63076=>"100111111",
  63077=>"010101011",
  63078=>"101011111",
  63079=>"101101111",
  63080=>"000000110",
  63081=>"101111000",
  63082=>"011111111",
  63083=>"000110001",
  63084=>"101111010",
  63085=>"010101001",
  63086=>"000111111",
  63087=>"011101111",
  63088=>"000110110",
  63089=>"100101010",
  63090=>"111001001",
  63091=>"011010100",
  63092=>"101101111",
  63093=>"111100010",
  63094=>"001000010",
  63095=>"000111011",
  63096=>"111101010",
  63097=>"000110100",
  63098=>"101110001",
  63099=>"000100010",
  63100=>"000001101",
  63101=>"101001000",
  63102=>"100101101",
  63103=>"011110101",
  63104=>"100000100",
  63105=>"110001111",
  63106=>"010011101",
  63107=>"000010011",
  63108=>"001010111",
  63109=>"000110010",
  63110=>"110111111",
  63111=>"011101000",
  63112=>"100001001",
  63113=>"001001111",
  63114=>"111101011",
  63115=>"100000010",
  63116=>"001101000",
  63117=>"100000000",
  63118=>"100000101",
  63119=>"110000111",
  63120=>"110110111",
  63121=>"111010000",
  63122=>"110010110",
  63123=>"010101100",
  63124=>"001101100",
  63125=>"111100001",
  63126=>"101100011",
  63127=>"110010110",
  63128=>"101000110",
  63129=>"101111010",
  63130=>"110101101",
  63131=>"001100000",
  63132=>"110101100",
  63133=>"010000100",
  63134=>"101110100",
  63135=>"110000101",
  63136=>"010101110",
  63137=>"111101101",
  63138=>"010011110",
  63139=>"100110101",
  63140=>"100110111",
  63141=>"000011111",
  63142=>"010011101",
  63143=>"001000001",
  63144=>"010000000",
  63145=>"000110001",
  63146=>"101101111",
  63147=>"101100011",
  63148=>"010101010",
  63149=>"001111111",
  63150=>"111000001",
  63151=>"110100000",
  63152=>"000110010",
  63153=>"011010011",
  63154=>"000111000",
  63155=>"010001010",
  63156=>"100101100",
  63157=>"010110011",
  63158=>"011010000",
  63159=>"011011010",
  63160=>"001000000",
  63161=>"001000100",
  63162=>"000100001",
  63163=>"110100101",
  63164=>"110100101",
  63165=>"100010110",
  63166=>"011001000",
  63167=>"101100100",
  63168=>"010110110",
  63169=>"000110110",
  63170=>"101101110",
  63171=>"010010101",
  63172=>"000001110",
  63173=>"010000110",
  63174=>"110111010",
  63175=>"000110111",
  63176=>"011010010",
  63177=>"111011100",
  63178=>"100111010",
  63179=>"100101111",
  63180=>"101100111",
  63181=>"010111110",
  63182=>"001110110",
  63183=>"101110011",
  63184=>"010001111",
  63185=>"000110100",
  63186=>"110100110",
  63187=>"100001011",
  63188=>"000011100",
  63189=>"000011110",
  63190=>"100100011",
  63191=>"100110001",
  63192=>"011101011",
  63193=>"010011010",
  63194=>"010010101",
  63195=>"111011001",
  63196=>"100010011",
  63197=>"001110101",
  63198=>"010101100",
  63199=>"001000000",
  63200=>"010001111",
  63201=>"110010101",
  63202=>"110100101",
  63203=>"001011110",
  63204=>"001101110",
  63205=>"011111111",
  63206=>"000101111",
  63207=>"000001000",
  63208=>"101000100",
  63209=>"010001010",
  63210=>"100011100",
  63211=>"100000101",
  63212=>"000000001",
  63213=>"001010101",
  63214=>"000101100",
  63215=>"000001000",
  63216=>"000110010",
  63217=>"110011001",
  63218=>"100110111",
  63219=>"001101100",
  63220=>"010001100",
  63221=>"011011010",
  63222=>"000011100",
  63223=>"101000011",
  63224=>"100001001",
  63225=>"110100001",
  63226=>"110011111",
  63227=>"001110001",
  63228=>"110101101",
  63229=>"000001101",
  63230=>"011001110",
  63231=>"010110000",
  63232=>"000011011",
  63233=>"010110010",
  63234=>"110010100",
  63235=>"001011111",
  63236=>"010011000",
  63237=>"111000001",
  63238=>"011100001",
  63239=>"011100010",
  63240=>"101111111",
  63241=>"101010001",
  63242=>"010011110",
  63243=>"111101001",
  63244=>"110010000",
  63245=>"100011011",
  63246=>"000110000",
  63247=>"011111000",
  63248=>"110101011",
  63249=>"011110111",
  63250=>"001000001",
  63251=>"110001101",
  63252=>"011010100",
  63253=>"101001010",
  63254=>"011010010",
  63255=>"001100011",
  63256=>"101101101",
  63257=>"000110000",
  63258=>"000011110",
  63259=>"011010010",
  63260=>"100110001",
  63261=>"110100000",
  63262=>"110100100",
  63263=>"011010001",
  63264=>"101100101",
  63265=>"001111111",
  63266=>"010011011",
  63267=>"101110101",
  63268=>"011001010",
  63269=>"100111010",
  63270=>"100000100",
  63271=>"011110010",
  63272=>"010111100",
  63273=>"100010111",
  63274=>"111011010",
  63275=>"101101010",
  63276=>"111011001",
  63277=>"111111111",
  63278=>"100000000",
  63279=>"010111011",
  63280=>"011010111",
  63281=>"000010001",
  63282=>"110001010",
  63283=>"000001010",
  63284=>"000100000",
  63285=>"111011001",
  63286=>"001111101",
  63287=>"101011001",
  63288=>"010101001",
  63289=>"011110011",
  63290=>"001000101",
  63291=>"110110100",
  63292=>"111010110",
  63293=>"101111110",
  63294=>"100011001",
  63295=>"100100100",
  63296=>"101100111",
  63297=>"100001001",
  63298=>"001001001",
  63299=>"010100001",
  63300=>"110110011",
  63301=>"010011111",
  63302=>"001000111",
  63303=>"111001011",
  63304=>"100011110",
  63305=>"000010011",
  63306=>"101000100",
  63307=>"110101110",
  63308=>"001111111",
  63309=>"011100110",
  63310=>"101011001",
  63311=>"100111100",
  63312=>"000000100",
  63313=>"111100010",
  63314=>"011010001",
  63315=>"010000001",
  63316=>"100110111",
  63317=>"101101000",
  63318=>"011011000",
  63319=>"111101001",
  63320=>"001001101",
  63321=>"000111111",
  63322=>"100101010",
  63323=>"010101011",
  63324=>"001010010",
  63325=>"011010010",
  63326=>"010000101",
  63327=>"000010110",
  63328=>"000011011",
  63329=>"010100000",
  63330=>"100000001",
  63331=>"101110111",
  63332=>"010000100",
  63333=>"011101000",
  63334=>"000001010",
  63335=>"001111100",
  63336=>"111010111",
  63337=>"110110000",
  63338=>"101000111",
  63339=>"100011111",
  63340=>"110001101",
  63341=>"111001101",
  63342=>"111100101",
  63343=>"101101101",
  63344=>"100001000",
  63345=>"001100111",
  63346=>"110110000",
  63347=>"111110100",
  63348=>"000001101",
  63349=>"010011111",
  63350=>"100001111",
  63351=>"001001100",
  63352=>"110000100",
  63353=>"011010011",
  63354=>"010110001",
  63355=>"000011110",
  63356=>"110100110",
  63357=>"100011101",
  63358=>"110110100",
  63359=>"110011110",
  63360=>"010101111",
  63361=>"100001001",
  63362=>"101111001",
  63363=>"101010011",
  63364=>"010001001",
  63365=>"111011011",
  63366=>"101001000",
  63367=>"110001111",
  63368=>"000000101",
  63369=>"100101010",
  63370=>"001111110",
  63371=>"111101001",
  63372=>"000111101",
  63373=>"111101110",
  63374=>"010110100",
  63375=>"100001101",
  63376=>"001011101",
  63377=>"000100010",
  63378=>"010000110",
  63379=>"001011011",
  63380=>"111110100",
  63381=>"011110111",
  63382=>"011010110",
  63383=>"001100111",
  63384=>"110010101",
  63385=>"001000100",
  63386=>"001011110",
  63387=>"001111101",
  63388=>"011000100",
  63389=>"011101001",
  63390=>"100100100",
  63391=>"011101101",
  63392=>"100000100",
  63393=>"111111101",
  63394=>"000011111",
  63395=>"111000011",
  63396=>"110001011",
  63397=>"111111111",
  63398=>"100001001",
  63399=>"010001110",
  63400=>"110011001",
  63401=>"111101111",
  63402=>"011110001",
  63403=>"001010101",
  63404=>"000000000",
  63405=>"010101100",
  63406=>"000101000",
  63407=>"101100101",
  63408=>"101001111",
  63409=>"100000100",
  63410=>"111010001",
  63411=>"100100100",
  63412=>"110111100",
  63413=>"101011100",
  63414=>"100001101",
  63415=>"010110111",
  63416=>"000000100",
  63417=>"000000110",
  63418=>"010011100",
  63419=>"110101101",
  63420=>"001110000",
  63421=>"000011000",
  63422=>"111001011",
  63423=>"110111111",
  63424=>"111111101",
  63425=>"111110111",
  63426=>"001100010",
  63427=>"101010110",
  63428=>"101101000",
  63429=>"110101111",
  63430=>"101011011",
  63431=>"110110000",
  63432=>"100010000",
  63433=>"110110000",
  63434=>"010101111",
  63435=>"101000101",
  63436=>"110001011",
  63437=>"101100100",
  63438=>"010001111",
  63439=>"110011010",
  63440=>"110010100",
  63441=>"111110011",
  63442=>"100100011",
  63443=>"000111111",
  63444=>"000000000",
  63445=>"000100010",
  63446=>"000100010",
  63447=>"100000110",
  63448=>"010001101",
  63449=>"101001001",
  63450=>"101111000",
  63451=>"101111001",
  63452=>"111111110",
  63453=>"000010100",
  63454=>"111111101",
  63455=>"010101111",
  63456=>"001001110",
  63457=>"111101010",
  63458=>"000111100",
  63459=>"100011000",
  63460=>"110011000",
  63461=>"100101000",
  63462=>"011101110",
  63463=>"111110001",
  63464=>"101100101",
  63465=>"001111000",
  63466=>"000111011",
  63467=>"111101111",
  63468=>"000110101",
  63469=>"110101100",
  63470=>"110100110",
  63471=>"001010010",
  63472=>"000000001",
  63473=>"100010010",
  63474=>"000101110",
  63475=>"001001101",
  63476=>"010100000",
  63477=>"111000110",
  63478=>"010010011",
  63479=>"111110111",
  63480=>"010010110",
  63481=>"100000111",
  63482=>"101001010",
  63483=>"011001100",
  63484=>"101100000",
  63485=>"000010010",
  63486=>"100110110",
  63487=>"001001000",
  63488=>"000000010",
  63489=>"110100000",
  63490=>"111110100",
  63491=>"110111010",
  63492=>"100011110",
  63493=>"001011010",
  63494=>"000001101",
  63495=>"111111101",
  63496=>"111001101",
  63497=>"000110000",
  63498=>"110110100",
  63499=>"101001011",
  63500=>"101011101",
  63501=>"000100101",
  63502=>"110000100",
  63503=>"000101010",
  63504=>"011100011",
  63505=>"100101101",
  63506=>"011101110",
  63507=>"010100000",
  63508=>"100100111",
  63509=>"111111111",
  63510=>"101111011",
  63511=>"011010000",
  63512=>"001110100",
  63513=>"001010110",
  63514=>"011001110",
  63515=>"001011011",
  63516=>"101101111",
  63517=>"100010110",
  63518=>"011011000",
  63519=>"001110011",
  63520=>"000001110",
  63521=>"100101111",
  63522=>"001100100",
  63523=>"110110100",
  63524=>"111011010",
  63525=>"100010001",
  63526=>"001010101",
  63527=>"011001110",
  63528=>"111100101",
  63529=>"000110100",
  63530=>"101000001",
  63531=>"100111011",
  63532=>"000000000",
  63533=>"011101010",
  63534=>"111011001",
  63535=>"010101000",
  63536=>"111100011",
  63537=>"010010110",
  63538=>"000001101",
  63539=>"100111111",
  63540=>"111001100",
  63541=>"100110000",
  63542=>"110100110",
  63543=>"110110010",
  63544=>"001001111",
  63545=>"011010100",
  63546=>"000001110",
  63547=>"000101011",
  63548=>"001110101",
  63549=>"100001010",
  63550=>"011110011",
  63551=>"111001111",
  63552=>"000001000",
  63553=>"011000110",
  63554=>"101111101",
  63555=>"101110110",
  63556=>"011001001",
  63557=>"001111111",
  63558=>"000011011",
  63559=>"000111101",
  63560=>"100110010",
  63561=>"001011000",
  63562=>"001110101",
  63563=>"000011101",
  63564=>"000011010",
  63565=>"000101011",
  63566=>"000010100",
  63567=>"000001011",
  63568=>"101001111",
  63569=>"000011011",
  63570=>"110100000",
  63571=>"010110010",
  63572=>"010100101",
  63573=>"101000111",
  63574=>"111111001",
  63575=>"010000010",
  63576=>"010001001",
  63577=>"010101101",
  63578=>"101001111",
  63579=>"101010110",
  63580=>"000101000",
  63581=>"101010001",
  63582=>"101111101",
  63583=>"010001110",
  63584=>"110100000",
  63585=>"000000000",
  63586=>"000111010",
  63587=>"001010011",
  63588=>"100111111",
  63589=>"100001000",
  63590=>"111111010",
  63591=>"111100111",
  63592=>"011001010",
  63593=>"101011001",
  63594=>"000100110",
  63595=>"100111010",
  63596=>"001001100",
  63597=>"100011011",
  63598=>"000101010",
  63599=>"100101101",
  63600=>"010001111",
  63601=>"000011101",
  63602=>"010111011",
  63603=>"001011110",
  63604=>"101011100",
  63605=>"001111011",
  63606=>"110000110",
  63607=>"011100111",
  63608=>"000000111",
  63609=>"011000001",
  63610=>"101110101",
  63611=>"000100011",
  63612=>"011000101",
  63613=>"010111010",
  63614=>"111111011",
  63615=>"010001001",
  63616=>"100110001",
  63617=>"101000111",
  63618=>"100000100",
  63619=>"111110100",
  63620=>"100100000",
  63621=>"101101011",
  63622=>"101011110",
  63623=>"101100100",
  63624=>"010010011",
  63625=>"100110110",
  63626=>"011000000",
  63627=>"111111100",
  63628=>"101100111",
  63629=>"101011000",
  63630=>"000101001",
  63631=>"101100110",
  63632=>"100101100",
  63633=>"001010001",
  63634=>"010100101",
  63635=>"111010100",
  63636=>"101101111",
  63637=>"011101001",
  63638=>"111111100",
  63639=>"101011110",
  63640=>"111000001",
  63641=>"101011010",
  63642=>"011110010",
  63643=>"111001111",
  63644=>"010100100",
  63645=>"000111001",
  63646=>"000001000",
  63647=>"000000011",
  63648=>"101110111",
  63649=>"101000011",
  63650=>"101100010",
  63651=>"010000101",
  63652=>"000110111",
  63653=>"001111100",
  63654=>"101001011",
  63655=>"000000001",
  63656=>"000011100",
  63657=>"000100000",
  63658=>"101100111",
  63659=>"000100000",
  63660=>"001011001",
  63661=>"111110111",
  63662=>"110010001",
  63663=>"110110100",
  63664=>"010010001",
  63665=>"010111010",
  63666=>"011011011",
  63667=>"001000111",
  63668=>"010100010",
  63669=>"100000111",
  63670=>"110100011",
  63671=>"110010110",
  63672=>"100000101",
  63673=>"000110000",
  63674=>"000011101",
  63675=>"111011001",
  63676=>"101100011",
  63677=>"101110111",
  63678=>"011001110",
  63679=>"110001000",
  63680=>"000010100",
  63681=>"010101101",
  63682=>"000110001",
  63683=>"111110111",
  63684=>"111110110",
  63685=>"111111011",
  63686=>"001110101",
  63687=>"000010001",
  63688=>"010101101",
  63689=>"001001101",
  63690=>"110000111",
  63691=>"111101011",
  63692=>"001111110",
  63693=>"110001010",
  63694=>"011000000",
  63695=>"001001111",
  63696=>"101110011",
  63697=>"000011011",
  63698=>"110001010",
  63699=>"101111010",
  63700=>"010110111",
  63701=>"110010100",
  63702=>"000110110",
  63703=>"110011101",
  63704=>"000011010",
  63705=>"010100100",
  63706=>"011101110",
  63707=>"010001000",
  63708=>"010100100",
  63709=>"000100000",
  63710=>"011001111",
  63711=>"000101010",
  63712=>"010010111",
  63713=>"000000101",
  63714=>"101101001",
  63715=>"000000010",
  63716=>"101111011",
  63717=>"010010111",
  63718=>"010010010",
  63719=>"101101011",
  63720=>"000000000",
  63721=>"101010111",
  63722=>"001110110",
  63723=>"011100000",
  63724=>"011101010",
  63725=>"010000010",
  63726=>"001100010",
  63727=>"101010101",
  63728=>"100011111",
  63729=>"001001100",
  63730=>"111001100",
  63731=>"110011010",
  63732=>"110111001",
  63733=>"011010011",
  63734=>"011101010",
  63735=>"010001101",
  63736=>"000000010",
  63737=>"111001010",
  63738=>"011111000",
  63739=>"000100011",
  63740=>"000101100",
  63741=>"010000001",
  63742=>"100100000",
  63743=>"000000110",
  63744=>"001110111",
  63745=>"111110001",
  63746=>"110101110",
  63747=>"001000011",
  63748=>"111011010",
  63749=>"000010010",
  63750=>"111111100",
  63751=>"010101110",
  63752=>"011100010",
  63753=>"001100100",
  63754=>"100101100",
  63755=>"100001111",
  63756=>"111000010",
  63757=>"111100111",
  63758=>"110010000",
  63759=>"011010110",
  63760=>"000011111",
  63761=>"001101101",
  63762=>"101100001",
  63763=>"110111011",
  63764=>"101100010",
  63765=>"100001110",
  63766=>"000110011",
  63767=>"010111100",
  63768=>"111000110",
  63769=>"110110110",
  63770=>"110100001",
  63771=>"111000011",
  63772=>"111100101",
  63773=>"001100101",
  63774=>"101100111",
  63775=>"111100011",
  63776=>"011001111",
  63777=>"001000110",
  63778=>"001001101",
  63779=>"001111111",
  63780=>"111101100",
  63781=>"111000001",
  63782=>"010111111",
  63783=>"000110010",
  63784=>"001101011",
  63785=>"101001101",
  63786=>"111011111",
  63787=>"100111000",
  63788=>"111101000",
  63789=>"110000000",
  63790=>"000101010",
  63791=>"010011110",
  63792=>"110110101",
  63793=>"000001001",
  63794=>"110110100",
  63795=>"101111001",
  63796=>"001000001",
  63797=>"100000000",
  63798=>"100110110",
  63799=>"110111000",
  63800=>"100111011",
  63801=>"011000001",
  63802=>"000010000",
  63803=>"010010010",
  63804=>"011010000",
  63805=>"000101100",
  63806=>"111111011",
  63807=>"101100000",
  63808=>"000111011",
  63809=>"110011010",
  63810=>"110100010",
  63811=>"011100101",
  63812=>"011010011",
  63813=>"101010011",
  63814=>"010000101",
  63815=>"001001010",
  63816=>"100110110",
  63817=>"101010010",
  63818=>"010100101",
  63819=>"011001100",
  63820=>"101101100",
  63821=>"000011111",
  63822=>"110101010",
  63823=>"000101001",
  63824=>"010000100",
  63825=>"100011111",
  63826=>"110001011",
  63827=>"100000000",
  63828=>"001011111",
  63829=>"101101101",
  63830=>"110100111",
  63831=>"100000100",
  63832=>"111110000",
  63833=>"100100011",
  63834=>"010111110",
  63835=>"111101101",
  63836=>"001100001",
  63837=>"100000101",
  63838=>"000000011",
  63839=>"111010011",
  63840=>"101011100",
  63841=>"000111000",
  63842=>"110100100",
  63843=>"011111011",
  63844=>"111110011",
  63845=>"110101100",
  63846=>"011010011",
  63847=>"000111100",
  63848=>"000100110",
  63849=>"110110000",
  63850=>"100001000",
  63851=>"001101010",
  63852=>"011110100",
  63853=>"110000001",
  63854=>"101010100",
  63855=>"110100001",
  63856=>"110010010",
  63857=>"101010010",
  63858=>"100100011",
  63859=>"001000101",
  63860=>"111101110",
  63861=>"100011111",
  63862=>"010100000",
  63863=>"111110010",
  63864=>"001001100",
  63865=>"000011110",
  63866=>"101011110",
  63867=>"000001011",
  63868=>"010111101",
  63869=>"100100010",
  63870=>"011111011",
  63871=>"100101011",
  63872=>"011100101",
  63873=>"011010010",
  63874=>"110110000",
  63875=>"100111100",
  63876=>"000100110",
  63877=>"101101111",
  63878=>"011010010",
  63879=>"001101001",
  63880=>"010111110",
  63881=>"010110001",
  63882=>"010011110",
  63883=>"000000010",
  63884=>"101110110",
  63885=>"100101101",
  63886=>"010000100",
  63887=>"010001001",
  63888=>"101101011",
  63889=>"100101011",
  63890=>"110111100",
  63891=>"000111001",
  63892=>"001001001",
  63893=>"011000000",
  63894=>"000011100",
  63895=>"011101001",
  63896=>"000111010",
  63897=>"000100000",
  63898=>"101000110",
  63899=>"000100010",
  63900=>"100010010",
  63901=>"011011111",
  63902=>"111001111",
  63903=>"010110101",
  63904=>"001010010",
  63905=>"011111111",
  63906=>"011001110",
  63907=>"011100101",
  63908=>"001001000",
  63909=>"111111011",
  63910=>"010110011",
  63911=>"101101110",
  63912=>"010011101",
  63913=>"000000000",
  63914=>"110001000",
  63915=>"111111101",
  63916=>"000110011",
  63917=>"111000011",
  63918=>"010111111",
  63919=>"110110110",
  63920=>"000101000",
  63921=>"100001000",
  63922=>"110110111",
  63923=>"000001101",
  63924=>"000100110",
  63925=>"111000111",
  63926=>"100100001",
  63927=>"011100100",
  63928=>"101011000",
  63929=>"000010011",
  63930=>"101000011",
  63931=>"010110000",
  63932=>"011011000",
  63933=>"111001110",
  63934=>"110111101",
  63935=>"111011110",
  63936=>"000010101",
  63937=>"101111101",
  63938=>"110011011",
  63939=>"110110000",
  63940=>"010101000",
  63941=>"011101000",
  63942=>"100000100",
  63943=>"011110111",
  63944=>"111011111",
  63945=>"110011110",
  63946=>"010001001",
  63947=>"110101111",
  63948=>"001011100",
  63949=>"000101101",
  63950=>"110111000",
  63951=>"111010010",
  63952=>"000110111",
  63953=>"101111110",
  63954=>"110011111",
  63955=>"011000110",
  63956=>"011100111",
  63957=>"011000000",
  63958=>"101000111",
  63959=>"011010101",
  63960=>"001100000",
  63961=>"011011000",
  63962=>"110101001",
  63963=>"111011100",
  63964=>"100011101",
  63965=>"111111001",
  63966=>"100001000",
  63967=>"000000001",
  63968=>"000111110",
  63969=>"110001110",
  63970=>"010011101",
  63971=>"110110011",
  63972=>"101010101",
  63973=>"100110000",
  63974=>"010111110",
  63975=>"010010101",
  63976=>"001110010",
  63977=>"000100110",
  63978=>"010100101",
  63979=>"000110111",
  63980=>"111101011",
  63981=>"001110111",
  63982=>"100100110",
  63983=>"101101011",
  63984=>"110101011",
  63985=>"011111100",
  63986=>"010111001",
  63987=>"001001001",
  63988=>"001101000",
  63989=>"000100111",
  63990=>"111111011",
  63991=>"100100100",
  63992=>"001011110",
  63993=>"100101100",
  63994=>"110000001",
  63995=>"011110100",
  63996=>"010110100",
  63997=>"001100111",
  63998=>"111110010",
  63999=>"111011010",
  64000=>"000010000",
  64001=>"101001010",
  64002=>"100000000",
  64003=>"100101111",
  64004=>"010010001",
  64005=>"100001000",
  64006=>"110010111",
  64007=>"000100111",
  64008=>"001100010",
  64009=>"101111111",
  64010=>"100010111",
  64011=>"101011001",
  64012=>"010001110",
  64013=>"110011000",
  64014=>"000000000",
  64015=>"001110001",
  64016=>"111011100",
  64017=>"000011111",
  64018=>"000101101",
  64019=>"111111010",
  64020=>"101100010",
  64021=>"110111100",
  64022=>"111100011",
  64023=>"000101010",
  64024=>"111110100",
  64025=>"000100000",
  64026=>"110001011",
  64027=>"111011110",
  64028=>"001000000",
  64029=>"011110011",
  64030=>"111110010",
  64031=>"011110011",
  64032=>"000010011",
  64033=>"000000111",
  64034=>"101111101",
  64035=>"000111000",
  64036=>"000110011",
  64037=>"100001110",
  64038=>"111111111",
  64039=>"011100011",
  64040=>"111111000",
  64041=>"100010110",
  64042=>"000100110",
  64043=>"110100000",
  64044=>"001001100",
  64045=>"011000011",
  64046=>"011010011",
  64047=>"111000101",
  64048=>"010010010",
  64049=>"010001101",
  64050=>"011101101",
  64051=>"000101111",
  64052=>"110001001",
  64053=>"000101101",
  64054=>"010010101",
  64055=>"101000000",
  64056=>"000111001",
  64057=>"101111011",
  64058=>"011010110",
  64059=>"110000111",
  64060=>"000110111",
  64061=>"111111100",
  64062=>"110010110",
  64063=>"000100000",
  64064=>"001010010",
  64065=>"100000011",
  64066=>"111110011",
  64067=>"010001100",
  64068=>"010111110",
  64069=>"011000100",
  64070=>"100100110",
  64071=>"111100011",
  64072=>"111111111",
  64073=>"001000101",
  64074=>"111011111",
  64075=>"010010011",
  64076=>"000001000",
  64077=>"100000001",
  64078=>"110111010",
  64079=>"001100010",
  64080=>"000011011",
  64081=>"100011001",
  64082=>"101010010",
  64083=>"001101100",
  64084=>"000100000",
  64085=>"101100001",
  64086=>"001001000",
  64087=>"000101001",
  64088=>"110111111",
  64089=>"111110001",
  64090=>"000100110",
  64091=>"111100111",
  64092=>"101001010",
  64093=>"000100010",
  64094=>"010100010",
  64095=>"000001010",
  64096=>"111001001",
  64097=>"000001010",
  64098=>"100011100",
  64099=>"001001001",
  64100=>"011101010",
  64101=>"000000010",
  64102=>"001010000",
  64103=>"111111111",
  64104=>"000111100",
  64105=>"010000100",
  64106=>"111111001",
  64107=>"110100000",
  64108=>"111101001",
  64109=>"101000111",
  64110=>"110011111",
  64111=>"100000001",
  64112=>"001100100",
  64113=>"111111111",
  64114=>"100000101",
  64115=>"101000010",
  64116=>"001011010",
  64117=>"101000001",
  64118=>"001000010",
  64119=>"011111001",
  64120=>"110100110",
  64121=>"100011010",
  64122=>"011001000",
  64123=>"011111100",
  64124=>"001100011",
  64125=>"111001111",
  64126=>"000100011",
  64127=>"110010100",
  64128=>"101101100",
  64129=>"011100000",
  64130=>"100001101",
  64131=>"111010000",
  64132=>"001001001",
  64133=>"011100100",
  64134=>"110010001",
  64135=>"100010001",
  64136=>"100110111",
  64137=>"110101001",
  64138=>"111001100",
  64139=>"000000000",
  64140=>"111111100",
  64141=>"110011001",
  64142=>"111000111",
  64143=>"110110101",
  64144=>"010000111",
  64145=>"010110000",
  64146=>"111111110",
  64147=>"111111001",
  64148=>"000110001",
  64149=>"010111001",
  64150=>"010011111",
  64151=>"010100101",
  64152=>"111110101",
  64153=>"100010111",
  64154=>"111101111",
  64155=>"010011100",
  64156=>"000001000",
  64157=>"001010100",
  64158=>"100011010",
  64159=>"101011011",
  64160=>"101001111",
  64161=>"100010011",
  64162=>"111110101",
  64163=>"111001100",
  64164=>"101101100",
  64165=>"000110010",
  64166=>"100111001",
  64167=>"101010110",
  64168=>"111111111",
  64169=>"100110001",
  64170=>"100000010",
  64171=>"001000000",
  64172=>"010010110",
  64173=>"010110011",
  64174=>"010001001",
  64175=>"010110101",
  64176=>"111110011",
  64177=>"011001001",
  64178=>"110111100",
  64179=>"110010010",
  64180=>"001001100",
  64181=>"100001011",
  64182=>"001010101",
  64183=>"100111011",
  64184=>"010100011",
  64185=>"110100000",
  64186=>"110101100",
  64187=>"010000000",
  64188=>"100100110",
  64189=>"010000000",
  64190=>"000010101",
  64191=>"011110100",
  64192=>"111100001",
  64193=>"010101111",
  64194=>"011110100",
  64195=>"111001101",
  64196=>"001111101",
  64197=>"011011011",
  64198=>"110110010",
  64199=>"000101110",
  64200=>"111011101",
  64201=>"001010001",
  64202=>"010000001",
  64203=>"011110110",
  64204=>"010001101",
  64205=>"100100000",
  64206=>"111001110",
  64207=>"001011111",
  64208=>"110001101",
  64209=>"101011101",
  64210=>"000101110",
  64211=>"001110011",
  64212=>"111111111",
  64213=>"010111011",
  64214=>"000100110",
  64215=>"001110001",
  64216=>"011110010",
  64217=>"111001101",
  64218=>"101101100",
  64219=>"001011001",
  64220=>"001011100",
  64221=>"100011000",
  64222=>"100101010",
  64223=>"110000000",
  64224=>"100110001",
  64225=>"001001100",
  64226=>"010001110",
  64227=>"110101101",
  64228=>"001010111",
  64229=>"101000010",
  64230=>"001010001",
  64231=>"000011010",
  64232=>"000000101",
  64233=>"111011101",
  64234=>"001000001",
  64235=>"101011010",
  64236=>"101100010",
  64237=>"000111110",
  64238=>"001101000",
  64239=>"000100011",
  64240=>"100010110",
  64241=>"000000110",
  64242=>"000111101",
  64243=>"011010011",
  64244=>"111101011",
  64245=>"001101100",
  64246=>"001100001",
  64247=>"111100000",
  64248=>"101001010",
  64249=>"011111001",
  64250=>"010011001",
  64251=>"111011100",
  64252=>"110001110",
  64253=>"001010011",
  64254=>"100011011",
  64255=>"010110010",
  64256=>"000010111",
  64257=>"110101001",
  64258=>"100000111",
  64259=>"011101100",
  64260=>"010011100",
  64261=>"111001110",
  64262=>"110111011",
  64263=>"101010000",
  64264=>"001110000",
  64265=>"010011111",
  64266=>"010001111",
  64267=>"011000110",
  64268=>"110110101",
  64269=>"011100101",
  64270=>"011100101",
  64271=>"100100010",
  64272=>"010000110",
  64273=>"100110010",
  64274=>"110000100",
  64275=>"100110010",
  64276=>"011110000",
  64277=>"111100111",
  64278=>"000111110",
  64279=>"110111110",
  64280=>"111011001",
  64281=>"100101111",
  64282=>"111000011",
  64283=>"110110011",
  64284=>"110110000",
  64285=>"010111011",
  64286=>"011010000",
  64287=>"101001100",
  64288=>"110010111",
  64289=>"010001000",
  64290=>"111110100",
  64291=>"001001011",
  64292=>"000110100",
  64293=>"101001110",
  64294=>"101011001",
  64295=>"111011000",
  64296=>"100001101",
  64297=>"101100010",
  64298=>"010010011",
  64299=>"000011101",
  64300=>"111101000",
  64301=>"100110111",
  64302=>"001000110",
  64303=>"010110101",
  64304=>"010010010",
  64305=>"001010000",
  64306=>"010001110",
  64307=>"101011101",
  64308=>"100100111",
  64309=>"000001011",
  64310=>"000001000",
  64311=>"000010111",
  64312=>"111111100",
  64313=>"101110001",
  64314=>"010111010",
  64315=>"100001001",
  64316=>"101110110",
  64317=>"000100100",
  64318=>"101010111",
  64319=>"010111101",
  64320=>"001001100",
  64321=>"111101010",
  64322=>"001100001",
  64323=>"001101000",
  64324=>"110110000",
  64325=>"101001100",
  64326=>"010111001",
  64327=>"000000001",
  64328=>"000100010",
  64329=>"011010111",
  64330=>"010001110",
  64331=>"011000101",
  64332=>"110011101",
  64333=>"100110000",
  64334=>"011001000",
  64335=>"010111100",
  64336=>"111011000",
  64337=>"001111101",
  64338=>"100001010",
  64339=>"110000100",
  64340=>"111010111",
  64341=>"011101100",
  64342=>"110011000",
  64343=>"000010110",
  64344=>"100000001",
  64345=>"000110100",
  64346=>"110100000",
  64347=>"000000110",
  64348=>"100100100",
  64349=>"000011111",
  64350=>"000000000",
  64351=>"100000000",
  64352=>"111011101",
  64353=>"110010000",
  64354=>"000100100",
  64355=>"111010010",
  64356=>"001100011",
  64357=>"101000111",
  64358=>"010001011",
  64359=>"101101011",
  64360=>"001010001",
  64361=>"101001010",
  64362=>"001001110",
  64363=>"100101110",
  64364=>"100000110",
  64365=>"011100100",
  64366=>"010110001",
  64367=>"101111001",
  64368=>"000100010",
  64369=>"010100101",
  64370=>"000000101",
  64371=>"100000100",
  64372=>"100011100",
  64373=>"101100000",
  64374=>"001100101",
  64375=>"001100101",
  64376=>"001101110",
  64377=>"000101101",
  64378=>"011010000",
  64379=>"001111101",
  64380=>"101100001",
  64381=>"111011101",
  64382=>"001101101",
  64383=>"100111110",
  64384=>"100011001",
  64385=>"101000010",
  64386=>"111101111",
  64387=>"000000110",
  64388=>"110111010",
  64389=>"111111001",
  64390=>"001111000",
  64391=>"111111000",
  64392=>"001011010",
  64393=>"101010001",
  64394=>"011011100",
  64395=>"011001011",
  64396=>"111010101",
  64397=>"000100111",
  64398=>"100010111",
  64399=>"110000011",
  64400=>"010011110",
  64401=>"111100011",
  64402=>"100100111",
  64403=>"110101000",
  64404=>"110000111",
  64405=>"101110100",
  64406=>"101000011",
  64407=>"001010010",
  64408=>"011001100",
  64409=>"111111111",
  64410=>"101001111",
  64411=>"000000000",
  64412=>"100010010",
  64413=>"101100101",
  64414=>"000011100",
  64415=>"001011001",
  64416=>"101100110",
  64417=>"001110010",
  64418=>"011011011",
  64419=>"001011101",
  64420=>"101000001",
  64421=>"001110011",
  64422=>"110000000",
  64423=>"001101100",
  64424=>"110101001",
  64425=>"101001010",
  64426=>"111011111",
  64427=>"111101111",
  64428=>"001010111",
  64429=>"010000010",
  64430=>"100011000",
  64431=>"101100001",
  64432=>"011111001",
  64433=>"100001110",
  64434=>"001001011",
  64435=>"000001001",
  64436=>"100111001",
  64437=>"110111101",
  64438=>"010001010",
  64439=>"011011001",
  64440=>"111101000",
  64441=>"001010011",
  64442=>"000100010",
  64443=>"010001001",
  64444=>"001110110",
  64445=>"100000100",
  64446=>"111111100",
  64447=>"000010001",
  64448=>"000101110",
  64449=>"000110100",
  64450=>"100010010",
  64451=>"101111111",
  64452=>"110100011",
  64453=>"010010101",
  64454=>"111100110",
  64455=>"011101011",
  64456=>"010001011",
  64457=>"101101111",
  64458=>"001011011",
  64459=>"101010111",
  64460=>"100000111",
  64461=>"001000011",
  64462=>"101111000",
  64463=>"110011001",
  64464=>"111001111",
  64465=>"100100111",
  64466=>"011101110",
  64467=>"001111111",
  64468=>"010111001",
  64469=>"111001011",
  64470=>"101011000",
  64471=>"101110001",
  64472=>"100011110",
  64473=>"011010111",
  64474=>"111011100",
  64475=>"100001010",
  64476=>"101101011",
  64477=>"000110000",
  64478=>"100111001",
  64479=>"110101110",
  64480=>"001111100",
  64481=>"011000110",
  64482=>"000001100",
  64483=>"001100001",
  64484=>"110111110",
  64485=>"000001000",
  64486=>"011001011",
  64487=>"011000001",
  64488=>"001011110",
  64489=>"000110101",
  64490=>"001111100",
  64491=>"111110001",
  64492=>"011001110",
  64493=>"000101001",
  64494=>"011011111",
  64495=>"001000111",
  64496=>"000101000",
  64497=>"110110110",
  64498=>"010101001",
  64499=>"010000001",
  64500=>"001001000",
  64501=>"100000100",
  64502=>"111001100",
  64503=>"111100111",
  64504=>"100110010",
  64505=>"100000100",
  64506=>"010011111",
  64507=>"100010110",
  64508=>"110010110",
  64509=>"101001011",
  64510=>"110011100",
  64511=>"011101110",
  64512=>"011100001",
  64513=>"101010011",
  64514=>"111000111",
  64515=>"100111100",
  64516=>"010101001",
  64517=>"110000110",
  64518=>"001000001",
  64519=>"010001111",
  64520=>"110111110",
  64521=>"111100100",
  64522=>"100110111",
  64523=>"010101101",
  64524=>"000000100",
  64525=>"010010011",
  64526=>"111101101",
  64527=>"000000010",
  64528=>"111001111",
  64529=>"110011011",
  64530=>"110111010",
  64531=>"001101001",
  64532=>"000010101",
  64533=>"001101000",
  64534=>"001111011",
  64535=>"000000110",
  64536=>"111111001",
  64537=>"000100000",
  64538=>"100110010",
  64539=>"101100011",
  64540=>"100111010",
  64541=>"100001111",
  64542=>"101011111",
  64543=>"000111010",
  64544=>"010010100",
  64545=>"010010110",
  64546=>"000010110",
  64547=>"010011111",
  64548=>"111101000",
  64549=>"100011011",
  64550=>"100110100",
  64551=>"110010011",
  64552=>"011101110",
  64553=>"010101000",
  64554=>"001011100",
  64555=>"011111000",
  64556=>"100010001",
  64557=>"010110100",
  64558=>"110110110",
  64559=>"011111010",
  64560=>"101100100",
  64561=>"000001000",
  64562=>"110101000",
  64563=>"001001010",
  64564=>"000100110",
  64565=>"101001011",
  64566=>"111010100",
  64567=>"011000010",
  64568=>"101100000",
  64569=>"110110110",
  64570=>"100100000",
  64571=>"100101100",
  64572=>"011000000",
  64573=>"101100111",
  64574=>"010001000",
  64575=>"000001010",
  64576=>"000111101",
  64577=>"101100111",
  64578=>"110101100",
  64579=>"011100101",
  64580=>"100100111",
  64581=>"110100010",
  64582=>"111101111",
  64583=>"110101001",
  64584=>"110001001",
  64585=>"101100100",
  64586=>"110111010",
  64587=>"010001110",
  64588=>"000010111",
  64589=>"001001001",
  64590=>"111100110",
  64591=>"101110111",
  64592=>"010010101",
  64593=>"110011100",
  64594=>"101011001",
  64595=>"001000010",
  64596=>"110101001",
  64597=>"010010101",
  64598=>"100010110",
  64599=>"001010100",
  64600=>"001010110",
  64601=>"100100110",
  64602=>"111110010",
  64603=>"010011100",
  64604=>"010001101",
  64605=>"001100110",
  64606=>"100101011",
  64607=>"011011011",
  64608=>"001010111",
  64609=>"111101110",
  64610=>"000000110",
  64611=>"001000000",
  64612=>"011110001",
  64613=>"000011110",
  64614=>"011100100",
  64615=>"100000000",
  64616=>"011111011",
  64617=>"011001101",
  64618=>"001110111",
  64619=>"111110001",
  64620=>"011111011",
  64621=>"011111010",
  64622=>"110110000",
  64623=>"000010101",
  64624=>"011011011",
  64625=>"000001000",
  64626=>"000010110",
  64627=>"010001101",
  64628=>"010010001",
  64629=>"010111011",
  64630=>"000010010",
  64631=>"111100000",
  64632=>"100110100",
  64633=>"111101000",
  64634=>"000001111",
  64635=>"000111011",
  64636=>"000000010",
  64637=>"111011001",
  64638=>"001001000",
  64639=>"111011100",
  64640=>"101001101",
  64641=>"000000011",
  64642=>"101101111",
  64643=>"101100100",
  64644=>"100010010",
  64645=>"111110111",
  64646=>"001000101",
  64647=>"110000011",
  64648=>"101101110",
  64649=>"101010001",
  64650=>"111110011",
  64651=>"000010100",
  64652=>"010111100",
  64653=>"001100101",
  64654=>"101110101",
  64655=>"111100011",
  64656=>"110010000",
  64657=>"111110110",
  64658=>"100110110",
  64659=>"010001000",
  64660=>"111110101",
  64661=>"110110010",
  64662=>"011110010",
  64663=>"101010110",
  64664=>"000010011",
  64665=>"111100110",
  64666=>"001110000",
  64667=>"001010011",
  64668=>"101101001",
  64669=>"011011111",
  64670=>"110100101",
  64671=>"111101010",
  64672=>"110000011",
  64673=>"100110100",
  64674=>"001010100",
  64675=>"100101110",
  64676=>"110110110",
  64677=>"001001100",
  64678=>"000010001",
  64679=>"001101111",
  64680=>"011000011",
  64681=>"010111110",
  64682=>"101010001",
  64683=>"110100100",
  64684=>"011110011",
  64685=>"101001100",
  64686=>"000000110",
  64687=>"111100000",
  64688=>"101100000",
  64689=>"111110010",
  64690=>"000010010",
  64691=>"110111101",
  64692=>"110000111",
  64693=>"010000110",
  64694=>"011111110",
  64695=>"011010011",
  64696=>"111010001",
  64697=>"110100101",
  64698=>"010100000",
  64699=>"110101111",
  64700=>"110101000",
  64701=>"010000110",
  64702=>"010011011",
  64703=>"110011010",
  64704=>"010000110",
  64705=>"101111010",
  64706=>"000111011",
  64707=>"000000011",
  64708=>"100011110",
  64709=>"011101100",
  64710=>"000010101",
  64711=>"011111011",
  64712=>"011001111",
  64713=>"111000101",
  64714=>"100101101",
  64715=>"001010111",
  64716=>"111010110",
  64717=>"100101101",
  64718=>"000011000",
  64719=>"101110011",
  64720=>"011110001",
  64721=>"101110100",
  64722=>"000110001",
  64723=>"100110100",
  64724=>"100000110",
  64725=>"011000011",
  64726=>"100001111",
  64727=>"000011101",
  64728=>"000101100",
  64729=>"110100010",
  64730=>"010111101",
  64731=>"010101000",
  64732=>"011000001",
  64733=>"111011001",
  64734=>"110111000",
  64735=>"010011100",
  64736=>"001000001",
  64737=>"000000000",
  64738=>"010111101",
  64739=>"100001100",
  64740=>"010100110",
  64741=>"110100110",
  64742=>"100000100",
  64743=>"000100100",
  64744=>"000010110",
  64745=>"001011001",
  64746=>"110000011",
  64747=>"000111101",
  64748=>"111101101",
  64749=>"011001001",
  64750=>"100011001",
  64751=>"100111011",
  64752=>"010001000",
  64753=>"111100101",
  64754=>"110010010",
  64755=>"111000100",
  64756=>"101100110",
  64757=>"111100110",
  64758=>"000000110",
  64759=>"111110010",
  64760=>"101110010",
  64761=>"101111011",
  64762=>"110101111",
  64763=>"101110101",
  64764=>"000001011",
  64765=>"000110010",
  64766=>"011001101",
  64767=>"110101010",
  64768=>"110100011",
  64769=>"001001010",
  64770=>"000100000",
  64771=>"010000011",
  64772=>"001001110",
  64773=>"101110111",
  64774=>"000000000",
  64775=>"110010001",
  64776=>"001110111",
  64777=>"011011001",
  64778=>"100111111",
  64779=>"000100001",
  64780=>"000000011",
  64781=>"101110010",
  64782=>"111111110",
  64783=>"000000001",
  64784=>"110000000",
  64785=>"100100011",
  64786=>"111010010",
  64787=>"110001110",
  64788=>"000110000",
  64789=>"000000110",
  64790=>"000101100",
  64791=>"001010110",
  64792=>"111010111",
  64793=>"100011001",
  64794=>"010001110",
  64795=>"111000011",
  64796=>"001000011",
  64797=>"010010010",
  64798=>"110001011",
  64799=>"100011010",
  64800=>"001111001",
  64801=>"001000111",
  64802=>"010100000",
  64803=>"000101001",
  64804=>"011110101",
  64805=>"111100111",
  64806=>"101110110",
  64807=>"001000001",
  64808=>"001011101",
  64809=>"111100111",
  64810=>"100101001",
  64811=>"110001000",
  64812=>"101001011",
  64813=>"000111011",
  64814=>"100101010",
  64815=>"101011111",
  64816=>"010001001",
  64817=>"011001000",
  64818=>"001101010",
  64819=>"101011110",
  64820=>"100011111",
  64821=>"100100111",
  64822=>"010111001",
  64823=>"101110101",
  64824=>"011001000",
  64825=>"111101111",
  64826=>"101001110",
  64827=>"100100010",
  64828=>"100100110",
  64829=>"101001000",
  64830=>"101110010",
  64831=>"111100100",
  64832=>"100010101",
  64833=>"010000010",
  64834=>"111110101",
  64835=>"101000001",
  64836=>"111001001",
  64837=>"111101100",
  64838=>"110000001",
  64839=>"111100001",
  64840=>"010110100",
  64841=>"011000011",
  64842=>"100001010",
  64843=>"000000001",
  64844=>"111111001",
  64845=>"001000110",
  64846=>"100110110",
  64847=>"101111111",
  64848=>"011010011",
  64849=>"111101110",
  64850=>"000101000",
  64851=>"010100001",
  64852=>"111000000",
  64853=>"110001001",
  64854=>"101001000",
  64855=>"011100010",
  64856=>"000100010",
  64857=>"000100101",
  64858=>"000111110",
  64859=>"011000101",
  64860=>"011100100",
  64861=>"110001110",
  64862=>"111011000",
  64863=>"111110001",
  64864=>"001110101",
  64865=>"111100011",
  64866=>"111101000",
  64867=>"000000000",
  64868=>"100001101",
  64869=>"110100001",
  64870=>"010100001",
  64871=>"011100111",
  64872=>"001000111",
  64873=>"001011011",
  64874=>"011000000",
  64875=>"000100110",
  64876=>"001100101",
  64877=>"101010110",
  64878=>"101001000",
  64879=>"011011000",
  64880=>"100100010",
  64881=>"110100111",
  64882=>"111001101",
  64883=>"110111100",
  64884=>"101111011",
  64885=>"011001001",
  64886=>"110100111",
  64887=>"111100100",
  64888=>"001010100",
  64889=>"101000100",
  64890=>"100010001",
  64891=>"011110110",
  64892=>"110100110",
  64893=>"100000011",
  64894=>"010101011",
  64895=>"101101101",
  64896=>"111110010",
  64897=>"011001010",
  64898=>"000001111",
  64899=>"000001010",
  64900=>"001011001",
  64901=>"010010011",
  64902=>"011101111",
  64903=>"110011100",
  64904=>"110001000",
  64905=>"000000000",
  64906=>"101011110",
  64907=>"010001110",
  64908=>"111010000",
  64909=>"101011000",
  64910=>"110011100",
  64911=>"110111111",
  64912=>"001110001",
  64913=>"101101101",
  64914=>"100111110",
  64915=>"111011001",
  64916=>"001010010",
  64917=>"110100100",
  64918=>"101110100",
  64919=>"110011101",
  64920=>"001011101",
  64921=>"100110100",
  64922=>"001010100",
  64923=>"100000000",
  64924=>"111100101",
  64925=>"000101000",
  64926=>"101011101",
  64927=>"001100111",
  64928=>"100110110",
  64929=>"111011101",
  64930=>"011100000",
  64931=>"100100000",
  64932=>"111101101",
  64933=>"011011001",
  64934=>"000000110",
  64935=>"011000011",
  64936=>"001111100",
  64937=>"001000000",
  64938=>"100111100",
  64939=>"010110010",
  64940=>"000010010",
  64941=>"101111110",
  64942=>"100110000",
  64943=>"101100011",
  64944=>"110100000",
  64945=>"010011100",
  64946=>"101001111",
  64947=>"100110010",
  64948=>"111010101",
  64949=>"000001001",
  64950=>"001111011",
  64951=>"110010100",
  64952=>"111011110",
  64953=>"010010110",
  64954=>"001011001",
  64955=>"001110111",
  64956=>"111011010",
  64957=>"110111100",
  64958=>"001111000",
  64959=>"110000100",
  64960=>"000110011",
  64961=>"100011110",
  64962=>"001111110",
  64963=>"010111010",
  64964=>"110010010",
  64965=>"011001011",
  64966=>"010011101",
  64967=>"111001000",
  64968=>"001101111",
  64969=>"110000101",
  64970=>"100101001",
  64971=>"100110111",
  64972=>"010000010",
  64973=>"111110100",
  64974=>"000000000",
  64975=>"100011110",
  64976=>"100001100",
  64977=>"000000000",
  64978=>"011101111",
  64979=>"010100111",
  64980=>"101011101",
  64981=>"111001010",
  64982=>"001110101",
  64983=>"100011010",
  64984=>"010000010",
  64985=>"111110101",
  64986=>"010110000",
  64987=>"111011111",
  64988=>"111011000",
  64989=>"011001100",
  64990=>"101000100",
  64991=>"011011010",
  64992=>"000100100",
  64993=>"110111011",
  64994=>"111101110",
  64995=>"011111101",
  64996=>"011101100",
  64997=>"110111000",
  64998=>"001010001",
  64999=>"100000101",
  65000=>"001111000",
  65001=>"000001111",
  65002=>"010000001",
  65003=>"001011111",
  65004=>"111111100",
  65005=>"100010011",
  65006=>"101000010",
  65007=>"011101011",
  65008=>"001101010",
  65009=>"011101111",
  65010=>"100100100",
  65011=>"110111001",
  65012=>"010110001",
  65013=>"001011010",
  65014=>"000001001",
  65015=>"100100000",
  65016=>"111001000",
  65017=>"011011010",
  65018=>"001101011",
  65019=>"001110011",
  65020=>"001110100",
  65021=>"110000100",
  65022=>"110011100",
  65023=>"110011011",
  65024=>"011001101",
  65025=>"101110000",
  65026=>"101101011",
  65027=>"111010000",
  65028=>"101101111",
  65029=>"111011000",
  65030=>"010001111",
  65031=>"111000010",
  65032=>"100011010",
  65033=>"000110110",
  65034=>"001100111",
  65035=>"111011001",
  65036=>"011110001",
  65037=>"001000001",
  65038=>"111110010",
  65039=>"001110000",
  65040=>"100100011",
  65041=>"110101001",
  65042=>"001011000",
  65043=>"111111110",
  65044=>"010000011",
  65045=>"000111010",
  65046=>"011101010",
  65047=>"110111001",
  65048=>"000001000",
  65049=>"010011010",
  65050=>"011011111",
  65051=>"011001110",
  65052=>"100101111",
  65053=>"100110100",
  65054=>"100011111",
  65055=>"110001100",
  65056=>"000010010",
  65057=>"111101000",
  65058=>"000001100",
  65059=>"110000100",
  65060=>"010111101",
  65061=>"100101111",
  65062=>"110000010",
  65063=>"101010001",
  65064=>"000111010",
  65065=>"110101101",
  65066=>"111010101",
  65067=>"001110001",
  65068=>"111010001",
  65069=>"100110101",
  65070=>"010011010",
  65071=>"011011110",
  65072=>"011110100",
  65073=>"110101111",
  65074=>"111101111",
  65075=>"001111000",
  65076=>"101011111",
  65077=>"110000000",
  65078=>"110111010",
  65079=>"001011001",
  65080=>"100110010",
  65081=>"110011001",
  65082=>"100000110",
  65083=>"111011110",
  65084=>"000111010",
  65085=>"001111010",
  65086=>"111101001",
  65087=>"101011111",
  65088=>"111111111",
  65089=>"111010000",
  65090=>"101101011",
  65091=>"001110010",
  65092=>"110000001",
  65093=>"001100101",
  65094=>"100010100",
  65095=>"011010010",
  65096=>"011100100",
  65097=>"010010111",
  65098=>"010111010",
  65099=>"000110100",
  65100=>"000110111",
  65101=>"000000011",
  65102=>"001111101",
  65103=>"011101000",
  65104=>"000111010",
  65105=>"000011111",
  65106=>"100011000",
  65107=>"000110110",
  65108=>"000110101",
  65109=>"011001000",
  65110=>"011000000",
  65111=>"111100111",
  65112=>"111011010",
  65113=>"001100010",
  65114=>"011110111",
  65115=>"110111011",
  65116=>"000011000",
  65117=>"001011111",
  65118=>"000111101",
  65119=>"111010111",
  65120=>"101011000",
  65121=>"101001011",
  65122=>"010101010",
  65123=>"000000001",
  65124=>"111111100",
  65125=>"110110110",
  65126=>"000111001",
  65127=>"100110010",
  65128=>"000000100",
  65129=>"111000001",
  65130=>"001000011",
  65131=>"101100111",
  65132=>"100101100",
  65133=>"111100000",
  65134=>"010000110",
  65135=>"010011011",
  65136=>"001000110",
  65137=>"001011011",
  65138=>"011110011",
  65139=>"111110100",
  65140=>"100001010",
  65141=>"111001000",
  65142=>"110111011",
  65143=>"110111001",
  65144=>"101100111",
  65145=>"011100111",
  65146=>"101000001",
  65147=>"100110111",
  65148=>"100000001",
  65149=>"011101110",
  65150=>"110110110",
  65151=>"001100010",
  65152=>"001100101",
  65153=>"010000010",
  65154=>"101100100",
  65155=>"000101001",
  65156=>"100001100",
  65157=>"110001000",
  65158=>"001100101",
  65159=>"110111111",
  65160=>"000001100",
  65161=>"101001100",
  65162=>"001011111",
  65163=>"100010101",
  65164=>"110000101",
  65165=>"111011110",
  65166=>"110111000",
  65167=>"101110111",
  65168=>"010010101",
  65169=>"100010111",
  65170=>"010111011",
  65171=>"001010011",
  65172=>"000000110",
  65173=>"001001011",
  65174=>"110001000",
  65175=>"000011001",
  65176=>"111001011",
  65177=>"010100011",
  65178=>"001010110",
  65179=>"100101100",
  65180=>"111010100",
  65181=>"011110101",
  65182=>"101000010",
  65183=>"111000001",
  65184=>"110110101",
  65185=>"110110011",
  65186=>"101001001",
  65187=>"001000111",
  65188=>"110100000",
  65189=>"000000111",
  65190=>"111100010",
  65191=>"000001110",
  65192=>"110000001",
  65193=>"001010000",
  65194=>"101101111",
  65195=>"101101110",
  65196=>"110001100",
  65197=>"010100001",
  65198=>"111111001",
  65199=>"011011111",
  65200=>"010000100",
  65201=>"001011110",
  65202=>"101101000",
  65203=>"110101010",
  65204=>"011101011",
  65205=>"110100001",
  65206=>"000010010",
  65207=>"010001100",
  65208=>"101000010",
  65209=>"101001011",
  65210=>"000110011",
  65211=>"101101101",
  65212=>"111010100",
  65213=>"010101000",
  65214=>"100011011",
  65215=>"100101100",
  65216=>"100011000",
  65217=>"010110100",
  65218=>"100000111",
  65219=>"010100010",
  65220=>"001011000",
  65221=>"110100000",
  65222=>"111100100",
  65223=>"001001110",
  65224=>"101111110",
  65225=>"010101010",
  65226=>"010011100",
  65227=>"101100011",
  65228=>"010010110",
  65229=>"110101011",
  65230=>"101011010",
  65231=>"001111011",
  65232=>"000110011",
  65233=>"111111000",
  65234=>"000000001",
  65235=>"111100100",
  65236=>"001101011",
  65237=>"101000000",
  65238=>"011000011",
  65239=>"010010010",
  65240=>"000000001",
  65241=>"000111010",
  65242=>"111100000",
  65243=>"111101111",
  65244=>"011001000",
  65245=>"110011101",
  65246=>"000000111",
  65247=>"010000101",
  65248=>"101001000",
  65249=>"011101101",
  65250=>"111000001",
  65251=>"001100101",
  65252=>"101100000",
  65253=>"111101111",
  65254=>"101111001",
  65255=>"100101000",
  65256=>"000100011",
  65257=>"101011100",
  65258=>"010010111",
  65259=>"001010100",
  65260=>"011011101",
  65261=>"000010100",
  65262=>"010100111",
  65263=>"000001011",
  65264=>"000010111",
  65265=>"000101101",
  65266=>"101101010",
  65267=>"111001000",
  65268=>"110011101",
  65269=>"010000100",
  65270=>"000101111",
  65271=>"000111111",
  65272=>"101011000",
  65273=>"101010000",
  65274=>"010010010",
  65275=>"111001101",
  65276=>"011011010",
  65277=>"111110110",
  65278=>"001110010",
  65279=>"111001110",
  65280=>"111001101",
  65281=>"101101011",
  65282=>"110011011",
  65283=>"111100111",
  65284=>"111001101",
  65285=>"010010001",
  65286=>"101111010",
  65287=>"111000101",
  65288=>"011001100",
  65289=>"100101101",
  65290=>"000001001",
  65291=>"100001000",
  65292=>"101011110",
  65293=>"000101001",
  65294=>"010000011",
  65295=>"010110000",
  65296=>"001001001",
  65297=>"000011010",
  65298=>"001111100",
  65299=>"001001110",
  65300=>"101100001",
  65301=>"111011110",
  65302=>"011011110",
  65303=>"111011100",
  65304=>"011010010",
  65305=>"110011110",
  65306=>"000111010",
  65307=>"011001000",
  65308=>"111111101",
  65309=>"111011100",
  65310=>"110100110",
  65311=>"000000111",
  65312=>"110111011",
  65313=>"111000001",
  65314=>"111110100",
  65315=>"101101101",
  65316=>"100000011",
  65317=>"101110000",
  65318=>"001000011",
  65319=>"110011110",
  65320=>"011100110",
  65321=>"011011011",
  65322=>"011111000",
  65323=>"000010011",
  65324=>"000100100",
  65325=>"001011011",
  65326=>"110110001",
  65327=>"000110011",
  65328=>"000010001",
  65329=>"001010011",
  65330=>"001100001",
  65331=>"111101101",
  65332=>"011101101",
  65333=>"111001110",
  65334=>"111110010",
  65335=>"101000001",
  65336=>"011100101",
  65337=>"101011110",
  65338=>"111110001",
  65339=>"111011011",
  65340=>"101001001",
  65341=>"111101101",
  65342=>"111001010",
  65343=>"110001010",
  65344=>"000010111",
  65345=>"111000111",
  65346=>"111100001",
  65347=>"011011011",
  65348=>"111100111",
  65349=>"010101000",
  65350=>"111111011",
  65351=>"000110111",
  65352=>"100111110",
  65353=>"101110011",
  65354=>"010101110",
  65355=>"001000111",
  65356=>"000110010",
  65357=>"001111001",
  65358=>"111000100",
  65359=>"010111010",
  65360=>"110100001",
  65361=>"000001101",
  65362=>"110011001",
  65363=>"111001011",
  65364=>"101010111",
  65365=>"001110101",
  65366=>"100001101",
  65367=>"011100110",
  65368=>"100000100",
  65369=>"000110100",
  65370=>"101110011",
  65371=>"000101001",
  65372=>"100000100",
  65373=>"101111101",
  65374=>"100011101",
  65375=>"001001000",
  65376=>"110111100",
  65377=>"110001000",
  65378=>"000101011",
  65379=>"001011110",
  65380=>"010001000",
  65381=>"111110000",
  65382=>"010000010",
  65383=>"111110010",
  65384=>"011011011",
  65385=>"000110110",
  65386=>"011000000",
  65387=>"000100000",
  65388=>"011110111",
  65389=>"110011000",
  65390=>"110101011",
  65391=>"010010000",
  65392=>"011010100",
  65393=>"001110010",
  65394=>"100111010",
  65395=>"010000000",
  65396=>"110000110",
  65397=>"100001010",
  65398=>"101001011",
  65399=>"110100100",
  65400=>"101100101",
  65401=>"100100111",
  65402=>"001010101",
  65403=>"111110000",
  65404=>"000000000",
  65405=>"100100010",
  65406=>"000110110",
  65407=>"010010011",
  65408=>"001110111",
  65409=>"010011010",
  65410=>"110010011",
  65411=>"100111101",
  65412=>"110101101",
  65413=>"010010111",
  65414=>"101011110",
  65415=>"010110100",
  65416=>"111011101",
  65417=>"001011101",
  65418=>"101010110",
  65419=>"110101000",
  65420=>"111001111",
  65421=>"101001101",
  65422=>"101100101",
  65423=>"101101011",
  65424=>"100011100",
  65425=>"101011101",
  65426=>"100001000",
  65427=>"111100001",
  65428=>"000011000",
  65429=>"011101111",
  65430=>"110110010",
  65431=>"011011001",
  65432=>"010010111",
  65433=>"110101110",
  65434=>"010010000",
  65435=>"100001111",
  65436=>"010100111",
  65437=>"010101001",
  65438=>"011000111",
  65439=>"011010101",
  65440=>"111101101",
  65441=>"101111111",
  65442=>"101010001",
  65443=>"001001001",
  65444=>"000010001",
  65445=>"011010100",
  65446=>"100111110",
  65447=>"011111101",
  65448=>"110111011",
  65449=>"011100010",
  65450=>"100001101",
  65451=>"001110010",
  65452=>"010101111",
  65453=>"000111101",
  65454=>"010100001",
  65455=>"101101111",
  65456=>"010011101",
  65457=>"111110111",
  65458=>"111110100",
  65459=>"110001001",
  65460=>"101010100",
  65461=>"011111000",
  65462=>"010110001",
  65463=>"011101011",
  65464=>"001111010",
  65465=>"011001111",
  65466=>"001100011",
  65467=>"010101111",
  65468=>"001011010",
  65469=>"011110100",
  65470=>"101011111",
  65471=>"101101010",
  65472=>"000011001",
  65473=>"011100011",
  65474=>"000100111",
  65475=>"111100101",
  65476=>"001000111",
  65477=>"100000101",
  65478=>"010100100",
  65479=>"110001000",
  65480=>"011010101",
  65481=>"110000000",
  65482=>"110100011",
  65483=>"111001101",
  65484=>"011111111",
  65485=>"101000110",
  65486=>"100101000",
  65487=>"000100101",
  65488=>"000110100",
  65489=>"111111101",
  65490=>"100110000",
  65491=>"000100000",
  65492=>"001000000",
  65493=>"000010010",
  65494=>"011101000",
  65495=>"000001100",
  65496=>"001011101",
  65497=>"000100000",
  65498=>"000101000",
  65499=>"000111011",
  65500=>"111101010",
  65501=>"001111010",
  65502=>"000001011",
  65503=>"011110000",
  65504=>"000001011",
  65505=>"000001110",
  65506=>"011101011",
  65507=>"101000111",
  65508=>"111001100",
  65509=>"111101001",
  65510=>"100001000",
  65511=>"111001001",
  65512=>"010001000",
  65513=>"000001011",
  65514=>"110011111",
  65515=>"000011010",
  65516=>"000011100",
  65517=>"111101101",
  65518=>"000011000",
  65519=>"011101000",
  65520=>"000011000",
  65521=>"110101101",
  65522=>"010101011",
  65523=>"100101010",
  65524=>"111010101",
  65525=>"010001001",
  65526=>"001011000",
  65527=>"001000000",
  65528=>"101011001",
  65529=>"000111000",
  65530=>"011010001",
  65531=>"110110001",
  65532=>"111100000",
  65533=>"010101111",
  65534=>"010101101",
  65535=>"000111100");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;