LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L5_1_WROM IS
    PORT (
        weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
        address : IN unsigned(weightsbitsAddress(5)-1 DOWNTO 0));
END L5_1_WROM;

ARCHITECTURE RTL OF L5_1_WROM IS

    TYPE ROM_mem IS ARRAY (0 TO 16383) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem := (0=>"000110111",
    1=>"011001100",
    2=>"011001000",
    3=>"000010011",
    4=>"010011001",
    5=>"010000100",
    6=>"000000111",
    7=>"001100000",
    8=>"110011111",
    9=>"000111000",
    10=>"010001001",
    11=>"110011000",
    12=>"000100110",
    13=>"010111111",
    14=>"000000111",
    15=>"001100110",
    16=>"010110000",
    17=>"011011010",
    18=>"110011001",
    19=>"000100101",
    20=>"000110110",
    21=>"011001000",
    22=>"110000110",
    23=>"100100110",
    24=>"010011001",
    25=>"101100000",
    26=>"010011101",
    27=>"110111111",
    28=>"000000000",
    29=>"010011101",
    30=>"010011001",
    31=>"100001001",
    32=>"010111001",
    33=>"100010001",
    34=>"111011001",
    35=>"010011011",
    36=>"110010111",
    37=>"010001000",
    38=>"000100110",
    39=>"010111111",
    40=>"110011001",
    41=>"000100101",
    42=>"001000001",
    43=>"110001001",
    44=>"110011100",
    45=>"010111011",
    46=>"110001000",
    47=>"110011000",
    48=>"110010111",
    49=>"001100000",
    50=>"110000000",
    51=>"100110111",
    52=>"110011111",
    53=>"100100011",
    54=>"110111100",
    55=>"011011010",
    56=>"100001101",
    57=>"110011001",
    58=>"110001001",
    59=>"001000010",
    60=>"101000000",
    61=>"100000000",
    62=>"000100000",
    63=>"110111101",
    64=>"011001001",
    65=>"101100111",
    66=>"110110000",
    67=>"100110111",
    68=>"010111100",
    69=>"100010011",
    70=>"100010010",
    71=>"100000110",
    72=>"100100110",
    73=>"000000111",
    74=>"110011000",
    75=>"000100100",
    76=>"100110000",
    77=>"110001000",
    78=>"110100110",
    79=>"001100110",
    80=>"100110110",
    81=>"001100110",
    82=>"000000000",
    83=>"000000011",
    84=>"100111110",
    85=>"001100010",
    86=>"000110010",
    87=>"000011011",
    88=>"010001101",
    89=>"010001111",
    90=>"110000111",
    91=>"000000110",
    92=>"010010011",
    93=>"110011001",
    94=>"010001111",
    95=>"001000000",
    96=>"010111111",
    97=>"100110110",
    98=>"101110111",
    99=>"110011100",
    100=>"110011000",
    101=>"000110011",
    102=>"000100010",
    103=>"010010100",
    104=>"000110110",
    105=>"001000000",
    106=>"010001001",
    107=>"000101111",
    108=>"000100010",
    109=>"000100110",
    110=>"010111011",
    111=>"010011001",
    112=>"110110000",
    113=>"000000100",
    114=>"000110110",
    115=>"010110100",
    116=>"011001100",
    117=>"001000110",
    118=>"001101111",
    119=>"100110110",
    120=>"110011111",
    121=>"101000101",
    122=>"001100100",
    123=>"111101100",
    124=>"001000100",
    125=>"111001000",
    126=>"110101000",
    127=>"101000111",
    128=>"000101101",
    129=>"000000001",
    130=>"000001111",
    131=>"010001010",
    132=>"000011011",
    133=>"010111110",
    134=>"000101101",
    135=>"111000000",
    136=>"111011011",
    137=>"000000000",
    138=>"000000110",
    139=>"001100010",
    140=>"010110101",
    141=>"110111100",
    142=>"101100000",
    143=>"110100100",
    144=>"110011000",
    145=>"110110111",
    146=>"000000000",
    147=>"110111110",
    148=>"101001101",
    149=>"010010000",
    150=>"000000000",
    151=>"110000000",
    152=>"000110100",
    153=>"100000010",
    154=>"000010011",
    155=>"111001000",
    156=>"101001001",
    157=>"000010110",
    158=>"011011011",
    159=>"101000010",
    160=>"100010111",
    161=>"111111111",
    162=>"001000110",
    163=>"010111101",
    164=>"111101000",
    165=>"001111001",
    166=>"111011000",
    167=>"001101111",
    168=>"001111111",
    169=>"111110100",
    170=>"000011101",
    171=>"001110110",
    172=>"010011001",
    173=>"111000000",
    174=>"111111001",
    175=>"110000000",
    176=>"001001000",
    177=>"000001111",
    178=>"100111001",
    179=>"001100100",
    180=>"001000010",
    181=>"011000010",
    182=>"000000010",
    183=>"111001010",
    184=>"000000000",
    185=>"010111111",
    186=>"001000000",
    187=>"101000011",
    188=>"001000000",
    189=>"010100101",
    190=>"111100000",
    191=>"000011001",
    192=>"000010110",
    193=>"000000000",
    194=>"110000000",
    195=>"001000000",
    196=>"111111001",
    197=>"000100101",
    198=>"111001000",
    199=>"000110000",
    200=>"110110100",
    201=>"000000110",
    202=>"000011011",
    203=>"000000010",
    204=>"111000001",
    205=>"000111011",
    206=>"111000000",
    207=>"101000011",
    208=>"000000010",
    209=>"100100001",
    210=>"001011000",
    211=>"001111011",
    212=>"110001101",
    213=>"001000000",
    214=>"001001000",
    215=>"011000000",
    216=>"110000001",
    217=>"111101000",
    218=>"010111110",
    219=>"111000111",
    220=>"000010111",
    221=>"111011001",
    222=>"000110110",
    223=>"010010010",
    224=>"100100100",
    225=>"100100001",
    226=>"101000111",
    227=>"100000011",
    228=>"111111000",
    229=>"111000001",
    230=>"011001100",
    231=>"011111000",
    232=>"111111000",
    233=>"000000011",
    234=>"000111111",
    235=>"111101000",
    236=>"000000000",
    237=>"111010010",
    238=>"001010111",
    239=>"111101100",
    240=>"111000000",
    241=>"100111111",
    242=>"100101011",
    243=>"001011111",
    244=>"000000111",
    245=>"101000101",
    246=>"101111100",
    247=>"001111110",
    248=>"001011000",
    249=>"000111111",
    250=>"111100100",
    251=>"100011110",
    252=>"010111011",
    253=>"111000000",
    254=>"010010010",
    255=>"000000110",
    256=>"110111110",
    257=>"000000000",
    258=>"111111111",
    259=>"111111111",
    260=>"000000000",
    261=>"001101000",
    262=>"001010111",
    263=>"000000000",
    264=>"000100100",
    265=>"000000000",
    266=>"111111111",
    267=>"111011111",
    268=>"111010101",
    269=>"111111100",
    270=>"000100000",
    271=>"001000100",
    272=>"111001101",
    273=>"100100000",
    274=>"000000000",
    275=>"000000000",
    276=>"000000000",
    277=>"110100010",
    278=>"000000000",
    279=>"000000000",
    280=>"000000000",
    281=>"011110101",
    282=>"000000000",
    283=>"000000000",
    284=>"110111111",
    285=>"000000000",
    286=>"000100000",
    287=>"000111010",
    288=>"111111111",
    289=>"100100100",
    290=>"111111111",
    291=>"101001000",
    292=>"001011000",
    293=>"000000000",
    294=>"000010000",
    295=>"111000000",
    296=>"000000000",
    297=>"000000000",
    298=>"111011101",
    299=>"000000000",
    300=>"000000000",
    301=>"000000000",
    302=>"000000011",
    303=>"000110101",
    304=>"000010010",
    305=>"111111111",
    306=>"111111011",
    307=>"000010111",
    308=>"000100101",
    309=>"101000001",
    310=>"101000101",
    311=>"010011110",
    312=>"111111111",
    313=>"000000000",
    314=>"000000000",
    315=>"111111111",
    316=>"111010001",
    317=>"000000001",
    318=>"000000000",
    319=>"001100011",
    320=>"110100101",
    321=>"111111111",
    322=>"001000000",
    323=>"111111111",
    324=>"111111111",
    325=>"000000000",
    326=>"100000000",
    327=>"111101001",
    328=>"111111111",
    329=>"100100100",
    330=>"000000000",
    331=>"111111111",
    332=>"000100000",
    333=>"111111111",
    334=>"000000000",
    335=>"111111111",
    336=>"011100000",
    337=>"010000000",
    338=>"000000000",
    339=>"111111111",
    340=>"010000000",
    341=>"111000000",
    342=>"000000000",
    343=>"000111010",
    344=>"001100000",
    345=>"000000100",
    346=>"101011110",
    347=>"111100000",
    348=>"000000000",
    349=>"000111110",
    350=>"111111101",
    351=>"111111111",
    352=>"001001001",
    353=>"000000000",
    354=>"111010111",
    355=>"000000100",
    356=>"000000000",
    357=>"000000000",
    358=>"010010001",
    359=>"000000000",
    360=>"111111111",
    361=>"000000100",
    362=>"000000001",
    363=>"000000000",
    364=>"111110000",
    365=>"000000000",
    366=>"111111111",
    367=>"001101001",
    368=>"000010010",
    369=>"000111111",
    370=>"010000000",
    371=>"111111111",
    372=>"111111101",
    373=>"000000000",
    374=>"011111111",
    375=>"111111111",
    376=>"000000000",
    377=>"111001101",
    378=>"110111111",
    379=>"111101111",
    380=>"111111011",
    381=>"110000000",
    382=>"000001011",
    383=>"011111110",
    384=>"111111111",
    385=>"100000011",
    386=>"001101111",
    387=>"100000000",
    388=>"000011000",
    389=>"000000001",
    390=>"011010000",
    391=>"000101101",
    392=>"100000001",
    393=>"000000000",
    394=>"000010111",
    395=>"100100000",
    396=>"000000100",
    397=>"000000101",
    398=>"100000011",
    399=>"010100111",
    400=>"001000000",
    401=>"000011011",
    402=>"000010111",
    403=>"000010000",
    404=>"011010000",
    405=>"000000000",
    406=>"010000000",
    407=>"001110110",
    408=>"100000000",
    409=>"100011010",
    410=>"001011001",
    411=>"101000100",
    412=>"110110000",
    413=>"101010010",
    414=>"100000000",
    415=>"000001111",
    416=>"110111111",
    417=>"100110110",
    418=>"111011001",
    419=>"111111101",
    420=>"000010010",
    421=>"000011100",
    422=>"100111111",
    423=>"110100010",
    424=>"111100100",
    425=>"111111110",
    426=>"111110000",
    427=>"101110110",
    428=>"111011111",
    429=>"000000011",
    430=>"111100000",
    431=>"000100100",
    432=>"111000000",
    433=>"101001011",
    434=>"111011000",
    435=>"000000000",
    436=>"100011000",
    437=>"000000000",
    438=>"100000000",
    439=>"111111111",
    440=>"000010111",
    441=>"111111111",
    442=>"000000000",
    443=>"000000000",
    444=>"000111111",
    445=>"011111111",
    446=>"100100011",
    447=>"110100000",
    448=>"010000111",
    449=>"000000000",
    450=>"011111111",
    451=>"000000111",
    452=>"000000000",
    453=>"110100000",
    454=>"000000000",
    455=>"010000000",
    456=>"000000000",
    457=>"000110000",
    458=>"111011100",
    459=>"100111001",
    460=>"011000110",
    461=>"011000000",
    462=>"111111011",
    463=>"111000000",
    464=>"111110000",
    465=>"110110100",
    466=>"111000000",
    467=>"111000000",
    468=>"001001000",
    469=>"000110110",
    470=>"111010100",
    471=>"000000000",
    472=>"111111111",
    473=>"001011000",
    474=>"000110101",
    475=>"000111110",
    476=>"111111000",
    477=>"011100110",
    478=>"100001001",
    479=>"001000010",
    480=>"001000000",
    481=>"010001001",
    482=>"010100110",
    483=>"000011111",
    484=>"010111010",
    485=>"001001010",
    486=>"000001000",
    487=>"100011001",
    488=>"000000001",
    489=>"101011010",
    490=>"011111001",
    491=>"011110000",
    492=>"000111111",
    493=>"000000000",
    494=>"000000000",
    495=>"100000100",
    496=>"000111111",
    497=>"111111111",
    498=>"000111011",
    499=>"111111000",
    500=>"100100111",
    501=>"000000001",
    502=>"111101111",
    503=>"111110100",
    504=>"011011000",
    505=>"010000000",
    506=>"000000110",
    507=>"000000111",
    508=>"100011111",
    509=>"100111110",
    510=>"001011111",
    511=>"011011100",
    512=>"011011011",
    513=>"010110000",
    514=>"110110000",
    515=>"000000000",
    516=>"000000100",
    517=>"110110100",
    518=>"001001001",
    519=>"101100101",
    520=>"100110100",
    521=>"111111011",
    522=>"100000000",
    523=>"001100000",
    524=>"100100000",
    525=>"111111110",
    526=>"000000000",
    527=>"000100111",
    528=>"010100000",
    529=>"000110000",
    530=>"111011011",
    531=>"110110100",
    532=>"110110000",
    533=>"001001011",
    534=>"000000001",
    535=>"000100111",
    536=>"000000000",
    537=>"110111111",
    538=>"001100100",
    539=>"001000000",
    540=>"000000101",
    541=>"001000001",
    542=>"111111111",
    543=>"011111111",
    544=>"110111111",
    545=>"001000000",
    546=>"110101000",
    547=>"000110100",
    548=>"001001000",
    549=>"100000101",
    550=>"110110000",
    551=>"001001001",
    552=>"100000001",
    553=>"001011111",
    554=>"110101111",
    555=>"111111011",
    556=>"001000101",
    557=>"001000001",
    558=>"100100100",
    559=>"001111111",
    560=>"100000000",
    561=>"110110110",
    562=>"111111100",
    563=>"100011011",
    564=>"111111111",
    565=>"001001001",
    566=>"001001001",
    567=>"000111000",
    568=>"100000010",
    569=>"100100110",
    570=>"110110100",
    571=>"010101000",
    572=>"111001011",
    573=>"100110010",
    574=>"000000100",
    575=>"110110110",
    576=>"110101000",
    577=>"100111111",
    578=>"011110110",
    579=>"000000000",
    580=>"100111000",
    581=>"100000010",
    582=>"001001000",
    583=>"110000000",
    584=>"100111010",
    585=>"011001001",
    586=>"000100110",
    587=>"001000001",
    588=>"000111110",
    589=>"011001000",
    590=>"111111110",
    591=>"001001111",
    592=>"110110010",
    593=>"001001001",
    594=>"110110100",
    595=>"111111111",
    596=>"111111111",
    597=>"110110000",
    598=>"000000000",
    599=>"110110110",
    600=>"000000000",
    601=>"110110110",
    602=>"000001101",
    603=>"001011011",
    604=>"100000000",
    605=>"111100000",
    606=>"101111111",
    607=>"100100100",
    608=>"100100001",
    609=>"010010000",
    610=>"110110111",
    611=>"001001001",
    612=>"010100000",
    613=>"100010001",
    614=>"001001001",
    615=>"000001001",
    616=>"110110000",
    617=>"010000100",
    618=>"111111011",
    619=>"111100111",
    620=>"000001001",
    621=>"001001001",
    622=>"100000001",
    623=>"110100100",
    624=>"100000111",
    625=>"000000100",
    626=>"000000110",
    627=>"011011000",
    628=>"100111110",
    629=>"000000000",
    630=>"110110000",
    631=>"100111111",
    632=>"110001101",
    633=>"001000111",
    634=>"011111111",
    635=>"011110100",
    636=>"101110111",
    637=>"101101111",
    638=>"110000000",
    639=>"100110000",
    640=>"000000111",
    641=>"100000101",
    642=>"001011100",
    643=>"100100000",
    644=>"111000001",
    645=>"000001011",
    646=>"000000101",
    647=>"000011010",
    648=>"111110110",
    649=>"111111110",
    650=>"111101000",
    651=>"001101100",
    652=>"101000000",
    653=>"010110111",
    654=>"111100100",
    655=>"110110000",
    656=>"100100100",
    657=>"101100000",
    658=>"000101011",
    659=>"111110110",
    660=>"111101111",
    661=>"010111011",
    662=>"101011100",
    663=>"111000000",
    664=>"110100100",
    665=>"101100001",
    666=>"110101000",
    667=>"000000000",
    668=>"000000000",
    669=>"010110100",
    670=>"000000000",
    671=>"011011000",
    672=>"000111011",
    673=>"100000100",
    674=>"111101011",
    675=>"000010110",
    676=>"011011001",
    677=>"000101001",
    678=>"111000010",
    679=>"000000111",
    680=>"111000000",
    681=>"111100000",
    682=>"000000100",
    683=>"000110110",
    684=>"011001000",
    685=>"011011111",
    686=>"010111111",
    687=>"111111111",
    688=>"110000111",
    689=>"000001110",
    690=>"001000100",
    691=>"110100011",
    692=>"000000100",
    693=>"001101100",
    694=>"101000000",
    695=>"000000010",
    696=>"100100000",
    697=>"111100000",
    698=>"100011011",
    699=>"101000000",
    700=>"000011011",
    701=>"001001010",
    702=>"000100110",
    703=>"010100001",
    704=>"001110010",
    705=>"000000100",
    706=>"111111001",
    707=>"000000000",
    708=>"110101011",
    709=>"000010100",
    710=>"000111011",
    711=>"011101111",
    712=>"000000000",
    713=>"000000111",
    714=>"111011000",
    715=>"100000011",
    716=>"011011000",
    717=>"000111111",
    718=>"011111000",
    719=>"000011111",
    720=>"111011000",
    721=>"110110100",
    722=>"110000111",
    723=>"000000011",
    724=>"000100000",
    725=>"100111000",
    726=>"101101000",
    727=>"000000111",
    728=>"001000100",
    729=>"011111111",
    730=>"110000000",
    731=>"111011011",
    732=>"000110101",
    733=>"000001011",
    734=>"110100000",
    735=>"111111100",
    736=>"100001011",
    737=>"001011111",
    738=>"010111111",
    739=>"010111100",
    740=>"001000010",
    741=>"000011000",
    742=>"001001001",
    743=>"011101111",
    744=>"000000001",
    745=>"111000000",
    746=>"010110001",
    747=>"111011000",
    748=>"000101101",
    749=>"000010111",
    750=>"100000001",
    751=>"101001001",
    752=>"111111001",
    753=>"011011011",
    754=>"111011011",
    755=>"100000000",
    756=>"000000000",
    757=>"000000111",
    758=>"101000010",
    759=>"010000000",
    760=>"011011001",
    761=>"101000100",
    762=>"000100100",
    763=>"000000000",
    764=>"001000110",
    765=>"100100111",
    766=>"111110100",
    767=>"111110101",
    768=>"111010111",
    769=>"111111111",
    770=>"010000000",
    771=>"000100000",
    772=>"011000000",
    773=>"101111100",
    774=>"010000100",
    775=>"111111010",
    776=>"000111000",
    777=>"111111100",
    778=>"101000000",
    779=>"001000100",
    780=>"000111011",
    781=>"000111100",
    782=>"000011000",
    783=>"000000011",
    784=>"001111101",
    785=>"111100111",
    786=>"000000000",
    787=>"000001001",
    788=>"010110010",
    789=>"010011000",
    790=>"000111111",
    791=>"010000000",
    792=>"001100111",
    793=>"110100000",
    794=>"000111000",
    795=>"000011111",
    796=>"000001111",
    797=>"100110100",
    798=>"111011001",
    799=>"000000001",
    800=>"100100100",
    801=>"000001000",
    802=>"001001000",
    803=>"111101010",
    804=>"001101111",
    805=>"000010000",
    806=>"000010111",
    807=>"000000100",
    808=>"000100110",
    809=>"100000000",
    810=>"011101001",
    811=>"011111011",
    812=>"111011001",
    813=>"000010000",
    814=>"000000000",
    815=>"111111111",
    816=>"101100110",
    817=>"010010000",
    818=>"011001100",
    819=>"000010111",
    820=>"000000000",
    821=>"010001001",
    822=>"000101001",
    823=>"111101111",
    824=>"000001001",
    825=>"010101111",
    826=>"010011010",
    827=>"000000100",
    828=>"000110000",
    829=>"111101111",
    830=>"001010111",
    831=>"010101111",
    832=>"111111000",
    833=>"111111011",
    834=>"111000001",
    835=>"111000101",
    836=>"101000011",
    837=>"010010010",
    838=>"000111000",
    839=>"110010001",
    840=>"100111001",
    841=>"010000010",
    842=>"000000110",
    843=>"010110010",
    844=>"101101000",
    845=>"111000100",
    846=>"100000100",
    847=>"101000001",
    848=>"000100010",
    849=>"000111110",
    850=>"000010010",
    851=>"111111010",
    852=>"110010010",
    853=>"100111110",
    854=>"100111000",
    855=>"101100111",
    856=>"111000000",
    857=>"111110001",
    858=>"001000000",
    859=>"111101101",
    860=>"110100100",
    861=>"010000010",
    862=>"001011111",
    863=>"111111111",
    864=>"100100111",
    865=>"001000100",
    866=>"000000000",
    867=>"000000000",
    868=>"100110001",
    869=>"111110110",
    870=>"100111011",
    871=>"001001111",
    872=>"000000010",
    873=>"000100100",
    874=>"000011011",
    875=>"111111000",
    876=>"111000101",
    877=>"000001000",
    878=>"010110110",
    879=>"111001100",
    880=>"000000000",
    881=>"111111001",
    882=>"101110000",
    883=>"000101000",
    884=>"111101111",
    885=>"111111000",
    886=>"000000000",
    887=>"111110000",
    888=>"111110000",
    889=>"100100000",
    890=>"100000000",
    891=>"000000000",
    892=>"001001001",
    893=>"000000001",
    894=>"111110110",
    895=>"110111111",
    896=>"010011100",
    897=>"000000111",
    898=>"000001111",
    899=>"010000000",
    900=>"110110001",
    901=>"110010000",
    902=>"010000000",
    903=>"000000000",
    904=>"111000000",
    905=>"000000000",
    906=>"000100110",
    907=>"000000111",
    908=>"011100100",
    909=>"111110111",
    910=>"010000000",
    911=>"000001111",
    912=>"111010000",
    913=>"111111000",
    914=>"111000000",
    915=>"001011111",
    916=>"000100111",
    917=>"001000111",
    918=>"000000000",
    919=>"100011101",
    920=>"101000000",
    921=>"100000111",
    922=>"100100011",
    923=>"110000110",
    924=>"001111010",
    925=>"111100000",
    926=>"011000000",
    927=>"111111010",
    928=>"111000000",
    929=>"110100000",
    930=>"111110010",
    931=>"010010000",
    932=>"010000000",
    933=>"110101111",
    934=>"110110000",
    935=>"000000101",
    936=>"001010111",
    937=>"110001111",
    938=>"001000000",
    939=>"011001000",
    940=>"110110111",
    941=>"011010000",
    942=>"111111000",
    943=>"111000000",
    944=>"001101001",
    945=>"100000000",
    946=>"111111001",
    947=>"011000000",
    948=>"011111100",
    949=>"101001000",
    950=>"000101011",
    951=>"111000000",
    952=>"000000101",
    953=>"111001101",
    954=>"000100000",
    955=>"000001111",
    956=>"000100101",
    957=>"111010000",
    958=>"110000001",
    959=>"101001000",
    960=>"001011101",
    961=>"111110000",
    962=>"010000000",
    963=>"000000111",
    964=>"011011100",
    965=>"111010000",
    966=>"101101000",
    967=>"011110001",
    968=>"111010000",
    969=>"101111010",
    970=>"100110000",
    971=>"111100000",
    972=>"110101000",
    973=>"111011001",
    974=>"010100000",
    975=>"100000111",
    976=>"100111010",
    977=>"000001011",
    978=>"000100111",
    979=>"110000000",
    980=>"011011000",
    981=>"000000101",
    982=>"111011000",
    983=>"000001001",
    984=>"011100110",
    985=>"111001000",
    986=>"000000100",
    987=>"111110001",
    988=>"111000000",
    989=>"100100111",
    990=>"000000001",
    991=>"111111101",
    992=>"111010000",
    993=>"011000101",
    994=>"000101111",
    995=>"000000000",
    996=>"010000000",
    997=>"000000101",
    998=>"000000110",
    999=>"101110110",
    1000=>"011011111",
    1001=>"000001011",
    1002=>"111011000",
    1003=>"110110000",
    1004=>"000000101",
    1005=>"000001111",
    1006=>"001001000",
    1007=>"110000000",
    1008=>"000000011",
    1009=>"000000100",
    1010=>"111111010",
    1011=>"000001111",
    1012=>"000000100",
    1013=>"001000101",
    1014=>"101010000",
    1015=>"100011100",
    1016=>"011000000",
    1017=>"001000000",
    1018=>"001000011",
    1019=>"111110000",
    1020=>"000000000",
    1021=>"010001010",
    1022=>"111101010",
    1023=>"111111110",
    1024=>"111100010",
    1025=>"000000111",
    1026=>"000110100",
    1027=>"000010000",
    1028=>"101101111",
    1029=>"111000000",
    1030=>"110100100",
    1031=>"010000000",
    1032=>"000000000",
    1033=>"100100100",
    1034=>"111101000",
    1035=>"011111010",
    1036=>"000000100",
    1037=>"111111100",
    1038=>"111001001",
    1039=>"110011001",
    1040=>"011011001",
    1041=>"000001011",
    1042=>"111111111",
    1043=>"110101001",
    1044=>"011011011",
    1045=>"010000000",
    1046=>"011100000",
    1047=>"010011010",
    1048=>"101111101",
    1049=>"111111001",
    1050=>"001101110",
    1051=>"001011111",
    1052=>"000000010",
    1053=>"110110111",
    1054=>"100100111",
    1055=>"011011011",
    1056=>"111000010",
    1057=>"000001001",
    1058=>"101100000",
    1059=>"011101101",
    1060=>"110001000",
    1061=>"101001010",
    1062=>"001110111",
    1063=>"011111111",
    1064=>"111010100",
    1065=>"111111111",
    1066=>"111011111",
    1067=>"110100011",
    1068=>"100100110",
    1069=>"001010100",
    1070=>"100000010",
    1071=>"101101111",
    1072=>"111011001",
    1073=>"010111100",
    1074=>"100111110",
    1075=>"011011011",
    1076=>"101101111",
    1077=>"000100110",
    1078=>"000000101",
    1079=>"101000000",
    1080=>"000001010",
    1081=>"101101111",
    1082=>"001000000",
    1083=>"000000000",
    1084=>"000000110",
    1085=>"100100111",
    1086=>"110111011",
    1087=>"011001011",
    1088=>"111101000",
    1089=>"000000000",
    1090=>"101011011",
    1091=>"000000000",
    1092=>"110001001",
    1093=>"110010010",
    1094=>"111110000",
    1095=>"000010011",
    1096=>"010110100",
    1097=>"001000000",
    1098=>"111110110",
    1099=>"000000100",
    1100=>"011010111",
    1101=>"010010001",
    1102=>"010010111",
    1103=>"011011000",
    1104=>"011011011",
    1105=>"110001001",
    1106=>"111110000",
    1107=>"110000000",
    1108=>"011001000",
    1109=>"001010000",
    1110=>"111111011",
    1111=>"101000000",
    1112=>"111110111",
    1113=>"000101100",
    1114=>"000001001",
    1115=>"110010010",
    1116=>"110011001",
    1117=>"001011101",
    1118=>"000000000",
    1119=>"100100000",
    1120=>"010011011",
    1121=>"111110110",
    1122=>"111011000",
    1123=>"000101000",
    1124=>"111111111",
    1125=>"011010100",
    1126=>"001000000",
    1127=>"000100000",
    1128=>"000000001",
    1129=>"000100100",
    1130=>"111101001",
    1131=>"000000001",
    1132=>"111100000",
    1133=>"011111111",
    1134=>"111001111",
    1135=>"100100100",
    1136=>"111000100",
    1137=>"100100111",
    1138=>"100000000",
    1139=>"000000000",
    1140=>"101100100",
    1141=>"000001011",
    1142=>"000000100",
    1143=>"000001010",
    1144=>"001111110",
    1145=>"000000000",
    1146=>"000000100",
    1147=>"110110111",
    1148=>"000110110",
    1149=>"100101111",
    1150=>"111111110",
    1151=>"000000001",
    1152=>"111111111",
    1153=>"010111111",
    1154=>"000111111",
    1155=>"110110111",
    1156=>"001000000",
    1157=>"000000000",
    1158=>"111111111",
    1159=>"000000000",
    1160=>"000001001",
    1161=>"000000101",
    1162=>"111101000",
    1163=>"011001100",
    1164=>"000111111",
    1165=>"010110000",
    1166=>"000100000",
    1167=>"110101010",
    1168=>"111111111",
    1169=>"000010000",
    1170=>"001000000",
    1171=>"000100000",
    1172=>"010000101",
    1173=>"111100000",
    1174=>"111101011",
    1175=>"000000010",
    1176=>"100000000",
    1177=>"100100000",
    1178=>"001000000",
    1179=>"111110000",
    1180=>"111111011",
    1181=>"111000000",
    1182=>"001000000",
    1183=>"011010000",
    1184=>"010000000",
    1185=>"111100100",
    1186=>"001000000",
    1187=>"011100111",
    1188=>"111111111",
    1189=>"010000000",
    1190=>"011111000",
    1191=>"111111111",
    1192=>"111111000",
    1193=>"111110001",
    1194=>"111110000",
    1195=>"100000000",
    1196=>"011000101",
    1197=>"011100111",
    1198=>"111000000",
    1199=>"000111010",
    1200=>"111000000",
    1201=>"001111111",
    1202=>"001000000",
    1203=>"000100010",
    1204=>"100000000",
    1205=>"100001000",
    1206=>"000000111",
    1207=>"000000111",
    1208=>"111111110",
    1209=>"111111110",
    1210=>"000000011",
    1211=>"000000000",
    1212=>"011111000",
    1213=>"000000000",
    1214=>"111000000",
    1215=>"010111111",
    1216=>"110111001",
    1217=>"000000101",
    1218=>"111001000",
    1219=>"000000000",
    1220=>"100111011",
    1221=>"000000001",
    1222=>"000111000",
    1223=>"111101000",
    1224=>"111111111",
    1225=>"001000000",
    1226=>"111001000",
    1227=>"111110010",
    1228=>"111100000",
    1229=>"111111101",
    1230=>"100000000",
    1231=>"000111111",
    1232=>"011111000",
    1233=>"110111110",
    1234=>"000000000",
    1235=>"111011111",
    1236=>"000000000",
    1237=>"000101000",
    1238=>"001000000",
    1239=>"000000110",
    1240=>"010000000",
    1241=>"100000010",
    1242=>"000000000",
    1243=>"000111111",
    1244=>"100100000",
    1245=>"001111111",
    1246=>"000001000",
    1247=>"000001000",
    1248=>"001100100",
    1249=>"111111101",
    1250=>"110111111",
    1251=>"100011011",
    1252=>"101111111",
    1253=>"111111111",
    1254=>"111111011",
    1255=>"111111111",
    1256=>"111111111",
    1257=>"100000000",
    1258=>"100100000",
    1259=>"111011111",
    1260=>"110110010",
    1261=>"111000000",
    1262=>"111111111",
    1263=>"000001000",
    1264=>"000001111",
    1265=>"000010010",
    1266=>"000101000",
    1267=>"001101111",
    1268=>"000111000",
    1269=>"001001000",
    1270=>"111111010",
    1271=>"100000000",
    1272=>"011111101",
    1273=>"111111000",
    1274=>"110111111",
    1275=>"111111111",
    1276=>"000000000",
    1277=>"011111101",
    1278=>"111110000",
    1279=>"000010000",
    1280=>"101001100",
    1281=>"100111001",
    1282=>"111111011",
    1283=>"110011100",
    1284=>"111000001",
    1285=>"110111000",
    1286=>"010010011",
    1287=>"011000110",
    1288=>"001111011",
    1289=>"110011011",
    1290=>"110000000",
    1291=>"111111111",
    1292=>"110110110",
    1293=>"111111100",
    1294=>"101100101",
    1295=>"000000000",
    1296=>"011010110",
    1297=>"100011111",
    1298=>"001110000",
    1299=>"110100100",
    1300=>"000000110",
    1301=>"100010000",
    1302=>"101100011",
    1303=>"001000011",
    1304=>"010011001",
    1305=>"000000000",
    1306=>"100001110",
    1307=>"110000000",
    1308=>"100001010",
    1309=>"100110100",
    1310=>"111110110",
    1311=>"111101111",
    1312=>"000000000",
    1313=>"000100000",
    1314=>"000000000",
    1315=>"000100000",
    1316=>"010011001",
    1317=>"110010110",
    1318=>"111110010",
    1319=>"100011001",
    1320=>"001011111",
    1321=>"111001011",
    1322=>"000000100",
    1323=>"100101001",
    1324=>"011001000",
    1325=>"011011000",
    1326=>"110000010",
    1327=>"111111111",
    1328=>"110011010",
    1329=>"001100001",
    1330=>"111111111",
    1331=>"110010010",
    1332=>"100111110",
    1333=>"000001000",
    1334=>"011000000",
    1335=>"010111010",
    1336=>"001000001",
    1337=>"111100100",
    1338=>"011001001",
    1339=>"000000000",
    1340=>"111111111",
    1341=>"100001101",
    1342=>"000101110",
    1343=>"001000100",
    1344=>"110111101",
    1345=>"000000001",
    1346=>"010010011",
    1347=>"110111011",
    1348=>"110101100",
    1349=>"110110010",
    1350=>"111111000",
    1351=>"000100110",
    1352=>"100111100",
    1353=>"100111101",
    1354=>"011000010",
    1355=>"000000000",
    1356=>"000000100",
    1357=>"001101101",
    1358=>"111111000",
    1359=>"001111000",
    1360=>"100110010",
    1361=>"100111001",
    1362=>"001100111",
    1363=>"111010110",
    1364=>"011010000",
    1365=>"110111010",
    1366=>"100111011",
    1367=>"011000101",
    1368=>"111111000",
    1369=>"110000001",
    1370=>"111111110",
    1371=>"110000000",
    1372=>"000100001",
    1373=>"011000010",
    1374=>"010011000",
    1375=>"100010011",
    1376=>"111111001",
    1377=>"000001000",
    1378=>"110111011",
    1379=>"010011010",
    1380=>"011110111",
    1381=>"000011000",
    1382=>"000000000",
    1383=>"011000010",
    1384=>"000000000",
    1385=>"111111001",
    1386=>"000101011",
    1387=>"111001010",
    1388=>"010010000",
    1389=>"011001111",
    1390=>"100100001",
    1391=>"110000100",
    1392=>"000000110",
    1393=>"011110111",
    1394=>"110110001",
    1395=>"000110000",
    1396=>"111101111",
    1397=>"000000000",
    1398=>"011001110",
    1399=>"000000000",
    1400=>"001000100",
    1401=>"010001000",
    1402=>"111111111",
    1403=>"011000000",
    1404=>"001100001",
    1405=>"111100111",
    1406=>"110011011",
    1407=>"111111111",
    1408=>"011101011",
    1409=>"000000000",
    1410=>"000000000",
    1411=>"111111101",
    1412=>"011011111",
    1413=>"111000101",
    1414=>"111111110",
    1415=>"111111111",
    1416=>"011011111",
    1417=>"011111111",
    1418=>"000111110",
    1419=>"011000110",
    1420=>"001000000",
    1421=>"010111111",
    1422=>"000010011",
    1423=>"000011011",
    1424=>"010111100",
    1425=>"010111000",
    1426=>"001010000",
    1427=>"110100101",
    1428=>"000111111",
    1429=>"111001101",
    1430=>"100000111",
    1431=>"100111111",
    1432=>"111100100",
    1433=>"100100111",
    1434=>"100101101",
    1435=>"001001011",
    1436=>"111110110",
    1437=>"001001110",
    1438=>"011111001",
    1439=>"011100010",
    1440=>"111101111",
    1441=>"010111110",
    1442=>"011001100",
    1443=>"001111110",
    1444=>"111000000",
    1445=>"001000100",
    1446=>"101000010",
    1447=>"111111101",
    1448=>"111100000",
    1449=>"110100111",
    1450=>"011001101",
    1451=>"100101011",
    1452=>"000110110",
    1453=>"000111010",
    1454=>"110111111",
    1455=>"111000000",
    1456=>"000100000",
    1457=>"101000101",
    1458=>"100100111",
    1459=>"011001000",
    1460=>"101101100",
    1461=>"010010000",
    1462=>"000111111",
    1463=>"000010100",
    1464=>"000000000",
    1465=>"000000110",
    1466=>"011001111",
    1467=>"111000101",
    1468=>"101000000",
    1469=>"000110010",
    1470=>"110111110",
    1471=>"001011101",
    1472=>"111001000",
    1473=>"111111000",
    1474=>"101111110",
    1475=>"110111111",
    1476=>"110111000",
    1477=>"011011101",
    1478=>"101100111",
    1479=>"000000010",
    1480=>"111000001",
    1481=>"010101001",
    1482=>"111001111",
    1483=>"100000000",
    1484=>"111100101",
    1485=>"001111010",
    1486=>"111111000",
    1487=>"101000000",
    1488=>"000110000",
    1489=>"111011011",
    1490=>"111111111",
    1491=>"000000000",
    1492=>"111110111",
    1493=>"001000000",
    1494=>"000111111",
    1495=>"000110010",
    1496=>"001110110",
    1497=>"101101100",
    1498=>"001001010",
    1499=>"000010000",
    1500=>"000101011",
    1501=>"011000100",
    1502=>"101001001",
    1503=>"101000000",
    1504=>"100111010",
    1505=>"111000000",
    1506=>"111111111",
    1507=>"000000000",
    1508=>"111010010",
    1509=>"110011000",
    1510=>"111110110",
    1511=>"010000111",
    1512=>"011011000",
    1513=>"100100100",
    1514=>"000101001",
    1515=>"010010011",
    1516=>"010000000",
    1517=>"111000101",
    1518=>"000000011",
    1519=>"000100100",
    1520=>"010010000",
    1521=>"101100010",
    1522=>"111010000",
    1523=>"001000001",
    1524=>"101000011",
    1525=>"000000000",
    1526=>"110000000",
    1527=>"011001000",
    1528=>"001000110",
    1529=>"000000111",
    1530=>"110110100",
    1531=>"111001100",
    1532=>"100100001",
    1533=>"001010010",
    1534=>"000000000",
    1535=>"110101101",
    1536=>"111001101",
    1537=>"000000000",
    1538=>"110111111",
    1539=>"111001000",
    1540=>"101100101",
    1541=>"111010100",
    1542=>"111111111",
    1543=>"111111100",
    1544=>"001000000",
    1545=>"111111100",
    1546=>"011000000",
    1547=>"001001001",
    1548=>"000000000",
    1549=>"010010010",
    1550=>"111111011",
    1551=>"110111011",
    1552=>"000000000",
    1553=>"011111000",
    1554=>"001111110",
    1555=>"111000000",
    1556=>"111111001",
    1557=>"110010101",
    1558=>"010000000",
    1559=>"011111110",
    1560=>"110011111",
    1561=>"100000101",
    1562=>"111111111",
    1563=>"111111111",
    1564=>"110101111",
    1565=>"111011110",
    1566=>"101111111",
    1567=>"000100111",
    1568=>"101000000",
    1569=>"111111110",
    1570=>"001100001",
    1571=>"111011111",
    1572=>"011001000",
    1573=>"111111111",
    1574=>"000000000",
    1575=>"111111001",
    1576=>"111111111",
    1577=>"000111111",
    1578=>"000000100",
    1579=>"111101000",
    1580=>"000110000",
    1581=>"000001000",
    1582=>"111111001",
    1583=>"010011111",
    1584=>"000000000",
    1585=>"000111111",
    1586=>"111000110",
    1587=>"000111111",
    1588=>"000110111",
    1589=>"000000000",
    1590=>"000000000",
    1591=>"100001001",
    1592=>"000000000",
    1593=>"011011110",
    1594=>"101101000",
    1595=>"000000000",
    1596=>"000001000",
    1597=>"111111010",
    1598=>"111111111",
    1599=>"111110011",
    1600=>"100101011",
    1601=>"111111111",
    1602=>"010101111",
    1603=>"000111111",
    1604=>"111001111",
    1605=>"110110110",
    1606=>"000110000",
    1607=>"111110000",
    1608=>"000000000",
    1609=>"111101111",
    1610=>"011101101",
    1611=>"111111111",
    1612=>"111010000",
    1613=>"000000000",
    1614=>"111110010",
    1615=>"111110000",
    1616=>"000000000",
    1617=>"110001000",
    1618=>"111111111",
    1619=>"111110110",
    1620=>"111001001",
    1621=>"100111111",
    1622=>"111101111",
    1623=>"010110101",
    1624=>"101100011",
    1625=>"010110110",
    1626=>"001010010",
    1627=>"111011000",
    1628=>"101101101",
    1629=>"011011001",
    1630=>"000000000",
    1631=>"111111010",
    1632=>"000000000",
    1633=>"000000010",
    1634=>"000000000",
    1635=>"001101110",
    1636=>"111111111",
    1637=>"000000111",
    1638=>"001100000",
    1639=>"110101111",
    1640=>"000000000",
    1641=>"101100110",
    1642=>"100100010",
    1643=>"000101001",
    1644=>"101000000",
    1645=>"010010101",
    1646=>"010111111",
    1647=>"110111111",
    1648=>"111111111",
    1649=>"011111111",
    1650=>"000000000",
    1651=>"010000100",
    1652=>"000000000",
    1653=>"000000000",
    1654=>"000000000",
    1655=>"110011011",
    1656=>"011010100",
    1657=>"000000000",
    1658=>"000000000",
    1659=>"000000000",
    1660=>"000100000",
    1661=>"000000000",
    1662=>"111111101",
    1663=>"110111111",
    1664=>"101101100",
    1665=>"101101111",
    1666=>"110111110",
    1667=>"010011111",
    1668=>"011001011",
    1669=>"101100111",
    1670=>"001101001",
    1671=>"111000101",
    1672=>"110111000",
    1673=>"111110000",
    1674=>"111010000",
    1675=>"010000000",
    1676=>"000000000",
    1677=>"111111010",
    1678=>"111101101",
    1679=>"110010000",
    1680=>"010011111",
    1681=>"111101111",
    1682=>"000000010",
    1683=>"110100100",
    1684=>"000111111",
    1685=>"101000111",
    1686=>"000000000",
    1687=>"010000001",
    1688=>"001001010",
    1689=>"110100000",
    1690=>"011101100",
    1691=>"000010100",
    1692=>"000000100",
    1693=>"011011011",
    1694=>"100110111",
    1695=>"101111111",
    1696=>"001101011",
    1697=>"100100101",
    1698=>"011101000",
    1699=>"111111111",
    1700=>"110011000",
    1701=>"010111110",
    1702=>"000011101",
    1703=>"010111111",
    1704=>"111000000",
    1705=>"000000011",
    1706=>"000001111",
    1707=>"110100101",
    1708=>"111001000",
    1709=>"111111101",
    1710=>"000000000",
    1711=>"100000000",
    1712=>"010111100",
    1713=>"000000000",
    1714=>"000100000",
    1715=>"010010010",
    1716=>"110100101",
    1717=>"001001000",
    1718=>"111111100",
    1719=>"000011000",
    1720=>"111100101",
    1721=>"001000111",
    1722=>"011011011",
    1723=>"111001101",
    1724=>"000000000",
    1725=>"000000111",
    1726=>"000110011",
    1727=>"000100011",
    1728=>"111110000",
    1729=>"000111111",
    1730=>"110111111",
    1731=>"000000110",
    1732=>"111101111",
    1733=>"010110111",
    1734=>"101101010",
    1735=>"110000010",
    1736=>"100111101",
    1737=>"010110110",
    1738=>"111001000",
    1739=>"000000101",
    1740=>"000011010",
    1741=>"000000001",
    1742=>"011100111",
    1743=>"111110010",
    1744=>"010111000",
    1745=>"100110100",
    1746=>"000100010",
    1747=>"000100111",
    1748=>"110110111",
    1749=>"111101100",
    1750=>"001110111",
    1751=>"101111111",
    1752=>"001101110",
    1753=>"110111111",
    1754=>"100011011",
    1755=>"000000000",
    1756=>"001011111",
    1757=>"001011001",
    1758=>"100101101",
    1759=>"000000000",
    1760=>"001111110",
    1761=>"110100001",
    1762=>"111010010",
    1763=>"110000000",
    1764=>"100111111",
    1765=>"111111111",
    1766=>"001010011",
    1767=>"010000100",
    1768=>"001000000",
    1769=>"100000101",
    1770=>"110110100",
    1771=>"101111110",
    1772=>"000110111",
    1773=>"001000101",
    1774=>"110100111",
    1775=>"000001111",
    1776=>"010010010",
    1777=>"000000111",
    1778=>"000010110",
    1779=>"111001000",
    1780=>"111111111",
    1781=>"000101000",
    1782=>"000000111",
    1783=>"000001111",
    1784=>"101111111",
    1785=>"110111101",
    1786=>"000101000",
    1787=>"000000111",
    1788=>"011101110",
    1789=>"000001000",
    1790=>"010000000",
    1791=>"110100010",
    1792=>"011001011",
    1793=>"111111100",
    1794=>"001001001",
    1795=>"001001001",
    1796=>"001001000",
    1797=>"000010101",
    1798=>"101000011",
    1799=>"110000110",
    1800=>"011001001",
    1801=>"000100000",
    1802=>"011100001",
    1803=>"000100001",
    1804=>"110110000",
    1805=>"100100011",
    1806=>"101101011",
    1807=>"110011111",
    1808=>"010011000",
    1809=>"000100000",
    1810=>"001001011",
    1811=>"000000011",
    1812=>"110110000",
    1813=>"110100000",
    1814=>"011000110",
    1815=>"110101110",
    1816=>"001001011",
    1817=>"110100000",
    1818=>"001001001",
    1819=>"101000101",
    1820=>"001101001",
    1821=>"000101001",
    1822=>"011000001",
    1823=>"110000001",
    1824=>"000000001",
    1825=>"000000001",
    1826=>"001100000",
    1827=>"110010100",
    1828=>"111110110",
    1829=>"111110100",
    1830=>"010010110",
    1831=>"011011110",
    1832=>"100100001",
    1833=>"000001011",
    1834=>"011101001",
    1835=>"001001011",
    1836=>"000000100",
    1837=>"000001000",
    1838=>"000000000",
    1839=>"001001111",
    1840=>"111101110",
    1841=>"010110110",
    1842=>"100000000",
    1843=>"000001011",
    1844=>"001011011",
    1845=>"111100100",
    1846=>"110100001",
    1847=>"111111000",
    1848=>"111011000",
    1849=>"111001011",
    1850=>"101110111",
    1851=>"011110010",
    1852=>"101000000",
    1853=>"110000000",
    1854=>"000000000",
    1855=>"110110011",
    1856=>"111111101",
    1857=>"110000111",
    1858=>"110111000",
    1859=>"011101100",
    1860=>"101001011",
    1861=>"111110010",
    1862=>"111110100",
    1863=>"100000110",
    1864=>"000001011",
    1865=>"011111000",
    1866=>"000000011",
    1867=>"110110000",
    1868=>"000000001",
    1869=>"111011010",
    1870=>"100100110",
    1871=>"110110110",
    1872=>"011010110",
    1873=>"000001110",
    1874=>"000000011",
    1875=>"011111011",
    1876=>"001001111",
    1877=>"110110110",
    1878=>"011011011",
    1879=>"101011101",
    1880=>"001001001",
    1881=>"000101011",
    1882=>"101101011",
    1883=>"001010100",
    1884=>"001001011",
    1885=>"111100100",
    1886=>"001001001",
    1887=>"000001011",
    1888=>"000001011",
    1889=>"100110110",
    1890=>"011111110",
    1891=>"111101001",
    1892=>"000001111",
    1893=>"111111111",
    1894=>"110110000",
    1895=>"100000011",
    1896=>"111110110",
    1897=>"100100000",
    1898=>"001001011",
    1899=>"110110111",
    1900=>"101000001",
    1901=>"100110100",
    1902=>"110110100",
    1903=>"001101001",
    1904=>"110110000",
    1905=>"000100100",
    1906=>"000000000",
    1907=>"111110010",
    1908=>"100110100",
    1909=>"000110100",
    1910=>"110000110",
    1911=>"110011011",
    1912=>"010000010",
    1913=>"110110010",
    1914=>"110100100",
    1915=>"110100111",
    1916=>"000100000",
    1917=>"001001111",
    1918=>"111111101",
    1919=>"000001011",
    1920=>"010010010",
    1921=>"000000001",
    1922=>"011000111",
    1923=>"111011111",
    1924=>"110100101",
    1925=>"001111111",
    1926=>"111111101",
    1927=>"011100101",
    1928=>"001111101",
    1929=>"010110100",
    1930=>"111101101",
    1931=>"101000000",
    1932=>"011001100",
    1933=>"111100000",
    1934=>"000100001",
    1935=>"000100101",
    1936=>"101111100",
    1937=>"100000000",
    1938=>"111111100",
    1939=>"011100100",
    1940=>"100000110",
    1941=>"000000000",
    1942=>"110000000",
    1943=>"111100101",
    1944=>"000101100",
    1945=>"111101000",
    1946=>"011010010",
    1947=>"001001011",
    1948=>"001001001",
    1949=>"011110100",
    1950=>"111001001",
    1951=>"110110101",
    1952=>"111101000",
    1953=>"000100001",
    1954=>"111111111",
    1955=>"000100111",
    1956=>"011011000",
    1957=>"101000000",
    1958=>"111100101",
    1959=>"011100000",
    1960=>"110000000",
    1961=>"111101111",
    1962=>"011100000",
    1963=>"000100001",
    1964=>"101101000",
    1965=>"111010100",
    1966=>"001111000",
    1967=>"111101101",
    1968=>"011100001",
    1969=>"000000000",
    1970=>"100011100",
    1971=>"011001001",
    1972=>"001000110",
    1973=>"000111100",
    1974=>"000011111",
    1975=>"000101111",
    1976=>"110111011",
    1977=>"000100001",
    1978=>"011100000",
    1979=>"000000001",
    1980=>"001000000",
    1981=>"000011111",
    1982=>"100100111",
    1983=>"101001001",
    1984=>"100011011",
    1985=>"100011111",
    1986=>"010101101",
    1987=>"001001111",
    1988=>"111011001",
    1989=>"001011100",
    1990=>"100100001",
    1991=>"000000000",
    1992=>"010011100",
    1993=>"000000011",
    1994=>"011000010",
    1995=>"011000001",
    1996=>"111111100",
    1997=>"111100010",
    1998=>"001000111",
    1999=>"111101101",
    2000=>"111101100",
    2001=>"001000000",
    2002=>"000000000",
    2003=>"111001101",
    2004=>"110110001",
    2005=>"101000100",
    2006=>"000101100",
    2007=>"000101111",
    2008=>"011011010",
    2009=>"111010100",
    2010=>"000111101",
    2011=>"110000010",
    2012=>"000010000",
    2013=>"000001101",
    2014=>"111101000",
    2015=>"000010111",
    2016=>"110110110",
    2017=>"101000110",
    2018=>"000011010",
    2019=>"000010110",
    2020=>"000011111",
    2021=>"011001000",
    2022=>"101000100",
    2023=>"111111111",
    2024=>"000100000",
    2025=>"100000110",
    2026=>"110100001",
    2027=>"111010000",
    2028=>"000000000",
    2029=>"000000010",
    2030=>"000011011",
    2031=>"001000010",
    2032=>"000000110",
    2033=>"111001101",
    2034=>"101111111",
    2035=>"001101000",
    2036=>"000010111",
    2037=>"100000000",
    2038=>"001000100",
    2039=>"000101101",
    2040=>"001011000",
    2041=>"011000000",
    2042=>"000100000",
    2043=>"111100100",
    2044=>"111111100",
    2045=>"000000100",
    2046=>"101011000",
    2047=>"110111010",
    2048=>"111111000",
    2049=>"000111111",
    2050=>"111000000",
    2051=>"000111111",
    2052=>"111100000",
    2053=>"011111111",
    2054=>"111010010",
    2055=>"000111111",
    2056=>"111000000",
    2057=>"000100111",
    2058=>"111000000",
    2059=>"011001100",
    2060=>"101111101",
    2061=>"010110110",
    2062=>"100001001",
    2063=>"000011010",
    2064=>"001011001",
    2065=>"010000110",
    2066=>"011111111",
    2067=>"111011000",
    2068=>"000000001",
    2069=>"001000000",
    2070=>"100000000",
    2071=>"011011111",
    2072=>"111001111",
    2073=>"111010000",
    2074=>"011011000",
    2075=>"101101101",
    2076=>"000001100",
    2077=>"000001001",
    2078=>"111100010",
    2079=>"010100111",
    2080=>"000010000",
    2081=>"000000000",
    2082=>"111011000",
    2083=>"100010000",
    2084=>"010101111",
    2085=>"000000111",
    2086=>"000100111",
    2087=>"101000000",
    2088=>"111110011",
    2089=>"000010011",
    2090=>"111000011",
    2091=>"111101001",
    2092=>"111100111",
    2093=>"000111000",
    2094=>"001111111",
    2095=>"111000001",
    2096=>"101111000",
    2097=>"000111011",
    2098=>"001110111",
    2099=>"111111001",
    2100=>"010100100",
    2101=>"000000001",
    2102=>"000111111",
    2103=>"000000111",
    2104=>"111000000",
    2105=>"101001111",
    2106=>"001001001",
    2107=>"101000000",
    2108=>"111000000",
    2109=>"111001101",
    2110=>"101101101",
    2111=>"011000011",
    2112=>"010010011",
    2113=>"111000000",
    2114=>"000111111",
    2115=>"000000000",
    2116=>"000001000",
    2117=>"111111111",
    2118=>"100010111",
    2119=>"100010111",
    2120=>"100110110",
    2121=>"000000000",
    2122=>"111010100",
    2123=>"001000000",
    2124=>"000010000",
    2125=>"010010100",
    2126=>"000000000",
    2127=>"100000111",
    2128=>"000111111",
    2129=>"111001001",
    2130=>"000000110",
    2131=>"000011111",
    2132=>"111111111",
    2133=>"000111111",
    2134=>"001110000",
    2135=>"111101001",
    2136=>"101110000",
    2137=>"010000110",
    2138=>"000101010",
    2139=>"111111011",
    2140=>"111001000",
    2141=>"100111011",
    2142=>"111000001",
    2143=>"111111011",
    2144=>"000001001",
    2145=>"100110100",
    2146=>"000010010",
    2147=>"111111111",
    2148=>"111000110",
    2149=>"100000000",
    2150=>"111100100",
    2151=>"011010100",
    2152=>"010111011",
    2153=>"111110100",
    2154=>"111101001",
    2155=>"000110111",
    2156=>"111000000",
    2157=>"000010000",
    2158=>"010110000",
    2159=>"011000100",
    2160=>"111000001",
    2161=>"101000111",
    2162=>"101000000",
    2163=>"000111110",
    2164=>"001001001",
    2165=>"101000000",
    2166=>"111000010",
    2167=>"110111111",
    2168=>"001110110",
    2169=>"000000000",
    2170=>"000110110",
    2171=>"111000000",
    2172=>"100001000",
    2173=>"000000111",
    2174=>"111110000",
    2175=>"010011110",
    2176=>"111101111",
    2177=>"000111000",
    2178=>"111000000",
    2179=>"100101111",
    2180=>"101000111",
    2181=>"010111111",
    2182=>"111110111",
    2183=>"101111111",
    2184=>"000000001",
    2185=>"000001101",
    2186=>"010010000",
    2187=>"000000000",
    2188=>"100010011",
    2189=>"010111000",
    2190=>"000000000",
    2191=>"111111111",
    2192=>"010111000",
    2193=>"111000000",
    2194=>"101001100",
    2195=>"010111111",
    2196=>"010000000",
    2197=>"111000100",
    2198=>"000000000",
    2199=>"111111111",
    2200=>"110000001",
    2201=>"000000000",
    2202=>"110111111",
    2203=>"101100110",
    2204=>"000011111",
    2205=>"000000000",
    2206=>"001000011",
    2207=>"010101111",
    2208=>"111111101",
    2209=>"100100100",
    2210=>"000100111",
    2211=>"001000010",
    2212=>"001111001",
    2213=>"110010000",
    2214=>"101111111",
    2215=>"111000001",
    2216=>"001101011",
    2217=>"111101111",
    2218=>"000001001",
    2219=>"110000100",
    2220=>"101111001",
    2221=>"000000101",
    2222=>"000000111",
    2223=>"111101010",
    2224=>"111111111",
    2225=>"000000000",
    2226=>"000000000",
    2227=>"000000111",
    2228=>"110101111",
    2229=>"110000000",
    2230=>"110110100",
    2231=>"111100000",
    2232=>"111111111",
    2233=>"110000000",
    2234=>"110100000",
    2235=>"000000111",
    2236=>"111110111",
    2237=>"001001101",
    2238=>"101011111",
    2239=>"111011111",
    2240=>"010111111",
    2241=>"011000101",
    2242=>"111011100",
    2243=>"111111111",
    2244=>"000000000",
    2245=>"011011111",
    2246=>"111000101",
    2247=>"101111011",
    2248=>"011111000",
    2249=>"000000001",
    2250=>"001001010",
    2251=>"101000100",
    2252=>"100000111",
    2253=>"000000111",
    2254=>"100101111",
    2255=>"000111111",
    2256=>"000100101",
    2257=>"000000000",
    2258=>"000000111",
    2259=>"111111010",
    2260=>"110110111",
    2261=>"000110010",
    2262=>"000000000",
    2263=>"000001111",
    2264=>"111100010",
    2265=>"000000000",
    2266=>"000100110",
    2267=>"011000010",
    2268=>"001001000",
    2269=>"000110010",
    2270=>"000100110",
    2271=>"110011011",
    2272=>"000100000",
    2273=>"000011011",
    2274=>"111111111",
    2275=>"111000000",
    2276=>"111111111",
    2277=>"001001011",
    2278=>"000000000",
    2279=>"000101011",
    2280=>"110111010",
    2281=>"011000000",
    2282=>"110000000",
    2283=>"011111111",
    2284=>"000000000",
    2285=>"001101111",
    2286=>"111111110",
    2287=>"000000000",
    2288=>"000000000",
    2289=>"010111111",
    2290=>"000000100",
    2291=>"000000100",
    2292=>"010000000",
    2293=>"100010000",
    2294=>"110101100",
    2295=>"100000000",
    2296=>"101100110",
    2297=>"111111111",
    2298=>"000111011",
    2299=>"000111110",
    2300=>"000001011",
    2301=>"101101000",
    2302=>"000000000",
    2303=>"110000111",
    2304=>"010010111",
    2305=>"010011110",
    2306=>"000010000",
    2307=>"000000000",
    2308=>"000110110",
    2309=>"000000000",
    2310=>"101001101",
    2311=>"011010010",
    2312=>"110110010",
    2313=>"001001000",
    2314=>"101000000",
    2315=>"000110111",
    2316=>"111111111",
    2317=>"000010000",
    2318=>"100110100",
    2319=>"100000000",
    2320=>"011011000",
    2321=>"010110000",
    2322=>"000011000",
    2323=>"000111111",
    2324=>"101000101",
    2325=>"000000110",
    2326=>"001100100",
    2327=>"000111111",
    2328=>"010011011",
    2329=>"001111111",
    2330=>"000101111",
    2331=>"110110100",
    2332=>"000000000",
    2333=>"011000111",
    2334=>"111100110",
    2335=>"111000000",
    2336=>"111111011",
    2337=>"110100100",
    2338=>"010110111",
    2339=>"000000010",
    2340=>"000000001",
    2341=>"101000000",
    2342=>"000011010",
    2343=>"000011000",
    2344=>"011111111",
    2345=>"011111111",
    2346=>"010111011",
    2347=>"010010010",
    2348=>"000001000",
    2349=>"000000000",
    2350=>"000100100",
    2351=>"010111010",
    2352=>"110100100",
    2353=>"000011000",
    2354=>"110111001",
    2355=>"110000000",
    2356=>"011011111",
    2357=>"110101101",
    2358=>"101100100",
    2359=>"111101001",
    2360=>"110110010",
    2361=>"111110111",
    2362=>"100100000",
    2363=>"000000010",
    2364=>"000110000",
    2365=>"000000000",
    2366=>"011001001",
    2367=>"111000111",
    2368=>"101100111",
    2369=>"111000001",
    2370=>"001000000",
    2371=>"111111111",
    2372=>"000000000",
    2373=>"000110100",
    2374=>"001000001",
    2375=>"010000001",
    2376=>"110010011",
    2377=>"111000000",
    2378=>"000110100",
    2379=>"000001010",
    2380=>"111111111",
    2381=>"010000000",
    2382=>"000000000",
    2383=>"000010000",
    2384=>"000000000",
    2385=>"000000001",
    2386=>"011000000",
    2387=>"000000000",
    2388=>"011001001",
    2389=>"001111100",
    2390=>"111100000",
    2391=>"111011111",
    2392=>"011001101",
    2393=>"000000010",
    2394=>"110111110",
    2395=>"111111010",
    2396=>"110110000",
    2397=>"000010110",
    2398=>"100110010",
    2399=>"010110000",
    2400=>"111001011",
    2401=>"000001000",
    2402=>"000010000",
    2403=>"000111111",
    2404=>"111001011",
    2405=>"010010110",
    2406=>"000000100",
    2407=>"011000000",
    2408=>"010111111",
    2409=>"000010110",
    2410=>"001001000",
    2411=>"000111010",
    2412=>"011111101",
    2413=>"000100111",
    2414=>"111000110",
    2415=>"000001001",
    2416=>"000000010",
    2417=>"010011111",
    2418=>"110111011",
    2419=>"110110010",
    2420=>"000000101",
    2421=>"110101111",
    2422=>"010010000",
    2423=>"010111110",
    2424=>"100111111",
    2425=>"000000110",
    2426=>"001111111",
    2427=>"011111110",
    2428=>"111001001",
    2429=>"111111001",
    2430=>"001111111",
    2431=>"011001011",
    2432=>"110101111",
    2433=>"111111000",
    2434=>"000000111",
    2435=>"111111101",
    2436=>"100100111",
    2437=>"111101110",
    2438=>"000000000",
    2439=>"111111000",
    2440=>"010011111",
    2441=>"111000010",
    2442=>"111110011",
    2443=>"110100111",
    2444=>"111110100",
    2445=>"110110110",
    2446=>"111100001",
    2447=>"010011001",
    2448=>"110111111",
    2449=>"110100000",
    2450=>"011001111",
    2451=>"010000111",
    2452=>"111111000",
    2453=>"000000111",
    2454=>"111000000",
    2455=>"010000101",
    2456=>"100011110",
    2457=>"100000110",
    2458=>"111011000",
    2459=>"111100000",
    2460=>"111101111",
    2461=>"000000001",
    2462=>"101110010",
    2463=>"111001000",
    2464=>"000111010",
    2465=>"111111111",
    2466=>"110000011",
    2467=>"000000000",
    2468=>"000100111",
    2469=>"111110000",
    2470=>"111111001",
    2471=>"000000111",
    2472=>"000010111",
    2473=>"000001111",
    2474=>"000000101",
    2475=>"000100010",
    2476=>"000111111",
    2477=>"111100001",
    2478=>"000111110",
    2479=>"111111000",
    2480=>"001111100",
    2481=>"001001111",
    2482=>"000100011",
    2483=>"000000100",
    2484=>"011001000",
    2485=>"000000000",
    2486=>"000000010",
    2487=>"000001111",
    2488=>"000000000",
    2489=>"000000010",
    2490=>"001010010",
    2491=>"100100000",
    2492=>"000000000",
    2493=>"000000110",
    2494=>"011001001",
    2495=>"110111000",
    2496=>"000011000",
    2497=>"001010000",
    2498=>"010000000",
    2499=>"111000010",
    2500=>"011110101",
    2501=>"000100110",
    2502=>"000000111",
    2503=>"000111000",
    2504=>"011110100",
    2505=>"000001111",
    2506=>"000110110",
    2507=>"111101000",
    2508=>"001101110",
    2509=>"000000111",
    2510=>"101111111",
    2511=>"100101111",
    2512=>"000100111",
    2513=>"000100001",
    2514=>"000111111",
    2515=>"111101000",
    2516=>"000000011",
    2517=>"000000000",
    2518=>"001001101",
    2519=>"000000000",
    2520=>"000100111",
    2521=>"001111101",
    2522=>"111000000",
    2523=>"110000000",
    2524=>"001011110",
    2525=>"100110101",
    2526=>"010000000",
    2527=>"000000101",
    2528=>"100100010",
    2529=>"001000111",
    2530=>"100001110",
    2531=>"111001000",
    2532=>"000110101",
    2533=>"011111000",
    2534=>"011001001",
    2535=>"001111111",
    2536=>"011111001",
    2537=>"100000000",
    2538=>"001001111",
    2539=>"000001111",
    2540=>"010000010",
    2541=>"111000000",
    2542=>"111001101",
    2543=>"111001101",
    2544=>"111001100",
    2545=>"000100000",
    2546=>"101000000",
    2547=>"111111001",
    2548=>"000000111",
    2549=>"100110000",
    2550=>"000111111",
    2551=>"001001100",
    2552=>"101111111",
    2553=>"100000010",
    2554=>"111100100",
    2555=>"000111110",
    2556=>"011001001",
    2557=>"111101101",
    2558=>"000000110",
    2559=>"111001111",
    2560=>"011001001",
    2561=>"111001101",
    2562=>"100010111",
    2563=>"111101001",
    2564=>"110001100",
    2565=>"110111110",
    2566=>"001100101",
    2567=>"000000000",
    2568=>"000011101",
    2569=>"001100100",
    2570=>"110101101",
    2571=>"011010000",
    2572=>"010101111",
    2573=>"110111110",
    2574=>"010001000",
    2575=>"010000011",
    2576=>"001001111",
    2577=>"010110000",
    2578=>"011100101",
    2579=>"111110001",
    2580=>"000000000",
    2581=>"000000001",
    2582=>"000011100",
    2583=>"010101001",
    2584=>"100001011",
    2585=>"110101000",
    2586=>"100011101",
    2587=>"100001001",
    2588=>"111111110",
    2589=>"010100101",
    2590=>"111111111",
    2591=>"000111111",
    2592=>"010111101",
    2593=>"000000100",
    2594=>"111111001",
    2595=>"111110000",
    2596=>"000111111",
    2597=>"000001000",
    2598=>"110000000",
    2599=>"000001111",
    2600=>"001010111",
    2601=>"111110000",
    2602=>"000001001",
    2603=>"000001010",
    2604=>"000001111",
    2605=>"000000000",
    2606=>"000000000",
    2607=>"101010000",
    2608=>"001010010",
    2609=>"000111000",
    2610=>"011001101",
    2611=>"000011011",
    2612=>"000000001",
    2613=>"001101111",
    2614=>"111110000",
    2615=>"000010010",
    2616=>"000000100",
    2617=>"110010001",
    2618=>"110101010",
    2619=>"111000000",
    2620=>"111000000",
    2621=>"111101101",
    2622=>"001101111",
    2623=>"100010000",
    2624=>"100100100",
    2625=>"011100000",
    2626=>"000100000",
    2627=>"000000000",
    2628=>"000100111",
    2629=>"100110001",
    2630=>"000110111",
    2631=>"111000101",
    2632=>"000100101",
    2633=>"000001101",
    2634=>"000000111",
    2635=>"001000000",
    2636=>"000111111",
    2637=>"000111000",
    2638=>"000000110",
    2639=>"101000111",
    2640=>"100000110",
    2641=>"000100000",
    2642=>"000000000",
    2643=>"000011010",
    2644=>"000101101",
    2645=>"000111010",
    2646=>"000000111",
    2647=>"010011111",
    2648=>"010001000",
    2649=>"101100000",
    2650=>"100000001",
    2651=>"000000010",
    2652=>"010100000",
    2653=>"001001100",
    2654=>"110101101",
    2655=>"111000000",
    2656=>"000100101",
    2657=>"000010110",
    2658=>"000000000",
    2659=>"000010000",
    2660=>"000000110",
    2661=>"001000011",
    2662=>"000011100",
    2663=>"001100000",
    2664=>"100000011",
    2665=>"111000000",
    2666=>"100001101",
    2667=>"111111000",
    2668=>"000010000",
    2669=>"000000000",
    2670=>"010111001",
    2671=>"100110011",
    2672=>"000110000",
    2673=>"111111100",
    2674=>"100101111",
    2675=>"111011000",
    2676=>"111100101",
    2677=>"000000111",
    2678=>"000000001",
    2679=>"110100001",
    2680=>"111011000",
    2681=>"101010000",
    2682=>"001000110",
    2683=>"011111110",
    2684=>"001001100",
    2685=>"111000000",
    2686=>"000000111",
    2687=>"111101101",
    2688=>"111101111",
    2689=>"100110111",
    2690=>"000000000",
    2691=>"000111000",
    2692=>"111101110",
    2693=>"111111000",
    2694=>"011111111",
    2695=>"001111100",
    2696=>"111011011",
    2697=>"011011110",
    2698=>"111111111",
    2699=>"100001111",
    2700=>"110110101",
    2701=>"111111110",
    2702=>"111010010",
    2703=>"000000010",
    2704=>"111110100",
    2705=>"000000000",
    2706=>"100100111",
    2707=>"100000001",
    2708=>"101001111",
    2709=>"000001111",
    2710=>"100000000",
    2711=>"111110110",
    2712=>"001001001",
    2713=>"010100001",
    2714=>"100000100",
    2715=>"110111111",
    2716=>"101011010",
    2717=>"110000000",
    2718=>"111111010",
    2719=>"011111110",
    2720=>"111110111",
    2721=>"111100110",
    2722=>"000111011",
    2723=>"011000110",
    2724=>"111110000",
    2725=>"000000000",
    2726=>"100100000",
    2727=>"110110000",
    2728=>"101100110",
    2729=>"000101111",
    2730=>"111001001",
    2731=>"000000000",
    2732=>"000000111",
    2733=>"011000000",
    2734=>"111011111",
    2735=>"111111000",
    2736=>"110001100",
    2737=>"111111000",
    2738=>"111111000",
    2739=>"000000000",
    2740=>"100100011",
    2741=>"000000000",
    2742=>"111111111",
    2743=>"000110111",
    2744=>"111110110",
    2745=>"111001011",
    2746=>"011110110",
    2747=>"111000000",
    2748=>"101000001",
    2749=>"011001011",
    2750=>"111111111",
    2751=>"000111111",
    2752=>"000000000",
    2753=>"000000000",
    2754=>"111001110",
    2755=>"001000110",
    2756=>"111110001",
    2757=>"111111111",
    2758=>"000110111",
    2759=>"101111011",
    2760=>"111011111",
    2761=>"111111111",
    2762=>"000000000",
    2763=>"000000000",
    2764=>"001010011",
    2765=>"111111011",
    2766=>"000111111",
    2767=>"111111111",
    2768=>"011000100",
    2769=>"000000100",
    2770=>"000000111",
    2771=>"010111011",
    2772=>"111111111",
    2773=>"110010000",
    2774=>"000000010",
    2775=>"111111011",
    2776=>"000001111",
    2777=>"101011101",
    2778=>"111011011",
    2779=>"111111110",
    2780=>"100100000",
    2781=>"000000101",
    2782=>"011111001",
    2783=>"111101011",
    2784=>"000001000",
    2785=>"000000000",
    2786=>"000011111",
    2787=>"100000000",
    2788=>"110100111",
    2789=>"000000011",
    2790=>"000000011",
    2791=>"100000000",
    2792=>"001001010",
    2793=>"000010111",
    2794=>"000100000",
    2795=>"110111110",
    2796=>"111110111",
    2797=>"001000111",
    2798=>"000000000",
    2799=>"111011100",
    2800=>"000000000",
    2801=>"001101111",
    2802=>"101111111",
    2803=>"000000000",
    2804=>"110000000",
    2805=>"101000110",
    2806=>"000001000",
    2807=>"111111110",
    2808=>"000000000",
    2809=>"111101010",
    2810=>"100000100",
    2811=>"000011111",
    2812=>"101010100",
    2813=>"100010100",
    2814=>"111111000",
    2815=>"000111010",
    2816=>"001001100",
    2817=>"011001100",
    2818=>"001000100",
    2819=>"111101000",
    2820=>"001011001",
    2821=>"011110000",
    2822=>"011011011",
    2823=>"011101000",
    2824=>"101001010",
    2825=>"000000001",
    2826=>"000001101",
    2827=>"100111111",
    2828=>"100110011",
    2829=>"100110011",
    2830=>"100111111",
    2831=>"111001100",
    2832=>"100110011",
    2833=>"011101100",
    2834=>"001001101",
    2835=>"011000100",
    2836=>"011001001",
    2837=>"010011000",
    2838=>"011001100",
    2839=>"100001110",
    2840=>"001001111",
    2841=>"110000010",
    2842=>"011001100",
    2843=>"000010001",
    2844=>"011111010",
    2845=>"111001011",
    2846=>"110111111",
    2847=>"011011110",
    2848=>"110101110",
    2849=>"110110011",
    2850=>"110011101",
    2851=>"000000100",
    2852=>"111000011",
    2853=>"110011110",
    2854=>"101111011",
    2855=>"011011011",
    2856=>"000001110",
    2857=>"000011000",
    2858=>"110100000",
    2859=>"010101101",
    2860=>"000100100",
    2861=>"000000001",
    2862=>"100010011",
    2863=>"110011000",
    2864=>"000100010",
    2865=>"001000000",
    2866=>"100110011",
    2867=>"001001011",
    2868=>"100100011",
    2869=>"100110011",
    2870=>"000100000",
    2871=>"010111101",
    2872=>"101011001",
    2873=>"100110110",
    2874=>"000001000",
    2875=>"100000000",
    2876=>"011001000",
    2877=>"000001001",
    2878=>"000000000",
    2879=>"111001001",
    2880=>"100110100",
    2881=>"000000000",
    2882=>"000000011",
    2883=>"001000100",
    2884=>"100110001",
    2885=>"011001001",
    2886=>"000010011",
    2887=>"110001000",
    2888=>"110100000",
    2889=>"101101010",
    2890=>"110000000",
    2891=>"000000100",
    2892=>"110000000",
    2893=>"111001101",
    2894=>"000100100",
    2895=>"011000100",
    2896=>"111101100",
    2897=>"001001101",
    2898=>"000000001",
    2899=>"011001011",
    2900=>"001001110",
    2901=>"001001010",
    2902=>"000000000",
    2903=>"101100000",
    2904=>"110111000",
    2905=>"100000001",
    2906=>"000101101",
    2907=>"000000000",
    2908=>"001000000",
    2909=>"001111011",
    2910=>"001101110",
    2911=>"010000110",
    2912=>"000000000",
    2913=>"001001010",
    2914=>"011001111",
    2915=>"111001001",
    2916=>"101100000",
    2917=>"001011110",
    2918=>"110010000",
    2919=>"101000001",
    2920=>"111000000",
    2921=>"000001000",
    2922=>"111001001",
    2923=>"010000000",
    2924=>"001001111",
    2925=>"011000100",
    2926=>"101111111",
    2927=>"000000001",
    2928=>"100100000",
    2929=>"011000110",
    2930=>"000000100",
    2931=>"100010000",
    2932=>"011001101",
    2933=>"011001000",
    2934=>"011100110",
    2935=>"111100000",
    2936=>"011001000",
    2937=>"011011101",
    2938=>"000110111",
    2939=>"110110110",
    2940=>"001011110",
    2941=>"111011000",
    2942=>"011011101",
    2943=>"001001001",
    2944=>"000010010",
    2945=>"111011000",
    2946=>"000000101",
    2947=>"000011101",
    2948=>"001001010",
    2949=>"111111000",
    2950=>"000000000",
    2951=>"000000010",
    2952=>"110011100",
    2953=>"001001000",
    2954=>"000100101",
    2955=>"011000100",
    2956=>"000010000",
    2957=>"111111010",
    2958=>"000011101",
    2959=>"110011011",
    2960=>"010010000",
    2961=>"111111001",
    2962=>"100011001",
    2963=>"000000011",
    2964=>"000001000",
    2965=>"100000010",
    2966=>"100000101",
    2967=>"000010111",
    2968=>"001110000",
    2969=>"110110000",
    2970=>"000100100",
    2971=>"000000100",
    2972=>"011111011",
    2973=>"000011001",
    2974=>"100011000",
    2975=>"000111011",
    2976=>"011100100",
    2977=>"011000000",
    2978=>"111111101",
    2979=>"000010011",
    2980=>"000000001",
    2981=>"010001000",
    2982=>"010010000",
    2983=>"000000101",
    2984=>"000000001",
    2985=>"111011010",
    2986=>"110000100",
    2987=>"000001000",
    2988=>"010111010",
    2989=>"010011010",
    2990=>"101000011",
    2991=>"010010000",
    2992=>"000000100",
    2993=>"001100101",
    2994=>"001100110",
    2995=>"000110100",
    2996=>"100111100",
    2997=>"011111000",
    2998=>"011111000",
    2999=>"011111000",
    3000=>"010000111",
    3001=>"001010111",
    3002=>"110110100",
    3003=>"111000000",
    3004=>"000000010",
    3005=>"101100101",
    3006=>"000000001",
    3007=>"111111000",
    3008=>"101101001",
    3009=>"000010011",
    3010=>"010010001",
    3011=>"000100101",
    3012=>"001111111",
    3013=>"001110101",
    3014=>"111000000",
    3015=>"010010000",
    3016=>"010111000",
    3017=>"000000000",
    3018=>"010000111",
    3019=>"001000001",
    3020=>"000000000",
    3021=>"000000111",
    3022=>"010010010",
    3023=>"100111000",
    3024=>"100000111",
    3025=>"100000111",
    3026=>"000111111",
    3027=>"000111011",
    3028=>"100001101",
    3029=>"000000000",
    3030=>"000010000",
    3031=>"000000111",
    3032=>"101110000",
    3033=>"000111010",
    3034=>"101000111",
    3035=>"101000000",
    3036=>"001001001",
    3037=>"110110110",
    3038=>"111101101",
    3039=>"011001111",
    3040=>"001111001",
    3041=>"001000101",
    3042=>"101010100",
    3043=>"111000100",
    3044=>"010010000",
    3045=>"000000101",
    3046=>"001100100",
    3047=>"010011010",
    3048=>"000010010",
    3049=>"000000001",
    3050=>"000101101",
    3051=>"111111111",
    3052=>"000000101",
    3053=>"010000011",
    3054=>"011111011",
    3055=>"000110010",
    3056=>"000000010",
    3057=>"101111111",
    3058=>"000000000",
    3059=>"010111000",
    3060=>"111101111",
    3061=>"000000000",
    3062=>"110000000",
    3063=>"000000000",
    3064=>"010111010",
    3065=>"000001010",
    3066=>"001010000",
    3067=>"010111010",
    3068=>"101111001",
    3069=>"011000111",
    3070=>"010100000",
    3071=>"110111001",
    3072=>"101100111",
    3073=>"010111111",
    3074=>"111000101",
    3075=>"000000000",
    3076=>"001000110",
    3077=>"000110111",
    3078=>"000100011",
    3079=>"101000000",
    3080=>"111111111",
    3081=>"111111110",
    3082=>"000000000",
    3083=>"100000110",
    3084=>"111111110",
    3085=>"000011000",
    3086=>"001011111",
    3087=>"111110000",
    3088=>"111111001",
    3089=>"110110010",
    3090=>"011111111",
    3091=>"100111111",
    3092=>"000000101",
    3093=>"011111111",
    3094=>"111000000",
    3095=>"001110110",
    3096=>"100011011",
    3097=>"100000001",
    3098=>"111111101",
    3099=>"010100000",
    3100=>"000010001",
    3101=>"010001001",
    3102=>"001111111",
    3103=>"100000000",
    3104=>"000000000",
    3105=>"000000000",
    3106=>"000000100",
    3107=>"000010110",
    3108=>"000000100",
    3109=>"000000110",
    3110=>"110011000",
    3111=>"011111111",
    3112=>"111110001",
    3113=>"111111111",
    3114=>"111111111",
    3115=>"001111111",
    3116=>"011011100",
    3117=>"000000000",
    3118=>"111111000",
    3119=>"001111111",
    3120=>"111111111",
    3121=>"111001000",
    3122=>"110110111",
    3123=>"100000001",
    3124=>"000101001",
    3125=>"000000000",
    3126=>"100010000",
    3127=>"000000010",
    3128=>"110101110",
    3129=>"000111111",
    3130=>"101111111",
    3131=>"000000100",
    3132=>"010111111",
    3133=>"000001111",
    3134=>"000001100",
    3135=>"100000111",
    3136=>"000110000",
    3137=>"001111000",
    3138=>"111110100",
    3139=>"000000000",
    3140=>"101000000",
    3141=>"100100100",
    3142=>"001011000",
    3143=>"010000111",
    3144=>"111111000",
    3145=>"000101101",
    3146=>"100110100",
    3147=>"010010000",
    3148=>"111111111",
    3149=>"111011000",
    3150=>"010010100",
    3151=>"011000000",
    3152=>"110000011",
    3153=>"100100111",
    3154=>"001000000",
    3155=>"111011111",
    3156=>"001101000",
    3157=>"001000000",
    3158=>"010100011",
    3159=>"001111111",
    3160=>"111010101",
    3161=>"110110001",
    3162=>"001011101",
    3163=>"000000000",
    3164=>"100111111",
    3165=>"111111111",
    3166=>"011111111",
    3167=>"010011100",
    3168=>"111111101",
    3169=>"001110100",
    3170=>"111111001",
    3171=>"000000111",
    3172=>"111110000",
    3173=>"010000000",
    3174=>"001000111",
    3175=>"111000000",
    3176=>"111111011",
    3177=>"000000111",
    3178=>"101111111",
    3179=>"011110101",
    3180=>"000101000",
    3181=>"001000111",
    3182=>"000000000",
    3183=>"101111111",
    3184=>"100000000",
    3185=>"111101101",
    3186=>"000000110",
    3187=>"111000111",
    3188=>"000000000",
    3189=>"000000000",
    3190=>"111111111",
    3191=>"100011111",
    3192=>"111000100",
    3193=>"000000110",
    3194=>"110111000",
    3195=>"111111000",
    3196=>"100100110",
    3197=>"111010111",
    3198=>"010000001",
    3199=>"101001001",
    3200=>"111111101",
    3201=>"101100101",
    3202=>"100100110",
    3203=>"111001000",
    3204=>"000001101",
    3205=>"011111000",
    3206=>"000111001",
    3207=>"000000111",
    3208=>"011111100",
    3209=>"111110100",
    3210=>"010001001",
    3211=>"011001001",
    3212=>"001000000",
    3213=>"110111110",
    3214=>"001011100",
    3215=>"110000111",
    3216=>"000100011",
    3217=>"101100111",
    3218=>"000000000",
    3219=>"110111111",
    3220=>"000001111",
    3221=>"011000000",
    3222=>"100000100",
    3223=>"000111011",
    3224=>"000100000",
    3225=>"110011100",
    3226=>"000111100",
    3227=>"001011111",
    3228=>"111001010",
    3229=>"001010000",
    3230=>"111101100",
    3231=>"011010010",
    3232=>"011000011",
    3233=>"000000001",
    3234=>"000110000",
    3235=>"000000101",
    3236=>"010010010",
    3237=>"100101100",
    3238=>"011111010",
    3239=>"101101000",
    3240=>"011010010",
    3241=>"000000000",
    3242=>"000110110",
    3243=>"100111101",
    3244=>"011000110",
    3245=>"010000000",
    3246=>"000000000",
    3247=>"111100000",
    3248=>"010001001",
    3249=>"001100111",
    3250=>"010110111",
    3251=>"100000000",
    3252=>"010000000",
    3253=>"000000000",
    3254=>"010111011",
    3255=>"111101101",
    3256=>"111000001",
    3257=>"000000010",
    3258=>"011001000",
    3259=>"100111101",
    3260=>"000111100",
    3261=>"010011000",
    3262=>"100110011",
    3263=>"011100101",
    3264=>"111001011",
    3265=>"000111011",
    3266=>"000000010",
    3267=>"111011011",
    3268=>"011110011",
    3269=>"100100101",
    3270=>"111111111",
    3271=>"100000000",
    3272=>"110001000",
    3273=>"100000000",
    3274=>"011000111",
    3275=>"000000000",
    3276=>"011011010",
    3277=>"000001111",
    3278=>"011010010",
    3279=>"100101001",
    3280=>"111011011",
    3281=>"100101001",
    3282=>"000000000",
    3283=>"011110110",
    3284=>"001000000",
    3285=>"100000101",
    3286=>"000011011",
    3287=>"000000001",
    3288=>"000100100",
    3289=>"111001000",
    3290=>"100101001",
    3291=>"011010101",
    3292=>"000010000",
    3293=>"011101110",
    3294=>"101001000",
    3295=>"010110110",
    3296=>"000111000",
    3297=>"000100110",
    3298=>"111001101",
    3299=>"010111010",
    3300=>"111010010",
    3301=>"000111010",
    3302=>"001100010",
    3303=>"111111010",
    3304=>"001000100",
    3305=>"101000100",
    3306=>"000101001",
    3307=>"111011111",
    3308=>"100100100",
    3309=>"000000000",
    3310=>"101110000",
    3311=>"010111000",
    3312=>"000000111",
    3313=>"011011010",
    3314=>"011000000",
    3315=>"010111000",
    3316=>"111101111",
    3317=>"100101100",
    3318=>"011111000",
    3319=>"110011111",
    3320=>"011000110",
    3321=>"100000011",
    3322=>"100000101",
    3323=>"111000111",
    3324=>"000110000",
    3325=>"000110011",
    3326=>"000010000",
    3327=>"110011000",
    3328=>"111110101",
    3329=>"101001001",
    3330=>"111111110",
    3331=>"111000011",
    3332=>"111011111",
    3333=>"011111111",
    3334=>"100101000",
    3335=>"111000000",
    3336=>"000111101",
    3337=>"011111111",
    3338=>"111001001",
    3339=>"011101101",
    3340=>"111000010",
    3341=>"000111111",
    3342=>"011011111",
    3343=>"000001011",
    3344=>"010111100",
    3345=>"001001001",
    3346=>"010000000",
    3347=>"111111001",
    3348=>"111001001",
    3349=>"000000100",
    3350=>"010100110",
    3351=>"110100111",
    3352=>"011000000",
    3353=>"111101110",
    3354=>"110001101",
    3355=>"111011011",
    3356=>"000000000",
    3357=>"001001000",
    3358=>"101000101",
    3359=>"110000000",
    3360=>"110100111",
    3361=>"110010110",
    3362=>"111101110",
    3363=>"110011001",
    3364=>"111111111",
    3365=>"101001001",
    3366=>"010110111",
    3367=>"101111111",
    3368=>"110001000",
    3369=>"001110111",
    3370=>"111000001",
    3371=>"001001111",
    3372=>"011001101",
    3373=>"011000000",
    3374=>"010000101",
    3375=>"001001001",
    3376=>"110110110",
    3377=>"010111110",
    3378=>"110000110",
    3379=>"001001011",
    3380=>"001101011",
    3381=>"101101111",
    3382=>"100000101",
    3383=>"000110110",
    3384=>"111000001",
    3385=>"001001000",
    3386=>"110111111",
    3387=>"101000001",
    3388=>"101000000",
    3389=>"000000000",
    3390=>"111100101",
    3391=>"001000000",
    3392=>"000000100",
    3393=>"110110011",
    3394=>"001000010",
    3395=>"000000000",
    3396=>"010100100",
    3397=>"110110110",
    3398=>"011111111",
    3399=>"000001101",
    3400=>"100111011",
    3401=>"110000000",
    3402=>"101110111",
    3403=>"001000000",
    3404=>"000111111",
    3405=>"110111000",
    3406=>"000000000",
    3407=>"000110110",
    3408=>"010010110",
    3409=>"000011010",
    3410=>"110110000",
    3411=>"001111111",
    3412=>"011011011",
    3413=>"101111010",
    3414=>"111000111",
    3415=>"001001000",
    3416=>"000100000",
    3417=>"111111111",
    3418=>"001001011",
    3419=>"111111110",
    3420=>"110111110",
    3421=>"010011100",
    3422=>"100101100",
    3423=>"001000100",
    3424=>"000111001",
    3425=>"100100100",
    3426=>"110111011",
    3427=>"000000000",
    3428=>"111111111",
    3429=>"011000000",
    3430=>"000000100",
    3431=>"010010000",
    3432=>"000000000",
    3433=>"001000000",
    3434=>"101001000",
    3435=>"101001110",
    3436=>"111101000",
    3437=>"110110111",
    3438=>"011000000",
    3439=>"101011111",
    3440=>"110000000",
    3441=>"000000000",
    3442=>"111110111",
    3443=>"000010000",
    3444=>"010010010",
    3445=>"000000000",
    3446=>"000111011",
    3447=>"110001011",
    3448=>"000000101",
    3449=>"111111000",
    3450=>"000000000",
    3451=>"000110111",
    3452=>"001101100",
    3453=>"000001111",
    3454=>"011001001",
    3455=>"001101001",
    3456=>"000111111",
    3457=>"111111111",
    3458=>"111111111",
    3459=>"001111110",
    3460=>"101001000",
    3461=>"000000000",
    3462=>"001111101",
    3463=>"000000111",
    3464=>"001011001",
    3465=>"111110010",
    3466=>"111011000",
    3467=>"111111110",
    3468=>"110111100",
    3469=>"110110110",
    3470=>"100001000",
    3471=>"000011111",
    3472=>"111011100",
    3473=>"110111111",
    3474=>"100110001",
    3475=>"000000000",
    3476=>"111111000",
    3477=>"001000000",
    3478=>"000000011",
    3479=>"001000000",
    3480=>"000101000",
    3481=>"111010001",
    3482=>"011100100",
    3483=>"011011111",
    3484=>"001000000",
    3485=>"111110000",
    3486=>"000000000",
    3487=>"000111111",
    3488=>"011101101",
    3489=>"111111111",
    3490=>"101110110",
    3491=>"011000011",
    3492=>"110111000",
    3493=>"001111000",
    3494=>"110111111",
    3495=>"001110000",
    3496=>"000000000",
    3497=>"100000001",
    3498=>"110001001",
    3499=>"100000101",
    3500=>"001000100",
    3501=>"011111000",
    3502=>"000000000",
    3503=>"000111111",
    3504=>"111101111",
    3505=>"000011100",
    3506=>"110111110",
    3507=>"000000000",
    3508=>"111111111",
    3509=>"111100000",
    3510=>"111111010",
    3511=>"000000000",
    3512=>"000001000",
    3513=>"001000000",
    3514=>"010010011",
    3515=>"010010010",
    3516=>"000000101",
    3517=>"101111111",
    3518=>"110111110",
    3519=>"111000100",
    3520=>"110111111",
    3521=>"110111111",
    3522=>"111111111",
    3523=>"111111111",
    3524=>"000111111",
    3525=>"011011000",
    3526=>"111100010",
    3527=>"111111111",
    3528=>"110111001",
    3529=>"111111111",
    3530=>"101000000",
    3531=>"111000000",
    3532=>"000000000",
    3533=>"101011010",
    3534=>"110100111",
    3535=>"110111111",
    3536=>"111011000",
    3537=>"000011001",
    3538=>"111000000",
    3539=>"000000000",
    3540=>"110010001",
    3541=>"110110000",
    3542=>"011000111",
    3543=>"000000000",
    3544=>"011001000",
    3545=>"111010001",
    3546=>"101111111",
    3547=>"000001011",
    3548=>"101100010",
    3549=>"001000000",
    3550=>"111111111",
    3551=>"000000000",
    3552=>"111100110",
    3553=>"100001000",
    3554=>"111111111",
    3555=>"000010000",
    3556=>"000000111",
    3557=>"001111101",
    3558=>"001111100",
    3559=>"001000001",
    3560=>"011111010",
    3561=>"100110011",
    3562=>"001000101",
    3563=>"000000000",
    3564=>"111111001",
    3565=>"000000000",
    3566=>"111111000",
    3567=>"000000000",
    3568=>"011011000",
    3569=>"111111111",
    3570=>"111110000",
    3571=>"101000000",
    3572=>"000111111",
    3573=>"101111000",
    3574=>"000000111",
    3575=>"111111111",
    3576=>"111000000",
    3577=>"111111111",
    3578=>"110111111",
    3579=>"111110110",
    3580=>"000100100",
    3581=>"101111111",
    3582=>"000000000",
    3583=>"000000011",
    3584=>"000001001",
    3585=>"111000101",
    3586=>"111111111",
    3587=>"000010010",
    3588=>"001000100",
    3589=>"100000100",
    3590=>"000110110",
    3591=>"010110110",
    3592=>"101011000",
    3593=>"111110100",
    3594=>"010110000",
    3595=>"010010000",
    3596=>"010111000",
    3597=>"110101000",
    3598=>"000000000",
    3599=>"110100011",
    3600=>"000011101",
    3601=>"000010000",
    3602=>"100111110",
    3603=>"100000000",
    3604=>"101000001",
    3605=>"110110000",
    3606=>"101000001",
    3607=>"110000000",
    3608=>"000111010",
    3609=>"110010010",
    3610=>"000011001",
    3611=>"001011011",
    3612=>"110001000",
    3613=>"010110111",
    3614=>"000011001",
    3615=>"110011111",
    3616=>"010111111",
    3617=>"000110100",
    3618=>"110111110",
    3619=>"000000111",
    3620=>"110010001",
    3621=>"000111111",
    3622=>"001010001",
    3623=>"000111110",
    3624=>"110010110",
    3625=>"000111000",
    3626=>"011100100",
    3627=>"000111011",
    3628=>"010011110",
    3629=>"000011111",
    3630=>"000000110",
    3631=>"000111111",
    3632=>"110111000",
    3633=>"001011010",
    3634=>"110111110",
    3635=>"000000010",
    3636=>"111111111",
    3637=>"110101010",
    3638=>"111000110",
    3639=>"111000111",
    3640=>"000000000",
    3641=>"100000000",
    3642=>"011011001",
    3643=>"100100100",
    3644=>"000110110",
    3645=>"000110110",
    3646=>"000100110",
    3647=>"010010101",
    3648=>"000011000",
    3649=>"000011001",
    3650=>"110110111",
    3651=>"111111010",
    3652=>"111111000",
    3653=>"000110001",
    3654=>"110101000",
    3655=>"111111111",
    3656=>"110110010",
    3657=>"000101101",
    3658=>"000000110",
    3659=>"000010000",
    3660=>"110110111",
    3661=>"000000000",
    3662=>"010110110",
    3663=>"000000000",
    3664=>"000000000",
    3665=>"100100110",
    3666=>"010010010",
    3667=>"111100000",
    3668=>"000010000",
    3669=>"101000100",
    3670=>"000000010",
    3671=>"001001011",
    3672=>"000111101",
    3673=>"111110000",
    3674=>"001111111",
    3675=>"001000000",
    3676=>"000110000",
    3677=>"011001100",
    3678=>"111011110",
    3679=>"011011111",
    3680=>"001101111",
    3681=>"000000000",
    3682=>"111100101",
    3683=>"101000010",
    3684=>"000000000",
    3685=>"010111010",
    3686=>"000011101",
    3687=>"110100011",
    3688=>"010011101",
    3689=>"000100110",
    3690=>"001111001",
    3691=>"010000000",
    3692=>"000000000",
    3693=>"100100001",
    3694=>"000000000",
    3695=>"100000100",
    3696=>"000101001",
    3697=>"111011011",
    3698=>"000111111",
    3699=>"100000000",
    3700=>"111001101",
    3701=>"010011000",
    3702=>"110010001",
    3703=>"111111010",
    3704=>"110011010",
    3705=>"111000000",
    3706=>"100000011",
    3707=>"111011111",
    3708=>"000111001",
    3709=>"111000000",
    3710=>"111110010",
    3711=>"010111011",
    3712=>"111101001",
    3713=>"000010010",
    3714=>"001000001",
    3715=>"011100000",
    3716=>"010001111",
    3717=>"111010100",
    3718=>"111110110",
    3719=>"101001000",
    3720=>"001100110",
    3721=>"101000101",
    3722=>"001001000",
    3723=>"001100110",
    3724=>"000101111",
    3725=>"010010010",
    3726=>"101111110",
    3727=>"110100000",
    3728=>"000000011",
    3729=>"111111010",
    3730=>"111001000",
    3731=>"100100110",
    3732=>"010010000",
    3733=>"111111111",
    3734=>"111000000",
    3735=>"000000000",
    3736=>"101001000",
    3737=>"000001011",
    3738=>"001001000",
    3739=>"101100000",
    3740=>"010111111",
    3741=>"001100110",
    3742=>"011001100",
    3743=>"001001000",
    3744=>"010101111",
    3745=>"100000001",
    3746=>"001101101",
    3747=>"111100111",
    3748=>"001111111",
    3749=>"010000010",
    3750=>"101100000",
    3751=>"000001111",
    3752=>"111111111",
    3753=>"000001001",
    3754=>"000001111",
    3755=>"111101001",
    3756=>"110000100",
    3757=>"111000000",
    3758=>"111111101",
    3759=>"011000000",
    3760=>"110010111",
    3761=>"101001000",
    3762=>"000110110",
    3763=>"111000111",
    3764=>"111100100",
    3765=>"001101101",
    3766=>"000000000",
    3767=>"111101001",
    3768=>"000000000",
    3769=>"110111101",
    3770=>"011000100",
    3771=>"000011001",
    3772=>"000000000",
    3773=>"011101101",
    3774=>"111010000",
    3775=>"111011111",
    3776=>"101110010",
    3777=>"101101111",
    3778=>"010010000",
    3779=>"010011111",
    3780=>"101101101",
    3781=>"110110110",
    3782=>"111000010",
    3783=>"000101111",
    3784=>"000100110",
    3785=>"010111111",
    3786=>"000000111",
    3787=>"101100000",
    3788=>"001101100",
    3789=>"010000000",
    3790=>"001001000",
    3791=>"111000000",
    3792=>"000000000",
    3793=>"100100110",
    3794=>"111110010",
    3795=>"000111101",
    3796=>"011011111",
    3797=>"000010000",
    3798=>"111111000",
    3799=>"111101001",
    3800=>"111100100",
    3801=>"111111001",
    3802=>"000001011",
    3803=>"110110100",
    3804=>"101001000",
    3805=>"011011011",
    3806=>"100000001",
    3807=>"111101001",
    3808=>"110001011",
    3809=>"001100100",
    3810=>"010010110",
    3811=>"001000001",
    3812=>"101001000",
    3813=>"001000101",
    3814=>"000001011",
    3815=>"111101010",
    3816=>"000011011",
    3817=>"101101001",
    3818=>"100001001",
    3819=>"010001000",
    3820=>"111111100",
    3821=>"111000101",
    3822=>"111110110",
    3823=>"110111011",
    3824=>"000001000",
    3825=>"011101101",
    3826=>"000010111",
    3827=>"000100100",
    3828=>"111011000",
    3829=>"000000010",
    3830=>"110111010",
    3831=>"000011011",
    3832=>"111000100",
    3833=>"011010111",
    3834=>"000111110",
    3835=>"000000000",
    3836=>"001000100",
    3837=>"100101111",
    3838=>"110000000",
    3839=>"110001000",
    3840=>"001000000",
    3841=>"000010000",
    3842=>"100000110",
    3843=>"000111111",
    3844=>"100010001",
    3845=>"000000011",
    3846=>"111100100",
    3847=>"000111110",
    3848=>"011100011",
    3849=>"000011011",
    3850=>"011111000",
    3851=>"100111111",
    3852=>"111000100",
    3853=>"101010110",
    3854=>"001110100",
    3855=>"001110100",
    3856=>"100000111",
    3857=>"111010000",
    3858=>"011000001",
    3859=>"001111100",
    3860=>"110000011",
    3861=>"110001000",
    3862=>"000110000",
    3863=>"001111111",
    3864=>"111000100",
    3865=>"011110100",
    3866=>"111000000",
    3867=>"100000000",
    3868=>"000100000",
    3869=>"001011100",
    3870=>"100110100",
    3871=>"000111111",
    3872=>"111111101",
    3873=>"000110100",
    3874=>"110000000",
    3875=>"001111100",
    3876=>"000011111",
    3877=>"110100000",
    3878=>"111111011",
    3879=>"111000000",
    3880=>"001111100",
    3881=>"001011010",
    3882=>"111000000",
    3883=>"011110100",
    3884=>"000111101",
    3885=>"000000111",
    3886=>"000111111",
    3887=>"111111000",
    3888=>"000011111",
    3889=>"111000011",
    3890=>"000101101",
    3891=>"000000111",
    3892=>"010001101",
    3893=>"000000111",
    3894=>"000001000",
    3895=>"111100111",
    3896=>"001110000",
    3897=>"000110000",
    3898=>"001011111",
    3899=>"111000000",
    3900=>"111011000",
    3901=>"100000011",
    3902=>"000000110",
    3903=>"010111010",
    3904=>"111000000",
    3905=>"111110000",
    3906=>"000111001",
    3907=>"000000100",
    3908=>"011100100",
    3909=>"000000011",
    3910=>"000010011",
    3911=>"001111011",
    3912=>"001010111",
    3913=>"111000111",
    3914=>"101111111",
    3915=>"110000000",
    3916=>"000101111",
    3917=>"010010001",
    3918=>"000111111",
    3919=>"111000111",
    3920=>"000000111",
    3921=>"011000110",
    3922=>"101000000",
    3923=>"101111000",
    3924=>"000000110",
    3925=>"100000111",
    3926=>"000000001",
    3927=>"000000111",
    3928=>"010110100",
    3929=>"100011100",
    3930=>"110000000",
    3931=>"110000011",
    3932=>"001110001",
    3933=>"110000011",
    3934=>"111000000",
    3935=>"011010000",
    3936=>"011001100",
    3937=>"000000111",
    3938=>"000011111",
    3939=>"000011000",
    3940=>"000111000",
    3941=>"000100111",
    3942=>"111000011",
    3943=>"000111100",
    3944=>"011110001",
    3945=>"111000000",
    3946=>"001111100",
    3947=>"000111000",
    3948=>"110000111",
    3949=>"000000111",
    3950=>"101000001",
    3951=>"110001001",
    3952=>"010000111",
    3953=>"100100000",
    3954=>"111101000",
    3955=>"111100010",
    3956=>"111100000",
    3957=>"110000000",
    3958=>"111000000",
    3959=>"010111101",
    3960=>"000111001",
    3961=>"000111110",
    3962=>"110000010",
    3963=>"000011000",
    3964=>"111000000",
    3965=>"000111000",
    3966=>"000000101",
    3967=>"001000100",
    3968=>"110001101",
    3969=>"000000101",
    3970=>"001101001",
    3971=>"111111111",
    3972=>"111100101",
    3973=>"010000000",
    3974=>"110000000",
    3975=>"001001101",
    3976=>"010100101",
    3977=>"100111001",
    3978=>"001101000",
    3979=>"011001000",
    3980=>"000000000",
    3981=>"111111110",
    3982=>"000001011",
    3983=>"100000101",
    3984=>"100110110",
    3985=>"001000000",
    3986=>"000100000",
    3987=>"000000000",
    3988=>"100100000",
    3989=>"111001111",
    3990=>"000000000",
    3991=>"000000110",
    3992=>"001001001",
    3993=>"100101001",
    3994=>"100100111",
    3995=>"111111111",
    3996=>"100000001",
    3997=>"101101011",
    3998=>"011011011",
    3999=>"000101000",
    4000=>"000001001",
    4001=>"111001000",
    4002=>"111001011",
    4003=>"010000000",
    4004=>"010010011",
    4005=>"010011010",
    4006=>"100110110",
    4007=>"110110010",
    4008=>"000100000",
    4009=>"100001010",
    4010=>"100001111",
    4011=>"111101101",
    4012=>"111000000",
    4013=>"011001000",
    4014=>"010010111",
    4015=>"101101100",
    4016=>"000000101",
    4017=>"000000101",
    4018=>"001001100",
    4019=>"000000000",
    4020=>"111011110",
    4021=>"001000000",
    4022=>"000000000",
    4023=>"101111111",
    4024=>"000000000",
    4025=>"110010000",
    4026=>"000111111",
    4027=>"000000000",
    4028=>"000000000",
    4029=>"111010000",
    4030=>"110011111",
    4031=>"111011010",
    4032=>"001111000",
    4033=>"010000010",
    4034=>"001000000",
    4035=>"000000000",
    4036=>"110111011",
    4037=>"111111111",
    4038=>"101111000",
    4039=>"000000011",
    4040=>"000011111",
    4041=>"111011010",
    4042=>"111011000",
    4043=>"000100111",
    4044=>"000000000",
    4045=>"111100100",
    4046=>"110010110",
    4047=>"000100111",
    4048=>"000000000",
    4049=>"100000001",
    4050=>"111000000",
    4051=>"011011011",
    4052=>"111011111",
    4053=>"000000000",
    4054=>"111000000",
    4055=>"000000000",
    4056=>"111111110",
    4057=>"000000001",
    4058=>"010100111",
    4059=>"000000000",
    4060=>"101101001",
    4061=>"000000100",
    4062=>"001100111",
    4063=>"001000000",
    4064=>"110011011",
    4065=>"001100100",
    4066=>"111000000",
    4067=>"001011010",
    4068=>"010000010",
    4069=>"001101000",
    4070=>"000000100",
    4071=>"000110111",
    4072=>"000000011",
    4073=>"101101101",
    4074=>"100100000",
    4075=>"000000001",
    4076=>"111101111",
    4077=>"000000000",
    4078=>"111110110",
    4079=>"001100100",
    4080=>"000000000",
    4081=>"110011111",
    4082=>"111111111",
    4083=>"000000110",
    4084=>"111111010",
    4085=>"000101101",
    4086=>"000000111",
    4087=>"000100001",
    4088=>"010000100",
    4089=>"000000000",
    4090=>"000000100",
    4091=>"000000101",
    4092=>"000000111",
    4093=>"101111111",
    4094=>"010010000",
    4095=>"111111111",
    4096=>"111110101",
    4097=>"010010011",
    4098=>"000000001",
    4099=>"100000101",
    4100=>"111011001",
    4101=>"000000000",
    4102=>"101101111",
    4103=>"111010111",
    4104=>"010011000",
    4105=>"010010000",
    4106=>"100001001",
    4107=>"111111011",
    4108=>"110111000",
    4109=>"110111000",
    4110=>"001000000",
    4111=>"100000111",
    4112=>"010110000",
    4113=>"000000000",
    4114=>"011010100",
    4115=>"110100101",
    4116=>"101001011",
    4117=>"010010001",
    4118=>"000000100",
    4119=>"000000000",
    4120=>"111111111",
    4121=>"111111010",
    4122=>"011001101",
    4123=>"100001101",
    4124=>"111111111",
    4125=>"011011011",
    4126=>"111011111",
    4127=>"000011101",
    4128=>"010111101",
    4129=>"011011110",
    4130=>"011111110",
    4131=>"000000000",
    4132=>"101101100",
    4133=>"111011111",
    4134=>"111000000",
    4135=>"101101000",
    4136=>"000000010",
    4137=>"000011110",
    4138=>"111011001",
    4139=>"111111001",
    4140=>"011001111",
    4141=>"111111101",
    4142=>"000000000",
    4143=>"111111011",
    4144=>"111101101",
    4145=>"011110010",
    4146=>"011111110",
    4147=>"101101001",
    4148=>"110111111",
    4149=>"000000010",
    4150=>"000011010",
    4151=>"000111111",
    4152=>"111111111",
    4153=>"111111111",
    4154=>"011010000",
    4155=>"111111111",
    4156=>"001000000",
    4157=>"001000000",
    4158=>"101111111",
    4159=>"100100101",
    4160=>"000100100",
    4161=>"000000000",
    4162=>"000110111",
    4163=>"000000000",
    4164=>"011100110",
    4165=>"100110001",
    4166=>"000001111",
    4167=>"111111101",
    4168=>"110010000",
    4169=>"000000000",
    4170=>"010111111",
    4171=>"000000000",
    4172=>"000110111",
    4173=>"111111000",
    4174=>"111111111",
    4175=>"010111110",
    4176=>"010011000",
    4177=>"101001001",
    4178=>"011000000",
    4179=>"100000000",
    4180=>"001001000",
    4181=>"000000000",
    4182=>"000011001",
    4183=>"101011111",
    4184=>"101111101",
    4185=>"111000100",
    4186=>"000000001",
    4187=>"011010000",
    4188=>"111111010",
    4189=>"001001101",
    4190=>"111011000",
    4191=>"000000001",
    4192=>"111110111",
    4193=>"011111110",
    4194=>"111111111",
    4195=>"000111111",
    4196=>"000000011",
    4197=>"010111000",
    4198=>"101100000",
    4199=>"111111101",
    4200=>"010010001",
    4201=>"011100011",
    4202=>"111111100",
    4203=>"000111100",
    4204=>"001000000",
    4205=>"000000000",
    4206=>"111001111",
    4207=>"000100110",
    4208=>"100100101",
    4209=>"000000000",
    4210=>"000101000",
    4211=>"010011000",
    4212=>"101000010",
    4213=>"000000000",
    4214=>"111010111",
    4215=>"110110000",
    4216=>"101111111",
    4217=>"111111000",
    4218=>"011111110",
    4219=>"111010001",
    4220=>"101101001",
    4221=>"000000000",
    4222=>"110111111",
    4223=>"111010010",
    4224=>"000011111",
    4225=>"101000101",
    4226=>"000111000",
    4227=>"110111001",
    4228=>"011011111",
    4229=>"111111101",
    4230=>"011111111",
    4231=>"001000111",
    4232=>"001001001",
    4233=>"011100100",
    4234=>"110010010",
    4235=>"011011000",
    4236=>"011000000",
    4237=>"111111101",
    4238=>"100000011",
    4239=>"000001011",
    4240=>"011111100",
    4241=>"010010111",
    4242=>"100110011",
    4243=>"110110001",
    4244=>"010011000",
    4245=>"101000000",
    4246=>"000000000",
    4247=>"011010010",
    4248=>"001111110",
    4249=>"110100000",
    4250=>"000101101",
    4251=>"111011011",
    4252=>"000000000",
    4253=>"000001000",
    4254=>"100001001",
    4255=>"000011110",
    4256=>"101100100",
    4257=>"111100101",
    4258=>"010001000",
    4259=>"111111110",
    4260=>"010010000",
    4261=>"110100100",
    4262=>"011000000",
    4263=>"001111111",
    4264=>"111111000",
    4265=>"100010111",
    4266=>"111111011",
    4267=>"000011001",
    4268=>"011111111",
    4269=>"000011010",
    4270=>"101000100",
    4271=>"111001101",
    4272=>"010011111",
    4273=>"100110111",
    4274=>"011100110",
    4275=>"000010000",
    4276=>"000100110",
    4277=>"000000000",
    4278=>"110111110",
    4279=>"110111001",
    4280=>"000111111",
    4281=>"010110111",
    4282=>"100001101",
    4283=>"000000000",
    4284=>"111000000",
    4285=>"000000101",
    4286=>"111111101",
    4287=>"111111010",
    4288=>"111011000",
    4289=>"111111111",
    4290=>"000111111",
    4291=>"000000000",
    4292=>"010111100",
    4293=>"010011011",
    4294=>"101111111",
    4295=>"111010000",
    4296=>"100100011",
    4297=>"000000000",
    4298=>"010010110",
    4299=>"100000100",
    4300=>"110111111",
    4301=>"000111010",
    4302=>"010111000",
    4303=>"101101000",
    4304=>"110010010",
    4305=>"111000111",
    4306=>"011111110",
    4307=>"100101111",
    4308=>"001010110",
    4309=>"000000000",
    4310=>"010010011",
    4311=>"110011111",
    4312=>"010110110",
    4313=>"111111000",
    4314=>"111011010",
    4315=>"000010101",
    4316=>"000110010",
    4317=>"001001100",
    4318=>"010100100",
    4319=>"111101000",
    4320=>"101101100",
    4321=>"000110100",
    4322=>"000111011",
    4323=>"010110110",
    4324=>"000010110",
    4325=>"000010010",
    4326=>"001100111",
    4327=>"111110000",
    4328=>"000000001",
    4329=>"111000001",
    4330=>"100111000",
    4331=>"100110111",
    4332=>"000000000",
    4333=>"010001000",
    4334=>"111111111",
    4335=>"000100100",
    4336=>"010111000",
    4337=>"001000010",
    4338=>"111111101",
    4339=>"000010010",
    4340=>"001000000",
    4341=>"000000000",
    4342=>"100000110",
    4343=>"100100011",
    4344=>"010010100",
    4345=>"111010011",
    4346=>"000000010",
    4347=>"111111111",
    4348=>"011111011",
    4349=>"111010010",
    4350=>"101111111",
    4351=>"100111001",
    4352=>"111111111",
    4353=>"110010000",
    4354=>"001001000",
    4355=>"011010000",
    4356=>"101001101",
    4357=>"111110111",
    4358=>"010101000",
    4359=>"000101101",
    4360=>"100101000",
    4361=>"001000000",
    4362=>"110011010",
    4363=>"011001100",
    4364=>"000011001",
    4365=>"111000011",
    4366=>"100001011",
    4367=>"000001111",
    4368=>"100100100",
    4369=>"111001000",
    4370=>"001111010",
    4371=>"000001101",
    4372=>"000000000",
    4373=>"000000101",
    4374=>"000000000",
    4375=>"100111111",
    4376=>"000001000",
    4377=>"111100000",
    4378=>"000100101",
    4379=>"000111011",
    4380=>"001001111",
    4381=>"000000111",
    4382=>"101001011",
    4383=>"111111011",
    4384=>"101010000",
    4385=>"111001111",
    4386=>"010101100",
    4387=>"000000100",
    4388=>"111111100",
    4389=>"000000001",
    4390=>"101000000",
    4391=>"111111101",
    4392=>"111000000",
    4393=>"110110100",
    4394=>"000000111",
    4395=>"100001000",
    4396=>"101110110",
    4397=>"000110010",
    4398=>"110000100",
    4399=>"101000000",
    4400=>"001101111",
    4401=>"111100100",
    4402=>"000010110",
    4403=>"000110010",
    4404=>"101101100",
    4405=>"010111110",
    4406=>"100100110",
    4407=>"010010010",
    4408=>"100000010",
    4409=>"111111111",
    4410=>"100000100",
    4411=>"010001000",
    4412=>"110000101",
    4413=>"101111111",
    4414=>"001011111",
    4415=>"000010111",
    4416=>"100000110",
    4417=>"010000000",
    4418=>"111000010",
    4419=>"000010101",
    4420=>"000000000",
    4421=>"001011110",
    4422=>"110110010",
    4423=>"111011110",
    4424=>"001001001",
    4425=>"111000111",
    4426=>"001111100",
    4427=>"000000100",
    4428=>"010011111",
    4429=>"111000000",
    4430=>"011000000",
    4431=>"001100000",
    4432=>"000000101",
    4433=>"000000001",
    4434=>"000000000",
    4435=>"111111011",
    4436=>"100110011",
    4437=>"010000000",
    4438=>"001010111",
    4439=>"111111111",
    4440=>"010011001",
    4441=>"000101110",
    4442=>"011111100",
    4443=>"001000101",
    4444=>"000000000",
    4445=>"100100100",
    4446=>"001000100",
    4447=>"000101111",
    4448=>"001000000",
    4449=>"000010100",
    4450=>"001000000",
    4451=>"000000000",
    4452=>"011000101",
    4453=>"001000101",
    4454=>"000000000",
    4455=>"000011011",
    4456=>"111001000",
    4457=>"111101001",
    4458=>"100110101",
    4459=>"000000110",
    4460=>"101101001",
    4461=>"111000111",
    4462=>"111110010",
    4463=>"001101110",
    4464=>"110010000",
    4465=>"101001001",
    4466=>"011101000",
    4467=>"111001000",
    4468=>"000000110",
    4469=>"000111000",
    4470=>"000000000",
    4471=>"100000011",
    4472=>"000010011",
    4473=>"010000110",
    4474=>"010000000",
    4475=>"000101101",
    4476=>"110101000",
    4477=>"000010011",
    4478=>"101010000",
    4479=>"111111001",
    4480=>"000000101",
    4481=>"000000010",
    4482=>"000100000",
    4483=>"000000001",
    4484=>"100100110",
    4485=>"000000000",
    4486=>"000100001",
    4487=>"111001001",
    4488=>"001001001",
    4489=>"010000100",
    4490=>"100001001",
    4491=>"000000000",
    4492=>"000000000",
    4493=>"111111110",
    4494=>"000011000",
    4495=>"000000000",
    4496=>"001111011",
    4497=>"111101101",
    4498=>"111110111",
    4499=>"001011111",
    4500=>"000000100",
    4501=>"010011000",
    4502=>"000010000",
    4503=>"110111010",
    4504=>"000111110",
    4505=>"000000000",
    4506=>"011100111",
    4507=>"011111110",
    4508=>"011001001",
    4509=>"111111100",
    4510=>"000111111",
    4511=>"000000110",
    4512=>"100101111",
    4513=>"100100100",
    4514=>"001100000",
    4515=>"000000001",
    4516=>"111111000",
    4517=>"001000000",
    4518=>"100100011",
    4519=>"101111011",
    4520=>"101111111",
    4521=>"110100000",
    4522=>"100101001",
    4523=>"001100000",
    4524=>"110011001",
    4525=>"101111010",
    4526=>"100000011",
    4527=>"110110010",
    4528=>"001000000",
    4529=>"010000000",
    4530=>"000111011",
    4531=>"011011111",
    4532=>"001001001",
    4533=>"110101000",
    4534=>"000000000",
    4535=>"010111100",
    4536=>"111111100",
    4537=>"110111111",
    4538=>"000000011",
    4539=>"011000111",
    4540=>"000000000",
    4541=>"000000001",
    4542=>"110111111",
    4543=>"111111010",
    4544=>"000001101",
    4545=>"000000000",
    4546=>"011011010",
    4547=>"000000000",
    4548=>"000000011",
    4549=>"000000000",
    4550=>"111110000",
    4551=>"100000110",
    4552=>"110001111",
    4553=>"101101100",
    4554=>"010000000",
    4555=>"111000100",
    4556=>"000000000",
    4557=>"000001000",
    4558=>"111111111",
    4559=>"110000000",
    4560=>"000110110",
    4561=>"011001011",
    4562=>"100111111",
    4563=>"100011010",
    4564=>"000000000",
    4565=>"010000000",
    4566=>"011011101",
    4567=>"110111101",
    4568=>"111011011",
    4569=>"000001111",
    4570=>"000001101",
    4571=>"011111111",
    4572=>"000000000",
    4573=>"011100010",
    4574=>"000000101",
    4575=>"111111111",
    4576=>"100000000",
    4577=>"100110110",
    4578=>"000000001",
    4579=>"000000000",
    4580=>"000000001",
    4581=>"010111011",
    4582=>"100000101",
    4583=>"010110000",
    4584=>"000000001",
    4585=>"000000100",
    4586=>"010011100",
    4587=>"110011111",
    4588=>"111111111",
    4589=>"100000000",
    4590=>"000000000",
    4591=>"000110100",
    4592=>"111110111",
    4593=>"111111111",
    4594=>"101101111",
    4595=>"000000001",
    4596=>"000000000",
    4597=>"001000001",
    4598=>"101111110",
    4599=>"000011110",
    4600=>"111111011",
    4601=>"100000000",
    4602=>"000000000",
    4603=>"111110111",
    4604=>"000100110",
    4605=>"000000000",
    4606=>"111111111",
    4607=>"000000100",
    4608=>"000000010",
    4609=>"001011001",
    4610=>"110110110",
    4611=>"000001001",
    4612=>"100000100",
    4613=>"001001010",
    4614=>"000011010",
    4615=>"100100101",
    4616=>"000000000",
    4617=>"010110100",
    4618=>"111100000",
    4619=>"010011100",
    4620=>"000001000",
    4621=>"001011000",
    4622=>"010001001",
    4623=>"110101010",
    4624=>"100110110",
    4625=>"110100100",
    4626=>"000000001",
    4627=>"100100100",
    4628=>"100100100",
    4629=>"100000000",
    4630=>"110010010",
    4631=>"100101011",
    4632=>"101111111",
    4633=>"000101010",
    4634=>"000100101",
    4635=>"100001101",
    4636=>"011110111",
    4637=>"000000000",
    4638=>"000000000",
    4639=>"100100001",
    4640=>"011101000",
    4641=>"001010101",
    4642=>"101100100",
    4643=>"010011001",
    4644=>"001000000",
    4645=>"000100000",
    4646=>"000011001",
    4647=>"100100100",
    4648=>"110011100",
    4649=>"011001011",
    4650=>"101100011",
    4651=>"111111111",
    4652=>"000001001",
    4653=>"001011011",
    4654=>"100000001",
    4655=>"110111001",
    4656=>"000000100",
    4657=>"000110100",
    4658=>"001111111",
    4659=>"010011010",
    4660=>"111111101",
    4661=>"011011011",
    4662=>"001011001",
    4663=>"011011000",
    4664=>"110100000",
    4665=>"100101011",
    4666=>"100110110",
    4667=>"000000011",
    4668=>"111111100",
    4669=>"100100000",
    4670=>"100111011",
    4671=>"100111011",
    4672=>"110110110",
    4673=>"100110110",
    4674=>"000011111",
    4675=>"000001110",
    4676=>"110110100",
    4677=>"001001001",
    4678=>"010110010",
    4679=>"111011010",
    4680=>"010111100",
    4681=>"000011001",
    4682=>"000000000",
    4683=>"011000000",
    4684=>"110110110",
    4685=>"100100110",
    4686=>"110001100",
    4687=>"001011001",
    4688=>"001100100",
    4689=>"010000000",
    4690=>"000001001",
    4691=>"100011010",
    4692=>"101101110",
    4693=>"010100011",
    4694=>"110000001",
    4695=>"111000101",
    4696=>"001011011",
    4697=>"000100110",
    4698=>"111010111",
    4699=>"010100100",
    4700=>"000000000",
    4701=>"001000001",
    4702=>"101000110",
    4703=>"100011010",
    4704=>"000111110",
    4705=>"100100111",
    4706=>"100100110",
    4707=>"110100110",
    4708=>"100100110",
    4709=>"010000000",
    4710=>"100100011",
    4711=>"001011011",
    4712=>"000011000",
    4713=>"111100000",
    4714=>"111111111",
    4715=>"111110001",
    4716=>"100100100",
    4717=>"001111000",
    4718=>"000100001",
    4719=>"001101111",
    4720=>"010110011",
    4721=>"001111111",
    4722=>"010110110",
    4723=>"001011001",
    4724=>"011111111",
    4725=>"101000001",
    4726=>"111011111",
    4727=>"110110010",
    4728=>"111111111",
    4729=>"011111101",
    4730=>"010001001",
    4731=>"000011001",
    4732=>"011000100",
    4733=>"001011010",
    4734=>"001001001",
    4735=>"010111111",
    4736=>"101000110",
    4737=>"111001000",
    4738=>"100100100",
    4739=>"000111001",
    4740=>"001000111",
    4741=>"110111100",
    4742=>"000110110",
    4743=>"101011000",
    4744=>"110100100",
    4745=>"111110101",
    4746=>"011100000",
    4747=>"100110110",
    4748=>"100110010",
    4749=>"011111011",
    4750=>"110100100",
    4751=>"011011001",
    4752=>"111100110",
    4753=>"011001011",
    4754=>"001101001",
    4755=>"110110101",
    4756=>"000000011",
    4757=>"100111010",
    4758=>"100000000",
    4759=>"011001011",
    4760=>"000110101",
    4761=>"110111000",
    4762=>"001000100",
    4763=>"000001000",
    4764=>"011111110",
    4765=>"000101001",
    4766=>"000000100",
    4767=>"000001011",
    4768=>"000110110",
    4769=>"100111110",
    4770=>"101000001",
    4771=>"010010011",
    4772=>"000110110",
    4773=>"100001011",
    4774=>"010111011",
    4775=>"100100110",
    4776=>"011000001",
    4777=>"111100001",
    4778=>"000000011",
    4779=>"000110100",
    4780=>"001001110",
    4781=>"010011011",
    4782=>"011111111",
    4783=>"111101000",
    4784=>"000011000",
    4785=>"110111000",
    4786=>"000100010",
    4787=>"110110111",
    4788=>"011100100",
    4789=>"000000100",
    4790=>"011011000",
    4791=>"110100111",
    4792=>"001011111",
    4793=>"011100100",
    4794=>"010100000",
    4795=>"101001000",
    4796=>"011001001",
    4797=>"000000000",
    4798=>"011111111",
    4799=>"111011001",
    4800=>"110111100",
    4801=>"000000101",
    4802=>"011000000",
    4803=>"100111110",
    4804=>"110110000",
    4805=>"000111111",
    4806=>"000101101",
    4807=>"011111001",
    4808=>"000110110",
    4809=>"000000101",
    4810=>"001000000",
    4811=>"000001011",
    4812=>"110111010",
    4813=>"000000111",
    4814=>"100001011",
    4815=>"100100100",
    4816=>"000000010",
    4817=>"000110110",
    4818=>"001100100",
    4819=>"111001100",
    4820=>"000010110",
    4821=>"100011010",
    4822=>"000100100",
    4823=>"100100100",
    4824=>"100110111",
    4825=>"111110000",
    4826=>"000000111",
    4827=>"100000000",
    4828=>"010110101",
    4829=>"100001000",
    4830=>"001000010",
    4831=>"100000101",
    4832=>"001111111",
    4833=>"000011111",
    4834=>"011110111",
    4835=>"110111011",
    4836=>"011111011",
    4837=>"000101000",
    4838=>"111000011",
    4839=>"001001001",
    4840=>"011011001",
    4841=>"011100100",
    4842=>"000110101",
    4843=>"010011111",
    4844=>"100000110",
    4845=>"000000001",
    4846=>"111110100",
    4847=>"000000001",
    4848=>"110110010",
    4849=>"100000010",
    4850=>"001010110",
    4851=>"110110010",
    4852=>"111100101",
    4853=>"000000010",
    4854=>"101011101",
    4855=>"111010010",
    4856=>"011000011",
    4857=>"001001011",
    4858=>"000101111",
    4859=>"011001101",
    4860=>"111001101",
    4861=>"011101001",
    4862=>"000000000",
    4863=>"000110111",
    4864=>"111011011",
    4865=>"011110111",
    4866=>"111111100",
    4867=>"001001101",
    4868=>"011001001",
    4869=>"010011000",
    4870=>"111101101",
    4871=>"000000000",
    4872=>"000000001",
    4873=>"101001000",
    4874=>"000000000",
    4875=>"011000000",
    4876=>"011000101",
    4877=>"110110110",
    4878=>"001111101",
    4879=>"111001001",
    4880=>"110110111",
    4881=>"111111111",
    4882=>"100000000",
    4883=>"110100000",
    4884=>"111000000",
    4885=>"000000000",
    4886=>"111000000",
    4887=>"010010010",
    4888=>"000100001",
    4889=>"110010101",
    4890=>"001101011",
    4891=>"011110110",
    4892=>"111110000",
    4893=>"100100100",
    4894=>"000011110",
    4895=>"000000111",
    4896=>"011000000",
    4897=>"111011111",
    4898=>"001010001",
    4899=>"111111111",
    4900=>"010110010",
    4901=>"111000001",
    4902=>"000100110",
    4903=>"111011000",
    4904=>"011101100",
    4905=>"111011111",
    4906=>"000010011",
    4907=>"000001001",
    4908=>"000000000",
    4909=>"001111100",
    4910=>"111011110",
    4911=>"110111111",
    4912=>"010011101",
    4913=>"111111111",
    4914=>"111100010",
    4915=>"011101001",
    4916=>"000100000",
    4917=>"000000110",
    4918=>"111110010",
    4919=>"000111111",
    4920=>"010010000",
    4921=>"000000000",
    4922=>"111010000",
    4923=>"101111110",
    4924=>"101000001",
    4925=>"111010111",
    4926=>"100110001",
    4927=>"000000000",
    4928=>"000000000",
    4929=>"100111110",
    4930=>"000000111",
    4931=>"111011010",
    4932=>"111010110",
    4933=>"101111111",
    4934=>"111101111",
    4935=>"010011000",
    4936=>"001001001",
    4937=>"000111001",
    4938=>"001000100",
    4939=>"111000000",
    4940=>"110010100",
    4941=>"110111111",
    4942=>"000000000",
    4943=>"010111110",
    4944=>"111101110",
    4945=>"101001000",
    4946=>"111010111",
    4947=>"000101111",
    4948=>"111111111",
    4949=>"011011001",
    4950=>"111111010",
    4951=>"111110010",
    4952=>"101110101",
    4953=>"000000000",
    4954=>"010111101",
    4955=>"110111111",
    4956=>"000101101",
    4957=>"011000000",
    4958=>"000001011",
    4959=>"000100000",
    4960=>"000101111",
    4961=>"001101101",
    4962=>"111111110",
    4963=>"100000000",
    4964=>"000110111",
    4965=>"111011100",
    4966=>"111000100",
    4967=>"000000000",
    4968=>"111111011",
    4969=>"100000110",
    4970=>"000001000",
    4971=>"010110011",
    4972=>"111110000",
    4973=>"111101101",
    4974=>"111000000",
    4975=>"101111111",
    4976=>"111001000",
    4977=>"100010000",
    4978=>"000010111",
    4979=>"001101000",
    4980=>"001000111",
    4981=>"000000000",
    4982=>"111111111",
    4983=>"100111100",
    4984=>"010000000",
    4985=>"011000111",
    4986=>"110010110",
    4987=>"000100000",
    4988=>"100110111",
    4989=>"110111010",
    4990=>"111100000",
    4991=>"010110000",
    4992=>"000000000",
    4993=>"111000000",
    4994=>"000000111",
    4995=>"111111111",
    4996=>"011011101",
    4997=>"010011101",
    4998=>"111001101",
    4999=>"101000000",
    5000=>"011000000",
    5001=>"110110111",
    5002=>"110101100",
    5003=>"111101010",
    5004=>"101111111",
    5005=>"110110010",
    5006=>"000010011",
    5007=>"100001001",
    5008=>"001100010",
    5009=>"000101011",
    5010=>"110000100",
    5011=>"111100111",
    5012=>"000001000",
    5013=>"010000000",
    5014=>"000000000",
    5015=>"111111111",
    5016=>"001100000",
    5017=>"111101110",
    5018=>"110100001",
    5019=>"010110111",
    5020=>"010000000",
    5021=>"000011000",
    5022=>"010001000",
    5023=>"000010010",
    5024=>"000000111",
    5025=>"000001100",
    5026=>"101000000",
    5027=>"100000001",
    5028=>"000011111",
    5029=>"000000000",
    5030=>"000111111",
    5031=>"100101000",
    5032=>"000000101",
    5033=>"111100000",
    5034=>"000001111",
    5035=>"100001001",
    5036=>"110110000",
    5037=>"111111000",
    5038=>"000000001",
    5039=>"111000111",
    5040=>"001000111",
    5041=>"111000010",
    5042=>"000100110",
    5043=>"010000001",
    5044=>"110110110",
    5045=>"011000000",
    5046=>"011111000",
    5047=>"000111000",
    5048=>"001011011",
    5049=>"000011111",
    5050=>"111011101",
    5051=>"000000000",
    5052=>"111000101",
    5053=>"111001111",
    5054=>"001011000",
    5055=>"111110000",
    5056=>"111111010",
    5057=>"101000110",
    5058=>"011111111",
    5059=>"010000001",
    5060=>"000001100",
    5061=>"001010100",
    5062=>"111111000",
    5063=>"111101000",
    5064=>"110001000",
    5065=>"000111110",
    5066=>"000000110",
    5067=>"000000001",
    5068=>"101001110",
    5069=>"100000111",
    5070=>"100111001",
    5071=>"000000111",
    5072=>"000010010",
    5073=>"011010000",
    5074=>"000111011",
    5075=>"000100111",
    5076=>"100000001",
    5077=>"111111011",
    5078=>"000011101",
    5079=>"101111010",
    5080=>"111111000",
    5081=>"000000100",
    5082=>"110100110",
    5083=>"000000000",
    5084=>"000100000",
    5085=>"001100111",
    5086=>"000100110",
    5087=>"000000010",
    5088=>"000100111",
    5089=>"110100111",
    5090=>"000000000",
    5091=>"011000000",
    5092=>"101111111",
    5093=>"000000000",
    5094=>"110110100",
    5095=>"011111111",
    5096=>"100001000",
    5097=>"111000101",
    5098=>"110001001",
    5099=>"011111000",
    5100=>"111000101",
    5101=>"000001000",
    5102=>"100111100",
    5103=>"000000100",
    5104=>"010000000",
    5105=>"000010111",
    5106=>"100000000",
    5107=>"010111111",
    5108=>"101001000",
    5109=>"000001111",
    5110=>"000000111",
    5111=>"000001011",
    5112=>"110010000",
    5113=>"111000111",
    5114=>"000000000",
    5115=>"011000111",
    5116=>"000000000",
    5117=>"111100111",
    5118=>"111111101",
    5119=>"110111000",
    5120=>"000000000",
    5121=>"010000111",
    5122=>"000111110",
    5123=>"000000000",
    5124=>"011001000",
    5125=>"010111111",
    5126=>"111110010",
    5127=>"100000110",
    5128=>"000111011",
    5129=>"010110000",
    5130=>"101000000",
    5131=>"000111100",
    5132=>"001000000",
    5133=>"110111110",
    5134=>"001101011",
    5135=>"000010011",
    5136=>"000111100",
    5137=>"101000000",
    5138=>"001000001",
    5139=>"110010000",
    5140=>"101000001",
    5141=>"100000000",
    5142=>"000000000",
    5143=>"011000110",
    5144=>"111001110",
    5145=>"010110000",
    5146=>"101101100",
    5147=>"011001011",
    5148=>"001011111",
    5149=>"011111001",
    5150=>"110110111",
    5151=>"000000000",
    5152=>"110100111",
    5153=>"111110111",
    5154=>"011101110",
    5155=>"100111110",
    5156=>"011001011",
    5157=>"111001001",
    5158=>"000000000",
    5159=>"000111011",
    5160=>"111000000",
    5161=>"000001011",
    5162=>"001001010",
    5163=>"011011011",
    5164=>"011001001",
    5165=>"111011001",
    5166=>"000000011",
    5167=>"000000000",
    5168=>"111011010",
    5169=>"000000000",
    5170=>"110111110",
    5171=>"000000110",
    5172=>"100100100",
    5173=>"001000010",
    5174=>"010110010",
    5175=>"000010000",
    5176=>"000000000",
    5177=>"111111110",
    5178=>"000011001",
    5179=>"000000001",
    5180=>"101000000",
    5181=>"101000101",
    5182=>"100100110",
    5183=>"111000100",
    5184=>"000110100",
    5185=>"000000011",
    5186=>"000000000",
    5187=>"101011000",
    5188=>"010110111",
    5189=>"001011001",
    5190=>"110111111",
    5191=>"100001000",
    5192=>"000110001",
    5193=>"111010010",
    5194=>"000110110",
    5195=>"000000000",
    5196=>"000111010",
    5197=>"011111011",
    5198=>"000000000",
    5199=>"000010010",
    5200=>"110011010",
    5201=>"000000000",
    5202=>"100000000",
    5203=>"110100110",
    5204=>"011110110",
    5205=>"100010010",
    5206=>"010011011",
    5207=>"110111011",
    5208=>"001100110",
    5209=>"111111010",
    5210=>"011001011",
    5211=>"000010000",
    5212=>"110100100",
    5213=>"000000100",
    5214=>"001001001",
    5215=>"101000010",
    5216=>"001001011",
    5217=>"100100011",
    5218=>"010011010",
    5219=>"010000000",
    5220=>"000111111",
    5221=>"000000000",
    5222=>"001000000",
    5223=>"011110000",
    5224=>"000011101",
    5225=>"101100000",
    5226=>"100100011",
    5227=>"111111110",
    5228=>"101000111",
    5229=>"010000000",
    5230=>"111000000",
    5231=>"100001110",
    5232=>"000000000",
    5233=>"000000010",
    5234=>"000000000",
    5235=>"010111111",
    5236=>"111001100",
    5237=>"000000101",
    5238=>"000001111",
    5239=>"100111011",
    5240=>"000001000",
    5241=>"111000000",
    5242=>"111000110",
    5243=>"110000111",
    5244=>"100110110",
    5245=>"001010110",
    5246=>"111001000",
    5247=>"111111011",
    5248=>"111101100",
    5249=>"101100111",
    5250=>"011011000",
    5251=>"111111110",
    5252=>"000000000",
    5253=>"111100111",
    5254=>"111111101",
    5255=>"000000000",
    5256=>"011001101",
    5257=>"110110010",
    5258=>"111000000",
    5259=>"111100101",
    5260=>"001100111",
    5261=>"100101111",
    5262=>"111100001",
    5263=>"100000011",
    5264=>"001100000",
    5265=>"000010000",
    5266=>"011011000",
    5267=>"110100000",
    5268=>"001000000",
    5269=>"000000000",
    5270=>"101001101",
    5271=>"000111111",
    5272=>"011110000",
    5273=>"111001111",
    5274=>"101101010",
    5275=>"000011001",
    5276=>"111111101",
    5277=>"111111001",
    5278=>"110111011",
    5279=>"000010010",
    5280=>"111001000",
    5281=>"111110010",
    5282=>"001101010",
    5283=>"000111011",
    5284=>"011011000",
    5285=>"000000000",
    5286=>"000010111",
    5287=>"011111000",
    5288=>"011000000",
    5289=>"001011011",
    5290=>"011000000",
    5291=>"000011000",
    5292=>"000110111",
    5293=>"010011010",
    5294=>"000110010",
    5295=>"111111001",
    5296=>"010010000",
    5297=>"010010000",
    5298=>"010100100",
    5299=>"000011000",
    5300=>"001101110",
    5301=>"000001011",
    5302=>"111100111",
    5303=>"000000000",
    5304=>"000100111",
    5305=>"010110011",
    5306=>"011000100",
    5307=>"101100111",
    5308=>"100100111",
    5309=>"010011000",
    5310=>"100111100",
    5311=>"100000100",
    5312=>"100100111",
    5313=>"000110000",
    5314=>"000101000",
    5315=>"100000110",
    5316=>"111011000",
    5317=>"011011000",
    5318=>"101101110",
    5319=>"111111111",
    5320=>"100000000",
    5321=>"101000101",
    5322=>"000110011",
    5323=>"000000101",
    5324=>"111000000",
    5325=>"010011000",
    5326=>"111111000",
    5327=>"100000100",
    5328=>"011010010",
    5329=>"000000001",
    5330=>"100100111",
    5331=>"111000100",
    5332=>"110110000",
    5333=>"001001101",
    5334=>"100000001",
    5335=>"111101000",
    5336=>"111100100",
    5337=>"111111010",
    5338=>"000001110",
    5339=>"101000000",
    5340=>"110110000",
    5341=>"001000100",
    5342=>"100110100",
    5343=>"100000101",
    5344=>"000010001",
    5345=>"100010000",
    5346=>"110011000",
    5347=>"000000000",
    5348=>"111110011",
    5349=>"010010001",
    5350=>"001100110",
    5351=>"110100101",
    5352=>"100000010",
    5353=>"101100101",
    5354=>"111111000",
    5355=>"111000010",
    5356=>"100000000",
    5357=>"101101100",
    5358=>"001000011",
    5359=>"010000100",
    5360=>"010110101",
    5361=>"100101111",
    5362=>"101101111",
    5363=>"101000111",
    5364=>"101100111",
    5365=>"000000100",
    5366=>"000000000",
    5367=>"010001111",
    5368=>"111000100",
    5369=>"110100111",
    5370=>"101000001",
    5371=>"111000001",
    5372=>"000100001",
    5373=>"011000100",
    5374=>"111111000",
    5375=>"000111111",
    5376=>"000000000",
    5377=>"000111010",
    5378=>"001000000",
    5379=>"011111111",
    5380=>"000111000",
    5381=>"111111111",
    5382=>"000000000",
    5383=>"000111100",
    5384=>"011111011",
    5385=>"111011010",
    5386=>"010101011",
    5387=>"011001000",
    5388=>"010010000",
    5389=>"110111010",
    5390=>"110111011",
    5391=>"110000000",
    5392=>"011001000",
    5393=>"100111101",
    5394=>"010000011",
    5395=>"000100010",
    5396=>"011111000",
    5397=>"000000000",
    5398=>"111011101",
    5399=>"011000111",
    5400=>"000110110",
    5401=>"110000000",
    5402=>"001111010",
    5403=>"000100110",
    5404=>"011111111",
    5405=>"111111000",
    5406=>"110111101",
    5407=>"000111111",
    5408=>"011000000",
    5409=>"110111010",
    5410=>"011000100",
    5411=>"010000010",
    5412=>"111111000",
    5413=>"110000100",
    5414=>"111111111",
    5415=>"001001001",
    5416=>"111000001",
    5417=>"110110111",
    5418=>"011001000",
    5419=>"110101011",
    5420=>"111111011",
    5421=>"000111111",
    5422=>"111111011",
    5423=>"111111111",
    5424=>"111000111",
    5425=>"011000001",
    5426=>"110000110",
    5427=>"001011111",
    5428=>"011111010",
    5429=>"111111000",
    5430=>"111111000",
    5431=>"000111000",
    5432=>"111101001",
    5433=>"110100111",
    5434=>"111110110",
    5435=>"111000001",
    5436=>"000000001",
    5437=>"000000000",
    5438=>"000000101",
    5439=>"011011000",
    5440=>"000100000",
    5441=>"111101000",
    5442=>"111101111",
    5443=>"000111111",
    5444=>"111111011",
    5445=>"001000100",
    5446=>"011111101",
    5447=>"110000000",
    5448=>"110000010",
    5449=>"000000101",
    5450=>"111000110",
    5451=>"111010111",
    5452=>"111111101",
    5453=>"111001101",
    5454=>"111111111",
    5455=>"001111111",
    5456=>"000111110",
    5457=>"111000100",
    5458=>"100101111",
    5459=>"100101101",
    5460=>"000000000",
    5461=>"000000001",
    5462=>"000000001",
    5463=>"111111111",
    5464=>"001000000",
    5465=>"100000110",
    5466=>"100110111",
    5467=>"000000000",
    5468=>"000001010",
    5469=>"001001010",
    5470=>"110111111",
    5471=>"000000000",
    5472=>"100111101",
    5473=>"110010001",
    5474=>"000000111",
    5475=>"111101000",
    5476=>"111010101",
    5477=>"001010000",
    5478=>"010000001",
    5479=>"000001111",
    5480=>"000111111",
    5481=>"000000000",
    5482=>"000000011",
    5483=>"111111011",
    5484=>"000000000",
    5485=>"101101101",
    5486=>"010111110",
    5487=>"000100100",
    5488=>"000000000",
    5489=>"000100010",
    5490=>"100000111",
    5491=>"111001001",
    5492=>"000000000",
    5493=>"100100001",
    5494=>"010000000",
    5495=>"110001011",
    5496=>"111111111",
    5497=>"111000010",
    5498=>"100111011",
    5499=>"011111110",
    5500=>"000111011",
    5501=>"111000001",
    5502=>"111101101",
    5503=>"110111111",
    5504=>"111111101",
    5505=>"101100101",
    5506=>"101000100",
    5507=>"011011000",
    5508=>"010110010",
    5509=>"000010000",
    5510=>"101101101",
    5511=>"011011111",
    5512=>"011000010",
    5513=>"110110000",
    5514=>"000110111",
    5515=>"000000110",
    5516=>"110101000",
    5517=>"110000100",
    5518=>"111111111",
    5519=>"110001011",
    5520=>"001100111",
    5521=>"000000000",
    5522=>"010011010",
    5523=>"000011011",
    5524=>"000000001",
    5525=>"111010000",
    5526=>"000000110",
    5527=>"000011110",
    5528=>"010110000",
    5529=>"000011010",
    5530=>"011011011",
    5531=>"001011011",
    5532=>"000010111",
    5533=>"110100000",
    5534=>"001101000",
    5535=>"000011011",
    5536=>"011011101",
    5537=>"111011101",
    5538=>"100010010",
    5539=>"010000111",
    5540=>"100100110",
    5541=>"000010001",
    5542=>"111111100",
    5543=>"111111100",
    5544=>"000010010",
    5545=>"000110110",
    5546=>"011110010",
    5547=>"110110001",
    5548=>"011001100",
    5549=>"000000011",
    5550=>"001101111",
    5551=>"111111111",
    5552=>"101001000",
    5553=>"001100101",
    5554=>"011011000",
    5555=>"010000000",
    5556=>"111011010",
    5557=>"000000000",
    5558=>"101000110",
    5559=>"000101111",
    5560=>"000011011",
    5561=>"111011000",
    5562=>"011000001",
    5563=>"000000110",
    5564=>"001111010",
    5565=>"000000010",
    5566=>"100111110",
    5567=>"001101000",
    5568=>"000011000",
    5569=>"010000000",
    5570=>"111111111",
    5571=>"111111110",
    5572=>"001110111",
    5573=>"100100001",
    5574=>"100000000",
    5575=>"000110000",
    5576=>"110101001",
    5577=>"000101101",
    5578=>"011000110",
    5579=>"010010000",
    5580=>"000000111",
    5581=>"111101111",
    5582=>"000000011",
    5583=>"101000000",
    5584=>"000000111",
    5585=>"110111011",
    5586=>"010000000",
    5587=>"100001000",
    5588=>"001001000",
    5589=>"000101111",
    5590=>"000111111",
    5591=>"101110101",
    5592=>"000110110",
    5593=>"111000000",
    5594=>"010110111",
    5595=>"000000000",
    5596=>"100011000",
    5597=>"011000100",
    5598=>"000010000",
    5599=>"110011010",
    5600=>"000110011",
    5601=>"001001011",
    5602=>"100000111",
    5603=>"000111111",
    5604=>"111100000",
    5605=>"000001000",
    5606=>"001111100",
    5607=>"000011011",
    5608=>"100000100",
    5609=>"001011011",
    5610=>"110101011",
    5611=>"100111000",
    5612=>"101101111",
    5613=>"111011000",
    5614=>"111111111",
    5615=>"100101000",
    5616=>"011000111",
    5617=>"011001000",
    5618=>"101101001",
    5619=>"010011000",
    5620=>"000100111",
    5621=>"111111000",
    5622=>"111110001",
    5623=>"111110000",
    5624=>"000000110",
    5625=>"111111000",
    5626=>"011000111",
    5627=>"100000001",
    5628=>"000011101",
    5629=>"000001000",
    5630=>"000010000",
    5631=>"000010000",
    5632=>"100110100",
    5633=>"001000100",
    5634=>"110110000",
    5635=>"111110000",
    5636=>"111111100",
    5637=>"011011110",
    5638=>"011110100",
    5639=>"100110100",
    5640=>"010001111",
    5641=>"001001011",
    5642=>"001001010",
    5643=>"111001111",
    5644=>"001001001",
    5645=>"111011110",
    5646=>"000001100",
    5647=>"100110100",
    5648=>"011001011",
    5649=>"000000101",
    5650=>"100100101",
    5651=>"100100100",
    5652=>"011001011",
    5653=>"111011001",
    5654=>"000000000",
    5655=>"110000011",
    5656=>"100100000",
    5657=>"100001110",
    5658=>"111011000",
    5659=>"001001011",
    5660=>"111110100",
    5661=>"000100000",
    5662=>"001001000",
    5663=>"111110000",
    5664=>"011001000",
    5665=>"100000000",
    5666=>"001001101",
    5667=>"001001111",
    5668=>"111110000",
    5669=>"100000011",
    5670=>"110110100",
    5671=>"011111011",
    5672=>"110100100",
    5673=>"110110111",
    5674=>"011001010",
    5675=>"100101111",
    5676=>"010110110",
    5677=>"110110010",
    5678=>"001111111",
    5679=>"110110000",
    5680=>"001001011",
    5681=>"101110111",
    5682=>"001001101",
    5683=>"110100000",
    5684=>"111000000",
    5685=>"001011011",
    5686=>"001000000",
    5687=>"100100000",
    5688=>"100100100",
    5689=>"000000000",
    5690=>"011000111",
    5691=>"001001001",
    5692=>"001000001",
    5693=>"001001011",
    5694=>"011011001",
    5695=>"110001111",
    5696=>"111111000",
    5697=>"101000000",
    5698=>"100110011",
    5699=>"000001010",
    5700=>"111110101",
    5701=>"110110000",
    5702=>"111100100",
    5703=>"101100110",
    5704=>"001001111",
    5705=>"001011010",
    5706=>"110100111",
    5707=>"101000000",
    5708=>"111110000",
    5709=>"001101110",
    5710=>"111110110",
    5711=>"001001001",
    5712=>"000100000",
    5713=>"110110110",
    5714=>"000001000",
    5715=>"111110100",
    5716=>"111111000",
    5717=>"000001011",
    5718=>"011011011",
    5719=>"011010000",
    5720=>"000000100",
    5721=>"011001100",
    5722=>"011110100",
    5723=>"011000000",
    5724=>"100100000",
    5725=>"111100100",
    5726=>"101101001",
    5727=>"101100100",
    5728=>"000001100",
    5729=>"000000000",
    5730=>"001111110",
    5731=>"100100000",
    5732=>"100110110",
    5733=>"110110000",
    5734=>"111111100",
    5735=>"110100100",
    5736=>"011010100",
    5737=>"000000000",
    5738=>"100111110",
    5739=>"001100110",
    5740=>"100000100",
    5741=>"101100111",
    5742=>"011011111",
    5743=>"011011110",
    5744=>"110110000",
    5745=>"000000110",
    5746=>"011011111",
    5747=>"100100100",
    5748=>"001001011",
    5749=>"000001101",
    5750=>"001001110",
    5751=>"001001011",
    5752=>"100100100",
    5753=>"110111110",
    5754=>"000100010",
    5755=>"001001111",
    5756=>"000000010",
    5757=>"001001111",
    5758=>"001000101",
    5759=>"001011011",
    5760=>"000000010",
    5761=>"101000111",
    5762=>"011101101",
    5763=>"010100111",
    5764=>"000100100",
    5765=>"010000000",
    5766=>"111110010",
    5767=>"010101101",
    5768=>"001011110",
    5769=>"010000001",
    5770=>"100101000",
    5771=>"011101100",
    5772=>"010000100",
    5773=>"111100110",
    5774=>"100001010",
    5775=>"010001100",
    5776=>"111100001",
    5777=>"000001011",
    5778=>"001111000",
    5779=>"100001001",
    5780=>"101110000",
    5781=>"011000000",
    5782=>"011101000",
    5783=>"111101100",
    5784=>"101001110",
    5785=>"110100101",
    5786=>"001111110",
    5787=>"100001111",
    5788=>"101011111",
    5789=>"000000011",
    5790=>"111011010",
    5791=>"000000100",
    5792=>"000000000",
    5793=>"100000011",
    5794=>"001001101",
    5795=>"000010101",
    5796=>"010111111",
    5797=>"110010110",
    5798=>"110000101",
    5799=>"101000010",
    5800=>"111111110",
    5801=>"010011111",
    5802=>"001100110",
    5803=>"100001010",
    5804=>"001110010",
    5805=>"000011001",
    5806=>"000011000",
    5807=>"010101101",
    5808=>"000000010",
    5809=>"111100000",
    5810=>"110111110",
    5811=>"011001001",
    5812=>"000000010",
    5813=>"000000100",
    5814=>"000010000",
    5815=>"010000100",
    5816=>"101001000",
    5817=>"000101001",
    5818=>"001010010",
    5819=>"101001110",
    5820=>"010100100",
    5821=>"000001100",
    5822=>"001111011",
    5823=>"000111101",
    5824=>"100011011",
    5825=>"101000000",
    5826=>"010010100",
    5827=>"000000000",
    5828=>"111011000",
    5829=>"000010110",
    5830=>"111110000",
    5831=>"100000000",
    5832=>"010010010",
    5833=>"101010110",
    5834=>"010110001",
    5835=>"000001000",
    5836=>"000010000",
    5837=>"001011000",
    5838=>"000101101",
    5839=>"111000001",
    5840=>"001100101",
    5841=>"111000000",
    5842=>"110111100",
    5843=>"011000000",
    5844=>"100001001",
    5845=>"111100000",
    5846=>"101011000",
    5847=>"111100000",
    5848=>"100111011",
    5849=>"000000001",
    5850=>"100000010",
    5851=>"010101100",
    5852=>"101001010",
    5853=>"010010110",
    5854=>"100100011",
    5855=>"101101000",
    5856=>"100010011",
    5857=>"111111000",
    5858=>"111011101",
    5859=>"000010011",
    5860=>"110110101",
    5861=>"111000100",
    5862=>"111000000",
    5863=>"000010000",
    5864=>"100001011",
    5865=>"000000100",
    5866=>"100000011",
    5867=>"011111111",
    5868=>"111111100",
    5869=>"111010000",
    5870=>"010010110",
    5871=>"001110110",
    5872=>"111111000",
    5873=>"001011110",
    5874=>"100000011",
    5875=>"101001111",
    5876=>"111100000",
    5877=>"010000000",
    5878=>"111010011",
    5879=>"000111011",
    5880=>"010111101",
    5881=>"010000110",
    5882=>"001100100",
    5883=>"000111101",
    5884=>"101000111",
    5885=>"111111111",
    5886=>"110000101",
    5887=>"000011111",
    5888=>"010111111",
    5889=>"000000000",
    5890=>"000111110",
    5891=>"111111110",
    5892=>"011011010",
    5893=>"101111011",
    5894=>"000100111",
    5895=>"111011010",
    5896=>"000101111",
    5897=>"111100000",
    5898=>"110000000",
    5899=>"011001010",
    5900=>"111100011",
    5901=>"010101111",
    5902=>"100111001",
    5903=>"110000011",
    5904=>"010110100",
    5905=>"011011000",
    5906=>"110001001",
    5907=>"100100011",
    5908=>"111000000",
    5909=>"010000001",
    5910=>"000001000",
    5911=>"111000110",
    5912=>"111100000",
    5913=>"110000010",
    5914=>"111111110",
    5915=>"000101100",
    5916=>"001000111",
    5917=>"100100000",
    5918=>"110100111",
    5919=>"111111000",
    5920=>"111101100",
    5921=>"100011000",
    5922=>"011001100",
    5923=>"001100001",
    5924=>"111101000",
    5925=>"010001101",
    5926=>"001011111",
    5927=>"000111111",
    5928=>"111000000",
    5929=>"110001000",
    5930=>"010101111",
    5931=>"001001110",
    5932=>"011001000",
    5933=>"111111000",
    5934=>"011111001",
    5935=>"111111000",
    5936=>"111000000",
    5937=>"000010111",
    5938=>"111001000",
    5939=>"000111011",
    5940=>"011100000",
    5941=>"001000000",
    5942=>"001000111",
    5943=>"000111111",
    5944=>"111000000",
    5945=>"111000000",
    5946=>"111000000",
    5947=>"000000001",
    5948=>"000000000",
    5949=>"000110111",
    5950=>"100101001",
    5951=>"001001011",
    5952=>"010100110",
    5953=>"000010110",
    5954=>"111000000",
    5955=>"000000000",
    5956=>"111100100",
    5957=>"000110110",
    5958=>"011001000",
    5959=>"111111000",
    5960=>"100111001",
    5961=>"000110110",
    5962=>"111000000",
    5963=>"000000000",
    5964=>"100000110",
    5965=>"110111000",
    5966=>"111000000",
    5967=>"000110111",
    5968=>"011000010",
    5969=>"000110011",
    5970=>"000010111",
    5971=>"111101000",
    5972=>"000011111",
    5973=>"000110111",
    5974=>"000000000",
    5975=>"111101101",
    5976=>"001110000",
    5977=>"100000000",
    5978=>"011011111",
    5979=>"110111000",
    5980=>"100100001",
    5981=>"011001000",
    5982=>"101111111",
    5983=>"000000110",
    5984=>"100100000",
    5985=>"000001110",
    5986=>"110000001",
    5987=>"111000000",
    5988=>"111001010",
    5989=>"010111000",
    5990=>"000011110",
    5991=>"010111111",
    5992=>"110101101",
    5993=>"111010111",
    5994=>"000101001",
    5995=>"111101000",
    5996=>"000111111",
    5997=>"000111111",
    5998=>"110101111",
    5999=>"000101111",
    6000=>"101001000",
    6001=>"000000110",
    6002=>"000111111",
    6003=>"000111011",
    6004=>"111001111",
    6005=>"000111001",
    6006=>"000000001",
    6007=>"100100111",
    6008=>"001000000",
    6009=>"111011001",
    6010=>"010101000",
    6011=>"010000000",
    6012=>"100110110",
    6013=>"000000010",
    6014=>"110000000",
    6015=>"100100011",
    6016=>"111000110",
    6017=>"101100011",
    6018=>"100000100",
    6019=>"110111000",
    6020=>"011001110",
    6021=>"101001000",
    6022=>"000000111",
    6023=>"111001111",
    6024=>"110110111",
    6025=>"101110100",
    6026=>"000010111",
    6027=>"010100100",
    6028=>"100110101",
    6029=>"111111111",
    6030=>"100000000",
    6031=>"110000100",
    6032=>"110110111",
    6033=>"100100111",
    6034=>"111001111",
    6035=>"110100000",
    6036=>"001000010",
    6037=>"100000000",
    6038=>"000000010",
    6039=>"011011011",
    6040=>"100100110",
    6041=>"010100101",
    6042=>"100000000",
    6043=>"011000000",
    6044=>"001111111",
    6045=>"110100100",
    6046=>"000001001",
    6047=>"000000101",
    6048=>"101111111",
    6049=>"000000100",
    6050=>"011001100",
    6051=>"010111010",
    6052=>"100100111",
    6053=>"000000101",
    6054=>"100000111",
    6055=>"010011010",
    6056=>"000100101",
    6057=>"000101001",
    6058=>"100100111",
    6059=>"100110111",
    6060=>"011001000",
    6061=>"011001000",
    6062=>"100100010",
    6063=>"111000100",
    6064=>"000111111",
    6065=>"001101110",
    6066=>"000010000",
    6067=>"110000000",
    6068=>"010110000",
    6069=>"100101111",
    6070=>"000010000",
    6071=>"000000010",
    6072=>"000011011",
    6073=>"111100100",
    6074=>"000001000",
    6075=>"111000000",
    6076=>"001101010",
    6077=>"011011011",
    6078=>"101100100",
    6079=>"000000000",
    6080=>"011011000",
    6081=>"100000011",
    6082=>"000011110",
    6083=>"100000000",
    6084=>"011010000",
    6085=>"110110111",
    6086=>"010100111",
    6087=>"010100010",
    6088=>"011111000",
    6089=>"000010010",
    6090=>"100101101",
    6091=>"100100111",
    6092=>"100010111",
    6093=>"100100111",
    6094=>"111011000",
    6095=>"111001001",
    6096=>"011011001",
    6097=>"100000000",
    6098=>"000111000",
    6099=>"100000100",
    6100=>"001001111",
    6101=>"011010000",
    6102=>"100000011",
    6103=>"010111100",
    6104=>"000100111",
    6105=>"001101000",
    6106=>"001000000",
    6107=>"101000000",
    6108=>"000001111",
    6109=>"000000000",
    6110=>"110100001",
    6111=>"111111111",
    6112=>"001001010",
    6113=>"100110011",
    6114=>"000111111",
    6115=>"000101111",
    6116=>"000000010",
    6117=>"100101101",
    6118=>"100100100",
    6119=>"000000000",
    6120=>"100000010",
    6121=>"000000010",
    6122=>"000001000",
    6123=>"111001010",
    6124=>"100100111",
    6125=>"110100001",
    6126=>"110101110",
    6127=>"100101110",
    6128=>"000010000",
    6129=>"000111111",
    6130=>"111000000",
    6131=>"111101110",
    6132=>"010001010",
    6133=>"100000000",
    6134=>"101000000",
    6135=>"100100100",
    6136=>"000101100",
    6137=>"101000100",
    6138=>"000000010",
    6139=>"101101000",
    6140=>"100000100",
    6141=>"010011010",
    6142=>"000110111",
    6143=>"000100111",
    6144=>"111010000",
    6145=>"101101111",
    6146=>"111010000",
    6147=>"000001111",
    6148=>"111100100",
    6149=>"101111111",
    6150=>"100101111",
    6151=>"000000001",
    6152=>"110000000",
    6153=>"100001110",
    6154=>"111111000",
    6155=>"100111111",
    6156=>"000000111",
    6157=>"100111111",
    6158=>"000000100",
    6159=>"110001100",
    6160=>"000110111",
    6161=>"000111111",
    6162=>"000000011",
    6163=>"110001001",
    6164=>"111000000",
    6165=>"000000000",
    6166=>"000100010",
    6167=>"000000111",
    6168=>"000110110",
    6169=>"101111101",
    6170=>"111000000",
    6171=>"000100101",
    6172=>"000110011",
    6173=>"000000110",
    6174=>"010011100",
    6175=>"000000001",
    6176=>"000101111",
    6177=>"000100111",
    6178=>"110010011",
    6179=>"100010000",
    6180=>"101111111",
    6181=>"000100010",
    6182=>"001000111",
    6183=>"111000000",
    6184=>"100000000",
    6185=>"101111101",
    6186=>"000111111",
    6187=>"001011110",
    6188=>"000100001",
    6189=>"000101111",
    6190=>"000000001",
    6191=>"000000111",
    6192=>"000110111",
    6193=>"111000000",
    6194=>"000000100",
    6195=>"100000111",
    6196=>"000010011",
    6197=>"000111111",
    6198=>"000111111",
    6199=>"110010000",
    6200=>"101111111",
    6201=>"100101000",
    6202=>"000111011",
    6203=>"000001010",
    6204=>"000000010",
    6205=>"110010111",
    6206=>"000000000",
    6207=>"001001000",
    6208=>"011000000",
    6209=>"111010000",
    6210=>"100111110",
    6211=>"000000000",
    6212=>"100110111",
    6213=>"000001111",
    6214=>"011111000",
    6215=>"000000000",
    6216=>"000011111",
    6217=>"100000001",
    6218=>"111111111",
    6219=>"000101111",
    6220=>"101000111",
    6221=>"111000000",
    6222=>"111001111",
    6223=>"111000100",
    6224=>"111101101",
    6225=>"101111001",
    6226=>"111000000",
    6227=>"111110111",
    6228=>"101100110",
    6229=>"001011010",
    6230=>"101011010",
    6231=>"000000000",
    6232=>"000111001",
    6233=>"000110110",
    6234=>"011000100",
    6235=>"000010000",
    6236=>"110000011",
    6237=>"010000001",
    6238=>"110000000",
    6239=>"001101000",
    6240=>"001001111",
    6241=>"011001111",
    6242=>"111010000",
    6243=>"000111010",
    6244=>"101000000",
    6245=>"000001111",
    6246=>"100100110",
    6247=>"000000111",
    6248=>"000000110",
    6249=>"000000000",
    6250=>"111011000",
    6251=>"001001111",
    6252=>"111111111",
    6253=>"101000000",
    6254=>"100110011",
    6255=>"111101100",
    6256=>"111000000",
    6257=>"110000000",
    6258=>"000000111",
    6259=>"000000100",
    6260=>"111111000",
    6261=>"000101010",
    6262=>"000111111",
    6263=>"000100000",
    6264=>"000000100",
    6265=>"000101011",
    6266=>"000000111",
    6267=>"000001111",
    6268=>"110100010",
    6269=>"101101111",
    6270=>"110000011",
    6271=>"111001000",
    6272=>"110110100",
    6273=>"111001001",
    6274=>"000001011",
    6275=>"000011011",
    6276=>"101111111",
    6277=>"100100001",
    6278=>"000110110",
    6279=>"101100100",
    6280=>"101011101",
    6281=>"010001001",
    6282=>"000001100",
    6283=>"100011111",
    6284=>"101110110",
    6285=>"000111001",
    6286=>"011011011",
    6287=>"000100001",
    6288=>"011011110",
    6289=>"000000111",
    6290=>"101111100",
    6291=>"000100000",
    6292=>"001001011",
    6293=>"100000000",
    6294=>"011001011",
    6295=>"001000111",
    6296=>"000000000",
    6297=>"110011011",
    6298=>"000100101",
    6299=>"111110100",
    6300=>"110101101",
    6301=>"100111110",
    6302=>"011111111",
    6303=>"111110100",
    6304=>"110101001",
    6305=>"010000000",
    6306=>"100000110",
    6307=>"000100100",
    6308=>"100100100",
    6309=>"001011011",
    6310=>"010011011",
    6311=>"100100100",
    6312=>"100100000",
    6313=>"110100100",
    6314=>"111111101",
    6315=>"111111101",
    6316=>"001000100",
    6317=>"100100101",
    6318=>"100000100",
    6319=>"011011011",
    6320=>"100110110",
    6321=>"001001011",
    6322=>"001001011",
    6323=>"000000000",
    6324=>"000000100",
    6325=>"000011000",
    6326=>"100110110",
    6327=>"101001000",
    6328=>"111110100",
    6329=>"000000100",
    6330=>"110011011",
    6331=>"000100100",
    6332=>"010010010",
    6333=>"111001011",
    6334=>"000000110",
    6335=>"010111101",
    6336=>"110110111",
    6337=>"011001011",
    6338=>"010100010",
    6339=>"101110110",
    6340=>"111110100",
    6341=>"001000000",
    6342=>"110010000",
    6343=>"011011011",
    6344=>"001011011",
    6345=>"000010000",
    6346=>"000000000",
    6347=>"001001001",
    6348=>"011000100",
    6349=>"110110110",
    6350=>"000000000",
    6351=>"110011010",
    6352=>"001110100",
    6353=>"001111001",
    6354=>"100100110",
    6355=>"001001001",
    6356=>"001111111",
    6357=>"001000011",
    6358=>"010000100",
    6359=>"100000001",
    6360=>"100000000",
    6361=>"110011010",
    6362=>"010110100",
    6363=>"011011011",
    6364=>"000100100",
    6365=>"000001010",
    6366=>"010001100",
    6367=>"010011010",
    6368=>"001001001",
    6369=>"100100100",
    6370=>"100100100",
    6371=>"001011011",
    6372=>"101100110",
    6373=>"000100000",
    6374=>"100101000",
    6375=>"100000011",
    6376=>"011111011",
    6377=>"011001010",
    6378=>"101111111",
    6379=>"011001011",
    6380=>"000000000",
    6381=>"000001000",
    6382=>"000100111",
    6383=>"000000000",
    6384=>"100100101",
    6385=>"001101111",
    6386=>"000010011",
    6387=>"110011011",
    6388=>"010111010",
    6389=>"001001000",
    6390=>"101110111",
    6391=>"111011011",
    6392=>"100100100",
    6393=>"011011011",
    6394=>"001101001",
    6395=>"001111100",
    6396=>"100000000",
    6397=>"010011011",
    6398=>"001000000",
    6399=>"001111101",
    6400=>"111110000",
    6401=>"000000001",
    6402=>"101111011",
    6403=>"110000111",
    6404=>"100011000",
    6405=>"101111100",
    6406=>"111101000",
    6407=>"001000111",
    6408=>"001100000",
    6409=>"100111001",
    6410=>"101001111",
    6411=>"000100100",
    6412=>"001000101",
    6413=>"111111111",
    6414=>"000001111",
    6415=>"000000111",
    6416=>"010011001",
    6417=>"101100111",
    6418=>"010110011",
    6419=>"001000000",
    6420=>"000000111",
    6421=>"000000000",
    6422=>"001000100",
    6423=>"000111111",
    6424=>"001001100",
    6425=>"110101011",
    6426=>"111100000",
    6427=>"110110110",
    6428=>"000100001",
    6429=>"000100000",
    6430=>"100101000",
    6431=>"101111111",
    6432=>"111111101",
    6433=>"111100000",
    6434=>"011101100",
    6435=>"011111000",
    6436=>"111010000",
    6437=>"111101111",
    6438=>"101101100",
    6439=>"111010000",
    6440=>"000000000",
    6441=>"111010000",
    6442=>"111000000",
    6443=>"111011000",
    6444=>"001110010",
    6445=>"101111000",
    6446=>"000010000",
    6447=>"000100111",
    6448=>"000010101",
    6449=>"101101101",
    6450=>"100100110",
    6451=>"011011000",
    6452=>"000100100",
    6453=>"011111000",
    6454=>"000000000",
    6455=>"000010010",
    6456=>"110111010",
    6457=>"111011000",
    6458=>"001011111",
    6459=>"010110101",
    6460=>"000000001",
    6461=>"101100101",
    6462=>"111011011",
    6463=>"101100010",
    6464=>"001100111",
    6465=>"111111110",
    6466=>"001101110",
    6467=>"000100101",
    6468=>"001111000",
    6469=>"111110000",
    6470=>"110110101",
    6471=>"001011011",
    6472=>"000000011",
    6473=>"110000000",
    6474=>"101100110",
    6475=>"000000000",
    6476=>"000000111",
    6477=>"011011000",
    6478=>"110110000",
    6479=>"000001000",
    6480=>"000010011",
    6481=>"001000001",
    6482=>"000000111",
    6483=>"100100011",
    6484=>"010011000",
    6485=>"000000101",
    6486=>"111110010",
    6487=>"000110010",
    6488=>"011011100",
    6489=>"110111101",
    6490=>"011001000",
    6491=>"111010000",
    6492=>"111111000",
    6493=>"010000110",
    6494=>"011001000",
    6495=>"010110111",
    6496=>"110011000",
    6497=>"110110000",
    6498=>"101001111",
    6499=>"111010000",
    6500=>"010001000",
    6501=>"000000010",
    6502=>"100000100",
    6503=>"010000000",
    6504=>"001000001",
    6505=>"101100111",
    6506=>"101001001",
    6507=>"101000000",
    6508=>"111111000",
    6509=>"101001100",
    6510=>"001111111",
    6511=>"000100100",
    6512=>"000000000",
    6513=>"100000000",
    6514=>"110000000",
    6515=>"101100111",
    6516=>"000100111",
    6517=>"001001001",
    6518=>"111000010",
    6519=>"101011111",
    6520=>"100111000",
    6521=>"000000111",
    6522=>"100100111",
    6523=>"000101111",
    6524=>"110110000",
    6525=>"000111110",
    6526=>"111111000",
    6527=>"111111000",
    6528=>"110011111",
    6529=>"000000010",
    6530=>"111011000",
    6531=>"100101000",
    6532=>"010010100",
    6533=>"110111010",
    6534=>"110111010",
    6535=>"000010111",
    6536=>"101001000",
    6537=>"010000000",
    6538=>"101101011",
    6539=>"101110010",
    6540=>"000000000",
    6541=>"111000110",
    6542=>"011110000",
    6543=>"000011111",
    6544=>"101000111",
    6545=>"111010000",
    6546=>"101111111",
    6547=>"111000000",
    6548=>"111110000",
    6549=>"010010100",
    6550=>"111101010",
    6551=>"000000100",
    6552=>"101111111",
    6553=>"110001001",
    6554=>"100111111",
    6555=>"110111111",
    6556=>"001111111",
    6557=>"111111000",
    6558=>"111111100",
    6559=>"000000111",
    6560=>"000010010",
    6561=>"000101111",
    6562=>"111000000",
    6563=>"001000000",
    6564=>"111000000",
    6565=>"111110010",
    6566=>"000111010",
    6567=>"111111000",
    6568=>"111100000",
    6569=>"100001111",
    6570=>"111111000",
    6571=>"111111101",
    6572=>"000000111",
    6573=>"000000010",
    6574=>"000000000",
    6575=>"110111110",
    6576=>"000000000",
    6577=>"111111000",
    6578=>"000100111",
    6579=>"001000001",
    6580=>"001011101",
    6581=>"000001111",
    6582=>"010000111",
    6583=>"110110010",
    6584=>"101111111",
    6585=>"000000010",
    6586=>"000000000",
    6587=>"011011000",
    6588=>"111111110",
    6589=>"111111000",
    6590=>"111111111",
    6591=>"101000101",
    6592=>"000010111",
    6593=>"000001010",
    6594=>"000000000",
    6595=>"000000100",
    6596=>"000000001",
    6597=>"010111000",
    6598=>"000000000",
    6599=>"001111111",
    6600=>"100000010",
    6601=>"111011000",
    6602=>"001000111",
    6603=>"010011000",
    6604=>"001001101",
    6605=>"000000111",
    6606=>"000111111",
    6607=>"111111111",
    6608=>"100100100",
    6609=>"111010000",
    6610=>"001001111",
    6611=>"101011010",
    6612=>"000011010",
    6613=>"100000000",
    6614=>"110111111",
    6615=>"111111000",
    6616=>"101110100",
    6617=>"000000000",
    6618=>"001001000",
    6619=>"010011000",
    6620=>"101111011",
    6621=>"001000100",
    6622=>"110111010",
    6623=>"000010000",
    6624=>"100100110",
    6625=>"000100000",
    6626=>"000000111",
    6627=>"000101111",
    6628=>"000111111",
    6629=>"100010011",
    6630=>"111011000",
    6631=>"000000110",
    6632=>"000001111",
    6633=>"101001011",
    6634=>"111111001",
    6635=>"000000000",
    6636=>"000000000",
    6637=>"111110000",
    6638=>"000000011",
    6639=>"011111100",
    6640=>"011010101",
    6641=>"000000010",
    6642=>"111000000",
    6643=>"111111000",
    6644=>"101101111",
    6645=>"000000000",
    6646=>"000001010",
    6647=>"000001101",
    6648=>"001001111",
    6649=>"000111111",
    6650=>"100000110",
    6651=>"000000111",
    6652=>"110110000",
    6653=>"000111111",
    6654=>"010011001",
    6655=>"010111101",
    6656=>"000000110",
    6657=>"111101111",
    6658=>"100101111",
    6659=>"001010001",
    6660=>"111111101",
    6661=>"111111111",
    6662=>"000000000",
    6663=>"000000000",
    6664=>"000000000",
    6665=>"010011011",
    6666=>"001001110",
    6667=>"111101110",
    6668=>"111111111",
    6669=>"111111010",
    6670=>"101000000",
    6671=>"001001000",
    6672=>"010100100",
    6673=>"111111011",
    6674=>"100111011",
    6675=>"100101110",
    6676=>"000000000",
    6677=>"111111111",
    6678=>"111001001",
    6679=>"000000010",
    6680=>"011111110",
    6681=>"110111011",
    6682=>"000000000",
    6683=>"011111100",
    6684=>"111100101",
    6685=>"110100010",
    6686=>"100101111",
    6687=>"000000000",
    6688=>"001101111",
    6689=>"000000000",
    6690=>"011101100",
    6691=>"011001010",
    6692=>"100000100",
    6693=>"111101010",
    6694=>"000010000",
    6695=>"001111111",
    6696=>"000000000",
    6697=>"110100000",
    6698=>"110110011",
    6699=>"110111010",
    6700=>"010100010",
    6701=>"111011011",
    6702=>"000101011",
    6703=>"110111111",
    6704=>"010000110",
    6705=>"001111011",
    6706=>"111111110",
    6707=>"001001111",
    6708=>"111100011",
    6709=>"000000000",
    6710=>"010000000",
    6711=>"000000000",
    6712=>"000000000",
    6713=>"111101000",
    6714=>"001010100",
    6715=>"100010101",
    6716=>"101000000",
    6717=>"000000000",
    6718=>"011110111",
    6719=>"111011000",
    6720=>"110110101",
    6721=>"000000000",
    6722=>"111011110",
    6723=>"111010101",
    6724=>"111111111",
    6725=>"100001110",
    6726=>"101010010",
    6727=>"010000000",
    6728=>"100001001",
    6729=>"100110001",
    6730=>"001000110",
    6731=>"000000010",
    6732=>"110100000",
    6733=>"000001100",
    6734=>"001000101",
    6735=>"111000101",
    6736=>"000000000",
    6737=>"000000110",
    6738=>"100111010",
    6739=>"111111111",
    6740=>"111000001",
    6741=>"011111111",
    6742=>"111111111",
    6743=>"000000000",
    6744=>"010011100",
    6745=>"111111111",
    6746=>"000101011",
    6747=>"111000100",
    6748=>"001011011",
    6749=>"000100110",
    6750=>"000000000",
    6751=>"011100000",
    6752=>"000000000",
    6753=>"000011001",
    6754=>"001100110",
    6755=>"010110111",
    6756=>"000010000",
    6757=>"000000000",
    6758=>"011000111",
    6759=>"110101011",
    6760=>"011011011",
    6761=>"110000001",
    6762=>"100101011",
    6763=>"010000010",
    6764=>"010000000",
    6765=>"000000100",
    6766=>"101110110",
    6767=>"000000000",
    6768=>"111111111",
    6769=>"011110110",
    6770=>"000100000",
    6771=>"111111111",
    6772=>"111001001",
    6773=>"100000000",
    6774=>"000000000",
    6775=>"111111011",
    6776=>"000000010",
    6777=>"000000000",
    6778=>"110110111",
    6779=>"111000000",
    6780=>"000000000",
    6781=>"000000000",
    6782=>"000000000",
    6783=>"000111010",
    6784=>"100011000",
    6785=>"011011011",
    6786=>"111101111",
    6787=>"110100100",
    6788=>"000001000",
    6789=>"000011001",
    6790=>"010010010",
    6791=>"101100101",
    6792=>"101111101",
    6793=>"100110010",
    6794=>"000010010",
    6795=>"111100101",
    6796=>"111010111",
    6797=>"111100111",
    6798=>"111111101",
    6799=>"000010010",
    6800=>"111001111",
    6801=>"000010011",
    6802=>"110101100",
    6803=>"100100001",
    6804=>"000001011",
    6805=>"100000000",
    6806=>"111100111",
    6807=>"011000010",
    6808=>"010111001",
    6809=>"110100101",
    6810=>"110100100",
    6811=>"011110100",
    6812=>"110010000",
    6813=>"000001011",
    6814=>"110111100",
    6815=>"111111010",
    6816=>"111011000",
    6817=>"000001001",
    6818=>"001001000",
    6819=>"010000011",
    6820=>"110100001",
    6821=>"010101000",
    6822=>"010101100",
    6823=>"111111010",
    6824=>"111010001",
    6825=>"110011111",
    6826=>"100000000",
    6827=>"001100000",
    6828=>"011000110",
    6829=>"001010001",
    6830=>"001000000",
    6831=>"111111111",
    6832=>"111101011",
    6833=>"111101111",
    6834=>"111100000",
    6835=>"110100000",
    6836=>"100110100",
    6837=>"000000000",
    6838=>"000000000",
    6839=>"101100111",
    6840=>"100011011",
    6841=>"011111010",
    6842=>"000001100",
    6843=>"000000100",
    6844=>"101100100",
    6845=>"000000100",
    6846=>"111011100",
    6847=>"000111011",
    6848=>"111011011",
    6849=>"011001100",
    6850=>"100000010",
    6851=>"000011111",
    6852=>"111111000",
    6853=>"101001000",
    6854=>"100000111",
    6855=>"010011111",
    6856=>"111111110",
    6857=>"000000000",
    6858=>"011011011",
    6859=>"010000000",
    6860=>"010101010",
    6861=>"001101100",
    6862=>"101111111",
    6863=>"000000001",
    6864=>"100000111",
    6865=>"000000000",
    6866=>"111011001",
    6867=>"001111101",
    6868=>"100100100",
    6869=>"000000000",
    6870=>"110100100",
    6871=>"000111010",
    6872=>"000011011",
    6873=>"111101100",
    6874=>"001000000",
    6875=>"010000000",
    6876=>"110101101",
    6877=>"001001000",
    6878=>"101000000",
    6879=>"111101001",
    6880=>"100111000",
    6881=>"001001000",
    6882=>"010110000",
    6883=>"000011010",
    6884=>"111001111",
    6885=>"101100111",
    6886=>"100000000",
    6887=>"011010001",
    6888=>"111111111",
    6889=>"000000000",
    6890=>"000101001",
    6891=>"111011010",
    6892=>"011001101",
    6893=>"111101111",
    6894=>"110000000",
    6895=>"010111000",
    6896=>"010011010",
    6897=>"100000011",
    6898=>"010001111",
    6899=>"001000000",
    6900=>"101000000",
    6901=>"101101100",
    6902=>"011000101",
    6903=>"111100010",
    6904=>"011111111",
    6905=>"001000111",
    6906=>"111111111",
    6907=>"100001000",
    6908=>"000000110",
    6909=>"101100101",
    6910=>"000111001",
    6911=>"010110000",
    6912=>"010101111",
    6913=>"100111111",
    6914=>"001000001",
    6915=>"111110100",
    6916=>"000001001",
    6917=>"111110100",
    6918=>"001111100",
    6919=>"000000000",
    6920=>"001000111",
    6921=>"001011100",
    6922=>"110000001",
    6923=>"000000000",
    6924=>"000110100",
    6925=>"110110100",
    6926=>"111111111",
    6927=>"111111111",
    6928=>"000000000",
    6929=>"100100000",
    6930=>"000001000",
    6931=>"111110110",
    6932=>"000100100",
    6933=>"100000001",
    6934=>"100001010",
    6935=>"101011001",
    6936=>"000111111",
    6937=>"100100111",
    6938=>"001001001",
    6939=>"000000011",
    6940=>"101111101",
    6941=>"111101111",
    6942=>"000000011",
    6943=>"100000000",
    6944=>"000000000",
    6945=>"110110100",
    6946=>"000000001",
    6947=>"000010010",
    6948=>"011111100",
    6949=>"001010100",
    6950=>"011110100",
    6951=>"000001011",
    6952=>"000000011",
    6953=>"111111111",
    6954=>"101111111",
    6955=>"110111111",
    6956=>"000000000",
    6957=>"001000001",
    6958=>"001011001",
    6959=>"010110000",
    6960=>"101101100",
    6961=>"000001011",
    6962=>"000000000",
    6963=>"001001101",
    6964=>"111101001",
    6965=>"010000000",
    6966=>"111100000",
    6967=>"010000000",
    6968=>"110111001",
    6969=>"100110011",
    6970=>"101101111",
    6971=>"000001011",
    6972=>"100101001",
    6973=>"000000000",
    6974=>"001000001",
    6975=>"111110100",
    6976=>"010000000",
    6977=>"010000010",
    6978=>"111000100",
    6979=>"110010100",
    6980=>"110101001",
    6981=>"110111111",
    6982=>"111100110",
    6983=>"100100000",
    6984=>"111111100",
    6985=>"101111111",
    6986=>"000000000",
    6987=>"100000010",
    6988=>"000100100",
    6989=>"000011011",
    6990=>"111110101",
    6991=>"001001000",
    6992=>"000010011",
    6993=>"111101101",
    6994=>"100000000",
    6995=>"011111010",
    6996=>"001001011",
    6997=>"000011000",
    6998=>"000000000",
    6999=>"111001001",
    7000=>"000000000",
    7001=>"000110111",
    7002=>"000001011",
    7003=>"000000000",
    7004=>"101111110",
    7005=>"000000000",
    7006=>"110101011",
    7007=>"000010000",
    7008=>"111011010",
    7009=>"000010000",
    7010=>"011110100",
    7011=>"011100000",
    7012=>"000010000",
    7013=>"100011110",
    7014=>"000000011",
    7015=>"110101011",
    7016=>"111110000",
    7017=>"100000001",
    7018=>"111111101",
    7019=>"110010111",
    7020=>"000000100",
    7021=>"000100000",
    7022=>"100100000",
    7023=>"011000000",
    7024=>"110100100",
    7025=>"000010110",
    7026=>"100011011",
    7027=>"000011011",
    7028=>"000111010",
    7029=>"100000001",
    7030=>"000010100",
    7031=>"111011011",
    7032=>"000000000",
    7033=>"110100010",
    7034=>"000000000",
    7035=>"110010000",
    7036=>"000111011",
    7037=>"111111010",
    7038=>"100001001",
    7039=>"110111110",
    7040=>"100000110",
    7041=>"111010010",
    7042=>"000000000",
    7043=>"110111110",
    7044=>"000000100",
    7045=>"010111011",
    7046=>"010101011",
    7047=>"000000101",
    7048=>"110111111",
    7049=>"010001000",
    7050=>"011001000",
    7051=>"011101100",
    7052=>"000111000",
    7053=>"010110010",
    7054=>"000010010",
    7055=>"000000101",
    7056=>"011111110",
    7057=>"110111110",
    7058=>"001101100",
    7059=>"000111001",
    7060=>"010000000",
    7061=>"000000111",
    7062=>"000000100",
    7063=>"000000111",
    7064=>"001001001",
    7065=>"110001001",
    7066=>"000000100",
    7067=>"011111110",
    7068=>"001001001",
    7069=>"111100111",
    7070=>"000100110",
    7071=>"000000000",
    7072=>"101111001",
    7073=>"111100100",
    7074=>"001000010",
    7075=>"111101001",
    7076=>"111111001",
    7077=>"011001000",
    7078=>"000011010",
    7079=>"111110010",
    7080=>"111101111",
    7081=>"101001111",
    7082=>"111111111",
    7083=>"011100110",
    7084=>"111001101",
    7085=>"111111101",
    7086=>"001001001",
    7087=>"110110110",
    7088=>"111111100",
    7089=>"000011000",
    7090=>"111110110",
    7091=>"001110100",
    7092=>"000000110",
    7093=>"001000000",
    7094=>"111001101",
    7095=>"100101111",
    7096=>"100000100",
    7097=>"111111101",
    7098=>"111000000",
    7099=>"000000000",
    7100=>"100000001",
    7101=>"100000000",
    7102=>"110111101",
    7103=>"011101011",
    7104=>"001000000",
    7105=>"000010010",
    7106=>"111101101",
    7107=>"000100111",
    7108=>"111111100",
    7109=>"001100100",
    7110=>"101000000",
    7111=>"101111111",
    7112=>"010111011",
    7113=>"001000000",
    7114=>"111111011",
    7115=>"000000000",
    7116=>"111100100",
    7117=>"000000001",
    7118=>"111010000",
    7119=>"000110010",
    7120=>"010010000",
    7121=>"111110111",
    7122=>"010100111",
    7123=>"110000000",
    7124=>"110001001",
    7125=>"000000000",
    7126=>"101110011",
    7127=>"100110111",
    7128=>"001000000",
    7129=>"110110101",
    7130=>"000000000",
    7131=>"110101101",
    7132=>"011011011",
    7133=>"001001001",
    7134=>"000000011",
    7135=>"100000000",
    7136=>"111111111",
    7137=>"110111011",
    7138=>"000000000",
    7139=>"111111111",
    7140=>"010011110",
    7141=>"101001000",
    7142=>"111011011",
    7143=>"000000101",
    7144=>"000010000",
    7145=>"000000000",
    7146=>"110101111",
    7147=>"101000111",
    7148=>"000000111",
    7149=>"101000111",
    7150=>"111001011",
    7151=>"001111111",
    7152=>"000000101",
    7153=>"000000111",
    7154=>"101111011",
    7155=>"001000101",
    7156=>"000000001",
    7157=>"001000000",
    7158=>"001000010",
    7159=>"110011111",
    7160=>"111111111",
    7161=>"011111111",
    7162=>"000100000",
    7163=>"101100111",
    7164=>"000110011",
    7165=>"110111111",
    7166=>"000000000",
    7167=>"000100110",
    7168=>"111011000",
    7169=>"101101100",
    7170=>"000000111",
    7171=>"111110000",
    7172=>"110110011",
    7173=>"000000100",
    7174=>"111111101",
    7175=>"111111000",
    7176=>"000101111",
    7177=>"001001001",
    7178=>"011000000",
    7179=>"011010001",
    7180=>"100000010",
    7181=>"110110010",
    7182=>"000001001",
    7183=>"011001000",
    7184=>"000010011",
    7185=>"111011000",
    7186=>"011001100",
    7187=>"011011110",
    7188=>"001001111",
    7189=>"010010000",
    7190=>"100000000",
    7191=>"000100111",
    7192=>"110100001",
    7193=>"101011111",
    7194=>"011001100",
    7195=>"100110111",
    7196=>"010000000",
    7197=>"111001000",
    7198=>"001000101",
    7199=>"000010111",
    7200=>"010000000",
    7201=>"000000000",
    7202=>"101110111",
    7203=>"111111111",
    7204=>"100001111",
    7205=>"111101000",
    7206=>"110111000",
    7207=>"111101000",
    7208=>"000000000",
    7209=>"111111111",
    7210=>"001000000",
    7211=>"011111110",
    7212=>"000111111",
    7213=>"000000000",
    7214=>"011111000",
    7215=>"111111000",
    7216=>"100100011",
    7217=>"111000000",
    7218=>"000010111",
    7219=>"110100001",
    7220=>"011001000",
    7221=>"000000000",
    7222=>"000000111",
    7223=>"100101111",
    7224=>"001111111",
    7225=>"100111111",
    7226=>"100100000",
    7227=>"111111111",
    7228=>"111010000",
    7229=>"111111000",
    7230=>"011000110",
    7231=>"000110110",
    7232=>"111011010",
    7233=>"111010011",
    7234=>"000000000",
    7235=>"011000001",
    7236=>"000000111",
    7237=>"011011100",
    7238=>"000000010",
    7239=>"111111000",
    7240=>"000010110",
    7241=>"100000111",
    7242=>"000000010",
    7243=>"111000000",
    7244=>"000100111",
    7245=>"000011110",
    7246=>"000100111",
    7247=>"000000000",
    7248=>"000000101",
    7249=>"111001000",
    7250=>"010011000",
    7251=>"100100000",
    7252=>"110000001",
    7253=>"111000000",
    7254=>"010011111",
    7255=>"001101101",
    7256=>"111111001",
    7257=>"111111111",
    7258=>"000100000",
    7259=>"000000111",
    7260=>"111011011",
    7261=>"110110010",
    7262=>"110110000",
    7263=>"001000111",
    7264=>"000000111",
    7265=>"010001100",
    7266=>"110000000",
    7267=>"000010111",
    7268=>"011000000",
    7269=>"101000000",
    7270=>"111100000",
    7271=>"111111110",
    7272=>"111100000",
    7273=>"000111011",
    7274=>"100000000",
    7275=>"110111111",
    7276=>"000000000",
    7277=>"011010000",
    7278=>"000111111",
    7279=>"000000100",
    7280=>"000000010",
    7281=>"111010010",
    7282=>"001000000",
    7283=>"011000000",
    7284=>"000010111",
    7285=>"011001000",
    7286=>"101101000",
    7287=>"000000000",
    7288=>"100000011",
    7289=>"000000010",
    7290=>"111000000",
    7291=>"010010111",
    7292=>"110100000",
    7293=>"101100111",
    7294=>"000000101",
    7295=>"001011001",
    7296=>"000000000",
    7297=>"101101000",
    7298=>"000000000",
    7299=>"111111111",
    7300=>"110110100",
    7301=>"000000000",
    7302=>"010011010",
    7303=>"111111111",
    7304=>"011111110",
    7305=>"010010010",
    7306=>"000000000",
    7307=>"000000000",
    7308=>"110111110",
    7309=>"010111010",
    7310=>"010110111",
    7311=>"000001001",
    7312=>"110110110",
    7313=>"110011110",
    7314=>"011111111",
    7315=>"000001001",
    7316=>"111000000",
    7317=>"000000101",
    7318=>"000000100",
    7319=>"111111111",
    7320=>"111101111",
    7321=>"110100101",
    7322=>"011001100",
    7323=>"011110011",
    7324=>"101000000",
    7325=>"110111111",
    7326=>"100111011",
    7327=>"111111010",
    7328=>"111001010",
    7329=>"110100100",
    7330=>"011111111",
    7331=>"101101101",
    7332=>"000000000",
    7333=>"111111011",
    7334=>"010010011",
    7335=>"111000000",
    7336=>"101111111",
    7337=>"110111111",
    7338=>"101111010",
    7339=>"111101111",
    7340=>"101110111",
    7341=>"100011111",
    7342=>"100000000",
    7343=>"010011011",
    7344=>"011111111",
    7345=>"010011000",
    7346=>"011111111",
    7347=>"011010000",
    7348=>"011011011",
    7349=>"111100000",
    7350=>"000000000",
    7351=>"000010000",
    7352=>"000000000",
    7353=>"010000000",
    7354=>"010001000",
    7355=>"000000000",
    7356=>"000000000",
    7357=>"111001111",
    7358=>"110110110",
    7359=>"101001110",
    7360=>"000000000",
    7361=>"111111011",
    7362=>"000000000",
    7363=>"001000000",
    7364=>"111011110",
    7365=>"111111110",
    7366=>"111111111",
    7367=>"000010001",
    7368=>"110111011",
    7369=>"101111000",
    7370=>"101110111",
    7371=>"101000000",
    7372=>"001111110",
    7373=>"000000000",
    7374=>"010010011",
    7375=>"110010000",
    7376=>"000000000",
    7377=>"110000000",
    7378=>"101110110",
    7379=>"000000000",
    7380=>"111111011",
    7381=>"000000000",
    7382=>"111011111",
    7383=>"000010110",
    7384=>"111111100",
    7385=>"011111101",
    7386=>"011111001",
    7387=>"000000000",
    7388=>"111111011",
    7389=>"001001100",
    7390=>"110111011",
    7391=>"000000000",
    7392=>"111111111",
    7393=>"000011001",
    7394=>"000000000",
    7395=>"111110000",
    7396=>"111111110",
    7397=>"010000111",
    7398=>"110000100",
    7399=>"110011111",
    7400=>"001001000",
    7401=>"000100100",
    7402=>"111111110",
    7403=>"000010000",
    7404=>"000111111",
    7405=>"000000100",
    7406=>"111101101",
    7407=>"001101100",
    7408=>"000000000",
    7409=>"000010010",
    7410=>"111011010",
    7411=>"111000100",
    7412=>"000000000",
    7413=>"010011000",
    7414=>"000011011",
    7415=>"011111111",
    7416=>"011111111",
    7417=>"000000010",
    7418=>"100110000",
    7419=>"111111111",
    7420=>"110011000",
    7421=>"111111111",
    7422=>"011111011",
    7423=>"111111111",
    7424=>"000000001",
    7425=>"111000000",
    7426=>"010111110",
    7427=>"101101111",
    7428=>"011001011",
    7429=>"111000001",
    7430=>"000000000",
    7431=>"111111111",
    7432=>"000001000",
    7433=>"001011011",
    7434=>"100110110",
    7435=>"000100010",
    7436=>"110100110",
    7437=>"111111100",
    7438=>"000110100",
    7439=>"110111111",
    7440=>"000001011",
    7441=>"101000000",
    7442=>"100110110",
    7443=>"000100111",
    7444=>"000001001",
    7445=>"000000000",
    7446=>"000100111",
    7447=>"111111001",
    7448=>"011011111",
    7449=>"000011111",
    7450=>"011011011",
    7451=>"101000111",
    7452=>"010100110",
    7453=>"111111000",
    7454=>"110111110",
    7455=>"111111111",
    7456=>"011100100",
    7457=>"000000110",
    7458=>"100100110",
    7459=>"001000000",
    7460=>"000000111",
    7461=>"101001001",
    7462=>"111111001",
    7463=>"000000001",
    7464=>"100000000",
    7465=>"001001011",
    7466=>"101111111",
    7467=>"101100101",
    7468=>"111011001",
    7469=>"111000000",
    7470=>"111001001",
    7471=>"110111110",
    7472=>"000101111",
    7473=>"100110110",
    7474=>"001001011",
    7475=>"111010001",
    7476=>"111011000",
    7477=>"100101001",
    7478=>"111100000",
    7479=>"001000000",
    7480=>"111111111",
    7481=>"111111101",
    7482=>"100100110",
    7483=>"000000000",
    7484=>"110000000",
    7485=>"101101111",
    7486=>"111111011",
    7487=>"001101001",
    7488=>"110110010",
    7489=>"000000000",
    7490=>"111101101",
    7491=>"000000001",
    7492=>"101110111",
    7493=>"001000001",
    7494=>"101100111",
    7495=>"001000000",
    7496=>"000000111",
    7497=>"111001000",
    7498=>"000000111",
    7499=>"000010111",
    7500=>"110010000",
    7501=>"110111111",
    7502=>"010010111",
    7503=>"110010110",
    7504=>"111110101",
    7505=>"000001000",
    7506=>"111001001",
    7507=>"100010000",
    7508=>"000000100",
    7509=>"001000001",
    7510=>"000000000",
    7511=>"111001111",
    7512=>"000100110",
    7513=>"001000001",
    7514=>"111110110",
    7515=>"000000111",
    7516=>"001000100",
    7517=>"000111110",
    7518=>"100110110",
    7519=>"111000001",
    7520=>"101000000",
    7521=>"101100000",
    7522=>"110110110",
    7523=>"000000000",
    7524=>"000000000",
    7525=>"000010010",
    7526=>"101000000",
    7527=>"000110100",
    7528=>"110100001",
    7529=>"110111111",
    7530=>"101001111",
    7531=>"110111000",
    7532=>"110000110",
    7533=>"110000100",
    7534=>"001001101",
    7535=>"000010010",
    7536=>"000110110",
    7537=>"011011011",
    7538=>"010111111",
    7539=>"010010010",
    7540=>"111111001",
    7541=>"000100111",
    7542=>"001001000",
    7543=>"000000100",
    7544=>"111101100",
    7545=>"101000000",
    7546=>"011011111",
    7547=>"111111111",
    7548=>"111011001",
    7549=>"111111001",
    7550=>"001000110",
    7551=>"101001100",
    7552=>"011111111",
    7553=>"000111000",
    7554=>"101000011",
    7555=>"110100100",
    7556=>"110011000",
    7557=>"000000100",
    7558=>"010111100",
    7559=>"001000100",
    7560=>"000001000",
    7561=>"100001000",
    7562=>"011000111",
    7563=>"100011101",
    7564=>"100110000",
    7565=>"000110000",
    7566=>"000011000",
    7567=>"000001011",
    7568=>"110111001",
    7569=>"100000111",
    7570=>"111111111",
    7571=>"011000111",
    7572=>"000000000",
    7573=>"010000000",
    7574=>"000000111",
    7575=>"111100100",
    7576=>"111101111",
    7577=>"011110011",
    7578=>"110000110",
    7579=>"110100110",
    7580=>"111011111",
    7581=>"110111111",
    7582=>"111111111",
    7583=>"010001111",
    7584=>"011001000",
    7585=>"000011011",
    7586=>"000000000",
    7587=>"000000011",
    7588=>"101101101",
    7589=>"111001100",
    7590=>"011000000",
    7591=>"111000011",
    7592=>"001000000",
    7593=>"101001110",
    7594=>"100011111",
    7595=>"111110011",
    7596=>"011000101",
    7597=>"101000000",
    7598=>"000000000",
    7599=>"010000000",
    7600=>"100111101",
    7601=>"001000001",
    7602=>"001111111",
    7603=>"111100111",
    7604=>"000111000",
    7605=>"101010000",
    7606=>"000111011",
    7607=>"111000111",
    7608=>"010000010",
    7609=>"111000100",
    7610=>"111000000",
    7611=>"001010000",
    7612=>"010010000",
    7613=>"000001110",
    7614=>"001001111",
    7615=>"101110000",
    7616=>"100111110",
    7617=>"000000000",
    7618=>"000111111",
    7619=>"100110000",
    7620=>"100100001",
    7621=>"000000001",
    7622=>"000001000",
    7623=>"111111000",
    7624=>"010111000",
    7625=>"001110000",
    7626=>"011000000",
    7627=>"111000111",
    7628=>"000000000",
    7629=>"111111111",
    7630=>"000000011",
    7631=>"011000000",
    7632=>"000000111",
    7633=>"100000000",
    7634=>"111111000",
    7635=>"001101111",
    7636=>"000000001",
    7637=>"100100000",
    7638=>"000000000",
    7639=>"111001000",
    7640=>"111101111",
    7641=>"000000000",
    7642=>"110000110",
    7643=>"111000110",
    7644=>"111011011",
    7645=>"001000111",
    7646=>"011010011",
    7647=>"110101110",
    7648=>"000101000",
    7649=>"011011110",
    7650=>"011111001",
    7651=>"000001111",
    7652=>"101000010",
    7653=>"000010000",
    7654=>"011000000",
    7655=>"111110101",
    7656=>"011111100",
    7657=>"111000000",
    7658=>"010000111",
    7659=>"101000100",
    7660=>"000110110",
    7661=>"010001000",
    7662=>"111111100",
    7663=>"011100110",
    7664=>"111000101",
    7665=>"011000011",
    7666=>"010000000",
    7667=>"010111000",
    7668=>"000111110",
    7669=>"111010001",
    7670=>"000000000",
    7671=>"100011111",
    7672=>"101000111",
    7673=>"000111111",
    7674=>"100111001",
    7675=>"000111110",
    7676=>"111000011",
    7677=>"010110000",
    7678=>"100101101",
    7679=>"011000000",
    7680=>"110111100",
    7681=>"000010000",
    7682=>"010111111",
    7683=>"011001111",
    7684=>"000110011",
    7685=>"110100111",
    7686=>"110111001",
    7687=>"100000100",
    7688=>"010011010",
    7689=>"111101010",
    7690=>"000100000",
    7691=>"100000000",
    7692=>"011001001",
    7693=>"111111100",
    7694=>"010011010",
    7695=>"111001101",
    7696=>"000100111",
    7697=>"110111111",
    7698=>"011000000",
    7699=>"111001000",
    7700=>"110110000",
    7701=>"111011001",
    7702=>"101110110",
    7703=>"000000011",
    7704=>"110000011",
    7705=>"000000010",
    7706=>"000110110",
    7707=>"000000100",
    7708=>"111111110",
    7709=>"111111011",
    7710=>"000110010",
    7711=>"110100100",
    7712=>"011001000",
    7713=>"000000000",
    7714=>"000001111",
    7715=>"100000001",
    7716=>"011000000",
    7717=>"010110100",
    7718=>"101011111",
    7719=>"111110010",
    7720=>"001001100",
    7721=>"000001000",
    7722=>"111111100",
    7723=>"011000000",
    7724=>"000101111",
    7725=>"000010011",
    7726=>"011000000",
    7727=>"011001111",
    7728=>"011000001",
    7729=>"100000111",
    7730=>"111101000",
    7731=>"011011000",
    7732=>"011001111",
    7733=>"000001101",
    7734=>"110100101",
    7735=>"000000000",
    7736=>"110100000",
    7737=>"100000000",
    7738=>"000000000",
    7739=>"001011101",
    7740=>"111011100",
    7741=>"000000001",
    7742=>"111111111",
    7743=>"111010000",
    7744=>"111101000",
    7745=>"000111011",
    7746=>"011000100",
    7747=>"101100100",
    7748=>"011001110",
    7749=>"110100101",
    7750=>"111100000",
    7751=>"100000100",
    7752=>"111001000",
    7753=>"001111000",
    7754=>"001000000",
    7755=>"110001000",
    7756=>"000000100",
    7757=>"000000111",
    7758=>"111111110",
    7759=>"100101111",
    7760=>"101000010",
    7761=>"111011000",
    7762=>"100100100",
    7763=>"011100111",
    7764=>"111011101",
    7765=>"100100100",
    7766=>"011000000",
    7767=>"110000100",
    7768=>"000010111",
    7769=>"100010010",
    7770=>"111110101",
    7771=>"000000110",
    7772=>"011001011",
    7773=>"000100111",
    7774=>"100111101",
    7775=>"010011001",
    7776=>"110000000",
    7777=>"011100110",
    7778=>"110111100",
    7779=>"011000000",
    7780=>"000001111",
    7781=>"011001001",
    7782=>"000101111",
    7783=>"100101010",
    7784=>"000011111",
    7785=>"000000000",
    7786=>"011000000",
    7787=>"000000000",
    7788=>"000011001",
    7789=>"000001110",
    7790=>"001011011",
    7791=>"010011111",
    7792=>"111000111",
    7793=>"001101100",
    7794=>"110110001",
    7795=>"010001011",
    7796=>"110110111",
    7797=>"000111000",
    7798=>"000110100",
    7799=>"000000111",
    7800=>"000000110",
    7801=>"110100110",
    7802=>"111010000",
    7803=>"000100100",
    7804=>"000110111",
    7805=>"100101011",
    7806=>"110010101",
    7807=>"111001000",
    7808=>"010111001",
    7809=>"000101000",
    7810=>"010000110",
    7811=>"000000010",
    7812=>"010111010",
    7813=>"110000010",
    7814=>"000110111",
    7815=>"001001111",
    7816=>"110111000",
    7817=>"100010110",
    7818=>"111000010",
    7819=>"011111010",
    7820=>"000010010",
    7821=>"111111111",
    7822=>"010011010",
    7823=>"100100011",
    7824=>"010011110",
    7825=>"010110010",
    7826=>"010011000",
    7827=>"110100110",
    7828=>"000011011",
    7829=>"010000011",
    7830=>"111101111",
    7831=>"010011010",
    7832=>"110111010",
    7833=>"110110010",
    7834=>"000111111",
    7835=>"011011111",
    7836=>"010101011",
    7837=>"010111010",
    7838=>"000111110",
    7839=>"000000010",
    7840=>"010111011",
    7841=>"000111001",
    7842=>"011111110",
    7843=>"010010010",
    7844=>"111111110",
    7845=>"000011010",
    7846=>"000001010",
    7847=>"000111000",
    7848=>"111010110",
    7849=>"010010011",
    7850=>"000111010",
    7851=>"010110100",
    7852=>"011100110",
    7853=>"010010110",
    7854=>"000000000",
    7855=>"010101010",
    7856=>"000111111",
    7857=>"001000110",
    7858=>"000010010",
    7859=>"110000011",
    7860=>"000111010",
    7861=>"000011010",
    7862=>"010000011",
    7863=>"000000001",
    7864=>"110000000",
    7865=>"010110010",
    7866=>"000000010",
    7867=>"101101111",
    7868=>"010000000",
    7869=>"111110101",
    7870=>"010111111",
    7871=>"000110011",
    7872=>"010011010",
    7873=>"000111111",
    7874=>"010110011",
    7875=>"110000000",
    7876=>"010110010",
    7877=>"000110000",
    7878=>"010010010",
    7879=>"010010010",
    7880=>"010110011",
    7881=>"000011000",
    7882=>"010001010",
    7883=>"000101010",
    7884=>"011000011",
    7885=>"010110010",
    7886=>"000010011",
    7887=>"000001010",
    7888=>"000011010",
    7889=>"010100011",
    7890=>"000111000",
    7891=>"000000000",
    7892=>"000111000",
    7893=>"000000011",
    7894=>"011011111",
    7895=>"111111111",
    7896=>"000111100",
    7897=>"111000110",
    7898=>"010011111",
    7899=>"011000010",
    7900=>"000111001",
    7901=>"000001010",
    7902=>"010011011",
    7903=>"000111000",
    7904=>"000111010",
    7905=>"110110110",
    7906=>"010010000",
    7907=>"010011010",
    7908=>"010111010",
    7909=>"010000010",
    7910=>"011011110",
    7911=>"110111011",
    7912=>"000110110",
    7913=>"111100110",
    7914=>"110111000",
    7915=>"000000010",
    7916=>"000100110",
    7917=>"101101101",
    7918=>"010110011",
    7919=>"010010110",
    7920=>"010000010",
    7921=>"000111110",
    7922=>"000111010",
    7923=>"010011010",
    7924=>"111000101",
    7925=>"101101101",
    7926=>"100111111",
    7927=>"010110111",
    7928=>"000111110",
    7929=>"000000110",
    7930=>"001011011",
    7931=>"000000111",
    7932=>"000110100",
    7933=>"000010010",
    7934=>"001000000",
    7935=>"010011010",
    7936=>"111100111",
    7937=>"111111000",
    7938=>"111111111",
    7939=>"111010000",
    7940=>"110011001",
    7941=>"110001000",
    7942=>"101111000",
    7943=>"111111111",
    7944=>"011010010",
    7945=>"110110000",
    7946=>"010010000",
    7947=>"110011000",
    7948=>"011010000",
    7949=>"000000000",
    7950=>"011111011",
    7951=>"111111111",
    7952=>"110111011",
    7953=>"000000100",
    7954=>"010110111",
    7955=>"011111000",
    7956=>"000111111",
    7957=>"010101000",
    7958=>"000000100",
    7959=>"010111111",
    7960=>"111011110",
    7961=>"110110100",
    7962=>"110110110",
    7963=>"001011011",
    7964=>"101111111",
    7965=>"011111111",
    7966=>"011011010",
    7967=>"011111111",
    7968=>"101111111",
    7969=>"111111111",
    7970=>"111011111",
    7971=>"101111100",
    7972=>"101111001",
    7973=>"010000101",
    7974=>"001011001",
    7975=>"111110111",
    7976=>"101111100",
    7977=>"111111100",
    7978=>"001111111",
    7979=>"011111111",
    7980=>"110111000",
    7981=>"001011110",
    7982=>"111111111",
    7983=>"110111111",
    7984=>"111111001",
    7985=>"000000011",
    7986=>"100111010",
    7987=>"010010000",
    7988=>"111110110",
    7989=>"111111111",
    7990=>"100111010",
    7991=>"000000000",
    7992=>"111111000",
    7993=>"111011111",
    7994=>"011011000",
    7995=>"000000000",
    7996=>"000110110",
    7997=>"111111110",
    7998=>"110110100",
    7999=>"000010001",
    8000=>"010010000",
    8001=>"000110010",
    8002=>"100111110",
    8003=>"010001000",
    8004=>"111111111",
    8005=>"001011111",
    8006=>"000111000",
    8007=>"111111000",
    8008=>"011111110",
    8009=>"111110111",
    8010=>"010111010",
    8011=>"010110011",
    8012=>"010010010",
    8013=>"100111111",
    8014=>"111111111",
    8015=>"000000111",
    8016=>"000000000",
    8017=>"111110100",
    8018=>"100111111",
    8019=>"110111111",
    8020=>"100110010",
    8021=>"000000111",
    8022=>"000111111",
    8023=>"110111000",
    8024=>"010010111",
    8025=>"010000000",
    8026=>"011011111",
    8027=>"000000000",
    8028=>"111111110",
    8029=>"011111111",
    8030=>"101011101",
    8031=>"010000000",
    8032=>"111111111",
    8033=>"100000111",
    8034=>"001000000",
    8035=>"010010000",
    8036=>"111111010",
    8037=>"111110010",
    8038=>"111111101",
    8039=>"010111000",
    8040=>"111111101",
    8041=>"111111110",
    8042=>"111111110",
    8043=>"010110000",
    8044=>"111001111",
    8045=>"000111010",
    8046=>"001010000",
    8047=>"110110110",
    8048=>"000000111",
    8049=>"110010101",
    8050=>"111111111",
    8051=>"000000100",
    8052=>"000000111",
    8053=>"001111111",
    8054=>"110111111",
    8055=>"001011010",
    8056=>"110111010",
    8057=>"000111111",
    8058=>"111111100",
    8059=>"000111111",
    8060=>"110110111",
    8061=>"000110011",
    8062=>"000010000",
    8063=>"000010110",
    8064=>"100111001",
    8065=>"000111100",
    8066=>"000100010",
    8067=>"001000000",
    8068=>"001000001",
    8069=>"001000011",
    8070=>"101100100",
    8071=>"101001101",
    8072=>"111111101",
    8073=>"100101111",
    8074=>"000000000",
    8075=>"001011001",
    8076=>"010010010",
    8077=>"100110110",
    8078=>"101000001",
    8079=>"111110001",
    8080=>"111010000",
    8081=>"000000111",
    8082=>"010001000",
    8083=>"111000001",
    8084=>"100010010",
    8085=>"001000100",
    8086=>"011010011",
    8087=>"011000000",
    8088=>"001001001",
    8089=>"100000000",
    8090=>"111101100",
    8091=>"010000010",
    8092=>"111011110",
    8093=>"000011011",
    8094=>"000000111",
    8095=>"010011011",
    8096=>"110000000",
    8097=>"111000000",
    8098=>"011100100",
    8099=>"011001001",
    8100=>"010011011",
    8101=>"001011000",
    8102=>"011011111",
    8103=>"011001011",
    8104=>"011010010",
    8105=>"111011111",
    8106=>"100100100",
    8107=>"100100000",
    8108=>"000001111",
    8109=>"011011011",
    8110=>"101010010",
    8111=>"111100101",
    8112=>"000100100",
    8113=>"110110110",
    8114=>"001000111",
    8115=>"111010000",
    8116=>"100101111",
    8117=>"001000000",
    8118=>"100100100",
    8119=>"100000001",
    8120=>"000001011",
    8121=>"110100111",
    8122=>"000000011",
    8123=>"100100000",
    8124=>"000001101",
    8125=>"000100100",
    8126=>"100100000",
    8127=>"000011001",
    8128=>"111000110",
    8129=>"100010001",
    8130=>"011001011",
    8131=>"111010000",
    8132=>"111000010",
    8133=>"100110000",
    8134=>"110011001",
    8135=>"110011011",
    8136=>"000100111",
    8137=>"111001100",
    8138=>"001000110",
    8139=>"111001111",
    8140=>"001011111",
    8141=>"111001000",
    8142=>"011011011",
    8143=>"011110010",
    8144=>"011001001",
    8145=>"110010000",
    8146=>"100001110",
    8147=>"000001011",
    8148=>"110111001",
    8149=>"011001001",
    8150=>"110110110",
    8151=>"001011111",
    8152=>"001001101",
    8153=>"110110110",
    8154=>"111001000",
    8155=>"011011011",
    8156=>"100100001",
    8157=>"011001000",
    8158=>"100000000",
    8159=>"000111001",
    8160=>"000000000",
    8161=>"000101111",
    8162=>"111111110",
    8163=>"011010000",
    8164=>"001001011",
    8165=>"110110011",
    8166=>"001100100",
    8167=>"100001001",
    8168=>"011101010",
    8169=>"100100100",
    8170=>"001000000",
    8171=>"011011111",
    8172=>"100110100",
    8173=>"011011011",
    8174=>"010011011",
    8175=>"000001001",
    8176=>"000010011",
    8177=>"001100110",
    8178=>"000010110",
    8179=>"001001001",
    8180=>"111100110",
    8181=>"000001100",
    8182=>"011001001",
    8183=>"011011001",
    8184=>"110001101",
    8185=>"011001001",
    8186=>"000011111",
    8187=>"100100100",
    8188=>"100100100",
    8189=>"011001001",
    8190=>"111100000",
    8191=>"100111111",
    8192=>"111011000",
    8193=>"000100111",
    8194=>"001101111",
    8195=>"000000010",
    8196=>"110100100",
    8197=>"111101111",
    8198=>"111110001",
    8199=>"000111110",
    8200=>"011001110",
    8201=>"000000001",
    8202=>"000111111",
    8203=>"000110111",
    8204=>"001101111",
    8205=>"000000110",
    8206=>"011011000",
    8207=>"010011000",
    8208=>"000100111",
    8209=>"000000000",
    8210=>"110101000",
    8211=>"111011000",
    8212=>"011000000",
    8213=>"111010000",
    8214=>"011101000",
    8215=>"111110000",
    8216=>"111100000",
    8217=>"001011111",
    8218=>"100000000",
    8219=>"000000000",
    8220=>"010000000",
    8221=>"111111000",
    8222=>"001101000",
    8223=>"111111000",
    8224=>"110101101",
    8225=>"100100110",
    8226=>"100100110",
    8227=>"000010001",
    8228=>"010010000",
    8229=>"110110000",
    8230=>"100111111",
    8231=>"111000000",
    8232=>"111111000",
    8233=>"100111010",
    8234=>"101000001",
    8235=>"011011000",
    8236=>"111110100",
    8237=>"000010000",
    8238=>"010000000",
    8239=>"101111110",
    8240=>"000100101",
    8241=>"000100110",
    8242=>"000100001",
    8243=>"011010000",
    8244=>"001001001",
    8245=>"000000000",
    8246=>"000000111",
    8247=>"111110100",
    8248=>"011010001",
    8249=>"100100000",
    8250=>"010000100",
    8251=>"001000111",
    8252=>"000110000",
    8253=>"111111100",
    8254=>"011000000",
    8255=>"111011000",
    8256=>"010010000",
    8257=>"000101111",
    8258=>"010000000",
    8259=>"111111001",
    8260=>"111111000",
    8261=>"011110100",
    8262=>"111111100",
    8263=>"010111111",
    8264=>"000001011",
    8265=>"111111101",
    8266=>"100110010",
    8267=>"001000000",
    8268=>"100110010",
    8269=>"111010000",
    8270=>"110010000",
    8271=>"000000110",
    8272=>"100100100",
    8273=>"101001000",
    8274=>"000101100",
    8275=>"010011000",
    8276=>"111111000",
    8277=>"010000111",
    8278=>"111000000",
    8279=>"001111101",
    8280=>"011000000",
    8281=>"010000101",
    8282=>"001000100",
    8283=>"010010000",
    8284=>"100001001",
    8285=>"011110100",
    8286=>"000000110",
    8287=>"100010000",
    8288=>"110100000",
    8289=>"110011011",
    8290=>"111111110",
    8291=>"000010010",
    8292=>"001101000",
    8293=>"101111110",
    8294=>"101100100",
    8295=>"011011111",
    8296=>"100101111",
    8297=>"000000010",
    8298=>"111001001",
    8299=>"000000110",
    8300=>"111000111",
    8301=>"001111110",
    8302=>"110110000",
    8303=>"111110000",
    8304=>"011010000",
    8305=>"000000000",
    8306=>"000000000",
    8307=>"000101111",
    8308=>"111010000",
    8309=>"000101100",
    8310=>"000000000",
    8311=>"000001000",
    8312=>"000110111",
    8313=>"000111010",
    8314=>"001100111",
    8315=>"000010111",
    8316=>"111001000",
    8317=>"000011101",
    8318=>"001101011",
    8319=>"010000001",
    8320=>"111111010",
    8321=>"000010010",
    8322=>"111100000",
    8323=>"111101111",
    8324=>"001001000",
    8325=>"101110000",
    8326=>"000101101",
    8327=>"000111011",
    8328=>"110001001",
    8329=>"111111001",
    8330=>"101000000",
    8331=>"001001001",
    8332=>"000100101",
    8333=>"010101010",
    8334=>"110100000",
    8335=>"110110110",
    8336=>"001001001",
    8337=>"110111010",
    8338=>"000000000",
    8339=>"000110111",
    8340=>"000000011",
    8341=>"000000110",
    8342=>"000000000",
    8343=>"111111011",
    8344=>"000000000",
    8345=>"000100011",
    8346=>"001000000",
    8347=>"000000001",
    8348=>"011110000",
    8349=>"000100000",
    8350=>"001001000",
    8351=>"011011111",
    8352=>"111000000",
    8353=>"010110100",
    8354=>"110110010",
    8355=>"000100110",
    8356=>"111000101",
    8357=>"110100011",
    8358=>"000001101",
    8359=>"111000000",
    8360=>"001011001",
    8361=>"110101000",
    8362=>"000000100",
    8363=>"101100100",
    8364=>"001011000",
    8365=>"011111011",
    8366=>"001011110",
    8367=>"100111001",
    8368=>"001111111",
    8369=>"111000010",
    8370=>"000001001",
    8371=>"111100100",
    8372=>"011001001",
    8373=>"000000001",
    8374=>"010110000",
    8375=>"000001110",
    8376=>"111110110",
    8377=>"000111000",
    8378=>"110100100",
    8379=>"010000000",
    8380=>"000010011",
    8381=>"000000000",
    8382=>"000100001",
    8383=>"000111100",
    8384=>"011111001",
    8385=>"101010111",
    8386=>"011111001",
    8387=>"111111010",
    8388=>"000100100",
    8389=>"110110110",
    8390=>"000010000",
    8391=>"110111000",
    8392=>"000110110",
    8393=>"101000100",
    8394=>"011111010",
    8395=>"011000000",
    8396=>"100000111",
    8397=>"111100010",
    8398=>"011010111",
    8399=>"111000000",
    8400=>"110010110",
    8401=>"101100111",
    8402=>"001000000",
    8403=>"111111000",
    8404=>"101110011",
    8405=>"110111111",
    8406=>"000000000",
    8407=>"101000000",
    8408=>"000001100",
    8409=>"101111111",
    8410=>"000001001",
    8411=>"111101111",
    8412=>"000100000",
    8413=>"001011011",
    8414=>"011011011",
    8415=>"000001111",
    8416=>"011000100",
    8417=>"001100100",
    8418=>"111111000",
    8419=>"001111100",
    8420=>"111111011",
    8421=>"000001101",
    8422=>"111100000",
    8423=>"001111111",
    8424=>"110110110",
    8425=>"100100010",
    8426=>"100100100",
    8427=>"111111111",
    8428=>"101001000",
    8429=>"001000011",
    8430=>"000100000",
    8431=>"011001000",
    8432=>"100100100",
    8433=>"111111111",
    8434=>"111111010",
    8435=>"100100110",
    8436=>"101010011",
    8437=>"001100000",
    8438=>"111010010",
    8439=>"100100100",
    8440=>"010011011",
    8441=>"110111010",
    8442=>"001011011",
    8443=>"000111011",
    8444=>"110000001",
    8445=>"010111011",
    8446=>"100111111",
    8447=>"011001000",
    8448=>"100101111",
    8449=>"101001101",
    8450=>"000111010",
    8451=>"000011011",
    8452=>"100110111",
    8453=>"100110110",
    8454=>"101111111",
    8455=>"101000000",
    8456=>"000110110",
    8457=>"110100100",
    8458=>"010001001",
    8459=>"011000110",
    8460=>"000000100",
    8461=>"000000111",
    8462=>"100111011",
    8463=>"111100101",
    8464=>"000100110",
    8465=>"110110111",
    8466=>"010101000",
    8467=>"011111111",
    8468=>"000000000",
    8469=>"000000000",
    8470=>"101000111",
    8471=>"011111111",
    8472=>"001001000",
    8473=>"110100101",
    8474=>"111111100",
    8475=>"001011110",
    8476=>"001001001",
    8477=>"110111111",
    8478=>"000110111",
    8479=>"000000000",
    8480=>"000100000",
    8481=>"000001000",
    8482=>"011001001",
    8483=>"010111101",
    8484=>"000010001",
    8485=>"111101000",
    8486=>"000110111",
    8487=>"000110110",
    8488=>"000000000",
    8489=>"110000001",
    8490=>"000000111",
    8491=>"000110011",
    8492=>"110111010",
    8493=>"010111110",
    8494=>"000010111",
    8495=>"111111111",
    8496=>"010110111",
    8497=>"001010110",
    8498=>"011000000",
    8499=>"000010111",
    8500=>"011011110",
    8501=>"000000000",
    8502=>"000000000",
    8503=>"000110010",
    8504=>"010000000",
    8505=>"011111111",
    8506=>"011011000",
    8507=>"000000000",
    8508=>"000000000",
    8509=>"101000000",
    8510=>"100010111",
    8511=>"010110111",
    8512=>"000000111",
    8513=>"000011110",
    8514=>"110000000",
    8515=>"000000000",
    8516=>"010011011",
    8517=>"000011000",
    8518=>"010010000",
    8519=>"010111110",
    8520=>"000000111",
    8521=>"001000111",
    8522=>"111100100",
    8523=>"110000000",
    8524=>"000000000",
    8525=>"000110111",
    8526=>"110000000",
    8527=>"000000010",
    8528=>"010010110",
    8529=>"110100000",
    8530=>"110101000",
    8531=>"000010111",
    8532=>"000110110",
    8533=>"001000101",
    8534=>"110101000",
    8535=>"000111110",
    8536=>"011001100",
    8537=>"111011111",
    8538=>"100001000",
    8539=>"000111111",
    8540=>"001111100",
    8541=>"110011000",
    8542=>"001001111",
    8543=>"111111000",
    8544=>"010011111",
    8545=>"000111111",
    8546=>"000000000",
    8547=>"111111000",
    8548=>"111010110",
    8549=>"010010010",
    8550=>"010000000",
    8551=>"010111110",
    8552=>"001000001",
    8553=>"101000000",
    8554=>"111111001",
    8555=>"000111111",
    8556=>"000000110",
    8557=>"111101000",
    8558=>"111000000",
    8559=>"001011011",
    8560=>"111110000",
    8561=>"111111111",
    8562=>"000000110",
    8563=>"010110111",
    8564=>"101101101",
    8565=>"010010000",
    8566=>"001001000",
    8567=>"110100110",
    8568=>"110111101",
    8569=>"111110000",
    8570=>"100100000",
    8571=>"001000001",
    8572=>"000100100",
    8573=>"101111111",
    8574=>"010000000",
    8575=>"110001010",
    8576=>"000000001",
    8577=>"101100100",
    8578=>"001011111",
    8579=>"010001010",
    8580=>"111111111",
    8581=>"000010000",
    8582=>"001000110",
    8583=>"001110100",
    8584=>"101100100",
    8585=>"110111111",
    8586=>"011001100",
    8587=>"111111110",
    8588=>"100010000",
    8589=>"110111000",
    8590=>"000000000",
    8591=>"000000100",
    8592=>"000000100",
    8593=>"000000100",
    8594=>"011001010",
    8595=>"000000000",
    8596=>"110001001",
    8597=>"001000100",
    8598=>"000000000",
    8599=>"110110000",
    8600=>"000000000",
    8601=>"000000000",
    8602=>"000100110",
    8603=>"111111001",
    8604=>"000000010",
    8605=>"000001100",
    8606=>"111111110",
    8607=>"110110000",
    8608=>"011101111",
    8609=>"000000000",
    8610=>"111111111",
    8611=>"100000011",
    8612=>"110011011",
    8613=>"100111100",
    8614=>"110110110",
    8615=>"110110110",
    8616=>"110011101",
    8617=>"000000000",
    8618=>"000000001",
    8619=>"000001000",
    8620=>"111111111",
    8621=>"110010110",
    8622=>"111001110",
    8623=>"111111100",
    8624=>"000011001",
    8625=>"110111101",
    8626=>"111111110",
    8627=>"000000100",
    8628=>"000011011",
    8629=>"000001011",
    8630=>"010001101",
    8631=>"001001101",
    8632=>"001000000",
    8633=>"110000000",
    8634=>"000000000",
    8635=>"000010000",
    8636=>"001100110",
    8637=>"000000101",
    8638=>"000000000",
    8639=>"011011001",
    8640=>"011000100",
    8641=>"000000100",
    8642=>"100111000",
    8643=>"100101000",
    8644=>"111111111",
    8645=>"100011011",
    8646=>"100000011",
    8647=>"001100000",
    8648=>"110111010",
    8649=>"000000001",
    8650=>"111110011",
    8651=>"101100111",
    8652=>"110111000",
    8653=>"000000001",
    8654=>"110100110",
    8655=>"000110110",
    8656=>"110110010",
    8657=>"001100111",
    8658=>"001000010",
    8659=>"000001101",
    8660=>"011111001",
    8661=>"110111000",
    8662=>"000011000",
    8663=>"001010000",
    8664=>"111111111",
    8665=>"100111011",
    8666=>"000000000",
    8667=>"010111100",
    8668=>"000000010",
    8669=>"111101101",
    8670=>"000000100",
    8671=>"000001011",
    8672=>"110110010",
    8673=>"110011011",
    8674=>"000111011",
    8675=>"000100000",
    8676=>"101011100",
    8677=>"000110111",
    8678=>"010011001",
    8679=>"111101100",
    8680=>"001101101",
    8681=>"001000110",
    8682=>"000000100",
    8683=>"010110011",
    8684=>"001000001",
    8685=>"011000000",
    8686=>"000001010",
    8687=>"110111011",
    8688=>"011011111",
    8689=>"110111111",
    8690=>"100110100",
    8691=>"000001010",
    8692=>"111011001",
    8693=>"001000110",
    8694=>"100100100",
    8695=>"000100101",
    8696=>"111111111",
    8697=>"100000000",
    8698=>"110110000",
    8699=>"011001110",
    8700=>"100110110",
    8701=>"110110110",
    8702=>"110000000",
    8703=>"010010010",
    8704=>"101001001",
    8705=>"000000000",
    8706=>"010111010",
    8707=>"111111111",
    8708=>"001001001",
    8709=>"010000000",
    8710=>"111111111",
    8711=>"001000101",
    8712=>"100110111",
    8713=>"001001101",
    8714=>"001000001",
    8715=>"001000110",
    8716=>"000000000",
    8717=>"111111100",
    8718=>"010000000",
    8719=>"011111011",
    8720=>"111111111",
    8721=>"010101111",
    8722=>"111111011",
    8723=>"110110100",
    8724=>"000111110",
    8725=>"000000001",
    8726=>"110000000",
    8727=>"101000000",
    8728=>"111111111",
    8729=>"101001010",
    8730=>"101001001",
    8731=>"111101110",
    8732=>"111111111",
    8733=>"000000001",
    8734=>"111110110",
    8735=>"111000000",
    8736=>"111111000",
    8737=>"111111010",
    8738=>"001101110",
    8739=>"000000000",
    8740=>"111101100",
    8741=>"001111010",
    8742=>"010110110",
    8743=>"000000000",
    8744=>"111101111",
    8745=>"001001101",
    8746=>"000001000",
    8747=>"111110110",
    8748=>"111000101",
    8749=>"000000011",
    8750=>"100001101",
    8751=>"111111111",
    8752=>"000000010",
    8753=>"000110110",
    8754=>"000000000",
    8755=>"110111011",
    8756=>"000000100",
    8757=>"000000110",
    8758=>"001111101",
    8759=>"000010010",
    8760=>"000000000",
    8761=>"111111101",
    8762=>"000000111",
    8763=>"011010010",
    8764=>"000000000",
    8765=>"000001000",
    8766=>"111100000",
    8767=>"000000110",
    8768=>"000100101",
    8769=>"011000000",
    8770=>"100000001",
    8771=>"000000000",
    8772=>"010101110",
    8773=>"001001001",
    8774=>"101000100",
    8775=>"110111111",
    8776=>"110011011",
    8777=>"000000001",
    8778=>"111000000",
    8779=>"000000000",
    8780=>"000000000",
    8781=>"111000000",
    8782=>"010000001",
    8783=>"010111010",
    8784=>"000010000",
    8785=>"001001001",
    8786=>"100100111",
    8787=>"011011101",
    8788=>"100100100",
    8789=>"000000000",
    8790=>"111101000",
    8791=>"111011111",
    8792=>"100100100",
    8793=>"101001111",
    8794=>"100000001",
    8795=>"110111110",
    8796=>"010011011",
    8797=>"010110000",
    8798=>"111010110",
    8799=>"000000000",
    8800=>"001111111",
    8801=>"011111111",
    8802=>"000010000",
    8803=>"000111111",
    8804=>"010111111",
    8805=>"111000001",
    8806=>"000100000",
    8807=>"111110000",
    8808=>"001000000",
    8809=>"101111111",
    8810=>"101100101",
    8811=>"000000111",
    8812=>"010111010",
    8813=>"000000000",
    8814=>"111111111",
    8815=>"011011001",
    8816=>"010111000",
    8817=>"000001100",
    8818=>"111111101",
    8819=>"000110000",
    8820=>"111000000",
    8821=>"011100101",
    8822=>"000001001",
    8823=>"010000000",
    8824=>"000100110",
    8825=>"111010000",
    8826=>"001000000",
    8827=>"010111111",
    8828=>"000000101",
    8829=>"111000000",
    8830=>"101001100",
    8831=>"010001110",
    8832=>"011111111",
    8833=>"101100100",
    8834=>"010010000",
    8835=>"011101111",
    8836=>"001011110",
    8837=>"111111000",
    8838=>"111110000",
    8839=>"101101111",
    8840=>"111010101",
    8841=>"110100111",
    8842=>"101001101",
    8843=>"100001011",
    8844=>"000000000",
    8845=>"110111010",
    8846=>"111000110",
    8847=>"000000000",
    8848=>"000000110",
    8849=>"000000111",
    8850=>"111000101",
    8851=>"111011100",
    8852=>"111101111",
    8853=>"101101000",
    8854=>"001000000",
    8855=>"000000010",
    8856=>"100001001",
    8857=>"000111111",
    8858=>"111100001",
    8859=>"011100001",
    8860=>"000111010",
    8861=>"011100101",
    8862=>"011111100",
    8863=>"111111011",
    8864=>"110000111",
    8865=>"110100000",
    8866=>"110110001",
    8867=>"000100001",
    8868=>"000000000",
    8869=>"000101110",
    8870=>"100010010",
    8871=>"101000101",
    8872=>"001111001",
    8873=>"101111111",
    8874=>"000110110",
    8875=>"011011000",
    8876=>"000110111",
    8877=>"000100101",
    8878=>"111000010",
    8879=>"101100111",
    8880=>"000000111",
    8881=>"111010000",
    8882=>"000101011",
    8883=>"000000111",
    8884=>"001111111",
    8885=>"001101001",
    8886=>"101000000",
    8887=>"010010000",
    8888=>"001100000",
    8889=>"111111110",
    8890=>"011000101",
    8891=>"000000000",
    8892=>"101001000",
    8893=>"111111010",
    8894=>"111000000",
    8895=>"100111001",
    8896=>"100101111",
    8897=>"000100100",
    8898=>"000100111",
    8899=>"000000000",
    8900=>"101100111",
    8901=>"011010100",
    8902=>"111000110",
    8903=>"001101101",
    8904=>"100000111",
    8905=>"000111111",
    8906=>"000001010",
    8907=>"001101101",
    8908=>"010000000",
    8909=>"111110000",
    8910=>"010011010",
    8911=>"101000111",
    8912=>"000100111",
    8913=>"000000101",
    8914=>"000101110",
    8915=>"000011010",
    8916=>"110010001",
    8917=>"000001000",
    8918=>"010111011",
    8919=>"111000001",
    8920=>"110111011",
    8921=>"111000001",
    8922=>"101001000",
    8923=>"111000110",
    8924=>"110110000",
    8925=>"001000001",
    8926=>"001100000",
    8927=>"010000000",
    8928=>"111111101",
    8929=>"100000001",
    8930=>"111011000",
    8931=>"000010111",
    8932=>"110111110",
    8933=>"101000101",
    8934=>"000000000",
    8935=>"101100101",
    8936=>"001100001",
    8937=>"100101100",
    8938=>"111101101",
    8939=>"010000101",
    8940=>"101010000",
    8941=>"111101100",
    8942=>"000010100",
    8943=>"110011001",
    8944=>"010100000",
    8945=>"111001100",
    8946=>"111000101",
    8947=>"000100111",
    8948=>"001101000",
    8949=>"101101100",
    8950=>"101001000",
    8951=>"000100110",
    8952=>"011001001",
    8953=>"101101100",
    8954=>"100001100",
    8955=>"101000000",
    8956=>"110010000",
    8957=>"101100111",
    8958=>"111111010",
    8959=>"111011010",
    8960=>"010010110",
    8961=>"000011000",
    8962=>"101000010",
    8963=>"100100000",
    8964=>"010001000",
    8965=>"010111111",
    8966=>"101111111",
    8967=>"000011000",
    8968=>"110001111",
    8969=>"111101001",
    8970=>"001000000",
    8971=>"001000000",
    8972=>"000000000",
    8973=>"010111010",
    8974=>"100100000",
    8975=>"000010010",
    8976=>"100000110",
    8977=>"111111111",
    8978=>"111110111",
    8979=>"000000010",
    8980=>"111111000",
    8981=>"000000000",
    8982=>"000000000",
    8983=>"110100110",
    8984=>"101001001",
    8985=>"110000000",
    8986=>"011011100",
    8987=>"000010001",
    8988=>"111111101",
    8989=>"111110111",
    8990=>"111110111",
    8991=>"100000000",
    8992=>"010000001",
    8993=>"000001001",
    8994=>"011111010",
    8995=>"100000000",
    8996=>"101100111",
    8997=>"000000000",
    8998=>"100111011",
    8999=>"000000100",
    9000=>"000000010",
    9001=>"100000001",
    9002=>"001110100",
    9003=>"001011011",
    9004=>"100110111",
    9005=>"111111111",
    9006=>"000000000",
    9007=>"111111111",
    9008=>"100101111",
    9009=>"000000000",
    9010=>"100000011",
    9011=>"110001011",
    9012=>"111001001",
    9013=>"111101111",
    9014=>"111111111",
    9015=>"101111011",
    9016=>"111001000",
    9017=>"100101111",
    9018=>"000100111",
    9019=>"111110010",
    9020=>"000010000",
    9021=>"000010000",
    9022=>"001100111",
    9023=>"011011000",
    9024=>"011111111",
    9025=>"010100111",
    9026=>"111001001",
    9027=>"111111111",
    9028=>"001001001",
    9029=>"110100110",
    9030=>"000010000",
    9031=>"010000000",
    9032=>"110100000",
    9033=>"000100111",
    9034=>"000110111",
    9035=>"010011000",
    9036=>"010000101",
    9037=>"000000000",
    9038=>"110101010",
    9039=>"101100111",
    9040=>"101101111",
    9041=>"000010100",
    9042=>"000010011",
    9043=>"101001011",
    9044=>"001000011",
    9045=>"000010010",
    9046=>"000000000",
    9047=>"111111111",
    9048=>"101000111",
    9049=>"000001110",
    9050=>"000000010",
    9051=>"000010100",
    9052=>"100111000",
    9053=>"010011000",
    9054=>"101111100",
    9055=>"000000001",
    9056=>"100100001",
    9057=>"100100110",
    9058=>"111101111",
    9059=>"000111001",
    9060=>"000001111",
    9061=>"010100000",
    9062=>"000000000",
    9063=>"111111111",
    9064=>"111111111",
    9065=>"000010010",
    9066=>"111101101",
    9067=>"010111011",
    9068=>"100000001",
    9069=>"000010011",
    9070=>"000111111",
    9071=>"011001001",
    9072=>"000010000",
    9073=>"000101000",
    9074=>"100100101",
    9075=>"011011000",
    9076=>"000010110",
    9077=>"100000101",
    9078=>"101001111",
    9079=>"001000000",
    9080=>"111111010",
    9081=>"111000000",
    9082=>"110010100",
    9083=>"000000111",
    9084=>"011001001",
    9085=>"110000111",
    9086=>"100111111",
    9087=>"110111100",
    9088=>"000000010",
    9089=>"111000010",
    9090=>"101101111",
    9091=>"111111110",
    9092=>"001100000",
    9093=>"000000000",
    9094=>"010010010",
    9095=>"101001101",
    9096=>"000100101",
    9097=>"011000010",
    9098=>"010111110",
    9099=>"100011001",
    9100=>"101111001",
    9101=>"101101101",
    9102=>"100000111",
    9103=>"111100100",
    9104=>"000010110",
    9105=>"101101101",
    9106=>"000000111",
    9107=>"100000111",
    9108=>"000000001",
    9109=>"000000001",
    9110=>"100000000",
    9111=>"111010010",
    9112=>"000101110",
    9113=>"000110011",
    9114=>"010110110",
    9115=>"011011010",
    9116=>"010111010",
    9117=>"000000001",
    9118=>"111111001",
    9119=>"101101101",
    9120=>"000111111",
    9121=>"000011100",
    9122=>"000011011",
    9123=>"000001000",
    9124=>"000011111",
    9125=>"001101010",
    9126=>"111100001",
    9127=>"100010010",
    9128=>"010111000",
    9129=>"010110101",
    9130=>"111111001",
    9131=>"000101111",
    9132=>"001001111",
    9133=>"111101101",
    9134=>"011000000",
    9135=>"111111001",
    9136=>"110100100",
    9137=>"101101000",
    9138=>"000000101",
    9139=>"011000010",
    9140=>"000010100",
    9141=>"000110000",
    9142=>"100000000",
    9143=>"000000111",
    9144=>"111101011",
    9145=>"000010011",
    9146=>"000000011",
    9147=>"000000000",
    9148=>"101101110",
    9149=>"100000111",
    9150=>"110111010",
    9151=>"011010010",
    9152=>"010111011",
    9153=>"101100101",
    9154=>"011010100",
    9155=>"000100010",
    9156=>"000111110",
    9157=>"011010111",
    9158=>"001100110",
    9159=>"000101011",
    9160=>"000000001",
    9161=>"000111010",
    9162=>"000011011",
    9163=>"000000100",
    9164=>"101000000",
    9165=>"010111001",
    9166=>"100011010",
    9167=>"101000001",
    9168=>"001001101",
    9169=>"100000111",
    9170=>"000011101",
    9171=>"011111100",
    9172=>"100000100",
    9173=>"001101110",
    9174=>"010010010",
    9175=>"000000100",
    9176=>"001011011",
    9177=>"000000111",
    9178=>"100011001",
    9179=>"000010000",
    9180=>"000101111",
    9181=>"011000101",
    9182=>"111111001",
    9183=>"001100010",
    9184=>"001011000",
    9185=>"000000110",
    9186=>"101100111",
    9187=>"111001010",
    9188=>"010111111",
    9189=>"011000101",
    9190=>"000000111",
    9191=>"000111100",
    9192=>"000001111",
    9193=>"110111100",
    9194=>"000000110",
    9195=>"111110000",
    9196=>"101101000",
    9197=>"000011000",
    9198=>"111111100",
    9199=>"001000000",
    9200=>"101000101",
    9201=>"000000110",
    9202=>"111111111",
    9203=>"011000000",
    9204=>"101101111",
    9205=>"000000010",
    9206=>"000000100",
    9207=>"100000101",
    9208=>"010011000",
    9209=>"111000000",
    9210=>"001000111",
    9211=>"101011000",
    9212=>"001110110",
    9213=>"011010010",
    9214=>"010000000",
    9215=>"010110010",
    9216=>"001100100",
    9217=>"001001111",
    9218=>"001001111",
    9219=>"011100001",
    9220=>"101000110",
    9221=>"010110110",
    9222=>"011110110",
    9223=>"100001011",
    9224=>"011100000",
    9225=>"000110111",
    9226=>"100001011",
    9227=>"010000001",
    9228=>"011000000",
    9229=>"101000101",
    9230=>"001101000",
    9231=>"100001001",
    9232=>"000001111",
    9233=>"100010011",
    9234=>"001000101",
    9235=>"100111011",
    9236=>"000000111",
    9237=>"110010111",
    9238=>"000000000",
    9239=>"110001001",
    9240=>"001001000",
    9241=>"101101001",
    9242=>"011100100",
    9243=>"011001100",
    9244=>"011110111",
    9245=>"001101110",
    9246=>"011100000",
    9247=>"100011001",
    9248=>"110011110",
    9249=>"011111110",
    9250=>"011000011",
    9251=>"111011001",
    9252=>"010010001",
    9253=>"101100111",
    9254=>"000001101",
    9255=>"011100110",
    9256=>"110011001",
    9257=>"100011101",
    9258=>"000001001",
    9259=>"001001100",
    9260=>"110000011",
    9261=>"110000001",
    9262=>"000010010",
    9263=>"100100101",
    9264=>"100100000",
    9265=>"100100111",
    9266=>"110010011",
    9267=>"100111000",
    9268=>"011010100",
    9269=>"010000011",
    9270=>"110110011",
    9271=>"010011110",
    9272=>"001001001",
    9273=>"111010001",
    9274=>"111100000",
    9275=>"000000000",
    9276=>"011101001",
    9277=>"111111001",
    9278=>"001011111",
    9279=>"010011101",
    9280=>"101001000",
    9281=>"010011100",
    9282=>"100011001",
    9283=>"000000000",
    9284=>"100111011",
    9285=>"111110100",
    9286=>"000000100",
    9287=>"100001001",
    9288=>"100101100",
    9289=>"001000110",
    9290=>"110011011",
    9291=>"101110100",
    9292=>"100100011",
    9293=>"000001001",
    9294=>"001001001",
    9295=>"101000011",
    9296=>"000001011",
    9297=>"001101100",
    9298=>"110001001",
    9299=>"111110101",
    9300=>"001000110",
    9301=>"111100111",
    9302=>"011011000",
    9303=>"000010100",
    9304=>"001000110",
    9305=>"100110011",
    9306=>"001101110",
    9307=>"101000011",
    9308=>"001101100",
    9309=>"110000010",
    9310=>"001100110",
    9311=>"001011111",
    9312=>"000101111",
    9313=>"000010000",
    9314=>"111101011",
    9315=>"011000001",
    9316=>"110010011",
    9317=>"011101110",
    9318=>"011010110",
    9319=>"110011001",
    9320=>"110010010",
    9321=>"001001100",
    9322=>"001101100",
    9323=>"110110011",
    9324=>"011110000",
    9325=>"100101001",
    9326=>"000001000",
    9327=>"001000110",
    9328=>"110100011",
    9329=>"110000000",
    9330=>"001100110",
    9331=>"110100100",
    9332=>"111001001",
    9333=>"110110001",
    9334=>"100110011",
    9335=>"110111101",
    9336=>"110011001",
    9337=>"100100011",
    9338=>"001111101",
    9339=>"100001001",
    9340=>"011100100",
    9341=>"111001111",
    9342=>"111111011",
    9343=>"101111101",
    9344=>"110010101",
    9345=>"111110111",
    9346=>"000111010",
    9347=>"000000000",
    9348=>"011111001",
    9349=>"000000000",
    9350=>"010010010",
    9351=>"010111010",
    9352=>"110111111",
    9353=>"111101111",
    9354=>"110000001",
    9355=>"011101110",
    9356=>"000011000",
    9357=>"010110010",
    9358=>"010011011",
    9359=>"000000000",
    9360=>"110111110",
    9361=>"000000010",
    9362=>"000111111",
    9363=>"111110000",
    9364=>"000111000",
    9365=>"001000000",
    9366=>"010010000",
    9367=>"111101001",
    9368=>"011101111",
    9369=>"111101011",
    9370=>"011111111",
    9371=>"011011110",
    9372=>"101000100",
    9373=>"000111101",
    9374=>"100101110",
    9375=>"101101000",
    9376=>"000000101",
    9377=>"000100100",
    9378=>"111101111",
    9379=>"111111111",
    9380=>"001000100",
    9381=>"101010000",
    9382=>"000110111",
    9383=>"100110111",
    9384=>"111111100",
    9385=>"111011111",
    9386=>"000001000",
    9387=>"011111101",
    9388=>"101111111",
    9389=>"010110000",
    9390=>"111000100",
    9391=>"111000000",
    9392=>"111111111",
    9393=>"110110000",
    9394=>"011101100",
    9395=>"011111111",
    9396=>"110110110",
    9397=>"000000010",
    9398=>"011001000",
    9399=>"000111111",
    9400=>"000110001",
    9401=>"011101001",
    9402=>"011000011",
    9403=>"100111011",
    9404=>"110000000",
    9405=>"010001001",
    9406=>"110110001",
    9407=>"100100101",
    9408=>"100100010",
    9409=>"000111000",
    9410=>"010111011",
    9411=>"010011111",
    9412=>"101000001",
    9413=>"000011011",
    9414=>"000011110",
    9415=>"111110000",
    9416=>"011011111",
    9417=>"001000111",
    9418=>"111110110",
    9419=>"000000010",
    9420=>"111111111",
    9421=>"010000011",
    9422=>"111100101",
    9423=>"000010010",
    9424=>"011011011",
    9425=>"000111010",
    9426=>"000010010",
    9427=>"111000000",
    9428=>"000110110",
    9429=>"010111111",
    9430=>"110111111",
    9431=>"101001001",
    9432=>"001100111",
    9433=>"111111111",
    9434=>"111011011",
    9435=>"000010010",
    9436=>"110111010",
    9437=>"000010000",
    9438=>"101110000",
    9439=>"000000000",
    9440=>"011111111",
    9441=>"010111111",
    9442=>"010111010",
    9443=>"111111111",
    9444=>"111111101",
    9445=>"111000000",
    9446=>"000111010",
    9447=>"111110000",
    9448=>"110110011",
    9449=>"110000111",
    9450=>"100101111",
    9451=>"111111111",
    9452=>"000111011",
    9453=>"010010000",
    9454=>"101001001",
    9455=>"011101100",
    9456=>"111000000",
    9457=>"111110110",
    9458=>"001011000",
    9459=>"111111001",
    9460=>"110010010",
    9461=>"000000101",
    9462=>"100000110",
    9463=>"101101011",
    9464=>"101011111",
    9465=>"001010000",
    9466=>"010110100",
    9467=>"000110010",
    9468=>"100100101",
    9469=>"111111111",
    9470=>"110111001",
    9471=>"000000001",
    9472=>"010000000",
    9473=>"001111111",
    9474=>"000000000",
    9475=>"011101100",
    9476=>"111110111",
    9477=>"011001000",
    9478=>"110010010",
    9479=>"111111011",
    9480=>"111100001",
    9481=>"110010100",
    9482=>"001111010",
    9483=>"111001001",
    9484=>"000001000",
    9485=>"000011010",
    9486=>"111111111",
    9487=>"001101110",
    9488=>"000000000",
    9489=>"000010000",
    9490=>"000000000",
    9491=>"011001111",
    9492=>"001000101",
    9493=>"000001010",
    9494=>"000000000",
    9495=>"101100010",
    9496=>"100000000",
    9497=>"110100100",
    9498=>"010100100",
    9499=>"000010001",
    9500=>"011100111",
    9501=>"111100100",
    9502=>"111011011",
    9503=>"000101000",
    9504=>"010000110",
    9505=>"011110100",
    9506=>"011001101",
    9507=>"011111111",
    9508=>"000010000",
    9509=>"110111111",
    9510=>"000100111",
    9511=>"000000000",
    9512=>"111101000",
    9513=>"000000100",
    9514=>"010001011",
    9515=>"011001111",
    9516=>"100111011",
    9517=>"101111111",
    9518=>"000010010",
    9519=>"111010101",
    9520=>"011000100",
    9521=>"000010000",
    9522=>"101100110",
    9523=>"001011000",
    9524=>"111111001",
    9525=>"000000000",
    9526=>"000000111",
    9527=>"000111000",
    9528=>"101000000",
    9529=>"011111001",
    9530=>"111000000",
    9531=>"001011000",
    9532=>"010111110",
    9533=>"111111111",
    9534=>"001010110",
    9535=>"010100101",
    9536=>"000000111",
    9537=>"111111111",
    9538=>"111111111",
    9539=>"000000000",
    9540=>"010111011",
    9541=>"111110110",
    9542=>"110111111",
    9543=>"100000010",
    9544=>"000000010",
    9545=>"111001110",
    9546=>"000101011",
    9547=>"011111010",
    9548=>"111111000",
    9549=>"010011000",
    9550=>"111111111",
    9551=>"000000001",
    9552=>"101101111",
    9553=>"111111111",
    9554=>"000100000",
    9555=>"101000000",
    9556=>"111010000",
    9557=>"111111111",
    9558=>"010010010",
    9559=>"011001000",
    9560=>"001001101",
    9561=>"011010000",
    9562=>"000011011",
    9563=>"111100101",
    9564=>"111110100",
    9565=>"000110111",
    9566=>"001000001",
    9567=>"100111110",
    9568=>"000000110",
    9569=>"100100001",
    9570=>"000000000",
    9571=>"111000000",
    9572=>"111111111",
    9573=>"101100100",
    9574=>"111011011",
    9575=>"110100010",
    9576=>"010000000",
    9577=>"111101111",
    9578=>"111000111",
    9579=>"111111001",
    9580=>"011000110",
    9581=>"000000000",
    9582=>"000000001",
    9583=>"110111110",
    9584=>"000000000",
    9585=>"001000000",
    9586=>"000000000",
    9587=>"100000000",
    9588=>"000000000",
    9589=>"011000011",
    9590=>"000101111",
    9591=>"111001011",
    9592=>"111001000",
    9593=>"010000110",
    9594=>"000011001",
    9595=>"000000000",
    9596=>"000010110",
    9597=>"111111111",
    9598=>"010001101",
    9599=>"111101101",
    9600=>"001010110",
    9601=>"010010000",
    9602=>"000000101",
    9603=>"111000100",
    9604=>"011111100",
    9605=>"111111011",
    9606=>"111101111",
    9607=>"110010101",
    9608=>"011111111",
    9609=>"011001111",
    9610=>"000000000",
    9611=>"011000001",
    9612=>"010110000",
    9613=>"111111000",
    9614=>"011011100",
    9615=>"010011001",
    9616=>"110111111",
    9617=>"111111010",
    9618=>"001100010",
    9619=>"110110010",
    9620=>"011011010",
    9621=>"100101111",
    9622=>"000000000",
    9623=>"010101000",
    9624=>"000011011",
    9625=>"000000100",
    9626=>"101111100",
    9627=>"110111111",
    9628=>"111111010",
    9629=>"100011001",
    9630=>"100100100",
    9631=>"101101100",
    9632=>"110001101",
    9633=>"000000001",
    9634=>"001000000",
    9635=>"000100101",
    9636=>"110110111",
    9637=>"111111010",
    9638=>"111111110",
    9639=>"101101101",
    9640=>"000000010",
    9641=>"110101010",
    9642=>"001000000",
    9643=>"111101011",
    9644=>"011100111",
    9645=>"100100000",
    9646=>"011111110",
    9647=>"001000111",
    9648=>"110000110",
    9649=>"010010000",
    9650=>"000000101",
    9651=>"000100000",
    9652=>"100110101",
    9653=>"000000010",
    9654=>"010010100",
    9655=>"011111010",
    9656=>"101000000",
    9657=>"110101101",
    9658=>"011010001",
    9659=>"000000000",
    9660=>"101000101",
    9661=>"011111000",
    9662=>"001011111",
    9663=>"111111011",
    9664=>"100100111",
    9665=>"101001100",
    9666=>"110010010",
    9667=>"111101101",
    9668=>"000100111",
    9669=>"001111011",
    9670=>"000010010",
    9671=>"111100011",
    9672=>"110110111",
    9673=>"000000101",
    9674=>"011000111",
    9675=>"100000010",
    9676=>"100000000",
    9677=>"000000101",
    9678=>"101011011",
    9679=>"110111011",
    9680=>"010010000",
    9681=>"000010000",
    9682=>"000100101",
    9683=>"111111011",
    9684=>"110001111",
    9685=>"000000000",
    9686=>"100001011",
    9687=>"111001000",
    9688=>"110101111",
    9689=>"001001111",
    9690=>"000100111",
    9691=>"000010010",
    9692=>"001001111",
    9693=>"001101000",
    9694=>"100001100",
    9695=>"111111011",
    9696=>"100101101",
    9697=>"011011001",
    9698=>"000000101",
    9699=>"010111010",
    9700=>"101010111",
    9701=>"001010000",
    9702=>"000110000",
    9703=>"010011011",
    9704=>"111111111",
    9705=>"100000000",
    9706=>"100101011",
    9707=>"101001010",
    9708=>"010010100",
    9709=>"000101100",
    9710=>"000001111",
    9711=>"111110000",
    9712=>"001000111",
    9713=>"011001000",
    9714=>"101101000",
    9715=>"010111000",
    9716=>"111111111",
    9717=>"000000100",
    9718=>"000000000",
    9719=>"100001111",
    9720=>"000000000",
    9721=>"001000011",
    9722=>"111111001",
    9723=>"111111111",
    9724=>"000111100",
    9725=>"000000000",
    9726=>"001000101",
    9727=>"000001011",
    9728=>"010010111",
    9729=>"111111111",
    9730=>"111111111",
    9731=>"010110110",
    9732=>"000000001",
    9733=>"000000000",
    9734=>"001110111",
    9735=>"111101000",
    9736=>"111111111",
    9737=>"111111111",
    9738=>"000100010",
    9739=>"001100001",
    9740=>"110111111",
    9741=>"010110010",
    9742=>"100100100",
    9743=>"111100000",
    9744=>"011111111",
    9745=>"100000000",
    9746=>"001001000",
    9747=>"100100101",
    9748=>"110111000",
    9749=>"000101111",
    9750=>"111000111",
    9751=>"000000000",
    9752=>"100001001",
    9753=>"001000100",
    9754=>"000000011",
    9755=>"000111111",
    9756=>"000000000",
    9757=>"000000001",
    9758=>"000000010",
    9759=>"000000000",
    9760=>"000111111",
    9761=>"111000101",
    9762=>"000011011",
    9763=>"000000001",
    9764=>"111110110",
    9765=>"000000000",
    9766=>"001000000",
    9767=>"000111111",
    9768=>"111000000",
    9769=>"001001001",
    9770=>"010010111",
    9771=>"000000101",
    9772=>"001001001",
    9773=>"011010111",
    9774=>"001011111",
    9775=>"111111000",
    9776=>"011111011",
    9777=>"001011000",
    9778=>"110111111",
    9779=>"001000000",
    9780=>"000100111",
    9781=>"000001111",
    9782=>"000101111",
    9783=>"110110100",
    9784=>"100100110",
    9785=>"111000000",
    9786=>"011111010",
    9787=>"110110111",
    9788=>"001111111",
    9789=>"000000101",
    9790=>"110111111",
    9791=>"000000101",
    9792=>"010000010",
    9793=>"000000000",
    9794=>"000000000",
    9795=>"000000000",
    9796=>"111111011",
    9797=>"000110110",
    9798=>"000000101",
    9799=>"001010000",
    9800=>"110111111",
    9801=>"000000111",
    9802=>"001000111",
    9803=>"000000000",
    9804=>"111111000",
    9805=>"110111000",
    9806=>"111111111",
    9807=>"010111110",
    9808=>"000111000",
    9809=>"111100100",
    9810=>"000000101",
    9811=>"000000000",
    9812=>"010111011",
    9813=>"110110110",
    9814=>"001111111",
    9815=>"111001101",
    9816=>"000000101",
    9817=>"111111111",
    9818=>"000000000",
    9819=>"000000000",
    9820=>"100000111",
    9821=>"011101111",
    9822=>"111011111",
    9823=>"101000000",
    9824=>"000100101",
    9825=>"000011011",
    9826=>"111111111",
    9827=>"000000100",
    9828=>"000000000",
    9829=>"100111010",
    9830=>"111001011",
    9831=>"101000000",
    9832=>"011111111",
    9833=>"111100000",
    9834=>"000000111",
    9835=>"011010011",
    9836=>"000000010",
    9837=>"111111111",
    9838=>"000000000",
    9839=>"001001001",
    9840=>"111111001",
    9841=>"000000000",
    9842=>"000111111",
    9843=>"000000000",
    9844=>"111100000",
    9845=>"100000011",
    9846=>"111000110",
    9847=>"010000000",
    9848=>"001000001",
    9849=>"000111111",
    9850=>"111111111",
    9851=>"111111111",
    9852=>"000101100",
    9853=>"000000000",
    9854=>"000000000",
    9855=>"000000000",
    9856=>"000111000",
    9857=>"100100000",
    9858=>"011111111",
    9859=>"110110110",
    9860=>"001100101",
    9861=>"110110110",
    9862=>"000000000",
    9863=>"000001100",
    9864=>"111111111",
    9865=>"000010111",
    9866=>"011111111",
    9867=>"011001000",
    9868=>"010110100",
    9869=>"010011000",
    9870=>"011001001",
    9871=>"100100111",
    9872=>"010010011",
    9873=>"000001001",
    9874=>"111111111",
    9875=>"100110011",
    9876=>"001001011",
    9877=>"011001001",
    9878=>"110000010",
    9879=>"111011000",
    9880=>"000000000",
    9881=>"000000001",
    9882=>"100001001",
    9883=>"001000111",
    9884=>"110110110",
    9885=>"111011011",
    9886=>"111111111",
    9887=>"110001110",
    9888=>"010001110",
    9889=>"110000000",
    9890=>"101001100",
    9891=>"000001100",
    9892=>"010000010",
    9893=>"000100100",
    9894=>"110110111",
    9895=>"000000010",
    9896=>"110000000",
    9897=>"101111110",
    9898=>"111011001",
    9899=>"000000000",
    9900=>"111011011",
    9901=>"010000000",
    9902=>"001101101",
    9903=>"010110110",
    9904=>"000110010",
    9905=>"000000000",
    9906=>"001000010",
    9907=>"000000001",
    9908=>"101110110",
    9909=>"010011011",
    9910=>"110011011",
    9911=>"000100101",
    9912=>"010001010",
    9913=>"001000001",
    9914=>"111111100",
    9915=>"100100110",
    9916=>"111011001",
    9917=>"011001001",
    9918=>"011001000",
    9919=>"100110101",
    9920=>"000001001",
    9921=>"110110110",
    9922=>"110101001",
    9923=>"110110110",
    9924=>"100111111",
    9925=>"000000110",
    9926=>"010001001",
    9927=>"111100000",
    9928=>"000000010",
    9929=>"011000011",
    9930=>"110111011",
    9931=>"010100000",
    9932=>"101000010",
    9933=>"011001001",
    9934=>"001100001",
    9935=>"110100000",
    9936=>"010100110",
    9937=>"000000010",
    9938=>"000000000",
    9939=>"011100001",
    9940=>"111110110",
    9941=>"010100110",
    9942=>"000010000",
    9943=>"100001011",
    9944=>"000000000",
    9945=>"000000001",
    9946=>"100111111",
    9947=>"101100111",
    9948=>"111111111",
    9949=>"010110100",
    9950=>"100101001",
    9951=>"011000011",
    9952=>"000001001",
    9953=>"111011000",
    9954=>"100110110",
    9955=>"011001011",
    9956=>"001000000",
    9957=>"110110000",
    9958=>"010001000",
    9959=>"110110100",
    9960=>"100110110",
    9961=>"001001000",
    9962=>"000000000",
    9963=>"011100111",
    9964=>"000010100",
    9965=>"001001001",
    9966=>"110110100",
    9967=>"010111010",
    9968=>"000000001",
    9969=>"000000000",
    9970=>"110110010",
    9971=>"110110110",
    9972=>"011111111",
    9973=>"000001110",
    9974=>"110110101",
    9975=>"000001111",
    9976=>"000000000",
    9977=>"110110011",
    9978=>"110000000",
    9979=>"000111111",
    9980=>"100100101",
    9981=>"111001111",
    9982=>"101000000",
    9983=>"110101111",
    9984=>"011001000",
    9985=>"001100100",
    9986=>"100110110",
    9987=>"001000011",
    9988=>"001101000",
    9989=>"011011010",
    9990=>"111011000",
    9991=>"001100000",
    9992=>"000001111",
    9993=>"010111110",
    9994=>"010101110",
    9995=>"111100010",
    9996=>"111100010",
    9997=>"110011000",
    9998=>"010001101",
    9999=>"001101110",
    10000=>"011011010",
    10001=>"011001011",
    10002=>"000000000",
    10003=>"001001000",
    10004=>"100110011",
    10005=>"000100010",
    10006=>"010000010",
    10007=>"000011101",
    10008=>"111111001",
    10009=>"010111111",
    10010=>"111101000",
    10011=>"110010001",
    10012=>"111001001",
    10013=>"001001000",
    10014=>"000000000",
    10015=>"011011001",
    10016=>"100101101",
    10017=>"000001001",
    10018=>"101101010",
    10019=>"000001000",
    10020=>"001001100",
    10021=>"110100100",
    10022=>"011111111",
    10023=>"000111000",
    10024=>"001000011",
    10025=>"001001000",
    10026=>"011010010",
    10027=>"001001000",
    10028=>"011011100",
    10029=>"001100001",
    10030=>"011001000",
    10031=>"000111111",
    10032=>"000000011",
    10033=>"000100111",
    10034=>"110111100",
    10035=>"001001001",
    10036=>"111100100",
    10037=>"100000000",
    10038=>"011010010",
    10039=>"000000000",
    10040=>"100000000",
    10041=>"001001011",
    10042=>"001000011",
    10043=>"001001001",
    10044=>"100100110",
    10045=>"001001001",
    10046=>"111111101",
    10047=>"101111100",
    10048=>"101100101",
    10049=>"100100010",
    10050=>"011100110",
    10051=>"001001001",
    10052=>"111111010",
    10053=>"011111011",
    10054=>"010010000",
    10055=>"111100000",
    10056=>"000110010",
    10057=>"010010000",
    10058=>"011011111",
    10059=>"000100001",
    10060=>"010011011",
    10061=>"000000101",
    10062=>"010000000",
    10063=>"100110010",
    10064=>"000001011",
    10065=>"001100110",
    10066=>"001001000",
    10067=>"110110111",
    10068=>"100000000",
    10069=>"010110110",
    10070=>"111001001",
    10071=>"110010101",
    10072=>"111111101",
    10073=>"011111001",
    10074=>"100001111",
    10075=>"100110110",
    10076=>"111101001",
    10077=>"010111100",
    10078=>"100101101",
    10079=>"010011011",
    10080=>"011001001",
    10081=>"001011000",
    10082=>"011011111",
    10083=>"100110110",
    10084=>"001001000",
    10085=>"000000000",
    10086=>"001001100",
    10087=>"001001000",
    10088=>"000100110",
    10089=>"100100111",
    10090=>"111001000",
    10091=>"110101100",
    10092=>"100100100",
    10093=>"000100011",
    10094=>"111011000",
    10095=>"101101111",
    10096=>"000001110",
    10097=>"111111111",
    10098=>"001000000",
    10099=>"111110010",
    10100=>"100110110",
    10101=>"000000110",
    10102=>"000001100",
    10103=>"000111111",
    10104=>"011011000",
    10105=>"001011011",
    10106=>"001001011",
    10107=>"011011001",
    10108=>"101111100",
    10109=>"110111010",
    10110=>"100000100",
    10111=>"100100011",
    10112=>"011001100",
    10113=>"111000000",
    10114=>"110010000",
    10115=>"111011111",
    10116=>"111000100",
    10117=>"000111010",
    10118=>"111111000",
    10119=>"110111001",
    10120=>"000001001",
    10121=>"001111111",
    10122=>"000000110",
    10123=>"100000100",
    10124=>"000001111",
    10125=>"101100010",
    10126=>"110001001",
    10127=>"111011000",
    10128=>"001100010",
    10129=>"000100000",
    10130=>"111111000",
    10131=>"011000000",
    10132=>"111001001",
    10133=>"010100101",
    10134=>"101000000",
    10135=>"000000011",
    10136=>"111000000",
    10137=>"000001001",
    10138=>"111000000",
    10139=>"110001001",
    10140=>"000111111",
    10141=>"110010001",
    10142=>"011111000",
    10143=>"010110100",
    10144=>"000000111",
    10145=>"000110011",
    10146=>"101100110",
    10147=>"000000000",
    10148=>"010010000",
    10149=>"111000000",
    10150=>"001001111",
    10151=>"111010000",
    10152=>"101000000",
    10153=>"110000001",
    10154=>"011000011",
    10155=>"110100001",
    10156=>"001100110",
    10157=>"000010010",
    10158=>"100111010",
    10159=>"111111111",
    10160=>"000000010",
    10161=>"111100001",
    10162=>"000110111",
    10163=>"110011000",
    10164=>"001001110",
    10165=>"000111011",
    10166=>"000000010",
    10167=>"110010000",
    10168=>"110010000",
    10169=>"000000000",
    10170=>"100101101",
    10171=>"100111011",
    10172=>"010000100",
    10173=>"000100000",
    10174=>"011100100",
    10175=>"101101010",
    10176=>"011000111",
    10177=>"000011111",
    10178=>"000000111",
    10179=>"000000010",
    10180=>"111111000",
    10181=>"001001111",
    10182=>"110111100",
    10183=>"100111111",
    10184=>"000001011",
    10185=>"100001011",
    10186=>"000000000",
    10187=>"111010101",
    10188=>"111111011",
    10189=>"000111010",
    10190=>"110111111",
    10191=>"110111110",
    10192=>"000000111",
    10193=>"111001001",
    10194=>"000100000",
    10195=>"000110111",
    10196=>"111110111",
    10197=>"101101011",
    10198=>"000011111",
    10199=>"101111111",
    10200=>"111000100",
    10201=>"100111111",
    10202=>"101001011",
    10203=>"000100111",
    10204=>"011011000",
    10205=>"110100000",
    10206=>"110111001",
    10207=>"010110100",
    10208=>"100100000",
    10209=>"110110100",
    10210=>"111001111",
    10211=>"111000001",
    10212=>"001110010",
    10213=>"111010000",
    10214=>"111100100",
    10215=>"111011010",
    10216=>"001010010",
    10217=>"101011000",
    10218=>"111110000",
    10219=>"110111100",
    10220=>"111010000",
    10221=>"010010111",
    10222=>"001111000",
    10223=>"011111100",
    10224=>"010000100",
    10225=>"011100111",
    10226=>"101101000",
    10227=>"000111111",
    10228=>"101001101",
    10229=>"000000000",
    10230=>"111101111",
    10231=>"000011011",
    10232=>"001000000",
    10233=>"000000111",
    10234=>"001010110",
    10235=>"000000000",
    10236=>"111100100",
    10237=>"000000110",
    10238=>"110000010",
    10239=>"100001111",
    10240=>"010111111",
    10241=>"000110000",
    10242=>"111111010",
    10243=>"010110111",
    10244=>"111001111",
    10245=>"111001001",
    10246=>"111111111",
    10247=>"000000000",
    10248=>"101101111",
    10249=>"000000100",
    10250=>"001101001",
    10251=>"000000000",
    10252=>"000000010",
    10253=>"110111111",
    10254=>"110111111",
    10255=>"000000000",
    10256=>"000100000",
    10257=>"100011010",
    10258=>"111111111",
    10259=>"110100111",
    10260=>"110100110",
    10261=>"101100000",
    10262=>"000000101",
    10263=>"000000000",
    10264=>"011111111",
    10265=>"100000000",
    10266=>"101101101",
    10267=>"000000000",
    10268=>"011011111",
    10269=>"101101101",
    10270=>"111111111",
    10271=>"000000000",
    10272=>"111101101",
    10273=>"110101101",
    10274=>"011101110",
    10275=>"100101101",
    10276=>"111111111",
    10277=>"111101111",
    10278=>"100101100",
    10279=>"111111111",
    10280=>"001000100",
    10281=>"101101001",
    10282=>"101001011",
    10283=>"111101101",
    10284=>"001100100",
    10285=>"100100000",
    10286=>"101000001",
    10287=>"110110111",
    10288=>"010001000",
    10289=>"000010000",
    10290=>"000000100",
    10291=>"011011011",
    10292=>"101111111",
    10293=>"000000000",
    10294=>"100000000",
    10295=>"010011111",
    10296=>"000000000",
    10297=>"000001000",
    10298=>"000000001",
    10299=>"000100000",
    10300=>"101100000",
    10301=>"000111110",
    10302=>"000000000",
    10303=>"100101101",
    10304=>"100100100",
    10305=>"011001111",
    10306=>"000000000",
    10307=>"000000101",
    10308=>"010001001",
    10309=>"011010000",
    10310=>"110010010",
    10311=>"000000000",
    10312=>"000101001",
    10313=>"111101001",
    10314=>"000000000",
    10315=>"100100101",
    10316=>"000001000",
    10317=>"100000100",
    10318=>"000000000",
    10319=>"010010011",
    10320=>"000000000",
    10321=>"011110110",
    10322=>"000000101",
    10323=>"111011010",
    10324=>"111110011",
    10325=>"000010011",
    10326=>"000000111",
    10327=>"111110111",
    10328=>"111111111",
    10329=>"111011111",
    10330=>"001001011",
    10331=>"010010010",
    10332=>"111111111",
    10333=>"011011011",
    10334=>"001111101",
    10335=>"100100101",
    10336=>"111110111",
    10337=>"110110110",
    10338=>"111111010",
    10339=>"110110010",
    10340=>"010000000",
    10341=>"100110110",
    10342=>"110110011",
    10343=>"100000000",
    10344=>"010001001",
    10345=>"101101101",
    10346=>"111101111",
    10347=>"010000000",
    10348=>"111011001",
    10349=>"001000011",
    10350=>"101001101",
    10351=>"111101111",
    10352=>"111000000",
    10353=>"100000000",
    10354=>"111100100",
    10355=>"111111110",
    10356=>"100000000",
    10357=>"111111111",
    10358=>"101101001",
    10359=>"000000000",
    10360=>"001001000",
    10361=>"000000000",
    10362=>"101101100",
    10363=>"000000000",
    10364=>"100110111",
    10365=>"000000000",
    10366=>"010111111",
    10367=>"110111111",
    10368=>"101111111",
    10369=>"000110111",
    10370=>"001111000",
    10371=>"101000000",
    10372=>"011011000",
    10373=>"111010000",
    10374=>"011101110",
    10375=>"111011000",
    10376=>"101110000",
    10377=>"000111111",
    10378=>"001000110",
    10379=>"001111001",
    10380=>"110111000",
    10381=>"101111101",
    10382=>"001111010",
    10383=>"111010000",
    10384=>"011111000",
    10385=>"000111000",
    10386=>"010111000",
    10387=>"101111000",
    10388=>"011000000",
    10389=>"100100001",
    10390=>"111100000",
    10391=>"000001001",
    10392=>"000100110",
    10393=>"000110000",
    10394=>"111111110",
    10395=>"110100000",
    10396=>"000001000",
    10397=>"001111011",
    10398=>"101011001",
    10399=>"101111111",
    10400=>"111111000",
    10401=>"101111000",
    10402=>"001010000",
    10403=>"000000000",
    10404=>"101101000",
    10405=>"111010000",
    10406=>"111111000",
    10407=>"001111111",
    10408=>"010111010",
    10409=>"010010000",
    10410=>"011111111",
    10411=>"101110011",
    10412=>"111110000",
    10413=>"010110000",
    10414=>"010100000",
    10415=>"010010000",
    10416=>"011001111",
    10417=>"000000000",
    10418=>"000111111",
    10419=>"111101000",
    10420=>"100100000",
    10421=>"010011000",
    10422=>"000010010",
    10423=>"111101000",
    10424=>"100011010",
    10425=>"000000000",
    10426=>"001111111",
    10427=>"111000000",
    10428=>"000000101",
    10429=>"110101100",
    10430=>"100011000",
    10431=>"001111000",
    10432=>"111110000",
    10433=>"001110010",
    10434=>"001111111",
    10435=>"000101000",
    10436=>"011111000",
    10437=>"011001001",
    10438=>"100010000",
    10439=>"011111000",
    10440=>"110111000",
    10441=>"111011000",
    10442=>"000011000",
    10443=>"111111010",
    10444=>"011000000",
    10445=>"000010000",
    10446=>"111111000",
    10447=>"011010000",
    10448=>"111010000",
    10449=>"111111111",
    10450=>"101000000",
    10451=>"011011100",
    10452=>"111100100",
    10453=>"011011010",
    10454=>"111010101",
    10455=>"111000111",
    10456=>"000111000",
    10457=>"111100111",
    10458=>"101111000",
    10459=>"101000000",
    10460=>"100110110",
    10461=>"001010100",
    10462=>"111010000",
    10463=>"000001000",
    10464=>"111001000",
    10465=>"110101000",
    10466=>"101111100",
    10467=>"000010000",
    10468=>"101001000",
    10469=>"101111010",
    10470=>"011011111",
    10471=>"010111000",
    10472=>"110000011",
    10473=>"000000000",
    10474=>"110110101",
    10475=>"010100010",
    10476=>"111000000",
    10477=>"011000010",
    10478=>"001101000",
    10479=>"100011010",
    10480=>"011000000",
    10481=>"010111000",
    10482=>"000010011",
    10483=>"111010000",
    10484=>"000010111",
    10485=>"001101001",
    10486=>"111101000",
    10487=>"000111111",
    10488=>"011010010",
    10489=>"011011000",
    10490=>"011111010",
    10491=>"000010000",
    10492=>"111100000",
    10493=>"000010000",
    10494=>"110100000",
    10495=>"101111000",
    10496=>"111000000",
    10497=>"111101001",
    10498=>"111000101",
    10499=>"000000111",
    10500=>"011100100",
    10501=>"001010111",
    10502=>"111011111",
    10503=>"000111111",
    10504=>"011011000",
    10505=>"010010110",
    10506=>"111001001",
    10507=>"110011001",
    10508=>"111111111",
    10509=>"110111010",
    10510=>"011100111",
    10511=>"001100100",
    10512=>"000000000",
    10513=>"111100000",
    10514=>"000011011",
    10515=>"000001111",
    10516=>"010000000",
    10517=>"000010011",
    10518=>"010010000",
    10519=>"001111111",
    10520=>"000110110",
    10521=>"011100000",
    10522=>"000111111",
    10523=>"000001011",
    10524=>"000111111",
    10525=>"000011010",
    10526=>"011011001",
    10527=>"111001101",
    10528=>"010000000",
    10529=>"000001001",
    10530=>"011001001",
    10531=>"000000010",
    10532=>"001010111",
    10533=>"000000000",
    10534=>"111000111",
    10535=>"101000011",
    10536=>"110111010",
    10537=>"001001011",
    10538=>"101000000",
    10539=>"011110100",
    10540=>"100110101",
    10541=>"001000101",
    10542=>"011001001",
    10543=>"010011000",
    10544=>"010011001",
    10545=>"110101111",
    10546=>"011001110",
    10547=>"011010000",
    10548=>"010011000",
    10549=>"111111000",
    10550=>"101000000",
    10551=>"111000001",
    10552=>"101000101",
    10553=>"000000011",
    10554=>"000000101",
    10555=>"101100111",
    10556=>"000000110",
    10557=>"111010111",
    10558=>"000000101",
    10559=>"100111011",
    10560=>"111011000",
    10561=>"110000000",
    10562=>"000010100",
    10563=>"111111111",
    10564=>"100100000",
    10565=>"111000000",
    10566=>"000010000",
    10567=>"111111000",
    10568=>"000000101",
    10569=>"010001001",
    10570=>"111111000",
    10571=>"000110011",
    10572=>"100000000",
    10573=>"111000000",
    10574=>"001101100",
    10575=>"011000111",
    10576=>"111101000",
    10577=>"011000110",
    10578=>"000011111",
    10579=>"011010000",
    10580=>"110000000",
    10581=>"111001111",
    10582=>"011010010",
    10583=>"000110110",
    10584=>"110110100",
    10585=>"110110000",
    10586=>"000001001",
    10587=>"111000000",
    10588=>"000000011",
    10589=>"000000111",
    10590=>"011111111",
    10591=>"001000001",
    10592=>"111000001",
    10593=>"100000010",
    10594=>"101000000",
    10595=>"111001000",
    10596=>"111111000",
    10597=>"000110111",
    10598=>"100000011",
    10599=>"000000000",
    10600=>"011011000",
    10601=>"001110100",
    10602=>"010110100",
    10603=>"101111000",
    10604=>"111000000",
    10605=>"000000000",
    10606=>"101111111",
    10607=>"110000000",
    10608=>"001000110",
    10609=>"001000100",
    10610=>"010100111",
    10611=>"000110011",
    10612=>"111001101",
    10613=>"000000110",
    10614=>"110110110",
    10615=>"111110010",
    10616=>"000110110",
    10617=>"001110010",
    10618=>"100000100",
    10619=>"000000001",
    10620=>"000000110",
    10621=>"010010101",
    10622=>"000111111",
    10623=>"000110110",
    10624=>"101111011",
    10625=>"111011001",
    10626=>"111111001",
    10627=>"000101100",
    10628=>"101110111",
    10629=>"000101110",
    10630=>"000000101",
    10631=>"100010011",
    10632=>"000100110",
    10633=>"000000111",
    10634=>"111111111",
    10635=>"000100111",
    10636=>"111011001",
    10637=>"101000111",
    10638=>"100100010",
    10639=>"111011001",
    10640=>"000100110",
    10641=>"110111010",
    10642=>"000000110",
    10643=>"000001001",
    10644=>"000000101",
    10645=>"000011001",
    10646=>"010011001",
    10647=>"000000111",
    10648=>"001100101",
    10649=>"000001001",
    10650=>"000000000",
    10651=>"100000100",
    10652=>"000001110",
    10653=>"000100110",
    10654=>"110110111",
    10655=>"001110110",
    10656=>"100100100",
    10657=>"101101110",
    10658=>"101100111",
    10659=>"100100110",
    10660=>"000000100",
    10661=>"111111011",
    10662=>"010000000",
    10663=>"011110011",
    10664=>"001000110",
    10665=>"001000111",
    10666=>"111011101",
    10667=>"000100110",
    10668=>"000100110",
    10669=>"000100000",
    10670=>"100110111",
    10671=>"001110011",
    10672=>"000000110",
    10673=>"111111001",
    10674=>"100100001",
    10675=>"111000000",
    10676=>"000000100",
    10677=>"000100110",
    10678=>"000100110",
    10679=>"110111111",
    10680=>"011011011",
    10681=>"000000100",
    10682=>"100100100",
    10683=>"111011001",
    10684=>"111111011",
    10685=>"110011111",
    10686=>"000000100",
    10687=>"100100100",
    10688=>"100110111",
    10689=>"011011001",
    10690=>"000000110",
    10691=>"011011001",
    10692=>"010001100",
    10693=>"001000100",
    10694=>"000110100",
    10695=>"100100111",
    10696=>"000000001",
    10697=>"000100100",
    10698=>"000100110",
    10699=>"000010000",
    10700=>"101000010",
    10701=>"010111111",
    10702=>"100001111",
    10703=>"111011001",
    10704=>"110111101",
    10705=>"000010011",
    10706=>"000100110",
    10707=>"000000111",
    10708=>"000000001",
    10709=>"111111001",
    10710=>"100110110",
    10711=>"000000000",
    10712=>"100100111",
    10713=>"000000111",
    10714=>"000001000",
    10715=>"010011000",
    10716=>"000000000",
    10717=>"100110111",
    10718=>"100100110",
    10719=>"111111011",
    10720=>"001100100",
    10721=>"010010000",
    10722=>"011011000",
    10723=>"001111001",
    10724=>"000100110",
    10725=>"000001001",
    10726=>"000001001",
    10727=>"000100111",
    10728=>"011011101",
    10729=>"101110111",
    10730=>"000100100",
    10731=>"000100111",
    10732=>"010011000",
    10733=>"000000100",
    10734=>"000101100",
    10735=>"100000000",
    10736=>"111011011",
    10737=>"111101001",
    10738=>"000010111",
    10739=>"000100110",
    10740=>"111011001",
    10741=>"100111001",
    10742=>"011011100",
    10743=>"000000000",
    10744=>"000100111",
    10745=>"000011101",
    10746=>"010011000",
    10747=>"100110110",
    10748=>"111111011",
    10749=>"000000110",
    10750=>"011000100",
    10751=>"001000000",
    10752=>"101000000",
    10753=>"000110000",
    10754=>"101111111",
    10755=>"111101111",
    10756=>"111000000",
    10757=>"111111111",
    10758=>"010000000",
    10759=>"111000000",
    10760=>"000000100",
    10761=>"000000101",
    10762=>"101000111",
    10763=>"011011010",
    10764=>"010011111",
    10765=>"011111010",
    10766=>"101111111",
    10767=>"111000000",
    10768=>"111111110",
    10769=>"111111110",
    10770=>"001101001",
    10771=>"000011011",
    10772=>"100000000",
    10773=>"011000000",
    10774=>"000000001",
    10775=>"111111110",
    10776=>"100000000",
    10777=>"110111011",
    10778=>"110101101",
    10779=>"000000000",
    10780=>"111111111",
    10781=>"000101100",
    10782=>"001000000",
    10783=>"000000010",
    10784=>"000010100",
    10785=>"000000000",
    10786=>"001111110",
    10787=>"000010100",
    10788=>"010011111",
    10789=>"000010000",
    10790=>"000001011",
    10791=>"101101100",
    10792=>"011111111",
    10793=>"111110011",
    10794=>"000001100",
    10795=>"000000000",
    10796=>"001000111",
    10797=>"000000001",
    10798=>"110101101",
    10799=>"100000000",
    10800=>"111100100",
    10801=>"000010000",
    10802=>"010011110",
    10803=>"100000111",
    10804=>"100101001",
    10805=>"000001001",
    10806=>"111111000",
    10807=>"000000000",
    10808=>"000000000",
    10809=>"000000000",
    10810=>"010000000",
    10811=>"000000000",
    10812=>"011011011",
    10813=>"000010000",
    10814=>"000000000",
    10815=>"000000111",
    10816=>"111011111",
    10817=>"000111111",
    10818=>"000000000",
    10819=>"111111111",
    10820=>"000000110",
    10821=>"000000001",
    10822=>"001000000",
    10823=>"111100000",
    10824=>"111111111",
    10825=>"010111110",
    10826=>"111000011",
    10827=>"111111000",
    10828=>"011000011",
    10829=>"000000000",
    10830=>"111000100",
    10831=>"001001000",
    10832=>"000110000",
    10833=>"111101001",
    10834=>"100111111",
    10835=>"000000000",
    10836=>"101000100",
    10837=>"010011010",
    10838=>"000000000",
    10839=>"000000000",
    10840=>"100000100",
    10841=>"001000111",
    10842=>"010111111",
    10843=>"111101111",
    10844=>"101000101",
    10845=>"111001100",
    10846=>"000011111",
    10847=>"000011011",
    10848=>"010100100",
    10849=>"011000011",
    10850=>"100000010",
    10851=>"100111111",
    10852=>"111101101",
    10853=>"011101100",
    10854=>"111101100",
    10855=>"110111010",
    10856=>"100110111",
    10857=>"100000000",
    10858=>"000000000",
    10859=>"111000100",
    10860=>"101101101",
    10861=>"000000000",
    10862=>"101100011",
    10863=>"100100101",
    10864=>"000000000",
    10865=>"111111111",
    10866=>"000101101",
    10867=>"010111110",
    10868=>"000000001",
    10869=>"001000010",
    10870=>"010010000",
    10871=>"111110011",
    10872=>"000010011",
    10873=>"001010010",
    10874=>"111100100",
    10875=>"111111100",
    10876=>"101111111",
    10877=>"000000111",
    10878=>"000000000",
    10879=>"101111111",
    10880=>"111011011",
    10881=>"011000111",
    10882=>"100101111",
    10883=>"100110010",
    10884=>"000110111",
    10885=>"111111000",
    10886=>"100111000",
    10887=>"100001111",
    10888=>"110000100",
    10889=>"111101000",
    10890=>"011001001",
    10891=>"011011111",
    10892=>"011011011",
    10893=>"000110111",
    10894=>"000000000",
    10895=>"111011000",
    10896=>"000101111",
    10897=>"100001101",
    10898=>"000110010",
    10899=>"111111000",
    10900=>"100111000",
    10901=>"100000000",
    10902=>"011000101",
    10903=>"011111111",
    10904=>"001100100",
    10905=>"111000010",
    10906=>"000100100",
    10907=>"011000100",
    10908=>"100011101",
    10909=>"100111011",
    10910=>"000000101",
    10911=>"111110100",
    10912=>"011001011",
    10913=>"001100111",
    10914=>"000011001",
    10915=>"111011011",
    10916=>"111010000",
    10917=>"000100111",
    10918=>"000010111",
    10919=>"000100111",
    10920=>"100000101",
    10921=>"101000000",
    10922=>"111001000",
    10923=>"111000000",
    10924=>"000100111",
    10925=>"000110000",
    10926=>"111110111",
    10927=>"111100101",
    10928=>"000000111",
    10929=>"000000100",
    10930=>"000000101",
    10931=>"001100011",
    10932=>"011100100",
    10933=>"000101000",
    10934=>"110011000",
    10935=>"110111011",
    10936=>"011001000",
    10937=>"000100111",
    10938=>"000000101",
    10939=>"000001000",
    10940=>"001000100",
    10941=>"001001100",
    10942=>"000110100",
    10943=>"111111111",
    10944=>"011100000",
    10945=>"000000000",
    10946=>"111011111",
    10947=>"000001101",
    10948=>"111111101",
    10949=>"100100000",
    10950=>"000110100",
    10951=>"011000100",
    10952=>"111011000",
    10953=>"001100110",
    10954=>"000000111",
    10955=>"000000000",
    10956=>"100001000",
    10957=>"000011111",
    10958=>"111100111",
    10959=>"100110000",
    10960=>"001001111",
    10961=>"111001000",
    10962=>"000110111",
    10963=>"000010111",
    10964=>"000011011",
    10965=>"100001101",
    10966=>"000010110",
    10967=>"110100110",
    10968=>"000000101",
    10969=>"100011010",
    10970=>"011011001",
    10971=>"110111111",
    10972=>"111110000",
    10973=>"000000111",
    10974=>"000000000",
    10975=>"001001110",
    10976=>"000111101",
    10977=>"111000000",
    10978=>"100010011",
    10979=>"100110001",
    10980=>"000000101",
    10981=>"101011101",
    10982=>"000001111",
    10983=>"111000010",
    10984=>"011001011",
    10985=>"111000100",
    10986=>"111100000",
    10987=>"111111011",
    10988=>"100001001",
    10989=>"001000101",
    10990=>"000111011",
    10991=>"000101101",
    10992=>"000000000",
    10993=>"001001011",
    10994=>"000000000",
    10995=>"100100110",
    10996=>"101101111",
    10997=>"001001001",
    10998=>"110001011",
    10999=>"101111011",
    11000=>"000000111",
    11001=>"110000011",
    11002=>"001011011",
    11003=>"100011001",
    11004=>"000100100",
    11005=>"110000010",
    11006=>"100100000",
    11007=>"110111110",
    11008=>"110001111",
    11009=>"101001011",
    11010=>"110110001",
    11011=>"001110011",
    11012=>"011101100",
    11013=>"011011100",
    11014=>"000110011",
    11015=>"000000111",
    11016=>"011101011",
    11017=>"101110111",
    11018=>"111011001",
    11019=>"111111111",
    11020=>"001001001",
    11021=>"100111000",
    11022=>"000000100",
    11023=>"011100100",
    11024=>"011001000",
    11025=>"011001001",
    11026=>"000100010",
    11027=>"000111010",
    11028=>"011001001",
    11029=>"000111111",
    11030=>"000000001",
    11031=>"100100000",
    11032=>"011110101",
    11033=>"011101000",
    11034=>"011001001",
    11035=>"111011111",
    11036=>"100010000",
    11037=>"111111111",
    11038=>"101101000",
    11039=>"100000111",
    11040=>"011011001",
    11041=>"000000100",
    11042=>"101011011",
    11043=>"100001110",
    11044=>"100110011",
    11045=>"011001001",
    11046=>"011011000",
    11047=>"001011010",
    11048=>"000110100",
    11049=>"000100110",
    11050=>"001011000",
    11051=>"000000001",
    11052=>"110011011",
    11053=>"000100110",
    11054=>"000000011",
    11055=>"110110110",
    11056=>"100001010",
    11057=>"001000000",
    11058=>"011001111",
    11059=>"000000110",
    11060=>"001100001",
    11061=>"110011001",
    11062=>"110110000",
    11063=>"100110110",
    11064=>"010110001",
    11065=>"100100101",
    11066=>"110110111",
    11067=>"110000000",
    11068=>"001011000",
    11069=>"010101011",
    11070=>"001111100",
    11071=>"000001010",
    11072=>"011001001",
    11073=>"001010000",
    11074=>"000110111",
    11075=>"100000000",
    11076=>"001000010",
    11077=>"100110110",
    11078=>"000110010",
    11079=>"011011111",
    11080=>"001001011",
    11081=>"000110110",
    11082=>"110111001",
    11083=>"111000110",
    11084=>"100100110",
    11085=>"100110100",
    11086=>"110110111",
    11087=>"100110110",
    11088=>"011010000",
    11089=>"011001110",
    11090=>"000001001",
    11091=>"110010111",
    11092=>"000100110",
    11093=>"001001001",
    11094=>"101111010",
    11095=>"001100110",
    11096=>"111111111",
    11097=>"011111110",
    11098=>"101000110",
    11099=>"110110000",
    11100=>"111011111",
    11101=>"110110110",
    11102=>"101011000",
    11103=>"110110110",
    11104=>"010000000",
    11105=>"110110100",
    11106=>"100110110",
    11107=>"000100110",
    11108=>"000000000",
    11109=>"011001001",
    11110=>"000000101",
    11111=>"100110100",
    11112=>"001111001",
    11113=>"111001001",
    11114=>"010011011",
    11115=>"100001110",
    11116=>"110000000",
    11117=>"000001001",
    11118=>"100011001",
    11119=>"000000000",
    11120=>"100100001",
    11121=>"000111111",
    11122=>"011001100",
    11123=>"111001001",
    11124=>"100111000",
    11125=>"001001001",
    11126=>"111011011",
    11127=>"001111111",
    11128=>"000100110",
    11129=>"100001001",
    11130=>"011001011",
    11131=>"000101100",
    11132=>"010100100",
    11133=>"110011011",
    11134=>"111110111",
    11135=>"001101010",
    11136=>"000000000",
    11137=>"000111010",
    11138=>"000000110",
    11139=>"111011111",
    11140=>"000000000",
    11141=>"000000000",
    11142=>"000000000",
    11143=>"010000000",
    11144=>"000000001",
    11145=>"011011111",
    11146=>"011001001",
    11147=>"101000010",
    11148=>"000011000",
    11149=>"111111010",
    11150=>"000000000",
    11151=>"110001011",
    11152=>"001101101",
    11153=>"110111110",
    11154=>"000000000",
    11155=>"000000000",
    11156=>"000010000",
    11157=>"100000110",
    11158=>"001010101",
    11159=>"001111111",
    11160=>"000000000",
    11161=>"000000000",
    11162=>"000000000",
    11163=>"111111111",
    11164=>"111111101",
    11165=>"000000000",
    11166=>"100000000",
    11167=>"011111010",
    11168=>"000000000",
    11169=>"000000000",
    11170=>"000000000",
    11171=>"100111000",
    11172=>"111111111",
    11173=>"000000000",
    11174=>"110111111",
    11175=>"010111110",
    11176=>"111001001",
    11177=>"111001111",
    11178=>"000000000",
    11179=>"100000000",
    11180=>"111100100",
    11181=>"111111000",
    11182=>"010111111",
    11183=>"101000000",
    11184=>"001000000",
    11185=>"000111000",
    11186=>"000000100",
    11187=>"110100000",
    11188=>"000000000",
    11189=>"000000110",
    11190=>"010101100",
    11191=>"010111111",
    11192=>"000000111",
    11193=>"111101111",
    11194=>"110110111",
    11195=>"010111110",
    11196=>"111000000",
    11197=>"111110011",
    11198=>"111011111",
    11199=>"011111111",
    11200=>"111001101",
    11201=>"100011000",
    11202=>"000100011",
    11203=>"111111111",
    11204=>"000000000",
    11205=>"110111001",
    11206=>"000000000",
    11207=>"111111111",
    11208=>"100101111",
    11209=>"000000000",
    11210=>"101101111",
    11211=>"111111111",
    11212=>"111111111",
    11213=>"000100000",
    11214=>"111110111",
    11215=>"000111000",
    11216=>"000100110",
    11217=>"010011001",
    11218=>"100000011",
    11219=>"001011111",
    11220=>"111111111",
    11221=>"010111010",
    11222=>"000000000",
    11223=>"111111111",
    11224=>"000000100",
    11225=>"000000100",
    11226=>"111000000",
    11227=>"111111110",
    11228=>"000000001",
    11229=>"101001100",
    11230=>"000000000",
    11231=>"111111111",
    11232=>"000000000",
    11233=>"001001001",
    11234=>"111111111",
    11235=>"000100000",
    11236=>"011101111",
    11237=>"000010000",
    11238=>"001111100",
    11239=>"101001011",
    11240=>"000010011",
    11241=>"010010010",
    11242=>"000000001",
    11243=>"111111010",
    11244=>"111111111",
    11245=>"111101001",
    11246=>"000000000",
    11247=>"001000000",
    11248=>"111111101",
    11249=>"111111110",
    11250=>"111111111",
    11251=>"111000101",
    11252=>"110111111",
    11253=>"001000000",
    11254=>"111011111",
    11255=>"011110001",
    11256=>"100111001",
    11257=>"111111111",
    11258=>"000000000",
    11259=>"111000000",
    11260=>"001000001",
    11261=>"111110011",
    11262=>"110111111",
    11263=>"111111011",
    11264=>"010011011",
    11265=>"100000000",
    11266=>"100101100",
    11267=>"111000101",
    11268=>"001001101",
    11269=>"101011011",
    11270=>"000000000",
    11271=>"101100111",
    11272=>"100110100",
    11273=>"000010000",
    11274=>"100100101",
    11275=>"001001010",
    11276=>"111001001",
    11277=>"111011010",
    11278=>"111111101",
    11279=>"100000101",
    11280=>"110100100",
    11281=>"100100000",
    11282=>"001001001",
    11283=>"001011000",
    11284=>"101101100",
    11285=>"011000000",
    11286=>"000011000",
    11287=>"000011011",
    11288=>"110110100",
    11289=>"110110110",
    11290=>"110110000",
    11291=>"000011111",
    11292=>"101110000",
    11293=>"000001011",
    11294=>"001000001",
    11295=>"101101100",
    11296=>"000100000",
    11297=>"100100100",
    11298=>"001001000",
    11299=>"000000000",
    11300=>"011011010",
    11301=>"011100101",
    11302=>"100000100",
    11303=>"011011011",
    11304=>"010111101",
    11305=>"101001010",
    11306=>"111111100",
    11307=>"010110100",
    11308=>"111101001",
    11309=>"111100100",
    11310=>"000011000",
    11311=>"111111110",
    11312=>"011010000",
    11313=>"000111011",
    11314=>"100100000",
    11315=>"000000000",
    11316=>"000010000",
    11317=>"000000000",
    11318=>"111101101",
    11319=>"111001011",
    11320=>"101111011",
    11321=>"100000010",
    11322=>"110101100",
    11323=>"101000111",
    11324=>"100100000",
    11325=>"101101000",
    11326=>"101010011",
    11327=>"011111101",
    11328=>"101100000",
    11329=>"100101000",
    11330=>"100100000",
    11331=>"100011011",
    11332=>"111111111",
    11333=>"011011100",
    11334=>"011000010",
    11335=>"100100000",
    11336=>"011001000",
    11337=>"011011010",
    11338=>"100101000",
    11339=>"111111111",
    11340=>"100101010",
    11341=>"100000111",
    11342=>"101100111",
    11343=>"001011011",
    11344=>"000000000",
    11345=>"011010010",
    11346=>"000000011",
    11347=>"011001001",
    11348=>"110010001",
    11349=>"000000101",
    11350=>"011010001",
    11351=>"000000110",
    11352=>"100100100",
    11353=>"001001100",
    11354=>"111111001",
    11355=>"101101100",
    11356=>"001001001",
    11357=>"101001110",
    11358=>"000101000",
    11359=>"001000100",
    11360=>"001011000",
    11361=>"010010110",
    11362=>"111011111",
    11363=>"100100100",
    11364=>"100101000",
    11365=>"111101000",
    11366=>"110001000",
    11367=>"011011010",
    11368=>"101101110",
    11369=>"110100000",
    11370=>"000110101",
    11371=>"011000000",
    11372=>"110100000",
    11373=>"000000000",
    11374=>"010110010",
    11375=>"001001100",
    11376=>"100000101",
    11377=>"111111110",
    11378=>"000000000",
    11379=>"111101000",
    11380=>"001001111",
    11381=>"000000111",
    11382=>"011011000",
    11383=>"000101110",
    11384=>"100000110",
    11385=>"110110111",
    11386=>"110100001",
    11387=>"100100101",
    11388=>"110110100",
    11389=>"000111111",
    11390=>"000011000",
    11391=>"110011001",
    11392=>"000000000",
    11393=>"101001111",
    11394=>"011111110",
    11395=>"111011011",
    11396=>"011011000",
    11397=>"111101011",
    11398=>"110110111",
    11399=>"011001111",
    11400=>"110010000",
    11401=>"100111010",
    11402=>"011011111",
    11403=>"100000010",
    11404=>"001011111",
    11405=>"111100100",
    11406=>"100110101",
    11407=>"011011011",
    11408=>"100100110",
    11409=>"011011011",
    11410=>"111011001",
    11411=>"011001111",
    11412=>"011011111",
    11413=>"000100000",
    11414=>"000010010",
    11415=>"011111101",
    11416=>"000000000",
    11417=>"000001110",
    11418=>"100000000",
    11419=>"011111100",
    11420=>"010000000",
    11421=>"111100100",
    11422=>"111110100",
    11423=>"011000001",
    11424=>"000100110",
    11425=>"111111111",
    11426=>"011011011",
    11427=>"000100101",
    11428=>"111011110",
    11429=>"001011111",
    11430=>"101101001",
    11431=>"111100010",
    11432=>"000000110",
    11433=>"011111111",
    11434=>"011010101",
    11435=>"101000001",
    11436=>"100000111",
    11437=>"111011011",
    11438=>"100100000",
    11439=>"111011011",
    11440=>"010010011",
    11441=>"000100111",
    11442=>"000000010",
    11443=>"010000000",
    11444=>"110100100",
    11445=>"100100000",
    11446=>"110100100",
    11447=>"000010000",
    11448=>"011011111",
    11449=>"010100100",
    11450=>"100110000",
    11451=>"001011111",
    11452=>"000001010",
    11453=>"000100000",
    11454=>"110111111",
    11455=>"011001000",
    11456=>"000000010",
    11457=>"000100100",
    11458=>"100110000",
    11459=>"001001001",
    11460=>"110000010",
    11461=>"011000101",
    11462=>"100000100",
    11463=>"100100000",
    11464=>"110100100",
    11465=>"100100100",
    11466=>"000011111",
    11467=>"010011100",
    11468=>"010010110",
    11469=>"011011111",
    11470=>"110100010",
    11471=>"110100000",
    11472=>"011011011",
    11473=>"010000100",
    11474=>"110110100",
    11475=>"110110000",
    11476=>"111110100",
    11477=>"001011011",
    11478=>"110100110",
    11479=>"100000000",
    11480=>"001001011",
    11481=>"100110001",
    11482=>"001010001",
    11483=>"011011011",
    11484=>"111111100",
    11485=>"000000010",
    11486=>"110110000",
    11487=>"100100100",
    11488=>"011111101",
    11489=>"011001011",
    11490=>"001001011",
    11491=>"011011011",
    11492=>"100100000",
    11493=>"000000100",
    11494=>"001110010",
    11495=>"110100000",
    11496=>"110100000",
    11497=>"000000110",
    11498=>"000101110",
    11499=>"101100000",
    11500=>"111001001",
    11501=>"001100100",
    11502=>"000010100",
    11503=>"100000000",
    11504=>"010011110",
    11505=>"100100000",
    11506=>"100100100",
    11507=>"100100000",
    11508=>"001001011",
    11509=>"001100000",
    11510=>"100100000",
    11511=>"010110111",
    11512=>"110100110",
    11513=>"101100100",
    11514=>"011001111",
    11515=>"110100100",
    11516=>"111000111",
    11517=>"111110001",
    11518=>"001001011",
    11519=>"110110000",
    11520=>"110110100",
    11521=>"100100100",
    11522=>"110110011",
    11523=>"001000000",
    11524=>"100100000",
    11525=>"110110111",
    11526=>"111100111",
    11527=>"011001001",
    11528=>"100001000",
    11529=>"010111111",
    11530=>"110011111",
    11531=>"000011011",
    11532=>"000000000",
    11533=>"100100100",
    11534=>"101000101",
    11535=>"001001001",
    11536=>"000000110",
    11537=>"010010000",
    11538=>"001100101",
    11539=>"110101111",
    11540=>"011011001",
    11541=>"110010000",
    11542=>"010000011",
    11543=>"011001011",
    11544=>"001000100",
    11545=>"110010000",
    11546=>"000000000",
    11547=>"000000000",
    11548=>"111111110",
    11549=>"101100100",
    11550=>"010010111",
    11551=>"011111000",
    11552=>"101101001",
    11553=>"101000100",
    11554=>"000000100",
    11555=>"000101011",
    11556=>"011011011",
    11557=>"011011111",
    11558=>"101101111",
    11559=>"100100100",
    11560=>"001011001",
    11561=>"011111111",
    11562=>"000000000",
    11563=>"100100000",
    11564=>"000011011",
    11565=>"001111001",
    11566=>"100110110",
    11567=>"001001101",
    11568=>"000000011",
    11569=>"001010011",
    11570=>"001011011",
    11571=>"011000000",
    11572=>"100000000",
    11573=>"000001100",
    11574=>"011001001",
    11575=>"111100111",
    11576=>"000010000",
    11577=>"111000100",
    11578=>"000000000",
    11579=>"011010000",
    11580=>"101000000",
    11581=>"011010101",
    11582=>"111111110",
    11583=>"001011001",
    11584=>"010111100",
    11585=>"011001011",
    11586=>"011011111",
    11587=>"000110110",
    11588=>"111111110",
    11589=>"101110100",
    11590=>"100110000",
    11591=>"011011011",
    11592=>"111010001",
    11593=>"100100100",
    11594=>"101111011",
    11595=>"011011001",
    11596=>"011011110",
    11597=>"000011111",
    11598=>"111111011",
    11599=>"100110100",
    11600=>"110110000",
    11601=>"111011001",
    11602=>"110110110",
    11603=>"110011111",
    11604=>"111010111",
    11605=>"001111011",
    11606=>"001000000",
    11607=>"110110011",
    11608=>"000000110",
    11609=>"110111111",
    11610=>"100000011",
    11611=>"111111011",
    11612=>"100100100",
    11613=>"000001100",
    11614=>"111111111",
    11615=>"100111101",
    11616=>"111111111",
    11617=>"111001001",
    11618=>"111111000",
    11619=>"011001000",
    11620=>"011001010",
    11621=>"011101101",
    11622=>"101100100",
    11623=>"111111011",
    11624=>"000000000",
    11625=>"010000000",
    11626=>"110100100",
    11627=>"011011111",
    11628=>"111000001",
    11629=>"001001101",
    11630=>"110110111",
    11631=>"111001000",
    11632=>"011011011",
    11633=>"100111100",
    11634=>"100110110",
    11635=>"011111101",
    11636=>"000000000",
    11637=>"000010111",
    11638=>"000011011",
    11639=>"011001000",
    11640=>"000011011",
    11641=>"011011011",
    11642=>"010000001",
    11643=>"001001001",
    11644=>"100001100",
    11645=>"100000010",
    11646=>"111011011",
    11647=>"111001001",
    11648=>"110010000",
    11649=>"011001011",
    11650=>"011001011",
    11651=>"110011001",
    11652=>"101111000",
    11653=>"000110110",
    11654=>"111000100",
    11655=>"111000100",
    11656=>"000011001",
    11657=>"111000010",
    11658=>"011111011",
    11659=>"011111101",
    11660=>"001011000",
    11661=>"100111110",
    11662=>"100111111",
    11663=>"100000100",
    11664=>"001000100",
    11665=>"000011110",
    11666=>"000000000",
    11667=>"011100001",
    11668=>"000111000",
    11669=>"100100110",
    11670=>"100100110",
    11671=>"000010110",
    11672=>"010001001",
    11673=>"100011010",
    11674=>"001001001",
    11675=>"111100110",
    11676=>"100000101",
    11677=>"000101101",
    11678=>"011101110",
    11679=>"001011001",
    11680=>"110111011",
    11681=>"110001001",
    11682=>"011011001",
    11683=>"111001101",
    11684=>"011001110",
    11685=>"000011000",
    11686=>"001001110",
    11687=>"011011011",
    11688=>"010001001",
    11689=>"000001000",
    11690=>"101010011",
    11691=>"110010001",
    11692=>"111101100",
    11693=>"000001001",
    11694=>"110110110",
    11695=>"111011000",
    11696=>"111111000",
    11697=>"011111010",
    11698=>"011011001",
    11699=>"111000000",
    11700=>"000100100",
    11701=>"000110110",
    11702=>"100100100",
    11703=>"000100110",
    11704=>"011011111",
    11705=>"111001110",
    11706=>"110001001",
    11707=>"010000001",
    11708=>"000001011",
    11709=>"000000000",
    11710=>"101001001",
    11711=>"111101011",
    11712=>"111001001",
    11713=>"011011001",
    11714=>"000100110",
    11715=>"000000001",
    11716=>"000001001",
    11717=>"111011001",
    11718=>"100111110",
    11719=>"010000001",
    11720=>"100101011",
    11721=>"000100100",
    11722=>"111011110",
    11723=>"010001001",
    11724=>"111011001",
    11725=>"111111100",
    11726=>"101011100",
    11727=>"000111110",
    11728=>"101100110",
    11729=>"001001101",
    11730=>"100100110",
    11731=>"100110110",
    11732=>"110000100",
    11733=>"100110110",
    11734=>"111001111",
    11735=>"110000110",
    11736=>"111111011",
    11737=>"111110000",
    11738=>"000001000",
    11739=>"000100110",
    11740=>"101001001",
    11741=>"111011000",
    11742=>"001011001",
    11743=>"000001101",
    11744=>"000111010",
    11745=>"110110010",
    11746=>"111011011",
    11747=>"001000001",
    11748=>"111001001",
    11749=>"011001000",
    11750=>"001001001",
    11751=>"011100001",
    11752=>"011010001",
    11753=>"111011011",
    11754=>"000000000",
    11755=>"110111110",
    11756=>"100111111",
    11757=>"100100010",
    11758=>"100100100",
    11759=>"000000000",
    11760=>"011001000",
    11761=>"111000011",
    11762=>"001001011",
    11763=>"100110100",
    11764=>"000110110",
    11765=>"110011011",
    11766=>"000000000",
    11767=>"001000001",
    11768=>"011001111",
    11769=>"001011000",
    11770=>"001101110",
    11771=>"100100110",
    11772=>"000010110",
    11773=>"001110110",
    11774=>"000000001",
    11775=>"100001000",
    11776=>"100000000",
    11777=>"011000000",
    11778=>"010111111",
    11779=>"000000000",
    11780=>"010011001",
    11781=>"010000101",
    11782=>"110100100",
    11783=>"101111111",
    11784=>"111011111",
    11785=>"101001111",
    11786=>"111111100",
    11787=>"111111000",
    11788=>"000111011",
    11789=>"010010000",
    11790=>"000001010",
    11791=>"110100000",
    11792=>"010110110",
    11793=>"101000101",
    11794=>"000110010",
    11795=>"111100100",
    11796=>"001000000",
    11797=>"000000000",
    11798=>"010101100",
    11799=>"111111010",
    11800=>"011011111",
    11801=>"011111001",
    11802=>"011011100",
    11803=>"111111111",
    11804=>"000000000",
    11805=>"100000000",
    11806=>"100100000",
    11807=>"000000000",
    11808=>"010111101",
    11809=>"101100111",
    11810=>"110111111",
    11811=>"111101000",
    11812=>"111111111",
    11813=>"111011101",
    11814=>"001000111",
    11815=>"001000111",
    11816=>"111111011",
    11817=>"010000000",
    11818=>"011011111",
    11819=>"000110110",
    11820=>"111011111",
    11821=>"010100101",
    11822=>"001000101",
    11823=>"001000000",
    11824=>"100111111",
    11825=>"001000010",
    11826=>"011111010",
    11827=>"001001101",
    11828=>"010100101",
    11829=>"000100000",
    11830=>"000000000",
    11831=>"001111111",
    11832=>"111111011",
    11833=>"101000101",
    11834=>"110000111",
    11835=>"111000110",
    11836=>"100000001",
    11837=>"101000000",
    11838=>"111111110",
    11839=>"010111000",
    11840=>"011011110",
    11841=>"111101000",
    11842=>"110000000",
    11843=>"000000000",
    11844=>"000100111",
    11845=>"110010000",
    11846=>"000110010",
    11847=>"111111100",
    11848=>"010011111",
    11849=>"000000000",
    11850=>"010111011",
    11851=>"000111011",
    11852=>"101010111",
    11853=>"101100111",
    11854=>"111111111",
    11855=>"001000111",
    11856=>"111110001",
    11857=>"000000001",
    11858=>"000000001",
    11859=>"111111111",
    11860=>"010010010",
    11861=>"000000011",
    11862=>"010111000",
    11863=>"000000101",
    11864=>"001001000",
    11865=>"110110010",
    11866=>"110010011",
    11867=>"111111111",
    11868=>"011011011",
    11869=>"000011000",
    11870=>"011001010",
    11871=>"101101100",
    11872=>"110111110",
    11873=>"100110111",
    11874=>"000000000",
    11875=>"111111110",
    11876=>"100111111",
    11877=>"001000111",
    11878=>"001010100",
    11879=>"010111000",
    11880=>"010110010",
    11881=>"111111000",
    11882=>"001111110",
    11883=>"111111101",
    11884=>"101001000",
    11885=>"001001111",
    11886=>"101010010",
    11887=>"000001000",
    11888=>"000000000",
    11889=>"000000000",
    11890=>"111001001",
    11891=>"011111000",
    11892=>"101000111",
    11893=>"101101111",
    11894=>"111101111",
    11895=>"111111111",
    11896=>"001111010",
    11897=>"111111000",
    11898=>"110000100",
    11899=>"111111100",
    11900=>"001001001",
    11901=>"000001010",
    11902=>"111001111",
    11903=>"111100111",
    11904=>"100100100",
    11905=>"011010000",
    11906=>"001011011",
    11907=>"111111111",
    11908=>"000100110",
    11909=>"110101100",
    11910=>"000000000",
    11911=>"011010010",
    11912=>"100100100",
    11913=>"000000000",
    11914=>"111111111",
    11915=>"000111111",
    11916=>"010000001",
    11917=>"111011001",
    11918=>"010000110",
    11919=>"011011011",
    11920=>"000000000",
    11921=>"011110000",
    11922=>"110100001",
    11923=>"110111111",
    11924=>"100100101",
    11925=>"000001110",
    11926=>"000000000",
    11927=>"001001000",
    11928=>"111100000",
    11929=>"001011011",
    11930=>"100000000",
    11931=>"110100110",
    11932=>"010011011",
    11933=>"110100100",
    11934=>"010110010",
    11935=>"111111111",
    11936=>"111110000",
    11937=>"111110110",
    11938=>"100110111",
    11939=>"100100100",
    11940=>"100100100",
    11941=>"110000101",
    11942=>"011000000",
    11943=>"101100100",
    11944=>"001111011",
    11945=>"110111100",
    11946=>"110100100",
    11947=>"110100000",
    11948=>"100001001",
    11949=>"010111101",
    11950=>"100100100",
    11951=>"011011011",
    11952=>"100000100",
    11953=>"001011011",
    11954=>"000000001",
    11955=>"100101100",
    11956=>"100100100",
    11957=>"000100110",
    11958=>"000000011",
    11959=>"111110110",
    11960=>"001111111",
    11961=>"111011101",
    11962=>"100100100",
    11963=>"001011001",
    11964=>"011011000",
    11965=>"101111100",
    11966=>"000000000",
    11967=>"110100000",
    11968=>"110010000",
    11969=>"001000000",
    11970=>"100101101",
    11971=>"000011011",
    11972=>"100100110",
    11973=>"100000000",
    11974=>"101001111",
    11975=>"001101100",
    11976=>"000110110",
    11977=>"100000000",
    11978=>"110111011",
    11979=>"010000000",
    11980=>"100010011",
    11981=>"111101100",
    11982=>"100110110",
    11983=>"001011011",
    11984=>"101000001",
    11985=>"100000000",
    11986=>"011000000",
    11987=>"001001111",
    11988=>"100100100",
    11989=>"001011001",
    11990=>"000000100",
    11991=>"000101100",
    11992=>"110110011",
    11993=>"000100000",
    11994=>"111111110",
    11995=>"011000000",
    11996=>"110110110",
    11997=>"101101111",
    11998=>"111110110",
    11999=>"101001011",
    12000=>"100100000",
    12001=>"000001000",
    12002=>"001011011",
    12003=>"110110011",
    12004=>"100100100",
    12005=>"100100100",
    12006=>"000100100",
    12007=>"000010110",
    12008=>"101110110",
    12009=>"001010010",
    12010=>"110110010",
    12011=>"001001000",
    12012=>"011011011",
    12013=>"011100110",
    12014=>"100100101",
    12015=>"010100111",
    12016=>"011011011",
    12017=>"000001101",
    12018=>"001011011",
    12019=>"000111111",
    12020=>"011011000",
    12021=>"000011011",
    12022=>"100000000",
    12023=>"111101111",
    12024=>"100010000",
    12025=>"000011001",
    12026=>"011011001",
    12027=>"001011011",
    12028=>"011101001",
    12029=>"101011111",
    12030=>"100111011",
    12031=>"110100100",
    12032=>"000010010",
    12033=>"111100000",
    12034=>"111010000",
    12035=>"011111111",
    12036=>"001101100",
    12037=>"111111111",
    12038=>"000010101",
    12039=>"000000000",
    12040=>"001101001",
    12041=>"100101100",
    12042=>"010000000",
    12043=>"011101101",
    12044=>"001001110",
    12045=>"010111110",
    12046=>"110100000",
    12047=>"100100100",
    12048=>"000111110",
    12049=>"000000111",
    12050=>"001001000",
    12051=>"100000000",
    12052=>"010010001",
    12053=>"000000000",
    12054=>"000000000",
    12055=>"000000111",
    12056=>"000000001",
    12057=>"100001101",
    12058=>"000000000",
    12059=>"111111111",
    12060=>"000110011",
    12061=>"011111011",
    12062=>"001000000",
    12063=>"001111100",
    12064=>"000011101",
    12065=>"011100100",
    12066=>"101101110",
    12067=>"000001100",
    12068=>"110111111",
    12069=>"011111111",
    12070=>"010111111",
    12071=>"000000000",
    12072=>"111101010",
    12073=>"000001001",
    12074=>"110110101",
    12075=>"001100000",
    12076=>"011011011",
    12077=>"111111111",
    12078=>"000000101",
    12079=>"010111111",
    12080=>"111111111",
    12081=>"111000000",
    12082=>"000111111",
    12083=>"100000000",
    12084=>"110111101",
    12085=>"000000001",
    12086=>"111111111",
    12087=>"000000000",
    12088=>"111100100",
    12089=>"000000000",
    12090=>"001001101",
    12091=>"000000000",
    12092=>"101000000",
    12093=>"000000000",
    12094=>"110011110",
    12095=>"011111011",
    12096=>"010100110",
    12097=>"001001100",
    12098=>"010010110",
    12099=>"000001110",
    12100=>"111111111",
    12101=>"110110110",
    12102=>"100000000",
    12103=>"111111010",
    12104=>"000100101",
    12105=>"110111101",
    12106=>"000000111",
    12107=>"000000000",
    12108=>"000110110",
    12109=>"000000000",
    12110=>"100000001",
    12111=>"000100100",
    12112=>"000101000",
    12113=>"000000000",
    12114=>"000000100",
    12115=>"111111101",
    12116=>"010011011",
    12117=>"000000000",
    12118=>"001111011",
    12119=>"111101000",
    12120=>"001000100",
    12121=>"010111111",
    12122=>"000000000",
    12123=>"000010000",
    12124=>"000001011",
    12125=>"011000001",
    12126=>"011100000",
    12127=>"101011111",
    12128=>"100111010",
    12129=>"000000001",
    12130=>"010111111",
    12131=>"010111010",
    12132=>"000001000",
    12133=>"001000001",
    12134=>"000000000",
    12135=>"111000010",
    12136=>"000000000",
    12137=>"000000000",
    12138=>"100101101",
    12139=>"010001111",
    12140=>"010000001",
    12141=>"000000000",
    12142=>"111111000",
    12143=>"100000001",
    12144=>"000000000",
    12145=>"010000000",
    12146=>"000000000",
    12147=>"001001101",
    12148=>"000000000",
    12149=>"000000000",
    12150=>"110111110",
    12151=>"011011111",
    12152=>"011011110",
    12153=>"111000111",
    12154=>"001000000",
    12155=>"011101111",
    12156=>"000000000",
    12157=>"111111010",
    12158=>"110000010",
    12159=>"111111111",
    12160=>"101000100",
    12161=>"100000001",
    12162=>"100000001",
    12163=>"011111111",
    12164=>"000000000",
    12165=>"001000000",
    12166=>"000000011",
    12167=>"100000000",
    12168=>"011111110",
    12169=>"000000000",
    12170=>"110100000",
    12171=>"000000001",
    12172=>"001011110",
    12173=>"011111000",
    12174=>"111111111",
    12175=>"111111111",
    12176=>"011111110",
    12177=>"101100001",
    12178=>"010000001",
    12179=>"111111111",
    12180=>"011110000",
    12181=>"010110100",
    12182=>"010000000",
    12183=>"111111110",
    12184=>"111111111",
    12185=>"111111111",
    12186=>"100100000",
    12187=>"000000000",
    12188=>"000000000",
    12189=>"010111111",
    12190=>"000000000",
    12191=>"000000000",
    12192=>"010111101",
    12193=>"111110111",
    12194=>"000000000",
    12195=>"011101111",
    12196=>"000010100",
    12197=>"011110100",
    12198=>"110000000",
    12199=>"011111011",
    12200=>"011100001",
    12201=>"111111111",
    12202=>"011110100",
    12203=>"111011111",
    12204=>"000000000",
    12205=>"001010100",
    12206=>"011100000",
    12207=>"010111000",
    12208=>"011110100",
    12209=>"000101010",
    12210=>"000000001",
    12211=>"011111111",
    12212=>"000010010",
    12213=>"010000100",
    12214=>"000000101",
    12215=>"010110101",
    12216=>"000100000",
    12217=>"110100000",
    12218=>"011111111",
    12219=>"100001000",
    12220=>"100000001",
    12221=>"000000000",
    12222=>"111111110",
    12223=>"001111110",
    12224=>"000000011",
    12225=>"101001001",
    12226=>"001111110",
    12227=>"100001000",
    12228=>"111111111",
    12229=>"111111110",
    12230=>"001110100",
    12231=>"111000000",
    12232=>"100000001",
    12233=>"000000111",
    12234=>"000000000",
    12235=>"110100111",
    12236=>"001111110",
    12237=>"000100000",
    12238=>"000101100",
    12239=>"000001010",
    12240=>"001111010",
    12241=>"001110100",
    12242=>"100000111",
    12243=>"000101000",
    12244=>"011111110",
    12245=>"011111100",
    12246=>"000000000",
    12247=>"110100100",
    12248=>"000000000",
    12249=>"100110100",
    12250=>"100001010",
    12251=>"001111000",
    12252=>"111111011",
    12253=>"000000001",
    12254=>"000000000",
    12255=>"111111001",
    12256=>"011010010",
    12257=>"000000001",
    12258=>"001111010",
    12259=>"010111000",
    12260=>"000000010",
    12261=>"010000001",
    12262=>"100000011",
    12263=>"111001000",
    12264=>"001011010",
    12265=>"110100001",
    12266=>"111111111",
    12267=>"011111000",
    12268=>"010010011",
    12269=>"000000000",
    12270=>"110000100",
    12271=>"000000000",
    12272=>"110110101",
    12273=>"000000000",
    12274=>"100000001",
    12275=>"011110101",
    12276=>"010111001",
    12277=>"000001011",
    12278=>"101001111",
    12279=>"111111010",
    12280=>"000000000",
    12281=>"101100000",
    12282=>"110110111",
    12283=>"111111011",
    12284=>"000000000",
    12285=>"111111111",
    12286=>"001100101",
    12287=>"111101111",
    12288=>"111111111",
    12289=>"000000000",
    12290=>"111111111",
    12291=>"001011001",
    12292=>"000000000",
    12293=>"000000000",
    12294=>"111111111",
    12295=>"111000000",
    12296=>"111111111",
    12297=>"001001111",
    12298=>"000000000",
    12299=>"001000000",
    12300=>"000000000",
    12301=>"010111110",
    12302=>"000000100",
    12303=>"100001001",
    12304=>"111100110",
    12305=>"010010111",
    12306=>"011001011",
    12307=>"110100100",
    12308=>"000000000",
    12309=>"000000010",
    12310=>"111011110",
    12311=>"000000000",
    12312=>"011010111",
    12313=>"100000001",
    12314=>"000000000",
    12315=>"110100100",
    12316=>"000000000",
    12317=>"100010000",
    12318=>"000110111",
    12319=>"010011001",
    12320=>"110111101",
    12321=>"000000000",
    12322=>"000100000",
    12323=>"000000001",
    12324=>"001001001",
    12325=>"010010000",
    12326=>"111111100",
    12327=>"111111011",
    12328=>"011001000",
    12329=>"001001111",
    12330=>"100000000",
    12331=>"000010110",
    12332=>"001001001",
    12333=>"010111111",
    12334=>"000001000",
    12335=>"010111111",
    12336=>"110111111",
    12337=>"011011000",
    12338=>"001000000",
    12339=>"000101111",
    12340=>"000000001",
    12341=>"001000111",
    12342=>"101101101",
    12343=>"000000000",
    12344=>"001011100",
    12345=>"011111101",
    12346=>"100100110",
    12347=>"000000000",
    12348=>"000000000",
    12349=>"000000010",
    12350=>"011001001",
    12351=>"001000001",
    12352=>"000000000",
    12353=>"000001111",
    12354=>"000000000",
    12355=>"000000000",
    12356=>"111111111",
    12357=>"111111011",
    12358=>"111111111",
    12359=>"000000000",
    12360=>"101000001",
    12361=>"111111000",
    12362=>"010111011",
    12363=>"111110000",
    12364=>"111110000",
    12365=>"111111111",
    12366=>"101111111",
    12367=>"111111000",
    12368=>"111110111",
    12369=>"111001111",
    12370=>"000100100",
    12371=>"000000000",
    12372=>"111110100",
    12373=>"100000000",
    12374=>"111111000",
    12375=>"001000000",
    12376=>"100100100",
    12377=>"000101111",
    12378=>"100000001",
    12379=>"000111000",
    12380=>"010110110",
    12381=>"001000000",
    12382=>"000010000",
    12383=>"000000000",
    12384=>"111111110",
    12385=>"111111111",
    12386=>"111111111",
    12387=>"000110000",
    12388=>"000011111",
    12389=>"000111001",
    12390=>"111100100",
    12391=>"110101000",
    12392=>"000000000",
    12393=>"110000000",
    12394=>"010000110",
    12395=>"000111110",
    12396=>"101101111",
    12397=>"111111111",
    12398=>"000000000",
    12399=>"010000001",
    12400=>"000101111",
    12401=>"100011001",
    12402=>"111111100",
    12403=>"110110000",
    12404=>"111111111",
    12405=>"101000101",
    12406=>"111001101",
    12407=>"110000000",
    12408=>"111111111",
    12409=>"001000000",
    12410=>"000000000",
    12411=>"111110111",
    12412=>"000000000",
    12413=>"110111010",
    12414=>"000000000",
    12415=>"000010000",
    12416=>"101111010",
    12417=>"110011010",
    12418=>"111010011",
    12419=>"111100111",
    12420=>"011111111",
    12421=>"010011110",
    12422=>"000000100",
    12423=>"000000111",
    12424=>"011011000",
    12425=>"011011001",
    12426=>"001101100",
    12427=>"111101101",
    12428=>"101000010",
    12429=>"111111000",
    12430=>"110110110",
    12431=>"001000111",
    12432=>"000000000",
    12433=>"101101100",
    12434=>"000000011",
    12435=>"100100101",
    12436=>"101000000",
    12437=>"000011111",
    12438=>"111111101",
    12439=>"100101111",
    12440=>"001001111",
    12441=>"110111111",
    12442=>"100000100",
    12443=>"101011111",
    12444=>"000000010",
    12445=>"011010101",
    12446=>"110110101",
    12447=>"111101111",
    12448=>"111001011",
    12449=>"011000111",
    12450=>"011101001",
    12451=>"100100000",
    12452=>"111000000",
    12453=>"000000101",
    12454=>"101000111",
    12455=>"011011000",
    12456=>"101101110",
    12457=>"101101001",
    12458=>"100000000",
    12459=>"111111000",
    12460=>"111001001",
    12461=>"111111111",
    12462=>"000001000",
    12463=>"101101111",
    12464=>"100111111",
    12465=>"011011011",
    12466=>"111100110",
    12467=>"000010101",
    12468=>"110111111",
    12469=>"001000100",
    12470=>"000010000",
    12471=>"111111111",
    12472=>"100100000",
    12473=>"111101111",
    12474=>"111110100",
    12475=>"000000100",
    12476=>"101101101",
    12477=>"000100000",
    12478=>"011010010",
    12479=>"100101000",
    12480=>"000010000",
    12481=>"101101101",
    12482=>"001000111",
    12483=>"000000100",
    12484=>"000000001",
    12485=>"000000000",
    12486=>"010010010",
    12487=>"000001101",
    12488=>"001000000",
    12489=>"111111010",
    12490=>"100111000",
    12491=>"000000110",
    12492=>"111101000",
    12493=>"011011000",
    12494=>"011111111",
    12495=>"000011011",
    12496=>"100100111",
    12497=>"111110010",
    12498=>"100101111",
    12499=>"010000000",
    12500=>"000010000",
    12501=>"001001000",
    12502=>"110001111",
    12503=>"000000000",
    12504=>"100110000",
    12505=>"110111110",
    12506=>"000000000",
    12507=>"111101000",
    12508=>"101111001",
    12509=>"111110110",
    12510=>"011001000",
    12511=>"001111111",
    12512=>"110110000",
    12513=>"010111110",
    12514=>"111111000",
    12515=>"000111111",
    12516=>"111111111",
    12517=>"010110000",
    12518=>"110111000",
    12519=>"100110100",
    12520=>"011011000",
    12521=>"101101100",
    12522=>"001001000",
    12523=>"001000000",
    12524=>"110111000",
    12525=>"111111100",
    12526=>"111011101",
    12527=>"111011001",
    12528=>"101100111",
    12529=>"000100101",
    12530=>"000000000",
    12531=>"010110000",
    12532=>"001000111",
    12533=>"001101100",
    12534=>"111001001",
    12535=>"011001111",
    12536=>"000000000",
    12537=>"111111101",
    12538=>"111110000",
    12539=>"000000000",
    12540=>"000000001",
    12541=>"000101000",
    12542=>"010011111",
    12543=>"111110111",
    12544=>"111111110",
    12545=>"000000000",
    12546=>"111010011",
    12547=>"101111111",
    12548=>"111001011",
    12549=>"000000000",
    12550=>"010010100",
    12551=>"000000000",
    12552=>"000000000",
    12553=>"000000000",
    12554=>"111111111",
    12555=>"011000000",
    12556=>"000000000",
    12557=>"100100100",
    12558=>"000001111",
    12559=>"101100110",
    12560=>"111111001",
    12561=>"111111111",
    12562=>"111111011",
    12563=>"111100101",
    12564=>"111001011",
    12565=>"000000000",
    12566=>"000000000",
    12567=>"000000000",
    12568=>"111111110",
    12569=>"000000000",
    12570=>"000000000",
    12571=>"000000000",
    12572=>"011101011",
    12573=>"011111011",
    12574=>"000000000",
    12575=>"111100011",
    12576=>"000000000",
    12577=>"100000000",
    12578=>"000000000",
    12579=>"001001101",
    12580=>"001000000",
    12581=>"111111111",
    12582=>"011111111",
    12583=>"111111111",
    12584=>"111111111",
    12585=>"111111000",
    12586=>"000000000",
    12587=>"011001001",
    12588=>"100001101",
    12589=>"100011111",
    12590=>"000000000",
    12591=>"000010010",
    12592=>"010000000",
    12593=>"111111111",
    12594=>"000000000",
    12595=>"110110100",
    12596=>"000000011",
    12597=>"000000000",
    12598=>"001000000",
    12599=>"111101101",
    12600=>"000000000",
    12601=>"001000000",
    12602=>"000000000",
    12603=>"000000000",
    12604=>"111010000",
    12605=>"000000000",
    12606=>"000000000",
    12607=>"000000000",
    12608=>"000000011",
    12609=>"000000000",
    12610=>"111111111",
    12611=>"000010010",
    12612=>"011111110",
    12613=>"111111111",
    12614=>"000000100",
    12615=>"000000000",
    12616=>"111111110",
    12617=>"011000000",
    12618=>"111111110",
    12619=>"000010000",
    12620=>"110111111",
    12621=>"001111111",
    12622=>"110010100",
    12623=>"110110111",
    12624=>"111111111",
    12625=>"111001100",
    12626=>"111001001",
    12627=>"111111111",
    12628=>"111111111",
    12629=>"111101101",
    12630=>"000000000",
    12631=>"000000000",
    12632=>"111101000",
    12633=>"000000000",
    12634=>"000000000",
    12635=>"111111111",
    12636=>"100100100",
    12637=>"001100010",
    12638=>"000000000",
    12639=>"111111111",
    12640=>"000000000",
    12641=>"111111111",
    12642=>"111111111",
    12643=>"000010110",
    12644=>"000000000",
    12645=>"010010000",
    12646=>"111100000",
    12647=>"111100000",
    12648=>"111001000",
    12649=>"001000000",
    12650=>"101100101",
    12651=>"000000011",
    12652=>"111111101",
    12653=>"111101111",
    12654=>"000000101",
    12655=>"000100111",
    12656=>"111111111",
    12657=>"100111000",
    12658=>"000010000",
    12659=>"010110001",
    12660=>"111101101",
    12661=>"000000000",
    12662=>"000000000",
    12663=>"000000000",
    12664=>"111111111",
    12665=>"010000000",
    12666=>"010000000",
    12667=>"111111000",
    12668=>"000000000",
    12669=>"000000000",
    12670=>"111111111",
    12671=>"000000110",
    12672=>"001001001",
    12673=>"001001001",
    12674=>"111110111",
    12675=>"100110101",
    12676=>"101000011",
    12677=>"001011010",
    12678=>"001001001",
    12679=>"110100110",
    12680=>"111101011",
    12681=>"000110000",
    12682=>"010010010",
    12683=>"111010010",
    12684=>"110110110",
    12685=>"100011100",
    12686=>"111001000",
    12687=>"110110110",
    12688=>"100000111",
    12689=>"010000001",
    12690=>"111100000",
    12691=>"000000000",
    12692=>"011010011",
    12693=>"010011000",
    12694=>"000000110",
    12695=>"100110100",
    12696=>"100010010",
    12697=>"000100010",
    12698=>"001001101",
    12699=>"011110001",
    12700=>"111011001",
    12701=>"011000100",
    12702=>"100000000",
    12703=>"010111111",
    12704=>"010111110",
    12705=>"010000000",
    12706=>"110010000",
    12707=>"000000001",
    12708=>"110110110",
    12709=>"100110011",
    12710=>"111011010",
    12711=>"011011001",
    12712=>"101101011",
    12713=>"111001111",
    12714=>"001001001",
    12715=>"011000000",
    12716=>"001110110",
    12717=>"000011111",
    12718=>"111110111",
    12719=>"110111110",
    12720=>"001001010",
    12721=>"100110110",
    12722=>"111110110",
    12723=>"110110110",
    12724=>"001101001",
    12725=>"000000001",
    12726=>"010110110",
    12727=>"110000010",
    12728=>"001010110",
    12729=>"001111100",
    12730=>"111100110",
    12731=>"010110110",
    12732=>"111001100",
    12733=>"111100000",
    12734=>"110000100",
    12735=>"001101001",
    12736=>"000011011",
    12737=>"110110000",
    12738=>"000100100",
    12739=>"001010000",
    12740=>"100110110",
    12741=>"010101111",
    12742=>"000111000",
    12743=>"001011001",
    12744=>"010010000",
    12745=>"001001001",
    12746=>"000110110",
    12747=>"100001000",
    12748=>"110110011",
    12749=>"101000000",
    12750=>"010110110",
    12751=>"110000110",
    12752=>"001001010",
    12753=>"111001100",
    12754=>"000100101",
    12755=>"001111011",
    12756=>"111001000",
    12757=>"100110110",
    12758=>"110100000",
    12759=>"110110110",
    12760=>"100000000",
    12761=>"111100010",
    12762=>"101001001",
    12763=>"100010100",
    12764=>"000000001",
    12765=>"001000101",
    12766=>"011001001",
    12767=>"000011001",
    12768=>"000000000",
    12769=>"111110010",
    12770=>"111111101",
    12771=>"000011001",
    12772=>"010100000",
    12773=>"011011111",
    12774=>"010010110",
    12775=>"111110111",
    12776=>"011001100",
    12777=>"100100100",
    12778=>"010000010",
    12779=>"001110111",
    12780=>"100010110",
    12781=>"010110010",
    12782=>"000000111",
    12783=>"001001111",
    12784=>"110110110",
    12785=>"001001100",
    12786=>"001001001",
    12787=>"100111111",
    12788=>"110110110",
    12789=>"100000000",
    12790=>"001001001",
    12791=>"110110110",
    12792=>"110110111",
    12793=>"000011111",
    12794=>"001011011",
    12795=>"110100110",
    12796=>"100101101",
    12797=>"110001001",
    12798=>"110110000",
    12799=>"110110111",
    12800=>"011011011",
    12801=>"000000001",
    12802=>"110110111",
    12803=>"110110110",
    12804=>"110011010",
    12805=>"011111101",
    12806=>"001011011",
    12807=>"001101101",
    12808=>"111001100",
    12809=>"011001111",
    12810=>"000000010",
    12811=>"100100100",
    12812=>"001001000",
    12813=>"000011000",
    12814=>"011010110",
    12815=>"001101100",
    12816=>"000111011",
    12817=>"000000100",
    12818=>"110110110",
    12819=>"011010010",
    12820=>"111110110",
    12821=>"111110111",
    12822=>"001000001",
    12823=>"001101000",
    12824=>"010010110",
    12825=>"011010111",
    12826=>"110110010",
    12827=>"100100000",
    12828=>"010000010",
    12829=>"011010010",
    12830=>"010011011",
    12831=>"111110110",
    12832=>"110000000",
    12833=>"010010111",
    12834=>"110010010",
    12835=>"010100101",
    12836=>"001001000",
    12837=>"001010011",
    12838=>"010101001",
    12839=>"010010010",
    12840=>"111110010",
    12841=>"010110111",
    12842=>"110110110",
    12843=>"010110010",
    12844=>"110010011",
    12845=>"000110110",
    12846=>"000000101",
    12847=>"110111110",
    12848=>"001011011",
    12849=>"000001000",
    12850=>"111011011",
    12851=>"000100000",
    12852=>"110011011",
    12853=>"101000100",
    12854=>"101100100",
    12855=>"110111111",
    12856=>"000100100",
    12857=>"111110010",
    12858=>"100100100",
    12859=>"000001100",
    12860=>"111100000",
    12861=>"010101101",
    12862=>"111010111",
    12863=>"010011010",
    12864=>"000000000",
    12865=>"100110111",
    12866=>"111101001",
    12867=>"000100000",
    12868=>"110110000",
    12869=>"101001111",
    12870=>"011011101",
    12871=>"101111001",
    12872=>"001001010",
    12873=>"000000000",
    12874=>"110011001",
    12875=>"000000000",
    12876=>"000100110",
    12877=>"010110000",
    12878=>"111111100",
    12879=>"001001101",
    12880=>"000111001",
    12881=>"001001001",
    12882=>"111010001",
    12883=>"000011100",
    12884=>"001101111",
    12885=>"101101101",
    12886=>"011001001",
    12887=>"001100000",
    12888=>"110010110",
    12889=>"001011111",
    12890=>"100100100",
    12891=>"001001001",
    12892=>"010010010",
    12893=>"100000000",
    12894=>"110111010",
    12895=>"001001000",
    12896=>"011001001",
    12897=>"001101000",
    12898=>"101101101",
    12899=>"111011010",
    12900=>"111000011",
    12901=>"001100010",
    12902=>"000001000",
    12903=>"000000111",
    12904=>"100000000",
    12905=>"010010010",
    12906=>"010010010",
    12907=>"001000001",
    12908=>"100001001",
    12909=>"100100000",
    12910=>"010010001",
    12911=>"111000010",
    12912=>"101101100",
    12913=>"000000001",
    12914=>"000000100",
    12915=>"001111110",
    12916=>"111100111",
    12917=>"000000000",
    12918=>"001000001",
    12919=>"111100100",
    12920=>"000000010",
    12921=>"101100101",
    12922=>"001000000",
    12923=>"101101011",
    12924=>"111011111",
    12925=>"000100101",
    12926=>"110110100",
    12927=>"011110111",
    12928=>"000000001",
    12929=>"000100100",
    12930=>"000110110",
    12931=>"101101000",
    12932=>"111011011",
    12933=>"100101100",
    12934=>"111000000",
    12935=>"111001100",
    12936=>"100001000",
    12937=>"001001010",
    12938=>"000101111",
    12939=>"011011100",
    12940=>"100110100",
    12941=>"101001000",
    12942=>"000111110",
    12943=>"001001101",
    12944=>"000101011",
    12945=>"000100000",
    12946=>"001001101",
    12947=>"100001101",
    12948=>"100100000",
    12949=>"101000000",
    12950=>"000001000",
    12951=>"001010010",
    12952=>"011001111",
    12953=>"001001101",
    12954=>"100101011",
    12955=>"110110100",
    12956=>"000101101",
    12957=>"001110111",
    12958=>"111110000",
    12959=>"011000101",
    12960=>"101011100",
    12961=>"100110000",
    12962=>"011011000",
    12963=>"111000111",
    12964=>"001110110",
    12965=>"000100100",
    12966=>"101001110",
    12967=>"111011101",
    12968=>"000000000",
    12969=>"001001001",
    12970=>"111011100",
    12971=>"111001001",
    12972=>"100101110",
    12973=>"111010011",
    12974=>"000010010",
    12975=>"100001111",
    12976=>"001011010",
    12977=>"000000001",
    12978=>"001100111",
    12979=>"101110010",
    12980=>"110100100",
    12981=>"100110100",
    12982=>"000110100",
    12983=>"111100100",
    12984=>"101111111",
    12985=>"000110111",
    12986=>"111001110",
    12987=>"101110110",
    12988=>"001001111",
    12989=>"110010011",
    12990=>"001110101",
    12991=>"110111011",
    12992=>"110110000",
    12993=>"111111011",
    12994=>"000011100",
    12995=>"001001001",
    12996=>"100110010",
    12997=>"110111111",
    12998=>"000000100",
    12999=>"101100010",
    13000=>"101011001",
    13001=>"111110110",
    13002=>"110010000",
    13003=>"001000000",
    13004=>"000111110",
    13005=>"011001111",
    13006=>"010000110",
    13007=>"001001011",
    13008=>"001001011",
    13009=>"110001001",
    13010=>"000000110",
    13011=>"111110000",
    13012=>"101111100",
    13013=>"110100110",
    13014=>"100110111",
    13015=>"100110111",
    13016=>"010110000",
    13017=>"111100001",
    13018=>"001010000",
    13019=>"001001001",
    13020=>"001001011",
    13021=>"111001010",
    13022=>"001000001",
    13023=>"001001111",
    13024=>"000000001",
    13025=>"100001101",
    13026=>"000101001",
    13027=>"100001000",
    13028=>"001000101",
    13029=>"000101010",
    13030=>"001000001",
    13031=>"001011111",
    13032=>"000101000",
    13033=>"001000000",
    13034=>"100111000",
    13035=>"110000001",
    13036=>"100000000",
    13037=>"011000000",
    13038=>"101011110",
    13039=>"111100100",
    13040=>"001000111",
    13041=>"011111111",
    13042=>"001001011",
    13043=>"000111100",
    13044=>"101001001",
    13045=>"001101111",
    13046=>"111001000",
    13047=>"001011111",
    13048=>"000000110",
    13049=>"000001111",
    13050=>"001101101",
    13051=>"111111111",
    13052=>"001001001",
    13053=>"001101110",
    13054=>"011000000",
    13055=>"101101100",
    13056=>"000000001",
    13057=>"000011011",
    13058=>"101101111",
    13059=>"001101111",
    13060=>"011011111",
    13061=>"011000110",
    13062=>"110100110",
    13063=>"111011000",
    13064=>"101101001",
    13065=>"111110110",
    13066=>"111110101",
    13067=>"110111101",
    13068=>"000011000",
    13069=>"010100111",
    13070=>"111110110",
    13071=>"000000000",
    13072=>"001100100",
    13073=>"000000101",
    13074=>"111001000",
    13075=>"000110100",
    13076=>"010100100",
    13077=>"000000000",
    13078=>"000001100",
    13079=>"011111011",
    13080=>"011000001",
    13081=>"111110100",
    13082=>"011011100",
    13083=>"000011111",
    13084=>"000000100",
    13085=>"000101000",
    13086=>"111110111",
    13087=>"000000100",
    13088=>"001111000",
    13089=>"000000000",
    13090=>"011101111",
    13091=>"000011011",
    13092=>"011011010",
    13093=>"000000000",
    13094=>"111100000",
    13095=>"000100100",
    13096=>"111000000",
    13097=>"111001011",
    13098=>"001000000",
    13099=>"001000000",
    13100=>"011000100",
    13101=>"010011000",
    13102=>"001000111",
    13103=>"000000101",
    13104=>"011111111",
    13105=>"000110111",
    13106=>"111101101",
    13107=>"000000000",
    13108=>"110110101",
    13109=>"111101011",
    13110=>"011111011",
    13111=>"111100000",
    13112=>"010000100",
    13113=>"001110111",
    13114=>"011011001",
    13115=>"110100000",
    13116=>"100100000",
    13117=>"011100101",
    13118=>"000011111",
    13119=>"011110100",
    13120=>"010110000",
    13121=>"000111111",
    13122=>"000111110",
    13123=>"100000000",
    13124=>"011010001",
    13125=>"110101010",
    13126=>"010111011",
    13127=>"010000000",
    13128=>"110100000",
    13129=>"011111111",
    13130=>"111000010",
    13131=>"000000000",
    13132=>"101111100",
    13133=>"011101111",
    13134=>"000100000",
    13135=>"000000101",
    13136=>"000011010",
    13137=>"111111100",
    13138=>"111100000",
    13139=>"101110000",
    13140=>"000011000",
    13141=>"101000000",
    13142=>"100111011",
    13143=>"011000001",
    13144=>"101111100",
    13145=>"111111110",
    13146=>"111101000",
    13147=>"110100111",
    13148=>"110001000",
    13149=>"001000110",
    13150=>"011001000",
    13151=>"110100111",
    13152=>"110110010",
    13153=>"000000000",
    13154=>"000000000",
    13155=>"111101111",
    13156=>"000011111",
    13157=>"000011011",
    13158=>"111111000",
    13159=>"010011101",
    13160=>"011011011",
    13161=>"111100100",
    13162=>"100101111",
    13163=>"000101111",
    13164=>"000010000",
    13165=>"010000000",
    13166=>"000000111",
    13167=>"111001011",
    13168=>"000000001",
    13169=>"111000111",
    13170=>"000100000",
    13171=>"000011010",
    13172=>"010000000",
    13173=>"100000000",
    13174=>"000000010",
    13175=>"111110011",
    13176=>"101000000",
    13177=>"000000101",
    13178=>"010110010",
    13179=>"111000000",
    13180=>"000110110",
    13181=>"010111110",
    13182=>"111111101",
    13183=>"110111111",
    13184=>"111101000",
    13185=>"101010100",
    13186=>"000000101",
    13187=>"000100011",
    13188=>"011111100",
    13189=>"101111000",
    13190=>"010010000",
    13191=>"111000000",
    13192=>"100110110",
    13193=>"000100000",
    13194=>"111001001",
    13195=>"111011011",
    13196=>"000000000",
    13197=>"110111110",
    13198=>"001110011",
    13199=>"111000000",
    13200=>"010010000",
    13201=>"010010000",
    13202=>"000111000",
    13203=>"100100000",
    13204=>"010010010",
    13205=>"110000000",
    13206=>"000000000",
    13207=>"011000000",
    13208=>"100111111",
    13209=>"110101011",
    13210=>"001000101",
    13211=>"001011011",
    13212=>"110111111",
    13213=>"110111111",
    13214=>"011111111",
    13215=>"010111111",
    13216=>"001011001",
    13217=>"000111011",
    13218=>"010001000",
    13219=>"111111111",
    13220=>"000111001",
    13221=>"011010000",
    13222=>"000001100",
    13223=>"000111111",
    13224=>"111010110",
    13225=>"110111111",
    13226=>"111000000",
    13227=>"000001111",
    13228=>"010100110",
    13229=>"011011010",
    13230=>"111100110",
    13231=>"101000101",
    13232=>"110011000",
    13233=>"001000110",
    13234=>"110011001",
    13235=>"000011110",
    13236=>"100100100",
    13237=>"010000000",
    13238=>"011000000",
    13239=>"000101111",
    13240=>"111001001",
    13241=>"010100000",
    13242=>"011011001",
    13243=>"111101000",
    13244=>"100000000",
    13245=>"100111101",
    13246=>"100100100",
    13247=>"110100001",
    13248=>"011000000",
    13249=>"000000010",
    13250=>"011111111",
    13251=>"101000000",
    13252=>"100001010",
    13253=>"000110100",
    13254=>"111000000",
    13255=>"111111110",
    13256=>"010110010",
    13257=>"010111111",
    13258=>"000000110",
    13259=>"000000001",
    13260=>"000000111",
    13261=>"111111000",
    13262=>"000010001",
    13263=>"000000111",
    13264=>"000011010",
    13265=>"100000001",
    13266=>"010010011",
    13267=>"011111011",
    13268=>"000011001",
    13269=>"011010010",
    13270=>"000110000",
    13271=>"111101101",
    13272=>"011111111",
    13273=>"000000000",
    13274=>"001001001",
    13275=>"000010010",
    13276=>"100101001",
    13277=>"011001100",
    13278=>"101000000",
    13279=>"001000000",
    13280=>"010011011",
    13281=>"010110000",
    13282=>"001010011",
    13283=>"011011101",
    13284=>"011001000",
    13285=>"000000000",
    13286=>"001000000",
    13287=>"001101011",
    13288=>"111100000",
    13289=>"111101000",
    13290=>"001101101",
    13291=>"000000010",
    13292=>"000000000",
    13293=>"100001001",
    13294=>"111100000",
    13295=>"001011111",
    13296=>"000000000",
    13297=>"000000111",
    13298=>"001111111",
    13299=>"110111011",
    13300=>"001000000",
    13301=>"000111011",
    13302=>"100101000",
    13303=>"011110001",
    13304=>"111111111",
    13305=>"111111101",
    13306=>"110101000",
    13307=>"000000000",
    13308=>"100100101",
    13309=>"000111111",
    13310=>"111010000",
    13311=>"100001011",
    13312=>"000111111",
    13313=>"000000111",
    13314=>"000100111",
    13315=>"001111111",
    13316=>"000001101",
    13317=>"010111100",
    13318=>"001010011",
    13319=>"011110100",
    13320=>"000001011",
    13321=>"100000000",
    13322=>"101111000",
    13323=>"011011000",
    13324=>"000110000",
    13325=>"100110110",
    13326=>"111110111",
    13327=>"111100001",
    13328=>"100110110",
    13329=>"111000111",
    13330=>"111111110",
    13331=>"000110111",
    13332=>"111001111",
    13333=>"111100000",
    13334=>"000001000",
    13335=>"110000000",
    13336=>"111011011",
    13337=>"101110100",
    13338=>"111111100",
    13339=>"011111111",
    13340=>"111110001",
    13341=>"100100110",
    13342=>"111110100",
    13343=>"111001000",
    13344=>"010010110",
    13345=>"001110100",
    13346=>"011001001",
    13347=>"110001101",
    13348=>"000011000",
    13349=>"000000111",
    13350=>"111001100",
    13351=>"111101000",
    13352=>"000000000",
    13353=>"110100111",
    13354=>"100101001",
    13355=>"001101101",
    13356=>"100000000",
    13357=>"010000110",
    13358=>"010000000",
    13359=>"000000110",
    13360=>"000000000",
    13361=>"011011111",
    13362=>"001001001",
    13363=>"100100110",
    13364=>"000100000",
    13365=>"000001101",
    13366=>"000000111",
    13367=>"000111111",
    13368=>"101111001",
    13369=>"000000111",
    13370=>"001000000",
    13371=>"111010000",
    13372=>"100000000",
    13373=>"010010100",
    13374=>"110110100",
    13375=>"001000000",
    13376=>"111010000",
    13377=>"111000000",
    13378=>"100100111",
    13379=>"101000000",
    13380=>"110101110",
    13381=>"001011010",
    13382=>"000001110",
    13383=>"111111110",
    13384=>"001011011",
    13385=>"110110000",
    13386=>"000010111",
    13387=>"001101000",
    13388=>"010001000",
    13389=>"111100100",
    13390=>"101101111",
    13391=>"000001111",
    13392=>"111100000",
    13393=>"100100111",
    13394=>"000000111",
    13395=>"000111001",
    13396=>"100110110",
    13397=>"111101001",
    13398=>"001001111",
    13399=>"011111010",
    13400=>"100111111",
    13401=>"000000000",
    13402=>"001001000",
    13403=>"101100011",
    13404=>"100110110",
    13405=>"000000100",
    13406=>"001001111",
    13407=>"000110010",
    13408=>"100110110",
    13409=>"011011011",
    13410=>"101111110",
    13411=>"001000100",
    13412=>"111001001",
    13413=>"100001111",
    13414=>"001001111",
    13415=>"100000010",
    13416=>"101010000",
    13417=>"100100110",
    13418=>"000111111",
    13419=>"111010010",
    13420=>"000000111",
    13421=>"100000100",
    13422=>"111010010",
    13423=>"100010111",
    13424=>"000000111",
    13425=>"010110001",
    13426=>"111111101",
    13427=>"100001111",
    13428=>"111111000",
    13429=>"000000000",
    13430=>"011001000",
    13431=>"110000100",
    13432=>"010000000",
    13433=>"001100000",
    13434=>"110000000",
    13435=>"000011111",
    13436=>"111011010",
    13437=>"111010111",
    13438=>"000000001",
    13439=>"111100010",
    13440=>"101000000",
    13441=>"111000000",
    13442=>"000111010",
    13443=>"101001010",
    13444=>"111100000",
    13445=>"111000000",
    13446=>"111000001",
    13447=>"001111110",
    13448=>"100000001",
    13449=>"001001011",
    13450=>"001001010",
    13451=>"111110111",
    13452=>"000000111",
    13453=>"110111100",
    13454=>"000011111",
    13455=>"100110110",
    13456=>"001011111",
    13457=>"111000000",
    13458=>"001011001",
    13459=>"011101100",
    13460=>"000100001",
    13461=>"000000111",
    13462=>"000000000",
    13463=>"111010110",
    13464=>"010110000",
    13465=>"001001111",
    13466=>"101001011",
    13467=>"110110100",
    13468=>"110010000",
    13469=>"011011110",
    13470=>"011011000",
    13471=>"111110111",
    13472=>"000000000",
    13473=>"001100100",
    13474=>"000100111",
    13475=>"000000101",
    13476=>"000000000",
    13477=>"100001101",
    13478=>"111001000",
    13479=>"110000001",
    13480=>"100000001",
    13481=>"101000000",
    13482=>"110001001",
    13483=>"111111000",
    13484=>"111011001",
    13485=>"101001001",
    13486=>"111001000",
    13487=>"101111110",
    13488=>"000000101",
    13489=>"000111111",
    13490=>"001111111",
    13491=>"000111001",
    13492=>"101001001",
    13493=>"000000101",
    13494=>"001001011",
    13495=>"001011000",
    13496=>"110010111",
    13497=>"110110010",
    13498=>"100100100",
    13499=>"000000110",
    13500=>"111000001",
    13501=>"000000000",
    13502=>"000110011",
    13503=>"100111111",
    13504=>"111001001",
    13505=>"010010101",
    13506=>"000010111",
    13507=>"111000000",
    13508=>"000110110",
    13509=>"110011111",
    13510=>"111101101",
    13511=>"110110000",
    13512=>"000100110",
    13513=>"110000000",
    13514=>"111110111",
    13515=>"001000100",
    13516=>"000111110",
    13517=>"111111101",
    13518=>"001111000",
    13519=>"000110010",
    13520=>"001001111",
    13521=>"101000111",
    13522=>"111110000",
    13523=>"100111000",
    13524=>"111111110",
    13525=>"000011101",
    13526=>"000000000",
    13527=>"000111111",
    13528=>"011100000",
    13529=>"000000000",
    13530=>"011101001",
    13531=>"110110000",
    13532=>"111101000",
    13533=>"000101010",
    13534=>"111110100",
    13535=>"111110000",
    13536=>"011000000",
    13537=>"100100101",
    13538=>"000111111",
    13539=>"101000110",
    13540=>"110000000",
    13541=>"001000100",
    13542=>"000000111",
    13543=>"110111111",
    13544=>"111100100",
    13545=>"000000010",
    13546=>"110000000",
    13547=>"111101001",
    13548=>"101001111",
    13549=>"101101111",
    13550=>"111111111",
    13551=>"111110011",
    13552=>"000101111",
    13553=>"011000000",
    13554=>"111000000",
    13555=>"000000010",
    13556=>"000000001",
    13557=>"001000110",
    13558=>"011001000",
    13559=>"000111110",
    13560=>"000010111",
    13561=>"001000100",
    13562=>"011001011",
    13563=>"001011110",
    13564=>"111011001",
    13565=>"111111101",
    13566=>"101101111",
    13567=>"111111111",
    13568=>"111111111",
    13569=>"010010000",
    13570=>"101111011",
    13571=>"110111000",
    13572=>"010000000",
    13573=>"000100010",
    13574=>"000000000",
    13575=>"000000000",
    13576=>"011111110",
    13577=>"011000000",
    13578=>"101101111",
    13579=>"110001110",
    13580=>"011110011",
    13581=>"110111111",
    13582=>"011111101",
    13583=>"011111111",
    13584=>"111000000",
    13585=>"000000100",
    13586=>"110001000",
    13587=>"000001000",
    13588=>"000000111",
    13589=>"111000000",
    13590=>"010000000",
    13591=>"111001101",
    13592=>"010100100",
    13593=>"111110101",
    13594=>"100000100",
    13595=>"110011011",
    13596=>"000000111",
    13597=>"011111010",
    13598=>"000110111",
    13599=>"111110111",
    13600=>"001101111",
    13601=>"110100100",
    13602=>"010001101",
    13603=>"000000100",
    13604=>"101001000",
    13605=>"111000000",
    13606=>"000011010",
    13607=>"100101111",
    13608=>"111111111",
    13609=>"100000000",
    13610=>"101110110",
    13611=>"011000000",
    13612=>"111111111",
    13613=>"111010010",
    13614=>"111000000",
    13615=>"000111111",
    13616=>"111000001",
    13617=>"000000111",
    13618=>"110000010",
    13619=>"100100111",
    13620=>"111101100",
    13621=>"111000000",
    13622=>"111000000",
    13623=>"110111010",
    13624=>"000000000",
    13625=>"100101111",
    13626=>"100100000",
    13627=>"000111111",
    13628=>"110110000",
    13629=>"111111000",
    13630=>"011101100",
    13631=>"010000101",
    13632=>"001011111",
    13633=>"011110000",
    13634=>"111001010",
    13635=>"111111001",
    13636=>"011111111",
    13637=>"010010000",
    13638=>"110000000",
    13639=>"001000000",
    13640=>"111010000",
    13641=>"111010000",
    13642=>"000000000",
    13643=>"111000000",
    13644=>"000000101",
    13645=>"101001111",
    13646=>"000000000",
    13647=>"000001111",
    13648=>"010000000",
    13649=>"000010001",
    13650=>"000100100",
    13651=>"111011111",
    13652=>"111110001",
    13653=>"101101000",
    13654=>"000000001",
    13655=>"101111111",
    13656=>"001100000",
    13657=>"111000000",
    13658=>"010101101",
    13659=>"111111000",
    13660=>"011111000",
    13661=>"000100000",
    13662=>"101100100",
    13663=>"111111010",
    13664=>"111101001",
    13665=>"011001110",
    13666=>"001111111",
    13667=>"111000000",
    13668=>"011111111",
    13669=>"110000000",
    13670=>"100000000",
    13671=>"010000000",
    13672=>"000010000",
    13673=>"100100111",
    13674=>"100000000",
    13675=>"101001111",
    13676=>"000000001",
    13677=>"011111000",
    13678=>"011100001",
    13679=>"110011101",
    13680=>"101000111",
    13681=>"000000000",
    13682=>"111000000",
    13683=>"010011010",
    13684=>"110101100",
    13685=>"000000000",
    13686=>"111111111",
    13687=>"011011000",
    13688=>"111111111",
    13689=>"111100000",
    13690=>"010111001",
    13691=>"011011000",
    13692=>"011111101",
    13693=>"000010111",
    13694=>"000001111",
    13695=>"000000101",
    13696=>"110010011",
    13697=>"101100100",
    13698=>"101101111",
    13699=>"000011110",
    13700=>"000011011",
    13701=>"101011010",
    13702=>"000011011",
    13703=>"111000101",
    13704=>"001011110",
    13705=>"110110111",
    13706=>"111001001",
    13707=>"111110111",
    13708=>"100111011",
    13709=>"111110100",
    13710=>"000100111",
    13711=>"100100101",
    13712=>"100101110",
    13713=>"111101000",
    13714=>"001001100",
    13715=>"100110111",
    13716=>"111001000",
    13717=>"111010000",
    13718=>"000000100",
    13719=>"110000110",
    13720=>"100100001",
    13721=>"111010100",
    13722=>"000101100",
    13723=>"000000100",
    13724=>"101001110",
    13725=>"011010001",
    13726=>"011111100",
    13727=>"011110101",
    13728=>"001111101",
    13729=>"000100001",
    13730=>"111011000",
    13731=>"000101101",
    13732=>"011011110",
    13733=>"110101000",
    13734=>"101101101",
    13735=>"101101111",
    13736=>"011010000",
    13737=>"110101101",
    13738=>"000000001",
    13739=>"100101110",
    13740=>"111001001",
    13741=>"010000000",
    13742=>"000010000",
    13743=>"111010101",
    13744=>"010111110",
    13745=>"010000111",
    13746=>"001001010",
    13747=>"010001010",
    13748=>"000001110",
    13749=>"000000000",
    13750=>"000000000",
    13751=>"111111001",
    13752=>"101101100",
    13753=>"000011101",
    13754=>"011011011",
    13755=>"000000000",
    13756=>"101000000",
    13757=>"000010011",
    13758=>"100000000",
    13759=>"001000011",
    13760=>"111000000",
    13761=>"000001011",
    13762=>"111101000",
    13763=>"001000100",
    13764=>"101111111",
    13765=>"001011110",
    13766=>"111101101",
    13767=>"000101000",
    13768=>"000100011",
    13769=>"101011010",
    13770=>"001001101",
    13771=>"111000101",
    13772=>"000010000",
    13773=>"111111111",
    13774=>"011010010",
    13775=>"100000011",
    13776=>"000000111",
    13777=>"100100000",
    13778=>"011101101",
    13779=>"011110011",
    13780=>"100010011",
    13781=>"100000101",
    13782=>"101100100",
    13783=>"000100000",
    13784=>"111100001",
    13785=>"111111111",
    13786=>"100101111",
    13787=>"111100000",
    13788=>"001110010",
    13789=>"000001100",
    13790=>"001001101",
    13791=>"111000000",
    13792=>"100101011",
    13793=>"100100010",
    13794=>"111001011",
    13795=>"111000100",
    13796=>"111111010",
    13797=>"110111000",
    13798=>"101001010",
    13799=>"010110110",
    13800=>"100001111",
    13801=>"000100000",
    13802=>"100101010",
    13803=>"010111101",
    13804=>"000011010",
    13805=>"000000100",
    13806=>"111111010",
    13807=>"110000001",
    13808=>"010000000",
    13809=>"011111111",
    13810=>"111110000",
    13811=>"111101000",
    13812=>"111101111",
    13813=>"100100111",
    13814=>"010000000",
    13815=>"000000000",
    13816=>"010000000",
    13817=>"010000100",
    13818=>"100100111",
    13819=>"100100000",
    13820=>"100110111",
    13821=>"011111110",
    13822=>"111011000",
    13823=>"110111000",
    13824=>"010010000",
    13825=>"100011000",
    13826=>"111101100",
    13827=>"100010000",
    13828=>"010000000",
    13829=>"000000000",
    13830=>"101101010",
    13831=>"101111111",
    13832=>"111111001",
    13833=>"111111111",
    13834=>"101101111",
    13835=>"111110010",
    13836=>"000000000",
    13837=>"111111110",
    13838=>"000000000",
    13839=>"000111110",
    13840=>"010000000",
    13841=>"010000000",
    13842=>"100110111",
    13843=>"000000010",
    13844=>"000000100",
    13845=>"000000111",
    13846=>"000000000",
    13847=>"000010010",
    13848=>"011111000",
    13849=>"110001001",
    13850=>"111110001",
    13851=>"100100110",
    13852=>"000000001",
    13853=>"100100111",
    13854=>"110111111",
    13855=>"011111111",
    13856=>"011000000",
    13857=>"111110111",
    13858=>"001101010",
    13859=>"111101011",
    13860=>"011011000",
    13861=>"000000000",
    13862=>"000000101",
    13863=>"000000000",
    13864=>"011000000",
    13865=>"000000000",
    13866=>"001000001",
    13867=>"011001000",
    13868=>"000001111",
    13869=>"111000111",
    13870=>"010010000",
    13871=>"111111111",
    13872=>"111110111",
    13873=>"000000000",
    13874=>"001000110",
    13875=>"001011010",
    13876=>"011001000",
    13877=>"101111111",
    13878=>"100000000",
    13879=>"001011101",
    13880=>"111101110",
    13881=>"011111111",
    13882=>"111111110",
    13883=>"001100101",
    13884=>"000100000",
    13885=>"000000111",
    13886=>"000001000",
    13887=>"100100111",
    13888=>"010000000",
    13889=>"011111111",
    13890=>"011000111",
    13891=>"000000101",
    13892=>"111111011",
    13893=>"110110101",
    13894=>"100000010",
    13895=>"111011111",
    13896=>"001011001",
    13897=>"000100111",
    13898=>"110011110",
    13899=>"000000101",
    13900=>"111111111",
    13901=>"011000000",
    13902=>"100011111",
    13903=>"000100111",
    13904=>"010000000",
    13905=>"000000010",
    13906=>"000000011",
    13907=>"100000000",
    13908=>"011011100",
    13909=>"000101101",
    13910=>"000000000",
    13911=>"111111111",
    13912=>"001001000",
    13913=>"010110110",
    13914=>"011011000",
    13915=>"010010000",
    13916=>"110100000",
    13917=>"001100010",
    13918=>"001100100",
    13919=>"100100111",
    13920=>"011000100",
    13921=>"000110111",
    13922=>"000000000",
    13923=>"010011010",
    13924=>"010001000",
    13925=>"011100000",
    13926=>"000000010",
    13927=>"110000010",
    13928=>"010111110",
    13929=>"100100011",
    13930=>"111011010",
    13931=>"111001100",
    13932=>"110100100",
    13933=>"101000011",
    13934=>"000000000",
    13935=>"001000110",
    13936=>"000000000",
    13937=>"001000011",
    13938=>"111011010",
    13939=>"001000111",
    13940=>"101101111",
    13941=>"010000000",
    13942=>"111111100",
    13943=>"000000111",
    13944=>"000000000",
    13945=>"111111011",
    13946=>"000111001",
    13947=>"111011010",
    13948=>"110100000",
    13949=>"110011011",
    13950=>"101100111",
    13951=>"100001011",
    13952=>"111111111",
    13953=>"010111000",
    13954=>"111111111",
    13955=>"111111011",
    13956=>"101100100",
    13957=>"010010000",
    13958=>"111111010",
    13959=>"110010110",
    13960=>"111111011",
    13961=>"111000111",
    13962=>"111001100",
    13963=>"000000000",
    13964=>"000000000",
    13965=>"110111110",
    13966=>"101111111",
    13967=>"010011011",
    13968=>"000000000",
    13969=>"010000111",
    13970=>"001110000",
    13971=>"110000110",
    13972=>"010011111",
    13973=>"100000010",
    13974=>"000100101",
    13975=>"010000110",
    13976=>"100100101",
    13977=>"000000000",
    13978=>"111101101",
    13979=>"100110100",
    13980=>"101000000",
    13981=>"000000101",
    13982=>"001111110",
    13983=>"110111111",
    13984=>"100001111",
    13985=>"110101000",
    13986=>"111111001",
    13987=>"111101101",
    13988=>"011111111",
    13989=>"001111111",
    13990=>"000110010",
    13991=>"101000101",
    13992=>"111010110",
    13993=>"110000001",
    13994=>"001001000",
    13995=>"100101101",
    13996=>"001010101",
    13997=>"000110110",
    13998=>"001000111",
    13999=>"101011000",
    14000=>"110111111",
    14001=>"011000111",
    14002=>"000000000",
    14003=>"110111000",
    14004=>"001101101",
    14005=>"000000100",
    14006=>"011110010",
    14007=>"101011111",
    14008=>"011011011",
    14009=>"010000000",
    14010=>"101000111",
    14011=>"101101101",
    14012=>"000100100",
    14013=>"001000100",
    14014=>"001001011",
    14015=>"011111000",
    14016=>"010011101",
    14017=>"000000000",
    14018=>"111010000",
    14019=>"000111010",
    14020=>"000000000",
    14021=>"011110000",
    14022=>"111010110",
    14023=>"111111110",
    14024=>"000000100",
    14025=>"100101001",
    14026=>"111000010",
    14027=>"111000000",
    14028=>"001001001",
    14029=>"111111101",
    14030=>"110111111",
    14031=>"001001001",
    14032=>"010011010",
    14033=>"001000101",
    14034=>"111100111",
    14035=>"011000000",
    14036=>"010010100",
    14037=>"000000000",
    14038=>"000011011",
    14039=>"101000000",
    14040=>"101100001",
    14041=>"100000000",
    14042=>"010111011",
    14043=>"001010101",
    14044=>"001001001",
    14045=>"011010010",
    14046=>"000110000",
    14047=>"101010000",
    14048=>"100110101",
    14049=>"000000100",
    14050=>"000111011",
    14051=>"000000010",
    14052=>"010010111",
    14053=>"001000101",
    14054=>"000000001",
    14055=>"000010010",
    14056=>"000000000",
    14057=>"100000000",
    14058=>"101101000",
    14059=>"110010001",
    14060=>"011000000",
    14061=>"000000010",
    14062=>"111111101",
    14063=>"111101111",
    14064=>"000000000",
    14065=>"011011000",
    14066=>"100111100",
    14067=>"000000000",
    14068=>"011010010",
    14069=>"000000000",
    14070=>"110111010",
    14071=>"000000000",
    14072=>"010000110",
    14073=>"011010110",
    14074=>"010010010",
    14075=>"010010010",
    14076=>"110110111",
    14077=>"111111111",
    14078=>"110110110",
    14079=>"111111111",
    14080=>"001101110",
    14081=>"111000000",
    14082=>"000010000",
    14083=>"000000000",
    14084=>"011000000",
    14085=>"000000100",
    14086=>"000001111",
    14087=>"111111111",
    14088=>"000111111",
    14089=>"010100000",
    14090=>"111111111",
    14091=>"110111100",
    14092=>"111111001",
    14093=>"000010010",
    14094=>"110101000",
    14095=>"110110111",
    14096=>"100100100",
    14097=>"010000001",
    14098=>"011000000",
    14099=>"100100001",
    14100=>"110111110",
    14101=>"110100111",
    14102=>"111011101",
    14103=>"110101111",
    14104=>"101001000",
    14105=>"111000001",
    14106=>"010011010",
    14107=>"111001001",
    14108=>"010000000",
    14109=>"111100100",
    14110=>"000100000",
    14111=>"000000000",
    14112=>"010000010",
    14113=>"011001111",
    14114=>"011011000",
    14115=>"011111111",
    14116=>"000000111",
    14117=>"000000000",
    14118=>"001100000",
    14119=>"111111110",
    14120=>"100001110",
    14121=>"010110000",
    14122=>"101000111",
    14123=>"100100101",
    14124=>"111101101",
    14125=>"111111000",
    14126=>"101000000",
    14127=>"000000000",
    14128=>"000010111",
    14129=>"001000000",
    14130=>"011000101",
    14131=>"101000111",
    14132=>"101100000",
    14133=>"000000000",
    14134=>"000000000",
    14135=>"111111111",
    14136=>"001111111",
    14137=>"001000111",
    14138=>"001001010",
    14139=>"111111111",
    14140=>"111111111",
    14141=>"001000001",
    14142=>"001110111",
    14143=>"111111111",
    14144=>"111100000",
    14145=>"000100111",
    14146=>"000111111",
    14147=>"000000101",
    14148=>"101001011",
    14149=>"000000100",
    14150=>"110110110",
    14151=>"110000000",
    14152=>"011001000",
    14153=>"010000000",
    14154=>"001001110",
    14155=>"111000000",
    14156=>"000000001",
    14157=>"000010100",
    14158=>"000000000",
    14159=>"111111111",
    14160=>"111111000",
    14161=>"111111110",
    14162=>"010101111",
    14163=>"100100001",
    14164=>"000011011",
    14165=>"111111011",
    14166=>"000010011",
    14167=>"000010000",
    14168=>"101101110",
    14169=>"000000000",
    14170=>"110000000",
    14171=>"111111111",
    14172=>"001001001",
    14173=>"001110100",
    14174=>"011011010",
    14175=>"101111111",
    14176=>"000010010",
    14177=>"001001111",
    14178=>"001000000",
    14179=>"001001000",
    14180=>"001101110",
    14181=>"100100000",
    14182=>"011111011",
    14183=>"000001111",
    14184=>"010110011",
    14185=>"010111111",
    14186=>"100001001",
    14187=>"000000111",
    14188=>"000000001",
    14189=>"111111111",
    14190=>"111111111",
    14191=>"111110011",
    14192=>"000111111",
    14193=>"111111000",
    14194=>"111000000",
    14195=>"111111000",
    14196=>"000000000",
    14197=>"000001101",
    14198=>"000000000",
    14199=>"100111011",
    14200=>"111111111",
    14201=>"000000110",
    14202=>"111100100",
    14203=>"000000001",
    14204=>"011101001",
    14205=>"111101010",
    14206=>"110111111",
    14207=>"010110011",
    14208=>"000000000",
    14209=>"101000101",
    14210=>"000111011",
    14211=>"111111111",
    14212=>"110011000",
    14213=>"111111111",
    14214=>"100110111",
    14215=>"111011000",
    14216=>"001001000",
    14217=>"111101011",
    14218=>"000001011",
    14219=>"000000000",
    14220=>"111101000",
    14221=>"010000111",
    14222=>"110110100",
    14223=>"010110110",
    14224=>"011001000",
    14225=>"100001101",
    14226=>"001011001",
    14227=>"111110100",
    14228=>"000001011",
    14229=>"011000000",
    14230=>"001010111",
    14231=>"111111000",
    14232=>"000000000",
    14233=>"000011000",
    14234=>"101011111",
    14235=>"101100101",
    14236=>"010011111",
    14237=>"011000101",
    14238=>"001000100",
    14239=>"111111000",
    14240=>"111111000",
    14241=>"100000000",
    14242=>"111010010",
    14243=>"000000111",
    14244=>"111101000",
    14245=>"000011111",
    14246=>"010010110",
    14247=>"000111111",
    14248=>"000000000",
    14249=>"001000000",
    14250=>"111001100",
    14251=>"111100100",
    14252=>"111001000",
    14253=>"100000101",
    14254=>"110000000",
    14255=>"011111111",
    14256=>"111111000",
    14257=>"000011111",
    14258=>"110011001",
    14259=>"000100000",
    14260=>"001001000",
    14261=>"111000010",
    14262=>"110111100",
    14263=>"110111111",
    14264=>"000000011",
    14265=>"111011000",
    14266=>"111001001",
    14267=>"011111111",
    14268=>"010110000",
    14269=>"101000100",
    14270=>"111000000",
    14271=>"111111111",
    14272=>"000100100",
    14273=>"010100110",
    14274=>"010000000",
    14275=>"111001001",
    14276=>"110100000",
    14277=>"110011011",
    14278=>"101110111",
    14279=>"000000000",
    14280=>"110100000",
    14281=>"100101111",
    14282=>"010010000",
    14283=>"000000111",
    14284=>"111111000",
    14285=>"000000000",
    14286=>"111111000",
    14287=>"000010111",
    14288=>"000010010",
    14289=>"000110111",
    14290=>"010000000",
    14291=>"101111110",
    14292=>"011110100",
    14293=>"000010111",
    14294=>"111000000",
    14295=>"111000000",
    14296=>"100100111",
    14297=>"111000000",
    14298=>"010110000",
    14299=>"000010111",
    14300=>"101000001",
    14301=>"111011011",
    14302=>"110111101",
    14303=>"111110000",
    14304=>"110000000",
    14305=>"000011001",
    14306=>"110111111",
    14307=>"000000111",
    14308=>"110000000",
    14309=>"000010111",
    14310=>"001011111",
    14311=>"111111000",
    14312=>"100000110",
    14313=>"000111111",
    14314=>"111110101",
    14315=>"001100000",
    14316=>"000110111",
    14317=>"000000011",
    14318=>"111100111",
    14319=>"010001101",
    14320=>"000110011",
    14321=>"110111001",
    14322=>"000101101",
    14323=>"000111111",
    14324=>"111000000",
    14325=>"010000111",
    14326=>"000111000",
    14327=>"111100000",
    14328=>"111000000",
    14329=>"110110110",
    14330=>"011001011",
    14331=>"111110000",
    14332=>"011111111",
    14333=>"111000000",
    14334=>"100110111",
    14335=>"011010011",
    14336=>"110010110",
    14337=>"001001001",
    14338=>"001011001",
    14339=>"000100010",
    14340=>"000000000",
    14341=>"111010100",
    14342=>"000100010",
    14343=>"110000100",
    14344=>"000000000",
    14345=>"000010111",
    14346=>"001011011",
    14347=>"000100100",
    14348=>"100100000",
    14349=>"101111100",
    14350=>"000000000",
    14351=>"001001001",
    14352=>"100100111",
    14353=>"000110110",
    14354=>"111110110",
    14355=>"111111011",
    14356=>"000010001",
    14357=>"100100110",
    14358=>"000100000",
    14359=>"111100110",
    14360=>"000000000",
    14361=>"111110100",
    14362=>"100100100",
    14363=>"000010010",
    14364=>"011011111",
    14365=>"110100110",
    14366=>"001111111",
    14367=>"010100010",
    14368=>"110110001",
    14369=>"000100101",
    14370=>"101000100",
    14371=>"111111101",
    14372=>"011010011",
    14373=>"111100100",
    14374=>"110100110",
    14375=>"100100100",
    14376=>"100100100",
    14377=>"100110110",
    14378=>"010100100",
    14379=>"001011101",
    14380=>"011000000",
    14381=>"110110110",
    14382=>"000000000",
    14383=>"110100110",
    14384=>"000000011",
    14385=>"010100111",
    14386=>"000100101",
    14387=>"111010110",
    14388=>"111111011",
    14389=>"010010001",
    14390=>"001001001",
    14391=>"000001000",
    14392=>"110111011",
    14393=>"010000110",
    14394=>"110010110",
    14395=>"011011110",
    14396=>"100100100",
    14397=>"110110110",
    14398=>"010000000",
    14399=>"011101001",
    14400=>"101001011",
    14401=>"110100100",
    14402=>"100001101",
    14403=>"011011001",
    14404=>"110010110",
    14405=>"000101100",
    14406=>"001001101",
    14407=>"000100110",
    14408=>"000000000",
    14409=>"001011010",
    14410=>"000001101",
    14411=>"110110110",
    14412=>"010011001",
    14413=>"001001001",
    14414=>"100100100",
    14415=>"011011001",
    14416=>"110100100",
    14417=>"110001000",
    14418=>"000100100",
    14419=>"000110101",
    14420=>"000110110",
    14421=>"011011001",
    14422=>"110100110",
    14423=>"011111111",
    14424=>"000010001",
    14425=>"010010000",
    14426=>"001011011",
    14427=>"000001001",
    14428=>"101100111",
    14429=>"010000001",
    14430=>"101011101",
    14431=>"000100100",
    14432=>"111110111",
    14433=>"001000000",
    14434=>"001011011",
    14435=>"001001001",
    14436=>"111101001",
    14437=>"110001111",
    14438=>"100000100",
    14439=>"100001100",
    14440=>"110100101",
    14441=>"001011001",
    14442=>"000000000",
    14443=>"100100111",
    14444=>"001011011",
    14445=>"000000000",
    14446=>"011011110",
    14447=>"011111111",
    14448=>"011011001",
    14449=>"100011000",
    14450=>"010000000",
    14451=>"011001001",
    14452=>"111100111",
    14453=>"100100000",
    14454=>"011000100",
    14455=>"110110000",
    14456=>"111110000",
    14457=>"110100100",
    14458=>"001001001",
    14459=>"011001001",
    14460=>"000000001",
    14461=>"010110100",
    14462=>"000100101",
    14463=>"100100111",
    14464=>"011000000",
    14465=>"000000101",
    14466=>"011101110",
    14467=>"111101100",
    14468=>"101110111",
    14469=>"111110111",
    14470=>"111000000",
    14471=>"000111000",
    14472=>"111111111",
    14473=>"001001111",
    14474=>"000101101",
    14475=>"110011011",
    14476=>"000000000",
    14477=>"111110000",
    14478=>"000000000",
    14479=>"001100111",
    14480=>"101001010",
    14481=>"000101000",
    14482=>"011100100",
    14483=>"011111111",
    14484=>"100000000",
    14485=>"000001000",
    14486=>"000111000",
    14487=>"111000000",
    14488=>"110010000",
    14489=>"110110100",
    14490=>"111010101",
    14491=>"100000000",
    14492=>"100000000",
    14493=>"111000000",
    14494=>"111000000",
    14495=>"110111101",
    14496=>"000000001",
    14497=>"001000000",
    14498=>"010010001",
    14499=>"111111101",
    14500=>"000000000",
    14501=>"000001111",
    14502=>"010100000",
    14503=>"111000000",
    14504=>"000001000",
    14505=>"111011100",
    14506=>"000010010",
    14507=>"001000000",
    14508=>"111010000",
    14509=>"010110000",
    14510=>"101000000",
    14511=>"000111111",
    14512=>"001000010",
    14513=>"100111111",
    14514=>"101001100",
    14515=>"111111100",
    14516=>"011001111",
    14517=>"101000000",
    14518=>"000100000",
    14519=>"010010111",
    14520=>"111111101",
    14521=>"111111000",
    14522=>"110111111",
    14523=>"111111111",
    14524=>"000111111",
    14525=>"000000000",
    14526=>"001000000",
    14527=>"000001101",
    14528=>"000110111",
    14529=>"111111000",
    14530=>"000101010",
    14531=>"111001101",
    14532=>"111101001",
    14533=>"111001110",
    14534=>"101000000",
    14535=>"111101000",
    14536=>"111110010",
    14537=>"000000111",
    14538=>"111100001",
    14539=>"101111111",
    14540=>"000000000",
    14541=>"100111111",
    14542=>"000000000",
    14543=>"010010000",
    14544=>"110111000",
    14545=>"000000011",
    14546=>"111011000",
    14547=>"000101000",
    14548=>"111100100",
    14549=>"000001111",
    14550=>"100000000",
    14551=>"100000000",
    14552=>"110101101",
    14553=>"000101101",
    14554=>"111100001",
    14555=>"000101111",
    14556=>"111001011",
    14557=>"100011110",
    14558=>"111110001",
    14559=>"000111111",
    14560=>"111000101",
    14561=>"011001101",
    14562=>"011000111",
    14563=>"000110111",
    14564=>"111101000",
    14565=>"110000000",
    14566=>"000000111",
    14567=>"000011010",
    14568=>"111100000",
    14569=>"000011011",
    14570=>"111000001",
    14571=>"000010000",
    14572=>"000000111",
    14573=>"000010111",
    14574=>"101001111",
    14575=>"000010011",
    14576=>"000000000",
    14577=>"000000000",
    14578=>"011001000",
    14579=>"000110111",
    14580=>"000011111",
    14581=>"000000000",
    14582=>"000000000",
    14583=>"101110111",
    14584=>"110000000",
    14585=>"110111011",
    14586=>"000011010",
    14587=>"000110000",
    14588=>"011001100",
    14589=>"111111111",
    14590=>"001001001",
    14591=>"011100111",
    14592=>"001100110",
    14593=>"011000111",
    14594=>"101000000",
    14595=>"000111001",
    14596=>"111011111",
    14597=>"100101101",
    14598=>"101100111",
    14599=>"000111110",
    14600=>"001000100",
    14601=>"101101101",
    14602=>"011001000",
    14603=>"111111110",
    14604=>"110110010",
    14605=>"010110000",
    14606=>"001000000",
    14607=>"000000000",
    14608=>"110111011",
    14609=>"010011011",
    14610=>"011001100",
    14611=>"000000100",
    14612=>"101001000",
    14613=>"000000100",
    14614=>"001010010",
    14615=>"110111101",
    14616=>"000000000",
    14617=>"000000000",
    14618=>"001000000",
    14619=>"111100000",
    14620=>"011110001",
    14621=>"000000000",
    14622=>"111111110",
    14623=>"111011000",
    14624=>"011110000",
    14625=>"001000100",
    14626=>"001011111",
    14627=>"011000101",
    14628=>"111111111",
    14629=>"110111011",
    14630=>"110111111",
    14631=>"000100110",
    14632=>"011000100",
    14633=>"000001000",
    14634=>"000000000",
    14635=>"000100000",
    14636=>"110111111",
    14637=>"010000110",
    14638=>"100100000",
    14639=>"110111010",
    14640=>"111110111",
    14641=>"000111011",
    14642=>"111101110",
    14643=>"000000000",
    14644=>"111111110",
    14645=>"111000000",
    14646=>"111001001",
    14647=>"001001100",
    14648=>"011000000",
    14649=>"110011100",
    14650=>"000100010",
    14651=>"001000101",
    14652=>"101000100",
    14653=>"000000000",
    14654=>"000001101",
    14655=>"010010011",
    14656=>"110010000",
    14657=>"000100100",
    14658=>"111011000",
    14659=>"011000010",
    14660=>"111111111",
    14661=>"000000100",
    14662=>"010100001",
    14663=>"001000000",
    14664=>"000000000",
    14665=>"100110110",
    14666=>"111111111",
    14667=>"001001111",
    14668=>"000000000",
    14669=>"101110111",
    14670=>"111011011",
    14671=>"000100000",
    14672=>"000011000",
    14673=>"000000000",
    14674=>"000000000",
    14675=>"110110111",
    14676=>"111111111",
    14677=>"000010000",
    14678=>"110100100",
    14679=>"110101100",
    14680=>"111110110",
    14681=>"000000111",
    14682=>"000000000",
    14683=>"000000000",
    14684=>"000000000",
    14685=>"111111011",
    14686=>"011111111",
    14687=>"001100000",
    14688=>"100100111",
    14689=>"101000101",
    14690=>"101111011",
    14691=>"010011000",
    14692=>"100110111",
    14693=>"001000100",
    14694=>"111100111",
    14695=>"111110001",
    14696=>"000000000",
    14697=>"001000000",
    14698=>"000000100",
    14699=>"001011011",
    14700=>"000000000",
    14701=>"010011001",
    14702=>"100111011",
    14703=>"011111111",
    14704=>"110011001",
    14705=>"001101011",
    14706=>"101100100",
    14707=>"110110001",
    14708=>"111111011",
    14709=>"001001000",
    14710=>"000001001",
    14711=>"000000000",
    14712=>"111111111",
    14713=>"001000000",
    14714=>"110111000",
    14715=>"110110000",
    14716=>"011001100",
    14717=>"111111000",
    14718=>"001000000",
    14719=>"000000001",
    14720=>"111111111",
    14721=>"100111111",
    14722=>"001000000",
    14723=>"101000111",
    14724=>"001111100",
    14725=>"111111111",
    14726=>"000111001",
    14727=>"011000000",
    14728=>"101100000",
    14729=>"111111111",
    14730=>"100000001",
    14731=>"011101011",
    14732=>"111011111",
    14733=>"000100110",
    14734=>"110010000",
    14735=>"110000011",
    14736=>"000000100",
    14737=>"101000000",
    14738=>"001000101",
    14739=>"100011000",
    14740=>"111000000",
    14741=>"111111011",
    14742=>"101000110",
    14743=>"111101100",
    14744=>"100001011",
    14745=>"100001010",
    14746=>"001000000",
    14747=>"100000011",
    14748=>"011111111",
    14749=>"100101110",
    14750=>"001111111",
    14751=>"010010100",
    14752=>"111000000",
    14753=>"000000000",
    14754=>"011100100",
    14755=>"000001000",
    14756=>"011111111",
    14757=>"000000010",
    14758=>"000000100",
    14759=>"000000101",
    14760=>"001000010",
    14761=>"000001100",
    14762=>"000000000",
    14763=>"001001001",
    14764=>"001000000",
    14765=>"111000101",
    14766=>"110110111",
    14767=>"111111111",
    14768=>"000000000",
    14769=>"001010101",
    14770=>"000000000",
    14771=>"000111111",
    14772=>"001101100",
    14773=>"000000110",
    14774=>"001000101",
    14775=>"000110010",
    14776=>"001111111",
    14777=>"010000000",
    14778=>"011111111",
    14779=>"011001111",
    14780=>"010001101",
    14781=>"100011111",
    14782=>"111001110",
    14783=>"110010110",
    14784=>"111000111",
    14785=>"000010000",
    14786=>"010000101",
    14787=>"111001111",
    14788=>"111110111",
    14789=>"000011111",
    14790=>"100101001",
    14791=>"001000010",
    14792=>"000000001",
    14793=>"010111111",
    14794=>"010000000",
    14795=>"101000001",
    14796=>"111010000",
    14797=>"010001100",
    14798=>"010111001",
    14799=>"001000000",
    14800=>"010000000",
    14801=>"100000000",
    14802=>"010010010",
    14803=>"111111111",
    14804=>"000100100",
    14805=>"000010011",
    14806=>"000000000",
    14807=>"110111010",
    14808=>"111101001",
    14809=>"111011111",
    14810=>"000001000",
    14811=>"111000000",
    14812=>"100101001",
    14813=>"011110100",
    14814=>"000000000",
    14815=>"100111101",
    14816=>"000001101",
    14817=>"000000101",
    14818=>"000000001",
    14819=>"001000000",
    14820=>"010010010",
    14821=>"111000001",
    14822=>"001000100",
    14823=>"111010000",
    14824=>"001001111",
    14825=>"101000000",
    14826=>"110101000",
    14827=>"111111010",
    14828=>"001001001",
    14829=>"100000001",
    14830=>"111111110",
    14831=>"101111001",
    14832=>"110000000",
    14833=>"011000110",
    14834=>"000000000",
    14835=>"001000001",
    14836=>"011010110",
    14837=>"001000010",
    14838=>"111111011",
    14839=>"000100000",
    14840=>"010000000",
    14841=>"110010010",
    14842=>"101100111",
    14843=>"000000000",
    14844=>"000000000",
    14845=>"101111111",
    14846=>"110111101",
    14847=>"110101001",
    14848=>"111111111",
    14849=>"010110000",
    14850=>"111000000",
    14851=>"000011001",
    14852=>"010101101",
    14853=>"110100101",
    14854=>"111101111",
    14855=>"000000101",
    14856=>"011011011",
    14857=>"111010101",
    14858=>"111111111",
    14859=>"010100011",
    14860=>"010110111",
    14861=>"110100010",
    14862=>"000001011",
    14863=>"010011000",
    14864=>"000111011",
    14865=>"000000111",
    14866=>"111000000",
    14867=>"010000001",
    14868=>"000000011",
    14869=>"100010100",
    14870=>"000111001",
    14871=>"000000110",
    14872=>"100110101",
    14873=>"110000110",
    14874=>"010000100",
    14875=>"000100111",
    14876=>"111111000",
    14877=>"111111101",
    14878=>"011111111",
    14879=>"000010000",
    14880=>"000010000",
    14881=>"000010001",
    14882=>"011000100",
    14883=>"000000110",
    14884=>"101111110",
    14885=>"000000000",
    14886=>"011100010",
    14887=>"110100100",
    14888=>"111111111",
    14889=>"111001000",
    14890=>"011111111",
    14891=>"000001011",
    14892=>"000000000",
    14893=>"111111011",
    14894=>"000000110",
    14895=>"110000000",
    14896=>"000000010",
    14897=>"111000000",
    14898=>"000000100",
    14899=>"011001111",
    14900=>"111101111",
    14901=>"100100001",
    14902=>"111010000",
    14903=>"111001010",
    14904=>"011111110",
    14905=>"000010110",
    14906=>"100110110",
    14907=>"111010001",
    14908=>"111000000",
    14909=>"100000000",
    14910=>"000100101",
    14911=>"000011111",
    14912=>"101111111",
    14913=>"110100000",
    14914=>"111011000",
    14915=>"000000000",
    14916=>"011111111",
    14917=>"100100111",
    14918=>"000000001",
    14919=>"011110101",
    14920=>"001011110",
    14921=>"100111000",
    14922=>"000000000",
    14923=>"111111001",
    14924=>"101001000",
    14925=>"000111111",
    14926=>"100001110",
    14927=>"111101000",
    14928=>"000000000",
    14929=>"000000000",
    14930=>"000000111",
    14931=>"111001101",
    14932=>"001001011",
    14933=>"101101011",
    14934=>"000010111",
    14935=>"011111101",
    14936=>"100000000",
    14937=>"000001111",
    14938=>"001110011",
    14939=>"000000000",
    14940=>"000111111",
    14941=>"010000000",
    14942=>"111100000",
    14943=>"010110101",
    14944=>"000000100",
    14945=>"011000111",
    14946=>"101000000",
    14947=>"011011000",
    14948=>"000111111",
    14949=>"000000000",
    14950=>"110000000",
    14951=>"110000000",
    14952=>"011011010",
    14953=>"010000101",
    14954=>"010001111",
    14955=>"110011111",
    14956=>"000110010",
    14957=>"010000000",
    14958=>"000000000",
    14959=>"010110110",
    14960=>"111111001",
    14961=>"111100000",
    14962=>"101111110",
    14963=>"010001101",
    14964=>"111110000",
    14965=>"000000100",
    14966=>"100000010",
    14967=>"000010011",
    14968=>"111111111",
    14969=>"000000000",
    14970=>"110101000",
    14971=>"000010110",
    14972=>"111111110",
    14973=>"100010111",
    14974=>"000000000",
    14975=>"011000010",
    14976=>"100011101",
    14977=>"111000010",
    14978=>"000010010",
    14979=>"110011001",
    14980=>"001001001",
    14981=>"101110110",
    14982=>"111111111",
    14983=>"111101101",
    14984=>"111111111",
    14985=>"111110100",
    14986=>"111001000",
    14987=>"111001001",
    14988=>"000000001",
    14989=>"000000000",
    14990=>"010101001",
    14991=>"000010010",
    14992=>"100100101",
    14993=>"001000100",
    14994=>"001101001",
    14995=>"110000001",
    14996=>"111111111",
    14997=>"111011000",
    14998=>"101000111",
    14999=>"110110100",
    15000=>"100001001",
    15001=>"110100100",
    15002=>"000001101",
    15003=>"001001111",
    15004=>"110111111",
    15005=>"100111001",
    15006=>"001001000",
    15007=>"010011111",
    15008=>"111000111",
    15009=>"000100100",
    15010=>"011001011",
    15011=>"101101101",
    15012=>"111111011",
    15013=>"001101100",
    15014=>"111111111",
    15015=>"000111111",
    15016=>"111000000",
    15017=>"110100000",
    15018=>"100000101",
    15019=>"111101001",
    15020=>"011001000",
    15021=>"111111111",
    15022=>"111110111",
    15023=>"011011010",
    15024=>"111111111",
    15025=>"001010000",
    15026=>"000000110",
    15027=>"001011111",
    15028=>"001101000",
    15029=>"000000000",
    15030=>"101111111",
    15031=>"111110110",
    15032=>"100100000",
    15033=>"110000000",
    15034=>"111011011",
    15035=>"100110111",
    15036=>"110111000",
    15037=>"111111111",
    15038=>"100110110",
    15039=>"111100000",
    15040=>"011111000",
    15041=>"111110101",
    15042=>"111101000",
    15043=>"010010001",
    15044=>"101100101",
    15045=>"000111111",
    15046=>"000010000",
    15047=>"111000000",
    15048=>"101101101",
    15049=>"000000111",
    15050=>"111001100",
    15051=>"110111101",
    15052=>"111111111",
    15053=>"000010010",
    15054=>"111111111",
    15055=>"000110111",
    15056=>"100101111",
    15057=>"110101111",
    15058=>"000000000",
    15059=>"011011011",
    15060=>"100111111",
    15061=>"111111111",
    15062=>"000011111",
    15063=>"111111110",
    15064=>"011001001",
    15065=>"111111101",
    15066=>"000001001",
    15067=>"010000101",
    15068=>"100100001",
    15069=>"001011001",
    15070=>"001000001",
    15071=>"100000000",
    15072=>"111110111",
    15073=>"111111111",
    15074=>"010111110",
    15075=>"100010111",
    15076=>"010001000",
    15077=>"011000101",
    15078=>"011101101",
    15079=>"111111101",
    15080=>"100100110",
    15081=>"111110000",
    15082=>"110101001",
    15083=>"010110000",
    15084=>"111111000",
    15085=>"000011000",
    15086=>"011000000",
    15087=>"000001001",
    15088=>"010111000",
    15089=>"010000010",
    15090=>"011101110",
    15091=>"110001001",
    15092=>"000010000",
    15093=>"111101111",
    15094=>"000000100",
    15095=>"100001001",
    15096=>"111011000",
    15097=>"111000100",
    15098=>"110000000",
    15099=>"000101001",
    15100=>"000100100",
    15101=>"111100000",
    15102=>"110010000",
    15103=>"000010000",
    15104=>"000000000",
    15105=>"111010000",
    15106=>"111111010",
    15107=>"111000000",
    15108=>"011000000",
    15109=>"111010000",
    15110=>"101000000",
    15111=>"000001101",
    15112=>"000010000",
    15113=>"010000000",
    15114=>"001101011",
    15115=>"000000000",
    15116=>"010011101",
    15117=>"111111010",
    15118=>"111111001",
    15119=>"111011001",
    15120=>"000110011",
    15121=>"010111100",
    15122=>"001101111",
    15123=>"000000000",
    15124=>"111010000",
    15125=>"001000000",
    15126=>"111000000",
    15127=>"010000111",
    15128=>"000101110",
    15129=>"100000100",
    15130=>"011100000",
    15131=>"111111101",
    15132=>"010000110",
    15133=>"111110001",
    15134=>"001100110",
    15135=>"000100111",
    15136=>"010000111",
    15137=>"000000000",
    15138=>"001100000",
    15139=>"000011110",
    15140=>"001000100",
    15141=>"111000001",
    15142=>"011111111",
    15143=>"111000000",
    15144=>"000000000",
    15145=>"000011111",
    15146=>"100100101",
    15147=>"100100100",
    15148=>"000110100",
    15149=>"111111110",
    15150=>"000000111",
    15151=>"111111111",
    15152=>"000000111",
    15153=>"111111111",
    15154=>"000100111",
    15155=>"100000011",
    15156=>"011111100",
    15157=>"001000000",
    15158=>"100100000",
    15159=>"101101000",
    15160=>"101000000",
    15161=>"011000011",
    15162=>"111000000",
    15163=>"101000111",
    15164=>"000000110",
    15165=>"011111110",
    15166=>"011011111",
    15167=>"010000100",
    15168=>"100111110",
    15169=>"000111110",
    15170=>"000110101",
    15171=>"010011000",
    15172=>"000001001",
    15173=>"111011111",
    15174=>"111000000",
    15175=>"000010011",
    15176=>"001011010",
    15177=>"111000000",
    15178=>"000000111",
    15179=>"111110111",
    15180=>"000000111",
    15181=>"001111111",
    15182=>"000010110",
    15183=>"011011000",
    15184=>"011000010",
    15185=>"100011001",
    15186=>"000100110",
    15187=>"111111100",
    15188=>"111110000",
    15189=>"111011000",
    15190=>"001101010",
    15191=>"111011000",
    15192=>"100110111",
    15193=>"010000000",
    15194=>"100101101",
    15195=>"111111000",
    15196=>"000011111",
    15197=>"000100110",
    15198=>"110011000",
    15199=>"000011010",
    15200=>"101111000",
    15201=>"001010000",
    15202=>"110111010",
    15203=>"111000000",
    15204=>"110111111",
    15205=>"111111000",
    15206=>"111110100",
    15207=>"000101111",
    15208=>"111000000",
    15209=>"001000001",
    15210=>"100001011",
    15211=>"010010111",
    15212=>"001111111",
    15213=>"001000000",
    15214=>"111011000",
    15215=>"111111000",
    15216=>"000100111",
    15217=>"000101101",
    15218=>"101000000",
    15219=>"111111000",
    15220=>"111001001",
    15221=>"111000000",
    15222=>"000000010",
    15223=>"000000111",
    15224=>"000000101",
    15225=>"000000111",
    15226=>"111011000",
    15227=>"000111111",
    15228=>"101101101",
    15229=>"000111111",
    15230=>"111011000",
    15231=>"000001111",
    15232=>"111000010",
    15233=>"000000000",
    15234=>"111000000",
    15235=>"111111111",
    15236=>"001011101",
    15237=>"111110010",
    15238=>"111010011",
    15239=>"000100010",
    15240=>"011011111",
    15241=>"111111110",
    15242=>"000000101",
    15243=>"000000000",
    15244=>"000000000",
    15245=>"010010000",
    15246=>"101011011",
    15247=>"000000010",
    15248=>"011001000",
    15249=>"111111010",
    15250=>"101100111",
    15251=>"000001101",
    15252=>"000001001",
    15253=>"101000000",
    15254=>"101100111",
    15255=>"111010010",
    15256=>"000000001",
    15257=>"000000000",
    15258=>"000000000",
    15259=>"100100010",
    15260=>"110110110",
    15261=>"000001010",
    15262=>"111011110",
    15263=>"110110110",
    15264=>"000000000",
    15265=>"000011011",
    15266=>"000000000",
    15267=>"100101111",
    15268=>"011111111",
    15269=>"000111111",
    15270=>"000111111",
    15271=>"000101111",
    15272=>"001000000",
    15273=>"000011111",
    15274=>"000000000",
    15275=>"000000001",
    15276=>"000100110",
    15277=>"010111111",
    15278=>"110000010",
    15279=>"111101111",
    15280=>"111010101",
    15281=>"000111110",
    15282=>"100000000",
    15283=>"011000111",
    15284=>"110101101",
    15285=>"000010000",
    15286=>"111100101",
    15287=>"000000000",
    15288=>"000000000",
    15289=>"101011010",
    15290=>"101010011",
    15291=>"000000100",
    15292=>"000110000",
    15293=>"000111010",
    15294=>"000001011",
    15295=>"000011111",
    15296=>"000000001",
    15297=>"001000000",
    15298=>"101101111",
    15299=>"000000010",
    15300=>"010111010",
    15301=>"001011111",
    15302=>"111111111",
    15303=>"000111011",
    15304=>"110110100",
    15305=>"000111111",
    15306=>"000111110",
    15307=>"000000000",
    15308=>"000111010",
    15309=>"111101011",
    15310=>"010111111",
    15311=>"111111000",
    15312=>"000000110",
    15313=>"110001110",
    15314=>"000000010",
    15315=>"111111110",
    15316=>"100100111",
    15317=>"000000110",
    15318=>"000000011",
    15319=>"111111111",
    15320=>"000100101",
    15321=>"101111111",
    15322=>"000000000",
    15323=>"101101000",
    15324=>"100100001",
    15325=>"011011011",
    15326=>"000000001",
    15327=>"000000000",
    15328=>"100100100",
    15329=>"100100000",
    15330=>"111100000",
    15331=>"000111100",
    15332=>"000000000",
    15333=>"000010110",
    15334=>"000000001",
    15335=>"010010000",
    15336=>"000010000",
    15337=>"000000000",
    15338=>"100101101",
    15339=>"101001111",
    15340=>"111000000",
    15341=>"001110000",
    15342=>"111111010",
    15343=>"001111110",
    15344=>"111111000",
    15345=>"000100110",
    15346=>"000100001",
    15347=>"000111111",
    15348=>"001101111",
    15349=>"000000111",
    15350=>"000000000",
    15351=>"101000001",
    15352=>"010000110",
    15353=>"110000000",
    15354=>"000010110",
    15355=>"100000000",
    15356=>"000000100",
    15357=>"000101011",
    15358=>"000000000",
    15359=>"000100111",
    15360=>"111000010",
    15361=>"010011010",
    15362=>"110111110",
    15363=>"100101000",
    15364=>"001001101",
    15365=>"001000111",
    15366=>"010000100",
    15367=>"101101100",
    15368=>"001000000",
    15369=>"000011010",
    15370=>"000101111",
    15371=>"001111111",
    15372=>"000110000",
    15373=>"110110000",
    15374=>"000000001",
    15375=>"100100100",
    15376=>"011010000",
    15377=>"001001100",
    15378=>"000000000",
    15379=>"000001101",
    15380=>"110000010",
    15381=>"000000000",
    15382=>"000000101",
    15383=>"100111111",
    15384=>"000000001",
    15385=>"000111111",
    15386=>"010110110",
    15387=>"011000000",
    15388=>"100010010",
    15389=>"001000000",
    15390=>"111101101",
    15391=>"110111111",
    15392=>"111111010",
    15393=>"000111011",
    15394=>"011111111",
    15395=>"000000100",
    15396=>"101100010",
    15397=>"100100000",
    15398=>"111111010",
    15399=>"001000011",
    15400=>"101101101",
    15401=>"101001111",
    15402=>"110010000",
    15403=>"001000001",
    15404=>"111101101",
    15405=>"101101111",
    15406=>"000000110",
    15407=>"110111111",
    15408=>"000000000",
    15409=>"110011010",
    15410=>"111110110",
    15411=>"001000101",
    15412=>"111111010",
    15413=>"111111111",
    15414=>"100110100",
    15415=>"000000000",
    15416=>"100000000",
    15417=>"111101111",
    15418=>"001001111",
    15419=>"000110111",
    15420=>"000111111",
    15421=>"100000000",
    15422=>"100110001",
    15423=>"010011001",
    15424=>"000000111",
    15425=>"101111010",
    15426=>"111111110",
    15427=>"000000101",
    15428=>"101001101",
    15429=>"101000100",
    15430=>"111110010",
    15431=>"111101101",
    15432=>"000010000",
    15433=>"110010010",
    15434=>"101101111",
    15435=>"101000001",
    15436=>"111111111",
    15437=>"001000111",
    15438=>"000101110",
    15439=>"010011010",
    15440=>"111101000",
    15441=>"100000111",
    15442=>"111001001",
    15443=>"111111111",
    15444=>"101100001",
    15445=>"100000000",
    15446=>"000100001",
    15447=>"111001011",
    15448=>"000000100",
    15449=>"100100101",
    15450=>"000110100",
    15451=>"000110110",
    15452=>"000000100",
    15453=>"000000000",
    15454=>"111111011",
    15455=>"011101000",
    15456=>"001000000",
    15457=>"101100101",
    15458=>"010111111",
    15459=>"010101111",
    15460=>"010101111",
    15461=>"011011000",
    15462=>"001000100",
    15463=>"100101101",
    15464=>"110110010",
    15465=>"110110110",
    15466=>"000000101",
    15467=>"111001000",
    15468=>"111000011",
    15469=>"000001010",
    15470=>"110010000",
    15471=>"000000000",
    15472=>"101001101",
    15473=>"111111111",
    15474=>"001011011",
    15475=>"010111010",
    15476=>"111111111",
    15477=>"000000000",
    15478=>"001101001",
    15479=>"111111011",
    15480=>"001101101",
    15481=>"010101111",
    15482=>"010110001",
    15483=>"111101101",
    15484=>"000011010",
    15485=>"000100110",
    15486=>"000000100",
    15487=>"011111110",
    15488=>"001011111",
    15489=>"111011000",
    15490=>"000111111",
    15491=>"101010001",
    15492=>"001000111",
    15493=>"111001101",
    15494=>"010010111",
    15495=>"111101000",
    15496=>"110111101",
    15497=>"011001100",
    15498=>"000100010",
    15499=>"010001001",
    15500=>"111001000",
    15501=>"111010000",
    15502=>"110110000",
    15503=>"000110111",
    15504=>"111001000",
    15505=>"000100111",
    15506=>"001011111",
    15507=>"011001101",
    15508=>"000010111",
    15509=>"111000000",
    15510=>"111101000",
    15511=>"000000111",
    15512=>"000001111",
    15513=>"010100100",
    15514=>"111000101",
    15515=>"011101001",
    15516=>"000111010",
    15517=>"000000010",
    15518=>"001000001",
    15519=>"100110111",
    15520=>"111010111",
    15521=>"111111110",
    15522=>"111101101",
    15523=>"000000110",
    15524=>"000111111",
    15525=>"110110001",
    15526=>"111000000",
    15527=>"001001010",
    15528=>"110011101",
    15529=>"110000110",
    15530=>"111110000",
    15531=>"000101111",
    15532=>"000011111",
    15533=>"000001111",
    15534=>"000000000",
    15535=>"000111111",
    15536=>"110000000",
    15537=>"100000000",
    15538=>"010010000",
    15539=>"000000110",
    15540=>"111000000",
    15541=>"110000000",
    15542=>"111000000",
    15543=>"111111000",
    15544=>"000000110",
    15545=>"111111111",
    15546=>"011110011",
    15547=>"110010000",
    15548=>"111000000",
    15549=>"011111111",
    15550=>"111110100",
    15551=>"111101000",
    15552=>"001101000",
    15553=>"000000000",
    15554=>"010000010",
    15555=>"110011111",
    15556=>"100111111",
    15557=>"000011110",
    15558=>"111111110",
    15559=>"000000001",
    15560=>"111000000",
    15561=>"111010000",
    15562=>"000000010",
    15563=>"111001000",
    15564=>"000010010",
    15565=>"000010111",
    15566=>"000110110",
    15567=>"101000111",
    15568=>"100000110",
    15569=>"010000000",
    15570=>"111010000",
    15571=>"010000000",
    15572=>"000111111",
    15573=>"111000000",
    15574=>"111010000",
    15575=>"000100000",
    15576=>"011110011",
    15577=>"011101111",
    15578=>"111011001",
    15579=>"000111110",
    15580=>"000110110",
    15581=>"001000011",
    15582=>"011001101",
    15583=>"111111110",
    15584=>"111101100",
    15585=>"000010000",
    15586=>"000110111",
    15587=>"000010110",
    15588=>"000000001",
    15589=>"011001000",
    15590=>"001000000",
    15591=>"001111111",
    15592=>"011000000",
    15593=>"100100100",
    15594=>"100011111",
    15595=>"010000000",
    15596=>"000111111",
    15597=>"111001000",
    15598=>"110000001",
    15599=>"111001100",
    15600=>"000110111",
    15601=>"000110110",
    15602=>"111101101",
    15603=>"111000000",
    15604=>"101000000",
    15605=>"101001101",
    15606=>"000001000",
    15607=>"000001000",
    15608=>"001010111",
    15609=>"000000000",
    15610=>"110001101",
    15611=>"111001000",
    15612=>"101111100",
    15613=>"110111101",
    15614=>"010000111",
    15615=>"011111111",
    15616=>"000000111",
    15617=>"000000010",
    15618=>"111010101",
    15619=>"010000000",
    15620=>"001001111",
    15621=>"111011000",
    15622=>"111111000",
    15623=>"000000111",
    15624=>"111001100",
    15625=>"010000000",
    15626=>"110100111",
    15627=>"001000100",
    15628=>"000101010",
    15629=>"111111010",
    15630=>"100101111",
    15631=>"100011111",
    15632=>"110110010",
    15633=>"100100000",
    15634=>"110110111",
    15635=>"110100011",
    15636=>"111000000",
    15637=>"000100111",
    15638=>"000100100",
    15639=>"000111111",
    15640=>"011111110",
    15641=>"100000100",
    15642=>"100100100",
    15643=>"101111100",
    15644=>"111001000",
    15645=>"101001111",
    15646=>"101101111",
    15647=>"011011111",
    15648=>"011101000",
    15649=>"000100000",
    15650=>"100000001",
    15651=>"111000001",
    15652=>"011000011",
    15653=>"110010000",
    15654=>"000000000",
    15655=>"111000101",
    15656=>"010111111",
    15657=>"100000000",
    15658=>"000101111",
    15659=>"111111011",
    15660=>"011011001",
    15661=>"000100101",
    15662=>"000000000",
    15663=>"100100111",
    15664=>"000111110",
    15665=>"000000111",
    15666=>"000110110",
    15667=>"000001111",
    15668=>"100100111",
    15669=>"110111010",
    15670=>"111011000",
    15671=>"011111000",
    15672=>"111010101",
    15673=>"111000111",
    15674=>"000000000",
    15675=>"101101110",
    15676=>"000000111",
    15677=>"000000111",
    15678=>"110110000",
    15679=>"011010000",
    15680=>"110010000",
    15681=>"010000000",
    15682=>"000111111",
    15683=>"111101010",
    15684=>"111111011",
    15685=>"000000111",
    15686=>"000010000",
    15687=>"000000000",
    15688=>"000011000",
    15689=>"111000000",
    15690=>"001100110",
    15691=>"000100111",
    15692=>"010000010",
    15693=>"111111000",
    15694=>"001001011",
    15695=>"100000101",
    15696=>"010101111",
    15697=>"100000001",
    15698=>"000100111",
    15699=>"001111000",
    15700=>"100110011",
    15701=>"000101000",
    15702=>"000111111",
    15703=>"101000101",
    15704=>"001001000",
    15705=>"000000000",
    15706=>"001101001",
    15707=>"000000000",
    15708=>"101011110",
    15709=>"001000010",
    15710=>"011111111",
    15711=>"000000111",
    15712=>"101100001",
    15713=>"001111110",
    15714=>"111011101",
    15715=>"011011000",
    15716=>"001111111",
    15717=>"000101111",
    15718=>"100100100",
    15719=>"000000101",
    15720=>"100011110",
    15721=>"100000000",
    15722=>"110001011",
    15723=>"000000000",
    15724=>"000010000",
    15725=>"101101110",
    15726=>"110111000",
    15727=>"101110110",
    15728=>"011000001",
    15729=>"111000110",
    15730=>"111101100",
    15731=>"111000001",
    15732=>"111111111",
    15733=>"000110000",
    15734=>"000111111",
    15735=>"010011111",
    15736=>"001111111",
    15737=>"010000111",
    15738=>"000111011",
    15739=>"000010000",
    15740=>"110011111",
    15741=>"111000000",
    15742=>"000000111",
    15743=>"111101101",
    15744=>"111111111",
    15745=>"001101101",
    15746=>"000001000",
    15747=>"100111111",
    15748=>"110011111",
    15749=>"000100000",
    15750=>"000011110",
    15751=>"101101111",
    15752=>"000000100",
    15753=>"011001011",
    15754=>"110011010",
    15755=>"110110111",
    15756=>"000000000",
    15757=>"111111100",
    15758=>"001001111",
    15759=>"001101100",
    15760=>"111100100",
    15761=>"101101111",
    15762=>"110110111",
    15763=>"001000110",
    15764=>"011011110",
    15765=>"001001000",
    15766=>"000000000",
    15767=>"001101111",
    15768=>"111110111",
    15769=>"000001010",
    15770=>"110110111",
    15771=>"110000000",
    15772=>"000111001",
    15773=>"010011110",
    15774=>"111011011",
    15775=>"111111001",
    15776=>"000000000",
    15777=>"001011011",
    15778=>"001010010",
    15779=>"100110000",
    15780=>"000000100",
    15781=>"110111110",
    15782=>"101000001",
    15783=>"010000000",
    15784=>"111111101",
    15785=>"111110100",
    15786=>"000000001",
    15787=>"010010110",
    15788=>"010010011",
    15789=>"001000000",
    15790=>"001000110",
    15791=>"000101111",
    15792=>"110101111",
    15793=>"101101101",
    15794=>"010000010",
    15795=>"110110110",
    15796=>"110110000",
    15797=>"000100110",
    15798=>"000001110",
    15799=>"000100000",
    15800=>"001100000",
    15801=>"010010000",
    15802=>"110100111",
    15803=>"000000100",
    15804=>"101101000",
    15805=>"000010010",
    15806=>"111000001",
    15807=>"010011000",
    15808=>"011010000",
    15809=>"001000000",
    15810=>"110110010",
    15811=>"000000000",
    15812=>"010010000",
    15813=>"011111011",
    15814=>"000110110",
    15815=>"110101100",
    15816=>"110000001",
    15817=>"010010000",
    15818=>"000011000",
    15819=>"101000100",
    15820=>"010011101",
    15821=>"011010110",
    15822=>"001011000",
    15823=>"111101100",
    15824=>"111111000",
    15825=>"000000000",
    15826=>"000000100",
    15827=>"100011011",
    15828=>"110110110",
    15829=>"001001111",
    15830=>"000100010",
    15831=>"001000001",
    15832=>"110011011",
    15833=>"101101001",
    15834=>"101000110",
    15835=>"001111010",
    15836=>"010010011",
    15837=>"100101101",
    15838=>"000000100",
    15839=>"110010110",
    15840=>"001110010",
    15841=>"011011011",
    15842=>"100101001",
    15843=>"010010010",
    15844=>"001001001",
    15845=>"000000001",
    15846=>"000000000",
    15847=>"010000000",
    15848=>"001000000",
    15849=>"001001001",
    15850=>"010010110",
    15851=>"111111000",
    15852=>"010010110",
    15853=>"011101001",
    15854=>"111111111",
    15855=>"110110111",
    15856=>"010110110",
    15857=>"101111011",
    15858=>"100000000",
    15859=>"010010110",
    15860=>"101101111",
    15861=>"000000000",
    15862=>"001001000",
    15863=>"111110100",
    15864=>"110110000",
    15865=>"000101001",
    15866=>"100000000",
    15867=>"101101001",
    15868=>"001001001",
    15869=>"111111111",
    15870=>"011111010",
    15871=>"111110111",
    15872=>"111111110",
    15873=>"110100100",
    15874=>"000011001",
    15875=>"001101110",
    15876=>"111110110",
    15877=>"000111110",
    15878=>"111000000",
    15879=>"000001101",
    15880=>"100100100",
    15881=>"110110110",
    15882=>"001100110",
    15883=>"001000001",
    15884=>"001111011",
    15885=>"100110011",
    15886=>"101000100",
    15887=>"000001100",
    15888=>"000011011",
    15889=>"100101100",
    15890=>"110111011",
    15891=>"001000000",
    15892=>"011000000",
    15893=>"010100000",
    15894=>"000000000",
    15895=>"101011110",
    15896=>"100110000",
    15897=>"111100100",
    15898=>"100100010",
    15899=>"001001011",
    15900=>"111101101",
    15901=>"110110000",
    15902=>"111110011",
    15903=>"000000000",
    15904=>"010110111",
    15905=>"000000000",
    15906=>"111110110",
    15907=>"000010001",
    15908=>"000001100",
    15909=>"100110110",
    15910=>"011011011",
    15911=>"111111010",
    15912=>"111111011",
    15913=>"001001011",
    15914=>"000000000",
    15915=>"100111000",
    15916=>"110111011",
    15917=>"011110011",
    15918=>"000000111",
    15919=>"110111011",
    15920=>"000000001",
    15921=>"010101110",
    15922=>"001111111",
    15923=>"011011100",
    15924=>"100110110",
    15925=>"000000011",
    15926=>"000001011",
    15927=>"010011000",
    15928=>"011000000",
    15929=>"001000010",
    15930=>"000000000",
    15931=>"011001101",
    15932=>"101001100",
    15933=>"001000100",
    15934=>"100111111",
    15935=>"001011011",
    15936=>"110110000",
    15937=>"001001000",
    15938=>"011000011",
    15939=>"011001100",
    15940=>"101111011",
    15941=>"000011110",
    15942=>"111100010",
    15943=>"111001101",
    15944=>"000000100",
    15945=>"110000000",
    15946=>"010110111",
    15947=>"100100000",
    15948=>"001011100",
    15949=>"100100011",
    15950=>"101001001",
    15951=>"011001000",
    15952=>"011011100",
    15953=>"011001100",
    15954=>"101000010",
    15955=>"100110110",
    15956=>"010010000",
    15957=>"011001101",
    15958=>"011110010",
    15959=>"110101100",
    15960=>"111110011",
    15961=>"001000000",
    15962=>"000001001",
    15963=>"001011100",
    15964=>"100100000",
    15965=>"011110011",
    15966=>"111000000",
    15967=>"010101100",
    15968=>"110010001",
    15969=>"101001001",
    15970=>"011011101",
    15971=>"111111000",
    15972=>"001000011",
    15973=>"001001000",
    15974=>"111011000",
    15975=>"001000001",
    15976=>"111111100",
    15977=>"100001110",
    15978=>"100110000",
    15979=>"001000111",
    15980=>"001001000",
    15981=>"001001100",
    15982=>"110111010",
    15983=>"111011001",
    15984=>"001111111",
    15985=>"100100000",
    15986=>"111001000",
    15987=>"000011010",
    15988=>"110100110",
    15989=>"000000000",
    15990=>"111100011",
    15991=>"011111101",
    15992=>"111110111",
    15993=>"101100000",
    15994=>"001001001",
    15995=>"000000111",
    15996=>"110110000",
    15997=>"101100001",
    15998=>"111010000",
    15999=>"000000001",
    16000=>"000001011",
    16001=>"111110100",
    16002=>"110110100",
    16003=>"111110110",
    16004=>"000001110",
    16005=>"101100011",
    16006=>"000001001",
    16007=>"111010000",
    16008=>"101011100",
    16009=>"001001111",
    16010=>"111111110",
    16011=>"000100100",
    16012=>"110100001",
    16013=>"111010100",
    16014=>"001011010",
    16015=>"111110110",
    16016=>"000000001",
    16017=>"111110010",
    16018=>"001011110",
    16019=>"101011110",
    16020=>"001001001",
    16021=>"000000110",
    16022=>"010000000",
    16023=>"000000000",
    16024=>"001001110",
    16025=>"001011111",
    16026=>"001011010",
    16027=>"000000001",
    16028=>"000110010",
    16029=>"001001010",
    16030=>"000000001",
    16031=>"011110101",
    16032=>"001001001",
    16033=>"001001000",
    16034=>"000000001",
    16035=>"001000011",
    16036=>"000001011",
    16037=>"111110011",
    16038=>"111000001",
    16039=>"101101101",
    16040=>"101011011",
    16041=>"001011110",
    16042=>"011111110",
    16043=>"001001011",
    16044=>"000001110",
    16045=>"000001011",
    16046=>"001011111",
    16047=>"110110110",
    16048=>"100001011",
    16049=>"110100000",
    16050=>"000000001",
    16051=>"110100000",
    16052=>"001011011",
    16053=>"000011111",
    16054=>"000001011",
    16055=>"011011111",
    16056=>"110111110",
    16057=>"000011100",
    16058=>"000000101",
    16059=>"111110000",
    16060=>"111111110",
    16061=>"101100000",
    16062=>"001001001",
    16063=>"000000000",
    16064=>"001001110",
    16065=>"110100000",
    16066=>"001001011",
    16067=>"110110000",
    16068=>"000001011",
    16069=>"000001001",
    16070=>"010010011",
    16071=>"100001011",
    16072=>"001001011",
    16073=>"011100010",
    16074=>"000001100",
    16075=>"000000000",
    16076=>"000010000",
    16077=>"100000110",
    16078=>"000001011",
    16079=>"110100000",
    16080=>"110100000",
    16081=>"000000000",
    16082=>"010000000",
    16083=>"100110111",
    16084=>"100100101",
    16085=>"110110110",
    16086=>"000000000",
    16087=>"000001111",
    16088=>"001001110",
    16089=>"000001111",
    16090=>"110100000",
    16091=>"110100100",
    16092=>"101001101",
    16093=>"110100100",
    16094=>"110111100",
    16095=>"111110100",
    16096=>"001001011",
    16097=>"000001001",
    16098=>"110110100",
    16099=>"100001010",
    16100=>"000001001",
    16101=>"010000000",
    16102=>"001110100",
    16103=>"001001011",
    16104=>"100100001",
    16105=>"001011110",
    16106=>"001001111",
    16107=>"100111111",
    16108=>"111110000",
    16109=>"110100010",
    16110=>"001001111",
    16111=>"101001110",
    16112=>"110110100",
    16113=>"110100001",
    16114=>"000110001",
    16115=>"000111110",
    16116=>"110110100",
    16117=>"010100100",
    16118=>"110110001",
    16119=>"000010100",
    16120=>"100001111",
    16121=>"010000101",
    16122=>"111100001",
    16123=>"011010011",
    16124=>"111101011",
    16125=>"111011110",
    16126=>"001100111",
    16127=>"001011111",
    16128=>"010000110",
    16129=>"010011000",
    16130=>"100000111",
    16131=>"011000001",
    16132=>"110011001",
    16133=>"000000000",
    16134=>"010010101",
    16135=>"101000000",
    16136=>"000100011",
    16137=>"101000000",
    16138=>"111101001",
    16139=>"000011000",
    16140=>"101010111",
    16141=>"111111111",
    16142=>"000000001",
    16143=>"000000010",
    16144=>"110110111",
    16145=>"110100000",
    16146=>"111100100",
    16147=>"011110100",
    16148=>"011111011",
    16149=>"110100000",
    16150=>"100000101",
    16151=>"111100000",
    16152=>"101001001",
    16153=>"011110101",
    16154=>"100100100",
    16155=>"000000100",
    16156=>"101001000",
    16157=>"011001101",
    16158=>"111101111",
    16159=>"111111111",
    16160=>"101101111",
    16161=>"000000000",
    16162=>"110011101",
    16163=>"110111110",
    16164=>"000001001",
    16165=>"111101101",
    16166=>"000000111",
    16167=>"000000010",
    16168=>"010000000",
    16169=>"110100000",
    16170=>"010000010",
    16171=>"000000001",
    16172=>"000101110",
    16173=>"000000000",
    16174=>"111000000",
    16175=>"111101100",
    16176=>"001111111",
    16177=>"101011010",
    16178=>"000100110",
    16179=>"111000011",
    16180=>"010110111",
    16181=>"111111101",
    16182=>"000111111",
    16183=>"011111011",
    16184=>"110110000",
    16185=>"111100011",
    16186=>"001100100",
    16187=>"111010011",
    16188=>"000000000",
    16189=>"111000001",
    16190=>"000000101",
    16191=>"010111010",
    16192=>"101000000",
    16193=>"101000111",
    16194=>"000111111",
    16195=>"000000000",
    16196=>"100001011",
    16197=>"001000001",
    16198=>"000000010",
    16199=>"011111000",
    16200=>"001011110",
    16201=>"010010010",
    16202=>"110011100",
    16203=>"100000000",
    16204=>"111000000",
    16205=>"000111000",
    16206=>"001110011",
    16207=>"000010111",
    16208=>"010010000",
    16209=>"101000000",
    16210=>"000000010",
    16211=>"110101101",
    16212=>"100000001",
    16213=>"000010010",
    16214=>"101000000",
    16215=>"001000000",
    16216=>"111001101",
    16217=>"000010110",
    16218=>"001001011",
    16219=>"000000110",
    16220=>"101100000",
    16221=>"000000000",
    16222=>"001001101",
    16223=>"100101111",
    16224=>"000011111",
    16225=>"001010110",
    16226=>"001011011",
    16227=>"011110000",
    16228=>"101001111",
    16229=>"111000000",
    16230=>"100000000",
    16231=>"011000000",
    16232=>"010011110",
    16233=>"111100000",
    16234=>"011100100",
    16235=>"111111100",
    16236=>"111000000",
    16237=>"010111000",
    16238=>"101111111",
    16239=>"100000000",
    16240=>"000010001",
    16241=>"000001110",
    16242=>"110000000",
    16243=>"010010110",
    16244=>"000111111",
    16245=>"000000000",
    16246=>"111101111",
    16247=>"000000011",
    16248=>"111011101",
    16249=>"000000101",
    16250=>"011110011",
    16251=>"000101111",
    16252=>"110000010",
    16253=>"010111000",
    16254=>"000000000",
    16255=>"111111101",
    16256=>"111111111",
    16257=>"000011000",
    16258=>"100000000",
    16259=>"101100011",
    16260=>"110100110",
    16261=>"001100010",
    16262=>"111111111",
    16263=>"000111001",
    16264=>"011001010",
    16265=>"000011011",
    16266=>"000000101",
    16267=>"000000000",
    16268=>"011010111",
    16269=>"010110010",
    16270=>"011011011",
    16271=>"011001001",
    16272=>"111111111",
    16273=>"010111010",
    16274=>"011111111",
    16275=>"000001101",
    16276=>"011010000",
    16277=>"001111011",
    16278=>"111111101",
    16279=>"000000000",
    16280=>"111101111",
    16281=>"000000000",
    16282=>"111111111",
    16283=>"000001001",
    16284=>"111111111",
    16285=>"111111111",
    16286=>"111111111",
    16287=>"000000000",
    16288=>"110000000",
    16289=>"100100100",
    16290=>"111101110",
    16291=>"111111111",
    16292=>"111111011",
    16293=>"100000001",
    16294=>"111111111",
    16295=>"101000000",
    16296=>"000000000",
    16297=>"000000001",
    16298=>"001101101",
    16299=>"111101111",
    16300=>"000000100",
    16301=>"000000000",
    16302=>"000000000",
    16303=>"000000001",
    16304=>"000000100",
    16305=>"000011000",
    16306=>"000000000",
    16307=>"011001000",
    16308=>"111111111",
    16309=>"010100111",
    16310=>"000000000",
    16311=>"111111110",
    16312=>"000000000",
    16313=>"000000000",
    16314=>"000000000",
    16315=>"010011000",
    16316=>"000000000",
    16317=>"101111011",
    16318=>"000000101",
    16319=>"010101011",
    16320=>"111100111",
    16321=>"101100000",
    16322=>"000000000",
    16323=>"011110000",
    16324=>"000000001",
    16325=>"110110111",
    16326=>"000101110",
    16327=>"000000000",
    16328=>"110111010",
    16329=>"111111111",
    16330=>"000000000",
    16331=>"111101111",
    16332=>"001101101",
    16333=>"000000000",
    16334=>"000000000",
    16335=>"010010010",
    16336=>"011111111",
    16337=>"000100000",
    16338=>"110100000",
    16339=>"111101111",
    16340=>"011011011",
    16341=>"010010010",
    16342=>"111111111",
    16343=>"101100001",
    16344=>"011011111",
    16345=>"111111111",
    16346=>"111011111",
    16347=>"010010000",
    16348=>"101111111",
    16349=>"000011011",
    16350=>"111111100",
    16351=>"000001001",
    16352=>"000100101",
    16353=>"100011111",
    16354=>"010010011",
    16355=>"000000000",
    16356=>"000000000",
    16357=>"101101100",
    16358=>"001000000",
    16359=>"000000000",
    16360=>"111111111",
    16361=>"000010000",
    16362=>"111111111",
    16363=>"000000000",
    16364=>"111010000",
    16365=>"000000000",
    16366=>"011001011",
    16367=>"111110111",
    16368=>"111111111",
    16369=>"000100000",
    16370=>"001001000",
    16371=>"101000101",
    16372=>"110010011",
    16373=>"000000000",
    16374=>"000000000",
    16375=>"000000000",
    16376=>"000000000",
    16377=>"000000000",
    16378=>"110111111",
    16379=>"010111010",
    16380=>"111110111",
    16381=>"000000000",
    16382=>"000011001",
    16383=>"111111111");
    BEGIN
    weight <= ROM_content(to_integer(address));
END RTL;