LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L9_2_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L9_2_BNROM;

ARCHITECTURE RTL OF L9_2_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 62) OF STD_LOGIC_VECTOR(15 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  (0=>"0000000010011011",
  1=>"1111111011110010",
  2=>"1111111111011010",
  3=>"0000000001101100",
  4=>"1111111101111110",
  5=>"1111111110010010",
  6=>"0000001101001000",
  7=>"0000000000010100",
  8=>"1111111101101011",
  9=>"1111111110111101",
  10=>"1111111111010001",
  11=>"1111111111110100",
  12=>"1111111111101010",
  13=>"1111111111110101",
  14=>"1111110101110100",
  15=>"1111111111010011",
  16=>"1111001100000010",
  17=>"0000000000000010",
  18=>"1111111110111101",
  19=>"1111111111011001",
  20=>"0000000001010111",
  21=>"1111111110101101",
  22=>"1111111110100001",
  23=>"0000000000111000",
  24=>"0000000000110011",
  25=>"0000000000010001",
  26=>"1111111101100001",
  27=>"0000000010110000",
  28=>"0000000001001100",
  29=>"1111111110010000",
  30=>"1111111110100100",
  31=>"0000000011111110",
  32=>"1111111111000011",
  33=>"1111111110001001",
  34=>"0000000000110101",
  35=>"0000000000010000",
  36=>"0000000000100110",
  37=>"1111111110011100",
  38=>"1111111110110100",
  39=>"1111110010100110",
  40=>"0000001001111111",
  41=>"1111001101011110",
  42=>"0000000000111010",
  43=>"0000000000101001",
  44=>"1111111101011001",
  45=>"0000000010011100",
  46=>"1111111101111101",
  47=>"1111111110101110",
  48=>"0000000000000100",
  49=>"0000000010011010",
  50=>"1111111111111100",
  51=>"1111111101111011",
  52=>"0000000001000011",
  53=>"0000000000110010",
  54=>"1111111111010000",
  55=>"1111111101000111",
  56=>"0000000101010100",
  57=>"1111111110001010",
  58=>"1111111101101011",
  59=>"0000000000111101",
  60=>"1111111111111000",
  61=>"0000000001011111",
  62=>"0000000000000000");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;